module basic_750_5000_1000_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_701,In_548);
nor U1 (N_1,In_668,In_12);
xnor U2 (N_2,In_192,In_11);
and U3 (N_3,In_529,In_107);
nor U4 (N_4,In_216,In_479);
xor U5 (N_5,In_532,In_525);
xnor U6 (N_6,In_109,In_318);
xor U7 (N_7,In_203,In_224);
nand U8 (N_8,In_636,In_475);
xnor U9 (N_9,In_616,In_162);
and U10 (N_10,In_561,In_491);
nor U11 (N_11,In_155,In_535);
or U12 (N_12,In_141,In_731);
nor U13 (N_13,In_632,In_703);
nor U14 (N_14,In_28,In_483);
nand U15 (N_15,In_380,In_176);
xnor U16 (N_16,In_56,In_426);
xor U17 (N_17,In_153,In_600);
or U18 (N_18,In_390,In_229);
nand U19 (N_19,In_283,In_424);
xnor U20 (N_20,In_193,In_39);
or U21 (N_21,In_101,In_586);
or U22 (N_22,In_628,In_106);
xor U23 (N_23,In_313,In_329);
or U24 (N_24,In_476,In_310);
nor U25 (N_25,In_412,In_667);
nand U26 (N_26,In_580,In_734);
nor U27 (N_27,In_740,In_385);
nor U28 (N_28,In_143,In_408);
nor U29 (N_29,In_414,In_705);
xnor U30 (N_30,In_625,In_123);
or U31 (N_31,In_641,In_403);
or U32 (N_32,In_607,In_376);
nor U33 (N_33,In_50,In_741);
or U34 (N_34,In_489,In_612);
nand U35 (N_35,In_320,In_236);
xnor U36 (N_36,In_443,In_265);
nand U37 (N_37,In_285,In_277);
nand U38 (N_38,In_199,In_630);
nand U39 (N_39,In_551,In_743);
nand U40 (N_40,In_344,In_558);
and U41 (N_41,In_732,In_67);
nand U42 (N_42,In_599,In_695);
or U43 (N_43,In_183,In_490);
nand U44 (N_44,In_437,In_299);
nor U45 (N_45,In_134,In_186);
xnor U46 (N_46,In_503,In_188);
or U47 (N_47,In_96,In_204);
xor U48 (N_48,In_161,In_32);
and U49 (N_49,In_677,In_685);
nor U50 (N_50,In_524,In_603);
and U51 (N_51,In_338,In_258);
xor U52 (N_52,In_650,In_635);
or U53 (N_53,In_480,In_230);
or U54 (N_54,In_547,In_418);
xor U55 (N_55,In_640,In_672);
nand U56 (N_56,In_5,In_332);
nor U57 (N_57,In_670,In_308);
or U58 (N_58,In_666,In_104);
or U59 (N_59,In_301,In_550);
nand U60 (N_60,In_737,In_3);
nor U61 (N_61,In_72,In_339);
nand U62 (N_62,In_178,In_516);
nand U63 (N_63,In_506,In_58);
nor U64 (N_64,In_202,In_191);
nand U65 (N_65,In_197,In_276);
nor U66 (N_66,In_453,In_92);
or U67 (N_67,In_127,In_281);
nand U68 (N_68,In_715,In_243);
or U69 (N_69,In_461,In_567);
and U70 (N_70,In_559,In_70);
xnor U71 (N_71,In_214,In_512);
nor U72 (N_72,In_302,In_352);
or U73 (N_73,In_664,In_268);
or U74 (N_74,In_98,In_458);
nor U75 (N_75,In_97,In_619);
and U76 (N_76,In_60,In_207);
nand U77 (N_77,In_404,In_520);
and U78 (N_78,In_564,In_704);
nor U79 (N_79,In_353,In_232);
nor U80 (N_80,In_169,In_38);
nand U81 (N_81,In_417,In_279);
xor U82 (N_82,In_24,In_263);
nor U83 (N_83,In_687,In_584);
nand U84 (N_84,In_570,In_721);
nor U85 (N_85,In_546,In_293);
and U86 (N_86,In_185,In_369);
nand U87 (N_87,In_656,In_87);
nand U88 (N_88,In_690,In_343);
and U89 (N_89,In_317,In_566);
or U90 (N_90,In_66,In_733);
xor U91 (N_91,In_723,In_306);
xor U92 (N_92,In_255,In_504);
or U93 (N_93,In_406,In_342);
nor U94 (N_94,In_45,In_307);
and U95 (N_95,In_365,In_444);
xnor U96 (N_96,In_634,In_341);
or U97 (N_97,In_719,In_442);
and U98 (N_98,In_26,In_747);
xnor U99 (N_99,In_136,In_717);
nand U100 (N_100,In_170,In_495);
xnor U101 (N_101,In_126,In_257);
or U102 (N_102,In_270,In_637);
nand U103 (N_103,In_234,In_439);
nand U104 (N_104,N_52,In_653);
xor U105 (N_105,In_448,In_595);
and U106 (N_106,N_75,In_590);
nor U107 (N_107,In_331,In_358);
and U108 (N_108,In_556,In_468);
xor U109 (N_109,In_608,In_83);
and U110 (N_110,In_118,In_43);
and U111 (N_111,In_614,In_510);
nand U112 (N_112,In_102,In_316);
nor U113 (N_113,In_691,In_288);
or U114 (N_114,In_633,In_400);
or U115 (N_115,In_583,N_60);
or U116 (N_116,N_90,In_541);
nor U117 (N_117,In_280,In_89);
nor U118 (N_118,In_182,In_706);
and U119 (N_119,In_275,In_7);
or U120 (N_120,In_484,In_722);
nand U121 (N_121,In_63,In_158);
xnor U122 (N_122,In_613,In_527);
nand U123 (N_123,In_659,In_91);
or U124 (N_124,In_488,In_111);
nor U125 (N_125,In_345,In_621);
and U126 (N_126,In_391,In_0);
and U127 (N_127,In_289,N_87);
or U128 (N_128,N_37,N_74);
xor U129 (N_129,N_32,In_330);
nor U130 (N_130,N_14,In_748);
and U131 (N_131,In_247,In_115);
or U132 (N_132,In_698,In_135);
nor U133 (N_133,In_233,In_356);
xor U134 (N_134,In_598,In_90);
xnor U135 (N_135,In_673,In_145);
nand U136 (N_136,In_166,N_76);
nor U137 (N_137,In_94,In_464);
or U138 (N_138,In_683,In_387);
and U139 (N_139,In_346,N_71);
xnor U140 (N_140,In_662,In_61);
nor U141 (N_141,In_411,In_511);
xor U142 (N_142,In_371,In_361);
nand U143 (N_143,N_2,In_381);
xor U144 (N_144,In_645,In_240);
or U145 (N_145,In_278,In_379);
and U146 (N_146,In_259,In_292);
nand U147 (N_147,N_33,N_48);
or U148 (N_148,In_62,N_93);
nor U149 (N_149,In_177,N_50);
nand U150 (N_150,In_472,In_474);
nor U151 (N_151,N_28,N_7);
nand U152 (N_152,In_73,In_206);
xnor U153 (N_153,In_565,In_602);
or U154 (N_154,In_364,In_696);
and U155 (N_155,In_648,In_42);
and U156 (N_156,In_374,In_351);
or U157 (N_157,In_618,In_322);
and U158 (N_158,In_296,In_99);
nand U159 (N_159,In_454,In_41);
nor U160 (N_160,In_187,In_700);
nand U161 (N_161,In_241,N_81);
nand U162 (N_162,N_64,In_429);
nand U163 (N_163,In_323,In_150);
or U164 (N_164,In_702,N_1);
nand U165 (N_165,In_446,In_738);
nand U166 (N_166,In_156,In_654);
nand U167 (N_167,In_425,In_457);
nand U168 (N_168,In_103,In_113);
or U169 (N_169,In_509,In_195);
or U170 (N_170,In_455,N_83);
nor U171 (N_171,In_609,In_451);
and U172 (N_172,In_16,In_534);
xnor U173 (N_173,In_321,In_264);
nor U174 (N_174,In_718,In_152);
nor U175 (N_175,In_427,In_496);
nor U176 (N_176,In_312,N_20);
or U177 (N_177,In_120,In_389);
nand U178 (N_178,In_410,In_250);
and U179 (N_179,In_742,In_368);
nor U180 (N_180,In_505,In_745);
and U181 (N_181,In_582,In_112);
and U182 (N_182,In_309,N_0);
xnor U183 (N_183,In_71,In_434);
nand U184 (N_184,In_724,In_522);
or U185 (N_185,In_746,In_646);
xor U186 (N_186,In_593,In_294);
nand U187 (N_187,In_736,In_626);
nand U188 (N_188,In_384,In_282);
and U189 (N_189,In_215,In_528);
and U190 (N_190,In_271,In_226);
and U191 (N_191,In_517,In_52);
nor U192 (N_192,In_601,In_225);
xnor U193 (N_193,In_431,In_65);
xnor U194 (N_194,In_217,In_340);
nor U195 (N_195,In_148,N_45);
and U196 (N_196,In_196,N_22);
xor U197 (N_197,In_508,N_94);
and U198 (N_198,In_712,In_560);
nand U199 (N_199,In_201,In_378);
nand U200 (N_200,In_75,In_370);
or U201 (N_201,In_487,In_69);
nor U202 (N_202,N_104,In_354);
and U203 (N_203,In_649,In_693);
or U204 (N_204,In_349,In_124);
nand U205 (N_205,In_34,In_573);
and U206 (N_206,In_68,N_195);
and U207 (N_207,N_3,In_679);
or U208 (N_208,N_107,N_150);
nand U209 (N_209,In_409,In_588);
xnor U210 (N_210,N_41,In_314);
nand U211 (N_211,In_327,In_594);
xnor U212 (N_212,N_95,N_184);
and U213 (N_213,In_382,In_692);
xor U214 (N_214,In_59,In_105);
nor U215 (N_215,N_192,N_144);
or U216 (N_216,In_671,In_304);
nor U217 (N_217,N_156,In_64);
xnor U218 (N_218,In_116,N_133);
nand U219 (N_219,In_48,N_165);
and U220 (N_220,N_55,In_235);
and U221 (N_221,N_125,In_171);
or U222 (N_222,In_147,In_184);
xnor U223 (N_223,In_518,N_84);
and U224 (N_224,In_728,In_337);
xnor U225 (N_225,N_47,N_198);
nor U226 (N_226,In_49,N_13);
xnor U227 (N_227,In_33,In_303);
xnor U228 (N_228,N_29,In_74);
or U229 (N_229,In_419,In_394);
or U230 (N_230,N_142,In_287);
or U231 (N_231,In_638,N_191);
nor U232 (N_232,In_544,In_173);
xor U233 (N_233,In_499,In_440);
xnor U234 (N_234,In_689,In_577);
nor U235 (N_235,N_62,In_441);
and U236 (N_236,In_575,In_27);
nor U237 (N_237,N_141,In_514);
xor U238 (N_238,In_8,N_91);
nor U239 (N_239,In_51,N_175);
nand U240 (N_240,In_13,N_10);
and U241 (N_241,In_328,In_413);
nand U242 (N_242,N_134,N_155);
xnor U243 (N_243,In_88,In_359);
nand U244 (N_244,N_77,In_729);
nand U245 (N_245,In_44,In_274);
xnor U246 (N_246,In_297,N_197);
and U247 (N_247,In_682,In_77);
and U248 (N_248,In_108,In_272);
nand U249 (N_249,In_80,In_167);
nand U250 (N_250,In_238,N_53);
nor U251 (N_251,In_205,N_42);
nand U252 (N_252,N_96,N_176);
xor U253 (N_253,In_622,In_357);
nor U254 (N_254,N_85,N_51);
nand U255 (N_255,In_699,In_149);
nand U256 (N_256,In_540,N_128);
and U257 (N_257,In_57,In_132);
or U258 (N_258,In_208,In_401);
and U259 (N_259,In_144,N_110);
nor U260 (N_260,In_326,In_194);
nor U261 (N_261,In_744,In_386);
and U262 (N_262,N_146,In_350);
nand U263 (N_263,In_311,N_161);
xor U264 (N_264,In_581,N_27);
nand U265 (N_265,In_174,In_139);
xnor U266 (N_266,In_200,In_131);
and U267 (N_267,In_471,In_642);
or U268 (N_268,In_53,In_663);
or U269 (N_269,N_35,In_360);
or U270 (N_270,In_397,In_17);
xor U271 (N_271,In_462,In_128);
xnor U272 (N_272,In_665,In_388);
xnor U273 (N_273,In_286,N_63);
and U274 (N_274,In_209,In_377);
and U275 (N_275,In_552,In_237);
and U276 (N_276,In_223,In_122);
xnor U277 (N_277,N_162,In_465);
or U278 (N_278,In_78,N_23);
nand U279 (N_279,N_180,In_163);
and U280 (N_280,N_159,In_450);
nor U281 (N_281,In_643,In_399);
nor U282 (N_282,In_325,In_611);
nand U283 (N_283,In_37,In_10);
nor U284 (N_284,In_709,In_597);
nand U285 (N_285,In_248,In_246);
and U286 (N_286,N_30,In_730);
or U287 (N_287,In_542,In_676);
xor U288 (N_288,In_267,N_157);
xor U289 (N_289,In_562,In_714);
nand U290 (N_290,In_231,N_66);
xor U291 (N_291,In_262,N_132);
or U292 (N_292,In_555,In_227);
xor U293 (N_293,N_189,In_298);
or U294 (N_294,In_54,In_355);
and U295 (N_295,N_108,N_173);
and U296 (N_296,N_168,In_130);
nor U297 (N_297,In_467,In_449);
nor U298 (N_298,In_261,In_735);
nor U299 (N_299,N_73,N_78);
or U300 (N_300,In_198,N_218);
nor U301 (N_301,In_578,In_416);
nand U302 (N_302,In_422,N_70);
and U303 (N_303,In_86,In_675);
xnor U304 (N_304,In_669,In_160);
or U305 (N_305,In_563,In_589);
nor U306 (N_306,In_30,N_240);
and U307 (N_307,N_265,In_658);
and U308 (N_308,In_605,N_167);
xnor U309 (N_309,In_435,In_6);
and U310 (N_310,In_222,N_235);
xor U311 (N_311,N_270,In_1);
nand U312 (N_312,In_686,N_171);
nor U313 (N_313,In_571,In_502);
and U314 (N_314,N_115,In_694);
nand U315 (N_315,N_109,N_247);
and U316 (N_316,In_291,In_610);
or U317 (N_317,N_160,In_697);
and U318 (N_318,N_206,N_181);
xnor U319 (N_319,N_231,In_300);
nand U320 (N_320,In_725,N_219);
xor U321 (N_321,In_568,In_15);
or U322 (N_322,N_224,N_82);
nand U323 (N_323,In_335,N_220);
xor U324 (N_324,In_716,N_59);
nor U325 (N_325,N_99,In_430);
or U326 (N_326,In_383,N_68);
xnor U327 (N_327,N_245,In_398);
or U328 (N_328,N_147,N_106);
xor U329 (N_329,In_459,N_130);
and U330 (N_330,N_44,In_9);
nor U331 (N_331,N_255,In_157);
or U332 (N_332,In_117,N_211);
nand U333 (N_333,N_253,N_251);
and U334 (N_334,In_604,In_657);
nor U335 (N_335,N_281,N_213);
nand U336 (N_336,In_55,In_639);
or U337 (N_337,N_223,In_168);
nand U338 (N_338,In_647,In_245);
and U339 (N_339,In_22,In_95);
nor U340 (N_340,N_241,N_89);
nand U341 (N_341,N_276,N_57);
nor U342 (N_342,In_4,N_212);
xnor U343 (N_343,N_88,In_707);
or U344 (N_344,N_120,N_216);
xnor U345 (N_345,In_2,In_129);
and U346 (N_346,N_283,N_280);
nand U347 (N_347,N_252,In_617);
or U348 (N_348,In_373,In_523);
nand U349 (N_349,In_681,N_6);
nor U350 (N_350,In_536,In_395);
nor U351 (N_351,N_153,N_228);
or U352 (N_352,N_183,N_268);
nand U353 (N_353,N_158,In_140);
nand U354 (N_354,In_84,In_624);
xor U355 (N_355,N_285,In_142);
nand U356 (N_356,N_124,N_193);
nand U357 (N_357,In_254,In_76);
or U358 (N_358,N_261,N_200);
nor U359 (N_359,N_49,In_739);
nor U360 (N_360,N_279,In_100);
or U361 (N_361,In_661,In_266);
or U362 (N_362,N_250,N_126);
nand U363 (N_363,In_498,N_293);
or U364 (N_364,N_177,N_119);
nor U365 (N_365,N_56,In_253);
and U366 (N_366,In_477,In_256);
and U367 (N_367,In_538,N_92);
xor U368 (N_368,In_500,N_246);
nor U369 (N_369,In_79,N_294);
or U370 (N_370,N_139,In_159);
nand U371 (N_371,N_272,In_501);
nor U372 (N_372,N_236,N_288);
xnor U373 (N_373,In_210,In_420);
xnor U374 (N_374,N_72,N_65);
xor U375 (N_375,N_221,N_101);
nand U376 (N_376,In_507,N_214);
and U377 (N_377,N_263,N_46);
xnor U378 (N_378,In_396,N_140);
xnor U379 (N_379,In_615,N_244);
and U380 (N_380,In_572,In_36);
nand U381 (N_381,In_574,N_154);
and U382 (N_382,In_596,In_249);
or U383 (N_383,In_366,N_164);
nand U384 (N_384,N_284,In_392);
nand U385 (N_385,In_469,N_103);
and U386 (N_386,N_137,N_258);
xor U387 (N_387,N_19,N_229);
nand U388 (N_388,N_100,N_112);
nand U389 (N_389,N_249,N_201);
xnor U390 (N_390,In_749,N_259);
nor U391 (N_391,In_543,In_220);
nand U392 (N_392,In_336,N_267);
xor U393 (N_393,N_145,N_260);
nor U394 (N_394,In_463,In_576);
xnor U395 (N_395,N_169,In_531);
nand U396 (N_396,N_117,In_260);
and U397 (N_397,N_170,N_287);
nand U398 (N_398,In_18,N_172);
nor U399 (N_399,N_15,In_154);
or U400 (N_400,N_289,In_515);
nand U401 (N_401,N_163,In_239);
nor U402 (N_402,N_316,N_271);
and U403 (N_403,N_38,In_539);
or U404 (N_404,In_433,N_182);
and U405 (N_405,N_123,In_81);
or U406 (N_406,N_273,N_310);
nand U407 (N_407,N_292,N_131);
nand U408 (N_408,N_395,In_362);
and U409 (N_409,N_269,In_553);
nand U410 (N_410,N_291,N_97);
nor U411 (N_411,N_203,N_39);
nand U412 (N_412,N_363,In_478);
or U413 (N_413,N_365,N_351);
nand U414 (N_414,N_24,In_151);
and U415 (N_415,In_466,N_186);
or U416 (N_416,N_31,N_54);
nand U417 (N_417,In_14,In_486);
or U418 (N_418,N_379,N_393);
nor U419 (N_419,In_652,In_591);
xor U420 (N_420,In_402,N_5);
xor U421 (N_421,N_396,In_726);
and U422 (N_422,N_366,In_375);
xor U423 (N_423,N_357,In_519);
nor U424 (N_424,N_69,N_326);
and U425 (N_425,N_98,N_323);
and U426 (N_426,N_313,N_345);
and U427 (N_427,In_219,N_8);
or U428 (N_428,In_172,N_359);
nand U429 (N_429,N_67,In_23);
nand U430 (N_430,In_549,In_213);
nor U431 (N_431,N_36,N_111);
nand U432 (N_432,N_327,N_382);
nand U433 (N_433,N_295,N_166);
xnor U434 (N_434,N_319,N_302);
nand U435 (N_435,In_333,In_557);
and U436 (N_436,In_315,In_252);
xnor U437 (N_437,In_473,In_432);
nand U438 (N_438,In_428,N_373);
nor U439 (N_439,N_341,In_85);
or U440 (N_440,N_335,N_300);
nor U441 (N_441,In_688,N_349);
nor U442 (N_442,In_319,N_356);
or U443 (N_443,In_526,N_187);
nand U444 (N_444,In_284,N_301);
or U445 (N_445,N_26,N_256);
or U446 (N_446,N_204,N_297);
nand U447 (N_447,In_19,In_620);
or U448 (N_448,N_391,In_29);
xnor U449 (N_449,N_304,N_143);
nand U450 (N_450,N_312,N_58);
and U451 (N_451,In_146,In_295);
and U452 (N_452,In_482,In_711);
xor U453 (N_453,N_378,N_339);
nand U454 (N_454,N_387,N_17);
nand U455 (N_455,In_585,In_460);
or U456 (N_456,In_513,N_232);
nor U457 (N_457,In_20,In_165);
and U458 (N_458,In_569,In_347);
xor U459 (N_459,N_369,N_372);
nor U460 (N_460,N_21,In_121);
nor U461 (N_461,N_194,N_209);
or U462 (N_462,In_720,N_306);
nand U463 (N_463,N_336,N_210);
or U464 (N_464,In_579,N_11);
or U465 (N_465,In_587,N_320);
or U466 (N_466,In_31,N_152);
nor U467 (N_467,N_334,N_399);
xnor U468 (N_468,In_114,In_494);
or U469 (N_469,In_393,N_242);
nor U470 (N_470,N_347,N_61);
nand U471 (N_471,In_708,N_348);
xnor U472 (N_472,In_119,N_381);
nand U473 (N_473,N_309,In_190);
and U474 (N_474,In_684,N_196);
or U475 (N_475,N_308,N_188);
nor U476 (N_476,N_376,N_80);
nand U477 (N_477,In_481,N_248);
nand U478 (N_478,In_242,N_370);
nand U479 (N_479,N_315,In_180);
and U480 (N_480,N_127,In_655);
and U481 (N_481,N_314,N_114);
nand U482 (N_482,N_113,N_25);
xor U483 (N_483,In_405,N_40);
xnor U484 (N_484,In_644,N_278);
and U485 (N_485,N_350,In_651);
and U486 (N_486,In_189,N_331);
and U487 (N_487,N_257,N_352);
and U488 (N_488,N_129,In_680);
and U489 (N_489,In_631,N_342);
and U490 (N_490,In_110,In_47);
nand U491 (N_491,N_274,N_374);
xor U492 (N_492,In_452,N_383);
xor U493 (N_493,N_385,In_138);
nand U494 (N_494,In_372,In_21);
nand U495 (N_495,N_18,N_227);
nand U496 (N_496,In_497,In_251);
and U497 (N_497,N_207,In_447);
or U498 (N_498,N_225,N_311);
and U499 (N_499,N_333,N_179);
and U500 (N_500,N_490,In_290);
xnor U501 (N_501,In_212,N_364);
nand U502 (N_502,N_234,N_430);
nor U503 (N_503,N_390,N_453);
xor U504 (N_504,N_459,N_264);
and U505 (N_505,In_678,In_133);
nand U506 (N_506,N_464,In_324);
and U507 (N_507,N_438,N_435);
and U508 (N_508,N_266,In_545);
xor U509 (N_509,N_427,N_398);
nor U510 (N_510,N_118,N_226);
nor U511 (N_511,N_299,N_151);
nand U512 (N_512,N_487,N_484);
or U513 (N_513,N_474,N_448);
or U514 (N_514,N_451,N_404);
xor U515 (N_515,N_405,N_16);
xor U516 (N_516,N_449,N_472);
xnor U517 (N_517,N_79,N_478);
or U518 (N_518,In_421,N_238);
xor U519 (N_519,N_442,In_493);
nor U520 (N_520,In_244,In_179);
xnor U521 (N_521,N_34,N_463);
xnor U522 (N_522,In_438,N_461);
xor U523 (N_523,N_237,N_475);
xor U524 (N_524,N_414,N_486);
nor U525 (N_525,N_424,N_222);
nor U526 (N_526,In_175,N_489);
xnor U527 (N_527,N_298,N_9);
xor U528 (N_528,In_363,N_185);
and U529 (N_529,N_230,In_485);
nand U530 (N_530,N_467,N_322);
nor U531 (N_531,N_441,N_468);
and U532 (N_532,N_494,N_12);
or U533 (N_533,N_215,In_164);
nand U534 (N_534,N_217,N_434);
or U535 (N_535,In_436,N_148);
nand U536 (N_536,N_321,N_135);
or U537 (N_537,N_317,In_407);
nor U538 (N_538,N_202,In_521);
xnor U539 (N_539,N_43,N_403);
or U540 (N_540,N_457,N_388);
nand U541 (N_541,N_425,N_422);
xor U542 (N_542,N_498,N_456);
xnor U543 (N_543,N_418,In_211);
or U544 (N_544,N_368,N_412);
or U545 (N_545,N_361,N_277);
or U546 (N_546,N_429,N_346);
nand U547 (N_547,N_481,In_35);
nor U548 (N_548,N_416,N_397);
nor U549 (N_549,N_324,In_40);
nand U550 (N_550,In_456,N_446);
nand U551 (N_551,In_537,N_375);
and U552 (N_552,N_466,In_218);
nand U553 (N_553,N_329,N_450);
xor U554 (N_554,In_623,N_389);
nor U555 (N_555,N_465,N_307);
and U556 (N_556,N_355,N_362);
nand U557 (N_557,N_86,N_421);
nor U558 (N_558,N_254,In_348);
and U559 (N_559,N_318,N_426);
or U560 (N_560,N_340,N_443);
nor U561 (N_561,N_121,In_554);
nand U562 (N_562,In_82,N_354);
and U563 (N_563,N_437,N_402);
and U564 (N_564,N_407,N_485);
xnor U565 (N_565,N_262,In_221);
nor U566 (N_566,N_330,N_439);
or U567 (N_567,N_410,In_367);
nand U568 (N_568,In_530,N_483);
or U569 (N_569,N_455,N_400);
and U570 (N_570,N_462,In_727);
and U571 (N_571,N_343,N_497);
nor U572 (N_572,In_228,In_592);
nor U573 (N_573,N_495,N_433);
or U574 (N_574,N_394,N_371);
or U575 (N_575,N_332,N_174);
xnor U576 (N_576,N_401,N_447);
xor U577 (N_577,In_674,N_190);
nor U578 (N_578,N_431,N_496);
and U579 (N_579,In_269,N_367);
xor U580 (N_580,In_492,N_305);
xor U581 (N_581,In_470,N_199);
or U582 (N_582,N_488,N_476);
xor U583 (N_583,In_710,In_46);
or U584 (N_584,N_415,N_205);
or U585 (N_585,N_471,In_423);
xnor U586 (N_586,N_477,In_25);
nand U587 (N_587,N_290,N_286);
and U588 (N_588,In_305,N_419);
or U589 (N_589,N_380,N_353);
nand U590 (N_590,N_469,In_629);
or U591 (N_591,In_273,In_606);
nor U592 (N_592,N_344,N_413);
nand U593 (N_593,N_296,N_432);
nand U594 (N_594,N_491,N_360);
nor U595 (N_595,N_444,N_138);
and U596 (N_596,N_377,N_411);
nand U597 (N_597,N_492,N_452);
or U598 (N_598,N_4,N_406);
and U599 (N_599,N_440,N_417);
nand U600 (N_600,N_545,N_579);
or U601 (N_601,N_116,N_544);
xor U602 (N_602,N_384,N_328);
or U603 (N_603,N_239,N_445);
xor U604 (N_604,N_566,N_420);
nand U605 (N_605,In_713,N_358);
or U606 (N_606,N_550,N_569);
nor U607 (N_607,N_516,N_565);
nor U608 (N_608,N_505,N_436);
xnor U609 (N_609,N_303,N_428);
nand U610 (N_610,N_500,N_325);
nor U611 (N_611,N_275,N_521);
nor U612 (N_612,N_558,In_415);
nor U613 (N_613,N_338,N_538);
xnor U614 (N_614,N_525,N_573);
nand U615 (N_615,N_535,N_512);
xor U616 (N_616,N_567,N_574);
xnor U617 (N_617,N_582,N_502);
and U618 (N_618,N_571,In_93);
xor U619 (N_619,N_122,N_564);
and U620 (N_620,N_233,In_533);
xor U621 (N_621,N_510,N_524);
nor U622 (N_622,N_529,N_557);
or U623 (N_623,N_515,N_597);
nand U624 (N_624,N_562,N_568);
nand U625 (N_625,N_585,N_460);
and U626 (N_626,In_125,N_243);
nor U627 (N_627,N_526,N_479);
xnor U628 (N_628,N_563,N_531);
nand U629 (N_629,N_480,N_556);
or U630 (N_630,N_540,N_530);
xor U631 (N_631,N_473,N_282);
xor U632 (N_632,N_482,N_553);
nand U633 (N_633,N_546,N_596);
and U634 (N_634,N_136,N_586);
xnor U635 (N_635,N_507,In_627);
nand U636 (N_636,N_337,N_509);
nor U637 (N_637,N_208,N_583);
nor U638 (N_638,N_386,N_547);
and U639 (N_639,N_551,N_409);
or U640 (N_640,N_408,N_454);
nor U641 (N_641,N_533,N_519);
nor U642 (N_642,N_548,N_523);
xnor U643 (N_643,N_552,N_105);
xor U644 (N_644,In_181,N_576);
or U645 (N_645,N_581,N_541);
nand U646 (N_646,N_584,N_578);
nor U647 (N_647,N_102,N_514);
nand U648 (N_648,N_149,N_537);
or U649 (N_649,In_660,N_518);
and U650 (N_650,N_392,N_588);
or U651 (N_651,N_458,N_572);
xnor U652 (N_652,N_511,N_527);
xor U653 (N_653,N_506,N_528);
xor U654 (N_654,In_445,N_577);
xnor U655 (N_655,N_592,N_587);
xor U656 (N_656,N_470,N_560);
xnor U657 (N_657,N_590,N_501);
nand U658 (N_658,In_334,N_595);
and U659 (N_659,N_534,N_593);
nand U660 (N_660,N_598,N_508);
or U661 (N_661,N_594,N_591);
xnor U662 (N_662,N_555,N_580);
or U663 (N_663,N_549,N_542);
or U664 (N_664,N_599,N_570);
nand U665 (N_665,N_561,N_493);
nor U666 (N_666,N_539,N_554);
nor U667 (N_667,N_513,In_137);
and U668 (N_668,N_517,N_423);
nor U669 (N_669,N_178,N_543);
nor U670 (N_670,N_532,N_520);
nand U671 (N_671,N_499,N_559);
nand U672 (N_672,N_575,N_589);
nand U673 (N_673,N_503,N_504);
nor U674 (N_674,N_522,N_536);
or U675 (N_675,N_502,In_334);
or U676 (N_676,N_542,N_358);
or U677 (N_677,N_517,N_558);
nand U678 (N_678,N_515,N_392);
and U679 (N_679,N_520,N_508);
or U680 (N_680,N_501,N_524);
nand U681 (N_681,N_597,N_567);
and U682 (N_682,N_420,N_384);
nand U683 (N_683,N_574,N_208);
nor U684 (N_684,N_445,N_543);
nand U685 (N_685,N_592,In_415);
and U686 (N_686,N_533,N_572);
nor U687 (N_687,N_510,N_499);
and U688 (N_688,N_558,N_509);
nor U689 (N_689,N_529,N_275);
nand U690 (N_690,N_579,N_520);
and U691 (N_691,N_545,N_537);
and U692 (N_692,N_574,N_571);
nor U693 (N_693,N_541,N_537);
or U694 (N_694,N_539,N_337);
xnor U695 (N_695,N_584,N_582);
xor U696 (N_696,N_479,N_592);
xor U697 (N_697,N_358,N_582);
xnor U698 (N_698,N_445,In_713);
nor U699 (N_699,In_93,N_552);
xor U700 (N_700,N_612,N_602);
and U701 (N_701,N_685,N_604);
and U702 (N_702,N_682,N_681);
or U703 (N_703,N_607,N_649);
nor U704 (N_704,N_621,N_666);
and U705 (N_705,N_673,N_640);
xnor U706 (N_706,N_661,N_695);
nand U707 (N_707,N_675,N_655);
or U708 (N_708,N_638,N_671);
or U709 (N_709,N_687,N_636);
and U710 (N_710,N_658,N_650);
nor U711 (N_711,N_644,N_656);
or U712 (N_712,N_698,N_635);
or U713 (N_713,N_611,N_680);
or U714 (N_714,N_679,N_603);
or U715 (N_715,N_696,N_631);
nand U716 (N_716,N_677,N_660);
nand U717 (N_717,N_665,N_615);
and U718 (N_718,N_618,N_668);
or U719 (N_719,N_624,N_657);
xnor U720 (N_720,N_625,N_630);
and U721 (N_721,N_689,N_647);
or U722 (N_722,N_676,N_648);
xor U723 (N_723,N_691,N_632);
and U724 (N_724,N_652,N_645);
nor U725 (N_725,N_606,N_667);
or U726 (N_726,N_654,N_684);
and U727 (N_727,N_626,N_659);
or U728 (N_728,N_651,N_646);
or U729 (N_729,N_692,N_608);
xnor U730 (N_730,N_669,N_664);
nand U731 (N_731,N_623,N_683);
nand U732 (N_732,N_616,N_633);
or U733 (N_733,N_663,N_617);
xor U734 (N_734,N_653,N_642);
nand U735 (N_735,N_619,N_641);
and U736 (N_736,N_622,N_699);
nor U737 (N_737,N_672,N_605);
nand U738 (N_738,N_600,N_627);
nand U739 (N_739,N_670,N_694);
nor U740 (N_740,N_614,N_674);
xor U741 (N_741,N_629,N_678);
and U742 (N_742,N_662,N_639);
xnor U743 (N_743,N_697,N_601);
and U744 (N_744,N_637,N_686);
nand U745 (N_745,N_688,N_610);
and U746 (N_746,N_690,N_643);
xor U747 (N_747,N_620,N_609);
xor U748 (N_748,N_613,N_634);
and U749 (N_749,N_693,N_628);
and U750 (N_750,N_627,N_680);
nand U751 (N_751,N_661,N_615);
nor U752 (N_752,N_682,N_602);
xnor U753 (N_753,N_671,N_632);
xnor U754 (N_754,N_642,N_662);
nand U755 (N_755,N_600,N_678);
or U756 (N_756,N_655,N_682);
xor U757 (N_757,N_651,N_655);
or U758 (N_758,N_648,N_681);
nor U759 (N_759,N_634,N_668);
xnor U760 (N_760,N_614,N_655);
nand U761 (N_761,N_642,N_677);
and U762 (N_762,N_620,N_699);
and U763 (N_763,N_650,N_641);
xor U764 (N_764,N_691,N_665);
xnor U765 (N_765,N_627,N_689);
or U766 (N_766,N_689,N_601);
nand U767 (N_767,N_679,N_601);
or U768 (N_768,N_657,N_655);
nand U769 (N_769,N_679,N_620);
xor U770 (N_770,N_653,N_675);
nor U771 (N_771,N_669,N_672);
and U772 (N_772,N_662,N_636);
xnor U773 (N_773,N_616,N_628);
or U774 (N_774,N_661,N_666);
nor U775 (N_775,N_672,N_609);
and U776 (N_776,N_646,N_614);
or U777 (N_777,N_607,N_676);
and U778 (N_778,N_648,N_686);
nor U779 (N_779,N_699,N_698);
nand U780 (N_780,N_608,N_684);
or U781 (N_781,N_624,N_675);
nor U782 (N_782,N_624,N_683);
and U783 (N_783,N_649,N_671);
or U784 (N_784,N_641,N_671);
xor U785 (N_785,N_678,N_672);
nand U786 (N_786,N_619,N_611);
or U787 (N_787,N_601,N_670);
or U788 (N_788,N_669,N_682);
and U789 (N_789,N_608,N_678);
nor U790 (N_790,N_603,N_647);
nor U791 (N_791,N_614,N_624);
nor U792 (N_792,N_646,N_664);
nand U793 (N_793,N_625,N_614);
nor U794 (N_794,N_681,N_646);
xnor U795 (N_795,N_681,N_668);
nand U796 (N_796,N_627,N_697);
nor U797 (N_797,N_615,N_631);
and U798 (N_798,N_615,N_668);
xor U799 (N_799,N_689,N_684);
and U800 (N_800,N_710,N_731);
and U801 (N_801,N_770,N_751);
and U802 (N_802,N_713,N_759);
xor U803 (N_803,N_747,N_795);
nor U804 (N_804,N_715,N_793);
and U805 (N_805,N_797,N_704);
and U806 (N_806,N_789,N_788);
nor U807 (N_807,N_727,N_722);
or U808 (N_808,N_737,N_721);
xor U809 (N_809,N_777,N_706);
or U810 (N_810,N_746,N_753);
and U811 (N_811,N_714,N_718);
xnor U812 (N_812,N_728,N_717);
or U813 (N_813,N_740,N_776);
or U814 (N_814,N_739,N_734);
and U815 (N_815,N_796,N_700);
xor U816 (N_816,N_732,N_744);
xnor U817 (N_817,N_768,N_754);
xor U818 (N_818,N_764,N_772);
and U819 (N_819,N_729,N_750);
nand U820 (N_820,N_765,N_798);
xor U821 (N_821,N_709,N_758);
and U822 (N_822,N_762,N_785);
and U823 (N_823,N_703,N_786);
xnor U824 (N_824,N_712,N_743);
nand U825 (N_825,N_749,N_752);
nand U826 (N_826,N_730,N_735);
xnor U827 (N_827,N_724,N_707);
xor U828 (N_828,N_711,N_792);
nor U829 (N_829,N_773,N_733);
xor U830 (N_830,N_779,N_726);
or U831 (N_831,N_736,N_799);
and U832 (N_832,N_720,N_738);
nand U833 (N_833,N_784,N_783);
nor U834 (N_834,N_767,N_719);
nand U835 (N_835,N_756,N_790);
xor U836 (N_836,N_725,N_769);
or U837 (N_837,N_701,N_774);
and U838 (N_838,N_761,N_771);
nor U839 (N_839,N_787,N_748);
and U840 (N_840,N_741,N_791);
xor U841 (N_841,N_708,N_760);
nor U842 (N_842,N_742,N_780);
and U843 (N_843,N_723,N_766);
xor U844 (N_844,N_763,N_755);
or U845 (N_845,N_775,N_702);
xor U846 (N_846,N_716,N_757);
nand U847 (N_847,N_745,N_778);
and U848 (N_848,N_782,N_794);
xor U849 (N_849,N_705,N_781);
nor U850 (N_850,N_767,N_700);
or U851 (N_851,N_729,N_710);
nor U852 (N_852,N_775,N_716);
xor U853 (N_853,N_738,N_742);
xnor U854 (N_854,N_777,N_707);
xor U855 (N_855,N_796,N_749);
nor U856 (N_856,N_755,N_772);
or U857 (N_857,N_747,N_721);
nand U858 (N_858,N_784,N_713);
xor U859 (N_859,N_791,N_769);
xor U860 (N_860,N_752,N_737);
or U861 (N_861,N_786,N_774);
nor U862 (N_862,N_733,N_757);
nor U863 (N_863,N_710,N_788);
or U864 (N_864,N_782,N_774);
and U865 (N_865,N_744,N_735);
and U866 (N_866,N_765,N_732);
and U867 (N_867,N_728,N_762);
and U868 (N_868,N_719,N_725);
or U869 (N_869,N_717,N_772);
nor U870 (N_870,N_758,N_759);
or U871 (N_871,N_755,N_762);
or U872 (N_872,N_790,N_737);
nor U873 (N_873,N_794,N_774);
nand U874 (N_874,N_778,N_701);
and U875 (N_875,N_743,N_714);
and U876 (N_876,N_710,N_714);
xnor U877 (N_877,N_788,N_741);
nand U878 (N_878,N_718,N_717);
and U879 (N_879,N_759,N_798);
xnor U880 (N_880,N_724,N_701);
or U881 (N_881,N_756,N_761);
nand U882 (N_882,N_748,N_751);
or U883 (N_883,N_735,N_777);
nor U884 (N_884,N_732,N_721);
nor U885 (N_885,N_775,N_760);
nor U886 (N_886,N_702,N_768);
and U887 (N_887,N_792,N_725);
nand U888 (N_888,N_732,N_707);
and U889 (N_889,N_707,N_749);
nor U890 (N_890,N_782,N_730);
nor U891 (N_891,N_792,N_785);
nand U892 (N_892,N_740,N_728);
nand U893 (N_893,N_768,N_791);
or U894 (N_894,N_703,N_729);
xor U895 (N_895,N_774,N_720);
nand U896 (N_896,N_759,N_799);
nor U897 (N_897,N_783,N_724);
nand U898 (N_898,N_729,N_783);
nand U899 (N_899,N_759,N_745);
nor U900 (N_900,N_842,N_809);
nor U901 (N_901,N_838,N_897);
or U902 (N_902,N_893,N_858);
nand U903 (N_903,N_856,N_810);
and U904 (N_904,N_837,N_877);
and U905 (N_905,N_881,N_863);
nor U906 (N_906,N_879,N_896);
nand U907 (N_907,N_872,N_825);
and U908 (N_908,N_873,N_841);
xor U909 (N_909,N_829,N_867);
or U910 (N_910,N_828,N_815);
nand U911 (N_911,N_851,N_826);
and U912 (N_912,N_862,N_824);
xor U913 (N_913,N_865,N_871);
xnor U914 (N_914,N_875,N_857);
xor U915 (N_915,N_866,N_860);
nand U916 (N_916,N_806,N_853);
xor U917 (N_917,N_822,N_868);
nand U918 (N_918,N_852,N_805);
nand U919 (N_919,N_861,N_820);
nand U920 (N_920,N_884,N_869);
nor U921 (N_921,N_899,N_814);
nor U922 (N_922,N_804,N_882);
nor U923 (N_923,N_887,N_812);
nand U924 (N_924,N_850,N_878);
xor U925 (N_925,N_808,N_874);
nand U926 (N_926,N_880,N_803);
nand U927 (N_927,N_885,N_895);
xor U928 (N_928,N_832,N_883);
xnor U929 (N_929,N_839,N_898);
or U930 (N_930,N_864,N_849);
nand U931 (N_931,N_876,N_807);
nor U932 (N_932,N_801,N_821);
or U933 (N_933,N_889,N_811);
xor U934 (N_934,N_890,N_848);
nand U935 (N_935,N_836,N_859);
and U936 (N_936,N_813,N_817);
nand U937 (N_937,N_854,N_802);
or U938 (N_938,N_891,N_855);
or U939 (N_939,N_886,N_892);
xnor U940 (N_940,N_830,N_846);
or U941 (N_941,N_894,N_840);
xor U942 (N_942,N_800,N_888);
or U943 (N_943,N_870,N_845);
xnor U944 (N_944,N_827,N_844);
nand U945 (N_945,N_816,N_819);
or U946 (N_946,N_834,N_847);
nand U947 (N_947,N_833,N_835);
or U948 (N_948,N_823,N_843);
nor U949 (N_949,N_831,N_818);
xor U950 (N_950,N_888,N_809);
xor U951 (N_951,N_874,N_889);
and U952 (N_952,N_885,N_864);
and U953 (N_953,N_811,N_861);
and U954 (N_954,N_874,N_878);
and U955 (N_955,N_863,N_809);
and U956 (N_956,N_852,N_863);
nor U957 (N_957,N_876,N_800);
nand U958 (N_958,N_846,N_832);
and U959 (N_959,N_867,N_834);
xor U960 (N_960,N_879,N_835);
and U961 (N_961,N_872,N_867);
or U962 (N_962,N_855,N_892);
and U963 (N_963,N_840,N_851);
xnor U964 (N_964,N_882,N_816);
xor U965 (N_965,N_885,N_897);
xor U966 (N_966,N_816,N_878);
nand U967 (N_967,N_877,N_847);
nor U968 (N_968,N_862,N_856);
or U969 (N_969,N_858,N_872);
or U970 (N_970,N_878,N_890);
or U971 (N_971,N_820,N_849);
xor U972 (N_972,N_812,N_835);
or U973 (N_973,N_819,N_810);
or U974 (N_974,N_895,N_826);
or U975 (N_975,N_832,N_875);
or U976 (N_976,N_801,N_897);
or U977 (N_977,N_868,N_853);
or U978 (N_978,N_859,N_864);
and U979 (N_979,N_834,N_801);
nand U980 (N_980,N_843,N_824);
nand U981 (N_981,N_874,N_866);
nor U982 (N_982,N_801,N_862);
and U983 (N_983,N_842,N_876);
nor U984 (N_984,N_803,N_861);
or U985 (N_985,N_861,N_830);
xnor U986 (N_986,N_851,N_815);
nor U987 (N_987,N_894,N_823);
nand U988 (N_988,N_824,N_864);
and U989 (N_989,N_879,N_885);
xor U990 (N_990,N_842,N_857);
and U991 (N_991,N_800,N_851);
nor U992 (N_992,N_870,N_895);
or U993 (N_993,N_880,N_816);
and U994 (N_994,N_831,N_879);
or U995 (N_995,N_810,N_869);
nor U996 (N_996,N_898,N_877);
nor U997 (N_997,N_811,N_804);
nand U998 (N_998,N_891,N_876);
or U999 (N_999,N_854,N_815);
xor U1000 (N_1000,N_990,N_914);
and U1001 (N_1001,N_969,N_919);
nor U1002 (N_1002,N_995,N_986);
and U1003 (N_1003,N_911,N_955);
nand U1004 (N_1004,N_976,N_987);
nand U1005 (N_1005,N_944,N_982);
xnor U1006 (N_1006,N_979,N_915);
or U1007 (N_1007,N_994,N_958);
nand U1008 (N_1008,N_943,N_967);
or U1009 (N_1009,N_968,N_903);
nor U1010 (N_1010,N_934,N_908);
nand U1011 (N_1011,N_907,N_930);
and U1012 (N_1012,N_929,N_912);
and U1013 (N_1013,N_946,N_950);
nand U1014 (N_1014,N_974,N_977);
xnor U1015 (N_1015,N_952,N_928);
nand U1016 (N_1016,N_953,N_961);
nor U1017 (N_1017,N_998,N_945);
and U1018 (N_1018,N_947,N_920);
xor U1019 (N_1019,N_931,N_988);
nor U1020 (N_1020,N_972,N_983);
nor U1021 (N_1021,N_923,N_993);
nor U1022 (N_1022,N_922,N_924);
xnor U1023 (N_1023,N_939,N_978);
nand U1024 (N_1024,N_999,N_933);
and U1025 (N_1025,N_949,N_992);
nand U1026 (N_1026,N_954,N_970);
or U1027 (N_1027,N_925,N_917);
or U1028 (N_1028,N_940,N_965);
nand U1029 (N_1029,N_900,N_918);
and U1030 (N_1030,N_938,N_962);
or U1031 (N_1031,N_981,N_913);
nor U1032 (N_1032,N_926,N_996);
or U1033 (N_1033,N_960,N_984);
and U1034 (N_1034,N_941,N_906);
nor U1035 (N_1035,N_909,N_905);
or U1036 (N_1036,N_956,N_980);
xor U1037 (N_1037,N_989,N_904);
or U1038 (N_1038,N_921,N_997);
nor U1039 (N_1039,N_991,N_932);
nor U1040 (N_1040,N_957,N_942);
and U1041 (N_1041,N_985,N_902);
or U1042 (N_1042,N_963,N_951);
xnor U1043 (N_1043,N_935,N_959);
nand U1044 (N_1044,N_936,N_910);
xor U1045 (N_1045,N_901,N_948);
nand U1046 (N_1046,N_937,N_971);
xor U1047 (N_1047,N_964,N_973);
and U1048 (N_1048,N_916,N_927);
or U1049 (N_1049,N_966,N_975);
xor U1050 (N_1050,N_939,N_973);
xnor U1051 (N_1051,N_925,N_957);
nor U1052 (N_1052,N_924,N_990);
nor U1053 (N_1053,N_965,N_935);
nand U1054 (N_1054,N_963,N_946);
nor U1055 (N_1055,N_914,N_946);
nand U1056 (N_1056,N_905,N_952);
and U1057 (N_1057,N_902,N_969);
and U1058 (N_1058,N_931,N_963);
nor U1059 (N_1059,N_943,N_984);
nand U1060 (N_1060,N_964,N_978);
and U1061 (N_1061,N_943,N_928);
nor U1062 (N_1062,N_903,N_956);
xnor U1063 (N_1063,N_933,N_989);
and U1064 (N_1064,N_951,N_982);
xor U1065 (N_1065,N_959,N_925);
or U1066 (N_1066,N_994,N_916);
and U1067 (N_1067,N_903,N_913);
nor U1068 (N_1068,N_967,N_954);
or U1069 (N_1069,N_928,N_929);
xnor U1070 (N_1070,N_984,N_972);
xnor U1071 (N_1071,N_915,N_946);
nand U1072 (N_1072,N_941,N_949);
and U1073 (N_1073,N_924,N_953);
nand U1074 (N_1074,N_905,N_963);
xor U1075 (N_1075,N_979,N_909);
nor U1076 (N_1076,N_918,N_915);
or U1077 (N_1077,N_972,N_994);
xnor U1078 (N_1078,N_934,N_994);
nor U1079 (N_1079,N_904,N_937);
and U1080 (N_1080,N_978,N_901);
or U1081 (N_1081,N_931,N_906);
and U1082 (N_1082,N_989,N_945);
and U1083 (N_1083,N_998,N_906);
xor U1084 (N_1084,N_924,N_986);
and U1085 (N_1085,N_916,N_940);
xor U1086 (N_1086,N_977,N_908);
and U1087 (N_1087,N_941,N_980);
nor U1088 (N_1088,N_937,N_911);
or U1089 (N_1089,N_953,N_988);
nand U1090 (N_1090,N_993,N_902);
xnor U1091 (N_1091,N_981,N_910);
xor U1092 (N_1092,N_965,N_968);
xor U1093 (N_1093,N_996,N_991);
or U1094 (N_1094,N_950,N_958);
xor U1095 (N_1095,N_978,N_916);
nor U1096 (N_1096,N_919,N_992);
nand U1097 (N_1097,N_992,N_905);
nor U1098 (N_1098,N_924,N_912);
and U1099 (N_1099,N_966,N_963);
nor U1100 (N_1100,N_1098,N_1002);
or U1101 (N_1101,N_1090,N_1009);
nand U1102 (N_1102,N_1060,N_1062);
nand U1103 (N_1103,N_1017,N_1069);
and U1104 (N_1104,N_1032,N_1046);
or U1105 (N_1105,N_1038,N_1013);
or U1106 (N_1106,N_1063,N_1048);
or U1107 (N_1107,N_1053,N_1083);
and U1108 (N_1108,N_1040,N_1051);
xnor U1109 (N_1109,N_1037,N_1054);
or U1110 (N_1110,N_1057,N_1097);
nor U1111 (N_1111,N_1079,N_1014);
and U1112 (N_1112,N_1024,N_1094);
and U1113 (N_1113,N_1036,N_1042);
xnor U1114 (N_1114,N_1049,N_1095);
xnor U1115 (N_1115,N_1044,N_1075);
or U1116 (N_1116,N_1096,N_1004);
nand U1117 (N_1117,N_1064,N_1021);
nor U1118 (N_1118,N_1065,N_1025);
nor U1119 (N_1119,N_1091,N_1022);
nand U1120 (N_1120,N_1047,N_1099);
and U1121 (N_1121,N_1039,N_1007);
xor U1122 (N_1122,N_1071,N_1061);
nand U1123 (N_1123,N_1029,N_1016);
nand U1124 (N_1124,N_1066,N_1005);
or U1125 (N_1125,N_1081,N_1068);
and U1126 (N_1126,N_1001,N_1010);
xor U1127 (N_1127,N_1019,N_1092);
xnor U1128 (N_1128,N_1052,N_1006);
nand U1129 (N_1129,N_1076,N_1035);
nand U1130 (N_1130,N_1018,N_1078);
and U1131 (N_1131,N_1067,N_1050);
nor U1132 (N_1132,N_1033,N_1086);
xor U1133 (N_1133,N_1056,N_1093);
or U1134 (N_1134,N_1027,N_1058);
nand U1135 (N_1135,N_1011,N_1088);
and U1136 (N_1136,N_1023,N_1031);
nor U1137 (N_1137,N_1000,N_1028);
or U1138 (N_1138,N_1077,N_1080);
nand U1139 (N_1139,N_1003,N_1084);
nand U1140 (N_1140,N_1026,N_1030);
nor U1141 (N_1141,N_1070,N_1087);
or U1142 (N_1142,N_1089,N_1072);
xor U1143 (N_1143,N_1012,N_1020);
nand U1144 (N_1144,N_1059,N_1043);
and U1145 (N_1145,N_1008,N_1073);
nand U1146 (N_1146,N_1074,N_1015);
and U1147 (N_1147,N_1085,N_1045);
xor U1148 (N_1148,N_1082,N_1041);
xnor U1149 (N_1149,N_1034,N_1055);
or U1150 (N_1150,N_1034,N_1098);
nand U1151 (N_1151,N_1061,N_1023);
nand U1152 (N_1152,N_1057,N_1000);
nor U1153 (N_1153,N_1061,N_1082);
or U1154 (N_1154,N_1087,N_1029);
or U1155 (N_1155,N_1030,N_1090);
nor U1156 (N_1156,N_1076,N_1007);
nor U1157 (N_1157,N_1011,N_1078);
or U1158 (N_1158,N_1011,N_1041);
nor U1159 (N_1159,N_1006,N_1076);
nor U1160 (N_1160,N_1051,N_1041);
nor U1161 (N_1161,N_1023,N_1008);
nor U1162 (N_1162,N_1022,N_1040);
nand U1163 (N_1163,N_1033,N_1088);
xor U1164 (N_1164,N_1004,N_1089);
xor U1165 (N_1165,N_1085,N_1086);
and U1166 (N_1166,N_1094,N_1090);
and U1167 (N_1167,N_1053,N_1012);
or U1168 (N_1168,N_1043,N_1017);
and U1169 (N_1169,N_1012,N_1089);
xnor U1170 (N_1170,N_1067,N_1066);
and U1171 (N_1171,N_1078,N_1060);
nor U1172 (N_1172,N_1058,N_1084);
nor U1173 (N_1173,N_1084,N_1077);
xnor U1174 (N_1174,N_1097,N_1080);
xnor U1175 (N_1175,N_1048,N_1003);
nand U1176 (N_1176,N_1067,N_1073);
nor U1177 (N_1177,N_1052,N_1089);
xor U1178 (N_1178,N_1010,N_1022);
nor U1179 (N_1179,N_1080,N_1089);
or U1180 (N_1180,N_1092,N_1013);
xnor U1181 (N_1181,N_1075,N_1034);
or U1182 (N_1182,N_1091,N_1076);
and U1183 (N_1183,N_1095,N_1050);
or U1184 (N_1184,N_1067,N_1043);
or U1185 (N_1185,N_1042,N_1076);
xnor U1186 (N_1186,N_1024,N_1063);
nand U1187 (N_1187,N_1037,N_1076);
xor U1188 (N_1188,N_1099,N_1062);
nor U1189 (N_1189,N_1042,N_1035);
nor U1190 (N_1190,N_1017,N_1047);
nor U1191 (N_1191,N_1091,N_1062);
and U1192 (N_1192,N_1035,N_1086);
and U1193 (N_1193,N_1030,N_1010);
nor U1194 (N_1194,N_1086,N_1004);
xnor U1195 (N_1195,N_1018,N_1017);
nand U1196 (N_1196,N_1084,N_1094);
and U1197 (N_1197,N_1061,N_1035);
nand U1198 (N_1198,N_1030,N_1098);
nor U1199 (N_1199,N_1025,N_1075);
xnor U1200 (N_1200,N_1166,N_1103);
and U1201 (N_1201,N_1167,N_1133);
nor U1202 (N_1202,N_1100,N_1124);
nand U1203 (N_1203,N_1188,N_1164);
nor U1204 (N_1204,N_1180,N_1175);
nor U1205 (N_1205,N_1158,N_1184);
xnor U1206 (N_1206,N_1195,N_1185);
xor U1207 (N_1207,N_1109,N_1106);
nand U1208 (N_1208,N_1126,N_1147);
xor U1209 (N_1209,N_1150,N_1186);
xor U1210 (N_1210,N_1128,N_1125);
xor U1211 (N_1211,N_1148,N_1138);
or U1212 (N_1212,N_1122,N_1153);
nand U1213 (N_1213,N_1119,N_1162);
or U1214 (N_1214,N_1104,N_1169);
xnor U1215 (N_1215,N_1140,N_1105);
nor U1216 (N_1216,N_1145,N_1190);
and U1217 (N_1217,N_1107,N_1194);
xnor U1218 (N_1218,N_1179,N_1120);
or U1219 (N_1219,N_1102,N_1135);
or U1220 (N_1220,N_1193,N_1172);
or U1221 (N_1221,N_1192,N_1155);
or U1222 (N_1222,N_1141,N_1123);
nand U1223 (N_1223,N_1114,N_1161);
nand U1224 (N_1224,N_1127,N_1146);
and U1225 (N_1225,N_1165,N_1181);
and U1226 (N_1226,N_1110,N_1177);
xnor U1227 (N_1227,N_1160,N_1115);
nand U1228 (N_1228,N_1189,N_1159);
nand U1229 (N_1229,N_1163,N_1121);
nor U1230 (N_1230,N_1199,N_1113);
or U1231 (N_1231,N_1131,N_1174);
nor U1232 (N_1232,N_1118,N_1132);
nand U1233 (N_1233,N_1134,N_1111);
or U1234 (N_1234,N_1170,N_1144);
or U1235 (N_1235,N_1149,N_1143);
and U1236 (N_1236,N_1187,N_1197);
xor U1237 (N_1237,N_1183,N_1101);
xnor U1238 (N_1238,N_1154,N_1182);
nor U1239 (N_1239,N_1198,N_1171);
xor U1240 (N_1240,N_1178,N_1173);
and U1241 (N_1241,N_1168,N_1191);
and U1242 (N_1242,N_1108,N_1152);
and U1243 (N_1243,N_1142,N_1117);
or U1244 (N_1244,N_1137,N_1129);
and U1245 (N_1245,N_1156,N_1157);
nor U1246 (N_1246,N_1116,N_1196);
xnor U1247 (N_1247,N_1136,N_1130);
nand U1248 (N_1248,N_1176,N_1151);
nand U1249 (N_1249,N_1112,N_1139);
and U1250 (N_1250,N_1171,N_1105);
nor U1251 (N_1251,N_1187,N_1175);
or U1252 (N_1252,N_1127,N_1131);
or U1253 (N_1253,N_1192,N_1142);
or U1254 (N_1254,N_1157,N_1180);
nor U1255 (N_1255,N_1127,N_1184);
nand U1256 (N_1256,N_1135,N_1118);
or U1257 (N_1257,N_1158,N_1132);
nand U1258 (N_1258,N_1158,N_1140);
nor U1259 (N_1259,N_1179,N_1142);
nor U1260 (N_1260,N_1101,N_1126);
nand U1261 (N_1261,N_1153,N_1199);
and U1262 (N_1262,N_1199,N_1121);
nand U1263 (N_1263,N_1120,N_1113);
nand U1264 (N_1264,N_1123,N_1109);
and U1265 (N_1265,N_1114,N_1129);
nor U1266 (N_1266,N_1115,N_1194);
xnor U1267 (N_1267,N_1100,N_1113);
or U1268 (N_1268,N_1127,N_1139);
nand U1269 (N_1269,N_1111,N_1117);
nor U1270 (N_1270,N_1193,N_1127);
nand U1271 (N_1271,N_1177,N_1189);
nor U1272 (N_1272,N_1181,N_1112);
or U1273 (N_1273,N_1174,N_1144);
and U1274 (N_1274,N_1155,N_1159);
nand U1275 (N_1275,N_1123,N_1188);
nand U1276 (N_1276,N_1104,N_1195);
and U1277 (N_1277,N_1154,N_1148);
nand U1278 (N_1278,N_1186,N_1188);
or U1279 (N_1279,N_1109,N_1194);
or U1280 (N_1280,N_1118,N_1126);
xor U1281 (N_1281,N_1146,N_1139);
and U1282 (N_1282,N_1105,N_1148);
and U1283 (N_1283,N_1172,N_1138);
nor U1284 (N_1284,N_1171,N_1160);
or U1285 (N_1285,N_1142,N_1149);
nor U1286 (N_1286,N_1139,N_1183);
xor U1287 (N_1287,N_1115,N_1100);
nand U1288 (N_1288,N_1189,N_1104);
or U1289 (N_1289,N_1183,N_1128);
and U1290 (N_1290,N_1194,N_1108);
or U1291 (N_1291,N_1161,N_1199);
and U1292 (N_1292,N_1105,N_1170);
nor U1293 (N_1293,N_1157,N_1115);
nor U1294 (N_1294,N_1191,N_1120);
and U1295 (N_1295,N_1157,N_1173);
nor U1296 (N_1296,N_1168,N_1142);
and U1297 (N_1297,N_1184,N_1102);
or U1298 (N_1298,N_1137,N_1114);
or U1299 (N_1299,N_1121,N_1172);
or U1300 (N_1300,N_1208,N_1266);
and U1301 (N_1301,N_1217,N_1204);
and U1302 (N_1302,N_1238,N_1292);
nand U1303 (N_1303,N_1299,N_1214);
nor U1304 (N_1304,N_1267,N_1232);
nand U1305 (N_1305,N_1212,N_1222);
xnor U1306 (N_1306,N_1264,N_1234);
nand U1307 (N_1307,N_1275,N_1270);
nor U1308 (N_1308,N_1290,N_1298);
nand U1309 (N_1309,N_1269,N_1221);
or U1310 (N_1310,N_1211,N_1236);
xor U1311 (N_1311,N_1268,N_1274);
xor U1312 (N_1312,N_1285,N_1242);
or U1313 (N_1313,N_1227,N_1278);
and U1314 (N_1314,N_1287,N_1202);
nor U1315 (N_1315,N_1282,N_1226);
or U1316 (N_1316,N_1240,N_1250);
and U1317 (N_1317,N_1207,N_1233);
xnor U1318 (N_1318,N_1209,N_1294);
nand U1319 (N_1319,N_1205,N_1296);
or U1320 (N_1320,N_1223,N_1284);
and U1321 (N_1321,N_1289,N_1277);
or U1322 (N_1322,N_1248,N_1244);
nor U1323 (N_1323,N_1247,N_1215);
or U1324 (N_1324,N_1271,N_1262);
or U1325 (N_1325,N_1297,N_1256);
nor U1326 (N_1326,N_1260,N_1257);
nand U1327 (N_1327,N_1263,N_1276);
and U1328 (N_1328,N_1224,N_1246);
nand U1329 (N_1329,N_1206,N_1210);
nand U1330 (N_1330,N_1200,N_1225);
and U1331 (N_1331,N_1281,N_1295);
or U1332 (N_1332,N_1245,N_1235);
xor U1333 (N_1333,N_1291,N_1216);
nand U1334 (N_1334,N_1288,N_1293);
nor U1335 (N_1335,N_1230,N_1203);
nand U1336 (N_1336,N_1237,N_1273);
or U1337 (N_1337,N_1255,N_1251);
xnor U1338 (N_1338,N_1286,N_1253);
xor U1339 (N_1339,N_1231,N_1279);
and U1340 (N_1340,N_1261,N_1258);
or U1341 (N_1341,N_1239,N_1213);
nand U1342 (N_1342,N_1280,N_1243);
and U1343 (N_1343,N_1220,N_1259);
and U1344 (N_1344,N_1219,N_1241);
nand U1345 (N_1345,N_1201,N_1283);
and U1346 (N_1346,N_1249,N_1229);
or U1347 (N_1347,N_1218,N_1272);
or U1348 (N_1348,N_1265,N_1254);
xor U1349 (N_1349,N_1228,N_1252);
xor U1350 (N_1350,N_1282,N_1265);
nand U1351 (N_1351,N_1272,N_1274);
or U1352 (N_1352,N_1202,N_1264);
xnor U1353 (N_1353,N_1233,N_1294);
nor U1354 (N_1354,N_1264,N_1274);
or U1355 (N_1355,N_1250,N_1276);
or U1356 (N_1356,N_1268,N_1237);
and U1357 (N_1357,N_1263,N_1278);
and U1358 (N_1358,N_1221,N_1250);
xor U1359 (N_1359,N_1230,N_1265);
or U1360 (N_1360,N_1262,N_1238);
and U1361 (N_1361,N_1278,N_1242);
nor U1362 (N_1362,N_1260,N_1269);
xor U1363 (N_1363,N_1233,N_1224);
or U1364 (N_1364,N_1214,N_1260);
xor U1365 (N_1365,N_1250,N_1244);
and U1366 (N_1366,N_1276,N_1235);
and U1367 (N_1367,N_1205,N_1223);
nand U1368 (N_1368,N_1287,N_1290);
and U1369 (N_1369,N_1274,N_1206);
xor U1370 (N_1370,N_1219,N_1273);
and U1371 (N_1371,N_1262,N_1257);
xor U1372 (N_1372,N_1293,N_1295);
nor U1373 (N_1373,N_1290,N_1235);
or U1374 (N_1374,N_1279,N_1237);
nand U1375 (N_1375,N_1285,N_1230);
nand U1376 (N_1376,N_1231,N_1267);
nor U1377 (N_1377,N_1240,N_1252);
nand U1378 (N_1378,N_1200,N_1244);
or U1379 (N_1379,N_1259,N_1240);
xor U1380 (N_1380,N_1238,N_1229);
nor U1381 (N_1381,N_1275,N_1226);
or U1382 (N_1382,N_1244,N_1296);
and U1383 (N_1383,N_1239,N_1276);
xor U1384 (N_1384,N_1292,N_1269);
or U1385 (N_1385,N_1252,N_1219);
nand U1386 (N_1386,N_1266,N_1285);
and U1387 (N_1387,N_1244,N_1223);
nand U1388 (N_1388,N_1253,N_1235);
nand U1389 (N_1389,N_1248,N_1231);
nand U1390 (N_1390,N_1260,N_1220);
xnor U1391 (N_1391,N_1210,N_1242);
xnor U1392 (N_1392,N_1216,N_1241);
xor U1393 (N_1393,N_1256,N_1219);
nor U1394 (N_1394,N_1210,N_1293);
and U1395 (N_1395,N_1239,N_1216);
nor U1396 (N_1396,N_1247,N_1267);
xor U1397 (N_1397,N_1294,N_1248);
or U1398 (N_1398,N_1253,N_1274);
nand U1399 (N_1399,N_1290,N_1227);
nand U1400 (N_1400,N_1336,N_1320);
nand U1401 (N_1401,N_1354,N_1396);
nor U1402 (N_1402,N_1344,N_1398);
and U1403 (N_1403,N_1345,N_1399);
xnor U1404 (N_1404,N_1316,N_1348);
nand U1405 (N_1405,N_1341,N_1352);
nand U1406 (N_1406,N_1379,N_1304);
xnor U1407 (N_1407,N_1378,N_1327);
nor U1408 (N_1408,N_1363,N_1333);
or U1409 (N_1409,N_1387,N_1315);
and U1410 (N_1410,N_1312,N_1305);
and U1411 (N_1411,N_1369,N_1380);
or U1412 (N_1412,N_1343,N_1306);
or U1413 (N_1413,N_1335,N_1361);
nor U1414 (N_1414,N_1368,N_1323);
nor U1415 (N_1415,N_1397,N_1371);
xnor U1416 (N_1416,N_1375,N_1374);
or U1417 (N_1417,N_1339,N_1365);
nor U1418 (N_1418,N_1337,N_1347);
xnor U1419 (N_1419,N_1389,N_1364);
nand U1420 (N_1420,N_1394,N_1351);
and U1421 (N_1421,N_1311,N_1388);
and U1422 (N_1422,N_1366,N_1362);
nor U1423 (N_1423,N_1360,N_1303);
or U1424 (N_1424,N_1330,N_1308);
and U1425 (N_1425,N_1307,N_1340);
nor U1426 (N_1426,N_1346,N_1310);
xnor U1427 (N_1427,N_1317,N_1372);
and U1428 (N_1428,N_1353,N_1301);
xor U1429 (N_1429,N_1329,N_1314);
and U1430 (N_1430,N_1332,N_1350);
or U1431 (N_1431,N_1391,N_1390);
nor U1432 (N_1432,N_1358,N_1325);
and U1433 (N_1433,N_1300,N_1370);
nor U1434 (N_1434,N_1393,N_1331);
nand U1435 (N_1435,N_1313,N_1318);
nand U1436 (N_1436,N_1384,N_1355);
xnor U1437 (N_1437,N_1334,N_1302);
nand U1438 (N_1438,N_1357,N_1367);
and U1439 (N_1439,N_1338,N_1342);
nand U1440 (N_1440,N_1383,N_1373);
and U1441 (N_1441,N_1328,N_1359);
and U1442 (N_1442,N_1309,N_1356);
and U1443 (N_1443,N_1377,N_1385);
nand U1444 (N_1444,N_1319,N_1322);
xnor U1445 (N_1445,N_1381,N_1382);
nor U1446 (N_1446,N_1392,N_1349);
and U1447 (N_1447,N_1376,N_1386);
xor U1448 (N_1448,N_1321,N_1395);
nand U1449 (N_1449,N_1326,N_1324);
nor U1450 (N_1450,N_1368,N_1366);
and U1451 (N_1451,N_1357,N_1355);
xor U1452 (N_1452,N_1391,N_1345);
xor U1453 (N_1453,N_1338,N_1391);
xnor U1454 (N_1454,N_1353,N_1358);
nor U1455 (N_1455,N_1376,N_1394);
or U1456 (N_1456,N_1395,N_1359);
nand U1457 (N_1457,N_1391,N_1394);
and U1458 (N_1458,N_1314,N_1363);
xor U1459 (N_1459,N_1325,N_1336);
nor U1460 (N_1460,N_1338,N_1354);
or U1461 (N_1461,N_1336,N_1300);
and U1462 (N_1462,N_1387,N_1332);
xnor U1463 (N_1463,N_1317,N_1341);
or U1464 (N_1464,N_1362,N_1307);
nor U1465 (N_1465,N_1300,N_1369);
nand U1466 (N_1466,N_1314,N_1398);
nand U1467 (N_1467,N_1322,N_1389);
nor U1468 (N_1468,N_1308,N_1317);
xnor U1469 (N_1469,N_1385,N_1327);
xnor U1470 (N_1470,N_1305,N_1398);
or U1471 (N_1471,N_1370,N_1388);
nand U1472 (N_1472,N_1396,N_1371);
or U1473 (N_1473,N_1366,N_1315);
and U1474 (N_1474,N_1388,N_1377);
nor U1475 (N_1475,N_1356,N_1338);
or U1476 (N_1476,N_1331,N_1309);
nand U1477 (N_1477,N_1311,N_1385);
or U1478 (N_1478,N_1375,N_1337);
xor U1479 (N_1479,N_1380,N_1323);
nor U1480 (N_1480,N_1337,N_1346);
nor U1481 (N_1481,N_1323,N_1334);
nor U1482 (N_1482,N_1326,N_1302);
or U1483 (N_1483,N_1396,N_1328);
or U1484 (N_1484,N_1361,N_1357);
nand U1485 (N_1485,N_1318,N_1322);
and U1486 (N_1486,N_1305,N_1320);
nor U1487 (N_1487,N_1397,N_1356);
or U1488 (N_1488,N_1331,N_1398);
nand U1489 (N_1489,N_1302,N_1392);
or U1490 (N_1490,N_1319,N_1382);
xor U1491 (N_1491,N_1329,N_1379);
or U1492 (N_1492,N_1345,N_1383);
nand U1493 (N_1493,N_1388,N_1379);
or U1494 (N_1494,N_1399,N_1317);
nand U1495 (N_1495,N_1384,N_1304);
xor U1496 (N_1496,N_1344,N_1347);
xor U1497 (N_1497,N_1301,N_1321);
xor U1498 (N_1498,N_1343,N_1370);
nor U1499 (N_1499,N_1371,N_1352);
nor U1500 (N_1500,N_1444,N_1467);
nor U1501 (N_1501,N_1468,N_1465);
and U1502 (N_1502,N_1482,N_1421);
or U1503 (N_1503,N_1457,N_1407);
and U1504 (N_1504,N_1486,N_1425);
and U1505 (N_1505,N_1454,N_1474);
or U1506 (N_1506,N_1430,N_1475);
nand U1507 (N_1507,N_1406,N_1404);
nor U1508 (N_1508,N_1495,N_1451);
nor U1509 (N_1509,N_1402,N_1471);
nor U1510 (N_1510,N_1490,N_1423);
and U1511 (N_1511,N_1401,N_1461);
nand U1512 (N_1512,N_1462,N_1440);
and U1513 (N_1513,N_1493,N_1408);
or U1514 (N_1514,N_1428,N_1481);
nand U1515 (N_1515,N_1419,N_1459);
or U1516 (N_1516,N_1400,N_1420);
and U1517 (N_1517,N_1417,N_1448);
nand U1518 (N_1518,N_1443,N_1405);
or U1519 (N_1519,N_1470,N_1447);
nor U1520 (N_1520,N_1441,N_1410);
xor U1521 (N_1521,N_1450,N_1445);
or U1522 (N_1522,N_1464,N_1496);
or U1523 (N_1523,N_1424,N_1427);
or U1524 (N_1524,N_1458,N_1411);
nor U1525 (N_1525,N_1416,N_1479);
and U1526 (N_1526,N_1491,N_1469);
or U1527 (N_1527,N_1484,N_1435);
nand U1528 (N_1528,N_1466,N_1473);
xor U1529 (N_1529,N_1485,N_1455);
or U1530 (N_1530,N_1472,N_1442);
xnor U1531 (N_1531,N_1437,N_1438);
nand U1532 (N_1532,N_1476,N_1414);
nor U1533 (N_1533,N_1432,N_1460);
or U1534 (N_1534,N_1480,N_1412);
nand U1535 (N_1535,N_1453,N_1494);
or U1536 (N_1536,N_1498,N_1433);
nand U1537 (N_1537,N_1456,N_1487);
xor U1538 (N_1538,N_1489,N_1499);
xor U1539 (N_1539,N_1418,N_1409);
nor U1540 (N_1540,N_1413,N_1429);
and U1541 (N_1541,N_1422,N_1436);
and U1542 (N_1542,N_1452,N_1431);
and U1543 (N_1543,N_1463,N_1415);
and U1544 (N_1544,N_1446,N_1477);
nand U1545 (N_1545,N_1403,N_1434);
nand U1546 (N_1546,N_1439,N_1426);
or U1547 (N_1547,N_1478,N_1449);
nand U1548 (N_1548,N_1483,N_1488);
and U1549 (N_1549,N_1492,N_1497);
and U1550 (N_1550,N_1407,N_1416);
nor U1551 (N_1551,N_1496,N_1449);
nand U1552 (N_1552,N_1481,N_1461);
xnor U1553 (N_1553,N_1455,N_1437);
nand U1554 (N_1554,N_1427,N_1421);
xor U1555 (N_1555,N_1484,N_1450);
xnor U1556 (N_1556,N_1469,N_1480);
and U1557 (N_1557,N_1453,N_1417);
nor U1558 (N_1558,N_1404,N_1493);
xnor U1559 (N_1559,N_1415,N_1492);
nand U1560 (N_1560,N_1488,N_1415);
nor U1561 (N_1561,N_1405,N_1479);
xnor U1562 (N_1562,N_1401,N_1481);
and U1563 (N_1563,N_1427,N_1451);
nand U1564 (N_1564,N_1437,N_1414);
and U1565 (N_1565,N_1448,N_1445);
and U1566 (N_1566,N_1415,N_1413);
nand U1567 (N_1567,N_1413,N_1476);
and U1568 (N_1568,N_1414,N_1484);
xnor U1569 (N_1569,N_1443,N_1467);
and U1570 (N_1570,N_1462,N_1474);
xnor U1571 (N_1571,N_1408,N_1448);
nand U1572 (N_1572,N_1403,N_1471);
xnor U1573 (N_1573,N_1498,N_1493);
xor U1574 (N_1574,N_1424,N_1481);
nand U1575 (N_1575,N_1443,N_1496);
and U1576 (N_1576,N_1424,N_1439);
nor U1577 (N_1577,N_1465,N_1433);
xor U1578 (N_1578,N_1466,N_1411);
or U1579 (N_1579,N_1454,N_1436);
nor U1580 (N_1580,N_1461,N_1428);
nor U1581 (N_1581,N_1473,N_1430);
and U1582 (N_1582,N_1420,N_1495);
nor U1583 (N_1583,N_1481,N_1449);
nand U1584 (N_1584,N_1490,N_1420);
nor U1585 (N_1585,N_1489,N_1457);
xnor U1586 (N_1586,N_1413,N_1463);
and U1587 (N_1587,N_1424,N_1429);
nor U1588 (N_1588,N_1438,N_1427);
xor U1589 (N_1589,N_1435,N_1406);
xor U1590 (N_1590,N_1408,N_1422);
or U1591 (N_1591,N_1444,N_1491);
or U1592 (N_1592,N_1414,N_1491);
nand U1593 (N_1593,N_1448,N_1493);
nand U1594 (N_1594,N_1484,N_1443);
and U1595 (N_1595,N_1430,N_1436);
nor U1596 (N_1596,N_1486,N_1407);
xnor U1597 (N_1597,N_1467,N_1451);
or U1598 (N_1598,N_1453,N_1491);
nor U1599 (N_1599,N_1479,N_1453);
and U1600 (N_1600,N_1511,N_1589);
xnor U1601 (N_1601,N_1572,N_1599);
or U1602 (N_1602,N_1578,N_1512);
nor U1603 (N_1603,N_1588,N_1574);
nor U1604 (N_1604,N_1500,N_1555);
and U1605 (N_1605,N_1590,N_1543);
or U1606 (N_1606,N_1584,N_1570);
and U1607 (N_1607,N_1529,N_1517);
nor U1608 (N_1608,N_1596,N_1550);
nand U1609 (N_1609,N_1553,N_1575);
and U1610 (N_1610,N_1506,N_1577);
or U1611 (N_1611,N_1546,N_1554);
and U1612 (N_1612,N_1597,N_1576);
nand U1613 (N_1613,N_1547,N_1592);
or U1614 (N_1614,N_1501,N_1504);
and U1615 (N_1615,N_1524,N_1552);
and U1616 (N_1616,N_1551,N_1549);
and U1617 (N_1617,N_1558,N_1523);
nor U1618 (N_1618,N_1594,N_1525);
or U1619 (N_1619,N_1568,N_1538);
nand U1620 (N_1620,N_1545,N_1527);
and U1621 (N_1621,N_1531,N_1565);
and U1622 (N_1622,N_1564,N_1593);
nand U1623 (N_1623,N_1528,N_1518);
nor U1624 (N_1624,N_1520,N_1513);
nor U1625 (N_1625,N_1522,N_1548);
nand U1626 (N_1626,N_1583,N_1539);
or U1627 (N_1627,N_1566,N_1580);
xor U1628 (N_1628,N_1562,N_1585);
and U1629 (N_1629,N_1557,N_1509);
and U1630 (N_1630,N_1507,N_1541);
or U1631 (N_1631,N_1586,N_1530);
and U1632 (N_1632,N_1540,N_1508);
or U1633 (N_1633,N_1563,N_1502);
and U1634 (N_1634,N_1514,N_1559);
nor U1635 (N_1635,N_1567,N_1534);
xnor U1636 (N_1636,N_1560,N_1544);
or U1637 (N_1637,N_1515,N_1526);
nor U1638 (N_1638,N_1571,N_1569);
and U1639 (N_1639,N_1595,N_1537);
and U1640 (N_1640,N_1536,N_1533);
nor U1641 (N_1641,N_1503,N_1591);
nor U1642 (N_1642,N_1510,N_1561);
or U1643 (N_1643,N_1535,N_1521);
and U1644 (N_1644,N_1582,N_1519);
nand U1645 (N_1645,N_1587,N_1532);
and U1646 (N_1646,N_1598,N_1505);
nor U1647 (N_1647,N_1579,N_1516);
nor U1648 (N_1648,N_1556,N_1573);
nor U1649 (N_1649,N_1542,N_1581);
nand U1650 (N_1650,N_1584,N_1599);
nand U1651 (N_1651,N_1505,N_1549);
or U1652 (N_1652,N_1503,N_1516);
nor U1653 (N_1653,N_1522,N_1521);
and U1654 (N_1654,N_1591,N_1568);
xor U1655 (N_1655,N_1587,N_1521);
xor U1656 (N_1656,N_1598,N_1542);
or U1657 (N_1657,N_1575,N_1572);
or U1658 (N_1658,N_1574,N_1502);
or U1659 (N_1659,N_1591,N_1544);
nor U1660 (N_1660,N_1508,N_1524);
xnor U1661 (N_1661,N_1545,N_1546);
xor U1662 (N_1662,N_1551,N_1541);
xnor U1663 (N_1663,N_1528,N_1522);
nand U1664 (N_1664,N_1548,N_1547);
or U1665 (N_1665,N_1539,N_1551);
xor U1666 (N_1666,N_1502,N_1586);
nor U1667 (N_1667,N_1549,N_1573);
or U1668 (N_1668,N_1573,N_1531);
xor U1669 (N_1669,N_1554,N_1591);
or U1670 (N_1670,N_1558,N_1542);
or U1671 (N_1671,N_1546,N_1516);
and U1672 (N_1672,N_1555,N_1575);
or U1673 (N_1673,N_1518,N_1524);
or U1674 (N_1674,N_1580,N_1524);
xor U1675 (N_1675,N_1529,N_1587);
or U1676 (N_1676,N_1567,N_1500);
xor U1677 (N_1677,N_1575,N_1550);
and U1678 (N_1678,N_1580,N_1505);
and U1679 (N_1679,N_1595,N_1552);
nand U1680 (N_1680,N_1582,N_1512);
nand U1681 (N_1681,N_1567,N_1515);
nor U1682 (N_1682,N_1553,N_1572);
and U1683 (N_1683,N_1593,N_1541);
nand U1684 (N_1684,N_1539,N_1582);
nand U1685 (N_1685,N_1526,N_1520);
nor U1686 (N_1686,N_1504,N_1577);
nand U1687 (N_1687,N_1516,N_1584);
or U1688 (N_1688,N_1598,N_1516);
and U1689 (N_1689,N_1507,N_1596);
or U1690 (N_1690,N_1515,N_1560);
or U1691 (N_1691,N_1542,N_1572);
and U1692 (N_1692,N_1536,N_1592);
nor U1693 (N_1693,N_1592,N_1576);
nor U1694 (N_1694,N_1503,N_1574);
or U1695 (N_1695,N_1564,N_1543);
and U1696 (N_1696,N_1561,N_1511);
nand U1697 (N_1697,N_1548,N_1557);
and U1698 (N_1698,N_1556,N_1584);
and U1699 (N_1699,N_1513,N_1568);
xor U1700 (N_1700,N_1613,N_1683);
nor U1701 (N_1701,N_1644,N_1620);
xor U1702 (N_1702,N_1604,N_1649);
xnor U1703 (N_1703,N_1660,N_1680);
and U1704 (N_1704,N_1616,N_1623);
or U1705 (N_1705,N_1691,N_1668);
nor U1706 (N_1706,N_1642,N_1614);
nor U1707 (N_1707,N_1694,N_1619);
or U1708 (N_1708,N_1600,N_1607);
or U1709 (N_1709,N_1622,N_1676);
nand U1710 (N_1710,N_1658,N_1646);
nand U1711 (N_1711,N_1678,N_1684);
nand U1712 (N_1712,N_1661,N_1654);
or U1713 (N_1713,N_1698,N_1672);
or U1714 (N_1714,N_1629,N_1695);
xnor U1715 (N_1715,N_1628,N_1652);
nand U1716 (N_1716,N_1690,N_1630);
xor U1717 (N_1717,N_1692,N_1674);
and U1718 (N_1718,N_1625,N_1665);
and U1719 (N_1719,N_1627,N_1631);
nor U1720 (N_1720,N_1656,N_1643);
and U1721 (N_1721,N_1697,N_1603);
xor U1722 (N_1722,N_1610,N_1602);
nand U1723 (N_1723,N_1662,N_1645);
xor U1724 (N_1724,N_1673,N_1618);
nor U1725 (N_1725,N_1696,N_1677);
nand U1726 (N_1726,N_1653,N_1638);
or U1727 (N_1727,N_1659,N_1617);
and U1728 (N_1728,N_1669,N_1647);
or U1729 (N_1729,N_1637,N_1611);
and U1730 (N_1730,N_1626,N_1687);
or U1731 (N_1731,N_1666,N_1624);
nand U1732 (N_1732,N_1675,N_1679);
nor U1733 (N_1733,N_1615,N_1664);
nand U1734 (N_1734,N_1667,N_1686);
nor U1735 (N_1735,N_1670,N_1641);
xnor U1736 (N_1736,N_1655,N_1699);
xnor U1737 (N_1737,N_1601,N_1606);
nand U1738 (N_1738,N_1657,N_1632);
or U1739 (N_1739,N_1639,N_1608);
nor U1740 (N_1740,N_1636,N_1640);
nor U1741 (N_1741,N_1621,N_1685);
or U1742 (N_1742,N_1650,N_1671);
nand U1743 (N_1743,N_1651,N_1648);
and U1744 (N_1744,N_1693,N_1605);
or U1745 (N_1745,N_1634,N_1681);
nand U1746 (N_1746,N_1663,N_1612);
nor U1747 (N_1747,N_1635,N_1688);
and U1748 (N_1748,N_1633,N_1682);
and U1749 (N_1749,N_1609,N_1689);
nor U1750 (N_1750,N_1615,N_1602);
and U1751 (N_1751,N_1648,N_1604);
nand U1752 (N_1752,N_1682,N_1655);
and U1753 (N_1753,N_1678,N_1616);
xor U1754 (N_1754,N_1635,N_1673);
nand U1755 (N_1755,N_1692,N_1650);
nand U1756 (N_1756,N_1646,N_1629);
nor U1757 (N_1757,N_1688,N_1698);
or U1758 (N_1758,N_1677,N_1687);
or U1759 (N_1759,N_1600,N_1651);
nand U1760 (N_1760,N_1612,N_1625);
nor U1761 (N_1761,N_1624,N_1625);
and U1762 (N_1762,N_1651,N_1640);
and U1763 (N_1763,N_1648,N_1621);
xnor U1764 (N_1764,N_1699,N_1683);
nand U1765 (N_1765,N_1667,N_1651);
or U1766 (N_1766,N_1660,N_1661);
nor U1767 (N_1767,N_1637,N_1668);
xnor U1768 (N_1768,N_1608,N_1651);
nand U1769 (N_1769,N_1685,N_1604);
and U1770 (N_1770,N_1676,N_1689);
nor U1771 (N_1771,N_1632,N_1677);
nor U1772 (N_1772,N_1647,N_1691);
nand U1773 (N_1773,N_1668,N_1605);
nand U1774 (N_1774,N_1667,N_1623);
nand U1775 (N_1775,N_1651,N_1693);
xor U1776 (N_1776,N_1669,N_1691);
and U1777 (N_1777,N_1618,N_1614);
and U1778 (N_1778,N_1666,N_1601);
nor U1779 (N_1779,N_1608,N_1653);
nand U1780 (N_1780,N_1638,N_1625);
xor U1781 (N_1781,N_1680,N_1625);
nand U1782 (N_1782,N_1626,N_1610);
and U1783 (N_1783,N_1642,N_1604);
nand U1784 (N_1784,N_1642,N_1693);
xnor U1785 (N_1785,N_1623,N_1666);
and U1786 (N_1786,N_1635,N_1627);
or U1787 (N_1787,N_1669,N_1605);
nand U1788 (N_1788,N_1632,N_1603);
and U1789 (N_1789,N_1617,N_1600);
nand U1790 (N_1790,N_1655,N_1609);
or U1791 (N_1791,N_1603,N_1627);
nor U1792 (N_1792,N_1629,N_1606);
or U1793 (N_1793,N_1672,N_1649);
xnor U1794 (N_1794,N_1633,N_1668);
or U1795 (N_1795,N_1604,N_1601);
and U1796 (N_1796,N_1677,N_1635);
and U1797 (N_1797,N_1665,N_1677);
or U1798 (N_1798,N_1627,N_1658);
xnor U1799 (N_1799,N_1606,N_1607);
nand U1800 (N_1800,N_1740,N_1721);
nor U1801 (N_1801,N_1774,N_1769);
nand U1802 (N_1802,N_1795,N_1754);
and U1803 (N_1803,N_1756,N_1718);
nand U1804 (N_1804,N_1724,N_1758);
nand U1805 (N_1805,N_1737,N_1750);
or U1806 (N_1806,N_1765,N_1705);
and U1807 (N_1807,N_1766,N_1785);
and U1808 (N_1808,N_1796,N_1728);
or U1809 (N_1809,N_1798,N_1727);
nor U1810 (N_1810,N_1794,N_1744);
or U1811 (N_1811,N_1784,N_1771);
nor U1812 (N_1812,N_1764,N_1745);
and U1813 (N_1813,N_1753,N_1770);
nor U1814 (N_1814,N_1702,N_1760);
or U1815 (N_1815,N_1713,N_1786);
and U1816 (N_1816,N_1719,N_1735);
xor U1817 (N_1817,N_1736,N_1788);
or U1818 (N_1818,N_1781,N_1720);
nand U1819 (N_1819,N_1777,N_1779);
nand U1820 (N_1820,N_1775,N_1704);
nor U1821 (N_1821,N_1717,N_1749);
and U1822 (N_1822,N_1793,N_1710);
nor U1823 (N_1823,N_1700,N_1755);
nand U1824 (N_1824,N_1741,N_1759);
xnor U1825 (N_1825,N_1733,N_1787);
nor U1826 (N_1826,N_1731,N_1712);
or U1827 (N_1827,N_1791,N_1751);
or U1828 (N_1828,N_1776,N_1761);
nand U1829 (N_1829,N_1742,N_1701);
or U1830 (N_1830,N_1734,N_1747);
and U1831 (N_1831,N_1783,N_1797);
and U1832 (N_1832,N_1738,N_1768);
xnor U1833 (N_1833,N_1709,N_1739);
or U1834 (N_1834,N_1790,N_1752);
nand U1835 (N_1835,N_1715,N_1792);
and U1836 (N_1836,N_1743,N_1714);
and U1837 (N_1837,N_1716,N_1748);
xor U1838 (N_1838,N_1703,N_1762);
xor U1839 (N_1839,N_1723,N_1726);
or U1840 (N_1840,N_1778,N_1725);
and U1841 (N_1841,N_1746,N_1732);
nand U1842 (N_1842,N_1757,N_1708);
or U1843 (N_1843,N_1711,N_1729);
and U1844 (N_1844,N_1782,N_1722);
xor U1845 (N_1845,N_1789,N_1780);
or U1846 (N_1846,N_1763,N_1707);
xor U1847 (N_1847,N_1772,N_1730);
nor U1848 (N_1848,N_1773,N_1767);
and U1849 (N_1849,N_1799,N_1706);
xnor U1850 (N_1850,N_1754,N_1702);
xor U1851 (N_1851,N_1739,N_1707);
nor U1852 (N_1852,N_1759,N_1722);
nand U1853 (N_1853,N_1765,N_1735);
or U1854 (N_1854,N_1753,N_1714);
nand U1855 (N_1855,N_1741,N_1782);
nand U1856 (N_1856,N_1755,N_1759);
xnor U1857 (N_1857,N_1773,N_1717);
nor U1858 (N_1858,N_1700,N_1754);
or U1859 (N_1859,N_1759,N_1707);
nor U1860 (N_1860,N_1704,N_1760);
nor U1861 (N_1861,N_1793,N_1776);
and U1862 (N_1862,N_1789,N_1709);
or U1863 (N_1863,N_1759,N_1782);
nor U1864 (N_1864,N_1763,N_1701);
nor U1865 (N_1865,N_1749,N_1727);
and U1866 (N_1866,N_1725,N_1789);
or U1867 (N_1867,N_1756,N_1720);
nor U1868 (N_1868,N_1779,N_1769);
nand U1869 (N_1869,N_1724,N_1736);
or U1870 (N_1870,N_1729,N_1753);
nor U1871 (N_1871,N_1703,N_1720);
nand U1872 (N_1872,N_1788,N_1756);
xnor U1873 (N_1873,N_1741,N_1704);
nor U1874 (N_1874,N_1776,N_1766);
nand U1875 (N_1875,N_1722,N_1747);
nand U1876 (N_1876,N_1764,N_1740);
or U1877 (N_1877,N_1760,N_1758);
xor U1878 (N_1878,N_1735,N_1713);
and U1879 (N_1879,N_1724,N_1749);
nor U1880 (N_1880,N_1795,N_1727);
xnor U1881 (N_1881,N_1755,N_1750);
xnor U1882 (N_1882,N_1798,N_1799);
or U1883 (N_1883,N_1712,N_1786);
nand U1884 (N_1884,N_1783,N_1704);
or U1885 (N_1885,N_1742,N_1731);
nand U1886 (N_1886,N_1726,N_1705);
xnor U1887 (N_1887,N_1799,N_1784);
nand U1888 (N_1888,N_1707,N_1740);
nor U1889 (N_1889,N_1789,N_1716);
or U1890 (N_1890,N_1708,N_1739);
and U1891 (N_1891,N_1769,N_1770);
or U1892 (N_1892,N_1765,N_1741);
xnor U1893 (N_1893,N_1799,N_1732);
xor U1894 (N_1894,N_1784,N_1758);
nand U1895 (N_1895,N_1727,N_1702);
nand U1896 (N_1896,N_1760,N_1756);
or U1897 (N_1897,N_1748,N_1767);
xnor U1898 (N_1898,N_1710,N_1749);
nor U1899 (N_1899,N_1745,N_1783);
or U1900 (N_1900,N_1828,N_1886);
nor U1901 (N_1901,N_1860,N_1858);
nor U1902 (N_1902,N_1809,N_1829);
nand U1903 (N_1903,N_1861,N_1887);
nand U1904 (N_1904,N_1875,N_1897);
and U1905 (N_1905,N_1814,N_1880);
nor U1906 (N_1906,N_1836,N_1841);
nand U1907 (N_1907,N_1800,N_1805);
and U1908 (N_1908,N_1889,N_1852);
and U1909 (N_1909,N_1826,N_1885);
xor U1910 (N_1910,N_1899,N_1878);
or U1911 (N_1911,N_1865,N_1874);
nor U1912 (N_1912,N_1862,N_1830);
nand U1913 (N_1913,N_1891,N_1843);
nor U1914 (N_1914,N_1844,N_1871);
nor U1915 (N_1915,N_1835,N_1842);
nor U1916 (N_1916,N_1833,N_1882);
or U1917 (N_1917,N_1846,N_1866);
nand U1918 (N_1918,N_1831,N_1847);
or U1919 (N_1919,N_1898,N_1817);
nand U1920 (N_1920,N_1822,N_1881);
xor U1921 (N_1921,N_1839,N_1893);
xor U1922 (N_1922,N_1832,N_1803);
nor U1923 (N_1923,N_1857,N_1851);
nor U1924 (N_1924,N_1868,N_1876);
xnor U1925 (N_1925,N_1834,N_1894);
and U1926 (N_1926,N_1849,N_1872);
nand U1927 (N_1927,N_1838,N_1824);
nand U1928 (N_1928,N_1816,N_1890);
and U1929 (N_1929,N_1879,N_1810);
and U1930 (N_1930,N_1856,N_1845);
or U1931 (N_1931,N_1820,N_1821);
nor U1932 (N_1932,N_1873,N_1807);
xor U1933 (N_1933,N_1837,N_1853);
xnor U1934 (N_1934,N_1801,N_1825);
and U1935 (N_1935,N_1808,N_1892);
or U1936 (N_1936,N_1813,N_1823);
xor U1937 (N_1937,N_1883,N_1896);
or U1938 (N_1938,N_1848,N_1863);
or U1939 (N_1939,N_1804,N_1840);
nand U1940 (N_1940,N_1811,N_1895);
nor U1941 (N_1941,N_1869,N_1864);
nand U1942 (N_1942,N_1859,N_1888);
nor U1943 (N_1943,N_1877,N_1819);
and U1944 (N_1944,N_1850,N_1815);
and U1945 (N_1945,N_1806,N_1818);
nand U1946 (N_1946,N_1812,N_1802);
nand U1947 (N_1947,N_1855,N_1870);
or U1948 (N_1948,N_1867,N_1854);
xor U1949 (N_1949,N_1827,N_1884);
nor U1950 (N_1950,N_1843,N_1886);
nand U1951 (N_1951,N_1861,N_1822);
nor U1952 (N_1952,N_1899,N_1806);
and U1953 (N_1953,N_1851,N_1892);
xor U1954 (N_1954,N_1814,N_1891);
or U1955 (N_1955,N_1832,N_1893);
or U1956 (N_1956,N_1808,N_1800);
nor U1957 (N_1957,N_1824,N_1847);
nor U1958 (N_1958,N_1847,N_1834);
or U1959 (N_1959,N_1874,N_1882);
and U1960 (N_1960,N_1890,N_1805);
xor U1961 (N_1961,N_1880,N_1898);
nand U1962 (N_1962,N_1820,N_1835);
nor U1963 (N_1963,N_1822,N_1826);
nand U1964 (N_1964,N_1872,N_1892);
nand U1965 (N_1965,N_1827,N_1886);
nand U1966 (N_1966,N_1894,N_1857);
or U1967 (N_1967,N_1887,N_1806);
or U1968 (N_1968,N_1897,N_1830);
and U1969 (N_1969,N_1824,N_1820);
and U1970 (N_1970,N_1861,N_1831);
nor U1971 (N_1971,N_1846,N_1822);
xor U1972 (N_1972,N_1842,N_1824);
nand U1973 (N_1973,N_1840,N_1812);
xnor U1974 (N_1974,N_1884,N_1829);
xor U1975 (N_1975,N_1876,N_1814);
or U1976 (N_1976,N_1817,N_1838);
xnor U1977 (N_1977,N_1898,N_1862);
xnor U1978 (N_1978,N_1842,N_1820);
nand U1979 (N_1979,N_1855,N_1875);
nand U1980 (N_1980,N_1845,N_1839);
xnor U1981 (N_1981,N_1884,N_1810);
nand U1982 (N_1982,N_1828,N_1842);
nand U1983 (N_1983,N_1826,N_1859);
xnor U1984 (N_1984,N_1870,N_1878);
or U1985 (N_1985,N_1856,N_1874);
and U1986 (N_1986,N_1818,N_1878);
or U1987 (N_1987,N_1800,N_1876);
or U1988 (N_1988,N_1855,N_1839);
or U1989 (N_1989,N_1877,N_1817);
or U1990 (N_1990,N_1866,N_1833);
xnor U1991 (N_1991,N_1822,N_1890);
nor U1992 (N_1992,N_1852,N_1805);
and U1993 (N_1993,N_1895,N_1864);
xnor U1994 (N_1994,N_1803,N_1858);
nand U1995 (N_1995,N_1832,N_1838);
or U1996 (N_1996,N_1853,N_1863);
nor U1997 (N_1997,N_1893,N_1858);
nand U1998 (N_1998,N_1870,N_1839);
or U1999 (N_1999,N_1827,N_1806);
and U2000 (N_2000,N_1912,N_1966);
nand U2001 (N_2001,N_1929,N_1924);
nand U2002 (N_2002,N_1986,N_1948);
nor U2003 (N_2003,N_1920,N_1991);
and U2004 (N_2004,N_1968,N_1916);
nor U2005 (N_2005,N_1970,N_1983);
nand U2006 (N_2006,N_1909,N_1995);
xor U2007 (N_2007,N_1939,N_1935);
and U2008 (N_2008,N_1954,N_1959);
nand U2009 (N_2009,N_1907,N_1947);
nor U2010 (N_2010,N_1952,N_1942);
xnor U2011 (N_2011,N_1904,N_1993);
nand U2012 (N_2012,N_1963,N_1956);
or U2013 (N_2013,N_1902,N_1931);
xnor U2014 (N_2014,N_1928,N_1925);
or U2015 (N_2015,N_1994,N_1955);
nor U2016 (N_2016,N_1914,N_1944);
nor U2017 (N_2017,N_1978,N_1974);
xnor U2018 (N_2018,N_1953,N_1972);
nor U2019 (N_2019,N_1915,N_1949);
and U2020 (N_2020,N_1982,N_1981);
nor U2021 (N_2021,N_1918,N_1961);
or U2022 (N_2022,N_1917,N_1997);
or U2023 (N_2023,N_1945,N_1927);
xnor U2024 (N_2024,N_1911,N_1937);
and U2025 (N_2025,N_1964,N_1932);
and U2026 (N_2026,N_1967,N_1969);
nand U2027 (N_2027,N_1976,N_1900);
and U2028 (N_2028,N_1975,N_1988);
nand U2029 (N_2029,N_1979,N_1951);
xor U2030 (N_2030,N_1987,N_1934);
and U2031 (N_2031,N_1940,N_1903);
or U2032 (N_2032,N_1990,N_1977);
xor U2033 (N_2033,N_1992,N_1960);
and U2034 (N_2034,N_1908,N_1973);
or U2035 (N_2035,N_1957,N_1980);
and U2036 (N_2036,N_1923,N_1921);
nand U2037 (N_2037,N_1933,N_1985);
xor U2038 (N_2038,N_1930,N_1905);
nand U2039 (N_2039,N_1910,N_1996);
and U2040 (N_2040,N_1962,N_1936);
nand U2041 (N_2041,N_1938,N_1971);
nand U2042 (N_2042,N_1958,N_1941);
xnor U2043 (N_2043,N_1946,N_1984);
nand U2044 (N_2044,N_1906,N_1999);
nor U2045 (N_2045,N_1965,N_1950);
nand U2046 (N_2046,N_1913,N_1943);
xor U2047 (N_2047,N_1926,N_1922);
nor U2048 (N_2048,N_1919,N_1989);
nand U2049 (N_2049,N_1998,N_1901);
nor U2050 (N_2050,N_1989,N_1955);
nor U2051 (N_2051,N_1979,N_1931);
and U2052 (N_2052,N_1929,N_1996);
nor U2053 (N_2053,N_1967,N_1909);
and U2054 (N_2054,N_1988,N_1973);
and U2055 (N_2055,N_1956,N_1974);
xor U2056 (N_2056,N_1941,N_1967);
nand U2057 (N_2057,N_1935,N_1969);
or U2058 (N_2058,N_1966,N_1977);
nand U2059 (N_2059,N_1998,N_1905);
nand U2060 (N_2060,N_1926,N_1925);
or U2061 (N_2061,N_1994,N_1928);
xor U2062 (N_2062,N_1961,N_1957);
or U2063 (N_2063,N_1974,N_1982);
xor U2064 (N_2064,N_1915,N_1935);
or U2065 (N_2065,N_1987,N_1954);
xnor U2066 (N_2066,N_1907,N_1915);
or U2067 (N_2067,N_1942,N_1930);
and U2068 (N_2068,N_1951,N_1946);
nand U2069 (N_2069,N_1950,N_1983);
and U2070 (N_2070,N_1973,N_1938);
nor U2071 (N_2071,N_1937,N_1976);
and U2072 (N_2072,N_1937,N_1939);
or U2073 (N_2073,N_1925,N_1936);
nor U2074 (N_2074,N_1960,N_1930);
and U2075 (N_2075,N_1918,N_1931);
or U2076 (N_2076,N_1906,N_1972);
nand U2077 (N_2077,N_1914,N_1933);
and U2078 (N_2078,N_1941,N_1912);
nor U2079 (N_2079,N_1944,N_1939);
or U2080 (N_2080,N_1917,N_1992);
and U2081 (N_2081,N_1931,N_1953);
or U2082 (N_2082,N_1993,N_1900);
xnor U2083 (N_2083,N_1949,N_1917);
nand U2084 (N_2084,N_1979,N_1915);
xor U2085 (N_2085,N_1973,N_1953);
nand U2086 (N_2086,N_1968,N_1951);
xor U2087 (N_2087,N_1943,N_1926);
nor U2088 (N_2088,N_1930,N_1997);
nor U2089 (N_2089,N_1963,N_1958);
or U2090 (N_2090,N_1946,N_1988);
or U2091 (N_2091,N_1995,N_1991);
nand U2092 (N_2092,N_1978,N_1915);
nand U2093 (N_2093,N_1928,N_1956);
nand U2094 (N_2094,N_1981,N_1916);
nor U2095 (N_2095,N_1945,N_1910);
and U2096 (N_2096,N_1936,N_1959);
xor U2097 (N_2097,N_1926,N_1997);
nor U2098 (N_2098,N_1985,N_1919);
nand U2099 (N_2099,N_1974,N_1977);
or U2100 (N_2100,N_2097,N_2049);
nand U2101 (N_2101,N_2074,N_2098);
xor U2102 (N_2102,N_2051,N_2055);
xnor U2103 (N_2103,N_2068,N_2048);
or U2104 (N_2104,N_2053,N_2042);
or U2105 (N_2105,N_2096,N_2092);
nor U2106 (N_2106,N_2031,N_2082);
and U2107 (N_2107,N_2009,N_2020);
or U2108 (N_2108,N_2046,N_2043);
nor U2109 (N_2109,N_2070,N_2095);
nor U2110 (N_2110,N_2091,N_2035);
xor U2111 (N_2111,N_2027,N_2099);
or U2112 (N_2112,N_2015,N_2047);
xor U2113 (N_2113,N_2073,N_2085);
or U2114 (N_2114,N_2018,N_2083);
nand U2115 (N_2115,N_2034,N_2078);
nor U2116 (N_2116,N_2054,N_2038);
nand U2117 (N_2117,N_2025,N_2029);
or U2118 (N_2118,N_2003,N_2081);
and U2119 (N_2119,N_2011,N_2077);
or U2120 (N_2120,N_2013,N_2044);
nand U2121 (N_2121,N_2017,N_2021);
nand U2122 (N_2122,N_2024,N_2030);
and U2123 (N_2123,N_2080,N_2069);
or U2124 (N_2124,N_2041,N_2088);
xor U2125 (N_2125,N_2045,N_2076);
xor U2126 (N_2126,N_2007,N_2010);
nor U2127 (N_2127,N_2059,N_2000);
or U2128 (N_2128,N_2057,N_2093);
and U2129 (N_2129,N_2062,N_2002);
or U2130 (N_2130,N_2016,N_2089);
nor U2131 (N_2131,N_2075,N_2004);
and U2132 (N_2132,N_2061,N_2040);
and U2133 (N_2133,N_2052,N_2028);
and U2134 (N_2134,N_2033,N_2063);
xnor U2135 (N_2135,N_2023,N_2090);
or U2136 (N_2136,N_2094,N_2008);
nand U2137 (N_2137,N_2079,N_2056);
and U2138 (N_2138,N_2037,N_2058);
nor U2139 (N_2139,N_2084,N_2066);
nor U2140 (N_2140,N_2022,N_2006);
xnor U2141 (N_2141,N_2065,N_2019);
nand U2142 (N_2142,N_2036,N_2032);
or U2143 (N_2143,N_2039,N_2087);
or U2144 (N_2144,N_2005,N_2001);
or U2145 (N_2145,N_2067,N_2071);
xnor U2146 (N_2146,N_2060,N_2012);
and U2147 (N_2147,N_2050,N_2086);
and U2148 (N_2148,N_2026,N_2072);
xor U2149 (N_2149,N_2064,N_2014);
nand U2150 (N_2150,N_2044,N_2016);
nand U2151 (N_2151,N_2034,N_2046);
and U2152 (N_2152,N_2012,N_2077);
and U2153 (N_2153,N_2071,N_2020);
nor U2154 (N_2154,N_2019,N_2024);
or U2155 (N_2155,N_2055,N_2026);
and U2156 (N_2156,N_2061,N_2016);
nand U2157 (N_2157,N_2090,N_2052);
nor U2158 (N_2158,N_2093,N_2026);
nor U2159 (N_2159,N_2021,N_2040);
nand U2160 (N_2160,N_2042,N_2028);
and U2161 (N_2161,N_2082,N_2003);
nor U2162 (N_2162,N_2055,N_2020);
nand U2163 (N_2163,N_2039,N_2037);
and U2164 (N_2164,N_2063,N_2094);
or U2165 (N_2165,N_2097,N_2041);
and U2166 (N_2166,N_2090,N_2053);
and U2167 (N_2167,N_2081,N_2034);
and U2168 (N_2168,N_2012,N_2066);
nor U2169 (N_2169,N_2065,N_2009);
nor U2170 (N_2170,N_2051,N_2050);
and U2171 (N_2171,N_2062,N_2079);
and U2172 (N_2172,N_2072,N_2057);
nor U2173 (N_2173,N_2003,N_2073);
nor U2174 (N_2174,N_2004,N_2048);
and U2175 (N_2175,N_2061,N_2047);
nor U2176 (N_2176,N_2078,N_2061);
nor U2177 (N_2177,N_2099,N_2040);
nand U2178 (N_2178,N_2005,N_2046);
and U2179 (N_2179,N_2011,N_2003);
nor U2180 (N_2180,N_2065,N_2057);
nand U2181 (N_2181,N_2045,N_2084);
or U2182 (N_2182,N_2071,N_2059);
xor U2183 (N_2183,N_2061,N_2054);
and U2184 (N_2184,N_2054,N_2032);
xor U2185 (N_2185,N_2055,N_2045);
nor U2186 (N_2186,N_2068,N_2051);
xnor U2187 (N_2187,N_2015,N_2035);
and U2188 (N_2188,N_2082,N_2026);
and U2189 (N_2189,N_2012,N_2057);
or U2190 (N_2190,N_2047,N_2052);
nand U2191 (N_2191,N_2073,N_2030);
nor U2192 (N_2192,N_2082,N_2045);
xnor U2193 (N_2193,N_2064,N_2016);
nor U2194 (N_2194,N_2013,N_2097);
xnor U2195 (N_2195,N_2063,N_2057);
or U2196 (N_2196,N_2014,N_2073);
nand U2197 (N_2197,N_2036,N_2092);
or U2198 (N_2198,N_2005,N_2071);
nand U2199 (N_2199,N_2044,N_2057);
nand U2200 (N_2200,N_2102,N_2147);
and U2201 (N_2201,N_2166,N_2149);
and U2202 (N_2202,N_2183,N_2124);
xor U2203 (N_2203,N_2164,N_2119);
and U2204 (N_2204,N_2181,N_2118);
nand U2205 (N_2205,N_2155,N_2128);
nor U2206 (N_2206,N_2191,N_2100);
nor U2207 (N_2207,N_2123,N_2109);
nor U2208 (N_2208,N_2170,N_2111);
xnor U2209 (N_2209,N_2121,N_2135);
or U2210 (N_2210,N_2130,N_2112);
or U2211 (N_2211,N_2178,N_2104);
xnor U2212 (N_2212,N_2154,N_2197);
nand U2213 (N_2213,N_2159,N_2167);
xor U2214 (N_2214,N_2140,N_2169);
nor U2215 (N_2215,N_2176,N_2175);
xor U2216 (N_2216,N_2157,N_2165);
nand U2217 (N_2217,N_2150,N_2168);
nor U2218 (N_2218,N_2137,N_2132);
and U2219 (N_2219,N_2127,N_2145);
and U2220 (N_2220,N_2125,N_2171);
or U2221 (N_2221,N_2141,N_2122);
and U2222 (N_2222,N_2177,N_2129);
and U2223 (N_2223,N_2195,N_2103);
nor U2224 (N_2224,N_2180,N_2173);
and U2225 (N_2225,N_2110,N_2158);
nand U2226 (N_2226,N_2126,N_2192);
xnor U2227 (N_2227,N_2186,N_2163);
nor U2228 (N_2228,N_2189,N_2120);
nand U2229 (N_2229,N_2179,N_2146);
xor U2230 (N_2230,N_2142,N_2152);
nor U2231 (N_2231,N_2156,N_2106);
nor U2232 (N_2232,N_2144,N_2136);
nor U2233 (N_2233,N_2198,N_2182);
and U2234 (N_2234,N_2138,N_2114);
xnor U2235 (N_2235,N_2131,N_2185);
and U2236 (N_2236,N_2116,N_2105);
and U2237 (N_2237,N_2184,N_2113);
or U2238 (N_2238,N_2194,N_2196);
and U2239 (N_2239,N_2115,N_2133);
nand U2240 (N_2240,N_2134,N_2143);
or U2241 (N_2241,N_2160,N_2193);
xnor U2242 (N_2242,N_2162,N_2199);
xnor U2243 (N_2243,N_2188,N_2148);
nor U2244 (N_2244,N_2101,N_2108);
xnor U2245 (N_2245,N_2187,N_2174);
and U2246 (N_2246,N_2151,N_2107);
and U2247 (N_2247,N_2190,N_2139);
and U2248 (N_2248,N_2117,N_2172);
nand U2249 (N_2249,N_2153,N_2161);
xnor U2250 (N_2250,N_2195,N_2105);
or U2251 (N_2251,N_2137,N_2152);
nor U2252 (N_2252,N_2106,N_2113);
or U2253 (N_2253,N_2180,N_2185);
and U2254 (N_2254,N_2174,N_2138);
nor U2255 (N_2255,N_2186,N_2131);
and U2256 (N_2256,N_2180,N_2199);
xnor U2257 (N_2257,N_2160,N_2136);
nand U2258 (N_2258,N_2196,N_2113);
and U2259 (N_2259,N_2130,N_2183);
nand U2260 (N_2260,N_2123,N_2126);
nand U2261 (N_2261,N_2110,N_2180);
xor U2262 (N_2262,N_2158,N_2167);
or U2263 (N_2263,N_2131,N_2187);
or U2264 (N_2264,N_2137,N_2150);
and U2265 (N_2265,N_2199,N_2160);
nand U2266 (N_2266,N_2103,N_2193);
or U2267 (N_2267,N_2144,N_2151);
and U2268 (N_2268,N_2198,N_2128);
xor U2269 (N_2269,N_2147,N_2187);
nand U2270 (N_2270,N_2189,N_2106);
xnor U2271 (N_2271,N_2193,N_2176);
nor U2272 (N_2272,N_2177,N_2145);
xnor U2273 (N_2273,N_2188,N_2193);
and U2274 (N_2274,N_2177,N_2134);
or U2275 (N_2275,N_2126,N_2169);
nor U2276 (N_2276,N_2150,N_2146);
and U2277 (N_2277,N_2173,N_2151);
nor U2278 (N_2278,N_2154,N_2100);
xnor U2279 (N_2279,N_2157,N_2170);
xnor U2280 (N_2280,N_2187,N_2190);
or U2281 (N_2281,N_2137,N_2101);
nor U2282 (N_2282,N_2143,N_2160);
and U2283 (N_2283,N_2132,N_2183);
or U2284 (N_2284,N_2130,N_2167);
or U2285 (N_2285,N_2166,N_2181);
and U2286 (N_2286,N_2195,N_2156);
and U2287 (N_2287,N_2109,N_2197);
nor U2288 (N_2288,N_2167,N_2100);
or U2289 (N_2289,N_2112,N_2185);
nand U2290 (N_2290,N_2186,N_2110);
nor U2291 (N_2291,N_2120,N_2139);
and U2292 (N_2292,N_2139,N_2100);
nor U2293 (N_2293,N_2116,N_2139);
or U2294 (N_2294,N_2185,N_2171);
nor U2295 (N_2295,N_2159,N_2119);
and U2296 (N_2296,N_2168,N_2156);
or U2297 (N_2297,N_2189,N_2126);
xor U2298 (N_2298,N_2178,N_2144);
or U2299 (N_2299,N_2155,N_2156);
nor U2300 (N_2300,N_2272,N_2203);
and U2301 (N_2301,N_2256,N_2259);
nand U2302 (N_2302,N_2285,N_2280);
nor U2303 (N_2303,N_2293,N_2257);
nor U2304 (N_2304,N_2268,N_2232);
nor U2305 (N_2305,N_2281,N_2238);
xnor U2306 (N_2306,N_2266,N_2299);
xnor U2307 (N_2307,N_2210,N_2263);
nor U2308 (N_2308,N_2284,N_2229);
nor U2309 (N_2309,N_2252,N_2271);
nor U2310 (N_2310,N_2243,N_2234);
nand U2311 (N_2311,N_2264,N_2213);
or U2312 (N_2312,N_2277,N_2289);
nand U2313 (N_2313,N_2212,N_2270);
and U2314 (N_2314,N_2221,N_2202);
or U2315 (N_2315,N_2286,N_2295);
nor U2316 (N_2316,N_2237,N_2254);
nand U2317 (N_2317,N_2251,N_2292);
nand U2318 (N_2318,N_2242,N_2208);
or U2319 (N_2319,N_2290,N_2246);
nand U2320 (N_2320,N_2247,N_2206);
nand U2321 (N_2321,N_2245,N_2227);
xor U2322 (N_2322,N_2216,N_2249);
nor U2323 (N_2323,N_2215,N_2217);
nand U2324 (N_2324,N_2276,N_2269);
nand U2325 (N_2325,N_2223,N_2297);
nor U2326 (N_2326,N_2248,N_2230);
or U2327 (N_2327,N_2273,N_2235);
nor U2328 (N_2328,N_2250,N_2241);
xnor U2329 (N_2329,N_2278,N_2267);
and U2330 (N_2330,N_2261,N_2236);
and U2331 (N_2331,N_2265,N_2294);
nor U2332 (N_2332,N_2287,N_2220);
xor U2333 (N_2333,N_2291,N_2231);
xnor U2334 (N_2334,N_2282,N_2226);
and U2335 (N_2335,N_2298,N_2224);
nor U2336 (N_2336,N_2209,N_2255);
and U2337 (N_2337,N_2225,N_2296);
nor U2338 (N_2338,N_2233,N_2274);
or U2339 (N_2339,N_2262,N_2283);
and U2340 (N_2340,N_2204,N_2222);
xnor U2341 (N_2341,N_2244,N_2240);
and U2342 (N_2342,N_2258,N_2239);
or U2343 (N_2343,N_2211,N_2228);
xnor U2344 (N_2344,N_2214,N_2218);
nor U2345 (N_2345,N_2219,N_2260);
xnor U2346 (N_2346,N_2253,N_2201);
nand U2347 (N_2347,N_2279,N_2200);
or U2348 (N_2348,N_2275,N_2205);
nor U2349 (N_2349,N_2207,N_2288);
nor U2350 (N_2350,N_2285,N_2251);
nor U2351 (N_2351,N_2243,N_2223);
and U2352 (N_2352,N_2284,N_2204);
nand U2353 (N_2353,N_2234,N_2247);
and U2354 (N_2354,N_2209,N_2295);
nand U2355 (N_2355,N_2206,N_2266);
nand U2356 (N_2356,N_2234,N_2231);
nor U2357 (N_2357,N_2262,N_2252);
nand U2358 (N_2358,N_2263,N_2291);
nor U2359 (N_2359,N_2284,N_2238);
nor U2360 (N_2360,N_2259,N_2204);
or U2361 (N_2361,N_2257,N_2272);
nand U2362 (N_2362,N_2250,N_2292);
nand U2363 (N_2363,N_2207,N_2268);
nand U2364 (N_2364,N_2274,N_2230);
or U2365 (N_2365,N_2215,N_2254);
and U2366 (N_2366,N_2239,N_2257);
xnor U2367 (N_2367,N_2238,N_2266);
or U2368 (N_2368,N_2250,N_2245);
nor U2369 (N_2369,N_2224,N_2277);
nand U2370 (N_2370,N_2284,N_2251);
and U2371 (N_2371,N_2205,N_2241);
xor U2372 (N_2372,N_2299,N_2245);
nand U2373 (N_2373,N_2274,N_2285);
nor U2374 (N_2374,N_2207,N_2245);
nor U2375 (N_2375,N_2259,N_2268);
xnor U2376 (N_2376,N_2285,N_2201);
xor U2377 (N_2377,N_2235,N_2288);
or U2378 (N_2378,N_2252,N_2243);
and U2379 (N_2379,N_2220,N_2299);
xor U2380 (N_2380,N_2246,N_2222);
xnor U2381 (N_2381,N_2217,N_2238);
or U2382 (N_2382,N_2295,N_2212);
xnor U2383 (N_2383,N_2204,N_2278);
nor U2384 (N_2384,N_2268,N_2293);
or U2385 (N_2385,N_2219,N_2299);
nor U2386 (N_2386,N_2298,N_2294);
nand U2387 (N_2387,N_2234,N_2272);
or U2388 (N_2388,N_2202,N_2248);
xnor U2389 (N_2389,N_2226,N_2254);
or U2390 (N_2390,N_2287,N_2218);
nor U2391 (N_2391,N_2288,N_2266);
or U2392 (N_2392,N_2289,N_2261);
and U2393 (N_2393,N_2269,N_2290);
xor U2394 (N_2394,N_2281,N_2262);
xnor U2395 (N_2395,N_2205,N_2278);
or U2396 (N_2396,N_2225,N_2299);
nand U2397 (N_2397,N_2248,N_2252);
nand U2398 (N_2398,N_2203,N_2299);
nor U2399 (N_2399,N_2294,N_2275);
xor U2400 (N_2400,N_2359,N_2304);
nor U2401 (N_2401,N_2384,N_2348);
xor U2402 (N_2402,N_2325,N_2358);
xnor U2403 (N_2403,N_2393,N_2366);
nor U2404 (N_2404,N_2318,N_2326);
xnor U2405 (N_2405,N_2330,N_2365);
nand U2406 (N_2406,N_2334,N_2383);
and U2407 (N_2407,N_2382,N_2399);
and U2408 (N_2408,N_2369,N_2345);
xnor U2409 (N_2409,N_2355,N_2332);
and U2410 (N_2410,N_2367,N_2335);
nor U2411 (N_2411,N_2306,N_2341);
xor U2412 (N_2412,N_2338,N_2324);
nor U2413 (N_2413,N_2347,N_2308);
xor U2414 (N_2414,N_2375,N_2360);
nand U2415 (N_2415,N_2328,N_2396);
nor U2416 (N_2416,N_2374,N_2313);
and U2417 (N_2417,N_2309,N_2370);
nor U2418 (N_2418,N_2314,N_2391);
nor U2419 (N_2419,N_2303,N_2379);
nor U2420 (N_2420,N_2322,N_2352);
and U2421 (N_2421,N_2316,N_2372);
xnor U2422 (N_2422,N_2398,N_2389);
xor U2423 (N_2423,N_2305,N_2300);
nand U2424 (N_2424,N_2315,N_2376);
or U2425 (N_2425,N_2356,N_2337);
nor U2426 (N_2426,N_2339,N_2350);
or U2427 (N_2427,N_2336,N_2354);
nand U2428 (N_2428,N_2397,N_2386);
nor U2429 (N_2429,N_2394,N_2371);
and U2430 (N_2430,N_2343,N_2310);
nor U2431 (N_2431,N_2368,N_2395);
xor U2432 (N_2432,N_2317,N_2319);
and U2433 (N_2433,N_2311,N_2373);
or U2434 (N_2434,N_2312,N_2392);
nand U2435 (N_2435,N_2351,N_2346);
or U2436 (N_2436,N_2385,N_2349);
and U2437 (N_2437,N_2353,N_2387);
xor U2438 (N_2438,N_2333,N_2380);
nand U2439 (N_2439,N_2364,N_2320);
xor U2440 (N_2440,N_2321,N_2357);
nand U2441 (N_2441,N_2329,N_2331);
xnor U2442 (N_2442,N_2381,N_2307);
nand U2443 (N_2443,N_2327,N_2363);
nor U2444 (N_2444,N_2390,N_2301);
nand U2445 (N_2445,N_2377,N_2340);
xnor U2446 (N_2446,N_2388,N_2344);
xnor U2447 (N_2447,N_2361,N_2342);
and U2448 (N_2448,N_2302,N_2323);
and U2449 (N_2449,N_2362,N_2378);
or U2450 (N_2450,N_2334,N_2375);
or U2451 (N_2451,N_2321,N_2345);
nor U2452 (N_2452,N_2394,N_2311);
nand U2453 (N_2453,N_2360,N_2336);
nand U2454 (N_2454,N_2366,N_2352);
and U2455 (N_2455,N_2308,N_2323);
nand U2456 (N_2456,N_2362,N_2321);
nor U2457 (N_2457,N_2395,N_2356);
nor U2458 (N_2458,N_2364,N_2399);
and U2459 (N_2459,N_2304,N_2392);
or U2460 (N_2460,N_2390,N_2347);
nor U2461 (N_2461,N_2379,N_2359);
or U2462 (N_2462,N_2367,N_2385);
nor U2463 (N_2463,N_2358,N_2347);
nand U2464 (N_2464,N_2313,N_2302);
and U2465 (N_2465,N_2310,N_2382);
nor U2466 (N_2466,N_2391,N_2335);
and U2467 (N_2467,N_2328,N_2302);
xor U2468 (N_2468,N_2388,N_2336);
or U2469 (N_2469,N_2385,N_2375);
or U2470 (N_2470,N_2348,N_2382);
nor U2471 (N_2471,N_2313,N_2300);
nor U2472 (N_2472,N_2360,N_2346);
nor U2473 (N_2473,N_2352,N_2389);
nand U2474 (N_2474,N_2381,N_2338);
or U2475 (N_2475,N_2356,N_2387);
and U2476 (N_2476,N_2365,N_2351);
and U2477 (N_2477,N_2325,N_2367);
or U2478 (N_2478,N_2355,N_2321);
nor U2479 (N_2479,N_2319,N_2328);
or U2480 (N_2480,N_2364,N_2390);
or U2481 (N_2481,N_2318,N_2348);
and U2482 (N_2482,N_2321,N_2398);
nand U2483 (N_2483,N_2329,N_2382);
nor U2484 (N_2484,N_2392,N_2313);
or U2485 (N_2485,N_2305,N_2307);
nand U2486 (N_2486,N_2362,N_2312);
and U2487 (N_2487,N_2383,N_2306);
and U2488 (N_2488,N_2304,N_2397);
or U2489 (N_2489,N_2355,N_2399);
and U2490 (N_2490,N_2300,N_2344);
xnor U2491 (N_2491,N_2301,N_2342);
xnor U2492 (N_2492,N_2399,N_2345);
and U2493 (N_2493,N_2324,N_2330);
and U2494 (N_2494,N_2305,N_2356);
or U2495 (N_2495,N_2371,N_2310);
xor U2496 (N_2496,N_2301,N_2373);
and U2497 (N_2497,N_2336,N_2362);
or U2498 (N_2498,N_2391,N_2329);
and U2499 (N_2499,N_2373,N_2318);
xor U2500 (N_2500,N_2430,N_2482);
nor U2501 (N_2501,N_2415,N_2427);
or U2502 (N_2502,N_2408,N_2406);
nor U2503 (N_2503,N_2485,N_2464);
nand U2504 (N_2504,N_2454,N_2491);
and U2505 (N_2505,N_2442,N_2473);
and U2506 (N_2506,N_2433,N_2448);
nor U2507 (N_2507,N_2405,N_2423);
nor U2508 (N_2508,N_2431,N_2460);
and U2509 (N_2509,N_2416,N_2435);
and U2510 (N_2510,N_2422,N_2474);
nor U2511 (N_2511,N_2436,N_2470);
xnor U2512 (N_2512,N_2471,N_2444);
xnor U2513 (N_2513,N_2469,N_2409);
and U2514 (N_2514,N_2490,N_2451);
or U2515 (N_2515,N_2489,N_2443);
nand U2516 (N_2516,N_2447,N_2429);
nand U2517 (N_2517,N_2499,N_2428);
and U2518 (N_2518,N_2493,N_2487);
nor U2519 (N_2519,N_2479,N_2484);
xnor U2520 (N_2520,N_2400,N_2440);
nor U2521 (N_2521,N_2478,N_2465);
xnor U2522 (N_2522,N_2411,N_2421);
or U2523 (N_2523,N_2401,N_2456);
nand U2524 (N_2524,N_2403,N_2466);
and U2525 (N_2525,N_2412,N_2404);
nor U2526 (N_2526,N_2407,N_2462);
nor U2527 (N_2527,N_2441,N_2492);
nor U2528 (N_2528,N_2481,N_2432);
nor U2529 (N_2529,N_2498,N_2449);
nor U2530 (N_2530,N_2410,N_2486);
and U2531 (N_2531,N_2495,N_2475);
xnor U2532 (N_2532,N_2467,N_2418);
nor U2533 (N_2533,N_2450,N_2426);
nand U2534 (N_2534,N_2476,N_2414);
xnor U2535 (N_2535,N_2434,N_2497);
or U2536 (N_2536,N_2461,N_2458);
xnor U2537 (N_2537,N_2480,N_2402);
nand U2538 (N_2538,N_2438,N_2496);
xor U2539 (N_2539,N_2459,N_2445);
nand U2540 (N_2540,N_2424,N_2439);
xor U2541 (N_2541,N_2453,N_2446);
nand U2542 (N_2542,N_2417,N_2419);
nand U2543 (N_2543,N_2483,N_2488);
and U2544 (N_2544,N_2477,N_2413);
xor U2545 (N_2545,N_2468,N_2463);
nand U2546 (N_2546,N_2455,N_2494);
nor U2547 (N_2547,N_2437,N_2457);
and U2548 (N_2548,N_2452,N_2425);
xor U2549 (N_2549,N_2420,N_2472);
nor U2550 (N_2550,N_2452,N_2470);
nand U2551 (N_2551,N_2475,N_2485);
xnor U2552 (N_2552,N_2490,N_2444);
xnor U2553 (N_2553,N_2415,N_2490);
and U2554 (N_2554,N_2461,N_2429);
and U2555 (N_2555,N_2410,N_2464);
or U2556 (N_2556,N_2437,N_2499);
nor U2557 (N_2557,N_2491,N_2412);
nand U2558 (N_2558,N_2435,N_2448);
and U2559 (N_2559,N_2411,N_2444);
or U2560 (N_2560,N_2448,N_2430);
or U2561 (N_2561,N_2436,N_2400);
and U2562 (N_2562,N_2413,N_2466);
nand U2563 (N_2563,N_2437,N_2426);
nor U2564 (N_2564,N_2479,N_2411);
and U2565 (N_2565,N_2409,N_2488);
nor U2566 (N_2566,N_2448,N_2434);
xor U2567 (N_2567,N_2460,N_2401);
or U2568 (N_2568,N_2468,N_2486);
nand U2569 (N_2569,N_2474,N_2459);
xnor U2570 (N_2570,N_2499,N_2497);
and U2571 (N_2571,N_2476,N_2461);
and U2572 (N_2572,N_2401,N_2414);
nor U2573 (N_2573,N_2455,N_2467);
and U2574 (N_2574,N_2410,N_2453);
nor U2575 (N_2575,N_2468,N_2405);
nand U2576 (N_2576,N_2464,N_2472);
or U2577 (N_2577,N_2471,N_2438);
and U2578 (N_2578,N_2414,N_2494);
xnor U2579 (N_2579,N_2424,N_2409);
or U2580 (N_2580,N_2427,N_2492);
nor U2581 (N_2581,N_2478,N_2477);
nand U2582 (N_2582,N_2406,N_2476);
or U2583 (N_2583,N_2415,N_2417);
xnor U2584 (N_2584,N_2411,N_2471);
and U2585 (N_2585,N_2491,N_2466);
xnor U2586 (N_2586,N_2493,N_2446);
xor U2587 (N_2587,N_2483,N_2493);
nand U2588 (N_2588,N_2478,N_2410);
nand U2589 (N_2589,N_2401,N_2410);
or U2590 (N_2590,N_2472,N_2481);
and U2591 (N_2591,N_2492,N_2429);
or U2592 (N_2592,N_2447,N_2463);
nor U2593 (N_2593,N_2444,N_2424);
nand U2594 (N_2594,N_2416,N_2477);
nor U2595 (N_2595,N_2474,N_2409);
and U2596 (N_2596,N_2477,N_2482);
nand U2597 (N_2597,N_2440,N_2493);
or U2598 (N_2598,N_2442,N_2436);
nand U2599 (N_2599,N_2415,N_2491);
nor U2600 (N_2600,N_2527,N_2599);
xor U2601 (N_2601,N_2522,N_2549);
or U2602 (N_2602,N_2539,N_2506);
nor U2603 (N_2603,N_2579,N_2546);
nor U2604 (N_2604,N_2524,N_2538);
or U2605 (N_2605,N_2528,N_2501);
or U2606 (N_2606,N_2519,N_2563);
or U2607 (N_2607,N_2583,N_2573);
nand U2608 (N_2608,N_2591,N_2584);
and U2609 (N_2609,N_2525,N_2564);
xnor U2610 (N_2610,N_2574,N_2545);
or U2611 (N_2611,N_2521,N_2594);
nor U2612 (N_2612,N_2532,N_2540);
nand U2613 (N_2613,N_2534,N_2566);
nor U2614 (N_2614,N_2548,N_2553);
nor U2615 (N_2615,N_2511,N_2567);
or U2616 (N_2616,N_2557,N_2533);
nor U2617 (N_2617,N_2570,N_2544);
nor U2618 (N_2618,N_2550,N_2581);
or U2619 (N_2619,N_2518,N_2585);
and U2620 (N_2620,N_2576,N_2569);
and U2621 (N_2621,N_2523,N_2530);
xnor U2622 (N_2622,N_2582,N_2565);
nand U2623 (N_2623,N_2556,N_2587);
nand U2624 (N_2624,N_2592,N_2526);
and U2625 (N_2625,N_2547,N_2589);
or U2626 (N_2626,N_2572,N_2529);
nor U2627 (N_2627,N_2500,N_2520);
nand U2628 (N_2628,N_2537,N_2571);
xnor U2629 (N_2629,N_2504,N_2580);
or U2630 (N_2630,N_2560,N_2505);
or U2631 (N_2631,N_2516,N_2512);
nand U2632 (N_2632,N_2515,N_2517);
and U2633 (N_2633,N_2510,N_2593);
nand U2634 (N_2634,N_2558,N_2577);
nand U2635 (N_2635,N_2503,N_2531);
and U2636 (N_2636,N_2554,N_2541);
nand U2637 (N_2637,N_2507,N_2555);
xnor U2638 (N_2638,N_2535,N_2597);
nand U2639 (N_2639,N_2568,N_2596);
nand U2640 (N_2640,N_2562,N_2514);
nand U2641 (N_2641,N_2575,N_2561);
nor U2642 (N_2642,N_2551,N_2559);
nand U2643 (N_2643,N_2509,N_2588);
nor U2644 (N_2644,N_2543,N_2536);
and U2645 (N_2645,N_2502,N_2598);
xnor U2646 (N_2646,N_2513,N_2590);
nor U2647 (N_2647,N_2552,N_2578);
and U2648 (N_2648,N_2508,N_2595);
and U2649 (N_2649,N_2542,N_2586);
nand U2650 (N_2650,N_2550,N_2520);
and U2651 (N_2651,N_2508,N_2583);
xor U2652 (N_2652,N_2502,N_2571);
and U2653 (N_2653,N_2508,N_2527);
and U2654 (N_2654,N_2502,N_2552);
xnor U2655 (N_2655,N_2543,N_2573);
and U2656 (N_2656,N_2555,N_2539);
or U2657 (N_2657,N_2576,N_2596);
nand U2658 (N_2658,N_2576,N_2533);
nand U2659 (N_2659,N_2554,N_2536);
and U2660 (N_2660,N_2505,N_2520);
xor U2661 (N_2661,N_2530,N_2536);
xnor U2662 (N_2662,N_2517,N_2556);
nor U2663 (N_2663,N_2521,N_2504);
and U2664 (N_2664,N_2576,N_2577);
or U2665 (N_2665,N_2559,N_2563);
and U2666 (N_2666,N_2543,N_2521);
or U2667 (N_2667,N_2510,N_2578);
xnor U2668 (N_2668,N_2503,N_2521);
nor U2669 (N_2669,N_2582,N_2519);
and U2670 (N_2670,N_2568,N_2509);
or U2671 (N_2671,N_2566,N_2592);
xor U2672 (N_2672,N_2575,N_2595);
xor U2673 (N_2673,N_2536,N_2593);
nor U2674 (N_2674,N_2589,N_2529);
or U2675 (N_2675,N_2501,N_2505);
or U2676 (N_2676,N_2571,N_2554);
xnor U2677 (N_2677,N_2569,N_2540);
nand U2678 (N_2678,N_2558,N_2518);
nor U2679 (N_2679,N_2582,N_2549);
xnor U2680 (N_2680,N_2544,N_2582);
or U2681 (N_2681,N_2548,N_2511);
and U2682 (N_2682,N_2526,N_2534);
nand U2683 (N_2683,N_2578,N_2523);
and U2684 (N_2684,N_2503,N_2520);
or U2685 (N_2685,N_2514,N_2579);
and U2686 (N_2686,N_2539,N_2543);
nand U2687 (N_2687,N_2543,N_2568);
xnor U2688 (N_2688,N_2570,N_2511);
nor U2689 (N_2689,N_2542,N_2524);
or U2690 (N_2690,N_2572,N_2521);
nor U2691 (N_2691,N_2528,N_2538);
xor U2692 (N_2692,N_2588,N_2505);
and U2693 (N_2693,N_2563,N_2565);
xor U2694 (N_2694,N_2500,N_2501);
or U2695 (N_2695,N_2585,N_2520);
and U2696 (N_2696,N_2540,N_2543);
or U2697 (N_2697,N_2542,N_2570);
nor U2698 (N_2698,N_2579,N_2548);
nor U2699 (N_2699,N_2526,N_2533);
nand U2700 (N_2700,N_2633,N_2661);
or U2701 (N_2701,N_2613,N_2641);
and U2702 (N_2702,N_2697,N_2695);
xnor U2703 (N_2703,N_2614,N_2630);
and U2704 (N_2704,N_2651,N_2663);
nor U2705 (N_2705,N_2639,N_2658);
nor U2706 (N_2706,N_2665,N_2669);
nand U2707 (N_2707,N_2635,N_2690);
xnor U2708 (N_2708,N_2657,N_2683);
and U2709 (N_2709,N_2654,N_2649);
and U2710 (N_2710,N_2625,N_2674);
xnor U2711 (N_2711,N_2682,N_2622);
or U2712 (N_2712,N_2659,N_2642);
and U2713 (N_2713,N_2624,N_2667);
and U2714 (N_2714,N_2668,N_2646);
nor U2715 (N_2715,N_2672,N_2660);
xnor U2716 (N_2716,N_2604,N_2609);
or U2717 (N_2717,N_2617,N_2638);
or U2718 (N_2718,N_2645,N_2670);
nor U2719 (N_2719,N_2685,N_2601);
xor U2720 (N_2720,N_2687,N_2684);
nand U2721 (N_2721,N_2629,N_2644);
or U2722 (N_2722,N_2626,N_2666);
nand U2723 (N_2723,N_2696,N_2691);
and U2724 (N_2724,N_2608,N_2621);
or U2725 (N_2725,N_2676,N_2636);
nand U2726 (N_2726,N_2652,N_2662);
xnor U2727 (N_2727,N_2640,N_2647);
and U2728 (N_2728,N_2610,N_2653);
nor U2729 (N_2729,N_2627,N_2673);
nor U2730 (N_2730,N_2616,N_2664);
xnor U2731 (N_2731,N_2620,N_2602);
nor U2732 (N_2732,N_2600,N_2628);
or U2733 (N_2733,N_2619,N_2678);
or U2734 (N_2734,N_2648,N_2671);
nor U2735 (N_2735,N_2650,N_2656);
or U2736 (N_2736,N_2693,N_2611);
and U2737 (N_2737,N_2615,N_2603);
xnor U2738 (N_2738,N_2612,N_2632);
or U2739 (N_2739,N_2689,N_2637);
and U2740 (N_2740,N_2677,N_2631);
xor U2741 (N_2741,N_2699,N_2680);
and U2742 (N_2742,N_2634,N_2607);
or U2743 (N_2743,N_2681,N_2623);
or U2744 (N_2744,N_2679,N_2655);
nor U2745 (N_2745,N_2643,N_2698);
and U2746 (N_2746,N_2686,N_2688);
and U2747 (N_2747,N_2694,N_2692);
or U2748 (N_2748,N_2675,N_2605);
nand U2749 (N_2749,N_2606,N_2618);
or U2750 (N_2750,N_2677,N_2609);
xnor U2751 (N_2751,N_2661,N_2654);
xor U2752 (N_2752,N_2669,N_2677);
nand U2753 (N_2753,N_2694,N_2606);
or U2754 (N_2754,N_2687,N_2628);
or U2755 (N_2755,N_2697,N_2609);
and U2756 (N_2756,N_2658,N_2694);
nor U2757 (N_2757,N_2617,N_2640);
nor U2758 (N_2758,N_2670,N_2638);
nor U2759 (N_2759,N_2692,N_2625);
xnor U2760 (N_2760,N_2643,N_2675);
and U2761 (N_2761,N_2638,N_2693);
and U2762 (N_2762,N_2600,N_2615);
or U2763 (N_2763,N_2662,N_2620);
xor U2764 (N_2764,N_2614,N_2696);
or U2765 (N_2765,N_2618,N_2614);
or U2766 (N_2766,N_2605,N_2645);
and U2767 (N_2767,N_2647,N_2673);
or U2768 (N_2768,N_2666,N_2674);
or U2769 (N_2769,N_2696,N_2621);
xor U2770 (N_2770,N_2685,N_2666);
nor U2771 (N_2771,N_2656,N_2639);
or U2772 (N_2772,N_2650,N_2688);
and U2773 (N_2773,N_2688,N_2697);
xnor U2774 (N_2774,N_2656,N_2630);
or U2775 (N_2775,N_2602,N_2688);
nand U2776 (N_2776,N_2665,N_2633);
xor U2777 (N_2777,N_2670,N_2628);
nor U2778 (N_2778,N_2683,N_2654);
xnor U2779 (N_2779,N_2652,N_2673);
and U2780 (N_2780,N_2693,N_2665);
nor U2781 (N_2781,N_2617,N_2677);
xnor U2782 (N_2782,N_2683,N_2686);
nand U2783 (N_2783,N_2696,N_2688);
and U2784 (N_2784,N_2654,N_2692);
nor U2785 (N_2785,N_2657,N_2643);
nand U2786 (N_2786,N_2602,N_2684);
or U2787 (N_2787,N_2676,N_2632);
xnor U2788 (N_2788,N_2656,N_2617);
or U2789 (N_2789,N_2631,N_2643);
or U2790 (N_2790,N_2609,N_2685);
xnor U2791 (N_2791,N_2617,N_2637);
and U2792 (N_2792,N_2624,N_2653);
nand U2793 (N_2793,N_2629,N_2643);
nor U2794 (N_2794,N_2693,N_2655);
xnor U2795 (N_2795,N_2635,N_2632);
xor U2796 (N_2796,N_2699,N_2682);
nand U2797 (N_2797,N_2628,N_2676);
nor U2798 (N_2798,N_2646,N_2670);
xor U2799 (N_2799,N_2639,N_2645);
and U2800 (N_2800,N_2799,N_2770);
or U2801 (N_2801,N_2733,N_2756);
nor U2802 (N_2802,N_2784,N_2778);
nor U2803 (N_2803,N_2772,N_2711);
nand U2804 (N_2804,N_2723,N_2701);
xor U2805 (N_2805,N_2707,N_2781);
nand U2806 (N_2806,N_2790,N_2785);
or U2807 (N_2807,N_2731,N_2729);
or U2808 (N_2808,N_2740,N_2724);
xnor U2809 (N_2809,N_2705,N_2715);
xnor U2810 (N_2810,N_2721,N_2759);
and U2811 (N_2811,N_2792,N_2787);
xor U2812 (N_2812,N_2764,N_2755);
nor U2813 (N_2813,N_2745,N_2762);
nand U2814 (N_2814,N_2719,N_2777);
and U2815 (N_2815,N_2752,N_2709);
and U2816 (N_2816,N_2774,N_2737);
or U2817 (N_2817,N_2749,N_2776);
xnor U2818 (N_2818,N_2779,N_2797);
or U2819 (N_2819,N_2798,N_2738);
xnor U2820 (N_2820,N_2753,N_2750);
or U2821 (N_2821,N_2718,N_2710);
or U2822 (N_2822,N_2717,N_2708);
nand U2823 (N_2823,N_2725,N_2766);
nand U2824 (N_2824,N_2754,N_2735);
xor U2825 (N_2825,N_2713,N_2795);
xor U2826 (N_2826,N_2722,N_2775);
xor U2827 (N_2827,N_2761,N_2742);
and U2828 (N_2828,N_2760,N_2732);
or U2829 (N_2829,N_2706,N_2703);
or U2830 (N_2830,N_2789,N_2773);
xor U2831 (N_2831,N_2714,N_2702);
and U2832 (N_2832,N_2736,N_2739);
and U2833 (N_2833,N_2743,N_2712);
nand U2834 (N_2834,N_2771,N_2783);
nand U2835 (N_2835,N_2794,N_2728);
nand U2836 (N_2836,N_2747,N_2730);
nand U2837 (N_2837,N_2748,N_2726);
nor U2838 (N_2838,N_2796,N_2780);
and U2839 (N_2839,N_2746,N_2716);
nand U2840 (N_2840,N_2704,N_2769);
or U2841 (N_2841,N_2734,N_2763);
nand U2842 (N_2842,N_2720,N_2757);
or U2843 (N_2843,N_2788,N_2793);
or U2844 (N_2844,N_2751,N_2741);
nor U2845 (N_2845,N_2727,N_2791);
or U2846 (N_2846,N_2767,N_2786);
and U2847 (N_2847,N_2758,N_2700);
xor U2848 (N_2848,N_2744,N_2782);
nor U2849 (N_2849,N_2768,N_2765);
nand U2850 (N_2850,N_2790,N_2756);
xnor U2851 (N_2851,N_2746,N_2743);
or U2852 (N_2852,N_2701,N_2745);
and U2853 (N_2853,N_2703,N_2767);
xor U2854 (N_2854,N_2705,N_2724);
nand U2855 (N_2855,N_2756,N_2749);
xnor U2856 (N_2856,N_2799,N_2726);
and U2857 (N_2857,N_2704,N_2751);
nor U2858 (N_2858,N_2760,N_2782);
nor U2859 (N_2859,N_2736,N_2703);
and U2860 (N_2860,N_2761,N_2796);
and U2861 (N_2861,N_2736,N_2727);
or U2862 (N_2862,N_2711,N_2758);
nor U2863 (N_2863,N_2723,N_2753);
xor U2864 (N_2864,N_2709,N_2736);
nor U2865 (N_2865,N_2743,N_2749);
xor U2866 (N_2866,N_2785,N_2713);
or U2867 (N_2867,N_2785,N_2712);
and U2868 (N_2868,N_2767,N_2710);
nor U2869 (N_2869,N_2790,N_2722);
nor U2870 (N_2870,N_2722,N_2759);
xnor U2871 (N_2871,N_2778,N_2723);
nor U2872 (N_2872,N_2734,N_2782);
or U2873 (N_2873,N_2736,N_2722);
nand U2874 (N_2874,N_2727,N_2797);
or U2875 (N_2875,N_2714,N_2788);
nand U2876 (N_2876,N_2735,N_2717);
nand U2877 (N_2877,N_2732,N_2796);
nor U2878 (N_2878,N_2763,N_2775);
nor U2879 (N_2879,N_2704,N_2780);
or U2880 (N_2880,N_2719,N_2750);
nand U2881 (N_2881,N_2751,N_2765);
nor U2882 (N_2882,N_2701,N_2773);
nor U2883 (N_2883,N_2780,N_2742);
nand U2884 (N_2884,N_2714,N_2733);
nand U2885 (N_2885,N_2783,N_2760);
nand U2886 (N_2886,N_2700,N_2742);
nand U2887 (N_2887,N_2724,N_2744);
and U2888 (N_2888,N_2711,N_2754);
nand U2889 (N_2889,N_2709,N_2749);
nand U2890 (N_2890,N_2764,N_2705);
nand U2891 (N_2891,N_2708,N_2780);
or U2892 (N_2892,N_2791,N_2795);
or U2893 (N_2893,N_2767,N_2709);
nor U2894 (N_2894,N_2754,N_2783);
and U2895 (N_2895,N_2728,N_2703);
nor U2896 (N_2896,N_2711,N_2743);
nand U2897 (N_2897,N_2762,N_2784);
xor U2898 (N_2898,N_2722,N_2727);
xor U2899 (N_2899,N_2786,N_2704);
xor U2900 (N_2900,N_2824,N_2884);
xnor U2901 (N_2901,N_2835,N_2854);
or U2902 (N_2902,N_2883,N_2876);
nor U2903 (N_2903,N_2826,N_2805);
nand U2904 (N_2904,N_2808,N_2864);
nand U2905 (N_2905,N_2809,N_2870);
nor U2906 (N_2906,N_2877,N_2848);
nand U2907 (N_2907,N_2889,N_2822);
and U2908 (N_2908,N_2800,N_2850);
nand U2909 (N_2909,N_2810,N_2862);
or U2910 (N_2910,N_2820,N_2879);
xor U2911 (N_2911,N_2863,N_2828);
nand U2912 (N_2912,N_2853,N_2859);
nor U2913 (N_2913,N_2843,N_2855);
or U2914 (N_2914,N_2841,N_2885);
or U2915 (N_2915,N_2894,N_2811);
and U2916 (N_2916,N_2827,N_2823);
and U2917 (N_2917,N_2892,N_2873);
nand U2918 (N_2918,N_2857,N_2807);
or U2919 (N_2919,N_2801,N_2819);
nor U2920 (N_2920,N_2878,N_2804);
nand U2921 (N_2921,N_2866,N_2893);
nand U2922 (N_2922,N_2875,N_2851);
or U2923 (N_2923,N_2890,N_2869);
nor U2924 (N_2924,N_2898,N_2840);
nand U2925 (N_2925,N_2882,N_2895);
nand U2926 (N_2926,N_2865,N_2856);
or U2927 (N_2927,N_2846,N_2815);
nand U2928 (N_2928,N_2887,N_2896);
xor U2929 (N_2929,N_2837,N_2881);
nand U2930 (N_2930,N_2842,N_2821);
nand U2931 (N_2931,N_2802,N_2868);
xnor U2932 (N_2932,N_2871,N_2814);
or U2933 (N_2933,N_2886,N_2838);
nor U2934 (N_2934,N_2839,N_2861);
nand U2935 (N_2935,N_2888,N_2834);
or U2936 (N_2936,N_2852,N_2899);
nand U2937 (N_2937,N_2816,N_2825);
or U2938 (N_2938,N_2836,N_2844);
xnor U2939 (N_2939,N_2806,N_2830);
and U2940 (N_2940,N_2803,N_2872);
nor U2941 (N_2941,N_2874,N_2880);
nor U2942 (N_2942,N_2845,N_2818);
and U2943 (N_2943,N_2829,N_2813);
nand U2944 (N_2944,N_2847,N_2860);
and U2945 (N_2945,N_2833,N_2867);
and U2946 (N_2946,N_2817,N_2832);
or U2947 (N_2947,N_2849,N_2891);
nand U2948 (N_2948,N_2897,N_2831);
nor U2949 (N_2949,N_2812,N_2858);
nor U2950 (N_2950,N_2877,N_2808);
xor U2951 (N_2951,N_2800,N_2895);
nand U2952 (N_2952,N_2802,N_2809);
and U2953 (N_2953,N_2817,N_2809);
nor U2954 (N_2954,N_2889,N_2874);
xor U2955 (N_2955,N_2824,N_2879);
or U2956 (N_2956,N_2884,N_2840);
or U2957 (N_2957,N_2882,N_2843);
and U2958 (N_2958,N_2825,N_2830);
or U2959 (N_2959,N_2881,N_2824);
nand U2960 (N_2960,N_2820,N_2808);
xor U2961 (N_2961,N_2847,N_2885);
nor U2962 (N_2962,N_2807,N_2878);
nor U2963 (N_2963,N_2866,N_2820);
and U2964 (N_2964,N_2828,N_2811);
nand U2965 (N_2965,N_2821,N_2814);
nand U2966 (N_2966,N_2869,N_2851);
and U2967 (N_2967,N_2830,N_2812);
nor U2968 (N_2968,N_2860,N_2820);
or U2969 (N_2969,N_2870,N_2898);
nand U2970 (N_2970,N_2841,N_2845);
xor U2971 (N_2971,N_2830,N_2860);
nor U2972 (N_2972,N_2830,N_2827);
or U2973 (N_2973,N_2826,N_2847);
xnor U2974 (N_2974,N_2860,N_2894);
xor U2975 (N_2975,N_2872,N_2801);
and U2976 (N_2976,N_2890,N_2814);
nor U2977 (N_2977,N_2874,N_2865);
or U2978 (N_2978,N_2842,N_2849);
nor U2979 (N_2979,N_2807,N_2860);
nor U2980 (N_2980,N_2892,N_2829);
and U2981 (N_2981,N_2826,N_2888);
or U2982 (N_2982,N_2882,N_2898);
xor U2983 (N_2983,N_2895,N_2814);
nand U2984 (N_2984,N_2892,N_2808);
xnor U2985 (N_2985,N_2826,N_2804);
nand U2986 (N_2986,N_2864,N_2848);
xor U2987 (N_2987,N_2887,N_2889);
and U2988 (N_2988,N_2898,N_2835);
or U2989 (N_2989,N_2877,N_2875);
nand U2990 (N_2990,N_2870,N_2872);
or U2991 (N_2991,N_2873,N_2871);
and U2992 (N_2992,N_2834,N_2815);
nor U2993 (N_2993,N_2843,N_2864);
nor U2994 (N_2994,N_2848,N_2835);
or U2995 (N_2995,N_2866,N_2804);
and U2996 (N_2996,N_2861,N_2890);
or U2997 (N_2997,N_2865,N_2813);
or U2998 (N_2998,N_2846,N_2803);
nor U2999 (N_2999,N_2865,N_2885);
nor U3000 (N_3000,N_2972,N_2990);
xor U3001 (N_3001,N_2973,N_2996);
xor U3002 (N_3002,N_2920,N_2968);
nand U3003 (N_3003,N_2924,N_2938);
or U3004 (N_3004,N_2934,N_2932);
nor U3005 (N_3005,N_2904,N_2929);
or U3006 (N_3006,N_2919,N_2918);
and U3007 (N_3007,N_2952,N_2933);
nor U3008 (N_3008,N_2905,N_2999);
or U3009 (N_3009,N_2981,N_2993);
and U3010 (N_3010,N_2946,N_2953);
or U3011 (N_3011,N_2963,N_2912);
nor U3012 (N_3012,N_2967,N_2984);
xnor U3013 (N_3013,N_2983,N_2980);
or U3014 (N_3014,N_2957,N_2978);
nand U3015 (N_3015,N_2945,N_2921);
or U3016 (N_3016,N_2931,N_2958);
nand U3017 (N_3017,N_2965,N_2900);
or U3018 (N_3018,N_2916,N_2987);
xnor U3019 (N_3019,N_2975,N_2928);
nand U3020 (N_3020,N_2913,N_2992);
or U3021 (N_3021,N_2955,N_2922);
nand U3022 (N_3022,N_2977,N_2944);
nand U3023 (N_3023,N_2956,N_2943);
or U3024 (N_3024,N_2903,N_2909);
or U3025 (N_3025,N_2985,N_2964);
or U3026 (N_3026,N_2988,N_2917);
nand U3027 (N_3027,N_2991,N_2901);
xor U3028 (N_3028,N_2982,N_2907);
nand U3029 (N_3029,N_2902,N_2998);
and U3030 (N_3030,N_2954,N_2962);
or U3031 (N_3031,N_2936,N_2960);
or U3032 (N_3032,N_2935,N_2950);
nor U3033 (N_3033,N_2994,N_2923);
nand U3034 (N_3034,N_2997,N_2970);
and U3035 (N_3035,N_2942,N_2914);
xor U3036 (N_3036,N_2974,N_2949);
nor U3037 (N_3037,N_2947,N_2979);
nor U3038 (N_3038,N_2910,N_2976);
nor U3039 (N_3039,N_2940,N_2908);
and U3040 (N_3040,N_2995,N_2951);
nor U3041 (N_3041,N_2969,N_2930);
and U3042 (N_3042,N_2927,N_2926);
nor U3043 (N_3043,N_2915,N_2925);
or U3044 (N_3044,N_2966,N_2911);
nor U3045 (N_3045,N_2906,N_2971);
nor U3046 (N_3046,N_2941,N_2948);
or U3047 (N_3047,N_2986,N_2989);
and U3048 (N_3048,N_2961,N_2939);
nand U3049 (N_3049,N_2959,N_2937);
and U3050 (N_3050,N_2921,N_2913);
nand U3051 (N_3051,N_2938,N_2994);
xor U3052 (N_3052,N_2971,N_2902);
or U3053 (N_3053,N_2994,N_2974);
or U3054 (N_3054,N_2960,N_2958);
xnor U3055 (N_3055,N_2966,N_2965);
xor U3056 (N_3056,N_2948,N_2953);
nand U3057 (N_3057,N_2975,N_2927);
nor U3058 (N_3058,N_2996,N_2946);
or U3059 (N_3059,N_2903,N_2926);
or U3060 (N_3060,N_2945,N_2959);
xor U3061 (N_3061,N_2924,N_2926);
and U3062 (N_3062,N_2988,N_2927);
nand U3063 (N_3063,N_2932,N_2968);
and U3064 (N_3064,N_2921,N_2922);
and U3065 (N_3065,N_2939,N_2925);
xnor U3066 (N_3066,N_2919,N_2942);
nor U3067 (N_3067,N_2932,N_2982);
or U3068 (N_3068,N_2968,N_2936);
nor U3069 (N_3069,N_2940,N_2931);
nand U3070 (N_3070,N_2947,N_2951);
xnor U3071 (N_3071,N_2975,N_2968);
or U3072 (N_3072,N_2967,N_2939);
or U3073 (N_3073,N_2976,N_2963);
or U3074 (N_3074,N_2950,N_2971);
nor U3075 (N_3075,N_2996,N_2953);
xor U3076 (N_3076,N_2921,N_2996);
nand U3077 (N_3077,N_2921,N_2944);
nand U3078 (N_3078,N_2905,N_2963);
or U3079 (N_3079,N_2939,N_2974);
and U3080 (N_3080,N_2947,N_2969);
xor U3081 (N_3081,N_2921,N_2905);
or U3082 (N_3082,N_2959,N_2980);
nor U3083 (N_3083,N_2954,N_2991);
xnor U3084 (N_3084,N_2933,N_2909);
xnor U3085 (N_3085,N_2913,N_2922);
nor U3086 (N_3086,N_2929,N_2969);
nand U3087 (N_3087,N_2982,N_2938);
or U3088 (N_3088,N_2988,N_2905);
and U3089 (N_3089,N_2998,N_2973);
xor U3090 (N_3090,N_2962,N_2990);
or U3091 (N_3091,N_2958,N_2943);
nand U3092 (N_3092,N_2927,N_2990);
and U3093 (N_3093,N_2907,N_2989);
nand U3094 (N_3094,N_2924,N_2964);
xnor U3095 (N_3095,N_2946,N_2938);
and U3096 (N_3096,N_2977,N_2961);
nor U3097 (N_3097,N_2901,N_2937);
or U3098 (N_3098,N_2912,N_2937);
and U3099 (N_3099,N_2971,N_2955);
and U3100 (N_3100,N_3025,N_3097);
nor U3101 (N_3101,N_3086,N_3035);
or U3102 (N_3102,N_3064,N_3085);
nand U3103 (N_3103,N_3082,N_3042);
and U3104 (N_3104,N_3090,N_3089);
xor U3105 (N_3105,N_3065,N_3006);
xor U3106 (N_3106,N_3037,N_3076);
xnor U3107 (N_3107,N_3016,N_3077);
nand U3108 (N_3108,N_3001,N_3060);
xnor U3109 (N_3109,N_3027,N_3032);
xnor U3110 (N_3110,N_3002,N_3050);
or U3111 (N_3111,N_3023,N_3028);
xor U3112 (N_3112,N_3048,N_3069);
or U3113 (N_3113,N_3079,N_3092);
nor U3114 (N_3114,N_3039,N_3044);
or U3115 (N_3115,N_3078,N_3004);
nand U3116 (N_3116,N_3072,N_3084);
or U3117 (N_3117,N_3067,N_3013);
xnor U3118 (N_3118,N_3029,N_3088);
and U3119 (N_3119,N_3036,N_3075);
or U3120 (N_3120,N_3024,N_3056);
xor U3121 (N_3121,N_3099,N_3012);
xnor U3122 (N_3122,N_3033,N_3031);
and U3123 (N_3123,N_3055,N_3052);
xor U3124 (N_3124,N_3017,N_3094);
or U3125 (N_3125,N_3009,N_3026);
or U3126 (N_3126,N_3010,N_3018);
or U3127 (N_3127,N_3068,N_3080);
xor U3128 (N_3128,N_3019,N_3030);
nand U3129 (N_3129,N_3087,N_3093);
nand U3130 (N_3130,N_3070,N_3049);
nor U3131 (N_3131,N_3046,N_3074);
nand U3132 (N_3132,N_3081,N_3047);
or U3133 (N_3133,N_3011,N_3045);
xnor U3134 (N_3134,N_3014,N_3051);
or U3135 (N_3135,N_3091,N_3083);
nor U3136 (N_3136,N_3073,N_3041);
xor U3137 (N_3137,N_3053,N_3054);
nand U3138 (N_3138,N_3021,N_3057);
or U3139 (N_3139,N_3008,N_3096);
nor U3140 (N_3140,N_3059,N_3034);
and U3141 (N_3141,N_3038,N_3003);
and U3142 (N_3142,N_3095,N_3022);
nor U3143 (N_3143,N_3061,N_3098);
nor U3144 (N_3144,N_3071,N_3066);
xor U3145 (N_3145,N_3058,N_3062);
xor U3146 (N_3146,N_3063,N_3007);
nor U3147 (N_3147,N_3000,N_3020);
nand U3148 (N_3148,N_3015,N_3040);
nand U3149 (N_3149,N_3043,N_3005);
nor U3150 (N_3150,N_3076,N_3032);
nand U3151 (N_3151,N_3023,N_3021);
xnor U3152 (N_3152,N_3033,N_3091);
nor U3153 (N_3153,N_3099,N_3001);
or U3154 (N_3154,N_3011,N_3013);
and U3155 (N_3155,N_3071,N_3047);
nand U3156 (N_3156,N_3093,N_3034);
xnor U3157 (N_3157,N_3035,N_3001);
xnor U3158 (N_3158,N_3074,N_3018);
nor U3159 (N_3159,N_3083,N_3025);
or U3160 (N_3160,N_3068,N_3037);
nand U3161 (N_3161,N_3096,N_3092);
nand U3162 (N_3162,N_3066,N_3082);
xor U3163 (N_3163,N_3093,N_3027);
or U3164 (N_3164,N_3019,N_3074);
nor U3165 (N_3165,N_3092,N_3012);
nor U3166 (N_3166,N_3072,N_3044);
nand U3167 (N_3167,N_3051,N_3001);
nor U3168 (N_3168,N_3008,N_3037);
and U3169 (N_3169,N_3048,N_3020);
and U3170 (N_3170,N_3020,N_3035);
nor U3171 (N_3171,N_3010,N_3054);
xnor U3172 (N_3172,N_3010,N_3082);
nor U3173 (N_3173,N_3031,N_3091);
nor U3174 (N_3174,N_3094,N_3002);
nand U3175 (N_3175,N_3023,N_3082);
xor U3176 (N_3176,N_3019,N_3005);
nand U3177 (N_3177,N_3062,N_3045);
nor U3178 (N_3178,N_3013,N_3027);
xnor U3179 (N_3179,N_3097,N_3053);
xor U3180 (N_3180,N_3092,N_3051);
nand U3181 (N_3181,N_3024,N_3053);
xor U3182 (N_3182,N_3059,N_3037);
nor U3183 (N_3183,N_3099,N_3087);
and U3184 (N_3184,N_3019,N_3083);
nand U3185 (N_3185,N_3016,N_3070);
xor U3186 (N_3186,N_3025,N_3074);
and U3187 (N_3187,N_3032,N_3046);
nor U3188 (N_3188,N_3046,N_3099);
or U3189 (N_3189,N_3019,N_3041);
xnor U3190 (N_3190,N_3050,N_3037);
nor U3191 (N_3191,N_3087,N_3024);
and U3192 (N_3192,N_3007,N_3073);
nor U3193 (N_3193,N_3097,N_3033);
xor U3194 (N_3194,N_3063,N_3081);
or U3195 (N_3195,N_3067,N_3078);
or U3196 (N_3196,N_3062,N_3015);
nand U3197 (N_3197,N_3077,N_3022);
or U3198 (N_3198,N_3023,N_3055);
nor U3199 (N_3199,N_3051,N_3018);
nor U3200 (N_3200,N_3102,N_3192);
nand U3201 (N_3201,N_3146,N_3125);
xnor U3202 (N_3202,N_3155,N_3141);
and U3203 (N_3203,N_3169,N_3195);
nand U3204 (N_3204,N_3119,N_3156);
or U3205 (N_3205,N_3111,N_3110);
and U3206 (N_3206,N_3174,N_3144);
nand U3207 (N_3207,N_3168,N_3161);
nor U3208 (N_3208,N_3186,N_3182);
xnor U3209 (N_3209,N_3173,N_3178);
xor U3210 (N_3210,N_3131,N_3172);
nor U3211 (N_3211,N_3181,N_3198);
and U3212 (N_3212,N_3108,N_3167);
or U3213 (N_3213,N_3147,N_3193);
nand U3214 (N_3214,N_3133,N_3189);
nor U3215 (N_3215,N_3117,N_3116);
nand U3216 (N_3216,N_3114,N_3162);
or U3217 (N_3217,N_3159,N_3140);
or U3218 (N_3218,N_3179,N_3143);
or U3219 (N_3219,N_3139,N_3199);
nand U3220 (N_3220,N_3153,N_3164);
nor U3221 (N_3221,N_3151,N_3120);
or U3222 (N_3222,N_3190,N_3197);
nand U3223 (N_3223,N_3104,N_3113);
and U3224 (N_3224,N_3124,N_3170);
nor U3225 (N_3225,N_3149,N_3165);
and U3226 (N_3226,N_3103,N_3171);
nand U3227 (N_3227,N_3152,N_3123);
nor U3228 (N_3228,N_3128,N_3100);
nor U3229 (N_3229,N_3109,N_3121);
and U3230 (N_3230,N_3132,N_3127);
and U3231 (N_3231,N_3177,N_3136);
nor U3232 (N_3232,N_3129,N_3183);
nand U3233 (N_3233,N_3196,N_3191);
xor U3234 (N_3234,N_3115,N_3126);
or U3235 (N_3235,N_3142,N_3180);
xor U3236 (N_3236,N_3135,N_3176);
nand U3237 (N_3237,N_3163,N_3101);
nand U3238 (N_3238,N_3118,N_3122);
nor U3239 (N_3239,N_3105,N_3188);
nor U3240 (N_3240,N_3134,N_3148);
or U3241 (N_3241,N_3150,N_3187);
and U3242 (N_3242,N_3145,N_3175);
or U3243 (N_3243,N_3160,N_3106);
nand U3244 (N_3244,N_3112,N_3154);
nand U3245 (N_3245,N_3107,N_3157);
nand U3246 (N_3246,N_3130,N_3137);
nor U3247 (N_3247,N_3185,N_3166);
and U3248 (N_3248,N_3184,N_3138);
xnor U3249 (N_3249,N_3194,N_3158);
and U3250 (N_3250,N_3121,N_3111);
and U3251 (N_3251,N_3127,N_3181);
and U3252 (N_3252,N_3106,N_3147);
nor U3253 (N_3253,N_3189,N_3116);
nor U3254 (N_3254,N_3132,N_3165);
nand U3255 (N_3255,N_3153,N_3187);
nand U3256 (N_3256,N_3128,N_3164);
nand U3257 (N_3257,N_3149,N_3130);
xnor U3258 (N_3258,N_3168,N_3107);
nand U3259 (N_3259,N_3156,N_3148);
or U3260 (N_3260,N_3141,N_3171);
nand U3261 (N_3261,N_3149,N_3172);
or U3262 (N_3262,N_3118,N_3147);
and U3263 (N_3263,N_3132,N_3182);
xor U3264 (N_3264,N_3173,N_3120);
nand U3265 (N_3265,N_3138,N_3171);
and U3266 (N_3266,N_3199,N_3168);
nand U3267 (N_3267,N_3145,N_3179);
and U3268 (N_3268,N_3182,N_3108);
and U3269 (N_3269,N_3133,N_3109);
xnor U3270 (N_3270,N_3180,N_3158);
or U3271 (N_3271,N_3172,N_3132);
and U3272 (N_3272,N_3148,N_3184);
xor U3273 (N_3273,N_3178,N_3150);
xnor U3274 (N_3274,N_3149,N_3104);
and U3275 (N_3275,N_3165,N_3191);
xnor U3276 (N_3276,N_3140,N_3126);
nand U3277 (N_3277,N_3181,N_3146);
and U3278 (N_3278,N_3193,N_3146);
and U3279 (N_3279,N_3158,N_3199);
xor U3280 (N_3280,N_3117,N_3189);
nand U3281 (N_3281,N_3115,N_3135);
nand U3282 (N_3282,N_3176,N_3175);
nand U3283 (N_3283,N_3148,N_3180);
nand U3284 (N_3284,N_3112,N_3179);
nor U3285 (N_3285,N_3161,N_3156);
nor U3286 (N_3286,N_3164,N_3156);
or U3287 (N_3287,N_3136,N_3127);
or U3288 (N_3288,N_3106,N_3130);
nor U3289 (N_3289,N_3104,N_3191);
nand U3290 (N_3290,N_3163,N_3147);
nand U3291 (N_3291,N_3192,N_3173);
and U3292 (N_3292,N_3175,N_3160);
nor U3293 (N_3293,N_3165,N_3172);
nand U3294 (N_3294,N_3181,N_3123);
nor U3295 (N_3295,N_3162,N_3170);
nor U3296 (N_3296,N_3166,N_3103);
or U3297 (N_3297,N_3123,N_3109);
nand U3298 (N_3298,N_3102,N_3199);
or U3299 (N_3299,N_3121,N_3145);
xor U3300 (N_3300,N_3250,N_3281);
nor U3301 (N_3301,N_3273,N_3259);
nand U3302 (N_3302,N_3290,N_3209);
and U3303 (N_3303,N_3239,N_3202);
nand U3304 (N_3304,N_3298,N_3266);
nand U3305 (N_3305,N_3293,N_3228);
xor U3306 (N_3306,N_3297,N_3208);
nor U3307 (N_3307,N_3275,N_3288);
and U3308 (N_3308,N_3243,N_3295);
and U3309 (N_3309,N_3242,N_3279);
xor U3310 (N_3310,N_3223,N_3217);
or U3311 (N_3311,N_3233,N_3232);
or U3312 (N_3312,N_3265,N_3292);
nor U3313 (N_3313,N_3231,N_3286);
nor U3314 (N_3314,N_3227,N_3268);
xor U3315 (N_3315,N_3226,N_3216);
nor U3316 (N_3316,N_3284,N_3274);
nor U3317 (N_3317,N_3285,N_3264);
nand U3318 (N_3318,N_3218,N_3282);
nor U3319 (N_3319,N_3289,N_3251);
nand U3320 (N_3320,N_3254,N_3252);
nor U3321 (N_3321,N_3219,N_3258);
xor U3322 (N_3322,N_3230,N_3276);
nor U3323 (N_3323,N_3229,N_3244);
xor U3324 (N_3324,N_3207,N_3291);
nand U3325 (N_3325,N_3211,N_3249);
or U3326 (N_3326,N_3205,N_3246);
and U3327 (N_3327,N_3215,N_3255);
nor U3328 (N_3328,N_3269,N_3224);
xor U3329 (N_3329,N_3278,N_3247);
nand U3330 (N_3330,N_3238,N_3222);
or U3331 (N_3331,N_3271,N_3299);
nand U3332 (N_3332,N_3294,N_3283);
xor U3333 (N_3333,N_3201,N_3253);
nor U3334 (N_3334,N_3212,N_3237);
or U3335 (N_3335,N_3200,N_3241);
nand U3336 (N_3336,N_3267,N_3260);
xnor U3337 (N_3337,N_3220,N_3248);
nand U3338 (N_3338,N_3236,N_3210);
nand U3339 (N_3339,N_3296,N_3277);
and U3340 (N_3340,N_3245,N_3221);
xnor U3341 (N_3341,N_3280,N_3272);
and U3342 (N_3342,N_3235,N_3263);
or U3343 (N_3343,N_3203,N_3206);
nor U3344 (N_3344,N_3257,N_3234);
and U3345 (N_3345,N_3256,N_3262);
xnor U3346 (N_3346,N_3287,N_3225);
and U3347 (N_3347,N_3270,N_3240);
nor U3348 (N_3348,N_3214,N_3204);
nor U3349 (N_3349,N_3261,N_3213);
and U3350 (N_3350,N_3216,N_3231);
and U3351 (N_3351,N_3241,N_3276);
xor U3352 (N_3352,N_3205,N_3237);
and U3353 (N_3353,N_3273,N_3277);
and U3354 (N_3354,N_3236,N_3246);
nand U3355 (N_3355,N_3204,N_3287);
nor U3356 (N_3356,N_3260,N_3262);
nor U3357 (N_3357,N_3294,N_3260);
or U3358 (N_3358,N_3213,N_3290);
xnor U3359 (N_3359,N_3224,N_3262);
xor U3360 (N_3360,N_3279,N_3233);
xnor U3361 (N_3361,N_3286,N_3229);
xnor U3362 (N_3362,N_3261,N_3220);
xnor U3363 (N_3363,N_3210,N_3257);
nand U3364 (N_3364,N_3253,N_3213);
nand U3365 (N_3365,N_3276,N_3263);
nand U3366 (N_3366,N_3260,N_3271);
xor U3367 (N_3367,N_3247,N_3235);
nor U3368 (N_3368,N_3260,N_3204);
and U3369 (N_3369,N_3260,N_3257);
nor U3370 (N_3370,N_3215,N_3299);
xnor U3371 (N_3371,N_3214,N_3294);
or U3372 (N_3372,N_3229,N_3275);
nor U3373 (N_3373,N_3289,N_3253);
nand U3374 (N_3374,N_3280,N_3205);
and U3375 (N_3375,N_3279,N_3247);
and U3376 (N_3376,N_3277,N_3254);
nor U3377 (N_3377,N_3236,N_3213);
nor U3378 (N_3378,N_3230,N_3251);
nand U3379 (N_3379,N_3245,N_3272);
xnor U3380 (N_3380,N_3263,N_3219);
nor U3381 (N_3381,N_3237,N_3206);
or U3382 (N_3382,N_3267,N_3273);
and U3383 (N_3383,N_3267,N_3280);
nor U3384 (N_3384,N_3228,N_3259);
nor U3385 (N_3385,N_3234,N_3206);
and U3386 (N_3386,N_3298,N_3231);
nand U3387 (N_3387,N_3230,N_3207);
xnor U3388 (N_3388,N_3284,N_3287);
and U3389 (N_3389,N_3283,N_3281);
and U3390 (N_3390,N_3282,N_3299);
and U3391 (N_3391,N_3271,N_3220);
nor U3392 (N_3392,N_3212,N_3265);
nor U3393 (N_3393,N_3220,N_3233);
xor U3394 (N_3394,N_3295,N_3299);
and U3395 (N_3395,N_3215,N_3287);
xor U3396 (N_3396,N_3233,N_3236);
xnor U3397 (N_3397,N_3242,N_3236);
nand U3398 (N_3398,N_3272,N_3242);
xnor U3399 (N_3399,N_3270,N_3214);
xnor U3400 (N_3400,N_3387,N_3367);
and U3401 (N_3401,N_3354,N_3306);
nand U3402 (N_3402,N_3304,N_3355);
or U3403 (N_3403,N_3330,N_3398);
and U3404 (N_3404,N_3390,N_3326);
and U3405 (N_3405,N_3301,N_3356);
and U3406 (N_3406,N_3334,N_3382);
xor U3407 (N_3407,N_3378,N_3329);
nand U3408 (N_3408,N_3389,N_3362);
nor U3409 (N_3409,N_3305,N_3360);
nor U3410 (N_3410,N_3399,N_3302);
nand U3411 (N_3411,N_3363,N_3365);
nor U3412 (N_3412,N_3357,N_3352);
or U3413 (N_3413,N_3377,N_3333);
nor U3414 (N_3414,N_3337,N_3309);
and U3415 (N_3415,N_3374,N_3397);
nor U3416 (N_3416,N_3351,N_3336);
or U3417 (N_3417,N_3376,N_3368);
xnor U3418 (N_3418,N_3335,N_3350);
xor U3419 (N_3419,N_3339,N_3380);
nand U3420 (N_3420,N_3372,N_3386);
xor U3421 (N_3421,N_3394,N_3388);
nor U3422 (N_3422,N_3321,N_3361);
xnor U3423 (N_3423,N_3379,N_3349);
xnor U3424 (N_3424,N_3308,N_3338);
nand U3425 (N_3425,N_3371,N_3348);
and U3426 (N_3426,N_3340,N_3303);
nor U3427 (N_3427,N_3327,N_3359);
and U3428 (N_3428,N_3316,N_3395);
and U3429 (N_3429,N_3393,N_3300);
xnor U3430 (N_3430,N_3347,N_3320);
and U3431 (N_3431,N_3307,N_3319);
nand U3432 (N_3432,N_3396,N_3384);
or U3433 (N_3433,N_3358,N_3381);
xnor U3434 (N_3434,N_3314,N_3392);
xor U3435 (N_3435,N_3344,N_3353);
nand U3436 (N_3436,N_3318,N_3342);
and U3437 (N_3437,N_3312,N_3324);
and U3438 (N_3438,N_3328,N_3370);
nor U3439 (N_3439,N_3310,N_3317);
and U3440 (N_3440,N_3345,N_3346);
nand U3441 (N_3441,N_3341,N_3322);
nand U3442 (N_3442,N_3364,N_3385);
nor U3443 (N_3443,N_3375,N_3311);
nand U3444 (N_3444,N_3366,N_3373);
nor U3445 (N_3445,N_3331,N_3332);
nand U3446 (N_3446,N_3323,N_3313);
nor U3447 (N_3447,N_3369,N_3383);
or U3448 (N_3448,N_3315,N_3391);
nand U3449 (N_3449,N_3343,N_3325);
and U3450 (N_3450,N_3331,N_3382);
and U3451 (N_3451,N_3315,N_3386);
and U3452 (N_3452,N_3303,N_3328);
nor U3453 (N_3453,N_3334,N_3331);
and U3454 (N_3454,N_3311,N_3338);
nor U3455 (N_3455,N_3330,N_3353);
nand U3456 (N_3456,N_3372,N_3304);
xnor U3457 (N_3457,N_3314,N_3321);
xnor U3458 (N_3458,N_3369,N_3337);
nand U3459 (N_3459,N_3345,N_3307);
xnor U3460 (N_3460,N_3349,N_3372);
nand U3461 (N_3461,N_3323,N_3334);
and U3462 (N_3462,N_3367,N_3302);
and U3463 (N_3463,N_3353,N_3358);
nor U3464 (N_3464,N_3304,N_3390);
or U3465 (N_3465,N_3327,N_3308);
and U3466 (N_3466,N_3361,N_3317);
and U3467 (N_3467,N_3321,N_3344);
and U3468 (N_3468,N_3351,N_3303);
nand U3469 (N_3469,N_3351,N_3386);
nor U3470 (N_3470,N_3344,N_3382);
or U3471 (N_3471,N_3385,N_3315);
nor U3472 (N_3472,N_3316,N_3352);
nor U3473 (N_3473,N_3395,N_3371);
xnor U3474 (N_3474,N_3342,N_3383);
nor U3475 (N_3475,N_3302,N_3356);
xor U3476 (N_3476,N_3392,N_3375);
xor U3477 (N_3477,N_3315,N_3310);
nor U3478 (N_3478,N_3345,N_3392);
or U3479 (N_3479,N_3316,N_3317);
or U3480 (N_3480,N_3350,N_3300);
nor U3481 (N_3481,N_3398,N_3357);
and U3482 (N_3482,N_3350,N_3327);
and U3483 (N_3483,N_3397,N_3381);
nor U3484 (N_3484,N_3344,N_3360);
or U3485 (N_3485,N_3341,N_3370);
nor U3486 (N_3486,N_3395,N_3317);
nand U3487 (N_3487,N_3330,N_3343);
nor U3488 (N_3488,N_3364,N_3321);
nand U3489 (N_3489,N_3337,N_3373);
nand U3490 (N_3490,N_3308,N_3368);
nor U3491 (N_3491,N_3394,N_3336);
or U3492 (N_3492,N_3391,N_3363);
or U3493 (N_3493,N_3338,N_3307);
xnor U3494 (N_3494,N_3374,N_3370);
nand U3495 (N_3495,N_3320,N_3310);
nor U3496 (N_3496,N_3317,N_3323);
xnor U3497 (N_3497,N_3334,N_3383);
or U3498 (N_3498,N_3331,N_3399);
xor U3499 (N_3499,N_3395,N_3394);
nand U3500 (N_3500,N_3445,N_3419);
xnor U3501 (N_3501,N_3402,N_3400);
nor U3502 (N_3502,N_3439,N_3476);
xnor U3503 (N_3503,N_3494,N_3435);
or U3504 (N_3504,N_3474,N_3489);
or U3505 (N_3505,N_3407,N_3473);
xor U3506 (N_3506,N_3410,N_3415);
or U3507 (N_3507,N_3456,N_3451);
or U3508 (N_3508,N_3432,N_3464);
xor U3509 (N_3509,N_3418,N_3416);
xor U3510 (N_3510,N_3452,N_3479);
nor U3511 (N_3511,N_3436,N_3457);
nor U3512 (N_3512,N_3408,N_3412);
and U3513 (N_3513,N_3427,N_3441);
xor U3514 (N_3514,N_3491,N_3455);
nand U3515 (N_3515,N_3475,N_3487);
and U3516 (N_3516,N_3490,N_3434);
xor U3517 (N_3517,N_3460,N_3438);
nand U3518 (N_3518,N_3428,N_3403);
nor U3519 (N_3519,N_3458,N_3466);
nor U3520 (N_3520,N_3430,N_3449);
and U3521 (N_3521,N_3498,N_3485);
nor U3522 (N_3522,N_3459,N_3463);
and U3523 (N_3523,N_3404,N_3480);
or U3524 (N_3524,N_3461,N_3495);
xor U3525 (N_3525,N_3401,N_3411);
xnor U3526 (N_3526,N_3453,N_3421);
or U3527 (N_3527,N_3440,N_3446);
nand U3528 (N_3528,N_3409,N_3417);
xor U3529 (N_3529,N_3413,N_3447);
nand U3530 (N_3530,N_3420,N_3465);
and U3531 (N_3531,N_3481,N_3423);
and U3532 (N_3532,N_3422,N_3454);
and U3533 (N_3533,N_3468,N_3443);
nand U3534 (N_3534,N_3484,N_3492);
nor U3535 (N_3535,N_3450,N_3470);
xnor U3536 (N_3536,N_3477,N_3426);
or U3537 (N_3537,N_3482,N_3442);
or U3538 (N_3538,N_3437,N_3486);
xnor U3539 (N_3539,N_3467,N_3425);
xor U3540 (N_3540,N_3488,N_3414);
and U3541 (N_3541,N_3499,N_3424);
nor U3542 (N_3542,N_3444,N_3448);
nor U3543 (N_3543,N_3431,N_3471);
and U3544 (N_3544,N_3469,N_3478);
xnor U3545 (N_3545,N_3497,N_3483);
or U3546 (N_3546,N_3496,N_3472);
and U3547 (N_3547,N_3405,N_3493);
xnor U3548 (N_3548,N_3433,N_3429);
nand U3549 (N_3549,N_3462,N_3406);
and U3550 (N_3550,N_3445,N_3478);
nand U3551 (N_3551,N_3421,N_3455);
or U3552 (N_3552,N_3480,N_3487);
nor U3553 (N_3553,N_3434,N_3494);
nand U3554 (N_3554,N_3434,N_3436);
xor U3555 (N_3555,N_3453,N_3471);
or U3556 (N_3556,N_3461,N_3429);
xnor U3557 (N_3557,N_3434,N_3421);
or U3558 (N_3558,N_3488,N_3444);
and U3559 (N_3559,N_3423,N_3419);
and U3560 (N_3560,N_3444,N_3485);
xor U3561 (N_3561,N_3464,N_3423);
nor U3562 (N_3562,N_3475,N_3467);
or U3563 (N_3563,N_3450,N_3438);
nor U3564 (N_3564,N_3406,N_3441);
nor U3565 (N_3565,N_3460,N_3425);
nand U3566 (N_3566,N_3426,N_3468);
xor U3567 (N_3567,N_3446,N_3441);
nor U3568 (N_3568,N_3422,N_3473);
nor U3569 (N_3569,N_3436,N_3427);
or U3570 (N_3570,N_3452,N_3490);
and U3571 (N_3571,N_3475,N_3430);
nand U3572 (N_3572,N_3422,N_3457);
xor U3573 (N_3573,N_3406,N_3488);
and U3574 (N_3574,N_3401,N_3430);
nor U3575 (N_3575,N_3469,N_3431);
xor U3576 (N_3576,N_3496,N_3417);
and U3577 (N_3577,N_3470,N_3455);
and U3578 (N_3578,N_3416,N_3432);
nor U3579 (N_3579,N_3459,N_3469);
xor U3580 (N_3580,N_3472,N_3489);
and U3581 (N_3581,N_3426,N_3452);
nand U3582 (N_3582,N_3446,N_3490);
nor U3583 (N_3583,N_3405,N_3413);
nand U3584 (N_3584,N_3454,N_3409);
or U3585 (N_3585,N_3471,N_3496);
nor U3586 (N_3586,N_3420,N_3484);
nand U3587 (N_3587,N_3445,N_3480);
or U3588 (N_3588,N_3408,N_3456);
xnor U3589 (N_3589,N_3405,N_3476);
nand U3590 (N_3590,N_3431,N_3458);
and U3591 (N_3591,N_3435,N_3461);
xnor U3592 (N_3592,N_3423,N_3400);
nand U3593 (N_3593,N_3486,N_3491);
nor U3594 (N_3594,N_3492,N_3428);
nand U3595 (N_3595,N_3464,N_3497);
nor U3596 (N_3596,N_3438,N_3463);
and U3597 (N_3597,N_3431,N_3405);
nand U3598 (N_3598,N_3419,N_3485);
nand U3599 (N_3599,N_3441,N_3437);
nor U3600 (N_3600,N_3593,N_3591);
nand U3601 (N_3601,N_3508,N_3557);
and U3602 (N_3602,N_3599,N_3569);
nor U3603 (N_3603,N_3559,N_3547);
xnor U3604 (N_3604,N_3501,N_3558);
and U3605 (N_3605,N_3580,N_3512);
nand U3606 (N_3606,N_3540,N_3553);
nor U3607 (N_3607,N_3521,N_3525);
nand U3608 (N_3608,N_3586,N_3589);
nand U3609 (N_3609,N_3554,N_3581);
or U3610 (N_3610,N_3597,N_3595);
nor U3611 (N_3611,N_3565,N_3520);
nor U3612 (N_3612,N_3590,N_3573);
xor U3613 (N_3613,N_3594,N_3523);
nor U3614 (N_3614,N_3555,N_3535);
and U3615 (N_3615,N_3542,N_3544);
and U3616 (N_3616,N_3539,N_3550);
and U3617 (N_3617,N_3507,N_3505);
and U3618 (N_3618,N_3506,N_3564);
and U3619 (N_3619,N_3503,N_3598);
nor U3620 (N_3620,N_3538,N_3504);
xor U3621 (N_3621,N_3588,N_3543);
nand U3622 (N_3622,N_3570,N_3560);
nand U3623 (N_3623,N_3510,N_3596);
nand U3624 (N_3624,N_3519,N_3548);
xnor U3625 (N_3625,N_3561,N_3568);
nor U3626 (N_3626,N_3584,N_3526);
nand U3627 (N_3627,N_3511,N_3567);
nor U3628 (N_3628,N_3587,N_3502);
and U3629 (N_3629,N_3577,N_3533);
nand U3630 (N_3630,N_3592,N_3585);
and U3631 (N_3631,N_3513,N_3562);
and U3632 (N_3632,N_3579,N_3551);
nor U3633 (N_3633,N_3530,N_3516);
or U3634 (N_3634,N_3556,N_3578);
nor U3635 (N_3635,N_3500,N_3546);
xnor U3636 (N_3636,N_3522,N_3545);
or U3637 (N_3637,N_3531,N_3532);
and U3638 (N_3638,N_3534,N_3563);
nand U3639 (N_3639,N_3537,N_3576);
and U3640 (N_3640,N_3524,N_3574);
nor U3641 (N_3641,N_3515,N_3552);
or U3642 (N_3642,N_3572,N_3571);
and U3643 (N_3643,N_3549,N_3582);
xor U3644 (N_3644,N_3518,N_3528);
nor U3645 (N_3645,N_3529,N_3536);
xor U3646 (N_3646,N_3527,N_3514);
or U3647 (N_3647,N_3575,N_3517);
nand U3648 (N_3648,N_3583,N_3541);
nand U3649 (N_3649,N_3566,N_3509);
xor U3650 (N_3650,N_3500,N_3587);
and U3651 (N_3651,N_3589,N_3566);
or U3652 (N_3652,N_3507,N_3575);
nor U3653 (N_3653,N_3537,N_3571);
xnor U3654 (N_3654,N_3528,N_3527);
xor U3655 (N_3655,N_3552,N_3501);
or U3656 (N_3656,N_3577,N_3580);
xor U3657 (N_3657,N_3595,N_3599);
nor U3658 (N_3658,N_3538,N_3555);
xor U3659 (N_3659,N_3532,N_3528);
or U3660 (N_3660,N_3579,N_3576);
nor U3661 (N_3661,N_3541,N_3549);
nand U3662 (N_3662,N_3589,N_3584);
nor U3663 (N_3663,N_3522,N_3558);
nor U3664 (N_3664,N_3569,N_3542);
and U3665 (N_3665,N_3521,N_3556);
nor U3666 (N_3666,N_3562,N_3592);
nand U3667 (N_3667,N_3576,N_3527);
or U3668 (N_3668,N_3597,N_3552);
or U3669 (N_3669,N_3528,N_3566);
nor U3670 (N_3670,N_3596,N_3581);
xnor U3671 (N_3671,N_3560,N_3563);
nand U3672 (N_3672,N_3516,N_3524);
or U3673 (N_3673,N_3516,N_3554);
or U3674 (N_3674,N_3585,N_3502);
or U3675 (N_3675,N_3599,N_3501);
xnor U3676 (N_3676,N_3564,N_3512);
xnor U3677 (N_3677,N_3570,N_3594);
nor U3678 (N_3678,N_3540,N_3515);
nor U3679 (N_3679,N_3595,N_3526);
and U3680 (N_3680,N_3557,N_3560);
nor U3681 (N_3681,N_3592,N_3520);
nor U3682 (N_3682,N_3517,N_3516);
nor U3683 (N_3683,N_3523,N_3556);
or U3684 (N_3684,N_3550,N_3548);
xor U3685 (N_3685,N_3561,N_3594);
or U3686 (N_3686,N_3519,N_3541);
or U3687 (N_3687,N_3532,N_3518);
nand U3688 (N_3688,N_3559,N_3588);
nand U3689 (N_3689,N_3591,N_3537);
nand U3690 (N_3690,N_3513,N_3586);
nand U3691 (N_3691,N_3509,N_3599);
nand U3692 (N_3692,N_3571,N_3509);
xor U3693 (N_3693,N_3561,N_3572);
and U3694 (N_3694,N_3538,N_3573);
or U3695 (N_3695,N_3535,N_3579);
nor U3696 (N_3696,N_3544,N_3579);
or U3697 (N_3697,N_3557,N_3529);
nor U3698 (N_3698,N_3528,N_3579);
and U3699 (N_3699,N_3540,N_3594);
nor U3700 (N_3700,N_3649,N_3627);
nor U3701 (N_3701,N_3663,N_3612);
nand U3702 (N_3702,N_3645,N_3676);
nand U3703 (N_3703,N_3609,N_3643);
nor U3704 (N_3704,N_3652,N_3666);
or U3705 (N_3705,N_3653,N_3637);
nor U3706 (N_3706,N_3646,N_3628);
xor U3707 (N_3707,N_3678,N_3619);
and U3708 (N_3708,N_3670,N_3698);
and U3709 (N_3709,N_3648,N_3686);
or U3710 (N_3710,N_3669,N_3680);
and U3711 (N_3711,N_3658,N_3668);
nor U3712 (N_3712,N_3626,N_3616);
or U3713 (N_3713,N_3615,N_3682);
and U3714 (N_3714,N_3654,N_3673);
or U3715 (N_3715,N_3699,N_3642);
nor U3716 (N_3716,N_3667,N_3629);
nor U3717 (N_3717,N_3679,N_3631);
nor U3718 (N_3718,N_3639,N_3688);
xor U3719 (N_3719,N_3632,N_3657);
or U3720 (N_3720,N_3690,N_3607);
nand U3721 (N_3721,N_3601,N_3618);
nor U3722 (N_3722,N_3697,N_3656);
nand U3723 (N_3723,N_3677,N_3692);
nand U3724 (N_3724,N_3659,N_3693);
nand U3725 (N_3725,N_3623,N_3603);
nor U3726 (N_3726,N_3696,N_3625);
xnor U3727 (N_3727,N_3602,N_3662);
xnor U3728 (N_3728,N_3641,N_3611);
xor U3729 (N_3729,N_3689,N_3681);
nor U3730 (N_3730,N_3672,N_3633);
xor U3731 (N_3731,N_3651,N_3665);
nand U3732 (N_3732,N_3640,N_3635);
or U3733 (N_3733,N_3630,N_3675);
nor U3734 (N_3734,N_3660,N_3621);
or U3735 (N_3735,N_3655,N_3685);
xor U3736 (N_3736,N_3614,N_3620);
and U3737 (N_3737,N_3691,N_3617);
nand U3738 (N_3738,N_3606,N_3647);
nor U3739 (N_3739,N_3694,N_3610);
nor U3740 (N_3740,N_3624,N_3638);
and U3741 (N_3741,N_3604,N_3687);
or U3742 (N_3742,N_3664,N_3695);
nor U3743 (N_3743,N_3613,N_3683);
xnor U3744 (N_3744,N_3684,N_3622);
nand U3745 (N_3745,N_3608,N_3671);
nor U3746 (N_3746,N_3605,N_3634);
and U3747 (N_3747,N_3661,N_3600);
nor U3748 (N_3748,N_3650,N_3636);
nor U3749 (N_3749,N_3644,N_3674);
nor U3750 (N_3750,N_3601,N_3659);
or U3751 (N_3751,N_3680,N_3652);
or U3752 (N_3752,N_3634,N_3631);
xnor U3753 (N_3753,N_3620,N_3645);
xor U3754 (N_3754,N_3624,N_3691);
nand U3755 (N_3755,N_3695,N_3612);
nor U3756 (N_3756,N_3675,N_3644);
xor U3757 (N_3757,N_3651,N_3611);
nor U3758 (N_3758,N_3641,N_3690);
and U3759 (N_3759,N_3624,N_3675);
or U3760 (N_3760,N_3602,N_3618);
and U3761 (N_3761,N_3622,N_3623);
nand U3762 (N_3762,N_3647,N_3643);
nor U3763 (N_3763,N_3676,N_3642);
nor U3764 (N_3764,N_3656,N_3660);
xor U3765 (N_3765,N_3647,N_3690);
nor U3766 (N_3766,N_3691,N_3654);
nand U3767 (N_3767,N_3647,N_3636);
or U3768 (N_3768,N_3604,N_3641);
and U3769 (N_3769,N_3637,N_3669);
nor U3770 (N_3770,N_3605,N_3692);
nand U3771 (N_3771,N_3609,N_3640);
nor U3772 (N_3772,N_3640,N_3628);
xor U3773 (N_3773,N_3661,N_3644);
and U3774 (N_3774,N_3602,N_3639);
xnor U3775 (N_3775,N_3602,N_3669);
xnor U3776 (N_3776,N_3694,N_3617);
and U3777 (N_3777,N_3689,N_3668);
nand U3778 (N_3778,N_3608,N_3642);
nor U3779 (N_3779,N_3664,N_3607);
nand U3780 (N_3780,N_3640,N_3637);
nor U3781 (N_3781,N_3662,N_3616);
xnor U3782 (N_3782,N_3682,N_3667);
nand U3783 (N_3783,N_3673,N_3602);
nand U3784 (N_3784,N_3697,N_3611);
nor U3785 (N_3785,N_3602,N_3634);
nand U3786 (N_3786,N_3679,N_3655);
or U3787 (N_3787,N_3675,N_3659);
or U3788 (N_3788,N_3692,N_3613);
and U3789 (N_3789,N_3638,N_3608);
nor U3790 (N_3790,N_3638,N_3648);
nand U3791 (N_3791,N_3632,N_3616);
and U3792 (N_3792,N_3611,N_3604);
nor U3793 (N_3793,N_3611,N_3668);
nand U3794 (N_3794,N_3687,N_3657);
and U3795 (N_3795,N_3669,N_3643);
or U3796 (N_3796,N_3609,N_3624);
or U3797 (N_3797,N_3628,N_3605);
xnor U3798 (N_3798,N_3622,N_3611);
or U3799 (N_3799,N_3664,N_3690);
or U3800 (N_3800,N_3716,N_3774);
nor U3801 (N_3801,N_3739,N_3747);
nand U3802 (N_3802,N_3767,N_3749);
nor U3803 (N_3803,N_3799,N_3702);
nand U3804 (N_3804,N_3719,N_3787);
nor U3805 (N_3805,N_3797,N_3731);
xnor U3806 (N_3806,N_3715,N_3790);
and U3807 (N_3807,N_3707,N_3772);
or U3808 (N_3808,N_3730,N_3743);
nand U3809 (N_3809,N_3779,N_3735);
nand U3810 (N_3810,N_3725,N_3785);
xnor U3811 (N_3811,N_3717,N_3718);
nor U3812 (N_3812,N_3709,N_3750);
and U3813 (N_3813,N_3741,N_3792);
or U3814 (N_3814,N_3766,N_3740);
or U3815 (N_3815,N_3728,N_3759);
nor U3816 (N_3816,N_3753,N_3788);
nand U3817 (N_3817,N_3712,N_3789);
nand U3818 (N_3818,N_3781,N_3757);
and U3819 (N_3819,N_3729,N_3761);
nand U3820 (N_3820,N_3714,N_3724);
and U3821 (N_3821,N_3700,N_3798);
nand U3822 (N_3822,N_3706,N_3733);
nand U3823 (N_3823,N_3771,N_3710);
and U3824 (N_3824,N_3737,N_3756);
and U3825 (N_3825,N_3704,N_3708);
xnor U3826 (N_3826,N_3703,N_3726);
nand U3827 (N_3827,N_3754,N_3770);
nor U3828 (N_3828,N_3721,N_3763);
nor U3829 (N_3829,N_3723,N_3745);
nand U3830 (N_3830,N_3722,N_3780);
xor U3831 (N_3831,N_3796,N_3768);
xor U3832 (N_3832,N_3778,N_3775);
or U3833 (N_3833,N_3762,N_3748);
nand U3834 (N_3834,N_3777,N_3793);
or U3835 (N_3835,N_3736,N_3794);
nor U3836 (N_3836,N_3746,N_3783);
or U3837 (N_3837,N_3755,N_3720);
nand U3838 (N_3838,N_3782,N_3769);
nor U3839 (N_3839,N_3795,N_3742);
or U3840 (N_3840,N_3752,N_3784);
or U3841 (N_3841,N_3711,N_3727);
xnor U3842 (N_3842,N_3705,N_3744);
xnor U3843 (N_3843,N_3786,N_3713);
or U3844 (N_3844,N_3734,N_3764);
or U3845 (N_3845,N_3760,N_3776);
nand U3846 (N_3846,N_3773,N_3765);
xor U3847 (N_3847,N_3758,N_3751);
xnor U3848 (N_3848,N_3732,N_3701);
nand U3849 (N_3849,N_3738,N_3791);
nand U3850 (N_3850,N_3732,N_3792);
or U3851 (N_3851,N_3767,N_3743);
nand U3852 (N_3852,N_3770,N_3792);
and U3853 (N_3853,N_3787,N_3765);
nor U3854 (N_3854,N_3749,N_3766);
nor U3855 (N_3855,N_3746,N_3708);
nand U3856 (N_3856,N_3780,N_3716);
nand U3857 (N_3857,N_3764,N_3718);
nand U3858 (N_3858,N_3764,N_3784);
and U3859 (N_3859,N_3780,N_3701);
xnor U3860 (N_3860,N_3754,N_3798);
nor U3861 (N_3861,N_3776,N_3739);
nor U3862 (N_3862,N_3743,N_3763);
and U3863 (N_3863,N_3789,N_3792);
xor U3864 (N_3864,N_3783,N_3784);
xor U3865 (N_3865,N_3771,N_3784);
nor U3866 (N_3866,N_3788,N_3789);
nand U3867 (N_3867,N_3788,N_3756);
or U3868 (N_3868,N_3786,N_3706);
and U3869 (N_3869,N_3748,N_3746);
nor U3870 (N_3870,N_3725,N_3744);
or U3871 (N_3871,N_3731,N_3755);
nand U3872 (N_3872,N_3792,N_3734);
and U3873 (N_3873,N_3778,N_3755);
nor U3874 (N_3874,N_3726,N_3704);
nand U3875 (N_3875,N_3701,N_3728);
or U3876 (N_3876,N_3798,N_3740);
nand U3877 (N_3877,N_3729,N_3758);
and U3878 (N_3878,N_3758,N_3778);
and U3879 (N_3879,N_3783,N_3735);
nor U3880 (N_3880,N_3778,N_3729);
nor U3881 (N_3881,N_3738,N_3740);
or U3882 (N_3882,N_3720,N_3764);
nand U3883 (N_3883,N_3744,N_3788);
nor U3884 (N_3884,N_3794,N_3761);
nand U3885 (N_3885,N_3774,N_3766);
or U3886 (N_3886,N_3700,N_3776);
and U3887 (N_3887,N_3785,N_3721);
or U3888 (N_3888,N_3721,N_3748);
nor U3889 (N_3889,N_3768,N_3735);
and U3890 (N_3890,N_3732,N_3768);
nand U3891 (N_3891,N_3724,N_3754);
nor U3892 (N_3892,N_3735,N_3712);
and U3893 (N_3893,N_3757,N_3766);
xnor U3894 (N_3894,N_3718,N_3755);
or U3895 (N_3895,N_3742,N_3778);
and U3896 (N_3896,N_3713,N_3796);
and U3897 (N_3897,N_3789,N_3742);
or U3898 (N_3898,N_3726,N_3718);
nand U3899 (N_3899,N_3777,N_3773);
and U3900 (N_3900,N_3822,N_3887);
nor U3901 (N_3901,N_3862,N_3898);
or U3902 (N_3902,N_3873,N_3835);
nor U3903 (N_3903,N_3874,N_3851);
nor U3904 (N_3904,N_3858,N_3808);
or U3905 (N_3905,N_3863,N_3859);
nor U3906 (N_3906,N_3839,N_3888);
xor U3907 (N_3907,N_3848,N_3801);
nor U3908 (N_3908,N_3814,N_3815);
nor U3909 (N_3909,N_3849,N_3896);
nor U3910 (N_3910,N_3866,N_3834);
or U3911 (N_3911,N_3807,N_3832);
nor U3912 (N_3912,N_3861,N_3878);
xor U3913 (N_3913,N_3838,N_3872);
nor U3914 (N_3914,N_3899,N_3893);
and U3915 (N_3915,N_3854,N_3833);
nand U3916 (N_3916,N_3842,N_3847);
nor U3917 (N_3917,N_3850,N_3800);
or U3918 (N_3918,N_3841,N_3802);
nand U3919 (N_3919,N_3870,N_3864);
and U3920 (N_3920,N_3875,N_3892);
xnor U3921 (N_3921,N_3827,N_3837);
xor U3922 (N_3922,N_3811,N_3824);
or U3923 (N_3923,N_3868,N_3828);
and U3924 (N_3924,N_3894,N_3881);
and U3925 (N_3925,N_3880,N_3810);
or U3926 (N_3926,N_3805,N_3867);
or U3927 (N_3927,N_3886,N_3879);
and U3928 (N_3928,N_3844,N_3853);
xor U3929 (N_3929,N_3845,N_3897);
nor U3930 (N_3930,N_3813,N_3884);
nand U3931 (N_3931,N_3817,N_3869);
or U3932 (N_3932,N_3819,N_3843);
and U3933 (N_3933,N_3806,N_3871);
xnor U3934 (N_3934,N_3856,N_3852);
nor U3935 (N_3935,N_3877,N_3818);
or U3936 (N_3936,N_3809,N_3860);
or U3937 (N_3937,N_3836,N_3804);
nor U3938 (N_3938,N_3820,N_3876);
xor U3939 (N_3939,N_3825,N_3830);
and U3940 (N_3940,N_3857,N_3889);
xnor U3941 (N_3941,N_3882,N_3816);
xor U3942 (N_3942,N_3812,N_3885);
and U3943 (N_3943,N_3823,N_3803);
or U3944 (N_3944,N_3821,N_3865);
xnor U3945 (N_3945,N_3829,N_3826);
and U3946 (N_3946,N_3831,N_3895);
and U3947 (N_3947,N_3855,N_3840);
or U3948 (N_3948,N_3883,N_3846);
and U3949 (N_3949,N_3890,N_3891);
and U3950 (N_3950,N_3821,N_3881);
and U3951 (N_3951,N_3850,N_3840);
nor U3952 (N_3952,N_3874,N_3883);
xor U3953 (N_3953,N_3878,N_3865);
nand U3954 (N_3954,N_3810,N_3806);
nand U3955 (N_3955,N_3803,N_3894);
xnor U3956 (N_3956,N_3873,N_3804);
or U3957 (N_3957,N_3809,N_3865);
xor U3958 (N_3958,N_3867,N_3850);
xnor U3959 (N_3959,N_3894,N_3880);
or U3960 (N_3960,N_3884,N_3888);
nand U3961 (N_3961,N_3816,N_3877);
and U3962 (N_3962,N_3805,N_3865);
nand U3963 (N_3963,N_3886,N_3880);
or U3964 (N_3964,N_3889,N_3878);
or U3965 (N_3965,N_3855,N_3801);
xnor U3966 (N_3966,N_3879,N_3878);
and U3967 (N_3967,N_3826,N_3895);
xor U3968 (N_3968,N_3815,N_3868);
xor U3969 (N_3969,N_3869,N_3894);
nand U3970 (N_3970,N_3852,N_3816);
xor U3971 (N_3971,N_3866,N_3809);
or U3972 (N_3972,N_3895,N_3813);
nor U3973 (N_3973,N_3876,N_3875);
and U3974 (N_3974,N_3851,N_3853);
nand U3975 (N_3975,N_3814,N_3898);
nor U3976 (N_3976,N_3802,N_3804);
and U3977 (N_3977,N_3822,N_3888);
or U3978 (N_3978,N_3852,N_3870);
xor U3979 (N_3979,N_3895,N_3821);
nor U3980 (N_3980,N_3812,N_3886);
and U3981 (N_3981,N_3836,N_3807);
or U3982 (N_3982,N_3840,N_3899);
nand U3983 (N_3983,N_3850,N_3813);
nand U3984 (N_3984,N_3875,N_3810);
xnor U3985 (N_3985,N_3825,N_3809);
nor U3986 (N_3986,N_3819,N_3870);
xor U3987 (N_3987,N_3828,N_3826);
xnor U3988 (N_3988,N_3821,N_3889);
xor U3989 (N_3989,N_3805,N_3842);
nand U3990 (N_3990,N_3867,N_3896);
xnor U3991 (N_3991,N_3843,N_3892);
and U3992 (N_3992,N_3891,N_3860);
xnor U3993 (N_3993,N_3880,N_3863);
nand U3994 (N_3994,N_3800,N_3863);
xnor U3995 (N_3995,N_3885,N_3889);
or U3996 (N_3996,N_3847,N_3866);
xor U3997 (N_3997,N_3874,N_3830);
nor U3998 (N_3998,N_3871,N_3863);
and U3999 (N_3999,N_3822,N_3897);
and U4000 (N_4000,N_3921,N_3983);
xnor U4001 (N_4001,N_3914,N_3985);
nand U4002 (N_4002,N_3980,N_3918);
xor U4003 (N_4003,N_3960,N_3979);
nor U4004 (N_4004,N_3930,N_3932);
and U4005 (N_4005,N_3969,N_3942);
or U4006 (N_4006,N_3948,N_3966);
and U4007 (N_4007,N_3944,N_3926);
or U4008 (N_4008,N_3964,N_3925);
xor U4009 (N_4009,N_3940,N_3997);
xnor U4010 (N_4010,N_3945,N_3965);
xnor U4011 (N_4011,N_3974,N_3988);
nor U4012 (N_4012,N_3976,N_3950);
or U4013 (N_4013,N_3919,N_3935);
nand U4014 (N_4014,N_3990,N_3920);
nor U4015 (N_4015,N_3994,N_3975);
nand U4016 (N_4016,N_3995,N_3906);
and U4017 (N_4017,N_3998,N_3991);
nor U4018 (N_4018,N_3913,N_3970);
or U4019 (N_4019,N_3917,N_3924);
nand U4020 (N_4020,N_3992,N_3996);
xor U4021 (N_4021,N_3951,N_3916);
or U4022 (N_4022,N_3981,N_3939);
or U4023 (N_4023,N_3987,N_3963);
xor U4024 (N_4024,N_3973,N_3989);
nand U4025 (N_4025,N_3923,N_3908);
or U4026 (N_4026,N_3900,N_3956);
and U4027 (N_4027,N_3943,N_3903);
or U4028 (N_4028,N_3911,N_3953);
and U4029 (N_4029,N_3901,N_3986);
or U4030 (N_4030,N_3931,N_3922);
and U4031 (N_4031,N_3928,N_3910);
nor U4032 (N_4032,N_3909,N_3927);
and U4033 (N_4033,N_3961,N_3904);
nor U4034 (N_4034,N_3912,N_3982);
nand U4035 (N_4035,N_3915,N_3936);
nand U4036 (N_4036,N_3962,N_3907);
or U4037 (N_4037,N_3947,N_3946);
nor U4038 (N_4038,N_3977,N_3933);
nor U4039 (N_4039,N_3968,N_3967);
xor U4040 (N_4040,N_3978,N_3949);
nor U4041 (N_4041,N_3955,N_3958);
nand U4042 (N_4042,N_3934,N_3938);
xor U4043 (N_4043,N_3937,N_3972);
or U4044 (N_4044,N_3902,N_3993);
nor U4045 (N_4045,N_3999,N_3905);
and U4046 (N_4046,N_3941,N_3952);
and U4047 (N_4047,N_3984,N_3971);
and U4048 (N_4048,N_3954,N_3929);
nand U4049 (N_4049,N_3957,N_3959);
or U4050 (N_4050,N_3949,N_3939);
nand U4051 (N_4051,N_3942,N_3916);
nor U4052 (N_4052,N_3914,N_3947);
nand U4053 (N_4053,N_3991,N_3965);
nor U4054 (N_4054,N_3998,N_3955);
nor U4055 (N_4055,N_3924,N_3901);
nand U4056 (N_4056,N_3967,N_3911);
nor U4057 (N_4057,N_3912,N_3998);
nor U4058 (N_4058,N_3987,N_3977);
nand U4059 (N_4059,N_3975,N_3935);
xnor U4060 (N_4060,N_3931,N_3909);
xor U4061 (N_4061,N_3942,N_3909);
or U4062 (N_4062,N_3990,N_3902);
nand U4063 (N_4063,N_3943,N_3941);
nand U4064 (N_4064,N_3991,N_3939);
nand U4065 (N_4065,N_3924,N_3943);
nand U4066 (N_4066,N_3970,N_3918);
nor U4067 (N_4067,N_3967,N_3915);
and U4068 (N_4068,N_3954,N_3909);
xor U4069 (N_4069,N_3967,N_3954);
nor U4070 (N_4070,N_3993,N_3911);
xnor U4071 (N_4071,N_3997,N_3964);
xnor U4072 (N_4072,N_3986,N_3970);
nand U4073 (N_4073,N_3975,N_3940);
and U4074 (N_4074,N_3965,N_3992);
or U4075 (N_4075,N_3983,N_3984);
and U4076 (N_4076,N_3963,N_3977);
nor U4077 (N_4077,N_3927,N_3993);
or U4078 (N_4078,N_3934,N_3992);
and U4079 (N_4079,N_3912,N_3929);
xnor U4080 (N_4080,N_3926,N_3991);
and U4081 (N_4081,N_3946,N_3936);
nand U4082 (N_4082,N_3979,N_3907);
or U4083 (N_4083,N_3959,N_3920);
nor U4084 (N_4084,N_3990,N_3926);
xor U4085 (N_4085,N_3940,N_3922);
or U4086 (N_4086,N_3911,N_3903);
nand U4087 (N_4087,N_3957,N_3926);
or U4088 (N_4088,N_3917,N_3970);
nor U4089 (N_4089,N_3902,N_3950);
xnor U4090 (N_4090,N_3990,N_3968);
or U4091 (N_4091,N_3987,N_3988);
nor U4092 (N_4092,N_3920,N_3985);
or U4093 (N_4093,N_3910,N_3948);
nor U4094 (N_4094,N_3974,N_3919);
nand U4095 (N_4095,N_3919,N_3970);
nor U4096 (N_4096,N_3940,N_3921);
or U4097 (N_4097,N_3923,N_3987);
and U4098 (N_4098,N_3995,N_3959);
and U4099 (N_4099,N_3903,N_3928);
xnor U4100 (N_4100,N_4057,N_4099);
nand U4101 (N_4101,N_4051,N_4085);
nor U4102 (N_4102,N_4069,N_4078);
xnor U4103 (N_4103,N_4015,N_4035);
nand U4104 (N_4104,N_4070,N_4072);
nor U4105 (N_4105,N_4005,N_4033);
nor U4106 (N_4106,N_4020,N_4062);
nor U4107 (N_4107,N_4058,N_4025);
nor U4108 (N_4108,N_4000,N_4011);
nor U4109 (N_4109,N_4083,N_4076);
xor U4110 (N_4110,N_4093,N_4013);
or U4111 (N_4111,N_4063,N_4071);
and U4112 (N_4112,N_4016,N_4045);
or U4113 (N_4113,N_4054,N_4049);
or U4114 (N_4114,N_4089,N_4024);
nor U4115 (N_4115,N_4046,N_4066);
or U4116 (N_4116,N_4075,N_4052);
or U4117 (N_4117,N_4034,N_4061);
nand U4118 (N_4118,N_4044,N_4021);
and U4119 (N_4119,N_4030,N_4048);
xnor U4120 (N_4120,N_4023,N_4001);
nand U4121 (N_4121,N_4038,N_4092);
xor U4122 (N_4122,N_4042,N_4002);
or U4123 (N_4123,N_4067,N_4014);
or U4124 (N_4124,N_4094,N_4032);
or U4125 (N_4125,N_4098,N_4018);
and U4126 (N_4126,N_4084,N_4055);
and U4127 (N_4127,N_4087,N_4037);
or U4128 (N_4128,N_4074,N_4047);
nand U4129 (N_4129,N_4040,N_4003);
and U4130 (N_4130,N_4012,N_4029);
or U4131 (N_4131,N_4019,N_4081);
nor U4132 (N_4132,N_4008,N_4004);
or U4133 (N_4133,N_4077,N_4068);
nand U4134 (N_4134,N_4031,N_4065);
nand U4135 (N_4135,N_4073,N_4027);
nand U4136 (N_4136,N_4060,N_4043);
nor U4137 (N_4137,N_4036,N_4050);
xor U4138 (N_4138,N_4064,N_4091);
xor U4139 (N_4139,N_4010,N_4026);
or U4140 (N_4140,N_4028,N_4096);
nor U4141 (N_4141,N_4080,N_4006);
nand U4142 (N_4142,N_4017,N_4082);
nor U4143 (N_4143,N_4009,N_4039);
nand U4144 (N_4144,N_4095,N_4022);
and U4145 (N_4145,N_4090,N_4086);
and U4146 (N_4146,N_4053,N_4088);
nand U4147 (N_4147,N_4041,N_4056);
or U4148 (N_4148,N_4079,N_4059);
or U4149 (N_4149,N_4097,N_4007);
nor U4150 (N_4150,N_4086,N_4092);
xor U4151 (N_4151,N_4048,N_4089);
and U4152 (N_4152,N_4029,N_4014);
xor U4153 (N_4153,N_4087,N_4006);
nand U4154 (N_4154,N_4057,N_4025);
and U4155 (N_4155,N_4002,N_4014);
xnor U4156 (N_4156,N_4093,N_4038);
or U4157 (N_4157,N_4019,N_4093);
nor U4158 (N_4158,N_4085,N_4095);
nand U4159 (N_4159,N_4054,N_4057);
or U4160 (N_4160,N_4026,N_4067);
or U4161 (N_4161,N_4015,N_4091);
nor U4162 (N_4162,N_4002,N_4050);
or U4163 (N_4163,N_4090,N_4091);
nor U4164 (N_4164,N_4019,N_4082);
nor U4165 (N_4165,N_4085,N_4072);
or U4166 (N_4166,N_4027,N_4017);
xor U4167 (N_4167,N_4043,N_4057);
xor U4168 (N_4168,N_4049,N_4063);
nor U4169 (N_4169,N_4052,N_4054);
nor U4170 (N_4170,N_4059,N_4069);
xnor U4171 (N_4171,N_4074,N_4026);
or U4172 (N_4172,N_4065,N_4012);
nor U4173 (N_4173,N_4048,N_4003);
nand U4174 (N_4174,N_4038,N_4071);
nand U4175 (N_4175,N_4087,N_4083);
and U4176 (N_4176,N_4083,N_4059);
xor U4177 (N_4177,N_4092,N_4079);
xor U4178 (N_4178,N_4098,N_4012);
nor U4179 (N_4179,N_4089,N_4012);
xor U4180 (N_4180,N_4093,N_4004);
nand U4181 (N_4181,N_4027,N_4090);
nor U4182 (N_4182,N_4082,N_4058);
and U4183 (N_4183,N_4019,N_4028);
nor U4184 (N_4184,N_4076,N_4054);
nor U4185 (N_4185,N_4094,N_4042);
nand U4186 (N_4186,N_4054,N_4027);
xnor U4187 (N_4187,N_4066,N_4031);
or U4188 (N_4188,N_4066,N_4053);
or U4189 (N_4189,N_4074,N_4059);
or U4190 (N_4190,N_4022,N_4016);
nand U4191 (N_4191,N_4075,N_4055);
nor U4192 (N_4192,N_4084,N_4012);
and U4193 (N_4193,N_4013,N_4003);
nor U4194 (N_4194,N_4051,N_4017);
nand U4195 (N_4195,N_4053,N_4090);
nand U4196 (N_4196,N_4009,N_4017);
or U4197 (N_4197,N_4093,N_4092);
or U4198 (N_4198,N_4015,N_4066);
nor U4199 (N_4199,N_4001,N_4025);
xor U4200 (N_4200,N_4105,N_4129);
xor U4201 (N_4201,N_4117,N_4110);
nand U4202 (N_4202,N_4190,N_4199);
and U4203 (N_4203,N_4162,N_4112);
or U4204 (N_4204,N_4160,N_4109);
nor U4205 (N_4205,N_4175,N_4139);
or U4206 (N_4206,N_4178,N_4195);
and U4207 (N_4207,N_4187,N_4186);
and U4208 (N_4208,N_4155,N_4168);
nand U4209 (N_4209,N_4191,N_4184);
or U4210 (N_4210,N_4165,N_4176);
xor U4211 (N_4211,N_4102,N_4100);
xnor U4212 (N_4212,N_4120,N_4136);
nor U4213 (N_4213,N_4137,N_4174);
or U4214 (N_4214,N_4138,N_4185);
or U4215 (N_4215,N_4140,N_4169);
or U4216 (N_4216,N_4170,N_4152);
nor U4217 (N_4217,N_4159,N_4127);
or U4218 (N_4218,N_4149,N_4189);
or U4219 (N_4219,N_4147,N_4132);
xnor U4220 (N_4220,N_4157,N_4115);
nand U4221 (N_4221,N_4193,N_4103);
nand U4222 (N_4222,N_4180,N_4131);
or U4223 (N_4223,N_4163,N_4153);
and U4224 (N_4224,N_4148,N_4177);
xnor U4225 (N_4225,N_4146,N_4167);
or U4226 (N_4226,N_4158,N_4106);
xnor U4227 (N_4227,N_4118,N_4124);
nand U4228 (N_4228,N_4183,N_4107);
nor U4229 (N_4229,N_4196,N_4114);
xor U4230 (N_4230,N_4182,N_4198);
or U4231 (N_4231,N_4135,N_4181);
or U4232 (N_4232,N_4104,N_4113);
nor U4233 (N_4233,N_4150,N_4142);
or U4234 (N_4234,N_4134,N_4164);
or U4235 (N_4235,N_4172,N_4122);
nor U4236 (N_4236,N_4161,N_4133);
nor U4237 (N_4237,N_4121,N_4128);
xor U4238 (N_4238,N_4154,N_4108);
and U4239 (N_4239,N_4125,N_4126);
and U4240 (N_4240,N_4151,N_4111);
nand U4241 (N_4241,N_4197,N_4130);
xor U4242 (N_4242,N_4116,N_4145);
xor U4243 (N_4243,N_4192,N_4119);
nand U4244 (N_4244,N_4166,N_4188);
nand U4245 (N_4245,N_4179,N_4194);
xnor U4246 (N_4246,N_4156,N_4123);
xor U4247 (N_4247,N_4171,N_4143);
xnor U4248 (N_4248,N_4101,N_4144);
and U4249 (N_4249,N_4141,N_4173);
nor U4250 (N_4250,N_4199,N_4187);
nor U4251 (N_4251,N_4131,N_4195);
xnor U4252 (N_4252,N_4127,N_4177);
and U4253 (N_4253,N_4127,N_4112);
and U4254 (N_4254,N_4147,N_4103);
nor U4255 (N_4255,N_4120,N_4158);
or U4256 (N_4256,N_4130,N_4193);
xor U4257 (N_4257,N_4145,N_4174);
and U4258 (N_4258,N_4195,N_4117);
or U4259 (N_4259,N_4144,N_4106);
nor U4260 (N_4260,N_4183,N_4179);
nand U4261 (N_4261,N_4117,N_4193);
nor U4262 (N_4262,N_4109,N_4171);
nor U4263 (N_4263,N_4119,N_4149);
or U4264 (N_4264,N_4138,N_4111);
or U4265 (N_4265,N_4129,N_4115);
nand U4266 (N_4266,N_4111,N_4135);
or U4267 (N_4267,N_4103,N_4184);
nor U4268 (N_4268,N_4169,N_4151);
or U4269 (N_4269,N_4144,N_4102);
nor U4270 (N_4270,N_4171,N_4100);
and U4271 (N_4271,N_4161,N_4138);
or U4272 (N_4272,N_4140,N_4155);
nor U4273 (N_4273,N_4196,N_4162);
nand U4274 (N_4274,N_4133,N_4148);
or U4275 (N_4275,N_4114,N_4160);
and U4276 (N_4276,N_4105,N_4126);
xor U4277 (N_4277,N_4179,N_4150);
xnor U4278 (N_4278,N_4151,N_4160);
nand U4279 (N_4279,N_4192,N_4153);
nor U4280 (N_4280,N_4172,N_4174);
xor U4281 (N_4281,N_4164,N_4173);
nand U4282 (N_4282,N_4169,N_4185);
xor U4283 (N_4283,N_4159,N_4141);
nor U4284 (N_4284,N_4185,N_4142);
nand U4285 (N_4285,N_4151,N_4125);
and U4286 (N_4286,N_4190,N_4187);
xnor U4287 (N_4287,N_4161,N_4121);
xnor U4288 (N_4288,N_4130,N_4107);
or U4289 (N_4289,N_4161,N_4120);
nand U4290 (N_4290,N_4176,N_4185);
or U4291 (N_4291,N_4134,N_4176);
xor U4292 (N_4292,N_4141,N_4185);
and U4293 (N_4293,N_4157,N_4193);
nor U4294 (N_4294,N_4106,N_4186);
nor U4295 (N_4295,N_4162,N_4152);
and U4296 (N_4296,N_4155,N_4123);
xnor U4297 (N_4297,N_4143,N_4127);
nand U4298 (N_4298,N_4127,N_4107);
nand U4299 (N_4299,N_4195,N_4177);
nand U4300 (N_4300,N_4281,N_4229);
xor U4301 (N_4301,N_4218,N_4206);
and U4302 (N_4302,N_4216,N_4266);
nor U4303 (N_4303,N_4238,N_4267);
nor U4304 (N_4304,N_4260,N_4217);
nor U4305 (N_4305,N_4273,N_4246);
nand U4306 (N_4306,N_4258,N_4274);
xor U4307 (N_4307,N_4295,N_4255);
nand U4308 (N_4308,N_4248,N_4240);
or U4309 (N_4309,N_4253,N_4270);
nor U4310 (N_4310,N_4294,N_4288);
nand U4311 (N_4311,N_4215,N_4230);
nor U4312 (N_4312,N_4282,N_4247);
xor U4313 (N_4313,N_4221,N_4239);
nor U4314 (N_4314,N_4223,N_4297);
nor U4315 (N_4315,N_4219,N_4234);
and U4316 (N_4316,N_4244,N_4202);
and U4317 (N_4317,N_4210,N_4211);
xor U4318 (N_4318,N_4222,N_4256);
nor U4319 (N_4319,N_4277,N_4205);
and U4320 (N_4320,N_4250,N_4241);
nand U4321 (N_4321,N_4226,N_4263);
nor U4322 (N_4322,N_4236,N_4291);
or U4323 (N_4323,N_4200,N_4299);
nand U4324 (N_4324,N_4235,N_4287);
or U4325 (N_4325,N_4220,N_4269);
or U4326 (N_4326,N_4237,N_4212);
and U4327 (N_4327,N_4257,N_4280);
nand U4328 (N_4328,N_4284,N_4224);
nand U4329 (N_4329,N_4271,N_4261);
xor U4330 (N_4330,N_4214,N_4213);
or U4331 (N_4331,N_4231,N_4298);
or U4332 (N_4332,N_4245,N_4276);
xor U4333 (N_4333,N_4251,N_4279);
nor U4334 (N_4334,N_4264,N_4228);
xor U4335 (N_4335,N_4259,N_4233);
and U4336 (N_4336,N_4243,N_4285);
and U4337 (N_4337,N_4296,N_4252);
nor U4338 (N_4338,N_4207,N_4292);
or U4339 (N_4339,N_4275,N_4278);
nor U4340 (N_4340,N_4254,N_4272);
and U4341 (N_4341,N_4201,N_4283);
and U4342 (N_4342,N_4242,N_4265);
xnor U4343 (N_4343,N_4289,N_4290);
nor U4344 (N_4344,N_4209,N_4268);
and U4345 (N_4345,N_4286,N_4227);
nor U4346 (N_4346,N_4262,N_4203);
nor U4347 (N_4347,N_4249,N_4232);
or U4348 (N_4348,N_4293,N_4225);
nand U4349 (N_4349,N_4208,N_4204);
xnor U4350 (N_4350,N_4225,N_4204);
nand U4351 (N_4351,N_4265,N_4283);
nand U4352 (N_4352,N_4216,N_4294);
nand U4353 (N_4353,N_4210,N_4255);
nor U4354 (N_4354,N_4277,N_4244);
or U4355 (N_4355,N_4255,N_4242);
xor U4356 (N_4356,N_4279,N_4260);
or U4357 (N_4357,N_4269,N_4242);
nor U4358 (N_4358,N_4269,N_4277);
nor U4359 (N_4359,N_4252,N_4220);
or U4360 (N_4360,N_4211,N_4257);
nor U4361 (N_4361,N_4267,N_4215);
or U4362 (N_4362,N_4299,N_4297);
xnor U4363 (N_4363,N_4285,N_4229);
nand U4364 (N_4364,N_4271,N_4257);
or U4365 (N_4365,N_4299,N_4257);
nand U4366 (N_4366,N_4297,N_4286);
and U4367 (N_4367,N_4238,N_4258);
xor U4368 (N_4368,N_4240,N_4243);
nor U4369 (N_4369,N_4273,N_4238);
or U4370 (N_4370,N_4239,N_4287);
nand U4371 (N_4371,N_4212,N_4242);
or U4372 (N_4372,N_4298,N_4264);
or U4373 (N_4373,N_4229,N_4275);
nor U4374 (N_4374,N_4245,N_4226);
nand U4375 (N_4375,N_4209,N_4210);
nand U4376 (N_4376,N_4288,N_4274);
nor U4377 (N_4377,N_4266,N_4255);
xnor U4378 (N_4378,N_4296,N_4292);
and U4379 (N_4379,N_4221,N_4292);
nand U4380 (N_4380,N_4294,N_4237);
nand U4381 (N_4381,N_4211,N_4264);
and U4382 (N_4382,N_4214,N_4281);
or U4383 (N_4383,N_4263,N_4224);
or U4384 (N_4384,N_4221,N_4230);
xnor U4385 (N_4385,N_4288,N_4247);
xor U4386 (N_4386,N_4209,N_4265);
or U4387 (N_4387,N_4258,N_4222);
or U4388 (N_4388,N_4206,N_4234);
or U4389 (N_4389,N_4202,N_4251);
nor U4390 (N_4390,N_4224,N_4200);
nand U4391 (N_4391,N_4218,N_4229);
and U4392 (N_4392,N_4260,N_4267);
xnor U4393 (N_4393,N_4281,N_4237);
nand U4394 (N_4394,N_4237,N_4298);
nand U4395 (N_4395,N_4241,N_4244);
xnor U4396 (N_4396,N_4298,N_4240);
and U4397 (N_4397,N_4202,N_4205);
nand U4398 (N_4398,N_4296,N_4215);
or U4399 (N_4399,N_4249,N_4226);
xnor U4400 (N_4400,N_4314,N_4335);
and U4401 (N_4401,N_4349,N_4391);
nor U4402 (N_4402,N_4393,N_4394);
xnor U4403 (N_4403,N_4380,N_4344);
or U4404 (N_4404,N_4332,N_4310);
or U4405 (N_4405,N_4334,N_4359);
xor U4406 (N_4406,N_4395,N_4304);
and U4407 (N_4407,N_4363,N_4374);
nand U4408 (N_4408,N_4318,N_4343);
or U4409 (N_4409,N_4301,N_4340);
or U4410 (N_4410,N_4312,N_4383);
or U4411 (N_4411,N_4371,N_4317);
and U4412 (N_4412,N_4341,N_4324);
nor U4413 (N_4413,N_4326,N_4373);
nor U4414 (N_4414,N_4339,N_4369);
nor U4415 (N_4415,N_4353,N_4355);
xor U4416 (N_4416,N_4364,N_4375);
xnor U4417 (N_4417,N_4336,N_4348);
and U4418 (N_4418,N_4356,N_4351);
nor U4419 (N_4419,N_4322,N_4307);
and U4420 (N_4420,N_4350,N_4362);
and U4421 (N_4421,N_4309,N_4366);
or U4422 (N_4422,N_4308,N_4382);
nand U4423 (N_4423,N_4305,N_4361);
nand U4424 (N_4424,N_4384,N_4365);
nand U4425 (N_4425,N_4320,N_4378);
or U4426 (N_4426,N_4397,N_4302);
nor U4427 (N_4427,N_4372,N_4370);
nand U4428 (N_4428,N_4300,N_4338);
nor U4429 (N_4429,N_4345,N_4377);
nand U4430 (N_4430,N_4311,N_4325);
or U4431 (N_4431,N_4390,N_4329);
or U4432 (N_4432,N_4346,N_4313);
and U4433 (N_4433,N_4368,N_4399);
or U4434 (N_4434,N_4327,N_4316);
xor U4435 (N_4435,N_4386,N_4303);
nor U4436 (N_4436,N_4354,N_4385);
xnor U4437 (N_4437,N_4360,N_4379);
nand U4438 (N_4438,N_4398,N_4306);
and U4439 (N_4439,N_4376,N_4342);
or U4440 (N_4440,N_4321,N_4323);
nand U4441 (N_4441,N_4381,N_4333);
and U4442 (N_4442,N_4392,N_4337);
nor U4443 (N_4443,N_4319,N_4388);
nor U4444 (N_4444,N_4352,N_4331);
or U4445 (N_4445,N_4389,N_4387);
nor U4446 (N_4446,N_4315,N_4347);
and U4447 (N_4447,N_4358,N_4396);
xor U4448 (N_4448,N_4330,N_4367);
or U4449 (N_4449,N_4328,N_4357);
xnor U4450 (N_4450,N_4329,N_4386);
nand U4451 (N_4451,N_4366,N_4328);
xnor U4452 (N_4452,N_4383,N_4392);
nand U4453 (N_4453,N_4392,N_4336);
nor U4454 (N_4454,N_4326,N_4325);
nand U4455 (N_4455,N_4329,N_4389);
nand U4456 (N_4456,N_4381,N_4357);
nand U4457 (N_4457,N_4399,N_4310);
and U4458 (N_4458,N_4348,N_4330);
nand U4459 (N_4459,N_4306,N_4393);
or U4460 (N_4460,N_4397,N_4335);
and U4461 (N_4461,N_4348,N_4315);
nor U4462 (N_4462,N_4340,N_4359);
nor U4463 (N_4463,N_4378,N_4334);
and U4464 (N_4464,N_4346,N_4369);
xnor U4465 (N_4465,N_4318,N_4348);
and U4466 (N_4466,N_4322,N_4349);
nor U4467 (N_4467,N_4327,N_4395);
and U4468 (N_4468,N_4307,N_4305);
and U4469 (N_4469,N_4373,N_4315);
or U4470 (N_4470,N_4349,N_4312);
xor U4471 (N_4471,N_4346,N_4308);
nand U4472 (N_4472,N_4382,N_4312);
and U4473 (N_4473,N_4358,N_4316);
or U4474 (N_4474,N_4368,N_4365);
and U4475 (N_4475,N_4374,N_4348);
or U4476 (N_4476,N_4359,N_4388);
nand U4477 (N_4477,N_4376,N_4356);
and U4478 (N_4478,N_4307,N_4378);
or U4479 (N_4479,N_4305,N_4363);
or U4480 (N_4480,N_4381,N_4383);
or U4481 (N_4481,N_4303,N_4324);
or U4482 (N_4482,N_4311,N_4300);
and U4483 (N_4483,N_4376,N_4328);
nand U4484 (N_4484,N_4355,N_4317);
nand U4485 (N_4485,N_4318,N_4321);
nor U4486 (N_4486,N_4330,N_4379);
and U4487 (N_4487,N_4387,N_4315);
and U4488 (N_4488,N_4305,N_4303);
and U4489 (N_4489,N_4301,N_4322);
xnor U4490 (N_4490,N_4394,N_4303);
nor U4491 (N_4491,N_4398,N_4330);
xor U4492 (N_4492,N_4303,N_4315);
nor U4493 (N_4493,N_4382,N_4338);
and U4494 (N_4494,N_4332,N_4353);
and U4495 (N_4495,N_4329,N_4365);
and U4496 (N_4496,N_4314,N_4387);
nor U4497 (N_4497,N_4397,N_4305);
nor U4498 (N_4498,N_4341,N_4332);
and U4499 (N_4499,N_4394,N_4351);
and U4500 (N_4500,N_4477,N_4444);
nand U4501 (N_4501,N_4401,N_4422);
nor U4502 (N_4502,N_4459,N_4463);
xor U4503 (N_4503,N_4436,N_4405);
xor U4504 (N_4504,N_4473,N_4440);
or U4505 (N_4505,N_4450,N_4455);
xor U4506 (N_4506,N_4487,N_4486);
and U4507 (N_4507,N_4439,N_4469);
or U4508 (N_4508,N_4404,N_4496);
and U4509 (N_4509,N_4482,N_4483);
and U4510 (N_4510,N_4433,N_4474);
or U4511 (N_4511,N_4411,N_4428);
or U4512 (N_4512,N_4408,N_4495);
and U4513 (N_4513,N_4475,N_4445);
xnor U4514 (N_4514,N_4493,N_4458);
nand U4515 (N_4515,N_4492,N_4490);
or U4516 (N_4516,N_4464,N_4431);
or U4517 (N_4517,N_4494,N_4441);
xnor U4518 (N_4518,N_4403,N_4400);
nand U4519 (N_4519,N_4468,N_4437);
xnor U4520 (N_4520,N_4413,N_4443);
nand U4521 (N_4521,N_4407,N_4456);
and U4522 (N_4522,N_4423,N_4457);
or U4523 (N_4523,N_4470,N_4489);
or U4524 (N_4524,N_4402,N_4452);
and U4525 (N_4525,N_4499,N_4447);
nor U4526 (N_4526,N_4479,N_4434);
nor U4527 (N_4527,N_4446,N_4467);
nand U4528 (N_4528,N_4485,N_4432);
or U4529 (N_4529,N_4449,N_4430);
nor U4530 (N_4530,N_4488,N_4419);
nor U4531 (N_4531,N_4465,N_4448);
nand U4532 (N_4532,N_4484,N_4497);
and U4533 (N_4533,N_4453,N_4466);
nor U4534 (N_4534,N_4410,N_4438);
or U4535 (N_4535,N_4454,N_4416);
nand U4536 (N_4536,N_4427,N_4406);
or U4537 (N_4537,N_4414,N_4476);
or U4538 (N_4538,N_4426,N_4471);
and U4539 (N_4539,N_4462,N_4425);
xnor U4540 (N_4540,N_4498,N_4418);
nand U4541 (N_4541,N_4478,N_4420);
and U4542 (N_4542,N_4421,N_4429);
nor U4543 (N_4543,N_4415,N_4412);
xor U4544 (N_4544,N_4435,N_4481);
xnor U4545 (N_4545,N_4472,N_4480);
xor U4546 (N_4546,N_4461,N_4491);
xnor U4547 (N_4547,N_4451,N_4460);
and U4548 (N_4548,N_4417,N_4424);
or U4549 (N_4549,N_4409,N_4442);
nor U4550 (N_4550,N_4488,N_4482);
nand U4551 (N_4551,N_4442,N_4495);
or U4552 (N_4552,N_4490,N_4474);
or U4553 (N_4553,N_4487,N_4485);
nor U4554 (N_4554,N_4443,N_4432);
nand U4555 (N_4555,N_4461,N_4403);
nor U4556 (N_4556,N_4448,N_4426);
or U4557 (N_4557,N_4445,N_4427);
nand U4558 (N_4558,N_4428,N_4439);
xnor U4559 (N_4559,N_4416,N_4470);
nor U4560 (N_4560,N_4432,N_4412);
nor U4561 (N_4561,N_4463,N_4499);
nor U4562 (N_4562,N_4498,N_4486);
nand U4563 (N_4563,N_4402,N_4446);
xnor U4564 (N_4564,N_4494,N_4483);
or U4565 (N_4565,N_4434,N_4470);
or U4566 (N_4566,N_4490,N_4463);
nand U4567 (N_4567,N_4482,N_4489);
nor U4568 (N_4568,N_4438,N_4461);
nor U4569 (N_4569,N_4433,N_4424);
nand U4570 (N_4570,N_4471,N_4462);
nand U4571 (N_4571,N_4491,N_4458);
nand U4572 (N_4572,N_4474,N_4403);
xnor U4573 (N_4573,N_4401,N_4457);
xnor U4574 (N_4574,N_4478,N_4486);
or U4575 (N_4575,N_4430,N_4460);
or U4576 (N_4576,N_4435,N_4405);
and U4577 (N_4577,N_4435,N_4489);
and U4578 (N_4578,N_4435,N_4418);
and U4579 (N_4579,N_4415,N_4450);
xnor U4580 (N_4580,N_4400,N_4483);
and U4581 (N_4581,N_4432,N_4464);
or U4582 (N_4582,N_4426,N_4408);
xor U4583 (N_4583,N_4429,N_4448);
and U4584 (N_4584,N_4497,N_4436);
or U4585 (N_4585,N_4455,N_4494);
or U4586 (N_4586,N_4403,N_4434);
nand U4587 (N_4587,N_4441,N_4491);
nand U4588 (N_4588,N_4427,N_4474);
xor U4589 (N_4589,N_4432,N_4473);
nor U4590 (N_4590,N_4410,N_4492);
nand U4591 (N_4591,N_4430,N_4414);
xor U4592 (N_4592,N_4433,N_4446);
nor U4593 (N_4593,N_4451,N_4444);
nor U4594 (N_4594,N_4476,N_4496);
or U4595 (N_4595,N_4409,N_4453);
and U4596 (N_4596,N_4466,N_4489);
nor U4597 (N_4597,N_4416,N_4459);
xor U4598 (N_4598,N_4406,N_4466);
xnor U4599 (N_4599,N_4465,N_4490);
nor U4600 (N_4600,N_4519,N_4580);
xnor U4601 (N_4601,N_4521,N_4551);
xor U4602 (N_4602,N_4575,N_4587);
nand U4603 (N_4603,N_4511,N_4569);
and U4604 (N_4604,N_4538,N_4531);
or U4605 (N_4605,N_4566,N_4527);
nand U4606 (N_4606,N_4568,N_4582);
and U4607 (N_4607,N_4516,N_4530);
xnor U4608 (N_4608,N_4505,N_4594);
nor U4609 (N_4609,N_4513,N_4560);
xor U4610 (N_4610,N_4549,N_4528);
xor U4611 (N_4611,N_4535,N_4576);
or U4612 (N_4612,N_4567,N_4509);
nor U4613 (N_4613,N_4507,N_4593);
nand U4614 (N_4614,N_4585,N_4537);
or U4615 (N_4615,N_4596,N_4597);
nand U4616 (N_4616,N_4591,N_4583);
and U4617 (N_4617,N_4573,N_4548);
and U4618 (N_4618,N_4559,N_4588);
or U4619 (N_4619,N_4578,N_4504);
and U4620 (N_4620,N_4502,N_4540);
or U4621 (N_4621,N_4541,N_4554);
xor U4622 (N_4622,N_4552,N_4544);
nand U4623 (N_4623,N_4561,N_4550);
xnor U4624 (N_4624,N_4553,N_4525);
and U4625 (N_4625,N_4565,N_4508);
or U4626 (N_4626,N_4574,N_4500);
nor U4627 (N_4627,N_4598,N_4546);
xnor U4628 (N_4628,N_4526,N_4517);
or U4629 (N_4629,N_4503,N_4514);
xnor U4630 (N_4630,N_4555,N_4510);
or U4631 (N_4631,N_4563,N_4572);
xnor U4632 (N_4632,N_4558,N_4520);
nor U4633 (N_4633,N_4547,N_4562);
nand U4634 (N_4634,N_4532,N_4556);
and U4635 (N_4635,N_4518,N_4586);
nor U4636 (N_4636,N_4599,N_4524);
nor U4637 (N_4637,N_4589,N_4534);
or U4638 (N_4638,N_4577,N_4506);
nor U4639 (N_4639,N_4545,N_4515);
or U4640 (N_4640,N_4536,N_4539);
xnor U4641 (N_4641,N_4512,N_4501);
nor U4642 (N_4642,N_4592,N_4529);
and U4643 (N_4643,N_4533,N_4542);
and U4644 (N_4644,N_4564,N_4570);
xnor U4645 (N_4645,N_4522,N_4579);
xor U4646 (N_4646,N_4584,N_4523);
xor U4647 (N_4647,N_4543,N_4581);
and U4648 (N_4648,N_4595,N_4571);
nand U4649 (N_4649,N_4590,N_4557);
or U4650 (N_4650,N_4571,N_4535);
xor U4651 (N_4651,N_4533,N_4582);
or U4652 (N_4652,N_4597,N_4538);
nor U4653 (N_4653,N_4521,N_4561);
xor U4654 (N_4654,N_4524,N_4511);
or U4655 (N_4655,N_4552,N_4571);
nand U4656 (N_4656,N_4597,N_4514);
nand U4657 (N_4657,N_4530,N_4562);
or U4658 (N_4658,N_4535,N_4565);
nand U4659 (N_4659,N_4564,N_4541);
xnor U4660 (N_4660,N_4546,N_4597);
nand U4661 (N_4661,N_4521,N_4537);
and U4662 (N_4662,N_4563,N_4570);
or U4663 (N_4663,N_4563,N_4557);
or U4664 (N_4664,N_4598,N_4560);
nand U4665 (N_4665,N_4541,N_4579);
xnor U4666 (N_4666,N_4579,N_4530);
and U4667 (N_4667,N_4550,N_4547);
or U4668 (N_4668,N_4595,N_4593);
or U4669 (N_4669,N_4599,N_4578);
xor U4670 (N_4670,N_4526,N_4582);
and U4671 (N_4671,N_4556,N_4558);
and U4672 (N_4672,N_4548,N_4554);
nand U4673 (N_4673,N_4510,N_4578);
nand U4674 (N_4674,N_4537,N_4562);
nand U4675 (N_4675,N_4539,N_4522);
xor U4676 (N_4676,N_4516,N_4576);
nand U4677 (N_4677,N_4574,N_4558);
and U4678 (N_4678,N_4540,N_4548);
xor U4679 (N_4679,N_4550,N_4562);
xor U4680 (N_4680,N_4534,N_4512);
and U4681 (N_4681,N_4531,N_4544);
xnor U4682 (N_4682,N_4541,N_4558);
nand U4683 (N_4683,N_4584,N_4514);
or U4684 (N_4684,N_4503,N_4533);
or U4685 (N_4685,N_4502,N_4566);
xor U4686 (N_4686,N_4509,N_4547);
xnor U4687 (N_4687,N_4508,N_4546);
xor U4688 (N_4688,N_4588,N_4522);
or U4689 (N_4689,N_4537,N_4551);
or U4690 (N_4690,N_4588,N_4528);
nor U4691 (N_4691,N_4582,N_4583);
xor U4692 (N_4692,N_4520,N_4556);
nor U4693 (N_4693,N_4546,N_4544);
and U4694 (N_4694,N_4556,N_4531);
xnor U4695 (N_4695,N_4589,N_4568);
xnor U4696 (N_4696,N_4598,N_4518);
xnor U4697 (N_4697,N_4587,N_4569);
nor U4698 (N_4698,N_4528,N_4577);
and U4699 (N_4699,N_4553,N_4521);
xnor U4700 (N_4700,N_4690,N_4669);
nand U4701 (N_4701,N_4695,N_4624);
xnor U4702 (N_4702,N_4648,N_4680);
nor U4703 (N_4703,N_4611,N_4620);
xor U4704 (N_4704,N_4638,N_4697);
or U4705 (N_4705,N_4677,N_4654);
nor U4706 (N_4706,N_4676,N_4653);
nor U4707 (N_4707,N_4686,N_4612);
nor U4708 (N_4708,N_4627,N_4601);
xor U4709 (N_4709,N_4658,N_4687);
nor U4710 (N_4710,N_4639,N_4636);
nand U4711 (N_4711,N_4643,N_4619);
nor U4712 (N_4712,N_4683,N_4659);
nand U4713 (N_4713,N_4657,N_4688);
or U4714 (N_4714,N_4663,N_4685);
nor U4715 (N_4715,N_4692,N_4649);
and U4716 (N_4716,N_4684,N_4641);
nor U4717 (N_4717,N_4610,N_4629);
and U4718 (N_4718,N_4630,N_4655);
and U4719 (N_4719,N_4660,N_4626);
nor U4720 (N_4720,N_4651,N_4696);
nor U4721 (N_4721,N_4614,N_4664);
or U4722 (N_4722,N_4602,N_4600);
xor U4723 (N_4723,N_4666,N_4640);
or U4724 (N_4724,N_4665,N_4622);
or U4725 (N_4725,N_4662,N_4644);
nor U4726 (N_4726,N_4615,N_4691);
or U4727 (N_4727,N_4642,N_4632);
or U4728 (N_4728,N_4667,N_4693);
nor U4729 (N_4729,N_4679,N_4661);
or U4730 (N_4730,N_4606,N_4608);
and U4731 (N_4731,N_4625,N_4674);
nor U4732 (N_4732,N_4670,N_4650);
and U4733 (N_4733,N_4689,N_4623);
and U4734 (N_4734,N_4678,N_4652);
xor U4735 (N_4735,N_4609,N_4672);
xnor U4736 (N_4736,N_4635,N_4628);
or U4737 (N_4737,N_4656,N_4618);
and U4738 (N_4738,N_4675,N_4617);
and U4739 (N_4739,N_4637,N_4647);
xor U4740 (N_4740,N_4673,N_4604);
or U4741 (N_4741,N_4633,N_4621);
and U4742 (N_4742,N_4699,N_4616);
nand U4743 (N_4743,N_4646,N_4698);
or U4744 (N_4744,N_4671,N_4668);
or U4745 (N_4745,N_4645,N_4634);
nor U4746 (N_4746,N_4607,N_4694);
nand U4747 (N_4747,N_4681,N_4605);
nor U4748 (N_4748,N_4603,N_4631);
xor U4749 (N_4749,N_4682,N_4613);
xnor U4750 (N_4750,N_4651,N_4680);
xnor U4751 (N_4751,N_4631,N_4646);
nor U4752 (N_4752,N_4651,N_4646);
and U4753 (N_4753,N_4694,N_4645);
xor U4754 (N_4754,N_4634,N_4641);
xor U4755 (N_4755,N_4656,N_4643);
or U4756 (N_4756,N_4651,N_4626);
and U4757 (N_4757,N_4681,N_4685);
and U4758 (N_4758,N_4668,N_4642);
xnor U4759 (N_4759,N_4606,N_4662);
nor U4760 (N_4760,N_4649,N_4650);
xnor U4761 (N_4761,N_4621,N_4609);
or U4762 (N_4762,N_4683,N_4654);
nand U4763 (N_4763,N_4673,N_4637);
or U4764 (N_4764,N_4653,N_4684);
xnor U4765 (N_4765,N_4697,N_4600);
or U4766 (N_4766,N_4630,N_4677);
or U4767 (N_4767,N_4634,N_4608);
and U4768 (N_4768,N_4632,N_4679);
and U4769 (N_4769,N_4695,N_4666);
nor U4770 (N_4770,N_4674,N_4629);
or U4771 (N_4771,N_4681,N_4655);
xnor U4772 (N_4772,N_4688,N_4632);
nand U4773 (N_4773,N_4661,N_4643);
nand U4774 (N_4774,N_4648,N_4632);
nand U4775 (N_4775,N_4626,N_4653);
or U4776 (N_4776,N_4647,N_4629);
or U4777 (N_4777,N_4642,N_4667);
nand U4778 (N_4778,N_4633,N_4602);
nand U4779 (N_4779,N_4677,N_4627);
or U4780 (N_4780,N_4632,N_4698);
nor U4781 (N_4781,N_4602,N_4601);
xnor U4782 (N_4782,N_4609,N_4657);
or U4783 (N_4783,N_4659,N_4692);
xor U4784 (N_4784,N_4644,N_4653);
xnor U4785 (N_4785,N_4675,N_4671);
and U4786 (N_4786,N_4601,N_4619);
and U4787 (N_4787,N_4699,N_4697);
nand U4788 (N_4788,N_4637,N_4667);
nor U4789 (N_4789,N_4632,N_4634);
xnor U4790 (N_4790,N_4617,N_4690);
nand U4791 (N_4791,N_4690,N_4639);
nand U4792 (N_4792,N_4688,N_4611);
and U4793 (N_4793,N_4602,N_4697);
nand U4794 (N_4794,N_4650,N_4618);
or U4795 (N_4795,N_4642,N_4657);
xor U4796 (N_4796,N_4633,N_4608);
nand U4797 (N_4797,N_4698,N_4656);
xnor U4798 (N_4798,N_4687,N_4647);
or U4799 (N_4799,N_4664,N_4659);
xor U4800 (N_4800,N_4766,N_4724);
or U4801 (N_4801,N_4785,N_4744);
nand U4802 (N_4802,N_4757,N_4734);
nor U4803 (N_4803,N_4726,N_4715);
nor U4804 (N_4804,N_4725,N_4768);
xnor U4805 (N_4805,N_4794,N_4771);
and U4806 (N_4806,N_4769,N_4780);
or U4807 (N_4807,N_4739,N_4707);
xor U4808 (N_4808,N_4776,N_4732);
nor U4809 (N_4809,N_4751,N_4772);
and U4810 (N_4810,N_4755,N_4763);
xor U4811 (N_4811,N_4798,N_4741);
or U4812 (N_4812,N_4719,N_4778);
nor U4813 (N_4813,N_4752,N_4703);
nor U4814 (N_4814,N_4765,N_4754);
xor U4815 (N_4815,N_4711,N_4756);
and U4816 (N_4816,N_4791,N_4745);
and U4817 (N_4817,N_4782,N_4721);
and U4818 (N_4818,N_4781,N_4784);
nand U4819 (N_4819,N_4738,N_4789);
nor U4820 (N_4820,N_4723,N_4701);
and U4821 (N_4821,N_4742,N_4767);
xor U4822 (N_4822,N_4720,N_4722);
nor U4823 (N_4823,N_4760,N_4728);
xor U4824 (N_4824,N_4758,N_4748);
xnor U4825 (N_4825,N_4717,N_4786);
and U4826 (N_4826,N_4777,N_4799);
xor U4827 (N_4827,N_4783,N_4774);
nand U4828 (N_4828,N_4796,N_4749);
nand U4829 (N_4829,N_4792,N_4716);
nor U4830 (N_4830,N_4790,N_4729);
xnor U4831 (N_4831,N_4704,N_4773);
or U4832 (N_4832,N_4797,N_4736);
xnor U4833 (N_4833,N_4714,N_4700);
xor U4834 (N_4834,N_4746,N_4753);
or U4835 (N_4835,N_4727,N_4708);
or U4836 (N_4836,N_4762,N_4710);
or U4837 (N_4837,N_4737,N_4759);
nor U4838 (N_4838,N_4743,N_4733);
or U4839 (N_4839,N_4793,N_4775);
and U4840 (N_4840,N_4788,N_4747);
and U4841 (N_4841,N_4709,N_4706);
xor U4842 (N_4842,N_4718,N_4787);
or U4843 (N_4843,N_4735,N_4764);
xnor U4844 (N_4844,N_4731,N_4730);
nor U4845 (N_4845,N_4713,N_4712);
nand U4846 (N_4846,N_4779,N_4770);
and U4847 (N_4847,N_4705,N_4761);
and U4848 (N_4848,N_4740,N_4702);
nor U4849 (N_4849,N_4750,N_4795);
xor U4850 (N_4850,N_4734,N_4728);
nor U4851 (N_4851,N_4780,N_4708);
or U4852 (N_4852,N_4704,N_4746);
nand U4853 (N_4853,N_4780,N_4730);
and U4854 (N_4854,N_4732,N_4707);
or U4855 (N_4855,N_4777,N_4790);
nand U4856 (N_4856,N_4765,N_4748);
nand U4857 (N_4857,N_4777,N_4733);
xnor U4858 (N_4858,N_4747,N_4750);
nand U4859 (N_4859,N_4723,N_4700);
nand U4860 (N_4860,N_4723,N_4705);
or U4861 (N_4861,N_4728,N_4757);
and U4862 (N_4862,N_4734,N_4781);
and U4863 (N_4863,N_4715,N_4799);
nor U4864 (N_4864,N_4768,N_4793);
xnor U4865 (N_4865,N_4722,N_4708);
and U4866 (N_4866,N_4773,N_4744);
and U4867 (N_4867,N_4792,N_4731);
nand U4868 (N_4868,N_4718,N_4793);
nand U4869 (N_4869,N_4770,N_4710);
nor U4870 (N_4870,N_4792,N_4752);
nand U4871 (N_4871,N_4753,N_4700);
nor U4872 (N_4872,N_4776,N_4780);
xor U4873 (N_4873,N_4768,N_4704);
or U4874 (N_4874,N_4760,N_4733);
xnor U4875 (N_4875,N_4756,N_4777);
nand U4876 (N_4876,N_4743,N_4717);
nor U4877 (N_4877,N_4765,N_4764);
and U4878 (N_4878,N_4706,N_4738);
nor U4879 (N_4879,N_4792,N_4798);
nand U4880 (N_4880,N_4793,N_4786);
nor U4881 (N_4881,N_4744,N_4736);
nand U4882 (N_4882,N_4761,N_4786);
and U4883 (N_4883,N_4773,N_4751);
or U4884 (N_4884,N_4794,N_4727);
and U4885 (N_4885,N_4751,N_4739);
nand U4886 (N_4886,N_4733,N_4721);
or U4887 (N_4887,N_4779,N_4750);
and U4888 (N_4888,N_4729,N_4798);
and U4889 (N_4889,N_4782,N_4717);
or U4890 (N_4890,N_4795,N_4772);
xor U4891 (N_4891,N_4773,N_4774);
nand U4892 (N_4892,N_4716,N_4741);
nand U4893 (N_4893,N_4716,N_4750);
xnor U4894 (N_4894,N_4752,N_4751);
xor U4895 (N_4895,N_4771,N_4769);
and U4896 (N_4896,N_4784,N_4736);
and U4897 (N_4897,N_4770,N_4790);
nand U4898 (N_4898,N_4703,N_4784);
or U4899 (N_4899,N_4788,N_4748);
and U4900 (N_4900,N_4801,N_4839);
xnor U4901 (N_4901,N_4842,N_4802);
xnor U4902 (N_4902,N_4862,N_4858);
xnor U4903 (N_4903,N_4844,N_4882);
nand U4904 (N_4904,N_4857,N_4825);
and U4905 (N_4905,N_4856,N_4833);
or U4906 (N_4906,N_4828,N_4838);
or U4907 (N_4907,N_4840,N_4818);
xnor U4908 (N_4908,N_4873,N_4837);
xnor U4909 (N_4909,N_4867,N_4861);
nor U4910 (N_4910,N_4822,N_4860);
nor U4911 (N_4911,N_4859,N_4863);
or U4912 (N_4912,N_4865,N_4881);
xnor U4913 (N_4913,N_4811,N_4812);
or U4914 (N_4914,N_4897,N_4866);
or U4915 (N_4915,N_4834,N_4829);
xnor U4916 (N_4916,N_4896,N_4852);
nand U4917 (N_4917,N_4823,N_4813);
nor U4918 (N_4918,N_4898,N_4864);
and U4919 (N_4919,N_4846,N_4819);
xor U4920 (N_4920,N_4890,N_4826);
or U4921 (N_4921,N_4894,N_4830);
and U4922 (N_4922,N_4885,N_4804);
or U4923 (N_4923,N_4879,N_4831);
nor U4924 (N_4924,N_4899,N_4835);
nand U4925 (N_4925,N_4806,N_4853);
or U4926 (N_4926,N_4871,N_4850);
nor U4927 (N_4927,N_4843,N_4887);
xor U4928 (N_4928,N_4816,N_4886);
nand U4929 (N_4929,N_4889,N_4832);
or U4930 (N_4930,N_4817,N_4809);
nor U4931 (N_4931,N_4895,N_4888);
nand U4932 (N_4932,N_4810,N_4851);
nand U4933 (N_4933,N_4876,N_4807);
nand U4934 (N_4934,N_4870,N_4827);
and U4935 (N_4935,N_4893,N_4814);
xnor U4936 (N_4936,N_4847,N_4878);
nor U4937 (N_4937,N_4848,N_4883);
xor U4938 (N_4938,N_4820,N_4880);
nand U4939 (N_4939,N_4815,N_4824);
or U4940 (N_4940,N_4803,N_4874);
nor U4941 (N_4941,N_4800,N_4849);
nand U4942 (N_4942,N_4854,N_4877);
nand U4943 (N_4943,N_4892,N_4891);
xnor U4944 (N_4944,N_4805,N_4855);
xor U4945 (N_4945,N_4808,N_4821);
or U4946 (N_4946,N_4872,N_4836);
nand U4947 (N_4947,N_4868,N_4869);
nor U4948 (N_4948,N_4875,N_4845);
nor U4949 (N_4949,N_4884,N_4841);
nand U4950 (N_4950,N_4817,N_4884);
nand U4951 (N_4951,N_4833,N_4895);
nand U4952 (N_4952,N_4894,N_4821);
nand U4953 (N_4953,N_4878,N_4843);
nor U4954 (N_4954,N_4817,N_4893);
and U4955 (N_4955,N_4891,N_4894);
or U4956 (N_4956,N_4871,N_4894);
or U4957 (N_4957,N_4842,N_4888);
and U4958 (N_4958,N_4832,N_4860);
nor U4959 (N_4959,N_4827,N_4876);
nand U4960 (N_4960,N_4851,N_4886);
nand U4961 (N_4961,N_4820,N_4807);
or U4962 (N_4962,N_4837,N_4840);
xnor U4963 (N_4963,N_4812,N_4879);
xor U4964 (N_4964,N_4898,N_4835);
or U4965 (N_4965,N_4801,N_4846);
and U4966 (N_4966,N_4896,N_4886);
xor U4967 (N_4967,N_4888,N_4830);
and U4968 (N_4968,N_4813,N_4881);
nand U4969 (N_4969,N_4809,N_4859);
xor U4970 (N_4970,N_4896,N_4895);
xnor U4971 (N_4971,N_4860,N_4886);
and U4972 (N_4972,N_4892,N_4858);
and U4973 (N_4973,N_4806,N_4854);
and U4974 (N_4974,N_4813,N_4844);
xor U4975 (N_4975,N_4897,N_4851);
and U4976 (N_4976,N_4881,N_4800);
xor U4977 (N_4977,N_4800,N_4806);
or U4978 (N_4978,N_4824,N_4892);
or U4979 (N_4979,N_4824,N_4897);
nor U4980 (N_4980,N_4891,N_4884);
or U4981 (N_4981,N_4856,N_4845);
and U4982 (N_4982,N_4847,N_4814);
xor U4983 (N_4983,N_4895,N_4887);
nor U4984 (N_4984,N_4841,N_4894);
xnor U4985 (N_4985,N_4802,N_4832);
and U4986 (N_4986,N_4891,N_4869);
nand U4987 (N_4987,N_4896,N_4826);
and U4988 (N_4988,N_4802,N_4852);
xor U4989 (N_4989,N_4826,N_4803);
nand U4990 (N_4990,N_4822,N_4819);
xnor U4991 (N_4991,N_4851,N_4871);
and U4992 (N_4992,N_4855,N_4801);
and U4993 (N_4993,N_4883,N_4853);
nand U4994 (N_4994,N_4817,N_4832);
and U4995 (N_4995,N_4804,N_4819);
nor U4996 (N_4996,N_4821,N_4838);
xor U4997 (N_4997,N_4822,N_4855);
nand U4998 (N_4998,N_4803,N_4819);
nor U4999 (N_4999,N_4814,N_4881);
xor UO_0 (O_0,N_4926,N_4941);
xor UO_1 (O_1,N_4978,N_4969);
nor UO_2 (O_2,N_4939,N_4971);
nand UO_3 (O_3,N_4919,N_4985);
nand UO_4 (O_4,N_4987,N_4995);
xnor UO_5 (O_5,N_4942,N_4960);
xor UO_6 (O_6,N_4902,N_4907);
or UO_7 (O_7,N_4948,N_4992);
nor UO_8 (O_8,N_4927,N_4972);
nand UO_9 (O_9,N_4909,N_4991);
xor UO_10 (O_10,N_4957,N_4940);
nor UO_11 (O_11,N_4914,N_4923);
xnor UO_12 (O_12,N_4951,N_4901);
nand UO_13 (O_13,N_4982,N_4928);
or UO_14 (O_14,N_4958,N_4936);
or UO_15 (O_15,N_4917,N_4952);
or UO_16 (O_16,N_4915,N_4916);
and UO_17 (O_17,N_4967,N_4906);
xor UO_18 (O_18,N_4988,N_4999);
nand UO_19 (O_19,N_4908,N_4932);
nor UO_20 (O_20,N_4946,N_4955);
and UO_21 (O_21,N_4997,N_4938);
xor UO_22 (O_22,N_4953,N_4924);
nand UO_23 (O_23,N_4912,N_4961);
or UO_24 (O_24,N_4983,N_4954);
nand UO_25 (O_25,N_4975,N_4973);
xor UO_26 (O_26,N_4943,N_4947);
and UO_27 (O_27,N_4937,N_4931);
nor UO_28 (O_28,N_4986,N_4996);
nand UO_29 (O_29,N_4920,N_4993);
or UO_30 (O_30,N_4903,N_4959);
nand UO_31 (O_31,N_4966,N_4935);
nor UO_32 (O_32,N_4984,N_4900);
nor UO_33 (O_33,N_4968,N_4994);
and UO_34 (O_34,N_4944,N_4964);
nor UO_35 (O_35,N_4911,N_4913);
and UO_36 (O_36,N_4998,N_4904);
nand UO_37 (O_37,N_4979,N_4925);
and UO_38 (O_38,N_4962,N_4989);
nand UO_39 (O_39,N_4929,N_4930);
nor UO_40 (O_40,N_4981,N_4976);
and UO_41 (O_41,N_4905,N_4910);
nor UO_42 (O_42,N_4922,N_4974);
or UO_43 (O_43,N_4918,N_4977);
nand UO_44 (O_44,N_4990,N_4980);
nand UO_45 (O_45,N_4956,N_4970);
nor UO_46 (O_46,N_4965,N_4934);
or UO_47 (O_47,N_4933,N_4945);
and UO_48 (O_48,N_4950,N_4963);
nor UO_49 (O_49,N_4921,N_4949);
nor UO_50 (O_50,N_4928,N_4931);
or UO_51 (O_51,N_4937,N_4959);
and UO_52 (O_52,N_4963,N_4902);
nand UO_53 (O_53,N_4909,N_4976);
xnor UO_54 (O_54,N_4957,N_4996);
nand UO_55 (O_55,N_4910,N_4925);
nand UO_56 (O_56,N_4986,N_4945);
xnor UO_57 (O_57,N_4973,N_4935);
nor UO_58 (O_58,N_4979,N_4927);
or UO_59 (O_59,N_4932,N_4900);
xor UO_60 (O_60,N_4931,N_4935);
nor UO_61 (O_61,N_4960,N_4902);
or UO_62 (O_62,N_4967,N_4964);
or UO_63 (O_63,N_4926,N_4903);
or UO_64 (O_64,N_4988,N_4954);
xnor UO_65 (O_65,N_4952,N_4991);
nand UO_66 (O_66,N_4954,N_4957);
and UO_67 (O_67,N_4928,N_4968);
nand UO_68 (O_68,N_4998,N_4926);
xnor UO_69 (O_69,N_4986,N_4987);
xnor UO_70 (O_70,N_4953,N_4949);
and UO_71 (O_71,N_4967,N_4936);
xor UO_72 (O_72,N_4909,N_4974);
nand UO_73 (O_73,N_4966,N_4929);
nor UO_74 (O_74,N_4900,N_4997);
nor UO_75 (O_75,N_4932,N_4982);
or UO_76 (O_76,N_4947,N_4978);
and UO_77 (O_77,N_4993,N_4996);
or UO_78 (O_78,N_4927,N_4987);
nor UO_79 (O_79,N_4947,N_4914);
and UO_80 (O_80,N_4933,N_4971);
xnor UO_81 (O_81,N_4965,N_4933);
and UO_82 (O_82,N_4986,N_4939);
and UO_83 (O_83,N_4999,N_4914);
xor UO_84 (O_84,N_4945,N_4925);
and UO_85 (O_85,N_4957,N_4969);
and UO_86 (O_86,N_4936,N_4907);
or UO_87 (O_87,N_4924,N_4999);
nand UO_88 (O_88,N_4965,N_4902);
xor UO_89 (O_89,N_4997,N_4905);
and UO_90 (O_90,N_4939,N_4996);
or UO_91 (O_91,N_4938,N_4942);
and UO_92 (O_92,N_4918,N_4908);
xnor UO_93 (O_93,N_4913,N_4967);
and UO_94 (O_94,N_4916,N_4997);
nand UO_95 (O_95,N_4912,N_4968);
nand UO_96 (O_96,N_4929,N_4993);
or UO_97 (O_97,N_4952,N_4940);
xnor UO_98 (O_98,N_4946,N_4985);
or UO_99 (O_99,N_4998,N_4957);
nor UO_100 (O_100,N_4977,N_4980);
nand UO_101 (O_101,N_4970,N_4931);
and UO_102 (O_102,N_4930,N_4935);
xnor UO_103 (O_103,N_4929,N_4900);
or UO_104 (O_104,N_4940,N_4956);
and UO_105 (O_105,N_4973,N_4917);
nand UO_106 (O_106,N_4906,N_4951);
nor UO_107 (O_107,N_4948,N_4924);
or UO_108 (O_108,N_4902,N_4920);
or UO_109 (O_109,N_4961,N_4974);
nor UO_110 (O_110,N_4943,N_4967);
or UO_111 (O_111,N_4900,N_4905);
or UO_112 (O_112,N_4921,N_4930);
or UO_113 (O_113,N_4932,N_4965);
xor UO_114 (O_114,N_4930,N_4966);
or UO_115 (O_115,N_4931,N_4968);
and UO_116 (O_116,N_4958,N_4974);
xor UO_117 (O_117,N_4988,N_4941);
and UO_118 (O_118,N_4904,N_4938);
xnor UO_119 (O_119,N_4947,N_4961);
or UO_120 (O_120,N_4951,N_4936);
or UO_121 (O_121,N_4959,N_4931);
and UO_122 (O_122,N_4989,N_4983);
nand UO_123 (O_123,N_4901,N_4992);
nand UO_124 (O_124,N_4912,N_4906);
or UO_125 (O_125,N_4973,N_4930);
xnor UO_126 (O_126,N_4968,N_4935);
nor UO_127 (O_127,N_4947,N_4908);
and UO_128 (O_128,N_4901,N_4963);
and UO_129 (O_129,N_4909,N_4914);
or UO_130 (O_130,N_4942,N_4950);
nand UO_131 (O_131,N_4937,N_4929);
and UO_132 (O_132,N_4992,N_4931);
xor UO_133 (O_133,N_4986,N_4985);
xnor UO_134 (O_134,N_4994,N_4954);
nor UO_135 (O_135,N_4952,N_4987);
xnor UO_136 (O_136,N_4941,N_4992);
or UO_137 (O_137,N_4964,N_4991);
xnor UO_138 (O_138,N_4971,N_4966);
and UO_139 (O_139,N_4926,N_4984);
and UO_140 (O_140,N_4982,N_4956);
xnor UO_141 (O_141,N_4979,N_4969);
nor UO_142 (O_142,N_4989,N_4904);
and UO_143 (O_143,N_4999,N_4919);
xor UO_144 (O_144,N_4900,N_4909);
and UO_145 (O_145,N_4933,N_4992);
xnor UO_146 (O_146,N_4959,N_4966);
xnor UO_147 (O_147,N_4961,N_4939);
nor UO_148 (O_148,N_4999,N_4948);
or UO_149 (O_149,N_4999,N_4954);
nor UO_150 (O_150,N_4942,N_4920);
xor UO_151 (O_151,N_4992,N_4928);
and UO_152 (O_152,N_4937,N_4924);
nand UO_153 (O_153,N_4917,N_4911);
xnor UO_154 (O_154,N_4990,N_4973);
nor UO_155 (O_155,N_4961,N_4955);
or UO_156 (O_156,N_4997,N_4930);
xor UO_157 (O_157,N_4978,N_4946);
and UO_158 (O_158,N_4907,N_4922);
and UO_159 (O_159,N_4956,N_4968);
xor UO_160 (O_160,N_4960,N_4933);
xor UO_161 (O_161,N_4935,N_4912);
or UO_162 (O_162,N_4932,N_4969);
xnor UO_163 (O_163,N_4989,N_4986);
and UO_164 (O_164,N_4904,N_4911);
nor UO_165 (O_165,N_4988,N_4918);
nor UO_166 (O_166,N_4951,N_4908);
or UO_167 (O_167,N_4989,N_4991);
xor UO_168 (O_168,N_4919,N_4913);
or UO_169 (O_169,N_4935,N_4961);
nand UO_170 (O_170,N_4908,N_4991);
or UO_171 (O_171,N_4992,N_4918);
or UO_172 (O_172,N_4927,N_4995);
nand UO_173 (O_173,N_4925,N_4902);
or UO_174 (O_174,N_4927,N_4933);
xnor UO_175 (O_175,N_4916,N_4942);
and UO_176 (O_176,N_4936,N_4933);
or UO_177 (O_177,N_4946,N_4982);
or UO_178 (O_178,N_4948,N_4915);
nor UO_179 (O_179,N_4923,N_4928);
nand UO_180 (O_180,N_4953,N_4976);
nand UO_181 (O_181,N_4943,N_4936);
nor UO_182 (O_182,N_4949,N_4943);
nor UO_183 (O_183,N_4938,N_4924);
nand UO_184 (O_184,N_4923,N_4995);
xor UO_185 (O_185,N_4911,N_4980);
xnor UO_186 (O_186,N_4994,N_4974);
nand UO_187 (O_187,N_4984,N_4974);
nor UO_188 (O_188,N_4920,N_4984);
or UO_189 (O_189,N_4961,N_4926);
xor UO_190 (O_190,N_4948,N_4978);
or UO_191 (O_191,N_4990,N_4981);
nand UO_192 (O_192,N_4999,N_4994);
or UO_193 (O_193,N_4953,N_4911);
or UO_194 (O_194,N_4954,N_4900);
and UO_195 (O_195,N_4971,N_4977);
nor UO_196 (O_196,N_4986,N_4930);
xor UO_197 (O_197,N_4966,N_4992);
and UO_198 (O_198,N_4929,N_4996);
nor UO_199 (O_199,N_4956,N_4977);
nand UO_200 (O_200,N_4953,N_4970);
nand UO_201 (O_201,N_4962,N_4953);
nand UO_202 (O_202,N_4968,N_4983);
xnor UO_203 (O_203,N_4961,N_4938);
or UO_204 (O_204,N_4940,N_4936);
nor UO_205 (O_205,N_4995,N_4973);
or UO_206 (O_206,N_4912,N_4951);
xnor UO_207 (O_207,N_4968,N_4903);
and UO_208 (O_208,N_4976,N_4944);
xor UO_209 (O_209,N_4982,N_4930);
and UO_210 (O_210,N_4956,N_4988);
xor UO_211 (O_211,N_4953,N_4995);
and UO_212 (O_212,N_4959,N_4944);
and UO_213 (O_213,N_4917,N_4977);
xor UO_214 (O_214,N_4939,N_4932);
nor UO_215 (O_215,N_4913,N_4988);
nand UO_216 (O_216,N_4956,N_4954);
nor UO_217 (O_217,N_4981,N_4930);
nor UO_218 (O_218,N_4914,N_4981);
xnor UO_219 (O_219,N_4924,N_4920);
xnor UO_220 (O_220,N_4930,N_4995);
xnor UO_221 (O_221,N_4949,N_4995);
or UO_222 (O_222,N_4918,N_4957);
nand UO_223 (O_223,N_4959,N_4921);
nand UO_224 (O_224,N_4902,N_4997);
nor UO_225 (O_225,N_4997,N_4908);
xor UO_226 (O_226,N_4921,N_4906);
nor UO_227 (O_227,N_4911,N_4984);
xor UO_228 (O_228,N_4953,N_4923);
or UO_229 (O_229,N_4994,N_4941);
nor UO_230 (O_230,N_4913,N_4924);
nor UO_231 (O_231,N_4916,N_4927);
and UO_232 (O_232,N_4977,N_4997);
or UO_233 (O_233,N_4957,N_4901);
nand UO_234 (O_234,N_4917,N_4994);
nand UO_235 (O_235,N_4975,N_4997);
xnor UO_236 (O_236,N_4923,N_4915);
nand UO_237 (O_237,N_4902,N_4946);
nand UO_238 (O_238,N_4904,N_4905);
nor UO_239 (O_239,N_4906,N_4966);
or UO_240 (O_240,N_4963,N_4939);
nand UO_241 (O_241,N_4936,N_4971);
nor UO_242 (O_242,N_4952,N_4913);
nor UO_243 (O_243,N_4921,N_4916);
nor UO_244 (O_244,N_4935,N_4932);
and UO_245 (O_245,N_4920,N_4966);
nor UO_246 (O_246,N_4931,N_4906);
nor UO_247 (O_247,N_4989,N_4954);
nor UO_248 (O_248,N_4981,N_4996);
and UO_249 (O_249,N_4972,N_4908);
nor UO_250 (O_250,N_4970,N_4917);
xnor UO_251 (O_251,N_4907,N_4916);
xor UO_252 (O_252,N_4955,N_4976);
nand UO_253 (O_253,N_4917,N_4983);
or UO_254 (O_254,N_4908,N_4980);
and UO_255 (O_255,N_4922,N_4968);
xnor UO_256 (O_256,N_4938,N_4981);
nor UO_257 (O_257,N_4981,N_4932);
xnor UO_258 (O_258,N_4925,N_4997);
or UO_259 (O_259,N_4956,N_4973);
nor UO_260 (O_260,N_4938,N_4909);
nand UO_261 (O_261,N_4935,N_4938);
nand UO_262 (O_262,N_4925,N_4947);
nor UO_263 (O_263,N_4939,N_4926);
or UO_264 (O_264,N_4961,N_4910);
nand UO_265 (O_265,N_4940,N_4960);
or UO_266 (O_266,N_4964,N_4906);
nor UO_267 (O_267,N_4956,N_4983);
or UO_268 (O_268,N_4927,N_4949);
nor UO_269 (O_269,N_4976,N_4908);
nor UO_270 (O_270,N_4982,N_4979);
xnor UO_271 (O_271,N_4905,N_4911);
nand UO_272 (O_272,N_4975,N_4992);
nor UO_273 (O_273,N_4963,N_4966);
xnor UO_274 (O_274,N_4922,N_4989);
or UO_275 (O_275,N_4978,N_4952);
or UO_276 (O_276,N_4923,N_4918);
xor UO_277 (O_277,N_4928,N_4937);
and UO_278 (O_278,N_4971,N_4952);
nor UO_279 (O_279,N_4972,N_4977);
or UO_280 (O_280,N_4959,N_4954);
xnor UO_281 (O_281,N_4949,N_4969);
nor UO_282 (O_282,N_4958,N_4947);
xor UO_283 (O_283,N_4948,N_4918);
nor UO_284 (O_284,N_4982,N_4990);
or UO_285 (O_285,N_4951,N_4949);
xnor UO_286 (O_286,N_4943,N_4985);
nand UO_287 (O_287,N_4978,N_4954);
xnor UO_288 (O_288,N_4944,N_4980);
or UO_289 (O_289,N_4979,N_4951);
xnor UO_290 (O_290,N_4992,N_4953);
or UO_291 (O_291,N_4985,N_4995);
or UO_292 (O_292,N_4981,N_4904);
and UO_293 (O_293,N_4932,N_4918);
xnor UO_294 (O_294,N_4969,N_4910);
or UO_295 (O_295,N_4942,N_4991);
or UO_296 (O_296,N_4972,N_4901);
nor UO_297 (O_297,N_4982,N_4972);
nor UO_298 (O_298,N_4939,N_4911);
xor UO_299 (O_299,N_4967,N_4949);
xnor UO_300 (O_300,N_4914,N_4935);
or UO_301 (O_301,N_4931,N_4986);
nor UO_302 (O_302,N_4955,N_4953);
xor UO_303 (O_303,N_4934,N_4999);
nand UO_304 (O_304,N_4966,N_4923);
or UO_305 (O_305,N_4948,N_4912);
nand UO_306 (O_306,N_4918,N_4999);
nor UO_307 (O_307,N_4911,N_4972);
or UO_308 (O_308,N_4933,N_4937);
nand UO_309 (O_309,N_4924,N_4906);
nor UO_310 (O_310,N_4903,N_4932);
or UO_311 (O_311,N_4954,N_4998);
or UO_312 (O_312,N_4905,N_4962);
and UO_313 (O_313,N_4934,N_4952);
or UO_314 (O_314,N_4914,N_4978);
xnor UO_315 (O_315,N_4982,N_4923);
nor UO_316 (O_316,N_4900,N_4953);
and UO_317 (O_317,N_4910,N_4913);
nor UO_318 (O_318,N_4931,N_4938);
xnor UO_319 (O_319,N_4961,N_4908);
nand UO_320 (O_320,N_4942,N_4998);
nand UO_321 (O_321,N_4959,N_4953);
and UO_322 (O_322,N_4994,N_4900);
or UO_323 (O_323,N_4902,N_4908);
xnor UO_324 (O_324,N_4911,N_4998);
nand UO_325 (O_325,N_4920,N_4962);
or UO_326 (O_326,N_4900,N_4991);
xor UO_327 (O_327,N_4965,N_4989);
nand UO_328 (O_328,N_4924,N_4975);
and UO_329 (O_329,N_4916,N_4995);
and UO_330 (O_330,N_4946,N_4947);
xnor UO_331 (O_331,N_4939,N_4924);
nand UO_332 (O_332,N_4963,N_4952);
or UO_333 (O_333,N_4978,N_4920);
nand UO_334 (O_334,N_4987,N_4912);
xor UO_335 (O_335,N_4968,N_4917);
nand UO_336 (O_336,N_4979,N_4970);
xor UO_337 (O_337,N_4959,N_4941);
or UO_338 (O_338,N_4951,N_4934);
and UO_339 (O_339,N_4976,N_4963);
nand UO_340 (O_340,N_4917,N_4935);
xor UO_341 (O_341,N_4968,N_4915);
nor UO_342 (O_342,N_4916,N_4923);
or UO_343 (O_343,N_4911,N_4957);
nor UO_344 (O_344,N_4919,N_4902);
xnor UO_345 (O_345,N_4936,N_4991);
or UO_346 (O_346,N_4976,N_4924);
nand UO_347 (O_347,N_4919,N_4997);
nor UO_348 (O_348,N_4967,N_4972);
xor UO_349 (O_349,N_4996,N_4946);
and UO_350 (O_350,N_4920,N_4964);
nand UO_351 (O_351,N_4931,N_4974);
nor UO_352 (O_352,N_4967,N_4930);
nand UO_353 (O_353,N_4931,N_4999);
or UO_354 (O_354,N_4956,N_4962);
xnor UO_355 (O_355,N_4946,N_4993);
and UO_356 (O_356,N_4972,N_4947);
nor UO_357 (O_357,N_4978,N_4917);
nor UO_358 (O_358,N_4943,N_4975);
nor UO_359 (O_359,N_4997,N_4904);
xor UO_360 (O_360,N_4942,N_4982);
or UO_361 (O_361,N_4945,N_4963);
or UO_362 (O_362,N_4902,N_4929);
and UO_363 (O_363,N_4984,N_4993);
xnor UO_364 (O_364,N_4981,N_4964);
nor UO_365 (O_365,N_4919,N_4974);
nand UO_366 (O_366,N_4937,N_4900);
xor UO_367 (O_367,N_4991,N_4934);
or UO_368 (O_368,N_4968,N_4909);
nand UO_369 (O_369,N_4942,N_4946);
xnor UO_370 (O_370,N_4912,N_4992);
nor UO_371 (O_371,N_4991,N_4977);
nand UO_372 (O_372,N_4948,N_4961);
xnor UO_373 (O_373,N_4927,N_4977);
nor UO_374 (O_374,N_4992,N_4964);
nor UO_375 (O_375,N_4905,N_4918);
and UO_376 (O_376,N_4921,N_4987);
xnor UO_377 (O_377,N_4950,N_4994);
nand UO_378 (O_378,N_4930,N_4946);
nand UO_379 (O_379,N_4938,N_4937);
nor UO_380 (O_380,N_4922,N_4983);
nand UO_381 (O_381,N_4971,N_4914);
and UO_382 (O_382,N_4980,N_4968);
or UO_383 (O_383,N_4922,N_4919);
nand UO_384 (O_384,N_4912,N_4917);
nor UO_385 (O_385,N_4929,N_4944);
nor UO_386 (O_386,N_4946,N_4972);
nor UO_387 (O_387,N_4972,N_4999);
and UO_388 (O_388,N_4955,N_4974);
nand UO_389 (O_389,N_4991,N_4990);
or UO_390 (O_390,N_4979,N_4976);
xnor UO_391 (O_391,N_4947,N_4904);
and UO_392 (O_392,N_4995,N_4924);
or UO_393 (O_393,N_4970,N_4933);
and UO_394 (O_394,N_4999,N_4937);
or UO_395 (O_395,N_4937,N_4912);
or UO_396 (O_396,N_4958,N_4996);
or UO_397 (O_397,N_4955,N_4997);
or UO_398 (O_398,N_4920,N_4990);
xor UO_399 (O_399,N_4930,N_4904);
nand UO_400 (O_400,N_4950,N_4916);
nand UO_401 (O_401,N_4957,N_4995);
and UO_402 (O_402,N_4949,N_4944);
nor UO_403 (O_403,N_4960,N_4962);
nand UO_404 (O_404,N_4954,N_4922);
or UO_405 (O_405,N_4959,N_4961);
xnor UO_406 (O_406,N_4979,N_4968);
nand UO_407 (O_407,N_4939,N_4991);
nor UO_408 (O_408,N_4948,N_4952);
and UO_409 (O_409,N_4996,N_4920);
xor UO_410 (O_410,N_4904,N_4985);
xnor UO_411 (O_411,N_4999,N_4970);
nand UO_412 (O_412,N_4904,N_4965);
xnor UO_413 (O_413,N_4966,N_4926);
or UO_414 (O_414,N_4944,N_4988);
nand UO_415 (O_415,N_4953,N_4930);
and UO_416 (O_416,N_4985,N_4968);
nand UO_417 (O_417,N_4906,N_4945);
nand UO_418 (O_418,N_4983,N_4978);
or UO_419 (O_419,N_4969,N_4943);
or UO_420 (O_420,N_4969,N_4924);
and UO_421 (O_421,N_4934,N_4967);
xor UO_422 (O_422,N_4957,N_4971);
and UO_423 (O_423,N_4921,N_4983);
or UO_424 (O_424,N_4931,N_4904);
and UO_425 (O_425,N_4969,N_4972);
xnor UO_426 (O_426,N_4994,N_4906);
or UO_427 (O_427,N_4946,N_4926);
nand UO_428 (O_428,N_4901,N_4959);
xnor UO_429 (O_429,N_4969,N_4970);
or UO_430 (O_430,N_4935,N_4983);
nand UO_431 (O_431,N_4918,N_4903);
nand UO_432 (O_432,N_4995,N_4912);
and UO_433 (O_433,N_4945,N_4953);
or UO_434 (O_434,N_4987,N_4953);
xnor UO_435 (O_435,N_4952,N_4938);
or UO_436 (O_436,N_4985,N_4909);
xor UO_437 (O_437,N_4950,N_4918);
xor UO_438 (O_438,N_4914,N_4991);
xor UO_439 (O_439,N_4963,N_4996);
or UO_440 (O_440,N_4992,N_4909);
or UO_441 (O_441,N_4935,N_4993);
and UO_442 (O_442,N_4976,N_4993);
xor UO_443 (O_443,N_4987,N_4951);
or UO_444 (O_444,N_4911,N_4947);
nor UO_445 (O_445,N_4958,N_4920);
nand UO_446 (O_446,N_4987,N_4963);
nor UO_447 (O_447,N_4909,N_4942);
or UO_448 (O_448,N_4962,N_4983);
or UO_449 (O_449,N_4945,N_4956);
xnor UO_450 (O_450,N_4992,N_4958);
xnor UO_451 (O_451,N_4931,N_4958);
nand UO_452 (O_452,N_4924,N_4964);
xor UO_453 (O_453,N_4956,N_4998);
and UO_454 (O_454,N_4981,N_4907);
or UO_455 (O_455,N_4969,N_4989);
nor UO_456 (O_456,N_4984,N_4998);
nand UO_457 (O_457,N_4930,N_4923);
or UO_458 (O_458,N_4983,N_4961);
nor UO_459 (O_459,N_4977,N_4922);
nor UO_460 (O_460,N_4901,N_4944);
nand UO_461 (O_461,N_4902,N_4922);
nor UO_462 (O_462,N_4910,N_4951);
nor UO_463 (O_463,N_4900,N_4957);
nand UO_464 (O_464,N_4953,N_4904);
nand UO_465 (O_465,N_4924,N_4988);
or UO_466 (O_466,N_4979,N_4944);
xor UO_467 (O_467,N_4975,N_4955);
xnor UO_468 (O_468,N_4929,N_4914);
or UO_469 (O_469,N_4901,N_4910);
or UO_470 (O_470,N_4911,N_4925);
nand UO_471 (O_471,N_4959,N_4922);
or UO_472 (O_472,N_4928,N_4965);
xnor UO_473 (O_473,N_4963,N_4992);
or UO_474 (O_474,N_4919,N_4925);
nand UO_475 (O_475,N_4955,N_4935);
nor UO_476 (O_476,N_4943,N_4995);
xor UO_477 (O_477,N_4940,N_4917);
nor UO_478 (O_478,N_4995,N_4913);
nand UO_479 (O_479,N_4969,N_4945);
or UO_480 (O_480,N_4920,N_4948);
nand UO_481 (O_481,N_4952,N_4967);
nor UO_482 (O_482,N_4967,N_4926);
xnor UO_483 (O_483,N_4965,N_4912);
or UO_484 (O_484,N_4947,N_4956);
or UO_485 (O_485,N_4938,N_4911);
xor UO_486 (O_486,N_4990,N_4934);
nor UO_487 (O_487,N_4993,N_4919);
xnor UO_488 (O_488,N_4972,N_4988);
or UO_489 (O_489,N_4975,N_4960);
xor UO_490 (O_490,N_4948,N_4974);
xor UO_491 (O_491,N_4932,N_4905);
nand UO_492 (O_492,N_4973,N_4934);
xor UO_493 (O_493,N_4927,N_4932);
or UO_494 (O_494,N_4996,N_4990);
and UO_495 (O_495,N_4998,N_4931);
xnor UO_496 (O_496,N_4952,N_4905);
or UO_497 (O_497,N_4961,N_4936);
or UO_498 (O_498,N_4945,N_4974);
or UO_499 (O_499,N_4929,N_4959);
or UO_500 (O_500,N_4923,N_4902);
xor UO_501 (O_501,N_4965,N_4999);
or UO_502 (O_502,N_4939,N_4929);
nand UO_503 (O_503,N_4937,N_4960);
nor UO_504 (O_504,N_4967,N_4994);
or UO_505 (O_505,N_4960,N_4930);
xor UO_506 (O_506,N_4936,N_4997);
and UO_507 (O_507,N_4908,N_4979);
nand UO_508 (O_508,N_4961,N_4952);
and UO_509 (O_509,N_4976,N_4947);
xnor UO_510 (O_510,N_4986,N_4934);
or UO_511 (O_511,N_4982,N_4975);
nor UO_512 (O_512,N_4999,N_4982);
nor UO_513 (O_513,N_4958,N_4960);
or UO_514 (O_514,N_4924,N_4956);
xnor UO_515 (O_515,N_4903,N_4941);
nand UO_516 (O_516,N_4976,N_4994);
xor UO_517 (O_517,N_4995,N_4945);
nand UO_518 (O_518,N_4937,N_4961);
xor UO_519 (O_519,N_4931,N_4955);
xor UO_520 (O_520,N_4925,N_4918);
nor UO_521 (O_521,N_4977,N_4946);
xor UO_522 (O_522,N_4947,N_4901);
xnor UO_523 (O_523,N_4972,N_4917);
xor UO_524 (O_524,N_4977,N_4970);
and UO_525 (O_525,N_4993,N_4992);
nor UO_526 (O_526,N_4947,N_4973);
nor UO_527 (O_527,N_4960,N_4914);
or UO_528 (O_528,N_4970,N_4925);
nand UO_529 (O_529,N_4976,N_4936);
or UO_530 (O_530,N_4952,N_4972);
and UO_531 (O_531,N_4900,N_4981);
nand UO_532 (O_532,N_4900,N_4934);
xnor UO_533 (O_533,N_4906,N_4909);
or UO_534 (O_534,N_4928,N_4938);
nand UO_535 (O_535,N_4953,N_4915);
and UO_536 (O_536,N_4931,N_4914);
nor UO_537 (O_537,N_4962,N_4993);
or UO_538 (O_538,N_4913,N_4945);
nor UO_539 (O_539,N_4987,N_4942);
xnor UO_540 (O_540,N_4969,N_4930);
and UO_541 (O_541,N_4994,N_4945);
or UO_542 (O_542,N_4933,N_4909);
nand UO_543 (O_543,N_4988,N_4968);
or UO_544 (O_544,N_4931,N_4971);
or UO_545 (O_545,N_4905,N_4929);
nor UO_546 (O_546,N_4915,N_4940);
and UO_547 (O_547,N_4968,N_4902);
xor UO_548 (O_548,N_4982,N_4974);
xor UO_549 (O_549,N_4914,N_4982);
and UO_550 (O_550,N_4921,N_4946);
and UO_551 (O_551,N_4989,N_4999);
nor UO_552 (O_552,N_4933,N_4943);
and UO_553 (O_553,N_4925,N_4971);
nor UO_554 (O_554,N_4908,N_4952);
nor UO_555 (O_555,N_4991,N_4918);
xnor UO_556 (O_556,N_4934,N_4916);
or UO_557 (O_557,N_4988,N_4981);
nand UO_558 (O_558,N_4979,N_4933);
and UO_559 (O_559,N_4994,N_4914);
or UO_560 (O_560,N_4926,N_4986);
or UO_561 (O_561,N_4944,N_4904);
or UO_562 (O_562,N_4989,N_4905);
or UO_563 (O_563,N_4941,N_4948);
nor UO_564 (O_564,N_4998,N_4967);
nand UO_565 (O_565,N_4934,N_4984);
nor UO_566 (O_566,N_4971,N_4974);
and UO_567 (O_567,N_4913,N_4986);
nor UO_568 (O_568,N_4988,N_4990);
nor UO_569 (O_569,N_4934,N_4924);
and UO_570 (O_570,N_4979,N_4940);
xnor UO_571 (O_571,N_4988,N_4987);
or UO_572 (O_572,N_4979,N_4939);
and UO_573 (O_573,N_4941,N_4930);
or UO_574 (O_574,N_4991,N_4920);
nor UO_575 (O_575,N_4997,N_4933);
nor UO_576 (O_576,N_4998,N_4932);
nand UO_577 (O_577,N_4990,N_4907);
and UO_578 (O_578,N_4922,N_4914);
nand UO_579 (O_579,N_4944,N_4971);
xnor UO_580 (O_580,N_4953,N_4982);
or UO_581 (O_581,N_4963,N_4961);
or UO_582 (O_582,N_4989,N_4953);
xor UO_583 (O_583,N_4923,N_4987);
nand UO_584 (O_584,N_4939,N_4918);
xnor UO_585 (O_585,N_4976,N_4967);
and UO_586 (O_586,N_4925,N_4977);
and UO_587 (O_587,N_4943,N_4991);
and UO_588 (O_588,N_4973,N_4936);
nand UO_589 (O_589,N_4935,N_4963);
nand UO_590 (O_590,N_4923,N_4993);
and UO_591 (O_591,N_4979,N_4934);
or UO_592 (O_592,N_4970,N_4998);
and UO_593 (O_593,N_4939,N_4915);
nand UO_594 (O_594,N_4956,N_4943);
nor UO_595 (O_595,N_4918,N_4955);
xnor UO_596 (O_596,N_4932,N_4921);
nand UO_597 (O_597,N_4963,N_4948);
or UO_598 (O_598,N_4904,N_4942);
or UO_599 (O_599,N_4995,N_4971);
xnor UO_600 (O_600,N_4968,N_4969);
nor UO_601 (O_601,N_4967,N_4944);
nor UO_602 (O_602,N_4923,N_4924);
and UO_603 (O_603,N_4901,N_4987);
and UO_604 (O_604,N_4920,N_4950);
or UO_605 (O_605,N_4951,N_4988);
or UO_606 (O_606,N_4982,N_4931);
and UO_607 (O_607,N_4961,N_4954);
or UO_608 (O_608,N_4957,N_4985);
and UO_609 (O_609,N_4938,N_4962);
and UO_610 (O_610,N_4971,N_4913);
xor UO_611 (O_611,N_4980,N_4989);
nand UO_612 (O_612,N_4981,N_4917);
nand UO_613 (O_613,N_4994,N_4995);
and UO_614 (O_614,N_4970,N_4980);
nor UO_615 (O_615,N_4905,N_4923);
nand UO_616 (O_616,N_4930,N_4915);
nor UO_617 (O_617,N_4943,N_4926);
xor UO_618 (O_618,N_4994,N_4933);
and UO_619 (O_619,N_4998,N_4952);
nand UO_620 (O_620,N_4965,N_4996);
nor UO_621 (O_621,N_4944,N_4940);
or UO_622 (O_622,N_4938,N_4948);
xor UO_623 (O_623,N_4952,N_4953);
nand UO_624 (O_624,N_4921,N_4965);
nand UO_625 (O_625,N_4916,N_4966);
and UO_626 (O_626,N_4907,N_4974);
nand UO_627 (O_627,N_4923,N_4937);
and UO_628 (O_628,N_4920,N_4983);
nor UO_629 (O_629,N_4981,N_4909);
nor UO_630 (O_630,N_4977,N_4900);
xor UO_631 (O_631,N_4920,N_4992);
and UO_632 (O_632,N_4944,N_4991);
nor UO_633 (O_633,N_4988,N_4907);
nand UO_634 (O_634,N_4931,N_4981);
and UO_635 (O_635,N_4999,N_4947);
and UO_636 (O_636,N_4936,N_4989);
or UO_637 (O_637,N_4980,N_4969);
xnor UO_638 (O_638,N_4942,N_4977);
nor UO_639 (O_639,N_4999,N_4987);
and UO_640 (O_640,N_4905,N_4938);
nand UO_641 (O_641,N_4961,N_4981);
and UO_642 (O_642,N_4932,N_4992);
xnor UO_643 (O_643,N_4915,N_4995);
and UO_644 (O_644,N_4988,N_4927);
nor UO_645 (O_645,N_4912,N_4919);
or UO_646 (O_646,N_4958,N_4995);
or UO_647 (O_647,N_4924,N_4961);
nand UO_648 (O_648,N_4957,N_4925);
nand UO_649 (O_649,N_4938,N_4976);
and UO_650 (O_650,N_4904,N_4988);
nand UO_651 (O_651,N_4944,N_4909);
or UO_652 (O_652,N_4911,N_4975);
xnor UO_653 (O_653,N_4903,N_4948);
or UO_654 (O_654,N_4958,N_4907);
or UO_655 (O_655,N_4973,N_4901);
and UO_656 (O_656,N_4974,N_4965);
xnor UO_657 (O_657,N_4923,N_4964);
xnor UO_658 (O_658,N_4979,N_4946);
or UO_659 (O_659,N_4937,N_4919);
nand UO_660 (O_660,N_4947,N_4996);
or UO_661 (O_661,N_4930,N_4958);
and UO_662 (O_662,N_4916,N_4920);
nand UO_663 (O_663,N_4960,N_4980);
nand UO_664 (O_664,N_4918,N_4915);
or UO_665 (O_665,N_4951,N_4964);
and UO_666 (O_666,N_4941,N_4962);
xor UO_667 (O_667,N_4979,N_4911);
and UO_668 (O_668,N_4900,N_4912);
nand UO_669 (O_669,N_4904,N_4958);
nand UO_670 (O_670,N_4943,N_4966);
nand UO_671 (O_671,N_4968,N_4911);
or UO_672 (O_672,N_4971,N_4901);
nor UO_673 (O_673,N_4992,N_4935);
or UO_674 (O_674,N_4980,N_4946);
xnor UO_675 (O_675,N_4927,N_4961);
nor UO_676 (O_676,N_4925,N_4988);
or UO_677 (O_677,N_4976,N_4983);
nand UO_678 (O_678,N_4962,N_4919);
xnor UO_679 (O_679,N_4950,N_4915);
and UO_680 (O_680,N_4916,N_4917);
xor UO_681 (O_681,N_4911,N_4919);
nor UO_682 (O_682,N_4950,N_4952);
or UO_683 (O_683,N_4984,N_4918);
nor UO_684 (O_684,N_4911,N_4960);
or UO_685 (O_685,N_4919,N_4934);
nor UO_686 (O_686,N_4982,N_4917);
xor UO_687 (O_687,N_4949,N_4977);
xnor UO_688 (O_688,N_4933,N_4959);
nand UO_689 (O_689,N_4982,N_4910);
or UO_690 (O_690,N_4951,N_4998);
nor UO_691 (O_691,N_4982,N_4964);
nand UO_692 (O_692,N_4973,N_4959);
nand UO_693 (O_693,N_4950,N_4960);
nand UO_694 (O_694,N_4994,N_4998);
and UO_695 (O_695,N_4950,N_4984);
xor UO_696 (O_696,N_4976,N_4926);
nand UO_697 (O_697,N_4923,N_4978);
xor UO_698 (O_698,N_4971,N_4955);
or UO_699 (O_699,N_4945,N_4992);
nand UO_700 (O_700,N_4973,N_4999);
or UO_701 (O_701,N_4927,N_4951);
or UO_702 (O_702,N_4968,N_4974);
nand UO_703 (O_703,N_4928,N_4929);
nor UO_704 (O_704,N_4935,N_4900);
or UO_705 (O_705,N_4925,N_4976);
and UO_706 (O_706,N_4911,N_4990);
nor UO_707 (O_707,N_4918,N_4967);
and UO_708 (O_708,N_4952,N_4994);
nand UO_709 (O_709,N_4969,N_4997);
nor UO_710 (O_710,N_4987,N_4914);
or UO_711 (O_711,N_4972,N_4971);
or UO_712 (O_712,N_4925,N_4953);
nor UO_713 (O_713,N_4982,N_4941);
nand UO_714 (O_714,N_4980,N_4985);
and UO_715 (O_715,N_4987,N_4934);
nor UO_716 (O_716,N_4972,N_4979);
xnor UO_717 (O_717,N_4944,N_4973);
nand UO_718 (O_718,N_4917,N_4947);
nor UO_719 (O_719,N_4982,N_4998);
nor UO_720 (O_720,N_4937,N_4995);
and UO_721 (O_721,N_4988,N_4942);
xnor UO_722 (O_722,N_4980,N_4910);
and UO_723 (O_723,N_4952,N_4986);
nand UO_724 (O_724,N_4917,N_4915);
nand UO_725 (O_725,N_4996,N_4976);
nor UO_726 (O_726,N_4941,N_4928);
and UO_727 (O_727,N_4963,N_4926);
and UO_728 (O_728,N_4952,N_4951);
and UO_729 (O_729,N_4910,N_4967);
xor UO_730 (O_730,N_4972,N_4922);
nand UO_731 (O_731,N_4979,N_4988);
and UO_732 (O_732,N_4991,N_4999);
or UO_733 (O_733,N_4973,N_4996);
nor UO_734 (O_734,N_4998,N_4933);
nand UO_735 (O_735,N_4906,N_4991);
and UO_736 (O_736,N_4914,N_4901);
or UO_737 (O_737,N_4987,N_4950);
xnor UO_738 (O_738,N_4935,N_4944);
nor UO_739 (O_739,N_4954,N_4939);
nand UO_740 (O_740,N_4930,N_4999);
xnor UO_741 (O_741,N_4961,N_4916);
and UO_742 (O_742,N_4965,N_4957);
nand UO_743 (O_743,N_4959,N_4904);
and UO_744 (O_744,N_4900,N_4928);
nand UO_745 (O_745,N_4954,N_4990);
nor UO_746 (O_746,N_4946,N_4971);
xor UO_747 (O_747,N_4986,N_4997);
and UO_748 (O_748,N_4962,N_4969);
and UO_749 (O_749,N_4959,N_4911);
xnor UO_750 (O_750,N_4956,N_4978);
nand UO_751 (O_751,N_4946,N_4938);
nor UO_752 (O_752,N_4964,N_4955);
nand UO_753 (O_753,N_4907,N_4984);
nor UO_754 (O_754,N_4994,N_4972);
nand UO_755 (O_755,N_4907,N_4913);
nor UO_756 (O_756,N_4989,N_4933);
or UO_757 (O_757,N_4990,N_4924);
and UO_758 (O_758,N_4972,N_4902);
nor UO_759 (O_759,N_4966,N_4988);
xor UO_760 (O_760,N_4994,N_4979);
nand UO_761 (O_761,N_4913,N_4957);
nor UO_762 (O_762,N_4981,N_4927);
or UO_763 (O_763,N_4980,N_4954);
and UO_764 (O_764,N_4963,N_4934);
or UO_765 (O_765,N_4905,N_4975);
or UO_766 (O_766,N_4932,N_4967);
or UO_767 (O_767,N_4990,N_4969);
nor UO_768 (O_768,N_4900,N_4914);
xor UO_769 (O_769,N_4930,N_4902);
nor UO_770 (O_770,N_4917,N_4934);
nor UO_771 (O_771,N_4974,N_4966);
xor UO_772 (O_772,N_4957,N_4938);
and UO_773 (O_773,N_4917,N_4924);
or UO_774 (O_774,N_4940,N_4908);
nand UO_775 (O_775,N_4990,N_4930);
and UO_776 (O_776,N_4907,N_4923);
xor UO_777 (O_777,N_4926,N_4948);
and UO_778 (O_778,N_4915,N_4944);
or UO_779 (O_779,N_4953,N_4967);
nand UO_780 (O_780,N_4913,N_4981);
nand UO_781 (O_781,N_4919,N_4901);
xor UO_782 (O_782,N_4934,N_4936);
and UO_783 (O_783,N_4932,N_4914);
nor UO_784 (O_784,N_4992,N_4940);
nand UO_785 (O_785,N_4927,N_4993);
nor UO_786 (O_786,N_4932,N_4926);
or UO_787 (O_787,N_4964,N_4962);
and UO_788 (O_788,N_4907,N_4931);
or UO_789 (O_789,N_4936,N_4903);
nor UO_790 (O_790,N_4966,N_4969);
and UO_791 (O_791,N_4962,N_4942);
or UO_792 (O_792,N_4950,N_4945);
nand UO_793 (O_793,N_4995,N_4991);
and UO_794 (O_794,N_4964,N_4968);
nand UO_795 (O_795,N_4929,N_4962);
nand UO_796 (O_796,N_4965,N_4916);
or UO_797 (O_797,N_4986,N_4981);
and UO_798 (O_798,N_4948,N_4995);
or UO_799 (O_799,N_4974,N_4925);
and UO_800 (O_800,N_4970,N_4919);
nor UO_801 (O_801,N_4995,N_4964);
xnor UO_802 (O_802,N_4937,N_4969);
xnor UO_803 (O_803,N_4959,N_4980);
xnor UO_804 (O_804,N_4906,N_4934);
xnor UO_805 (O_805,N_4995,N_4951);
nor UO_806 (O_806,N_4929,N_4927);
or UO_807 (O_807,N_4935,N_4990);
nand UO_808 (O_808,N_4985,N_4913);
or UO_809 (O_809,N_4924,N_4933);
nor UO_810 (O_810,N_4937,N_4917);
or UO_811 (O_811,N_4932,N_4930);
and UO_812 (O_812,N_4987,N_4909);
or UO_813 (O_813,N_4907,N_4999);
nand UO_814 (O_814,N_4945,N_4976);
xor UO_815 (O_815,N_4930,N_4977);
and UO_816 (O_816,N_4905,N_4993);
or UO_817 (O_817,N_4943,N_4931);
or UO_818 (O_818,N_4943,N_4958);
xnor UO_819 (O_819,N_4921,N_4967);
and UO_820 (O_820,N_4987,N_4962);
xor UO_821 (O_821,N_4978,N_4951);
and UO_822 (O_822,N_4937,N_4914);
or UO_823 (O_823,N_4970,N_4963);
nand UO_824 (O_824,N_4999,N_4923);
or UO_825 (O_825,N_4934,N_4932);
xor UO_826 (O_826,N_4940,N_4925);
xnor UO_827 (O_827,N_4991,N_4941);
nand UO_828 (O_828,N_4963,N_4947);
nor UO_829 (O_829,N_4981,N_4980);
and UO_830 (O_830,N_4952,N_4993);
nand UO_831 (O_831,N_4904,N_4925);
or UO_832 (O_832,N_4966,N_4903);
or UO_833 (O_833,N_4994,N_4980);
nor UO_834 (O_834,N_4964,N_4945);
nand UO_835 (O_835,N_4912,N_4962);
nand UO_836 (O_836,N_4913,N_4914);
nor UO_837 (O_837,N_4992,N_4984);
xor UO_838 (O_838,N_4953,N_4909);
xor UO_839 (O_839,N_4926,N_4923);
xnor UO_840 (O_840,N_4978,N_4929);
or UO_841 (O_841,N_4959,N_4947);
nand UO_842 (O_842,N_4942,N_4986);
nor UO_843 (O_843,N_4972,N_4956);
and UO_844 (O_844,N_4998,N_4900);
nor UO_845 (O_845,N_4919,N_4990);
and UO_846 (O_846,N_4974,N_4987);
or UO_847 (O_847,N_4941,N_4939);
and UO_848 (O_848,N_4923,N_4967);
nor UO_849 (O_849,N_4995,N_4986);
nor UO_850 (O_850,N_4954,N_4941);
nor UO_851 (O_851,N_4972,N_4949);
nand UO_852 (O_852,N_4977,N_4933);
or UO_853 (O_853,N_4912,N_4923);
or UO_854 (O_854,N_4977,N_4947);
or UO_855 (O_855,N_4978,N_4901);
xnor UO_856 (O_856,N_4986,N_4906);
or UO_857 (O_857,N_4964,N_4921);
nor UO_858 (O_858,N_4922,N_4909);
nand UO_859 (O_859,N_4950,N_4959);
and UO_860 (O_860,N_4932,N_4990);
xnor UO_861 (O_861,N_4985,N_4900);
and UO_862 (O_862,N_4948,N_4988);
nor UO_863 (O_863,N_4956,N_4981);
nor UO_864 (O_864,N_4935,N_4941);
xnor UO_865 (O_865,N_4936,N_4978);
xnor UO_866 (O_866,N_4940,N_4964);
and UO_867 (O_867,N_4916,N_4901);
xor UO_868 (O_868,N_4934,N_4958);
and UO_869 (O_869,N_4926,N_4992);
or UO_870 (O_870,N_4954,N_4997);
nor UO_871 (O_871,N_4903,N_4906);
nor UO_872 (O_872,N_4920,N_4922);
xor UO_873 (O_873,N_4966,N_4907);
or UO_874 (O_874,N_4939,N_4977);
nor UO_875 (O_875,N_4972,N_4983);
or UO_876 (O_876,N_4968,N_4955);
and UO_877 (O_877,N_4962,N_4914);
or UO_878 (O_878,N_4976,N_4920);
xnor UO_879 (O_879,N_4943,N_4928);
xnor UO_880 (O_880,N_4966,N_4952);
or UO_881 (O_881,N_4956,N_4917);
nand UO_882 (O_882,N_4964,N_4996);
xnor UO_883 (O_883,N_4989,N_4913);
nand UO_884 (O_884,N_4969,N_4953);
nor UO_885 (O_885,N_4912,N_4959);
xor UO_886 (O_886,N_4941,N_4974);
nor UO_887 (O_887,N_4928,N_4986);
xor UO_888 (O_888,N_4917,N_4959);
and UO_889 (O_889,N_4953,N_4905);
nand UO_890 (O_890,N_4992,N_4943);
nand UO_891 (O_891,N_4974,N_4915);
nand UO_892 (O_892,N_4975,N_4926);
nand UO_893 (O_893,N_4999,N_4938);
or UO_894 (O_894,N_4963,N_4921);
nand UO_895 (O_895,N_4957,N_4990);
or UO_896 (O_896,N_4916,N_4984);
nand UO_897 (O_897,N_4939,N_4984);
nand UO_898 (O_898,N_4966,N_4985);
nor UO_899 (O_899,N_4970,N_4948);
or UO_900 (O_900,N_4946,N_4966);
or UO_901 (O_901,N_4939,N_4960);
nand UO_902 (O_902,N_4978,N_4944);
or UO_903 (O_903,N_4977,N_4957);
nor UO_904 (O_904,N_4911,N_4909);
nor UO_905 (O_905,N_4961,N_4904);
or UO_906 (O_906,N_4908,N_4938);
nor UO_907 (O_907,N_4954,N_4951);
nand UO_908 (O_908,N_4919,N_4921);
and UO_909 (O_909,N_4998,N_4977);
nor UO_910 (O_910,N_4971,N_4964);
nor UO_911 (O_911,N_4931,N_4996);
nor UO_912 (O_912,N_4981,N_4947);
nor UO_913 (O_913,N_4919,N_4931);
xor UO_914 (O_914,N_4928,N_4922);
or UO_915 (O_915,N_4960,N_4953);
xor UO_916 (O_916,N_4958,N_4971);
nor UO_917 (O_917,N_4919,N_4952);
and UO_918 (O_918,N_4918,N_4975);
and UO_919 (O_919,N_4929,N_4986);
xnor UO_920 (O_920,N_4949,N_4930);
xnor UO_921 (O_921,N_4986,N_4909);
xnor UO_922 (O_922,N_4990,N_4994);
xnor UO_923 (O_923,N_4931,N_4901);
xor UO_924 (O_924,N_4984,N_4952);
nand UO_925 (O_925,N_4954,N_4970);
xnor UO_926 (O_926,N_4928,N_4978);
and UO_927 (O_927,N_4942,N_4943);
or UO_928 (O_928,N_4935,N_4975);
nand UO_929 (O_929,N_4980,N_4920);
xor UO_930 (O_930,N_4915,N_4969);
nor UO_931 (O_931,N_4983,N_4960);
or UO_932 (O_932,N_4966,N_4962);
nor UO_933 (O_933,N_4949,N_4985);
nor UO_934 (O_934,N_4985,N_4914);
nor UO_935 (O_935,N_4948,N_4944);
and UO_936 (O_936,N_4904,N_4973);
and UO_937 (O_937,N_4978,N_4967);
or UO_938 (O_938,N_4979,N_4930);
nand UO_939 (O_939,N_4971,N_4956);
xnor UO_940 (O_940,N_4949,N_4912);
nand UO_941 (O_941,N_4906,N_4900);
nand UO_942 (O_942,N_4993,N_4912);
or UO_943 (O_943,N_4942,N_4933);
nand UO_944 (O_944,N_4933,N_4991);
nor UO_945 (O_945,N_4957,N_4941);
nor UO_946 (O_946,N_4910,N_4966);
nor UO_947 (O_947,N_4902,N_4957);
nand UO_948 (O_948,N_4928,N_4901);
or UO_949 (O_949,N_4902,N_4989);
or UO_950 (O_950,N_4937,N_4947);
xnor UO_951 (O_951,N_4919,N_4965);
or UO_952 (O_952,N_4919,N_4955);
xor UO_953 (O_953,N_4932,N_4953);
nand UO_954 (O_954,N_4928,N_4936);
and UO_955 (O_955,N_4928,N_4948);
or UO_956 (O_956,N_4905,N_4955);
nand UO_957 (O_957,N_4982,N_4916);
nor UO_958 (O_958,N_4983,N_4936);
nand UO_959 (O_959,N_4949,N_4970);
nor UO_960 (O_960,N_4903,N_4984);
or UO_961 (O_961,N_4907,N_4949);
xor UO_962 (O_962,N_4962,N_4911);
and UO_963 (O_963,N_4927,N_4944);
nor UO_964 (O_964,N_4940,N_4912);
and UO_965 (O_965,N_4900,N_4922);
or UO_966 (O_966,N_4900,N_4982);
xor UO_967 (O_967,N_4962,N_4959);
xnor UO_968 (O_968,N_4980,N_4904);
xor UO_969 (O_969,N_4940,N_4932);
and UO_970 (O_970,N_4995,N_4911);
nor UO_971 (O_971,N_4950,N_4996);
and UO_972 (O_972,N_4940,N_4959);
nand UO_973 (O_973,N_4969,N_4908);
and UO_974 (O_974,N_4975,N_4962);
nand UO_975 (O_975,N_4960,N_4908);
nand UO_976 (O_976,N_4916,N_4910);
nand UO_977 (O_977,N_4928,N_4924);
nor UO_978 (O_978,N_4984,N_4970);
or UO_979 (O_979,N_4974,N_4910);
nand UO_980 (O_980,N_4941,N_4996);
or UO_981 (O_981,N_4901,N_4942);
or UO_982 (O_982,N_4996,N_4960);
or UO_983 (O_983,N_4965,N_4935);
nand UO_984 (O_984,N_4946,N_4927);
and UO_985 (O_985,N_4995,N_4921);
and UO_986 (O_986,N_4914,N_4974);
or UO_987 (O_987,N_4941,N_4961);
and UO_988 (O_988,N_4907,N_4937);
or UO_989 (O_989,N_4952,N_4999);
and UO_990 (O_990,N_4900,N_4923);
nor UO_991 (O_991,N_4990,N_4927);
or UO_992 (O_992,N_4909,N_4917);
nor UO_993 (O_993,N_4901,N_4977);
xor UO_994 (O_994,N_4905,N_4976);
xor UO_995 (O_995,N_4978,N_4985);
nand UO_996 (O_996,N_4924,N_4947);
and UO_997 (O_997,N_4996,N_4998);
or UO_998 (O_998,N_4992,N_4967);
xnor UO_999 (O_999,N_4931,N_4997);
endmodule