module basic_2000_20000_2500_4_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1793,In_743);
or U1 (N_1,In_1234,In_1761);
or U2 (N_2,In_1445,In_466);
or U3 (N_3,In_11,In_853);
nand U4 (N_4,In_154,In_696);
or U5 (N_5,In_1739,In_960);
nand U6 (N_6,In_704,In_1668);
or U7 (N_7,In_1901,In_160);
nand U8 (N_8,In_1695,In_1674);
or U9 (N_9,In_1794,In_1880);
and U10 (N_10,In_1660,In_1856);
nor U11 (N_11,In_360,In_1920);
nor U12 (N_12,In_1106,In_1904);
nor U13 (N_13,In_1449,In_818);
and U14 (N_14,In_1529,In_580);
nor U15 (N_15,In_468,In_321);
or U16 (N_16,In_238,In_1231);
nand U17 (N_17,In_234,In_66);
and U18 (N_18,In_871,In_1972);
nand U19 (N_19,In_1614,In_1775);
nand U20 (N_20,In_210,In_431);
and U21 (N_21,In_576,In_366);
nor U22 (N_22,In_1437,In_139);
nand U23 (N_23,In_10,In_215);
nor U24 (N_24,In_1531,In_994);
and U25 (N_25,In_1135,In_1889);
and U26 (N_26,In_569,In_1276);
or U27 (N_27,In_1405,In_485);
nor U28 (N_28,In_379,In_1894);
and U29 (N_29,In_971,In_1390);
or U30 (N_30,In_371,In_1457);
and U31 (N_31,In_243,In_1357);
or U32 (N_32,In_456,In_342);
nand U33 (N_33,In_1962,In_136);
nor U34 (N_34,In_896,In_1267);
or U35 (N_35,In_983,In_59);
xnor U36 (N_36,In_1283,In_931);
nand U37 (N_37,In_1485,In_1341);
nor U38 (N_38,In_959,In_1333);
xor U39 (N_39,In_623,In_605);
nand U40 (N_40,In_1151,In_51);
or U41 (N_41,In_1062,In_1646);
nor U42 (N_42,In_1912,In_1483);
nand U43 (N_43,In_1490,In_1410);
or U44 (N_44,In_308,In_462);
nor U45 (N_45,In_1535,In_1050);
and U46 (N_46,In_748,In_7);
and U47 (N_47,In_268,In_1762);
or U48 (N_48,In_1564,In_716);
nor U49 (N_49,In_1905,In_1902);
or U50 (N_50,In_740,In_547);
and U51 (N_51,In_1145,In_311);
nor U52 (N_52,In_1781,In_251);
or U53 (N_53,In_247,In_588);
nor U54 (N_54,In_546,In_669);
nor U55 (N_55,In_1201,In_200);
nor U56 (N_56,In_1651,In_1324);
or U57 (N_57,In_843,In_369);
and U58 (N_58,In_1935,In_339);
nor U59 (N_59,In_447,In_214);
or U60 (N_60,In_1286,In_524);
or U61 (N_61,In_276,In_1077);
and U62 (N_62,In_1492,In_285);
and U63 (N_63,In_1611,In_1577);
nand U64 (N_64,In_1427,In_1165);
or U65 (N_65,In_831,In_1828);
or U66 (N_66,In_883,In_387);
nor U67 (N_67,In_1021,In_1732);
or U68 (N_68,In_1868,In_1735);
or U69 (N_69,In_1583,In_1008);
nor U70 (N_70,In_176,In_1501);
nand U71 (N_71,In_675,In_162);
nor U72 (N_72,In_718,In_350);
and U73 (N_73,In_956,In_315);
nand U74 (N_74,In_938,In_543);
nand U75 (N_75,In_1710,In_1945);
and U76 (N_76,In_309,In_497);
and U77 (N_77,In_312,In_1970);
or U78 (N_78,In_1161,In_1840);
and U79 (N_79,In_1619,In_1111);
or U80 (N_80,In_663,In_1884);
nand U81 (N_81,In_1585,In_1228);
nor U82 (N_82,In_691,In_758);
nand U83 (N_83,In_1398,In_594);
and U84 (N_84,In_448,In_1486);
nor U85 (N_85,In_1040,In_728);
nor U86 (N_86,In_1192,In_152);
nor U87 (N_87,In_884,In_1745);
nand U88 (N_88,In_392,In_1310);
and U89 (N_89,In_271,In_1957);
nor U90 (N_90,In_377,In_211);
nand U91 (N_91,In_1003,In_231);
nand U92 (N_92,In_157,In_689);
nand U93 (N_93,In_1353,In_954);
nand U94 (N_94,In_600,In_63);
or U95 (N_95,In_1691,In_49);
or U96 (N_96,In_1302,In_1463);
and U97 (N_97,In_964,In_292);
and U98 (N_98,In_278,In_1934);
nand U99 (N_99,In_1584,In_1843);
nor U100 (N_100,In_1787,In_1963);
nor U101 (N_101,In_750,In_1751);
nor U102 (N_102,In_341,In_1654);
nor U103 (N_103,In_1223,In_979);
nor U104 (N_104,In_374,In_1561);
nand U105 (N_105,In_1769,In_1924);
or U106 (N_106,In_627,In_1573);
nand U107 (N_107,In_1400,In_1084);
and U108 (N_108,In_1742,In_1725);
or U109 (N_109,In_1811,In_472);
nor U110 (N_110,In_1058,In_1607);
nand U111 (N_111,In_610,In_898);
nor U112 (N_112,In_1768,In_1314);
or U113 (N_113,In_572,In_1472);
or U114 (N_114,In_50,In_1612);
nand U115 (N_115,In_1892,In_1630);
nand U116 (N_116,In_1361,In_1337);
or U117 (N_117,In_1988,In_901);
nand U118 (N_118,In_1103,In_779);
or U119 (N_119,In_1647,In_1622);
or U120 (N_120,In_146,In_87);
or U121 (N_121,In_1331,In_1676);
and U122 (N_122,In_1504,In_286);
nor U123 (N_123,In_719,In_1296);
or U124 (N_124,In_1100,In_1915);
and U125 (N_125,In_1493,In_422);
or U126 (N_126,In_1347,In_1886);
nor U127 (N_127,In_895,In_1566);
and U128 (N_128,In_595,In_209);
and U129 (N_129,In_27,In_56);
nand U130 (N_130,In_226,In_1125);
nand U131 (N_131,In_1608,In_1044);
nor U132 (N_132,In_780,In_17);
nand U133 (N_133,In_403,In_1562);
nand U134 (N_134,In_294,In_1956);
or U135 (N_135,In_1034,In_1866);
nor U136 (N_136,In_1325,In_782);
nor U137 (N_137,In_1232,In_1443);
nand U138 (N_138,In_464,In_1329);
nor U139 (N_139,In_1266,In_463);
nor U140 (N_140,In_582,In_1086);
and U141 (N_141,In_842,In_941);
or U142 (N_142,In_1613,In_1638);
and U143 (N_143,In_969,In_1042);
and U144 (N_144,In_1248,In_654);
and U145 (N_145,In_736,In_705);
nor U146 (N_146,In_1699,In_90);
or U147 (N_147,In_1805,In_57);
nand U148 (N_148,In_764,In_245);
and U149 (N_149,In_331,In_180);
or U150 (N_150,In_746,In_1785);
xor U151 (N_151,In_833,In_5);
nand U152 (N_152,In_1830,In_1670);
or U153 (N_153,In_1079,In_679);
nor U154 (N_154,In_1547,In_1243);
nor U155 (N_155,In_281,In_1984);
and U156 (N_156,In_423,In_855);
nand U157 (N_157,In_989,In_601);
and U158 (N_158,In_1168,In_436);
and U159 (N_159,In_1429,In_1865);
nand U160 (N_160,In_1206,In_510);
nor U161 (N_161,In_1051,In_1662);
nand U162 (N_162,In_351,In_427);
or U163 (N_163,In_1899,In_401);
and U164 (N_164,In_1096,In_535);
and U165 (N_165,In_1539,In_1969);
and U166 (N_166,In_310,In_1839);
and U167 (N_167,In_95,In_202);
or U168 (N_168,In_1820,In_688);
and U169 (N_169,In_438,In_1250);
or U170 (N_170,In_1261,In_1610);
or U171 (N_171,In_1778,In_89);
or U172 (N_172,In_1747,In_1910);
and U173 (N_173,In_1394,In_265);
nand U174 (N_174,In_972,In_1404);
or U175 (N_175,In_163,In_106);
nor U176 (N_176,In_693,In_241);
or U177 (N_177,In_1278,In_1530);
nor U178 (N_178,In_900,In_246);
nor U179 (N_179,In_1795,In_706);
nand U180 (N_180,In_625,In_1727);
nand U181 (N_181,In_391,In_655);
nor U182 (N_182,In_71,In_1533);
nand U183 (N_183,In_1028,In_1881);
or U184 (N_184,In_807,In_1254);
or U185 (N_185,In_1665,In_213);
nor U186 (N_186,In_613,In_1133);
nand U187 (N_187,In_1696,In_1351);
or U188 (N_188,In_1025,In_41);
and U189 (N_189,In_1435,In_1401);
xor U190 (N_190,In_1444,In_1757);
nand U191 (N_191,In_336,In_1537);
or U192 (N_192,In_975,In_881);
and U193 (N_193,In_757,In_1797);
xnor U194 (N_194,In_399,In_1164);
and U195 (N_195,In_1152,In_306);
or U196 (N_196,In_1053,In_658);
nand U197 (N_197,In_97,In_1167);
and U198 (N_198,In_1627,In_1759);
and U199 (N_199,In_778,In_1569);
nand U200 (N_200,In_222,In_483);
and U201 (N_201,In_1246,In_493);
nor U202 (N_202,In_1122,In_1678);
nor U203 (N_203,In_1703,In_1076);
nand U204 (N_204,In_1551,In_861);
and U205 (N_205,In_927,In_1687);
or U206 (N_206,In_815,In_1527);
nor U207 (N_207,In_1697,In_1540);
or U208 (N_208,In_1194,In_1536);
nor U209 (N_209,In_496,In_1626);
and U210 (N_210,In_457,In_854);
or U211 (N_211,In_888,In_1059);
and U212 (N_212,In_859,In_648);
nor U213 (N_213,In_824,In_917);
nand U214 (N_214,In_1624,In_729);
nor U215 (N_215,In_1354,In_1301);
nor U216 (N_216,In_1581,In_1116);
nor U217 (N_217,In_1766,In_1862);
nand U218 (N_218,In_0,In_1603);
or U219 (N_219,In_1321,In_257);
xor U220 (N_220,In_1211,In_799);
or U221 (N_221,In_943,In_1016);
nand U222 (N_222,In_334,In_187);
or U223 (N_223,In_287,In_77);
or U224 (N_224,In_1235,In_512);
xor U225 (N_225,In_277,In_1744);
and U226 (N_226,In_414,In_987);
or U227 (N_227,In_849,In_1604);
or U228 (N_228,In_358,In_1383);
xor U229 (N_229,In_792,In_1731);
nand U230 (N_230,In_1502,In_385);
nand U231 (N_231,In_587,In_1944);
and U232 (N_232,In_1989,In_318);
and U233 (N_233,In_1519,In_1015);
nand U234 (N_234,In_284,In_958);
nand U235 (N_235,In_1796,In_1618);
nand U236 (N_236,In_1487,In_1085);
nor U237 (N_237,In_1222,In_1525);
and U238 (N_238,In_1875,In_936);
nand U239 (N_239,In_1774,In_362);
and U240 (N_240,In_409,In_539);
and U241 (N_241,In_1149,In_1440);
nand U242 (N_242,In_788,In_380);
nor U243 (N_243,In_1682,In_1422);
nand U244 (N_244,In_225,In_1157);
or U245 (N_245,In_1356,In_745);
nor U246 (N_246,In_1066,In_194);
and U247 (N_247,In_1433,In_459);
nand U248 (N_248,In_1092,In_1397);
nor U249 (N_249,In_1163,In_279);
or U250 (N_250,In_1426,In_538);
nor U251 (N_251,In_617,In_394);
and U252 (N_252,In_96,In_1458);
and U253 (N_253,In_1236,In_1661);
nor U254 (N_254,In_1032,In_1000);
and U255 (N_255,In_872,In_1464);
nor U256 (N_256,In_258,In_1863);
nand U257 (N_257,In_1045,In_1590);
or U258 (N_258,In_1808,In_505);
xor U259 (N_259,In_869,In_862);
or U260 (N_260,In_957,In_1565);
or U261 (N_261,In_1755,In_174);
nand U262 (N_262,In_1366,In_1848);
and U263 (N_263,In_698,In_1360);
nor U264 (N_264,In_1280,In_791);
or U265 (N_265,In_806,In_184);
or U266 (N_266,In_674,In_1128);
or U267 (N_267,In_100,In_1995);
or U268 (N_268,In_1249,In_252);
nand U269 (N_269,In_1481,In_786);
nor U270 (N_270,In_1144,In_619);
nor U271 (N_271,In_1495,In_1409);
xnor U272 (N_272,In_981,In_1037);
or U273 (N_273,In_12,In_420);
or U274 (N_274,In_879,In_1009);
nand U275 (N_275,In_13,In_660);
nand U276 (N_276,In_783,In_1600);
nor U277 (N_277,In_935,In_1098);
nand U278 (N_278,In_1245,In_34);
and U279 (N_279,In_632,In_646);
and U280 (N_280,In_1749,In_1210);
nor U281 (N_281,In_487,In_1575);
or U282 (N_282,In_255,In_518);
nand U283 (N_283,In_1279,In_1802);
and U284 (N_284,In_529,In_240);
nand U285 (N_285,In_460,In_249);
or U286 (N_286,In_1017,In_1977);
nand U287 (N_287,In_189,In_320);
or U288 (N_288,In_274,In_416);
nand U289 (N_289,In_1338,In_474);
nand U290 (N_290,In_282,In_1099);
nand U291 (N_291,In_1473,In_978);
nor U292 (N_292,In_1883,In_145);
or U293 (N_293,In_1968,In_1849);
or U294 (N_294,In_302,In_891);
and U295 (N_295,In_451,In_1983);
nor U296 (N_296,In_1406,In_577);
nand U297 (N_297,In_852,In_79);
and U298 (N_298,In_1430,In_1171);
nand U299 (N_299,In_733,In_1132);
nor U300 (N_300,In_695,In_1669);
nand U301 (N_301,In_1358,In_1809);
and U302 (N_302,In_440,In_1393);
or U303 (N_303,In_525,In_657);
nand U304 (N_304,In_633,In_823);
nor U305 (N_305,In_98,In_1538);
and U306 (N_306,In_322,In_647);
nand U307 (N_307,In_620,In_795);
and U308 (N_308,In_94,In_768);
nand U309 (N_309,In_982,In_785);
nor U310 (N_310,In_937,In_349);
nor U311 (N_311,In_819,In_1065);
nor U312 (N_312,In_353,In_47);
nor U313 (N_313,In_597,In_1907);
or U314 (N_314,In_1684,In_640);
or U315 (N_315,In_1973,In_1764);
nand U316 (N_316,In_630,In_589);
nor U317 (N_317,In_1195,In_110);
nand U318 (N_318,In_494,In_363);
nor U319 (N_319,In_1292,In_770);
and U320 (N_320,In_612,In_450);
or U321 (N_321,In_1655,In_1216);
nor U322 (N_322,In_624,In_1847);
or U323 (N_323,In_178,In_105);
and U324 (N_324,In_313,In_712);
or U325 (N_325,In_473,In_356);
or U326 (N_326,In_502,In_682);
or U327 (N_327,In_760,In_874);
nor U328 (N_328,In_398,In_1318);
or U329 (N_329,In_571,In_1287);
nor U330 (N_330,In_1162,In_680);
and U331 (N_331,In_45,In_1418);
and U332 (N_332,In_92,In_1829);
or U333 (N_333,In_511,In_16);
or U334 (N_334,In_886,In_1233);
nor U335 (N_335,In_1158,In_307);
nor U336 (N_336,In_429,In_1688);
or U337 (N_337,In_1947,In_383);
xnor U338 (N_338,In_1859,In_314);
nor U339 (N_339,In_1861,In_372);
nor U340 (N_340,In_1306,In_75);
and U341 (N_341,In_1469,In_1312);
nand U342 (N_342,In_1258,In_1002);
or U343 (N_343,In_501,In_685);
nor U344 (N_344,In_1371,In_1870);
or U345 (N_345,In_1416,In_254);
nor U346 (N_346,In_386,In_607);
xor U347 (N_347,In_1960,In_573);
xor U348 (N_348,In_1589,In_708);
and U349 (N_349,In_428,In_498);
or U350 (N_350,In_944,In_1153);
xor U351 (N_351,In_354,In_986);
nand U352 (N_352,In_1677,In_1885);
or U353 (N_353,In_335,In_919);
nand U354 (N_354,In_122,In_229);
and U355 (N_355,In_1184,In_121);
or U356 (N_356,In_1139,In_889);
nand U357 (N_357,In_35,In_1352);
xnor U358 (N_358,In_78,In_1365);
nor U359 (N_359,In_1202,In_444);
nand U360 (N_360,In_915,In_1679);
and U361 (N_361,In_1552,In_128);
nor U362 (N_362,In_230,In_875);
nor U363 (N_363,In_1081,In_641);
and U364 (N_364,In_1514,In_33);
nor U365 (N_365,In_435,In_1215);
or U366 (N_366,In_83,In_730);
and U367 (N_367,In_649,In_1175);
nand U368 (N_368,In_482,In_1137);
and U369 (N_369,In_291,In_490);
or U370 (N_370,In_1556,In_904);
or U371 (N_371,In_1240,In_1064);
and U372 (N_372,In_1737,In_1568);
and U373 (N_373,In_1411,In_382);
nand U374 (N_374,In_1497,In_1498);
nand U375 (N_375,In_1403,In_24);
or U376 (N_376,In_1980,In_26);
nor U377 (N_377,In_1996,In_1091);
and U378 (N_378,In_856,In_1982);
or U379 (N_379,In_40,In_1997);
nor U380 (N_380,In_906,In_1523);
nor U381 (N_381,In_329,In_1185);
nand U382 (N_382,In_1822,In_1951);
or U383 (N_383,In_947,In_1779);
nand U384 (N_384,In_1369,In_754);
or U385 (N_385,In_1466,In_364);
or U386 (N_386,In_916,In_1524);
nor U387 (N_387,In_541,In_190);
nor U388 (N_388,In_23,In_727);
or U389 (N_389,In_1928,In_1958);
or U390 (N_390,In_81,In_1906);
xnor U391 (N_391,In_344,In_950);
xor U392 (N_392,In_530,In_581);
and U393 (N_393,In_1105,In_1543);
nand U394 (N_394,In_1644,In_134);
nand U395 (N_395,In_404,In_1705);
and U396 (N_396,In_533,In_651);
nand U397 (N_397,In_52,In_1078);
nor U398 (N_398,In_1917,In_1707);
and U399 (N_399,In_319,In_540);
or U400 (N_400,In_1818,In_1726);
and U401 (N_401,In_1389,In_191);
nand U402 (N_402,In_1606,In_1491);
and U403 (N_403,In_347,In_108);
nand U404 (N_404,In_1072,In_559);
xnor U405 (N_405,In_1113,In_1966);
and U406 (N_406,In_455,In_1290);
nor U407 (N_407,In_28,In_1685);
nor U408 (N_408,In_101,In_638);
nor U409 (N_409,In_1323,In_949);
nor U410 (N_410,In_301,In_1038);
and U411 (N_411,In_1663,In_439);
or U412 (N_412,In_1650,In_1635);
nor U413 (N_413,In_825,In_1515);
and U414 (N_414,In_1681,In_596);
or U415 (N_415,In_147,In_1967);
or U416 (N_416,In_183,In_953);
nor U417 (N_417,In_711,In_132);
nor U418 (N_418,In_542,In_1061);
or U419 (N_419,In_32,In_809);
and U420 (N_420,In_699,In_1919);
or U421 (N_421,In_1871,In_296);
nand U422 (N_422,In_1760,In_150);
nand U423 (N_423,In_1238,In_1455);
and U424 (N_424,In_980,In_1642);
and U425 (N_425,In_68,In_1272);
nor U426 (N_426,In_609,In_531);
xnor U427 (N_427,In_1505,In_1680);
or U428 (N_428,In_902,In_378);
nand U429 (N_429,In_549,In_774);
nand U430 (N_430,In_1929,In_1499);
or U431 (N_431,In_1414,In_1134);
nand U432 (N_432,In_870,In_1571);
and U433 (N_433,In_1986,In_844);
or U434 (N_434,In_393,In_1667);
nand U435 (N_435,In_188,In_634);
and U436 (N_436,In_198,In_621);
nor U437 (N_437,In_1579,In_1548);
nor U438 (N_438,In_266,In_553);
nor U439 (N_439,In_1054,In_1582);
nor U440 (N_440,In_725,In_673);
nor U441 (N_441,In_556,In_637);
nor U442 (N_442,In_626,In_317);
or U443 (N_443,In_1916,In_939);
nor U444 (N_444,In_1262,In_264);
and U445 (N_445,In_1392,In_261);
and U446 (N_446,In_141,In_650);
nand U447 (N_447,In_1056,In_1842);
and U448 (N_448,In_1253,In_1189);
nor U449 (N_449,In_1110,In_491);
or U450 (N_450,In_1023,In_1067);
nand U451 (N_451,In_1036,In_527);
nand U452 (N_452,In_1070,In_645);
and U453 (N_453,In_926,In_1297);
or U454 (N_454,In_263,In_1940);
or U455 (N_455,In_109,In_585);
and U456 (N_456,In_1219,In_810);
nand U457 (N_457,In_1448,In_3);
nand U458 (N_458,In_1992,In_1227);
nor U459 (N_459,In_678,In_453);
nor U460 (N_460,In_461,In_811);
and U461 (N_461,In_44,In_945);
and U462 (N_462,In_1309,In_1709);
or U463 (N_463,In_1355,In_1180);
or U464 (N_464,In_397,In_1399);
and U465 (N_465,In_1922,In_1855);
or U466 (N_466,In_913,In_873);
nor U467 (N_467,In_118,In_933);
or U468 (N_468,In_1746,In_1178);
nor U469 (N_469,In_1478,In_1819);
and U470 (N_470,In_446,In_812);
nor U471 (N_471,In_1335,In_1615);
and U472 (N_472,In_199,In_169);
nor U473 (N_473,In_484,In_218);
and U474 (N_474,In_102,In_677);
nor U475 (N_475,In_413,In_1415);
and U476 (N_476,In_1273,In_561);
and U477 (N_477,In_421,In_478);
and U478 (N_478,In_1801,In_390);
or U479 (N_479,In_910,In_1269);
nand U480 (N_480,In_887,In_1198);
nor U481 (N_481,In_14,In_1419);
nand U482 (N_482,In_1150,In_1837);
and U483 (N_483,In_709,In_1792);
or U484 (N_484,In_999,In_1348);
nor U485 (N_485,In_653,In_272);
nand U486 (N_486,In_290,In_985);
nand U487 (N_487,In_1126,In_1169);
nor U488 (N_488,In_1570,In_239);
nor U489 (N_489,In_348,In_137);
nor U490 (N_490,In_828,In_161);
nor U491 (N_491,In_1317,In_1623);
nor U492 (N_492,In_742,In_1937);
nor U493 (N_493,In_995,In_1720);
nand U494 (N_494,In_1197,In_988);
and U495 (N_495,In_1639,In_721);
nand U496 (N_496,In_692,In_1740);
nor U497 (N_497,In_123,In_1702);
and U498 (N_498,In_1823,In_1686);
xnor U499 (N_499,In_814,In_479);
nand U500 (N_500,In_1363,In_1462);
nand U501 (N_501,In_1832,In_796);
nor U502 (N_502,In_76,In_475);
or U503 (N_503,In_111,In_1456);
or U504 (N_504,In_326,In_175);
nor U505 (N_505,In_29,In_963);
nand U506 (N_506,In_838,In_6);
or U507 (N_507,In_1782,In_1256);
nand U508 (N_508,In_1713,In_1729);
or U509 (N_509,In_1207,In_1388);
and U510 (N_510,In_973,In_1593);
or U511 (N_511,In_250,In_1391);
nor U512 (N_512,In_602,In_976);
nand U513 (N_513,In_74,In_1131);
and U514 (N_514,In_1019,In_1874);
or U515 (N_515,In_1738,In_603);
nand U516 (N_516,In_1181,In_835);
nor U517 (N_517,In_1716,In_1182);
and U518 (N_518,In_1773,In_1666);
or U519 (N_519,In_1109,In_179);
nor U520 (N_520,In_1226,In_593);
or U521 (N_521,In_1438,In_1313);
or U522 (N_522,In_1700,In_690);
and U523 (N_523,In_1193,In_702);
nor U524 (N_524,In_445,In_402);
and U525 (N_525,In_155,In_1328);
nor U526 (N_526,In_993,In_1734);
nor U527 (N_527,In_1550,In_1208);
and U528 (N_528,In_65,In_412);
nand U529 (N_529,In_470,In_1748);
and U530 (N_530,In_452,In_1482);
xor U531 (N_531,In_1020,In_848);
nand U532 (N_532,In_1041,In_299);
nor U533 (N_533,In_1965,In_1252);
nor U534 (N_534,In_686,In_1123);
and U535 (N_535,In_672,In_1563);
or U536 (N_536,In_1631,In_506);
and U537 (N_537,In_477,In_1102);
nand U538 (N_538,In_1893,In_1368);
and U539 (N_539,In_1402,In_1701);
and U540 (N_540,In_1806,In_583);
and U541 (N_541,In_373,In_1717);
and U542 (N_542,In_295,In_1814);
nand U543 (N_543,In_256,In_878);
and U544 (N_544,In_1683,In_1765);
nand U545 (N_545,In_1294,In_850);
nand U546 (N_546,In_813,In_753);
nor U547 (N_547,In_1345,In_499);
nand U548 (N_548,In_262,In_1380);
or U549 (N_549,In_676,In_1359);
or U550 (N_550,In_1452,In_1932);
nor U551 (N_551,In_1148,In_797);
nor U552 (N_552,In_1247,In_1601);
and U553 (N_553,In_1909,In_1914);
nand U554 (N_554,In_1378,In_652);
or U555 (N_555,In_273,In_1867);
xnor U556 (N_556,In_1616,In_1200);
nor U557 (N_557,In_1580,In_1447);
nor U558 (N_558,In_604,In_558);
or U559 (N_559,In_1659,In_611);
nor U560 (N_560,In_1555,In_1022);
nand U561 (N_561,In_1509,In_375);
nor U562 (N_562,In_196,In_43);
and U563 (N_563,In_469,In_1719);
nor U564 (N_564,In_237,In_773);
or U565 (N_565,In_130,In_1954);
and U566 (N_566,In_1844,In_1942);
or U567 (N_567,In_370,In_1320);
nor U568 (N_568,In_771,In_2);
or U569 (N_569,In_922,In_1362);
or U570 (N_570,In_1653,In_9);
and U571 (N_571,In_885,In_575);
or U572 (N_572,In_1784,In_1459);
nand U573 (N_573,In_384,In_739);
nor U574 (N_574,In_1350,In_1974);
and U575 (N_575,In_167,In_907);
nand U576 (N_576,In_925,In_903);
nor U577 (N_577,In_233,In_1229);
and U578 (N_578,In_777,In_1291);
or U579 (N_579,In_1836,In_1251);
and U580 (N_580,In_528,In_1791);
nand U581 (N_581,In_735,In_599);
and U582 (N_582,In_1159,In_1255);
nand U583 (N_583,In_928,In_909);
or U584 (N_584,In_359,In_1948);
or U585 (N_585,In_967,In_877);
nand U586 (N_586,In_1263,In_509);
nand U587 (N_587,In_298,In_1625);
nand U588 (N_588,In_616,In_803);
nor U589 (N_589,In_1521,In_1218);
and U590 (N_590,In_156,In_267);
or U591 (N_591,In_1209,In_955);
nand U592 (N_592,In_1424,In_346);
nor U593 (N_593,In_1692,In_866);
nand U594 (N_594,In_1783,In_1981);
and U595 (N_595,In_1943,In_1069);
nor U596 (N_596,In_212,In_1999);
or U597 (N_597,In_1187,In_1926);
nor U598 (N_598,In_1408,In_72);
and U599 (N_599,In_1330,In_968);
xnor U600 (N_600,In_288,In_1741);
nand U601 (N_601,In_67,In_495);
and U602 (N_602,In_1274,In_236);
nor U603 (N_603,In_1074,In_952);
or U604 (N_604,In_42,In_1304);
and U605 (N_605,In_164,In_775);
and U606 (N_606,In_1572,In_1450);
or U607 (N_607,In_701,In_1576);
or U608 (N_608,In_343,In_1810);
or U609 (N_609,In_1196,In_260);
nor U610 (N_610,In_1264,In_381);
nand U611 (N_611,In_1628,In_827);
nor U612 (N_612,In_1441,In_1033);
nor U613 (N_613,In_1179,In_1068);
and U614 (N_614,In_1071,In_1117);
nor U615 (N_615,In_283,In_1374);
nor U616 (N_616,In_432,In_908);
or U617 (N_617,In_905,In_1018);
and U618 (N_618,In_1242,In_668);
and U619 (N_619,In_1637,In_186);
nand U620 (N_620,In_1082,In_1629);
nand U621 (N_621,In_1174,In_1528);
nor U622 (N_622,In_269,In_1477);
nand U623 (N_623,In_1641,In_1672);
nor U624 (N_624,In_504,In_665);
nor U625 (N_625,In_1484,In_1598);
or U626 (N_626,In_400,In_1277);
and U627 (N_627,In_93,In_562);
and U628 (N_628,In_333,In_787);
and U629 (N_629,In_643,In_125);
nand U630 (N_630,In_1270,In_642);
nor U631 (N_631,In_1722,In_126);
nor U632 (N_632,In_703,In_1834);
nand U633 (N_633,In_1461,In_666);
nor U634 (N_634,In_1706,In_345);
nand U635 (N_635,In_514,In_946);
xor U636 (N_636,In_1854,In_598);
or U637 (N_637,In_192,In_361);
and U638 (N_638,In_430,In_635);
or U639 (N_639,In_914,In_1933);
nand U640 (N_640,In_1632,In_1442);
nor U641 (N_641,In_1396,In_858);
nor U642 (N_642,In_1094,In_1767);
and U643 (N_643,In_297,In_1088);
or U644 (N_644,In_1878,In_1512);
nor U645 (N_645,In_1756,In_830);
nand U646 (N_646,In_934,In_1694);
xnor U647 (N_647,In_1160,In_974);
and U648 (N_648,In_1812,In_536);
nor U649 (N_649,In_1640,In_840);
nand U650 (N_650,In_644,In_998);
and U651 (N_651,In_1494,In_54);
nor U652 (N_652,In_1888,In_636);
nor U653 (N_653,In_103,In_684);
or U654 (N_654,In_1154,In_124);
and U655 (N_655,In_1239,In_82);
nand U656 (N_656,In_60,In_30);
and U657 (N_657,In_1941,In_91);
and U658 (N_658,In_755,In_1114);
or U659 (N_659,In_557,In_1453);
or U660 (N_660,In_628,In_1872);
or U661 (N_661,In_722,In_116);
or U662 (N_662,In_38,In_1609);
and U663 (N_663,In_1621,In_723);
nand U664 (N_664,In_710,In_424);
or U665 (N_665,In_1282,In_25);
or U666 (N_666,In_1420,In_1853);
nand U667 (N_667,In_1326,In_1718);
nor U668 (N_668,In_513,In_182);
nand U669 (N_669,In_395,In_1089);
and U670 (N_670,In_789,In_1895);
xnor U671 (N_671,In_1474,In_1772);
and U672 (N_672,In_1516,In_1322);
or U673 (N_673,In_454,In_1377);
and U674 (N_674,In_1454,In_1652);
nor U675 (N_675,In_732,In_804);
and U676 (N_676,In_1188,In_738);
and U677 (N_677,In_1858,In_330);
nor U678 (N_678,In_114,In_88);
nand U679 (N_679,In_324,In_1799);
or U680 (N_680,In_327,In_1617);
or U681 (N_681,In_550,In_1750);
and U682 (N_682,In_1063,In_1307);
nand U683 (N_683,In_73,In_700);
nand U684 (N_684,In_177,In_991);
and U685 (N_685,In_1384,In_1097);
or U686 (N_686,In_534,In_216);
xnor U687 (N_687,In_70,In_1083);
nand U688 (N_688,In_368,In_962);
xor U689 (N_689,In_1387,In_1857);
nor U690 (N_690,In_1852,In_405);
nand U691 (N_691,In_1118,In_794);
nor U692 (N_692,In_1119,In_148);
or U693 (N_693,In_195,In_434);
and U694 (N_694,In_492,In_1827);
or U695 (N_695,In_707,In_1923);
nand U696 (N_696,In_1507,In_1446);
or U697 (N_697,In_1012,In_671);
and U698 (N_698,In_752,In_1578);
xor U699 (N_699,In_1284,In_1824);
nand U700 (N_700,In_1417,In_304);
and U701 (N_701,In_1434,In_1714);
and U702 (N_702,In_1826,In_741);
and U703 (N_703,In_220,In_1994);
and U704 (N_704,In_1346,In_567);
nor U705 (N_705,In_173,In_820);
nand U706 (N_706,In_1177,In_300);
or U707 (N_707,In_508,In_1203);
and U708 (N_708,In_734,In_115);
and U709 (N_709,In_1953,In_417);
and U710 (N_710,In_1860,In_143);
or U711 (N_711,In_338,In_1964);
and U712 (N_712,In_1903,In_1343);
nor U713 (N_713,In_568,In_1770);
nor U714 (N_714,In_131,In_578);
nand U715 (N_715,In_1244,In_151);
nor U716 (N_716,In_1877,In_790);
nor U717 (N_717,In_737,In_1221);
and U718 (N_718,In_1560,In_1813);
nor U719 (N_719,In_1349,In_1804);
or U720 (N_720,In_1436,In_744);
nand U721 (N_721,In_1108,In_253);
nand U722 (N_722,In_1534,In_756);
or U723 (N_723,In_119,In_1961);
or U724 (N_724,In_515,In_18);
and U725 (N_725,In_407,In_227);
nand U726 (N_726,In_1039,In_1319);
nand U727 (N_727,In_1927,In_376);
nand U728 (N_728,In_847,In_769);
and U729 (N_729,In_142,In_845);
and U730 (N_730,In_486,In_235);
nor U731 (N_731,In_1645,In_1803);
nor U732 (N_732,In_113,In_1558);
nor U733 (N_733,In_893,In_170);
nor U734 (N_734,In_1170,In_1300);
or U735 (N_735,In_1978,In_1011);
nor U736 (N_736,In_15,In_467);
or U737 (N_737,In_1120,In_1890);
and U738 (N_738,In_1816,In_920);
nand U739 (N_739,In_1055,In_171);
nor U740 (N_740,In_62,In_1753);
nand U741 (N_741,In_1882,In_629);
nor U742 (N_742,In_104,In_990);
nand U743 (N_743,In_418,In_232);
nand U744 (N_744,In_323,In_1596);
nor U745 (N_745,In_1790,In_458);
or U746 (N_746,In_1257,In_1728);
and U747 (N_747,In_1217,In_1379);
and U748 (N_748,In_1344,In_352);
or U749 (N_749,In_713,In_681);
nor U750 (N_750,In_822,In_1225);
nand U751 (N_751,In_1026,In_1115);
nor U752 (N_752,In_662,In_1913);
nand U753 (N_753,In_389,In_1993);
or U754 (N_754,In_85,In_1643);
nor U755 (N_755,In_867,In_570);
nor U756 (N_756,In_1147,In_293);
xnor U757 (N_757,In_1891,In_1298);
xnor U758 (N_758,In_388,In_1831);
or U759 (N_759,In_1671,In_396);
nand U760 (N_760,In_816,In_1898);
or U761 (N_761,In_522,In_140);
nor U762 (N_762,In_1939,In_1421);
and U763 (N_763,In_328,In_1190);
and U764 (N_764,In_259,In_117);
nand U765 (N_765,In_1532,In_1522);
and U766 (N_766,In_1771,In_860);
nor U767 (N_767,In_1090,In_1316);
nand U768 (N_768,In_1364,In_664);
or U769 (N_769,In_1293,In_766);
and U770 (N_770,In_1675,In_201);
or U771 (N_771,In_1835,In_921);
nor U772 (N_772,In_221,In_1468);
nor U773 (N_773,In_731,In_489);
and U774 (N_774,In_69,In_325);
and U775 (N_775,In_443,In_516);
nor U776 (N_776,In_1990,In_1595);
nand U777 (N_777,In_1689,In_1721);
and U778 (N_778,In_144,In_846);
nor U779 (N_779,In_1987,In_1873);
nand U780 (N_780,In_1520,In_275);
nand U781 (N_781,In_899,In_4);
nand U782 (N_782,In_1043,In_86);
or U783 (N_783,In_1711,In_1288);
nand U784 (N_784,In_762,In_948);
or U785 (N_785,In_1124,In_1979);
or U786 (N_786,In_1510,In_1004);
xor U787 (N_787,In_1780,In_1080);
nor U788 (N_788,In_1129,In_1156);
and U789 (N_789,In_425,In_1073);
and U790 (N_790,In_1095,In_208);
or U791 (N_791,In_1199,In_798);
nand U792 (N_792,In_1191,In_1467);
or U793 (N_793,In_270,In_1372);
nor U794 (N_794,In_1386,In_217);
or U795 (N_795,In_614,In_1104);
nand U796 (N_796,In_1237,In_223);
nor U797 (N_797,In_1800,In_1938);
and U798 (N_798,In_48,In_1599);
or U799 (N_799,In_1730,In_584);
and U800 (N_800,In_720,In_207);
and U801 (N_801,In_305,In_1476);
nand U802 (N_802,In_1864,In_39);
nand U803 (N_803,In_656,In_1432);
and U804 (N_804,In_1271,In_1541);
xnor U805 (N_805,In_1698,In_996);
and U806 (N_806,In_1605,In_715);
nor U807 (N_807,In_1112,In_1931);
nand U808 (N_808,In_1587,In_923);
nor U809 (N_809,In_1142,In_911);
nor U810 (N_810,In_1030,In_159);
and U811 (N_811,In_761,In_552);
nand U812 (N_812,In_1946,In_1846);
and U813 (N_813,In_1299,In_1308);
or U814 (N_814,In_924,In_591);
and U815 (N_815,In_1395,In_1841);
nor U816 (N_816,In_1704,In_1475);
and U817 (N_817,In_521,In_1712);
or U818 (N_818,In_172,In_133);
nand U819 (N_819,In_476,In_1648);
nor U820 (N_820,In_406,In_1673);
nand U821 (N_821,In_365,In_670);
or U822 (N_822,In_1815,In_1289);
or U823 (N_823,In_1075,In_863);
nand U824 (N_824,In_802,In_1281);
nand U825 (N_825,In_410,In_942);
nor U826 (N_826,In_1489,In_1260);
or U827 (N_827,In_1586,In_242);
nor U828 (N_828,In_1305,In_586);
nand U829 (N_829,In_1327,In_1908);
xnor U830 (N_830,In_449,In_1763);
or U831 (N_831,In_1027,In_930);
nand U832 (N_832,In_1048,In_837);
nor U833 (N_833,In_836,In_781);
and U834 (N_834,In_970,In_55);
xnor U835 (N_835,In_1205,In_1817);
or U836 (N_836,In_639,In_426);
nand U837 (N_837,In_1057,In_615);
and U838 (N_838,In_1649,In_1010);
or U839 (N_839,In_767,In_1006);
or U840 (N_840,In_1559,In_724);
nand U841 (N_841,In_1367,In_1046);
or U842 (N_842,In_687,In_1897);
nor U843 (N_843,In_1332,In_1991);
or U844 (N_844,In_1155,In_1107);
or U845 (N_845,In_829,In_1949);
nor U846 (N_846,In_1127,In_1413);
or U847 (N_847,In_1936,In_127);
xor U848 (N_848,In_940,In_1342);
or U849 (N_849,In_1851,In_1);
nor U850 (N_850,In_1921,In_1789);
and U851 (N_851,In_1544,In_793);
xor U852 (N_852,In_763,In_1439);
and U853 (N_853,In_488,In_747);
or U854 (N_854,In_1173,In_1658);
nor U855 (N_855,In_1005,In_433);
or U856 (N_856,In_1479,In_193);
nor U857 (N_857,In_1425,In_1887);
nor U858 (N_858,In_726,In_500);
or U859 (N_859,In_1876,In_21);
nor U860 (N_860,In_1385,In_316);
or U861 (N_861,In_1336,In_1007);
nand U862 (N_862,In_37,In_303);
and U863 (N_863,In_228,In_1758);
nand U864 (N_864,In_1511,In_357);
or U865 (N_865,In_1465,In_694);
nand U866 (N_866,In_205,In_1141);
and U867 (N_867,In_1428,In_1423);
and U868 (N_868,In_526,In_58);
xnor U869 (N_869,In_1971,In_1014);
and U870 (N_870,In_892,In_966);
nand U871 (N_871,In_1549,In_1807);
nor U872 (N_872,In_784,In_1373);
or U873 (N_873,In_1303,In_1998);
or U874 (N_874,In_697,In_367);
nor U875 (N_875,In_1754,In_1950);
or U876 (N_876,In_248,In_1334);
and U877 (N_877,In_1955,In_667);
xor U878 (N_878,In_1592,In_977);
or U879 (N_879,In_46,In_880);
and U880 (N_880,In_876,In_659);
and U881 (N_881,In_1121,In_1850);
or U882 (N_882,In_834,In_1295);
or U883 (N_883,In_1723,In_120);
nor U884 (N_884,In_1259,In_1715);
and U885 (N_885,In_759,In_503);
nor U886 (N_886,In_1285,In_1500);
or U887 (N_887,In_1896,In_1339);
nand U888 (N_888,In_841,In_1176);
nand U889 (N_889,In_1752,In_1376);
nand U890 (N_890,In_560,In_826);
or U891 (N_891,In_1985,In_1470);
nand U892 (N_892,In_1412,In_1657);
and U893 (N_893,In_442,In_1031);
and U894 (N_894,In_1591,In_894);
nand U895 (N_895,In_1001,In_1724);
nor U896 (N_896,In_1557,In_918);
and U897 (N_897,In_206,In_1172);
nor U898 (N_898,In_890,In_537);
nor U899 (N_899,In_1690,In_337);
and U900 (N_900,In_1513,In_961);
and U901 (N_901,In_1777,In_1838);
and U902 (N_902,In_204,In_554);
nand U903 (N_903,In_929,In_897);
and U904 (N_904,In_565,In_1597);
or U905 (N_905,In_1060,In_1375);
nor U906 (N_906,In_555,In_868);
and U907 (N_907,In_1382,In_280);
nor U908 (N_908,In_566,In_471);
or U909 (N_909,In_551,In_1140);
nor U910 (N_910,In_1186,In_1407);
nor U911 (N_911,In_1213,In_1594);
nor U912 (N_912,In_80,In_912);
nor U913 (N_913,In_1845,In_1093);
nand U914 (N_914,In_1733,In_1480);
and U915 (N_915,In_1542,In_563);
nand U916 (N_916,In_805,In_107);
nand U917 (N_917,In_1381,In_158);
or U918 (N_918,In_149,In_1736);
and U919 (N_919,In_1265,In_1230);
and U920 (N_920,In_821,In_1146);
or U921 (N_921,In_1471,In_22);
or U922 (N_922,In_532,In_1183);
and U923 (N_923,In_1488,In_135);
xnor U924 (N_924,In_1620,In_1825);
nand U925 (N_925,In_1503,In_84);
nand U926 (N_926,In_618,In_1029);
nor U927 (N_927,In_1496,In_1130);
and U928 (N_928,In_882,In_1821);
or U929 (N_929,In_185,In_808);
and U930 (N_930,In_1311,In_1553);
or U931 (N_931,In_1664,In_992);
or U932 (N_932,In_1786,In_480);
and U933 (N_933,In_832,In_592);
and U934 (N_934,In_1588,In_523);
and U935 (N_935,In_203,In_574);
nand U936 (N_936,In_1087,In_1224);
and U937 (N_937,In_1634,In_1024);
nand U938 (N_938,In_1275,In_138);
or U939 (N_939,In_1574,In_1220);
nand U940 (N_940,In_61,In_411);
xor U941 (N_941,In_1900,In_355);
and U942 (N_942,In_168,In_608);
nand U943 (N_943,In_717,In_408);
nor U944 (N_944,In_1214,In_1518);
or U945 (N_945,In_564,In_340);
xnor U946 (N_946,In_1602,In_776);
and U947 (N_947,In_1633,In_800);
nor U948 (N_948,In_419,In_1975);
xnor U949 (N_949,In_166,In_31);
nor U950 (N_950,In_1204,In_1212);
nand U951 (N_951,In_1879,In_181);
nor U952 (N_952,In_683,In_817);
and U953 (N_953,In_751,In_197);
xnor U954 (N_954,In_1166,In_1656);
and U955 (N_955,In_1545,In_631);
nor U956 (N_956,In_984,In_1047);
or U957 (N_957,In_53,In_965);
or U958 (N_958,In_839,In_219);
nand U959 (N_959,In_289,In_441);
or U960 (N_960,In_165,In_507);
nor U961 (N_961,In_1138,In_465);
or U962 (N_962,In_1833,In_1546);
nor U963 (N_963,In_1952,In_8);
and U964 (N_964,In_520,In_1013);
or U965 (N_965,In_153,In_951);
nor U966 (N_966,In_437,In_1554);
and U967 (N_967,In_579,In_1869);
and U968 (N_968,In_244,In_1340);
and U969 (N_969,In_765,In_865);
nand U970 (N_970,In_1708,In_1370);
or U971 (N_971,In_1460,In_1506);
nand U972 (N_972,In_1143,In_606);
or U973 (N_973,In_1136,In_19);
nor U974 (N_974,In_1925,In_481);
or U975 (N_975,In_661,In_1567);
and U976 (N_976,In_622,In_517);
and U977 (N_977,In_1268,In_1788);
or U978 (N_978,In_1636,In_772);
xor U979 (N_979,In_1976,In_64);
nor U980 (N_980,In_1241,In_1101);
nand U981 (N_981,In_20,In_1693);
or U982 (N_982,In_1049,In_544);
or U983 (N_983,In_851,In_1798);
nand U984 (N_984,In_1526,In_1959);
and U985 (N_985,In_1517,In_1508);
nor U986 (N_986,In_415,In_1743);
nor U987 (N_987,In_1918,In_1431);
and U988 (N_988,In_545,In_864);
nand U989 (N_989,In_1052,In_99);
nor U990 (N_990,In_932,In_857);
nor U991 (N_991,In_714,In_36);
nor U992 (N_992,In_1911,In_1035);
and U993 (N_993,In_590,In_801);
nand U994 (N_994,In_519,In_112);
and U995 (N_995,In_1776,In_1451);
and U996 (N_996,In_749,In_1315);
nand U997 (N_997,In_224,In_332);
nor U998 (N_998,In_129,In_1930);
nand U999 (N_999,In_997,In_548);
xor U1000 (N_1000,In_133,In_1633);
nand U1001 (N_1001,In_1577,In_88);
nand U1002 (N_1002,In_334,In_1773);
and U1003 (N_1003,In_1763,In_1210);
nand U1004 (N_1004,In_807,In_1693);
nor U1005 (N_1005,In_135,In_106);
or U1006 (N_1006,In_362,In_1300);
and U1007 (N_1007,In_712,In_1067);
nand U1008 (N_1008,In_1488,In_1152);
nor U1009 (N_1009,In_516,In_246);
xnor U1010 (N_1010,In_173,In_1898);
nand U1011 (N_1011,In_1583,In_286);
nand U1012 (N_1012,In_809,In_1538);
nor U1013 (N_1013,In_1653,In_221);
or U1014 (N_1014,In_1070,In_1064);
or U1015 (N_1015,In_185,In_1039);
and U1016 (N_1016,In_166,In_438);
and U1017 (N_1017,In_1146,In_1838);
or U1018 (N_1018,In_1427,In_786);
or U1019 (N_1019,In_716,In_1740);
or U1020 (N_1020,In_576,In_830);
nand U1021 (N_1021,In_748,In_498);
nand U1022 (N_1022,In_1991,In_1678);
or U1023 (N_1023,In_1919,In_417);
and U1024 (N_1024,In_1984,In_1887);
nor U1025 (N_1025,In_1637,In_1014);
nor U1026 (N_1026,In_735,In_970);
nor U1027 (N_1027,In_490,In_208);
or U1028 (N_1028,In_1591,In_1515);
nor U1029 (N_1029,In_200,In_1177);
nor U1030 (N_1030,In_1877,In_448);
nor U1031 (N_1031,In_500,In_362);
or U1032 (N_1032,In_648,In_1694);
and U1033 (N_1033,In_490,In_389);
nor U1034 (N_1034,In_1103,In_601);
or U1035 (N_1035,In_578,In_110);
and U1036 (N_1036,In_721,In_1959);
or U1037 (N_1037,In_1825,In_451);
nor U1038 (N_1038,In_466,In_1714);
and U1039 (N_1039,In_624,In_187);
or U1040 (N_1040,In_71,In_109);
nand U1041 (N_1041,In_962,In_1471);
nand U1042 (N_1042,In_830,In_777);
nand U1043 (N_1043,In_1675,In_1756);
nand U1044 (N_1044,In_1487,In_1367);
and U1045 (N_1045,In_832,In_1481);
nand U1046 (N_1046,In_198,In_812);
nor U1047 (N_1047,In_1415,In_310);
and U1048 (N_1048,In_800,In_88);
and U1049 (N_1049,In_1915,In_1549);
or U1050 (N_1050,In_1223,In_1416);
nand U1051 (N_1051,In_1495,In_1821);
and U1052 (N_1052,In_1106,In_317);
nand U1053 (N_1053,In_1267,In_1529);
or U1054 (N_1054,In_389,In_494);
nor U1055 (N_1055,In_877,In_1062);
and U1056 (N_1056,In_559,In_992);
or U1057 (N_1057,In_315,In_1567);
and U1058 (N_1058,In_1846,In_1572);
nand U1059 (N_1059,In_1229,In_704);
or U1060 (N_1060,In_575,In_1685);
nand U1061 (N_1061,In_192,In_418);
or U1062 (N_1062,In_112,In_366);
or U1063 (N_1063,In_1784,In_1663);
nor U1064 (N_1064,In_76,In_1709);
and U1065 (N_1065,In_530,In_140);
and U1066 (N_1066,In_363,In_1635);
and U1067 (N_1067,In_1967,In_953);
nor U1068 (N_1068,In_553,In_500);
nand U1069 (N_1069,In_1853,In_367);
and U1070 (N_1070,In_330,In_452);
or U1071 (N_1071,In_1281,In_1300);
or U1072 (N_1072,In_1521,In_1615);
nor U1073 (N_1073,In_1049,In_927);
or U1074 (N_1074,In_1278,In_1740);
nand U1075 (N_1075,In_636,In_1852);
nor U1076 (N_1076,In_1842,In_588);
xor U1077 (N_1077,In_792,In_1363);
and U1078 (N_1078,In_800,In_793);
and U1079 (N_1079,In_1727,In_1453);
nor U1080 (N_1080,In_1722,In_655);
nand U1081 (N_1081,In_600,In_353);
nand U1082 (N_1082,In_1881,In_49);
and U1083 (N_1083,In_1766,In_1557);
nand U1084 (N_1084,In_150,In_187);
nor U1085 (N_1085,In_1190,In_763);
nand U1086 (N_1086,In_1189,In_441);
and U1087 (N_1087,In_1893,In_218);
and U1088 (N_1088,In_1784,In_500);
nor U1089 (N_1089,In_333,In_1717);
and U1090 (N_1090,In_640,In_1406);
or U1091 (N_1091,In_1603,In_1403);
or U1092 (N_1092,In_847,In_452);
or U1093 (N_1093,In_300,In_1381);
or U1094 (N_1094,In_703,In_1032);
or U1095 (N_1095,In_1094,In_328);
or U1096 (N_1096,In_1318,In_1419);
nand U1097 (N_1097,In_73,In_1968);
nor U1098 (N_1098,In_1155,In_1627);
and U1099 (N_1099,In_1005,In_1046);
or U1100 (N_1100,In_672,In_1916);
nand U1101 (N_1101,In_894,In_868);
nor U1102 (N_1102,In_659,In_1426);
nor U1103 (N_1103,In_1849,In_291);
or U1104 (N_1104,In_168,In_1762);
nand U1105 (N_1105,In_351,In_1155);
or U1106 (N_1106,In_1232,In_529);
and U1107 (N_1107,In_1362,In_552);
nor U1108 (N_1108,In_1866,In_302);
nor U1109 (N_1109,In_282,In_661);
nor U1110 (N_1110,In_1099,In_1853);
nor U1111 (N_1111,In_1765,In_634);
nand U1112 (N_1112,In_316,In_1565);
nor U1113 (N_1113,In_760,In_1350);
or U1114 (N_1114,In_941,In_197);
nor U1115 (N_1115,In_59,In_1448);
nand U1116 (N_1116,In_210,In_653);
nand U1117 (N_1117,In_451,In_1171);
nand U1118 (N_1118,In_1873,In_136);
nand U1119 (N_1119,In_1340,In_473);
nor U1120 (N_1120,In_243,In_749);
nor U1121 (N_1121,In_552,In_765);
nor U1122 (N_1122,In_1453,In_1489);
and U1123 (N_1123,In_1799,In_356);
nand U1124 (N_1124,In_231,In_958);
or U1125 (N_1125,In_1842,In_381);
and U1126 (N_1126,In_515,In_8);
nand U1127 (N_1127,In_102,In_1983);
nor U1128 (N_1128,In_822,In_1062);
nor U1129 (N_1129,In_1807,In_1007);
and U1130 (N_1130,In_630,In_363);
and U1131 (N_1131,In_1785,In_1142);
and U1132 (N_1132,In_394,In_1830);
and U1133 (N_1133,In_252,In_1781);
or U1134 (N_1134,In_666,In_460);
nor U1135 (N_1135,In_1216,In_288);
and U1136 (N_1136,In_1855,In_1156);
nor U1137 (N_1137,In_546,In_150);
and U1138 (N_1138,In_845,In_603);
nor U1139 (N_1139,In_90,In_24);
nor U1140 (N_1140,In_1148,In_1695);
or U1141 (N_1141,In_1089,In_833);
nand U1142 (N_1142,In_1027,In_769);
and U1143 (N_1143,In_1559,In_20);
and U1144 (N_1144,In_659,In_675);
and U1145 (N_1145,In_998,In_652);
nor U1146 (N_1146,In_1815,In_975);
nand U1147 (N_1147,In_254,In_1989);
nor U1148 (N_1148,In_627,In_1022);
nor U1149 (N_1149,In_835,In_853);
nor U1150 (N_1150,In_775,In_1806);
xor U1151 (N_1151,In_920,In_666);
nand U1152 (N_1152,In_1336,In_136);
or U1153 (N_1153,In_1770,In_64);
or U1154 (N_1154,In_1070,In_225);
and U1155 (N_1155,In_1298,In_568);
nor U1156 (N_1156,In_30,In_1026);
nor U1157 (N_1157,In_732,In_54);
and U1158 (N_1158,In_831,In_904);
and U1159 (N_1159,In_707,In_838);
or U1160 (N_1160,In_516,In_1479);
and U1161 (N_1161,In_1741,In_374);
nor U1162 (N_1162,In_1749,In_483);
and U1163 (N_1163,In_988,In_1416);
or U1164 (N_1164,In_971,In_1450);
and U1165 (N_1165,In_524,In_1572);
nor U1166 (N_1166,In_790,In_131);
and U1167 (N_1167,In_1983,In_625);
or U1168 (N_1168,In_173,In_675);
and U1169 (N_1169,In_1923,In_1204);
nor U1170 (N_1170,In_56,In_69);
or U1171 (N_1171,In_576,In_496);
or U1172 (N_1172,In_1763,In_1563);
or U1173 (N_1173,In_45,In_439);
nor U1174 (N_1174,In_1772,In_420);
nand U1175 (N_1175,In_845,In_465);
nand U1176 (N_1176,In_1209,In_167);
and U1177 (N_1177,In_1764,In_258);
nand U1178 (N_1178,In_678,In_252);
or U1179 (N_1179,In_1752,In_1508);
nand U1180 (N_1180,In_166,In_989);
and U1181 (N_1181,In_1826,In_1541);
nand U1182 (N_1182,In_882,In_207);
or U1183 (N_1183,In_1987,In_1054);
nor U1184 (N_1184,In_1610,In_16);
nand U1185 (N_1185,In_789,In_469);
nand U1186 (N_1186,In_1630,In_658);
nor U1187 (N_1187,In_1211,In_1390);
nor U1188 (N_1188,In_1467,In_1049);
and U1189 (N_1189,In_554,In_898);
nor U1190 (N_1190,In_358,In_1977);
nor U1191 (N_1191,In_137,In_832);
nand U1192 (N_1192,In_1227,In_1020);
nand U1193 (N_1193,In_1684,In_745);
or U1194 (N_1194,In_1655,In_1950);
nand U1195 (N_1195,In_613,In_94);
nand U1196 (N_1196,In_551,In_1490);
or U1197 (N_1197,In_451,In_23);
and U1198 (N_1198,In_1741,In_760);
nand U1199 (N_1199,In_147,In_1139);
nor U1200 (N_1200,In_543,In_248);
and U1201 (N_1201,In_1694,In_1398);
nor U1202 (N_1202,In_667,In_472);
and U1203 (N_1203,In_32,In_759);
or U1204 (N_1204,In_1249,In_1490);
or U1205 (N_1205,In_674,In_781);
nand U1206 (N_1206,In_935,In_1944);
or U1207 (N_1207,In_438,In_1193);
nor U1208 (N_1208,In_85,In_1491);
nor U1209 (N_1209,In_419,In_1979);
nand U1210 (N_1210,In_1737,In_1045);
and U1211 (N_1211,In_1686,In_648);
or U1212 (N_1212,In_1856,In_957);
or U1213 (N_1213,In_181,In_911);
nand U1214 (N_1214,In_480,In_746);
nor U1215 (N_1215,In_70,In_943);
nor U1216 (N_1216,In_1936,In_139);
nor U1217 (N_1217,In_731,In_1512);
nor U1218 (N_1218,In_1934,In_258);
or U1219 (N_1219,In_378,In_1156);
and U1220 (N_1220,In_592,In_1);
and U1221 (N_1221,In_1482,In_1405);
or U1222 (N_1222,In_1778,In_1169);
nand U1223 (N_1223,In_172,In_509);
nand U1224 (N_1224,In_1398,In_1249);
nand U1225 (N_1225,In_1077,In_541);
nand U1226 (N_1226,In_1130,In_1104);
nand U1227 (N_1227,In_1041,In_672);
nor U1228 (N_1228,In_894,In_460);
or U1229 (N_1229,In_1794,In_1356);
nand U1230 (N_1230,In_395,In_819);
nand U1231 (N_1231,In_1279,In_1170);
and U1232 (N_1232,In_1684,In_1876);
nor U1233 (N_1233,In_1268,In_620);
nand U1234 (N_1234,In_762,In_415);
nand U1235 (N_1235,In_239,In_100);
nor U1236 (N_1236,In_941,In_1155);
nor U1237 (N_1237,In_1657,In_1165);
nor U1238 (N_1238,In_366,In_1534);
nor U1239 (N_1239,In_1624,In_452);
and U1240 (N_1240,In_1905,In_736);
or U1241 (N_1241,In_1252,In_1232);
nand U1242 (N_1242,In_1166,In_1300);
nor U1243 (N_1243,In_29,In_1971);
nand U1244 (N_1244,In_1586,In_707);
and U1245 (N_1245,In_1705,In_1640);
nand U1246 (N_1246,In_1620,In_1126);
nor U1247 (N_1247,In_1327,In_1622);
or U1248 (N_1248,In_621,In_1216);
and U1249 (N_1249,In_552,In_1678);
and U1250 (N_1250,In_1254,In_1005);
xnor U1251 (N_1251,In_1643,In_105);
xnor U1252 (N_1252,In_811,In_773);
nand U1253 (N_1253,In_1341,In_462);
nand U1254 (N_1254,In_12,In_1394);
nor U1255 (N_1255,In_60,In_47);
nand U1256 (N_1256,In_12,In_51);
nand U1257 (N_1257,In_1634,In_1333);
nor U1258 (N_1258,In_1905,In_1863);
nor U1259 (N_1259,In_856,In_1531);
and U1260 (N_1260,In_1344,In_813);
and U1261 (N_1261,In_1610,In_862);
or U1262 (N_1262,In_1411,In_774);
xnor U1263 (N_1263,In_125,In_913);
nor U1264 (N_1264,In_455,In_1840);
nor U1265 (N_1265,In_1420,In_401);
nor U1266 (N_1266,In_758,In_1846);
or U1267 (N_1267,In_1520,In_1404);
or U1268 (N_1268,In_13,In_708);
nor U1269 (N_1269,In_1889,In_1015);
nand U1270 (N_1270,In_1584,In_1099);
nor U1271 (N_1271,In_1998,In_1230);
and U1272 (N_1272,In_52,In_221);
or U1273 (N_1273,In_1334,In_959);
nand U1274 (N_1274,In_846,In_838);
and U1275 (N_1275,In_872,In_1352);
and U1276 (N_1276,In_1586,In_1987);
and U1277 (N_1277,In_1634,In_1688);
and U1278 (N_1278,In_204,In_1582);
or U1279 (N_1279,In_548,In_1641);
or U1280 (N_1280,In_1315,In_1696);
nand U1281 (N_1281,In_926,In_171);
or U1282 (N_1282,In_1317,In_1465);
or U1283 (N_1283,In_1801,In_1493);
nor U1284 (N_1284,In_168,In_1037);
or U1285 (N_1285,In_292,In_1687);
and U1286 (N_1286,In_1055,In_1532);
nor U1287 (N_1287,In_556,In_1173);
or U1288 (N_1288,In_1981,In_357);
nand U1289 (N_1289,In_1839,In_1337);
nor U1290 (N_1290,In_841,In_1507);
or U1291 (N_1291,In_1748,In_276);
and U1292 (N_1292,In_923,In_660);
or U1293 (N_1293,In_1637,In_1089);
or U1294 (N_1294,In_1732,In_363);
or U1295 (N_1295,In_1661,In_404);
or U1296 (N_1296,In_1822,In_1126);
and U1297 (N_1297,In_1851,In_531);
nor U1298 (N_1298,In_958,In_1145);
or U1299 (N_1299,In_536,In_1056);
or U1300 (N_1300,In_916,In_230);
and U1301 (N_1301,In_419,In_1698);
nand U1302 (N_1302,In_67,In_332);
nand U1303 (N_1303,In_326,In_803);
nand U1304 (N_1304,In_662,In_1367);
and U1305 (N_1305,In_406,In_856);
nand U1306 (N_1306,In_1207,In_1906);
nor U1307 (N_1307,In_129,In_1684);
and U1308 (N_1308,In_580,In_1775);
and U1309 (N_1309,In_287,In_1218);
nand U1310 (N_1310,In_1874,In_952);
or U1311 (N_1311,In_1059,In_485);
nor U1312 (N_1312,In_378,In_1888);
nand U1313 (N_1313,In_167,In_1431);
nor U1314 (N_1314,In_1371,In_1937);
and U1315 (N_1315,In_1230,In_446);
or U1316 (N_1316,In_209,In_1875);
nand U1317 (N_1317,In_236,In_341);
nand U1318 (N_1318,In_1029,In_1521);
and U1319 (N_1319,In_1211,In_1662);
nand U1320 (N_1320,In_581,In_1760);
nor U1321 (N_1321,In_1850,In_1646);
or U1322 (N_1322,In_1852,In_303);
and U1323 (N_1323,In_988,In_845);
or U1324 (N_1324,In_39,In_724);
nor U1325 (N_1325,In_680,In_1851);
or U1326 (N_1326,In_548,In_1964);
nand U1327 (N_1327,In_1401,In_734);
or U1328 (N_1328,In_702,In_1497);
and U1329 (N_1329,In_1986,In_1134);
xnor U1330 (N_1330,In_780,In_1364);
nand U1331 (N_1331,In_761,In_860);
nor U1332 (N_1332,In_1913,In_1805);
and U1333 (N_1333,In_1254,In_1179);
and U1334 (N_1334,In_953,In_1557);
and U1335 (N_1335,In_769,In_621);
nor U1336 (N_1336,In_124,In_1379);
nor U1337 (N_1337,In_315,In_1659);
nor U1338 (N_1338,In_1871,In_882);
nand U1339 (N_1339,In_1073,In_1087);
and U1340 (N_1340,In_1566,In_1761);
nand U1341 (N_1341,In_6,In_1117);
nor U1342 (N_1342,In_1001,In_1330);
and U1343 (N_1343,In_1493,In_998);
and U1344 (N_1344,In_822,In_1493);
nand U1345 (N_1345,In_636,In_1548);
nand U1346 (N_1346,In_384,In_1977);
nand U1347 (N_1347,In_1125,In_1526);
and U1348 (N_1348,In_254,In_586);
or U1349 (N_1349,In_1800,In_1112);
nand U1350 (N_1350,In_852,In_1594);
nor U1351 (N_1351,In_187,In_1444);
nor U1352 (N_1352,In_1542,In_1048);
xor U1353 (N_1353,In_354,In_983);
and U1354 (N_1354,In_880,In_43);
nor U1355 (N_1355,In_51,In_1433);
nor U1356 (N_1356,In_727,In_1884);
or U1357 (N_1357,In_1260,In_332);
nor U1358 (N_1358,In_21,In_705);
nand U1359 (N_1359,In_1195,In_471);
nor U1360 (N_1360,In_294,In_56);
and U1361 (N_1361,In_1624,In_1938);
nand U1362 (N_1362,In_119,In_555);
or U1363 (N_1363,In_972,In_1130);
nor U1364 (N_1364,In_1000,In_488);
nor U1365 (N_1365,In_1206,In_62);
or U1366 (N_1366,In_1532,In_191);
nor U1367 (N_1367,In_126,In_698);
nand U1368 (N_1368,In_251,In_1883);
nor U1369 (N_1369,In_1783,In_981);
nor U1370 (N_1370,In_467,In_1300);
nand U1371 (N_1371,In_1106,In_668);
nand U1372 (N_1372,In_400,In_776);
and U1373 (N_1373,In_1849,In_194);
nand U1374 (N_1374,In_562,In_1891);
or U1375 (N_1375,In_973,In_430);
nand U1376 (N_1376,In_573,In_1923);
nand U1377 (N_1377,In_1210,In_1875);
nor U1378 (N_1378,In_1654,In_422);
nor U1379 (N_1379,In_1014,In_616);
or U1380 (N_1380,In_957,In_1700);
or U1381 (N_1381,In_386,In_1794);
nand U1382 (N_1382,In_624,In_1651);
and U1383 (N_1383,In_1611,In_199);
or U1384 (N_1384,In_1345,In_1241);
and U1385 (N_1385,In_1770,In_39);
nor U1386 (N_1386,In_42,In_1132);
nand U1387 (N_1387,In_86,In_1955);
or U1388 (N_1388,In_1452,In_1087);
nor U1389 (N_1389,In_909,In_1883);
nand U1390 (N_1390,In_1443,In_824);
or U1391 (N_1391,In_655,In_499);
and U1392 (N_1392,In_1532,In_998);
and U1393 (N_1393,In_1910,In_454);
nand U1394 (N_1394,In_256,In_236);
or U1395 (N_1395,In_227,In_1664);
or U1396 (N_1396,In_1138,In_597);
and U1397 (N_1397,In_1698,In_925);
and U1398 (N_1398,In_300,In_961);
nor U1399 (N_1399,In_861,In_480);
or U1400 (N_1400,In_296,In_558);
and U1401 (N_1401,In_580,In_1959);
or U1402 (N_1402,In_264,In_1401);
or U1403 (N_1403,In_1127,In_721);
nand U1404 (N_1404,In_330,In_760);
nor U1405 (N_1405,In_1956,In_622);
nand U1406 (N_1406,In_90,In_784);
nand U1407 (N_1407,In_817,In_1526);
nor U1408 (N_1408,In_550,In_1142);
nand U1409 (N_1409,In_1166,In_428);
xnor U1410 (N_1410,In_921,In_1823);
nand U1411 (N_1411,In_1968,In_342);
nand U1412 (N_1412,In_1155,In_182);
or U1413 (N_1413,In_506,In_1491);
and U1414 (N_1414,In_528,In_1979);
nor U1415 (N_1415,In_55,In_735);
nand U1416 (N_1416,In_1751,In_1812);
or U1417 (N_1417,In_1807,In_163);
nor U1418 (N_1418,In_992,In_101);
nor U1419 (N_1419,In_1524,In_530);
nor U1420 (N_1420,In_1902,In_462);
and U1421 (N_1421,In_43,In_793);
nand U1422 (N_1422,In_333,In_1112);
and U1423 (N_1423,In_1960,In_114);
nor U1424 (N_1424,In_686,In_1932);
nor U1425 (N_1425,In_1800,In_1772);
nand U1426 (N_1426,In_1381,In_703);
nand U1427 (N_1427,In_1667,In_1476);
nand U1428 (N_1428,In_255,In_599);
and U1429 (N_1429,In_842,In_769);
nand U1430 (N_1430,In_1435,In_1252);
and U1431 (N_1431,In_1069,In_998);
xor U1432 (N_1432,In_285,In_1998);
or U1433 (N_1433,In_1563,In_324);
and U1434 (N_1434,In_1236,In_85);
and U1435 (N_1435,In_1731,In_1760);
or U1436 (N_1436,In_1013,In_333);
nor U1437 (N_1437,In_749,In_537);
nor U1438 (N_1438,In_1740,In_902);
nand U1439 (N_1439,In_272,In_1728);
or U1440 (N_1440,In_175,In_412);
and U1441 (N_1441,In_1574,In_320);
nor U1442 (N_1442,In_1482,In_1186);
and U1443 (N_1443,In_1098,In_273);
and U1444 (N_1444,In_497,In_23);
and U1445 (N_1445,In_1385,In_538);
and U1446 (N_1446,In_1572,In_1533);
and U1447 (N_1447,In_1456,In_761);
nor U1448 (N_1448,In_1191,In_1239);
or U1449 (N_1449,In_1122,In_611);
or U1450 (N_1450,In_1775,In_1099);
nand U1451 (N_1451,In_1559,In_919);
or U1452 (N_1452,In_1788,In_20);
nand U1453 (N_1453,In_736,In_518);
nand U1454 (N_1454,In_1189,In_1791);
and U1455 (N_1455,In_1604,In_1704);
xor U1456 (N_1456,In_1143,In_1793);
and U1457 (N_1457,In_1867,In_794);
and U1458 (N_1458,In_1510,In_1414);
or U1459 (N_1459,In_1972,In_1216);
or U1460 (N_1460,In_354,In_969);
and U1461 (N_1461,In_1452,In_1994);
or U1462 (N_1462,In_506,In_1105);
nor U1463 (N_1463,In_432,In_116);
or U1464 (N_1464,In_40,In_794);
or U1465 (N_1465,In_577,In_175);
nand U1466 (N_1466,In_1553,In_1720);
xor U1467 (N_1467,In_1308,In_765);
nor U1468 (N_1468,In_1047,In_1662);
and U1469 (N_1469,In_446,In_143);
or U1470 (N_1470,In_1320,In_1739);
nand U1471 (N_1471,In_1446,In_1076);
or U1472 (N_1472,In_761,In_1349);
nand U1473 (N_1473,In_1004,In_1211);
and U1474 (N_1474,In_1176,In_1058);
or U1475 (N_1475,In_196,In_430);
and U1476 (N_1476,In_1352,In_519);
nand U1477 (N_1477,In_281,In_651);
nor U1478 (N_1478,In_1665,In_1022);
nor U1479 (N_1479,In_1416,In_308);
nor U1480 (N_1480,In_1411,In_1163);
or U1481 (N_1481,In_1861,In_1516);
nor U1482 (N_1482,In_1987,In_529);
or U1483 (N_1483,In_1099,In_1334);
or U1484 (N_1484,In_949,In_79);
and U1485 (N_1485,In_157,In_510);
and U1486 (N_1486,In_1373,In_123);
nor U1487 (N_1487,In_1247,In_1958);
and U1488 (N_1488,In_432,In_1773);
xnor U1489 (N_1489,In_111,In_1340);
and U1490 (N_1490,In_455,In_1413);
nor U1491 (N_1491,In_916,In_1528);
nor U1492 (N_1492,In_1393,In_1869);
or U1493 (N_1493,In_1016,In_1968);
nand U1494 (N_1494,In_1603,In_430);
nor U1495 (N_1495,In_1284,In_299);
nand U1496 (N_1496,In_1504,In_1893);
and U1497 (N_1497,In_1566,In_1970);
nand U1498 (N_1498,In_166,In_608);
nand U1499 (N_1499,In_599,In_884);
nand U1500 (N_1500,In_1609,In_982);
nor U1501 (N_1501,In_1940,In_756);
and U1502 (N_1502,In_1571,In_1058);
nand U1503 (N_1503,In_331,In_268);
and U1504 (N_1504,In_457,In_1146);
nor U1505 (N_1505,In_1308,In_37);
nand U1506 (N_1506,In_1941,In_1533);
nor U1507 (N_1507,In_28,In_1721);
or U1508 (N_1508,In_186,In_1960);
nand U1509 (N_1509,In_1473,In_1301);
or U1510 (N_1510,In_373,In_1929);
or U1511 (N_1511,In_1155,In_1339);
nand U1512 (N_1512,In_296,In_1686);
or U1513 (N_1513,In_679,In_243);
or U1514 (N_1514,In_197,In_1853);
and U1515 (N_1515,In_1235,In_927);
nand U1516 (N_1516,In_23,In_155);
xor U1517 (N_1517,In_590,In_1893);
and U1518 (N_1518,In_618,In_472);
nand U1519 (N_1519,In_710,In_138);
nand U1520 (N_1520,In_143,In_759);
or U1521 (N_1521,In_782,In_866);
nand U1522 (N_1522,In_935,In_1592);
or U1523 (N_1523,In_257,In_864);
or U1524 (N_1524,In_1216,In_1004);
or U1525 (N_1525,In_1569,In_217);
nand U1526 (N_1526,In_568,In_948);
and U1527 (N_1527,In_34,In_584);
nand U1528 (N_1528,In_1927,In_1111);
nor U1529 (N_1529,In_63,In_1791);
or U1530 (N_1530,In_529,In_1905);
nand U1531 (N_1531,In_344,In_184);
or U1532 (N_1532,In_268,In_1455);
nand U1533 (N_1533,In_1305,In_1426);
nand U1534 (N_1534,In_8,In_918);
or U1535 (N_1535,In_1182,In_1871);
nand U1536 (N_1536,In_997,In_1455);
nand U1537 (N_1537,In_1695,In_1277);
and U1538 (N_1538,In_1598,In_1569);
nor U1539 (N_1539,In_1610,In_1053);
nand U1540 (N_1540,In_400,In_770);
nand U1541 (N_1541,In_570,In_796);
xor U1542 (N_1542,In_163,In_1948);
or U1543 (N_1543,In_920,In_1349);
and U1544 (N_1544,In_1840,In_1343);
or U1545 (N_1545,In_577,In_943);
nand U1546 (N_1546,In_1785,In_1318);
and U1547 (N_1547,In_1425,In_1014);
or U1548 (N_1548,In_569,In_1938);
and U1549 (N_1549,In_274,In_90);
nor U1550 (N_1550,In_573,In_1473);
nand U1551 (N_1551,In_1822,In_324);
or U1552 (N_1552,In_1294,In_220);
and U1553 (N_1553,In_998,In_476);
or U1554 (N_1554,In_1530,In_784);
nor U1555 (N_1555,In_1780,In_242);
or U1556 (N_1556,In_985,In_1183);
or U1557 (N_1557,In_1485,In_133);
nor U1558 (N_1558,In_1668,In_807);
or U1559 (N_1559,In_1939,In_1206);
nand U1560 (N_1560,In_1949,In_1228);
nand U1561 (N_1561,In_1173,In_212);
and U1562 (N_1562,In_1974,In_948);
and U1563 (N_1563,In_1143,In_249);
nor U1564 (N_1564,In_1358,In_245);
or U1565 (N_1565,In_1980,In_845);
nand U1566 (N_1566,In_230,In_1920);
nand U1567 (N_1567,In_1911,In_1061);
nor U1568 (N_1568,In_1943,In_260);
and U1569 (N_1569,In_1441,In_1103);
nor U1570 (N_1570,In_526,In_1467);
nand U1571 (N_1571,In_1459,In_1122);
nand U1572 (N_1572,In_1100,In_174);
nand U1573 (N_1573,In_229,In_223);
and U1574 (N_1574,In_1966,In_1590);
and U1575 (N_1575,In_560,In_670);
and U1576 (N_1576,In_637,In_1280);
and U1577 (N_1577,In_630,In_207);
or U1578 (N_1578,In_1739,In_1945);
or U1579 (N_1579,In_416,In_202);
or U1580 (N_1580,In_1819,In_135);
or U1581 (N_1581,In_1334,In_1669);
nand U1582 (N_1582,In_1662,In_973);
or U1583 (N_1583,In_1332,In_18);
and U1584 (N_1584,In_1440,In_1895);
or U1585 (N_1585,In_1856,In_1027);
or U1586 (N_1586,In_1875,In_1044);
nand U1587 (N_1587,In_1240,In_33);
nor U1588 (N_1588,In_433,In_1403);
nand U1589 (N_1589,In_782,In_35);
and U1590 (N_1590,In_505,In_1176);
or U1591 (N_1591,In_1620,In_672);
or U1592 (N_1592,In_1846,In_1492);
nand U1593 (N_1593,In_1318,In_1340);
nor U1594 (N_1594,In_515,In_1617);
nand U1595 (N_1595,In_396,In_322);
xnor U1596 (N_1596,In_1973,In_1841);
nand U1597 (N_1597,In_902,In_212);
or U1598 (N_1598,In_357,In_1391);
or U1599 (N_1599,In_1566,In_1801);
or U1600 (N_1600,In_1625,In_1913);
and U1601 (N_1601,In_116,In_894);
xor U1602 (N_1602,In_313,In_1416);
and U1603 (N_1603,In_1626,In_1027);
nor U1604 (N_1604,In_937,In_1444);
or U1605 (N_1605,In_974,In_1013);
nor U1606 (N_1606,In_292,In_487);
or U1607 (N_1607,In_890,In_358);
and U1608 (N_1608,In_1629,In_1098);
and U1609 (N_1609,In_1284,In_1526);
nand U1610 (N_1610,In_1371,In_610);
nand U1611 (N_1611,In_644,In_6);
or U1612 (N_1612,In_77,In_914);
nor U1613 (N_1613,In_378,In_38);
nand U1614 (N_1614,In_1835,In_1853);
nor U1615 (N_1615,In_194,In_1003);
nor U1616 (N_1616,In_864,In_730);
nand U1617 (N_1617,In_258,In_1585);
or U1618 (N_1618,In_437,In_1177);
nand U1619 (N_1619,In_1940,In_248);
nand U1620 (N_1620,In_1559,In_1820);
nand U1621 (N_1621,In_169,In_825);
nor U1622 (N_1622,In_585,In_764);
nor U1623 (N_1623,In_1633,In_1614);
or U1624 (N_1624,In_731,In_940);
nand U1625 (N_1625,In_494,In_536);
nor U1626 (N_1626,In_794,In_1417);
nor U1627 (N_1627,In_706,In_525);
nand U1628 (N_1628,In_1233,In_488);
or U1629 (N_1629,In_1617,In_1579);
nor U1630 (N_1630,In_1565,In_1311);
or U1631 (N_1631,In_794,In_319);
and U1632 (N_1632,In_182,In_7);
nand U1633 (N_1633,In_1096,In_1711);
or U1634 (N_1634,In_426,In_1622);
nor U1635 (N_1635,In_718,In_307);
and U1636 (N_1636,In_862,In_504);
and U1637 (N_1637,In_1521,In_916);
nand U1638 (N_1638,In_602,In_1143);
and U1639 (N_1639,In_1194,In_1867);
and U1640 (N_1640,In_1596,In_1518);
nor U1641 (N_1641,In_227,In_6);
or U1642 (N_1642,In_1731,In_1286);
nand U1643 (N_1643,In_1822,In_862);
nor U1644 (N_1644,In_1774,In_1133);
nor U1645 (N_1645,In_1374,In_38);
nand U1646 (N_1646,In_256,In_1500);
nor U1647 (N_1647,In_1312,In_125);
and U1648 (N_1648,In_387,In_1370);
nor U1649 (N_1649,In_1969,In_201);
and U1650 (N_1650,In_1046,In_1470);
nor U1651 (N_1651,In_1485,In_1062);
nand U1652 (N_1652,In_143,In_1262);
nor U1653 (N_1653,In_237,In_399);
nand U1654 (N_1654,In_1530,In_1212);
nand U1655 (N_1655,In_1959,In_1706);
nand U1656 (N_1656,In_872,In_1553);
nand U1657 (N_1657,In_1897,In_1858);
nand U1658 (N_1658,In_1280,In_1831);
nor U1659 (N_1659,In_690,In_600);
nor U1660 (N_1660,In_775,In_253);
nand U1661 (N_1661,In_577,In_300);
or U1662 (N_1662,In_481,In_1624);
and U1663 (N_1663,In_1497,In_108);
nand U1664 (N_1664,In_821,In_220);
or U1665 (N_1665,In_397,In_1895);
and U1666 (N_1666,In_759,In_683);
and U1667 (N_1667,In_124,In_1968);
or U1668 (N_1668,In_521,In_230);
nand U1669 (N_1669,In_220,In_1978);
or U1670 (N_1670,In_225,In_108);
and U1671 (N_1671,In_549,In_1927);
and U1672 (N_1672,In_311,In_1304);
or U1673 (N_1673,In_1781,In_325);
and U1674 (N_1674,In_155,In_222);
nand U1675 (N_1675,In_1389,In_71);
nor U1676 (N_1676,In_1354,In_763);
and U1677 (N_1677,In_1536,In_199);
and U1678 (N_1678,In_30,In_1396);
or U1679 (N_1679,In_47,In_61);
or U1680 (N_1680,In_1037,In_1154);
nand U1681 (N_1681,In_1442,In_1181);
nor U1682 (N_1682,In_211,In_943);
and U1683 (N_1683,In_1341,In_695);
or U1684 (N_1684,In_1300,In_1358);
or U1685 (N_1685,In_1118,In_401);
nand U1686 (N_1686,In_1861,In_480);
nand U1687 (N_1687,In_639,In_450);
and U1688 (N_1688,In_281,In_319);
or U1689 (N_1689,In_727,In_215);
and U1690 (N_1690,In_592,In_474);
nand U1691 (N_1691,In_1574,In_246);
and U1692 (N_1692,In_223,In_1754);
nor U1693 (N_1693,In_1895,In_1183);
and U1694 (N_1694,In_731,In_1641);
and U1695 (N_1695,In_1179,In_1102);
nor U1696 (N_1696,In_523,In_335);
nand U1697 (N_1697,In_382,In_178);
nor U1698 (N_1698,In_1202,In_1324);
nor U1699 (N_1699,In_435,In_1361);
nand U1700 (N_1700,In_1409,In_1823);
nand U1701 (N_1701,In_1538,In_524);
or U1702 (N_1702,In_1712,In_757);
or U1703 (N_1703,In_1647,In_1918);
or U1704 (N_1704,In_1131,In_1346);
nand U1705 (N_1705,In_191,In_1171);
xnor U1706 (N_1706,In_971,In_1153);
and U1707 (N_1707,In_1085,In_1647);
or U1708 (N_1708,In_1355,In_1956);
nor U1709 (N_1709,In_499,In_309);
or U1710 (N_1710,In_568,In_1904);
nor U1711 (N_1711,In_144,In_362);
nor U1712 (N_1712,In_1864,In_1852);
xnor U1713 (N_1713,In_1884,In_1774);
nand U1714 (N_1714,In_1539,In_1104);
or U1715 (N_1715,In_994,In_1007);
nand U1716 (N_1716,In_1363,In_827);
nor U1717 (N_1717,In_1860,In_810);
and U1718 (N_1718,In_1600,In_557);
or U1719 (N_1719,In_524,In_1712);
and U1720 (N_1720,In_357,In_918);
nor U1721 (N_1721,In_877,In_1107);
nor U1722 (N_1722,In_1627,In_1432);
xnor U1723 (N_1723,In_419,In_1428);
or U1724 (N_1724,In_581,In_1831);
or U1725 (N_1725,In_122,In_346);
or U1726 (N_1726,In_421,In_1641);
or U1727 (N_1727,In_558,In_761);
nand U1728 (N_1728,In_1980,In_711);
and U1729 (N_1729,In_695,In_344);
nor U1730 (N_1730,In_735,In_327);
nand U1731 (N_1731,In_1505,In_56);
or U1732 (N_1732,In_1321,In_1986);
or U1733 (N_1733,In_397,In_155);
nor U1734 (N_1734,In_841,In_1734);
nand U1735 (N_1735,In_1294,In_639);
or U1736 (N_1736,In_1187,In_1953);
nor U1737 (N_1737,In_755,In_675);
nand U1738 (N_1738,In_452,In_1652);
nand U1739 (N_1739,In_879,In_59);
or U1740 (N_1740,In_1153,In_788);
xor U1741 (N_1741,In_139,In_1700);
or U1742 (N_1742,In_605,In_1842);
xnor U1743 (N_1743,In_568,In_1439);
xnor U1744 (N_1744,In_1279,In_968);
and U1745 (N_1745,In_1703,In_1549);
or U1746 (N_1746,In_585,In_402);
nand U1747 (N_1747,In_1914,In_1911);
or U1748 (N_1748,In_1953,In_331);
or U1749 (N_1749,In_1426,In_1227);
nand U1750 (N_1750,In_1735,In_862);
or U1751 (N_1751,In_798,In_956);
and U1752 (N_1752,In_1226,In_1789);
or U1753 (N_1753,In_235,In_1097);
nor U1754 (N_1754,In_697,In_257);
and U1755 (N_1755,In_779,In_1669);
nor U1756 (N_1756,In_219,In_1961);
or U1757 (N_1757,In_451,In_442);
and U1758 (N_1758,In_27,In_79);
xnor U1759 (N_1759,In_1667,In_1326);
nand U1760 (N_1760,In_1361,In_1508);
nor U1761 (N_1761,In_337,In_407);
nand U1762 (N_1762,In_1532,In_507);
and U1763 (N_1763,In_1270,In_1080);
nor U1764 (N_1764,In_1870,In_1474);
xnor U1765 (N_1765,In_1004,In_1285);
and U1766 (N_1766,In_1404,In_1195);
and U1767 (N_1767,In_1816,In_1858);
nand U1768 (N_1768,In_304,In_1377);
and U1769 (N_1769,In_469,In_658);
or U1770 (N_1770,In_519,In_1279);
nand U1771 (N_1771,In_1916,In_1370);
and U1772 (N_1772,In_926,In_511);
or U1773 (N_1773,In_1192,In_1339);
or U1774 (N_1774,In_1168,In_718);
and U1775 (N_1775,In_901,In_1227);
nand U1776 (N_1776,In_1547,In_382);
nor U1777 (N_1777,In_1822,In_1007);
nand U1778 (N_1778,In_319,In_146);
nand U1779 (N_1779,In_1483,In_1313);
and U1780 (N_1780,In_1781,In_379);
nor U1781 (N_1781,In_235,In_905);
nand U1782 (N_1782,In_49,In_447);
or U1783 (N_1783,In_1418,In_1360);
nor U1784 (N_1784,In_1187,In_1022);
nor U1785 (N_1785,In_447,In_101);
nand U1786 (N_1786,In_1537,In_384);
and U1787 (N_1787,In_849,In_1223);
nand U1788 (N_1788,In_798,In_346);
or U1789 (N_1789,In_1647,In_545);
nor U1790 (N_1790,In_1903,In_1368);
and U1791 (N_1791,In_411,In_1733);
nand U1792 (N_1792,In_1660,In_1957);
nor U1793 (N_1793,In_1944,In_389);
nor U1794 (N_1794,In_1954,In_1583);
and U1795 (N_1795,In_1990,In_1189);
or U1796 (N_1796,In_43,In_1483);
or U1797 (N_1797,In_1095,In_790);
nand U1798 (N_1798,In_976,In_639);
and U1799 (N_1799,In_1061,In_67);
and U1800 (N_1800,In_1472,In_1494);
or U1801 (N_1801,In_1415,In_1692);
or U1802 (N_1802,In_824,In_738);
and U1803 (N_1803,In_1721,In_744);
nand U1804 (N_1804,In_1739,In_1360);
nand U1805 (N_1805,In_1950,In_755);
or U1806 (N_1806,In_718,In_712);
nand U1807 (N_1807,In_1564,In_489);
and U1808 (N_1808,In_1507,In_1962);
or U1809 (N_1809,In_30,In_454);
and U1810 (N_1810,In_910,In_1784);
nor U1811 (N_1811,In_592,In_1955);
or U1812 (N_1812,In_27,In_864);
nand U1813 (N_1813,In_0,In_762);
nor U1814 (N_1814,In_439,In_600);
nand U1815 (N_1815,In_126,In_564);
and U1816 (N_1816,In_1511,In_171);
nor U1817 (N_1817,In_1796,In_1841);
nor U1818 (N_1818,In_1312,In_699);
or U1819 (N_1819,In_105,In_1478);
or U1820 (N_1820,In_363,In_414);
nor U1821 (N_1821,In_742,In_1290);
or U1822 (N_1822,In_1863,In_636);
nor U1823 (N_1823,In_1576,In_371);
and U1824 (N_1824,In_1743,In_1690);
nand U1825 (N_1825,In_1968,In_1770);
xnor U1826 (N_1826,In_438,In_1470);
and U1827 (N_1827,In_597,In_1995);
or U1828 (N_1828,In_1487,In_3);
and U1829 (N_1829,In_231,In_1119);
or U1830 (N_1830,In_761,In_1372);
nand U1831 (N_1831,In_339,In_561);
or U1832 (N_1832,In_1047,In_689);
nand U1833 (N_1833,In_197,In_1737);
nand U1834 (N_1834,In_705,In_1810);
and U1835 (N_1835,In_1915,In_46);
nor U1836 (N_1836,In_156,In_1269);
or U1837 (N_1837,In_1149,In_1757);
or U1838 (N_1838,In_1497,In_1012);
and U1839 (N_1839,In_580,In_776);
nand U1840 (N_1840,In_621,In_1340);
nor U1841 (N_1841,In_357,In_1462);
nor U1842 (N_1842,In_1443,In_35);
nor U1843 (N_1843,In_867,In_815);
and U1844 (N_1844,In_98,In_839);
or U1845 (N_1845,In_1731,In_729);
or U1846 (N_1846,In_1456,In_134);
nand U1847 (N_1847,In_165,In_1608);
nand U1848 (N_1848,In_408,In_1094);
or U1849 (N_1849,In_897,In_1748);
or U1850 (N_1850,In_1963,In_1357);
or U1851 (N_1851,In_1298,In_634);
nor U1852 (N_1852,In_72,In_1900);
xnor U1853 (N_1853,In_1840,In_1110);
or U1854 (N_1854,In_969,In_1217);
or U1855 (N_1855,In_349,In_273);
nand U1856 (N_1856,In_1397,In_634);
and U1857 (N_1857,In_1577,In_797);
and U1858 (N_1858,In_1751,In_1966);
and U1859 (N_1859,In_410,In_171);
nor U1860 (N_1860,In_663,In_1322);
or U1861 (N_1861,In_271,In_726);
nand U1862 (N_1862,In_256,In_1425);
and U1863 (N_1863,In_1452,In_792);
nand U1864 (N_1864,In_510,In_809);
nor U1865 (N_1865,In_998,In_1398);
nand U1866 (N_1866,In_1305,In_465);
and U1867 (N_1867,In_1415,In_1080);
and U1868 (N_1868,In_924,In_1317);
or U1869 (N_1869,In_776,In_1097);
and U1870 (N_1870,In_720,In_1786);
xnor U1871 (N_1871,In_1377,In_579);
nor U1872 (N_1872,In_1675,In_800);
nor U1873 (N_1873,In_1395,In_1659);
nor U1874 (N_1874,In_1679,In_199);
nor U1875 (N_1875,In_1375,In_1233);
xnor U1876 (N_1876,In_7,In_548);
nor U1877 (N_1877,In_1532,In_1556);
nand U1878 (N_1878,In_1987,In_419);
and U1879 (N_1879,In_956,In_1551);
nand U1880 (N_1880,In_1331,In_1470);
nor U1881 (N_1881,In_990,In_776);
nand U1882 (N_1882,In_956,In_1015);
nand U1883 (N_1883,In_1121,In_626);
and U1884 (N_1884,In_1033,In_1848);
nor U1885 (N_1885,In_671,In_1292);
or U1886 (N_1886,In_877,In_746);
or U1887 (N_1887,In_1455,In_1981);
or U1888 (N_1888,In_122,In_251);
and U1889 (N_1889,In_1600,In_1258);
nand U1890 (N_1890,In_1659,In_1617);
or U1891 (N_1891,In_158,In_613);
nor U1892 (N_1892,In_1792,In_1469);
or U1893 (N_1893,In_1736,In_1663);
nand U1894 (N_1894,In_55,In_450);
and U1895 (N_1895,In_1672,In_399);
or U1896 (N_1896,In_716,In_308);
nand U1897 (N_1897,In_957,In_321);
nand U1898 (N_1898,In_1494,In_1888);
nand U1899 (N_1899,In_870,In_1157);
and U1900 (N_1900,In_269,In_1590);
nor U1901 (N_1901,In_439,In_1551);
or U1902 (N_1902,In_546,In_970);
nand U1903 (N_1903,In_805,In_908);
nor U1904 (N_1904,In_655,In_198);
and U1905 (N_1905,In_1400,In_300);
nor U1906 (N_1906,In_910,In_804);
nand U1907 (N_1907,In_63,In_1623);
nand U1908 (N_1908,In_1067,In_717);
nand U1909 (N_1909,In_1677,In_1078);
or U1910 (N_1910,In_104,In_442);
nand U1911 (N_1911,In_1019,In_1541);
nor U1912 (N_1912,In_189,In_1486);
or U1913 (N_1913,In_65,In_1405);
nor U1914 (N_1914,In_992,In_1467);
and U1915 (N_1915,In_242,In_1822);
nand U1916 (N_1916,In_1961,In_641);
nor U1917 (N_1917,In_787,In_1307);
or U1918 (N_1918,In_1699,In_1580);
nor U1919 (N_1919,In_723,In_941);
or U1920 (N_1920,In_957,In_1943);
nor U1921 (N_1921,In_1181,In_1464);
nor U1922 (N_1922,In_335,In_899);
or U1923 (N_1923,In_547,In_1034);
nor U1924 (N_1924,In_1572,In_1268);
and U1925 (N_1925,In_1440,In_291);
nor U1926 (N_1926,In_1049,In_1119);
nand U1927 (N_1927,In_459,In_204);
xnor U1928 (N_1928,In_695,In_15);
nor U1929 (N_1929,In_1820,In_1578);
nor U1930 (N_1930,In_1261,In_965);
nand U1931 (N_1931,In_1221,In_502);
xnor U1932 (N_1932,In_60,In_1244);
nor U1933 (N_1933,In_1551,In_1851);
and U1934 (N_1934,In_1236,In_1767);
and U1935 (N_1935,In_538,In_1674);
and U1936 (N_1936,In_204,In_387);
and U1937 (N_1937,In_1989,In_1853);
nand U1938 (N_1938,In_1056,In_286);
nor U1939 (N_1939,In_1965,In_946);
and U1940 (N_1940,In_1200,In_672);
nand U1941 (N_1941,In_1517,In_464);
nand U1942 (N_1942,In_1133,In_172);
nand U1943 (N_1943,In_64,In_274);
and U1944 (N_1944,In_1029,In_1272);
or U1945 (N_1945,In_1238,In_1957);
nand U1946 (N_1946,In_738,In_1552);
nor U1947 (N_1947,In_809,In_1561);
and U1948 (N_1948,In_1839,In_1694);
and U1949 (N_1949,In_923,In_1061);
nor U1950 (N_1950,In_366,In_1198);
nor U1951 (N_1951,In_849,In_1310);
nand U1952 (N_1952,In_780,In_226);
nand U1953 (N_1953,In_690,In_351);
nor U1954 (N_1954,In_1822,In_805);
and U1955 (N_1955,In_850,In_177);
xor U1956 (N_1956,In_1381,In_1728);
and U1957 (N_1957,In_1430,In_1658);
xor U1958 (N_1958,In_98,In_1575);
nor U1959 (N_1959,In_518,In_654);
and U1960 (N_1960,In_1517,In_569);
or U1961 (N_1961,In_458,In_1285);
or U1962 (N_1962,In_248,In_1319);
and U1963 (N_1963,In_1270,In_1553);
and U1964 (N_1964,In_1901,In_1294);
and U1965 (N_1965,In_1147,In_96);
nor U1966 (N_1966,In_938,In_1997);
and U1967 (N_1967,In_379,In_152);
and U1968 (N_1968,In_932,In_278);
nand U1969 (N_1969,In_92,In_298);
xnor U1970 (N_1970,In_841,In_1396);
nor U1971 (N_1971,In_624,In_1830);
and U1972 (N_1972,In_350,In_1534);
nor U1973 (N_1973,In_340,In_797);
nand U1974 (N_1974,In_1384,In_1129);
or U1975 (N_1975,In_1848,In_1305);
nand U1976 (N_1976,In_580,In_864);
nor U1977 (N_1977,In_1404,In_1800);
or U1978 (N_1978,In_936,In_1642);
nor U1979 (N_1979,In_1644,In_1119);
nor U1980 (N_1980,In_1311,In_593);
nand U1981 (N_1981,In_976,In_1252);
and U1982 (N_1982,In_1435,In_806);
or U1983 (N_1983,In_389,In_1253);
and U1984 (N_1984,In_47,In_1650);
nand U1985 (N_1985,In_940,In_67);
and U1986 (N_1986,In_1345,In_480);
nor U1987 (N_1987,In_1268,In_575);
or U1988 (N_1988,In_1221,In_3);
nand U1989 (N_1989,In_588,In_695);
and U1990 (N_1990,In_936,In_683);
nand U1991 (N_1991,In_737,In_6);
nor U1992 (N_1992,In_285,In_1739);
nor U1993 (N_1993,In_923,In_1259);
and U1994 (N_1994,In_1721,In_237);
and U1995 (N_1995,In_528,In_957);
nor U1996 (N_1996,In_299,In_188);
and U1997 (N_1997,In_1172,In_1986);
or U1998 (N_1998,In_632,In_517);
and U1999 (N_1999,In_1524,In_1533);
nand U2000 (N_2000,In_1447,In_616);
nor U2001 (N_2001,In_1349,In_116);
or U2002 (N_2002,In_625,In_1017);
and U2003 (N_2003,In_25,In_1153);
and U2004 (N_2004,In_1486,In_1544);
or U2005 (N_2005,In_1641,In_581);
or U2006 (N_2006,In_1840,In_1938);
xnor U2007 (N_2007,In_1540,In_1760);
or U2008 (N_2008,In_1734,In_721);
and U2009 (N_2009,In_359,In_796);
nor U2010 (N_2010,In_393,In_1264);
nor U2011 (N_2011,In_561,In_628);
nand U2012 (N_2012,In_1062,In_165);
nor U2013 (N_2013,In_692,In_22);
nor U2014 (N_2014,In_365,In_1729);
or U2015 (N_2015,In_865,In_1359);
nor U2016 (N_2016,In_402,In_381);
and U2017 (N_2017,In_1288,In_940);
xnor U2018 (N_2018,In_1541,In_217);
and U2019 (N_2019,In_589,In_134);
xnor U2020 (N_2020,In_1239,In_1279);
and U2021 (N_2021,In_515,In_1050);
nor U2022 (N_2022,In_1696,In_518);
nand U2023 (N_2023,In_52,In_21);
or U2024 (N_2024,In_923,In_732);
or U2025 (N_2025,In_1300,In_1805);
or U2026 (N_2026,In_1734,In_1244);
nor U2027 (N_2027,In_1093,In_1728);
and U2028 (N_2028,In_431,In_1033);
nand U2029 (N_2029,In_218,In_1475);
or U2030 (N_2030,In_1879,In_418);
nand U2031 (N_2031,In_1848,In_1103);
nor U2032 (N_2032,In_1207,In_660);
nand U2033 (N_2033,In_1946,In_867);
nor U2034 (N_2034,In_1821,In_1405);
or U2035 (N_2035,In_478,In_601);
or U2036 (N_2036,In_935,In_1411);
or U2037 (N_2037,In_540,In_1454);
and U2038 (N_2038,In_842,In_69);
nor U2039 (N_2039,In_541,In_104);
or U2040 (N_2040,In_91,In_448);
xnor U2041 (N_2041,In_1821,In_726);
nor U2042 (N_2042,In_626,In_1430);
nor U2043 (N_2043,In_450,In_1149);
nand U2044 (N_2044,In_695,In_1227);
nand U2045 (N_2045,In_1172,In_1163);
nor U2046 (N_2046,In_1592,In_779);
nand U2047 (N_2047,In_1950,In_1968);
nor U2048 (N_2048,In_1170,In_1160);
xnor U2049 (N_2049,In_240,In_542);
and U2050 (N_2050,In_105,In_1349);
and U2051 (N_2051,In_430,In_759);
and U2052 (N_2052,In_87,In_1637);
and U2053 (N_2053,In_1407,In_1845);
nor U2054 (N_2054,In_1108,In_822);
and U2055 (N_2055,In_907,In_959);
or U2056 (N_2056,In_367,In_1797);
nor U2057 (N_2057,In_792,In_1762);
or U2058 (N_2058,In_1610,In_790);
nand U2059 (N_2059,In_257,In_1947);
nor U2060 (N_2060,In_817,In_1601);
nor U2061 (N_2061,In_1309,In_1864);
nor U2062 (N_2062,In_1993,In_22);
nor U2063 (N_2063,In_1778,In_665);
nand U2064 (N_2064,In_186,In_645);
nand U2065 (N_2065,In_1867,In_536);
or U2066 (N_2066,In_859,In_1550);
and U2067 (N_2067,In_1326,In_358);
and U2068 (N_2068,In_1310,In_498);
nand U2069 (N_2069,In_15,In_605);
nand U2070 (N_2070,In_635,In_367);
nand U2071 (N_2071,In_1499,In_1840);
or U2072 (N_2072,In_129,In_351);
or U2073 (N_2073,In_1603,In_200);
or U2074 (N_2074,In_796,In_918);
nand U2075 (N_2075,In_1712,In_1975);
and U2076 (N_2076,In_111,In_1576);
or U2077 (N_2077,In_1384,In_981);
nand U2078 (N_2078,In_1721,In_465);
or U2079 (N_2079,In_617,In_577);
nand U2080 (N_2080,In_949,In_890);
or U2081 (N_2081,In_1876,In_365);
or U2082 (N_2082,In_1126,In_858);
nor U2083 (N_2083,In_968,In_637);
nor U2084 (N_2084,In_655,In_1510);
and U2085 (N_2085,In_1424,In_119);
xnor U2086 (N_2086,In_608,In_803);
or U2087 (N_2087,In_675,In_171);
and U2088 (N_2088,In_291,In_403);
and U2089 (N_2089,In_1136,In_1976);
and U2090 (N_2090,In_1363,In_1739);
or U2091 (N_2091,In_931,In_591);
or U2092 (N_2092,In_781,In_1026);
nand U2093 (N_2093,In_580,In_419);
and U2094 (N_2094,In_1676,In_364);
or U2095 (N_2095,In_207,In_398);
and U2096 (N_2096,In_1053,In_867);
or U2097 (N_2097,In_719,In_1442);
nand U2098 (N_2098,In_1272,In_506);
or U2099 (N_2099,In_1536,In_1619);
nand U2100 (N_2100,In_1297,In_199);
nand U2101 (N_2101,In_776,In_274);
or U2102 (N_2102,In_1855,In_1177);
nand U2103 (N_2103,In_1802,In_1535);
or U2104 (N_2104,In_1756,In_1356);
and U2105 (N_2105,In_1663,In_515);
nand U2106 (N_2106,In_191,In_224);
or U2107 (N_2107,In_1065,In_414);
xnor U2108 (N_2108,In_1163,In_1973);
nand U2109 (N_2109,In_181,In_1375);
nand U2110 (N_2110,In_914,In_915);
or U2111 (N_2111,In_1729,In_142);
or U2112 (N_2112,In_1049,In_330);
and U2113 (N_2113,In_1663,In_1577);
or U2114 (N_2114,In_1680,In_1184);
nand U2115 (N_2115,In_53,In_1909);
nand U2116 (N_2116,In_1850,In_1355);
nor U2117 (N_2117,In_1403,In_459);
and U2118 (N_2118,In_1131,In_1464);
nand U2119 (N_2119,In_1219,In_1117);
or U2120 (N_2120,In_995,In_603);
nand U2121 (N_2121,In_790,In_1069);
nand U2122 (N_2122,In_1760,In_968);
nand U2123 (N_2123,In_1009,In_1629);
or U2124 (N_2124,In_1357,In_613);
nor U2125 (N_2125,In_476,In_843);
or U2126 (N_2126,In_1231,In_1192);
or U2127 (N_2127,In_272,In_1586);
or U2128 (N_2128,In_1478,In_855);
nand U2129 (N_2129,In_847,In_109);
nor U2130 (N_2130,In_877,In_1857);
or U2131 (N_2131,In_1489,In_744);
xnor U2132 (N_2132,In_993,In_1823);
nor U2133 (N_2133,In_673,In_1769);
or U2134 (N_2134,In_469,In_1728);
nand U2135 (N_2135,In_437,In_1280);
and U2136 (N_2136,In_1112,In_855);
nor U2137 (N_2137,In_1461,In_1988);
and U2138 (N_2138,In_446,In_367);
and U2139 (N_2139,In_197,In_778);
nor U2140 (N_2140,In_1072,In_788);
nand U2141 (N_2141,In_206,In_932);
or U2142 (N_2142,In_1785,In_1770);
and U2143 (N_2143,In_211,In_829);
xor U2144 (N_2144,In_1847,In_365);
or U2145 (N_2145,In_1686,In_513);
nor U2146 (N_2146,In_124,In_1743);
nor U2147 (N_2147,In_1016,In_58);
nand U2148 (N_2148,In_564,In_217);
nor U2149 (N_2149,In_329,In_340);
and U2150 (N_2150,In_810,In_551);
nand U2151 (N_2151,In_174,In_1051);
or U2152 (N_2152,In_1236,In_1633);
or U2153 (N_2153,In_1659,In_787);
or U2154 (N_2154,In_1099,In_643);
nor U2155 (N_2155,In_1568,In_1444);
xnor U2156 (N_2156,In_744,In_193);
or U2157 (N_2157,In_753,In_126);
nor U2158 (N_2158,In_543,In_22);
nand U2159 (N_2159,In_1014,In_337);
nor U2160 (N_2160,In_670,In_1126);
nand U2161 (N_2161,In_1049,In_212);
nor U2162 (N_2162,In_836,In_1027);
nand U2163 (N_2163,In_545,In_1419);
and U2164 (N_2164,In_1938,In_779);
xnor U2165 (N_2165,In_1695,In_788);
and U2166 (N_2166,In_1165,In_1600);
and U2167 (N_2167,In_727,In_523);
or U2168 (N_2168,In_1093,In_1659);
nor U2169 (N_2169,In_1927,In_1918);
or U2170 (N_2170,In_874,In_505);
nand U2171 (N_2171,In_1204,In_142);
xnor U2172 (N_2172,In_1115,In_698);
or U2173 (N_2173,In_1436,In_1584);
or U2174 (N_2174,In_787,In_373);
nor U2175 (N_2175,In_1671,In_605);
or U2176 (N_2176,In_1058,In_982);
nand U2177 (N_2177,In_134,In_102);
nor U2178 (N_2178,In_654,In_665);
and U2179 (N_2179,In_900,In_1024);
nor U2180 (N_2180,In_1474,In_1460);
or U2181 (N_2181,In_1088,In_922);
or U2182 (N_2182,In_534,In_535);
and U2183 (N_2183,In_597,In_921);
nand U2184 (N_2184,In_310,In_1824);
xor U2185 (N_2185,In_1605,In_764);
and U2186 (N_2186,In_972,In_1363);
nand U2187 (N_2187,In_560,In_1835);
and U2188 (N_2188,In_1373,In_1086);
nor U2189 (N_2189,In_182,In_1523);
and U2190 (N_2190,In_1579,In_1261);
or U2191 (N_2191,In_32,In_1842);
or U2192 (N_2192,In_1120,In_169);
and U2193 (N_2193,In_238,In_49);
nor U2194 (N_2194,In_731,In_1881);
nor U2195 (N_2195,In_968,In_1060);
or U2196 (N_2196,In_4,In_1031);
xnor U2197 (N_2197,In_812,In_1334);
nor U2198 (N_2198,In_376,In_192);
and U2199 (N_2199,In_672,In_159);
xnor U2200 (N_2200,In_227,In_804);
and U2201 (N_2201,In_1458,In_1012);
xor U2202 (N_2202,In_1500,In_1966);
nor U2203 (N_2203,In_275,In_1158);
and U2204 (N_2204,In_1052,In_707);
nand U2205 (N_2205,In_447,In_814);
and U2206 (N_2206,In_1841,In_214);
xor U2207 (N_2207,In_1749,In_1285);
and U2208 (N_2208,In_548,In_391);
nand U2209 (N_2209,In_1859,In_765);
or U2210 (N_2210,In_1383,In_1513);
and U2211 (N_2211,In_1155,In_145);
or U2212 (N_2212,In_853,In_1455);
nand U2213 (N_2213,In_205,In_168);
or U2214 (N_2214,In_1974,In_70);
nand U2215 (N_2215,In_280,In_455);
and U2216 (N_2216,In_651,In_1583);
and U2217 (N_2217,In_882,In_1551);
nor U2218 (N_2218,In_148,In_708);
or U2219 (N_2219,In_1710,In_221);
xnor U2220 (N_2220,In_1670,In_1194);
or U2221 (N_2221,In_301,In_1033);
nor U2222 (N_2222,In_1694,In_21);
and U2223 (N_2223,In_1386,In_1461);
nor U2224 (N_2224,In_693,In_130);
or U2225 (N_2225,In_868,In_898);
nand U2226 (N_2226,In_1440,In_472);
nand U2227 (N_2227,In_943,In_776);
or U2228 (N_2228,In_1616,In_531);
and U2229 (N_2229,In_43,In_1619);
and U2230 (N_2230,In_437,In_1105);
nor U2231 (N_2231,In_1769,In_973);
nand U2232 (N_2232,In_1766,In_1237);
or U2233 (N_2233,In_1237,In_1550);
or U2234 (N_2234,In_52,In_110);
nand U2235 (N_2235,In_1452,In_799);
and U2236 (N_2236,In_1865,In_1662);
or U2237 (N_2237,In_784,In_155);
and U2238 (N_2238,In_425,In_1368);
xnor U2239 (N_2239,In_1701,In_895);
and U2240 (N_2240,In_772,In_1304);
nand U2241 (N_2241,In_608,In_30);
nor U2242 (N_2242,In_1644,In_234);
nor U2243 (N_2243,In_1448,In_1617);
xor U2244 (N_2244,In_23,In_1518);
xor U2245 (N_2245,In_1945,In_115);
or U2246 (N_2246,In_1510,In_989);
nand U2247 (N_2247,In_806,In_1265);
nor U2248 (N_2248,In_1520,In_8);
nand U2249 (N_2249,In_1749,In_1955);
xnor U2250 (N_2250,In_1440,In_1556);
nand U2251 (N_2251,In_234,In_679);
or U2252 (N_2252,In_126,In_1758);
and U2253 (N_2253,In_1690,In_652);
xor U2254 (N_2254,In_1600,In_1811);
nand U2255 (N_2255,In_318,In_1779);
nor U2256 (N_2256,In_1609,In_404);
and U2257 (N_2257,In_526,In_318);
or U2258 (N_2258,In_93,In_1638);
and U2259 (N_2259,In_205,In_772);
or U2260 (N_2260,In_924,In_810);
and U2261 (N_2261,In_872,In_161);
or U2262 (N_2262,In_586,In_1404);
and U2263 (N_2263,In_1585,In_1718);
nor U2264 (N_2264,In_351,In_603);
nand U2265 (N_2265,In_1882,In_1499);
and U2266 (N_2266,In_1282,In_310);
nor U2267 (N_2267,In_1219,In_1226);
or U2268 (N_2268,In_993,In_1296);
nor U2269 (N_2269,In_896,In_770);
and U2270 (N_2270,In_186,In_323);
nor U2271 (N_2271,In_1871,In_881);
nor U2272 (N_2272,In_1046,In_1066);
or U2273 (N_2273,In_1874,In_1968);
nand U2274 (N_2274,In_296,In_107);
and U2275 (N_2275,In_643,In_1881);
and U2276 (N_2276,In_1156,In_956);
nor U2277 (N_2277,In_1410,In_845);
or U2278 (N_2278,In_721,In_698);
xnor U2279 (N_2279,In_673,In_748);
or U2280 (N_2280,In_943,In_1555);
or U2281 (N_2281,In_458,In_1181);
and U2282 (N_2282,In_687,In_482);
and U2283 (N_2283,In_268,In_1183);
nor U2284 (N_2284,In_1,In_557);
nor U2285 (N_2285,In_1044,In_619);
nor U2286 (N_2286,In_1303,In_240);
nor U2287 (N_2287,In_1439,In_1647);
and U2288 (N_2288,In_1228,In_403);
and U2289 (N_2289,In_1857,In_896);
xnor U2290 (N_2290,In_1593,In_1324);
or U2291 (N_2291,In_461,In_1699);
and U2292 (N_2292,In_1344,In_1714);
nor U2293 (N_2293,In_1479,In_1395);
or U2294 (N_2294,In_864,In_533);
nor U2295 (N_2295,In_960,In_1498);
or U2296 (N_2296,In_1865,In_717);
or U2297 (N_2297,In_641,In_1607);
xor U2298 (N_2298,In_1206,In_407);
or U2299 (N_2299,In_1601,In_425);
nor U2300 (N_2300,In_1910,In_1597);
and U2301 (N_2301,In_662,In_1954);
and U2302 (N_2302,In_955,In_672);
nor U2303 (N_2303,In_953,In_1852);
and U2304 (N_2304,In_782,In_1407);
and U2305 (N_2305,In_1126,In_659);
nand U2306 (N_2306,In_1392,In_1012);
and U2307 (N_2307,In_1354,In_1255);
nor U2308 (N_2308,In_85,In_1122);
nand U2309 (N_2309,In_1161,In_1031);
nand U2310 (N_2310,In_823,In_1444);
nor U2311 (N_2311,In_29,In_103);
nand U2312 (N_2312,In_200,In_735);
and U2313 (N_2313,In_1692,In_174);
nor U2314 (N_2314,In_837,In_1855);
nor U2315 (N_2315,In_1103,In_630);
nor U2316 (N_2316,In_356,In_928);
nand U2317 (N_2317,In_81,In_1688);
nand U2318 (N_2318,In_733,In_662);
or U2319 (N_2319,In_485,In_1422);
nor U2320 (N_2320,In_333,In_495);
or U2321 (N_2321,In_817,In_1379);
nor U2322 (N_2322,In_1249,In_801);
and U2323 (N_2323,In_663,In_1083);
nand U2324 (N_2324,In_878,In_127);
nor U2325 (N_2325,In_954,In_1260);
nor U2326 (N_2326,In_697,In_753);
nand U2327 (N_2327,In_689,In_842);
nor U2328 (N_2328,In_728,In_1705);
and U2329 (N_2329,In_427,In_1564);
and U2330 (N_2330,In_325,In_991);
nor U2331 (N_2331,In_691,In_65);
or U2332 (N_2332,In_1193,In_1427);
or U2333 (N_2333,In_385,In_1992);
or U2334 (N_2334,In_388,In_344);
xor U2335 (N_2335,In_977,In_1092);
nand U2336 (N_2336,In_1010,In_653);
and U2337 (N_2337,In_1664,In_1229);
nor U2338 (N_2338,In_1936,In_1539);
nor U2339 (N_2339,In_1219,In_1653);
nand U2340 (N_2340,In_1602,In_235);
and U2341 (N_2341,In_693,In_183);
nand U2342 (N_2342,In_1515,In_1365);
and U2343 (N_2343,In_712,In_1535);
and U2344 (N_2344,In_28,In_182);
nor U2345 (N_2345,In_367,In_1074);
and U2346 (N_2346,In_1955,In_1256);
nor U2347 (N_2347,In_284,In_1313);
nand U2348 (N_2348,In_1467,In_1399);
nor U2349 (N_2349,In_315,In_928);
and U2350 (N_2350,In_922,In_858);
and U2351 (N_2351,In_543,In_1976);
nand U2352 (N_2352,In_64,In_1281);
nor U2353 (N_2353,In_1036,In_1479);
and U2354 (N_2354,In_999,In_480);
nand U2355 (N_2355,In_311,In_5);
or U2356 (N_2356,In_1692,In_128);
nand U2357 (N_2357,In_355,In_835);
nor U2358 (N_2358,In_159,In_92);
nand U2359 (N_2359,In_296,In_1360);
or U2360 (N_2360,In_249,In_1189);
nand U2361 (N_2361,In_1632,In_254);
nand U2362 (N_2362,In_1247,In_1979);
and U2363 (N_2363,In_1978,In_268);
nor U2364 (N_2364,In_1674,In_1410);
and U2365 (N_2365,In_65,In_1603);
xor U2366 (N_2366,In_604,In_107);
or U2367 (N_2367,In_492,In_1665);
or U2368 (N_2368,In_1173,In_64);
or U2369 (N_2369,In_1335,In_440);
nor U2370 (N_2370,In_1578,In_1034);
xor U2371 (N_2371,In_44,In_108);
nand U2372 (N_2372,In_279,In_1227);
nand U2373 (N_2373,In_878,In_407);
or U2374 (N_2374,In_534,In_1054);
nor U2375 (N_2375,In_1340,In_1148);
and U2376 (N_2376,In_1676,In_1918);
nor U2377 (N_2377,In_418,In_1541);
and U2378 (N_2378,In_691,In_733);
nand U2379 (N_2379,In_1094,In_247);
or U2380 (N_2380,In_1764,In_1600);
nor U2381 (N_2381,In_1630,In_909);
or U2382 (N_2382,In_158,In_787);
nor U2383 (N_2383,In_1621,In_204);
nand U2384 (N_2384,In_42,In_1098);
nor U2385 (N_2385,In_1310,In_492);
and U2386 (N_2386,In_1418,In_1447);
and U2387 (N_2387,In_1711,In_677);
or U2388 (N_2388,In_1369,In_1320);
nor U2389 (N_2389,In_876,In_698);
and U2390 (N_2390,In_945,In_101);
nand U2391 (N_2391,In_1400,In_1160);
nand U2392 (N_2392,In_522,In_1472);
and U2393 (N_2393,In_135,In_588);
and U2394 (N_2394,In_1366,In_616);
and U2395 (N_2395,In_1867,In_1134);
and U2396 (N_2396,In_1879,In_2);
and U2397 (N_2397,In_22,In_503);
or U2398 (N_2398,In_1436,In_396);
and U2399 (N_2399,In_757,In_888);
or U2400 (N_2400,In_1211,In_1427);
nor U2401 (N_2401,In_846,In_1595);
or U2402 (N_2402,In_1336,In_232);
nor U2403 (N_2403,In_272,In_366);
nor U2404 (N_2404,In_83,In_1287);
or U2405 (N_2405,In_426,In_1066);
nor U2406 (N_2406,In_466,In_1090);
or U2407 (N_2407,In_425,In_1056);
nor U2408 (N_2408,In_118,In_987);
nand U2409 (N_2409,In_158,In_103);
or U2410 (N_2410,In_138,In_671);
or U2411 (N_2411,In_466,In_994);
nand U2412 (N_2412,In_882,In_986);
and U2413 (N_2413,In_1998,In_436);
nor U2414 (N_2414,In_1714,In_592);
and U2415 (N_2415,In_546,In_149);
nor U2416 (N_2416,In_1129,In_252);
or U2417 (N_2417,In_1654,In_1467);
and U2418 (N_2418,In_1462,In_941);
or U2419 (N_2419,In_1316,In_133);
and U2420 (N_2420,In_1112,In_1744);
nor U2421 (N_2421,In_1218,In_951);
nor U2422 (N_2422,In_1175,In_1696);
and U2423 (N_2423,In_1211,In_1057);
nand U2424 (N_2424,In_613,In_1310);
and U2425 (N_2425,In_789,In_1580);
and U2426 (N_2426,In_1175,In_1261);
and U2427 (N_2427,In_1161,In_103);
nor U2428 (N_2428,In_1426,In_976);
and U2429 (N_2429,In_148,In_31);
and U2430 (N_2430,In_1708,In_1091);
nand U2431 (N_2431,In_1437,In_677);
nand U2432 (N_2432,In_154,In_1041);
or U2433 (N_2433,In_1696,In_657);
or U2434 (N_2434,In_1223,In_1244);
or U2435 (N_2435,In_1886,In_1505);
and U2436 (N_2436,In_861,In_347);
or U2437 (N_2437,In_522,In_929);
or U2438 (N_2438,In_61,In_355);
and U2439 (N_2439,In_1634,In_104);
nand U2440 (N_2440,In_775,In_957);
nand U2441 (N_2441,In_929,In_724);
and U2442 (N_2442,In_91,In_1507);
nor U2443 (N_2443,In_104,In_484);
or U2444 (N_2444,In_214,In_925);
nor U2445 (N_2445,In_1608,In_998);
and U2446 (N_2446,In_1786,In_891);
and U2447 (N_2447,In_1846,In_787);
nor U2448 (N_2448,In_1866,In_76);
nor U2449 (N_2449,In_310,In_1523);
and U2450 (N_2450,In_1029,In_1206);
nor U2451 (N_2451,In_1199,In_336);
and U2452 (N_2452,In_1759,In_307);
and U2453 (N_2453,In_1928,In_1933);
or U2454 (N_2454,In_1442,In_653);
nand U2455 (N_2455,In_480,In_574);
nor U2456 (N_2456,In_1110,In_585);
nand U2457 (N_2457,In_199,In_1633);
or U2458 (N_2458,In_1736,In_1721);
nand U2459 (N_2459,In_1929,In_1430);
and U2460 (N_2460,In_89,In_545);
and U2461 (N_2461,In_267,In_416);
and U2462 (N_2462,In_91,In_300);
or U2463 (N_2463,In_1298,In_1525);
and U2464 (N_2464,In_1997,In_784);
or U2465 (N_2465,In_779,In_90);
and U2466 (N_2466,In_325,In_1187);
and U2467 (N_2467,In_399,In_1947);
and U2468 (N_2468,In_3,In_1181);
nand U2469 (N_2469,In_1244,In_673);
or U2470 (N_2470,In_1909,In_1531);
nor U2471 (N_2471,In_866,In_715);
nor U2472 (N_2472,In_30,In_1233);
nor U2473 (N_2473,In_1157,In_1378);
and U2474 (N_2474,In_1253,In_1976);
nand U2475 (N_2475,In_559,In_1821);
nor U2476 (N_2476,In_776,In_1263);
nor U2477 (N_2477,In_1551,In_875);
and U2478 (N_2478,In_1748,In_1893);
or U2479 (N_2479,In_1866,In_165);
nand U2480 (N_2480,In_271,In_360);
nor U2481 (N_2481,In_997,In_1063);
or U2482 (N_2482,In_1776,In_973);
nor U2483 (N_2483,In_254,In_1286);
and U2484 (N_2484,In_1434,In_1572);
nand U2485 (N_2485,In_702,In_1587);
nand U2486 (N_2486,In_617,In_952);
nand U2487 (N_2487,In_622,In_66);
nor U2488 (N_2488,In_1329,In_882);
nor U2489 (N_2489,In_954,In_1149);
nand U2490 (N_2490,In_1827,In_947);
and U2491 (N_2491,In_1618,In_1301);
and U2492 (N_2492,In_1639,In_1544);
or U2493 (N_2493,In_317,In_1510);
nor U2494 (N_2494,In_307,In_512);
or U2495 (N_2495,In_1049,In_906);
nand U2496 (N_2496,In_265,In_673);
nand U2497 (N_2497,In_1810,In_1218);
or U2498 (N_2498,In_949,In_1430);
nand U2499 (N_2499,In_1276,In_1896);
nor U2500 (N_2500,In_1881,In_113);
nand U2501 (N_2501,In_1313,In_1012);
and U2502 (N_2502,In_481,In_484);
xor U2503 (N_2503,In_1708,In_1363);
nand U2504 (N_2504,In_1014,In_576);
and U2505 (N_2505,In_958,In_88);
or U2506 (N_2506,In_950,In_1878);
nand U2507 (N_2507,In_922,In_1199);
nand U2508 (N_2508,In_226,In_396);
and U2509 (N_2509,In_1590,In_1492);
nand U2510 (N_2510,In_494,In_153);
and U2511 (N_2511,In_650,In_1447);
and U2512 (N_2512,In_614,In_8);
and U2513 (N_2513,In_88,In_1136);
or U2514 (N_2514,In_1088,In_886);
nand U2515 (N_2515,In_764,In_264);
or U2516 (N_2516,In_573,In_100);
nand U2517 (N_2517,In_844,In_1628);
nand U2518 (N_2518,In_673,In_1081);
or U2519 (N_2519,In_1962,In_330);
or U2520 (N_2520,In_1375,In_485);
and U2521 (N_2521,In_473,In_1657);
or U2522 (N_2522,In_1153,In_1179);
nand U2523 (N_2523,In_1740,In_1598);
or U2524 (N_2524,In_501,In_1820);
or U2525 (N_2525,In_266,In_298);
and U2526 (N_2526,In_1590,In_1564);
nor U2527 (N_2527,In_926,In_1981);
nor U2528 (N_2528,In_1792,In_1262);
or U2529 (N_2529,In_1987,In_1284);
xnor U2530 (N_2530,In_1022,In_387);
and U2531 (N_2531,In_1199,In_1475);
or U2532 (N_2532,In_1320,In_1414);
or U2533 (N_2533,In_68,In_1755);
and U2534 (N_2534,In_1164,In_1876);
or U2535 (N_2535,In_370,In_1744);
or U2536 (N_2536,In_743,In_1791);
nor U2537 (N_2537,In_447,In_24);
and U2538 (N_2538,In_524,In_309);
or U2539 (N_2539,In_63,In_1891);
nand U2540 (N_2540,In_162,In_373);
nand U2541 (N_2541,In_494,In_297);
or U2542 (N_2542,In_791,In_1922);
nor U2543 (N_2543,In_902,In_1618);
and U2544 (N_2544,In_559,In_897);
nand U2545 (N_2545,In_1348,In_216);
nand U2546 (N_2546,In_542,In_1659);
or U2547 (N_2547,In_451,In_1826);
and U2548 (N_2548,In_1908,In_1799);
nand U2549 (N_2549,In_1186,In_1364);
and U2550 (N_2550,In_1562,In_604);
nor U2551 (N_2551,In_490,In_1346);
nand U2552 (N_2552,In_896,In_150);
nor U2553 (N_2553,In_1890,In_471);
or U2554 (N_2554,In_451,In_1059);
nand U2555 (N_2555,In_1000,In_1139);
nor U2556 (N_2556,In_975,In_1403);
nor U2557 (N_2557,In_1958,In_1966);
and U2558 (N_2558,In_181,In_1695);
nand U2559 (N_2559,In_1602,In_1632);
nand U2560 (N_2560,In_1505,In_1594);
and U2561 (N_2561,In_323,In_322);
nand U2562 (N_2562,In_78,In_1283);
nand U2563 (N_2563,In_186,In_80);
or U2564 (N_2564,In_1101,In_379);
nor U2565 (N_2565,In_1885,In_1512);
nor U2566 (N_2566,In_533,In_1166);
nor U2567 (N_2567,In_1947,In_1857);
or U2568 (N_2568,In_1033,In_1752);
nand U2569 (N_2569,In_120,In_1027);
or U2570 (N_2570,In_1471,In_124);
nand U2571 (N_2571,In_583,In_1599);
and U2572 (N_2572,In_1433,In_1267);
nand U2573 (N_2573,In_1373,In_1461);
nand U2574 (N_2574,In_1411,In_193);
and U2575 (N_2575,In_648,In_387);
and U2576 (N_2576,In_1137,In_450);
and U2577 (N_2577,In_948,In_601);
nand U2578 (N_2578,In_1346,In_1304);
nor U2579 (N_2579,In_815,In_723);
nor U2580 (N_2580,In_1905,In_786);
and U2581 (N_2581,In_89,In_790);
nand U2582 (N_2582,In_264,In_947);
nor U2583 (N_2583,In_1991,In_516);
nand U2584 (N_2584,In_1617,In_1783);
nor U2585 (N_2585,In_1283,In_1923);
and U2586 (N_2586,In_1476,In_985);
nand U2587 (N_2587,In_293,In_209);
nor U2588 (N_2588,In_1319,In_559);
nand U2589 (N_2589,In_1229,In_720);
and U2590 (N_2590,In_967,In_772);
nand U2591 (N_2591,In_228,In_1069);
and U2592 (N_2592,In_410,In_155);
and U2593 (N_2593,In_1330,In_357);
nand U2594 (N_2594,In_545,In_1211);
or U2595 (N_2595,In_1046,In_1561);
or U2596 (N_2596,In_696,In_217);
and U2597 (N_2597,In_803,In_145);
nand U2598 (N_2598,In_669,In_672);
and U2599 (N_2599,In_1915,In_179);
xnor U2600 (N_2600,In_1622,In_1312);
or U2601 (N_2601,In_1043,In_374);
nor U2602 (N_2602,In_1930,In_1355);
or U2603 (N_2603,In_1068,In_1045);
and U2604 (N_2604,In_948,In_6);
and U2605 (N_2605,In_957,In_1979);
and U2606 (N_2606,In_1422,In_959);
nand U2607 (N_2607,In_78,In_130);
and U2608 (N_2608,In_323,In_845);
or U2609 (N_2609,In_1068,In_594);
or U2610 (N_2610,In_11,In_1043);
nand U2611 (N_2611,In_1550,In_1961);
or U2612 (N_2612,In_1679,In_1046);
or U2613 (N_2613,In_125,In_1354);
or U2614 (N_2614,In_1631,In_1305);
nor U2615 (N_2615,In_735,In_539);
and U2616 (N_2616,In_1751,In_1775);
or U2617 (N_2617,In_3,In_1068);
nand U2618 (N_2618,In_159,In_1818);
and U2619 (N_2619,In_1887,In_1069);
or U2620 (N_2620,In_1493,In_1914);
and U2621 (N_2621,In_161,In_1587);
and U2622 (N_2622,In_23,In_1293);
or U2623 (N_2623,In_514,In_57);
nand U2624 (N_2624,In_127,In_1510);
and U2625 (N_2625,In_1267,In_1044);
nor U2626 (N_2626,In_1379,In_1200);
and U2627 (N_2627,In_1011,In_809);
nor U2628 (N_2628,In_559,In_1364);
nor U2629 (N_2629,In_917,In_1756);
nand U2630 (N_2630,In_1299,In_994);
and U2631 (N_2631,In_1759,In_1429);
nand U2632 (N_2632,In_614,In_183);
or U2633 (N_2633,In_1438,In_631);
nor U2634 (N_2634,In_1747,In_1513);
xnor U2635 (N_2635,In_334,In_1395);
nor U2636 (N_2636,In_300,In_1086);
or U2637 (N_2637,In_399,In_1990);
nand U2638 (N_2638,In_1323,In_1806);
nor U2639 (N_2639,In_127,In_1656);
nand U2640 (N_2640,In_605,In_1102);
nor U2641 (N_2641,In_1905,In_1961);
and U2642 (N_2642,In_1074,In_1830);
and U2643 (N_2643,In_798,In_1480);
and U2644 (N_2644,In_120,In_1321);
and U2645 (N_2645,In_121,In_793);
and U2646 (N_2646,In_1833,In_894);
nor U2647 (N_2647,In_1639,In_416);
and U2648 (N_2648,In_1721,In_831);
or U2649 (N_2649,In_528,In_1901);
nand U2650 (N_2650,In_1991,In_426);
and U2651 (N_2651,In_599,In_1748);
nor U2652 (N_2652,In_121,In_670);
or U2653 (N_2653,In_870,In_996);
nand U2654 (N_2654,In_299,In_1898);
or U2655 (N_2655,In_950,In_1737);
or U2656 (N_2656,In_1382,In_1328);
nor U2657 (N_2657,In_969,In_185);
nand U2658 (N_2658,In_822,In_691);
nand U2659 (N_2659,In_1188,In_25);
or U2660 (N_2660,In_1874,In_1461);
nor U2661 (N_2661,In_1264,In_1762);
nand U2662 (N_2662,In_1039,In_1475);
nor U2663 (N_2663,In_248,In_757);
nand U2664 (N_2664,In_12,In_683);
nand U2665 (N_2665,In_1521,In_1696);
or U2666 (N_2666,In_1135,In_89);
nand U2667 (N_2667,In_1502,In_77);
nor U2668 (N_2668,In_1614,In_352);
nor U2669 (N_2669,In_939,In_1472);
and U2670 (N_2670,In_392,In_1496);
nor U2671 (N_2671,In_1843,In_1616);
nor U2672 (N_2672,In_1379,In_1869);
or U2673 (N_2673,In_1467,In_554);
and U2674 (N_2674,In_530,In_160);
nand U2675 (N_2675,In_599,In_1435);
nand U2676 (N_2676,In_1148,In_1721);
nand U2677 (N_2677,In_508,In_631);
and U2678 (N_2678,In_870,In_1591);
nor U2679 (N_2679,In_48,In_1801);
and U2680 (N_2680,In_1436,In_1056);
and U2681 (N_2681,In_80,In_1367);
and U2682 (N_2682,In_1932,In_1790);
nand U2683 (N_2683,In_278,In_972);
nor U2684 (N_2684,In_808,In_627);
nor U2685 (N_2685,In_1715,In_912);
and U2686 (N_2686,In_1788,In_267);
nor U2687 (N_2687,In_1133,In_372);
nor U2688 (N_2688,In_492,In_939);
xor U2689 (N_2689,In_60,In_109);
nor U2690 (N_2690,In_1064,In_320);
nand U2691 (N_2691,In_151,In_306);
xnor U2692 (N_2692,In_702,In_1202);
nand U2693 (N_2693,In_729,In_1343);
or U2694 (N_2694,In_1382,In_287);
nor U2695 (N_2695,In_1541,In_684);
nor U2696 (N_2696,In_529,In_1077);
nand U2697 (N_2697,In_1559,In_757);
and U2698 (N_2698,In_1724,In_1786);
nand U2699 (N_2699,In_339,In_1939);
nor U2700 (N_2700,In_881,In_666);
nor U2701 (N_2701,In_1619,In_139);
nand U2702 (N_2702,In_578,In_1705);
nand U2703 (N_2703,In_1273,In_290);
and U2704 (N_2704,In_1678,In_668);
nand U2705 (N_2705,In_1985,In_120);
and U2706 (N_2706,In_170,In_932);
nand U2707 (N_2707,In_1032,In_276);
and U2708 (N_2708,In_622,In_304);
nor U2709 (N_2709,In_61,In_1809);
nand U2710 (N_2710,In_1041,In_457);
and U2711 (N_2711,In_1894,In_462);
or U2712 (N_2712,In_901,In_1217);
nor U2713 (N_2713,In_1829,In_658);
or U2714 (N_2714,In_923,In_233);
and U2715 (N_2715,In_198,In_1357);
nand U2716 (N_2716,In_1914,In_1205);
nor U2717 (N_2717,In_877,In_23);
or U2718 (N_2718,In_1230,In_842);
nor U2719 (N_2719,In_1435,In_704);
and U2720 (N_2720,In_1923,In_1052);
or U2721 (N_2721,In_813,In_1848);
and U2722 (N_2722,In_1049,In_1047);
and U2723 (N_2723,In_1846,In_622);
nand U2724 (N_2724,In_1398,In_1122);
nor U2725 (N_2725,In_690,In_19);
nand U2726 (N_2726,In_1683,In_748);
or U2727 (N_2727,In_658,In_611);
and U2728 (N_2728,In_1885,In_1614);
nand U2729 (N_2729,In_1213,In_252);
or U2730 (N_2730,In_1397,In_569);
nand U2731 (N_2731,In_806,In_1315);
xor U2732 (N_2732,In_524,In_1397);
nor U2733 (N_2733,In_374,In_238);
nand U2734 (N_2734,In_1165,In_914);
or U2735 (N_2735,In_276,In_656);
and U2736 (N_2736,In_938,In_483);
nand U2737 (N_2737,In_1606,In_1009);
xor U2738 (N_2738,In_236,In_0);
and U2739 (N_2739,In_1373,In_962);
and U2740 (N_2740,In_802,In_56);
and U2741 (N_2741,In_1403,In_1193);
nand U2742 (N_2742,In_1691,In_2);
nor U2743 (N_2743,In_101,In_81);
nor U2744 (N_2744,In_1964,In_159);
nor U2745 (N_2745,In_1574,In_356);
nor U2746 (N_2746,In_1941,In_1786);
and U2747 (N_2747,In_1072,In_966);
nand U2748 (N_2748,In_1666,In_1814);
and U2749 (N_2749,In_1538,In_99);
or U2750 (N_2750,In_1570,In_1111);
or U2751 (N_2751,In_21,In_671);
or U2752 (N_2752,In_1204,In_1933);
and U2753 (N_2753,In_1530,In_377);
or U2754 (N_2754,In_903,In_1964);
or U2755 (N_2755,In_717,In_507);
nor U2756 (N_2756,In_859,In_197);
nor U2757 (N_2757,In_168,In_248);
nand U2758 (N_2758,In_89,In_353);
nand U2759 (N_2759,In_1180,In_1688);
xor U2760 (N_2760,In_1382,In_1684);
and U2761 (N_2761,In_1887,In_149);
nand U2762 (N_2762,In_1367,In_1987);
nor U2763 (N_2763,In_1970,In_1999);
and U2764 (N_2764,In_500,In_327);
xnor U2765 (N_2765,In_1751,In_784);
nor U2766 (N_2766,In_569,In_924);
or U2767 (N_2767,In_1496,In_1615);
nand U2768 (N_2768,In_187,In_1628);
and U2769 (N_2769,In_351,In_1154);
or U2770 (N_2770,In_309,In_1420);
and U2771 (N_2771,In_1759,In_324);
or U2772 (N_2772,In_1524,In_1838);
nand U2773 (N_2773,In_472,In_1625);
or U2774 (N_2774,In_1959,In_1996);
nand U2775 (N_2775,In_1942,In_455);
nand U2776 (N_2776,In_1560,In_1646);
and U2777 (N_2777,In_408,In_1090);
or U2778 (N_2778,In_257,In_1283);
nand U2779 (N_2779,In_352,In_923);
nor U2780 (N_2780,In_914,In_1197);
and U2781 (N_2781,In_964,In_84);
or U2782 (N_2782,In_932,In_1043);
nand U2783 (N_2783,In_1030,In_458);
and U2784 (N_2784,In_657,In_908);
nor U2785 (N_2785,In_1789,In_925);
nand U2786 (N_2786,In_1476,In_1516);
and U2787 (N_2787,In_1537,In_756);
nand U2788 (N_2788,In_237,In_741);
and U2789 (N_2789,In_1259,In_1254);
nor U2790 (N_2790,In_1390,In_1142);
or U2791 (N_2791,In_1287,In_1320);
nor U2792 (N_2792,In_1194,In_782);
nand U2793 (N_2793,In_717,In_1232);
nor U2794 (N_2794,In_607,In_400);
nand U2795 (N_2795,In_1335,In_1382);
nand U2796 (N_2796,In_1322,In_1525);
nand U2797 (N_2797,In_63,In_191);
nor U2798 (N_2798,In_1097,In_1255);
or U2799 (N_2799,In_1384,In_1817);
or U2800 (N_2800,In_537,In_1983);
nand U2801 (N_2801,In_707,In_1490);
or U2802 (N_2802,In_206,In_1859);
nand U2803 (N_2803,In_1,In_358);
nand U2804 (N_2804,In_96,In_1079);
or U2805 (N_2805,In_1731,In_1825);
nor U2806 (N_2806,In_959,In_24);
nor U2807 (N_2807,In_969,In_1454);
and U2808 (N_2808,In_1353,In_833);
and U2809 (N_2809,In_454,In_687);
nand U2810 (N_2810,In_558,In_1139);
and U2811 (N_2811,In_1251,In_327);
or U2812 (N_2812,In_1437,In_524);
and U2813 (N_2813,In_370,In_1470);
or U2814 (N_2814,In_1195,In_695);
nand U2815 (N_2815,In_1266,In_1770);
nor U2816 (N_2816,In_1016,In_1286);
nor U2817 (N_2817,In_491,In_1687);
nor U2818 (N_2818,In_1657,In_745);
nand U2819 (N_2819,In_1267,In_944);
or U2820 (N_2820,In_957,In_784);
and U2821 (N_2821,In_715,In_1451);
nand U2822 (N_2822,In_761,In_1227);
nand U2823 (N_2823,In_211,In_321);
nand U2824 (N_2824,In_654,In_255);
and U2825 (N_2825,In_915,In_992);
or U2826 (N_2826,In_1664,In_748);
nor U2827 (N_2827,In_916,In_264);
and U2828 (N_2828,In_754,In_95);
or U2829 (N_2829,In_1731,In_1755);
nor U2830 (N_2830,In_284,In_621);
or U2831 (N_2831,In_520,In_64);
and U2832 (N_2832,In_553,In_127);
nand U2833 (N_2833,In_1692,In_753);
nand U2834 (N_2834,In_1824,In_1073);
nor U2835 (N_2835,In_813,In_1584);
nand U2836 (N_2836,In_1936,In_1589);
nand U2837 (N_2837,In_1345,In_1520);
or U2838 (N_2838,In_1788,In_1781);
nand U2839 (N_2839,In_983,In_827);
nor U2840 (N_2840,In_1221,In_780);
or U2841 (N_2841,In_154,In_1803);
and U2842 (N_2842,In_169,In_1240);
and U2843 (N_2843,In_1307,In_1824);
or U2844 (N_2844,In_748,In_837);
and U2845 (N_2845,In_770,In_1887);
or U2846 (N_2846,In_147,In_1067);
nor U2847 (N_2847,In_793,In_640);
nor U2848 (N_2848,In_1417,In_1861);
nor U2849 (N_2849,In_211,In_764);
or U2850 (N_2850,In_413,In_1267);
nand U2851 (N_2851,In_831,In_164);
nand U2852 (N_2852,In_1289,In_420);
nand U2853 (N_2853,In_1959,In_1942);
or U2854 (N_2854,In_1585,In_537);
and U2855 (N_2855,In_1078,In_131);
or U2856 (N_2856,In_1208,In_1568);
nand U2857 (N_2857,In_1409,In_1216);
nor U2858 (N_2858,In_721,In_525);
and U2859 (N_2859,In_1341,In_1337);
nand U2860 (N_2860,In_1222,In_1134);
nor U2861 (N_2861,In_388,In_1976);
nand U2862 (N_2862,In_1383,In_773);
nor U2863 (N_2863,In_865,In_42);
nand U2864 (N_2864,In_966,In_1268);
and U2865 (N_2865,In_505,In_913);
and U2866 (N_2866,In_368,In_401);
xnor U2867 (N_2867,In_1831,In_322);
and U2868 (N_2868,In_365,In_1790);
nand U2869 (N_2869,In_6,In_793);
or U2870 (N_2870,In_311,In_1510);
and U2871 (N_2871,In_1712,In_1066);
and U2872 (N_2872,In_1751,In_298);
nand U2873 (N_2873,In_1250,In_1208);
and U2874 (N_2874,In_1583,In_1230);
nand U2875 (N_2875,In_567,In_552);
and U2876 (N_2876,In_146,In_1892);
or U2877 (N_2877,In_1845,In_227);
and U2878 (N_2878,In_1506,In_661);
nor U2879 (N_2879,In_780,In_127);
nand U2880 (N_2880,In_376,In_739);
and U2881 (N_2881,In_418,In_1554);
and U2882 (N_2882,In_305,In_648);
nand U2883 (N_2883,In_1633,In_811);
or U2884 (N_2884,In_466,In_495);
or U2885 (N_2885,In_1147,In_1459);
nand U2886 (N_2886,In_1300,In_1072);
nand U2887 (N_2887,In_1477,In_336);
or U2888 (N_2888,In_1889,In_1960);
or U2889 (N_2889,In_1835,In_1221);
nand U2890 (N_2890,In_1944,In_1233);
and U2891 (N_2891,In_1452,In_1161);
and U2892 (N_2892,In_142,In_1384);
or U2893 (N_2893,In_1586,In_1084);
and U2894 (N_2894,In_824,In_12);
or U2895 (N_2895,In_1959,In_1212);
nor U2896 (N_2896,In_217,In_1447);
and U2897 (N_2897,In_847,In_1869);
nor U2898 (N_2898,In_634,In_982);
and U2899 (N_2899,In_1426,In_1986);
or U2900 (N_2900,In_140,In_1280);
and U2901 (N_2901,In_242,In_79);
nand U2902 (N_2902,In_369,In_1100);
nand U2903 (N_2903,In_192,In_1638);
nor U2904 (N_2904,In_1992,In_862);
nor U2905 (N_2905,In_1759,In_1727);
and U2906 (N_2906,In_554,In_528);
or U2907 (N_2907,In_1140,In_733);
nand U2908 (N_2908,In_299,In_1654);
nor U2909 (N_2909,In_894,In_702);
or U2910 (N_2910,In_102,In_1888);
or U2911 (N_2911,In_1620,In_1107);
and U2912 (N_2912,In_922,In_1352);
nor U2913 (N_2913,In_572,In_1437);
nor U2914 (N_2914,In_126,In_391);
nor U2915 (N_2915,In_1994,In_1336);
nand U2916 (N_2916,In_602,In_1905);
and U2917 (N_2917,In_1854,In_1340);
nor U2918 (N_2918,In_1252,In_394);
nand U2919 (N_2919,In_1687,In_350);
nand U2920 (N_2920,In_1080,In_1190);
or U2921 (N_2921,In_1910,In_1804);
and U2922 (N_2922,In_1805,In_933);
or U2923 (N_2923,In_1615,In_1678);
nand U2924 (N_2924,In_447,In_404);
and U2925 (N_2925,In_475,In_1543);
nor U2926 (N_2926,In_1370,In_331);
or U2927 (N_2927,In_659,In_1705);
and U2928 (N_2928,In_487,In_879);
or U2929 (N_2929,In_373,In_1004);
nand U2930 (N_2930,In_1847,In_166);
nor U2931 (N_2931,In_1785,In_1259);
nor U2932 (N_2932,In_1727,In_1865);
and U2933 (N_2933,In_1850,In_567);
or U2934 (N_2934,In_1180,In_1915);
xnor U2935 (N_2935,In_1322,In_928);
nand U2936 (N_2936,In_512,In_1174);
or U2937 (N_2937,In_1173,In_1785);
and U2938 (N_2938,In_954,In_1835);
xnor U2939 (N_2939,In_1493,In_361);
and U2940 (N_2940,In_287,In_767);
or U2941 (N_2941,In_1532,In_975);
nand U2942 (N_2942,In_34,In_532);
nand U2943 (N_2943,In_287,In_1287);
or U2944 (N_2944,In_1778,In_1548);
nor U2945 (N_2945,In_1641,In_263);
and U2946 (N_2946,In_1126,In_331);
nand U2947 (N_2947,In_1181,In_1660);
and U2948 (N_2948,In_1667,In_1591);
and U2949 (N_2949,In_1924,In_1632);
and U2950 (N_2950,In_291,In_1547);
or U2951 (N_2951,In_99,In_1719);
or U2952 (N_2952,In_1228,In_908);
nand U2953 (N_2953,In_556,In_239);
or U2954 (N_2954,In_1597,In_1125);
nor U2955 (N_2955,In_1120,In_373);
nor U2956 (N_2956,In_1016,In_615);
and U2957 (N_2957,In_1115,In_996);
and U2958 (N_2958,In_1625,In_738);
or U2959 (N_2959,In_228,In_1144);
nor U2960 (N_2960,In_1234,In_1071);
xor U2961 (N_2961,In_378,In_762);
or U2962 (N_2962,In_1575,In_650);
nand U2963 (N_2963,In_1471,In_1028);
nand U2964 (N_2964,In_763,In_120);
or U2965 (N_2965,In_646,In_927);
and U2966 (N_2966,In_1710,In_854);
nand U2967 (N_2967,In_631,In_75);
nor U2968 (N_2968,In_436,In_1004);
nand U2969 (N_2969,In_1461,In_1029);
and U2970 (N_2970,In_201,In_1511);
or U2971 (N_2971,In_1480,In_194);
nand U2972 (N_2972,In_1361,In_871);
nand U2973 (N_2973,In_1800,In_113);
and U2974 (N_2974,In_494,In_1824);
and U2975 (N_2975,In_435,In_1038);
or U2976 (N_2976,In_1610,In_318);
nand U2977 (N_2977,In_235,In_118);
or U2978 (N_2978,In_1566,In_555);
and U2979 (N_2979,In_138,In_1537);
nand U2980 (N_2980,In_1460,In_937);
and U2981 (N_2981,In_577,In_1351);
and U2982 (N_2982,In_86,In_1094);
and U2983 (N_2983,In_1535,In_1010);
and U2984 (N_2984,In_1278,In_1823);
and U2985 (N_2985,In_1931,In_56);
and U2986 (N_2986,In_1803,In_1666);
or U2987 (N_2987,In_1318,In_536);
and U2988 (N_2988,In_1296,In_1505);
nand U2989 (N_2989,In_316,In_1509);
and U2990 (N_2990,In_688,In_1533);
nor U2991 (N_2991,In_1407,In_284);
and U2992 (N_2992,In_391,In_1500);
nand U2993 (N_2993,In_1613,In_760);
nand U2994 (N_2994,In_1342,In_1504);
nor U2995 (N_2995,In_1990,In_1181);
and U2996 (N_2996,In_1311,In_1421);
or U2997 (N_2997,In_1239,In_1924);
and U2998 (N_2998,In_1202,In_583);
nand U2999 (N_2999,In_1853,In_882);
or U3000 (N_3000,In_1536,In_1124);
nor U3001 (N_3001,In_1915,In_1597);
nand U3002 (N_3002,In_1713,In_744);
and U3003 (N_3003,In_55,In_1273);
nand U3004 (N_3004,In_1141,In_1319);
and U3005 (N_3005,In_506,In_1585);
nand U3006 (N_3006,In_497,In_1187);
nand U3007 (N_3007,In_1553,In_1734);
and U3008 (N_3008,In_1066,In_721);
nor U3009 (N_3009,In_1277,In_578);
or U3010 (N_3010,In_221,In_1722);
nand U3011 (N_3011,In_655,In_1896);
nor U3012 (N_3012,In_1527,In_1468);
nand U3013 (N_3013,In_892,In_1683);
nand U3014 (N_3014,In_224,In_862);
xor U3015 (N_3015,In_1830,In_1453);
nor U3016 (N_3016,In_1091,In_1185);
nor U3017 (N_3017,In_1401,In_1275);
nand U3018 (N_3018,In_1283,In_183);
nor U3019 (N_3019,In_1215,In_1235);
nor U3020 (N_3020,In_1913,In_1173);
xnor U3021 (N_3021,In_281,In_40);
and U3022 (N_3022,In_1155,In_1725);
or U3023 (N_3023,In_265,In_9);
and U3024 (N_3024,In_540,In_1543);
or U3025 (N_3025,In_1039,In_1424);
nand U3026 (N_3026,In_1157,In_41);
or U3027 (N_3027,In_645,In_1733);
or U3028 (N_3028,In_1194,In_889);
or U3029 (N_3029,In_1660,In_476);
and U3030 (N_3030,In_1668,In_207);
nand U3031 (N_3031,In_453,In_1559);
or U3032 (N_3032,In_681,In_1702);
or U3033 (N_3033,In_1631,In_1976);
and U3034 (N_3034,In_303,In_1381);
xor U3035 (N_3035,In_1651,In_43);
and U3036 (N_3036,In_771,In_1993);
nand U3037 (N_3037,In_1350,In_1219);
xor U3038 (N_3038,In_889,In_493);
xnor U3039 (N_3039,In_1234,In_1842);
nand U3040 (N_3040,In_1782,In_1594);
nand U3041 (N_3041,In_244,In_762);
or U3042 (N_3042,In_1966,In_134);
or U3043 (N_3043,In_1535,In_978);
or U3044 (N_3044,In_1045,In_1427);
nor U3045 (N_3045,In_1467,In_1626);
nor U3046 (N_3046,In_393,In_734);
nor U3047 (N_3047,In_253,In_950);
or U3048 (N_3048,In_1941,In_447);
and U3049 (N_3049,In_1396,In_575);
and U3050 (N_3050,In_107,In_264);
nand U3051 (N_3051,In_41,In_622);
or U3052 (N_3052,In_1608,In_744);
and U3053 (N_3053,In_1304,In_687);
nor U3054 (N_3054,In_222,In_785);
nand U3055 (N_3055,In_169,In_1573);
xnor U3056 (N_3056,In_113,In_1722);
and U3057 (N_3057,In_125,In_1013);
nand U3058 (N_3058,In_745,In_90);
nor U3059 (N_3059,In_371,In_224);
nand U3060 (N_3060,In_645,In_438);
nand U3061 (N_3061,In_162,In_556);
nor U3062 (N_3062,In_1490,In_148);
and U3063 (N_3063,In_1710,In_1112);
nor U3064 (N_3064,In_689,In_165);
and U3065 (N_3065,In_461,In_379);
or U3066 (N_3066,In_1946,In_146);
and U3067 (N_3067,In_394,In_911);
nor U3068 (N_3068,In_642,In_449);
and U3069 (N_3069,In_174,In_423);
nor U3070 (N_3070,In_1339,In_163);
nand U3071 (N_3071,In_1950,In_1332);
nor U3072 (N_3072,In_329,In_1580);
and U3073 (N_3073,In_171,In_496);
nand U3074 (N_3074,In_1831,In_686);
or U3075 (N_3075,In_749,In_944);
or U3076 (N_3076,In_1202,In_1281);
nand U3077 (N_3077,In_1206,In_1420);
and U3078 (N_3078,In_1192,In_1362);
nor U3079 (N_3079,In_1195,In_1207);
nor U3080 (N_3080,In_895,In_147);
nand U3081 (N_3081,In_1897,In_627);
and U3082 (N_3082,In_1011,In_1164);
nor U3083 (N_3083,In_1188,In_699);
nand U3084 (N_3084,In_301,In_1605);
nor U3085 (N_3085,In_3,In_1725);
or U3086 (N_3086,In_1636,In_1782);
xnor U3087 (N_3087,In_1309,In_946);
nor U3088 (N_3088,In_1781,In_1196);
or U3089 (N_3089,In_1411,In_349);
nand U3090 (N_3090,In_113,In_984);
or U3091 (N_3091,In_669,In_826);
and U3092 (N_3092,In_1273,In_252);
nand U3093 (N_3093,In_490,In_502);
or U3094 (N_3094,In_353,In_1221);
nand U3095 (N_3095,In_680,In_91);
or U3096 (N_3096,In_1770,In_1278);
nand U3097 (N_3097,In_1029,In_226);
or U3098 (N_3098,In_396,In_1049);
or U3099 (N_3099,In_851,In_620);
nor U3100 (N_3100,In_195,In_969);
nor U3101 (N_3101,In_1123,In_919);
and U3102 (N_3102,In_187,In_1305);
nand U3103 (N_3103,In_786,In_233);
nor U3104 (N_3104,In_1847,In_1987);
nand U3105 (N_3105,In_1635,In_1079);
and U3106 (N_3106,In_1019,In_644);
nand U3107 (N_3107,In_992,In_1763);
nand U3108 (N_3108,In_1129,In_1081);
and U3109 (N_3109,In_718,In_619);
or U3110 (N_3110,In_1294,In_333);
or U3111 (N_3111,In_995,In_297);
and U3112 (N_3112,In_504,In_1134);
nor U3113 (N_3113,In_1000,In_1114);
xor U3114 (N_3114,In_409,In_1584);
nand U3115 (N_3115,In_489,In_517);
and U3116 (N_3116,In_1980,In_1520);
and U3117 (N_3117,In_16,In_1327);
and U3118 (N_3118,In_1007,In_1641);
nand U3119 (N_3119,In_25,In_951);
and U3120 (N_3120,In_1849,In_363);
and U3121 (N_3121,In_440,In_651);
nor U3122 (N_3122,In_1954,In_1154);
nor U3123 (N_3123,In_279,In_641);
nor U3124 (N_3124,In_680,In_24);
nor U3125 (N_3125,In_109,In_1745);
nand U3126 (N_3126,In_90,In_1374);
nand U3127 (N_3127,In_1091,In_1656);
nor U3128 (N_3128,In_1365,In_597);
and U3129 (N_3129,In_251,In_335);
and U3130 (N_3130,In_751,In_236);
nor U3131 (N_3131,In_1608,In_734);
or U3132 (N_3132,In_417,In_1623);
and U3133 (N_3133,In_115,In_411);
and U3134 (N_3134,In_141,In_406);
and U3135 (N_3135,In_1475,In_1643);
or U3136 (N_3136,In_552,In_1109);
nand U3137 (N_3137,In_1863,In_1792);
or U3138 (N_3138,In_1277,In_1534);
or U3139 (N_3139,In_670,In_1613);
and U3140 (N_3140,In_703,In_1531);
nor U3141 (N_3141,In_261,In_194);
and U3142 (N_3142,In_1692,In_125);
nor U3143 (N_3143,In_498,In_905);
nor U3144 (N_3144,In_42,In_848);
nand U3145 (N_3145,In_653,In_1663);
nor U3146 (N_3146,In_1213,In_1164);
nand U3147 (N_3147,In_830,In_492);
or U3148 (N_3148,In_1151,In_1059);
nor U3149 (N_3149,In_432,In_747);
nand U3150 (N_3150,In_372,In_589);
nand U3151 (N_3151,In_1322,In_1958);
and U3152 (N_3152,In_1846,In_326);
or U3153 (N_3153,In_464,In_83);
or U3154 (N_3154,In_1614,In_1981);
nand U3155 (N_3155,In_1907,In_1628);
or U3156 (N_3156,In_264,In_883);
nor U3157 (N_3157,In_1905,In_1144);
and U3158 (N_3158,In_1270,In_328);
and U3159 (N_3159,In_173,In_1788);
nor U3160 (N_3160,In_1502,In_1704);
nor U3161 (N_3161,In_253,In_940);
and U3162 (N_3162,In_1655,In_1728);
and U3163 (N_3163,In_710,In_162);
nand U3164 (N_3164,In_710,In_1907);
xor U3165 (N_3165,In_1450,In_1773);
nand U3166 (N_3166,In_1559,In_240);
nand U3167 (N_3167,In_1090,In_336);
nand U3168 (N_3168,In_1565,In_105);
or U3169 (N_3169,In_682,In_968);
nand U3170 (N_3170,In_1651,In_288);
or U3171 (N_3171,In_97,In_1467);
and U3172 (N_3172,In_1269,In_1725);
and U3173 (N_3173,In_1495,In_893);
nor U3174 (N_3174,In_1420,In_1112);
and U3175 (N_3175,In_1561,In_26);
nand U3176 (N_3176,In_1749,In_606);
and U3177 (N_3177,In_1996,In_1955);
nor U3178 (N_3178,In_1009,In_648);
nand U3179 (N_3179,In_1829,In_335);
and U3180 (N_3180,In_60,In_1130);
nand U3181 (N_3181,In_1958,In_1582);
nand U3182 (N_3182,In_1053,In_13);
or U3183 (N_3183,In_1380,In_308);
or U3184 (N_3184,In_1389,In_1561);
nand U3185 (N_3185,In_1003,In_433);
and U3186 (N_3186,In_496,In_145);
and U3187 (N_3187,In_1557,In_1467);
and U3188 (N_3188,In_1077,In_83);
nor U3189 (N_3189,In_1396,In_371);
and U3190 (N_3190,In_1293,In_1191);
and U3191 (N_3191,In_1515,In_508);
or U3192 (N_3192,In_654,In_693);
nand U3193 (N_3193,In_506,In_15);
nand U3194 (N_3194,In_1600,In_223);
nor U3195 (N_3195,In_1349,In_1524);
and U3196 (N_3196,In_1430,In_1300);
xor U3197 (N_3197,In_557,In_956);
nand U3198 (N_3198,In_821,In_1821);
nor U3199 (N_3199,In_1838,In_478);
and U3200 (N_3200,In_41,In_302);
and U3201 (N_3201,In_736,In_479);
nor U3202 (N_3202,In_1934,In_418);
nor U3203 (N_3203,In_1218,In_464);
nand U3204 (N_3204,In_55,In_204);
and U3205 (N_3205,In_1960,In_1821);
nor U3206 (N_3206,In_916,In_1721);
nor U3207 (N_3207,In_775,In_792);
or U3208 (N_3208,In_1240,In_714);
nand U3209 (N_3209,In_1780,In_282);
and U3210 (N_3210,In_1277,In_624);
or U3211 (N_3211,In_220,In_1742);
or U3212 (N_3212,In_1520,In_389);
nor U3213 (N_3213,In_1465,In_792);
and U3214 (N_3214,In_1793,In_1063);
nor U3215 (N_3215,In_1000,In_1726);
and U3216 (N_3216,In_1434,In_1742);
and U3217 (N_3217,In_10,In_1785);
nor U3218 (N_3218,In_10,In_1618);
nor U3219 (N_3219,In_729,In_1890);
nor U3220 (N_3220,In_1045,In_1375);
nand U3221 (N_3221,In_508,In_17);
nand U3222 (N_3222,In_12,In_1285);
nand U3223 (N_3223,In_867,In_1457);
nor U3224 (N_3224,In_818,In_423);
or U3225 (N_3225,In_492,In_987);
and U3226 (N_3226,In_235,In_1937);
or U3227 (N_3227,In_1145,In_1633);
and U3228 (N_3228,In_1861,In_834);
nand U3229 (N_3229,In_833,In_278);
nand U3230 (N_3230,In_1292,In_1147);
nand U3231 (N_3231,In_958,In_1732);
and U3232 (N_3232,In_1664,In_722);
or U3233 (N_3233,In_1149,In_1869);
nand U3234 (N_3234,In_1108,In_295);
nor U3235 (N_3235,In_1043,In_1821);
nor U3236 (N_3236,In_620,In_174);
or U3237 (N_3237,In_1488,In_1258);
nand U3238 (N_3238,In_1804,In_634);
and U3239 (N_3239,In_306,In_93);
and U3240 (N_3240,In_1674,In_1477);
or U3241 (N_3241,In_1630,In_1641);
and U3242 (N_3242,In_986,In_1359);
and U3243 (N_3243,In_209,In_139);
nor U3244 (N_3244,In_495,In_1757);
nor U3245 (N_3245,In_284,In_1668);
and U3246 (N_3246,In_1089,In_602);
and U3247 (N_3247,In_602,In_161);
or U3248 (N_3248,In_1338,In_308);
or U3249 (N_3249,In_878,In_668);
or U3250 (N_3250,In_1211,In_106);
nand U3251 (N_3251,In_1200,In_372);
and U3252 (N_3252,In_960,In_993);
nand U3253 (N_3253,In_1373,In_1948);
xnor U3254 (N_3254,In_32,In_1353);
nand U3255 (N_3255,In_792,In_1143);
nand U3256 (N_3256,In_1974,In_515);
and U3257 (N_3257,In_1887,In_739);
and U3258 (N_3258,In_1640,In_434);
or U3259 (N_3259,In_1598,In_69);
nor U3260 (N_3260,In_1186,In_1242);
and U3261 (N_3261,In_188,In_711);
or U3262 (N_3262,In_314,In_1204);
nand U3263 (N_3263,In_1991,In_1369);
nand U3264 (N_3264,In_1094,In_1586);
and U3265 (N_3265,In_188,In_971);
xor U3266 (N_3266,In_265,In_1778);
nor U3267 (N_3267,In_833,In_668);
and U3268 (N_3268,In_453,In_1009);
nor U3269 (N_3269,In_1495,In_805);
nor U3270 (N_3270,In_1319,In_602);
and U3271 (N_3271,In_1729,In_447);
nor U3272 (N_3272,In_661,In_1634);
nor U3273 (N_3273,In_631,In_711);
and U3274 (N_3274,In_952,In_589);
and U3275 (N_3275,In_9,In_1698);
nor U3276 (N_3276,In_725,In_1261);
or U3277 (N_3277,In_509,In_1305);
or U3278 (N_3278,In_624,In_1861);
nand U3279 (N_3279,In_1682,In_1517);
and U3280 (N_3280,In_742,In_1461);
nand U3281 (N_3281,In_1275,In_1638);
or U3282 (N_3282,In_186,In_1995);
nand U3283 (N_3283,In_1779,In_220);
and U3284 (N_3284,In_1930,In_19);
nor U3285 (N_3285,In_295,In_1276);
and U3286 (N_3286,In_1714,In_1215);
or U3287 (N_3287,In_1766,In_293);
nor U3288 (N_3288,In_503,In_880);
and U3289 (N_3289,In_436,In_335);
nor U3290 (N_3290,In_1974,In_1677);
or U3291 (N_3291,In_817,In_1222);
nand U3292 (N_3292,In_1780,In_1844);
or U3293 (N_3293,In_773,In_1245);
or U3294 (N_3294,In_809,In_4);
nor U3295 (N_3295,In_916,In_1487);
nand U3296 (N_3296,In_1548,In_952);
nor U3297 (N_3297,In_706,In_1144);
nand U3298 (N_3298,In_1754,In_353);
and U3299 (N_3299,In_1035,In_898);
nor U3300 (N_3300,In_258,In_497);
and U3301 (N_3301,In_147,In_1904);
nor U3302 (N_3302,In_1350,In_1439);
or U3303 (N_3303,In_1332,In_1094);
xnor U3304 (N_3304,In_215,In_1865);
and U3305 (N_3305,In_49,In_1544);
or U3306 (N_3306,In_806,In_69);
or U3307 (N_3307,In_182,In_1432);
or U3308 (N_3308,In_1967,In_900);
nor U3309 (N_3309,In_1256,In_1499);
nor U3310 (N_3310,In_199,In_150);
or U3311 (N_3311,In_1291,In_1967);
or U3312 (N_3312,In_610,In_921);
or U3313 (N_3313,In_1473,In_1637);
or U3314 (N_3314,In_869,In_932);
and U3315 (N_3315,In_1813,In_234);
or U3316 (N_3316,In_864,In_838);
nor U3317 (N_3317,In_718,In_873);
nand U3318 (N_3318,In_1476,In_1729);
or U3319 (N_3319,In_588,In_1805);
xor U3320 (N_3320,In_1463,In_55);
nor U3321 (N_3321,In_529,In_756);
or U3322 (N_3322,In_554,In_823);
nor U3323 (N_3323,In_663,In_930);
or U3324 (N_3324,In_506,In_1926);
and U3325 (N_3325,In_1702,In_1230);
or U3326 (N_3326,In_1584,In_671);
xor U3327 (N_3327,In_605,In_1133);
nor U3328 (N_3328,In_1269,In_1977);
and U3329 (N_3329,In_1357,In_1128);
nor U3330 (N_3330,In_417,In_1640);
or U3331 (N_3331,In_70,In_180);
nand U3332 (N_3332,In_1026,In_64);
nor U3333 (N_3333,In_1505,In_1400);
nor U3334 (N_3334,In_1463,In_1297);
and U3335 (N_3335,In_1099,In_1186);
or U3336 (N_3336,In_1489,In_1625);
and U3337 (N_3337,In_1487,In_1386);
or U3338 (N_3338,In_591,In_1615);
or U3339 (N_3339,In_1313,In_1153);
and U3340 (N_3340,In_172,In_1435);
nand U3341 (N_3341,In_28,In_1715);
nand U3342 (N_3342,In_1873,In_1338);
nand U3343 (N_3343,In_904,In_840);
nor U3344 (N_3344,In_682,In_1023);
nor U3345 (N_3345,In_1821,In_184);
nand U3346 (N_3346,In_809,In_933);
xor U3347 (N_3347,In_816,In_756);
or U3348 (N_3348,In_14,In_982);
or U3349 (N_3349,In_777,In_1901);
nor U3350 (N_3350,In_1262,In_1313);
nand U3351 (N_3351,In_1356,In_488);
or U3352 (N_3352,In_1148,In_403);
nor U3353 (N_3353,In_1590,In_6);
or U3354 (N_3354,In_1143,In_691);
or U3355 (N_3355,In_609,In_279);
or U3356 (N_3356,In_1021,In_58);
and U3357 (N_3357,In_747,In_1294);
nor U3358 (N_3358,In_1410,In_180);
nor U3359 (N_3359,In_1005,In_229);
nand U3360 (N_3360,In_1945,In_253);
and U3361 (N_3361,In_628,In_1905);
or U3362 (N_3362,In_57,In_1507);
nand U3363 (N_3363,In_1326,In_1921);
or U3364 (N_3364,In_1095,In_1043);
nor U3365 (N_3365,In_1699,In_423);
nand U3366 (N_3366,In_880,In_898);
nand U3367 (N_3367,In_1779,In_1195);
nor U3368 (N_3368,In_1521,In_1393);
or U3369 (N_3369,In_1192,In_1745);
and U3370 (N_3370,In_779,In_1343);
and U3371 (N_3371,In_1511,In_1898);
nor U3372 (N_3372,In_1438,In_130);
nor U3373 (N_3373,In_972,In_888);
and U3374 (N_3374,In_1737,In_1139);
nand U3375 (N_3375,In_1272,In_674);
nand U3376 (N_3376,In_698,In_276);
or U3377 (N_3377,In_893,In_1907);
nor U3378 (N_3378,In_1509,In_1829);
nor U3379 (N_3379,In_1349,In_127);
nand U3380 (N_3380,In_1603,In_773);
or U3381 (N_3381,In_1250,In_1220);
or U3382 (N_3382,In_1520,In_64);
nand U3383 (N_3383,In_1829,In_1904);
nand U3384 (N_3384,In_451,In_568);
nor U3385 (N_3385,In_658,In_375);
and U3386 (N_3386,In_801,In_34);
nor U3387 (N_3387,In_18,In_208);
nand U3388 (N_3388,In_1028,In_578);
nor U3389 (N_3389,In_656,In_1375);
and U3390 (N_3390,In_1294,In_1665);
nor U3391 (N_3391,In_1804,In_186);
nor U3392 (N_3392,In_472,In_1455);
and U3393 (N_3393,In_704,In_483);
or U3394 (N_3394,In_1683,In_1237);
or U3395 (N_3395,In_1973,In_116);
nor U3396 (N_3396,In_1411,In_1890);
and U3397 (N_3397,In_1104,In_1244);
or U3398 (N_3398,In_1716,In_1727);
nor U3399 (N_3399,In_34,In_1209);
and U3400 (N_3400,In_484,In_1044);
nand U3401 (N_3401,In_447,In_739);
xnor U3402 (N_3402,In_113,In_1244);
or U3403 (N_3403,In_1209,In_100);
nor U3404 (N_3404,In_1553,In_702);
or U3405 (N_3405,In_159,In_475);
nor U3406 (N_3406,In_1020,In_861);
nor U3407 (N_3407,In_1578,In_700);
nand U3408 (N_3408,In_1595,In_1579);
nand U3409 (N_3409,In_1381,In_1870);
nor U3410 (N_3410,In_1776,In_1932);
nor U3411 (N_3411,In_908,In_918);
nor U3412 (N_3412,In_1590,In_1870);
or U3413 (N_3413,In_1485,In_163);
nor U3414 (N_3414,In_72,In_1737);
nor U3415 (N_3415,In_1365,In_730);
and U3416 (N_3416,In_1790,In_1505);
nand U3417 (N_3417,In_1866,In_1383);
nor U3418 (N_3418,In_618,In_1310);
or U3419 (N_3419,In_1525,In_1305);
nand U3420 (N_3420,In_1616,In_1798);
nand U3421 (N_3421,In_878,In_960);
nor U3422 (N_3422,In_236,In_1884);
nor U3423 (N_3423,In_98,In_1932);
or U3424 (N_3424,In_898,In_643);
nor U3425 (N_3425,In_975,In_1037);
nand U3426 (N_3426,In_973,In_6);
or U3427 (N_3427,In_1567,In_1650);
xor U3428 (N_3428,In_1886,In_1733);
or U3429 (N_3429,In_439,In_344);
or U3430 (N_3430,In_1150,In_1228);
nor U3431 (N_3431,In_1928,In_429);
and U3432 (N_3432,In_525,In_1957);
nor U3433 (N_3433,In_606,In_5);
nand U3434 (N_3434,In_1107,In_1977);
nand U3435 (N_3435,In_869,In_118);
or U3436 (N_3436,In_1219,In_872);
or U3437 (N_3437,In_1285,In_1105);
or U3438 (N_3438,In_1134,In_104);
and U3439 (N_3439,In_236,In_547);
or U3440 (N_3440,In_864,In_1059);
or U3441 (N_3441,In_1723,In_1109);
or U3442 (N_3442,In_1741,In_241);
xor U3443 (N_3443,In_1502,In_1461);
nand U3444 (N_3444,In_173,In_1866);
and U3445 (N_3445,In_1233,In_1429);
or U3446 (N_3446,In_661,In_1393);
nor U3447 (N_3447,In_872,In_595);
nand U3448 (N_3448,In_1512,In_1209);
nand U3449 (N_3449,In_851,In_1249);
nor U3450 (N_3450,In_496,In_1809);
or U3451 (N_3451,In_1730,In_1106);
and U3452 (N_3452,In_1618,In_164);
nand U3453 (N_3453,In_328,In_1855);
nor U3454 (N_3454,In_492,In_877);
and U3455 (N_3455,In_609,In_287);
nor U3456 (N_3456,In_1087,In_1849);
and U3457 (N_3457,In_454,In_1878);
and U3458 (N_3458,In_1291,In_1507);
and U3459 (N_3459,In_563,In_240);
and U3460 (N_3460,In_558,In_1894);
nand U3461 (N_3461,In_1338,In_575);
and U3462 (N_3462,In_737,In_659);
and U3463 (N_3463,In_371,In_330);
and U3464 (N_3464,In_658,In_646);
xnor U3465 (N_3465,In_646,In_24);
nor U3466 (N_3466,In_936,In_1724);
nor U3467 (N_3467,In_371,In_261);
nand U3468 (N_3468,In_458,In_1465);
and U3469 (N_3469,In_839,In_1794);
and U3470 (N_3470,In_1334,In_461);
nor U3471 (N_3471,In_918,In_665);
or U3472 (N_3472,In_1033,In_792);
nor U3473 (N_3473,In_12,In_900);
nand U3474 (N_3474,In_468,In_1993);
nand U3475 (N_3475,In_1767,In_1613);
nor U3476 (N_3476,In_1442,In_1210);
nor U3477 (N_3477,In_1396,In_487);
or U3478 (N_3478,In_999,In_1574);
or U3479 (N_3479,In_152,In_1493);
nor U3480 (N_3480,In_625,In_699);
nor U3481 (N_3481,In_990,In_1571);
nand U3482 (N_3482,In_16,In_1575);
and U3483 (N_3483,In_1203,In_1842);
nor U3484 (N_3484,In_1006,In_1857);
and U3485 (N_3485,In_1297,In_1);
and U3486 (N_3486,In_1742,In_732);
nand U3487 (N_3487,In_1557,In_1861);
and U3488 (N_3488,In_1918,In_572);
nand U3489 (N_3489,In_1295,In_425);
and U3490 (N_3490,In_1482,In_50);
and U3491 (N_3491,In_908,In_1290);
nor U3492 (N_3492,In_1609,In_1602);
or U3493 (N_3493,In_558,In_1895);
or U3494 (N_3494,In_535,In_525);
nor U3495 (N_3495,In_1533,In_1084);
nor U3496 (N_3496,In_475,In_1421);
or U3497 (N_3497,In_140,In_929);
or U3498 (N_3498,In_1236,In_497);
nand U3499 (N_3499,In_1811,In_584);
nor U3500 (N_3500,In_991,In_1818);
and U3501 (N_3501,In_1200,In_650);
nor U3502 (N_3502,In_1219,In_1709);
or U3503 (N_3503,In_1077,In_1328);
or U3504 (N_3504,In_777,In_1823);
nor U3505 (N_3505,In_1746,In_1257);
nor U3506 (N_3506,In_827,In_624);
nand U3507 (N_3507,In_1274,In_472);
and U3508 (N_3508,In_327,In_746);
nor U3509 (N_3509,In_344,In_1534);
nand U3510 (N_3510,In_1032,In_1275);
nand U3511 (N_3511,In_78,In_714);
or U3512 (N_3512,In_1435,In_1266);
nand U3513 (N_3513,In_619,In_1709);
nor U3514 (N_3514,In_36,In_1504);
nor U3515 (N_3515,In_1159,In_1892);
and U3516 (N_3516,In_1449,In_251);
nor U3517 (N_3517,In_326,In_131);
and U3518 (N_3518,In_1981,In_1427);
or U3519 (N_3519,In_1232,In_108);
nor U3520 (N_3520,In_1793,In_1941);
nor U3521 (N_3521,In_1321,In_464);
or U3522 (N_3522,In_1858,In_1369);
nor U3523 (N_3523,In_1682,In_119);
nor U3524 (N_3524,In_1574,In_819);
nor U3525 (N_3525,In_333,In_275);
nand U3526 (N_3526,In_961,In_924);
nand U3527 (N_3527,In_1131,In_1490);
nor U3528 (N_3528,In_1444,In_1771);
nor U3529 (N_3529,In_1843,In_50);
nor U3530 (N_3530,In_264,In_555);
and U3531 (N_3531,In_1757,In_1678);
nand U3532 (N_3532,In_1530,In_478);
and U3533 (N_3533,In_793,In_127);
nand U3534 (N_3534,In_1763,In_1798);
nor U3535 (N_3535,In_977,In_1170);
and U3536 (N_3536,In_467,In_1383);
and U3537 (N_3537,In_985,In_1448);
nand U3538 (N_3538,In_184,In_1165);
or U3539 (N_3539,In_1321,In_1462);
nand U3540 (N_3540,In_1193,In_1904);
or U3541 (N_3541,In_1572,In_830);
and U3542 (N_3542,In_1160,In_470);
nor U3543 (N_3543,In_311,In_243);
xnor U3544 (N_3544,In_1149,In_1081);
and U3545 (N_3545,In_1177,In_653);
xor U3546 (N_3546,In_1962,In_616);
nand U3547 (N_3547,In_848,In_838);
xnor U3548 (N_3548,In_1308,In_1219);
nand U3549 (N_3549,In_1277,In_1083);
or U3550 (N_3550,In_1161,In_1717);
or U3551 (N_3551,In_962,In_1525);
nor U3552 (N_3552,In_1546,In_1900);
and U3553 (N_3553,In_1943,In_1346);
or U3554 (N_3554,In_818,In_550);
nor U3555 (N_3555,In_462,In_1890);
or U3556 (N_3556,In_28,In_396);
and U3557 (N_3557,In_1856,In_1503);
and U3558 (N_3558,In_147,In_1664);
nor U3559 (N_3559,In_1613,In_657);
nor U3560 (N_3560,In_1336,In_1826);
nand U3561 (N_3561,In_708,In_249);
and U3562 (N_3562,In_762,In_784);
or U3563 (N_3563,In_481,In_1818);
nand U3564 (N_3564,In_19,In_795);
or U3565 (N_3565,In_1163,In_1987);
nor U3566 (N_3566,In_308,In_916);
and U3567 (N_3567,In_1558,In_688);
nand U3568 (N_3568,In_1563,In_192);
and U3569 (N_3569,In_1724,In_318);
or U3570 (N_3570,In_1922,In_604);
nor U3571 (N_3571,In_241,In_590);
nand U3572 (N_3572,In_868,In_1297);
or U3573 (N_3573,In_356,In_1547);
nand U3574 (N_3574,In_1865,In_1867);
nand U3575 (N_3575,In_1889,In_755);
xor U3576 (N_3576,In_1503,In_1538);
and U3577 (N_3577,In_1146,In_556);
or U3578 (N_3578,In_678,In_1728);
nor U3579 (N_3579,In_1628,In_908);
nor U3580 (N_3580,In_1095,In_985);
nand U3581 (N_3581,In_1949,In_1279);
nand U3582 (N_3582,In_1897,In_874);
or U3583 (N_3583,In_802,In_675);
nand U3584 (N_3584,In_1349,In_1890);
and U3585 (N_3585,In_1682,In_1186);
or U3586 (N_3586,In_248,In_853);
nor U3587 (N_3587,In_1713,In_21);
nand U3588 (N_3588,In_1738,In_370);
and U3589 (N_3589,In_219,In_1145);
nor U3590 (N_3590,In_146,In_144);
and U3591 (N_3591,In_872,In_977);
or U3592 (N_3592,In_288,In_39);
nor U3593 (N_3593,In_1039,In_61);
and U3594 (N_3594,In_1344,In_258);
nor U3595 (N_3595,In_1702,In_1933);
or U3596 (N_3596,In_1890,In_1502);
nor U3597 (N_3597,In_206,In_1196);
or U3598 (N_3598,In_1801,In_1726);
or U3599 (N_3599,In_1518,In_568);
nor U3600 (N_3600,In_896,In_424);
or U3601 (N_3601,In_1554,In_559);
and U3602 (N_3602,In_1714,In_96);
and U3603 (N_3603,In_1972,In_390);
or U3604 (N_3604,In_153,In_504);
nor U3605 (N_3605,In_97,In_213);
and U3606 (N_3606,In_1022,In_1761);
nor U3607 (N_3607,In_960,In_694);
nor U3608 (N_3608,In_48,In_393);
nand U3609 (N_3609,In_596,In_1738);
or U3610 (N_3610,In_571,In_1702);
nor U3611 (N_3611,In_678,In_1172);
or U3612 (N_3612,In_1301,In_726);
or U3613 (N_3613,In_1533,In_660);
nor U3614 (N_3614,In_1815,In_387);
nor U3615 (N_3615,In_617,In_780);
or U3616 (N_3616,In_839,In_1924);
nor U3617 (N_3617,In_1261,In_876);
and U3618 (N_3618,In_800,In_492);
and U3619 (N_3619,In_1723,In_1560);
nor U3620 (N_3620,In_1053,In_1058);
and U3621 (N_3621,In_1287,In_741);
nor U3622 (N_3622,In_1664,In_590);
nand U3623 (N_3623,In_283,In_1997);
and U3624 (N_3624,In_1425,In_282);
and U3625 (N_3625,In_1625,In_1320);
or U3626 (N_3626,In_252,In_894);
nor U3627 (N_3627,In_1783,In_1520);
xor U3628 (N_3628,In_1108,In_791);
or U3629 (N_3629,In_1953,In_1540);
or U3630 (N_3630,In_820,In_750);
or U3631 (N_3631,In_1406,In_1036);
nand U3632 (N_3632,In_1600,In_875);
or U3633 (N_3633,In_1828,In_1685);
nand U3634 (N_3634,In_748,In_1175);
and U3635 (N_3635,In_393,In_246);
nand U3636 (N_3636,In_1352,In_1486);
nor U3637 (N_3637,In_1224,In_843);
or U3638 (N_3638,In_122,In_1225);
nor U3639 (N_3639,In_125,In_1876);
nand U3640 (N_3640,In_1655,In_1830);
or U3641 (N_3641,In_1223,In_838);
and U3642 (N_3642,In_1570,In_533);
or U3643 (N_3643,In_599,In_736);
nor U3644 (N_3644,In_728,In_1607);
nand U3645 (N_3645,In_761,In_583);
nor U3646 (N_3646,In_397,In_262);
nand U3647 (N_3647,In_941,In_1954);
nand U3648 (N_3648,In_500,In_236);
or U3649 (N_3649,In_1809,In_1643);
or U3650 (N_3650,In_586,In_544);
or U3651 (N_3651,In_1951,In_187);
nor U3652 (N_3652,In_1100,In_1853);
and U3653 (N_3653,In_589,In_1445);
or U3654 (N_3654,In_891,In_271);
nor U3655 (N_3655,In_1301,In_431);
nand U3656 (N_3656,In_1321,In_967);
nand U3657 (N_3657,In_381,In_209);
and U3658 (N_3658,In_1562,In_1511);
nand U3659 (N_3659,In_1123,In_690);
nand U3660 (N_3660,In_642,In_1419);
nand U3661 (N_3661,In_1362,In_88);
and U3662 (N_3662,In_311,In_1997);
and U3663 (N_3663,In_224,In_519);
nor U3664 (N_3664,In_1034,In_923);
and U3665 (N_3665,In_202,In_1188);
nand U3666 (N_3666,In_1476,In_1016);
or U3667 (N_3667,In_1925,In_248);
nor U3668 (N_3668,In_1755,In_1931);
or U3669 (N_3669,In_149,In_931);
or U3670 (N_3670,In_1217,In_804);
and U3671 (N_3671,In_500,In_913);
xnor U3672 (N_3672,In_1722,In_1981);
nand U3673 (N_3673,In_1179,In_1876);
or U3674 (N_3674,In_1607,In_785);
or U3675 (N_3675,In_588,In_1629);
nand U3676 (N_3676,In_1185,In_1094);
nor U3677 (N_3677,In_499,In_417);
nor U3678 (N_3678,In_1148,In_1466);
xnor U3679 (N_3679,In_799,In_479);
or U3680 (N_3680,In_1903,In_1252);
or U3681 (N_3681,In_152,In_745);
nor U3682 (N_3682,In_1822,In_1828);
or U3683 (N_3683,In_1463,In_1944);
nand U3684 (N_3684,In_609,In_1352);
and U3685 (N_3685,In_1355,In_623);
and U3686 (N_3686,In_652,In_1518);
nand U3687 (N_3687,In_443,In_1223);
nand U3688 (N_3688,In_1209,In_699);
or U3689 (N_3689,In_1067,In_1030);
nand U3690 (N_3690,In_1718,In_1728);
nor U3691 (N_3691,In_1926,In_842);
nand U3692 (N_3692,In_1697,In_1693);
and U3693 (N_3693,In_1237,In_1125);
nor U3694 (N_3694,In_1150,In_1590);
and U3695 (N_3695,In_765,In_1517);
or U3696 (N_3696,In_623,In_1282);
nor U3697 (N_3697,In_927,In_734);
and U3698 (N_3698,In_76,In_683);
or U3699 (N_3699,In_1544,In_1562);
or U3700 (N_3700,In_1466,In_1411);
nor U3701 (N_3701,In_1117,In_1029);
or U3702 (N_3702,In_321,In_1082);
nand U3703 (N_3703,In_1576,In_1973);
or U3704 (N_3704,In_371,In_90);
nor U3705 (N_3705,In_1471,In_259);
nor U3706 (N_3706,In_282,In_799);
nor U3707 (N_3707,In_1803,In_1445);
nand U3708 (N_3708,In_1300,In_1643);
or U3709 (N_3709,In_524,In_1383);
nor U3710 (N_3710,In_481,In_955);
nand U3711 (N_3711,In_1003,In_1470);
nand U3712 (N_3712,In_847,In_1479);
nand U3713 (N_3713,In_1497,In_69);
nor U3714 (N_3714,In_1884,In_354);
nand U3715 (N_3715,In_804,In_1722);
and U3716 (N_3716,In_1496,In_1550);
or U3717 (N_3717,In_1186,In_905);
nand U3718 (N_3718,In_1212,In_1298);
nand U3719 (N_3719,In_1627,In_234);
nor U3720 (N_3720,In_1180,In_1577);
or U3721 (N_3721,In_108,In_1249);
xnor U3722 (N_3722,In_617,In_776);
and U3723 (N_3723,In_1178,In_547);
nor U3724 (N_3724,In_554,In_416);
nand U3725 (N_3725,In_396,In_331);
or U3726 (N_3726,In_1305,In_1468);
and U3727 (N_3727,In_432,In_1877);
nand U3728 (N_3728,In_760,In_1475);
nand U3729 (N_3729,In_145,In_1957);
xnor U3730 (N_3730,In_0,In_549);
nand U3731 (N_3731,In_545,In_944);
nand U3732 (N_3732,In_392,In_1094);
nor U3733 (N_3733,In_1314,In_833);
or U3734 (N_3734,In_1611,In_1311);
nor U3735 (N_3735,In_1851,In_115);
nor U3736 (N_3736,In_624,In_733);
nor U3737 (N_3737,In_196,In_669);
nor U3738 (N_3738,In_178,In_310);
and U3739 (N_3739,In_132,In_1844);
and U3740 (N_3740,In_748,In_396);
nand U3741 (N_3741,In_1544,In_1419);
and U3742 (N_3742,In_1222,In_1624);
or U3743 (N_3743,In_1432,In_1431);
nor U3744 (N_3744,In_680,In_166);
nand U3745 (N_3745,In_88,In_258);
nor U3746 (N_3746,In_516,In_1220);
nand U3747 (N_3747,In_1200,In_1054);
or U3748 (N_3748,In_973,In_1373);
xnor U3749 (N_3749,In_1878,In_724);
nor U3750 (N_3750,In_688,In_393);
and U3751 (N_3751,In_1177,In_1128);
or U3752 (N_3752,In_840,In_1726);
nand U3753 (N_3753,In_1865,In_44);
and U3754 (N_3754,In_393,In_1365);
and U3755 (N_3755,In_1827,In_1192);
xor U3756 (N_3756,In_945,In_1423);
xor U3757 (N_3757,In_196,In_322);
and U3758 (N_3758,In_178,In_776);
nor U3759 (N_3759,In_582,In_1958);
nor U3760 (N_3760,In_1087,In_344);
nand U3761 (N_3761,In_1448,In_962);
nand U3762 (N_3762,In_1022,In_465);
nand U3763 (N_3763,In_1349,In_1874);
nor U3764 (N_3764,In_799,In_1783);
and U3765 (N_3765,In_1774,In_100);
nor U3766 (N_3766,In_975,In_143);
and U3767 (N_3767,In_84,In_365);
and U3768 (N_3768,In_409,In_104);
or U3769 (N_3769,In_466,In_1157);
nand U3770 (N_3770,In_1933,In_627);
and U3771 (N_3771,In_1959,In_1928);
nand U3772 (N_3772,In_545,In_1713);
nand U3773 (N_3773,In_465,In_1266);
nor U3774 (N_3774,In_758,In_1559);
and U3775 (N_3775,In_1488,In_138);
or U3776 (N_3776,In_492,In_918);
nand U3777 (N_3777,In_1495,In_476);
nor U3778 (N_3778,In_510,In_1689);
or U3779 (N_3779,In_1000,In_1959);
and U3780 (N_3780,In_386,In_1905);
nand U3781 (N_3781,In_1909,In_514);
nor U3782 (N_3782,In_900,In_340);
nor U3783 (N_3783,In_1034,In_187);
or U3784 (N_3784,In_1120,In_223);
or U3785 (N_3785,In_1629,In_1085);
nor U3786 (N_3786,In_1966,In_127);
and U3787 (N_3787,In_632,In_1387);
and U3788 (N_3788,In_1271,In_209);
and U3789 (N_3789,In_1293,In_206);
nor U3790 (N_3790,In_627,In_324);
or U3791 (N_3791,In_1123,In_1924);
or U3792 (N_3792,In_768,In_1066);
or U3793 (N_3793,In_836,In_271);
and U3794 (N_3794,In_810,In_1019);
and U3795 (N_3795,In_1030,In_558);
nor U3796 (N_3796,In_1399,In_730);
and U3797 (N_3797,In_1810,In_1889);
and U3798 (N_3798,In_782,In_733);
nand U3799 (N_3799,In_113,In_610);
and U3800 (N_3800,In_1140,In_1872);
xnor U3801 (N_3801,In_270,In_59);
nand U3802 (N_3802,In_1086,In_875);
or U3803 (N_3803,In_1418,In_1621);
nor U3804 (N_3804,In_35,In_874);
or U3805 (N_3805,In_1116,In_1154);
nor U3806 (N_3806,In_1894,In_1644);
or U3807 (N_3807,In_1344,In_1206);
nand U3808 (N_3808,In_1147,In_978);
nor U3809 (N_3809,In_325,In_228);
nand U3810 (N_3810,In_1548,In_225);
or U3811 (N_3811,In_1249,In_110);
xnor U3812 (N_3812,In_1047,In_1620);
xor U3813 (N_3813,In_373,In_1701);
xor U3814 (N_3814,In_1746,In_168);
xnor U3815 (N_3815,In_1557,In_722);
and U3816 (N_3816,In_545,In_392);
nor U3817 (N_3817,In_153,In_120);
nor U3818 (N_3818,In_1317,In_184);
and U3819 (N_3819,In_1715,In_280);
or U3820 (N_3820,In_1397,In_35);
nor U3821 (N_3821,In_559,In_1627);
nand U3822 (N_3822,In_681,In_1061);
nor U3823 (N_3823,In_1609,In_1141);
or U3824 (N_3824,In_390,In_451);
nand U3825 (N_3825,In_184,In_13);
xor U3826 (N_3826,In_1018,In_775);
nor U3827 (N_3827,In_572,In_651);
nand U3828 (N_3828,In_429,In_1431);
and U3829 (N_3829,In_828,In_491);
nand U3830 (N_3830,In_415,In_1833);
or U3831 (N_3831,In_1415,In_1091);
and U3832 (N_3832,In_1506,In_1580);
nand U3833 (N_3833,In_1540,In_775);
nor U3834 (N_3834,In_1424,In_1108);
and U3835 (N_3835,In_1656,In_797);
and U3836 (N_3836,In_1234,In_410);
nand U3837 (N_3837,In_393,In_1886);
xor U3838 (N_3838,In_334,In_1477);
and U3839 (N_3839,In_1767,In_1210);
and U3840 (N_3840,In_367,In_1415);
and U3841 (N_3841,In_1246,In_1666);
and U3842 (N_3842,In_656,In_1178);
nand U3843 (N_3843,In_1756,In_867);
nor U3844 (N_3844,In_1949,In_199);
nand U3845 (N_3845,In_964,In_402);
nand U3846 (N_3846,In_368,In_1831);
nand U3847 (N_3847,In_1424,In_639);
or U3848 (N_3848,In_68,In_822);
nor U3849 (N_3849,In_334,In_1895);
or U3850 (N_3850,In_1078,In_1269);
or U3851 (N_3851,In_821,In_105);
nand U3852 (N_3852,In_961,In_1212);
nor U3853 (N_3853,In_233,In_1168);
nor U3854 (N_3854,In_451,In_1377);
nand U3855 (N_3855,In_701,In_280);
xor U3856 (N_3856,In_708,In_886);
and U3857 (N_3857,In_338,In_168);
and U3858 (N_3858,In_307,In_1384);
or U3859 (N_3859,In_862,In_1072);
or U3860 (N_3860,In_169,In_1734);
nand U3861 (N_3861,In_1549,In_1734);
and U3862 (N_3862,In_1065,In_255);
nand U3863 (N_3863,In_591,In_1625);
and U3864 (N_3864,In_1813,In_1203);
or U3865 (N_3865,In_1244,In_146);
and U3866 (N_3866,In_111,In_1895);
nand U3867 (N_3867,In_43,In_2);
and U3868 (N_3868,In_573,In_1619);
nor U3869 (N_3869,In_1341,In_1065);
and U3870 (N_3870,In_5,In_1416);
or U3871 (N_3871,In_349,In_1797);
or U3872 (N_3872,In_1196,In_1263);
nor U3873 (N_3873,In_43,In_930);
nor U3874 (N_3874,In_1199,In_815);
or U3875 (N_3875,In_1527,In_413);
or U3876 (N_3876,In_94,In_1809);
nor U3877 (N_3877,In_1056,In_40);
nor U3878 (N_3878,In_830,In_946);
or U3879 (N_3879,In_1802,In_1700);
nand U3880 (N_3880,In_1148,In_93);
nor U3881 (N_3881,In_1824,In_341);
nor U3882 (N_3882,In_658,In_960);
or U3883 (N_3883,In_1163,In_1763);
nand U3884 (N_3884,In_90,In_1465);
or U3885 (N_3885,In_1722,In_1813);
nand U3886 (N_3886,In_767,In_332);
nor U3887 (N_3887,In_538,In_1026);
or U3888 (N_3888,In_1836,In_1946);
or U3889 (N_3889,In_573,In_137);
and U3890 (N_3890,In_526,In_1224);
and U3891 (N_3891,In_1748,In_489);
nand U3892 (N_3892,In_1756,In_1421);
or U3893 (N_3893,In_747,In_1119);
and U3894 (N_3894,In_432,In_1554);
xnor U3895 (N_3895,In_1060,In_419);
and U3896 (N_3896,In_195,In_1675);
or U3897 (N_3897,In_129,In_632);
and U3898 (N_3898,In_568,In_960);
nand U3899 (N_3899,In_83,In_251);
and U3900 (N_3900,In_40,In_857);
or U3901 (N_3901,In_785,In_1213);
and U3902 (N_3902,In_1677,In_1362);
or U3903 (N_3903,In_1754,In_944);
and U3904 (N_3904,In_1322,In_727);
nand U3905 (N_3905,In_1488,In_147);
nand U3906 (N_3906,In_515,In_1210);
nand U3907 (N_3907,In_823,In_873);
nor U3908 (N_3908,In_513,In_1560);
or U3909 (N_3909,In_264,In_497);
or U3910 (N_3910,In_326,In_1024);
or U3911 (N_3911,In_59,In_411);
and U3912 (N_3912,In_1838,In_925);
nand U3913 (N_3913,In_1753,In_1310);
and U3914 (N_3914,In_709,In_247);
or U3915 (N_3915,In_653,In_956);
xnor U3916 (N_3916,In_1628,In_1519);
or U3917 (N_3917,In_1648,In_1237);
nor U3918 (N_3918,In_886,In_1041);
and U3919 (N_3919,In_1923,In_621);
nor U3920 (N_3920,In_702,In_1205);
or U3921 (N_3921,In_805,In_654);
and U3922 (N_3922,In_1931,In_1859);
xnor U3923 (N_3923,In_1085,In_795);
and U3924 (N_3924,In_386,In_233);
and U3925 (N_3925,In_1842,In_26);
or U3926 (N_3926,In_930,In_1479);
xnor U3927 (N_3927,In_5,In_213);
and U3928 (N_3928,In_474,In_29);
or U3929 (N_3929,In_544,In_582);
and U3930 (N_3930,In_1986,In_479);
nand U3931 (N_3931,In_427,In_588);
and U3932 (N_3932,In_1903,In_1749);
nand U3933 (N_3933,In_699,In_108);
xor U3934 (N_3934,In_252,In_1671);
nand U3935 (N_3935,In_1166,In_1755);
or U3936 (N_3936,In_593,In_1824);
and U3937 (N_3937,In_967,In_397);
or U3938 (N_3938,In_830,In_339);
and U3939 (N_3939,In_1718,In_1556);
and U3940 (N_3940,In_1204,In_554);
nor U3941 (N_3941,In_468,In_93);
and U3942 (N_3942,In_1071,In_1565);
nand U3943 (N_3943,In_36,In_1013);
or U3944 (N_3944,In_332,In_447);
nor U3945 (N_3945,In_1425,In_601);
or U3946 (N_3946,In_1364,In_1994);
and U3947 (N_3947,In_1742,In_1429);
and U3948 (N_3948,In_1227,In_997);
and U3949 (N_3949,In_1589,In_881);
and U3950 (N_3950,In_425,In_1997);
or U3951 (N_3951,In_1567,In_1884);
nor U3952 (N_3952,In_741,In_1533);
and U3953 (N_3953,In_872,In_41);
and U3954 (N_3954,In_1223,In_92);
nand U3955 (N_3955,In_1206,In_258);
nor U3956 (N_3956,In_1057,In_1327);
and U3957 (N_3957,In_574,In_138);
or U3958 (N_3958,In_1395,In_690);
nand U3959 (N_3959,In_211,In_734);
nand U3960 (N_3960,In_184,In_42);
nand U3961 (N_3961,In_594,In_102);
or U3962 (N_3962,In_548,In_1578);
or U3963 (N_3963,In_384,In_1016);
nand U3964 (N_3964,In_1285,In_1018);
nor U3965 (N_3965,In_331,In_1201);
or U3966 (N_3966,In_1132,In_197);
nor U3967 (N_3967,In_1218,In_361);
or U3968 (N_3968,In_1932,In_982);
or U3969 (N_3969,In_1162,In_168);
or U3970 (N_3970,In_1823,In_1337);
and U3971 (N_3971,In_1434,In_114);
or U3972 (N_3972,In_620,In_1531);
nand U3973 (N_3973,In_1151,In_40);
or U3974 (N_3974,In_1790,In_1373);
nor U3975 (N_3975,In_428,In_1267);
nor U3976 (N_3976,In_36,In_1967);
nand U3977 (N_3977,In_1265,In_705);
nor U3978 (N_3978,In_1069,In_1179);
nand U3979 (N_3979,In_612,In_534);
nand U3980 (N_3980,In_933,In_300);
and U3981 (N_3981,In_1955,In_793);
or U3982 (N_3982,In_1851,In_55);
or U3983 (N_3983,In_1857,In_124);
xnor U3984 (N_3984,In_1301,In_1452);
nor U3985 (N_3985,In_1637,In_277);
nor U3986 (N_3986,In_1645,In_16);
nand U3987 (N_3987,In_1203,In_1670);
nand U3988 (N_3988,In_1401,In_1088);
nand U3989 (N_3989,In_1812,In_265);
nand U3990 (N_3990,In_910,In_48);
and U3991 (N_3991,In_1223,In_1715);
nand U3992 (N_3992,In_16,In_1767);
or U3993 (N_3993,In_1809,In_1124);
nand U3994 (N_3994,In_1927,In_1794);
and U3995 (N_3995,In_455,In_944);
and U3996 (N_3996,In_1518,In_800);
xor U3997 (N_3997,In_1691,In_575);
nor U3998 (N_3998,In_1831,In_1309);
or U3999 (N_3999,In_1655,In_1153);
xnor U4000 (N_4000,In_509,In_216);
nor U4001 (N_4001,In_1856,In_1491);
xnor U4002 (N_4002,In_1950,In_1475);
nor U4003 (N_4003,In_126,In_1492);
nand U4004 (N_4004,In_549,In_980);
nor U4005 (N_4005,In_1874,In_545);
nor U4006 (N_4006,In_536,In_1299);
or U4007 (N_4007,In_1404,In_1741);
nor U4008 (N_4008,In_1701,In_900);
or U4009 (N_4009,In_73,In_1171);
nor U4010 (N_4010,In_1478,In_91);
or U4011 (N_4011,In_1611,In_1341);
and U4012 (N_4012,In_885,In_1130);
nor U4013 (N_4013,In_1204,In_1535);
nor U4014 (N_4014,In_987,In_1892);
and U4015 (N_4015,In_1116,In_1210);
and U4016 (N_4016,In_1577,In_1122);
nand U4017 (N_4017,In_775,In_857);
or U4018 (N_4018,In_492,In_326);
and U4019 (N_4019,In_26,In_755);
and U4020 (N_4020,In_1463,In_274);
nand U4021 (N_4021,In_795,In_142);
and U4022 (N_4022,In_1243,In_1858);
nand U4023 (N_4023,In_1827,In_1617);
and U4024 (N_4024,In_1867,In_790);
or U4025 (N_4025,In_1599,In_1917);
or U4026 (N_4026,In_351,In_1941);
nor U4027 (N_4027,In_1543,In_1822);
nor U4028 (N_4028,In_266,In_1762);
nor U4029 (N_4029,In_1422,In_826);
nor U4030 (N_4030,In_1098,In_1413);
or U4031 (N_4031,In_263,In_213);
nand U4032 (N_4032,In_334,In_506);
or U4033 (N_4033,In_522,In_1961);
nand U4034 (N_4034,In_1340,In_1126);
nand U4035 (N_4035,In_1045,In_405);
xnor U4036 (N_4036,In_1333,In_1505);
and U4037 (N_4037,In_1414,In_1780);
nand U4038 (N_4038,In_282,In_1343);
and U4039 (N_4039,In_1560,In_1811);
nand U4040 (N_4040,In_995,In_1580);
nand U4041 (N_4041,In_676,In_898);
and U4042 (N_4042,In_20,In_1448);
and U4043 (N_4043,In_89,In_611);
nor U4044 (N_4044,In_1384,In_174);
nor U4045 (N_4045,In_1190,In_396);
nand U4046 (N_4046,In_1812,In_1586);
nand U4047 (N_4047,In_60,In_1809);
or U4048 (N_4048,In_850,In_1641);
nand U4049 (N_4049,In_1549,In_1794);
nand U4050 (N_4050,In_285,In_270);
nand U4051 (N_4051,In_1183,In_1616);
and U4052 (N_4052,In_661,In_1892);
or U4053 (N_4053,In_1777,In_1878);
or U4054 (N_4054,In_714,In_1606);
nor U4055 (N_4055,In_1665,In_1614);
nand U4056 (N_4056,In_1367,In_1807);
nor U4057 (N_4057,In_1482,In_1816);
nor U4058 (N_4058,In_471,In_285);
and U4059 (N_4059,In_212,In_732);
and U4060 (N_4060,In_1779,In_1938);
or U4061 (N_4061,In_302,In_1548);
nor U4062 (N_4062,In_336,In_827);
and U4063 (N_4063,In_436,In_1839);
and U4064 (N_4064,In_941,In_581);
nand U4065 (N_4065,In_772,In_416);
and U4066 (N_4066,In_708,In_45);
or U4067 (N_4067,In_707,In_1049);
nand U4068 (N_4068,In_172,In_320);
or U4069 (N_4069,In_1490,In_1127);
or U4070 (N_4070,In_272,In_1191);
nor U4071 (N_4071,In_1965,In_1231);
nor U4072 (N_4072,In_336,In_1301);
and U4073 (N_4073,In_245,In_1494);
or U4074 (N_4074,In_1330,In_1919);
nor U4075 (N_4075,In_166,In_95);
and U4076 (N_4076,In_975,In_446);
nand U4077 (N_4077,In_1275,In_41);
or U4078 (N_4078,In_1455,In_803);
nor U4079 (N_4079,In_1381,In_1427);
nand U4080 (N_4080,In_1767,In_1569);
nor U4081 (N_4081,In_1512,In_1164);
nand U4082 (N_4082,In_664,In_1600);
nand U4083 (N_4083,In_883,In_265);
nand U4084 (N_4084,In_451,In_947);
nand U4085 (N_4085,In_288,In_1381);
nor U4086 (N_4086,In_1504,In_1120);
or U4087 (N_4087,In_727,In_1017);
nand U4088 (N_4088,In_1006,In_1836);
or U4089 (N_4089,In_1351,In_1535);
or U4090 (N_4090,In_1415,In_1541);
nor U4091 (N_4091,In_96,In_439);
nand U4092 (N_4092,In_1576,In_1374);
nand U4093 (N_4093,In_1240,In_32);
or U4094 (N_4094,In_61,In_1828);
nand U4095 (N_4095,In_228,In_1074);
nor U4096 (N_4096,In_688,In_1933);
nor U4097 (N_4097,In_1650,In_386);
nand U4098 (N_4098,In_453,In_906);
and U4099 (N_4099,In_902,In_1804);
nand U4100 (N_4100,In_1610,In_1963);
xnor U4101 (N_4101,In_1100,In_1704);
nor U4102 (N_4102,In_509,In_1652);
nor U4103 (N_4103,In_1541,In_181);
nor U4104 (N_4104,In_45,In_1547);
nand U4105 (N_4105,In_685,In_699);
nand U4106 (N_4106,In_1557,In_444);
or U4107 (N_4107,In_1747,In_1926);
or U4108 (N_4108,In_1983,In_837);
nor U4109 (N_4109,In_655,In_719);
nor U4110 (N_4110,In_935,In_1416);
nor U4111 (N_4111,In_659,In_652);
nand U4112 (N_4112,In_1670,In_1289);
or U4113 (N_4113,In_243,In_24);
and U4114 (N_4114,In_1400,In_626);
nor U4115 (N_4115,In_1763,In_1941);
or U4116 (N_4116,In_44,In_1247);
nor U4117 (N_4117,In_105,In_1265);
nand U4118 (N_4118,In_321,In_626);
and U4119 (N_4119,In_1494,In_1509);
and U4120 (N_4120,In_491,In_1523);
nor U4121 (N_4121,In_145,In_1149);
and U4122 (N_4122,In_457,In_74);
and U4123 (N_4123,In_944,In_486);
xor U4124 (N_4124,In_1038,In_679);
and U4125 (N_4125,In_1194,In_748);
and U4126 (N_4126,In_1502,In_1541);
or U4127 (N_4127,In_946,In_1657);
and U4128 (N_4128,In_1044,In_577);
or U4129 (N_4129,In_793,In_1688);
nand U4130 (N_4130,In_1295,In_1556);
nor U4131 (N_4131,In_1156,In_1497);
nor U4132 (N_4132,In_610,In_1208);
or U4133 (N_4133,In_1438,In_837);
or U4134 (N_4134,In_1853,In_852);
nand U4135 (N_4135,In_85,In_615);
nand U4136 (N_4136,In_658,In_86);
and U4137 (N_4137,In_1339,In_1133);
or U4138 (N_4138,In_208,In_801);
nand U4139 (N_4139,In_270,In_696);
nor U4140 (N_4140,In_194,In_961);
nor U4141 (N_4141,In_123,In_1622);
and U4142 (N_4142,In_930,In_441);
and U4143 (N_4143,In_1639,In_94);
and U4144 (N_4144,In_413,In_490);
nor U4145 (N_4145,In_1062,In_1401);
and U4146 (N_4146,In_77,In_1915);
nor U4147 (N_4147,In_1573,In_435);
nor U4148 (N_4148,In_161,In_217);
nand U4149 (N_4149,In_728,In_1855);
nand U4150 (N_4150,In_1239,In_309);
nor U4151 (N_4151,In_1590,In_1481);
nand U4152 (N_4152,In_737,In_1992);
nand U4153 (N_4153,In_1039,In_1337);
nor U4154 (N_4154,In_1623,In_525);
nor U4155 (N_4155,In_299,In_1619);
and U4156 (N_4156,In_1940,In_1153);
and U4157 (N_4157,In_1881,In_177);
nand U4158 (N_4158,In_1010,In_390);
nor U4159 (N_4159,In_39,In_1863);
or U4160 (N_4160,In_1938,In_663);
nor U4161 (N_4161,In_946,In_467);
nor U4162 (N_4162,In_749,In_133);
and U4163 (N_4163,In_1988,In_1404);
nor U4164 (N_4164,In_159,In_507);
or U4165 (N_4165,In_1617,In_1507);
nand U4166 (N_4166,In_1111,In_134);
and U4167 (N_4167,In_1746,In_540);
and U4168 (N_4168,In_673,In_1887);
and U4169 (N_4169,In_952,In_918);
nand U4170 (N_4170,In_1900,In_1645);
nor U4171 (N_4171,In_215,In_1725);
or U4172 (N_4172,In_111,In_114);
nand U4173 (N_4173,In_1545,In_764);
or U4174 (N_4174,In_703,In_116);
nand U4175 (N_4175,In_1380,In_1606);
and U4176 (N_4176,In_366,In_1963);
nand U4177 (N_4177,In_951,In_828);
nand U4178 (N_4178,In_701,In_1537);
or U4179 (N_4179,In_1675,In_1811);
or U4180 (N_4180,In_277,In_1175);
nor U4181 (N_4181,In_1059,In_430);
or U4182 (N_4182,In_245,In_713);
and U4183 (N_4183,In_829,In_1007);
and U4184 (N_4184,In_505,In_162);
nor U4185 (N_4185,In_132,In_1089);
nand U4186 (N_4186,In_223,In_1403);
or U4187 (N_4187,In_301,In_157);
nand U4188 (N_4188,In_1801,In_195);
nor U4189 (N_4189,In_716,In_77);
or U4190 (N_4190,In_7,In_1638);
nand U4191 (N_4191,In_893,In_82);
or U4192 (N_4192,In_803,In_1268);
or U4193 (N_4193,In_1600,In_605);
and U4194 (N_4194,In_187,In_886);
and U4195 (N_4195,In_886,In_589);
nor U4196 (N_4196,In_983,In_1186);
or U4197 (N_4197,In_592,In_477);
nor U4198 (N_4198,In_453,In_246);
nor U4199 (N_4199,In_1009,In_517);
nand U4200 (N_4200,In_909,In_88);
nand U4201 (N_4201,In_1547,In_302);
nand U4202 (N_4202,In_718,In_1521);
nand U4203 (N_4203,In_1288,In_1489);
or U4204 (N_4204,In_573,In_1318);
or U4205 (N_4205,In_1925,In_1937);
nor U4206 (N_4206,In_299,In_1796);
nand U4207 (N_4207,In_1597,In_83);
or U4208 (N_4208,In_470,In_1179);
or U4209 (N_4209,In_1129,In_297);
nand U4210 (N_4210,In_905,In_58);
and U4211 (N_4211,In_1826,In_1387);
nor U4212 (N_4212,In_726,In_1843);
and U4213 (N_4213,In_75,In_929);
and U4214 (N_4214,In_1862,In_773);
nor U4215 (N_4215,In_787,In_818);
nand U4216 (N_4216,In_362,In_1084);
and U4217 (N_4217,In_896,In_1236);
nor U4218 (N_4218,In_607,In_215);
nand U4219 (N_4219,In_76,In_498);
nor U4220 (N_4220,In_1321,In_1733);
and U4221 (N_4221,In_34,In_1378);
nand U4222 (N_4222,In_439,In_1089);
and U4223 (N_4223,In_331,In_702);
or U4224 (N_4224,In_1358,In_909);
nor U4225 (N_4225,In_1549,In_1601);
or U4226 (N_4226,In_1311,In_1823);
or U4227 (N_4227,In_1429,In_1887);
or U4228 (N_4228,In_28,In_596);
or U4229 (N_4229,In_390,In_261);
nor U4230 (N_4230,In_1661,In_1398);
or U4231 (N_4231,In_1853,In_704);
and U4232 (N_4232,In_19,In_455);
nand U4233 (N_4233,In_687,In_1644);
nand U4234 (N_4234,In_776,In_1684);
or U4235 (N_4235,In_1083,In_1938);
xnor U4236 (N_4236,In_140,In_921);
or U4237 (N_4237,In_913,In_1065);
and U4238 (N_4238,In_614,In_1088);
nor U4239 (N_4239,In_1424,In_807);
nor U4240 (N_4240,In_1903,In_1023);
nand U4241 (N_4241,In_1341,In_1323);
nor U4242 (N_4242,In_1945,In_628);
and U4243 (N_4243,In_631,In_1454);
nor U4244 (N_4244,In_1987,In_524);
nand U4245 (N_4245,In_215,In_1913);
nand U4246 (N_4246,In_1885,In_969);
nand U4247 (N_4247,In_1801,In_875);
or U4248 (N_4248,In_619,In_1074);
and U4249 (N_4249,In_1801,In_1932);
and U4250 (N_4250,In_1081,In_784);
nand U4251 (N_4251,In_625,In_1598);
or U4252 (N_4252,In_188,In_983);
or U4253 (N_4253,In_1233,In_1501);
and U4254 (N_4254,In_1041,In_833);
nor U4255 (N_4255,In_1233,In_915);
nor U4256 (N_4256,In_871,In_999);
nor U4257 (N_4257,In_251,In_1567);
nor U4258 (N_4258,In_1648,In_1791);
or U4259 (N_4259,In_1952,In_412);
and U4260 (N_4260,In_1702,In_255);
or U4261 (N_4261,In_535,In_1902);
and U4262 (N_4262,In_956,In_1519);
nand U4263 (N_4263,In_1043,In_1925);
nand U4264 (N_4264,In_1991,In_390);
or U4265 (N_4265,In_698,In_1493);
nand U4266 (N_4266,In_1725,In_1187);
or U4267 (N_4267,In_249,In_1053);
nor U4268 (N_4268,In_932,In_1554);
or U4269 (N_4269,In_1191,In_1621);
and U4270 (N_4270,In_1723,In_1065);
nand U4271 (N_4271,In_1122,In_1141);
nand U4272 (N_4272,In_1322,In_54);
or U4273 (N_4273,In_1203,In_1980);
and U4274 (N_4274,In_1412,In_1487);
nor U4275 (N_4275,In_703,In_990);
nand U4276 (N_4276,In_991,In_302);
nor U4277 (N_4277,In_1942,In_431);
nor U4278 (N_4278,In_1280,In_1180);
or U4279 (N_4279,In_1998,In_1497);
nor U4280 (N_4280,In_1300,In_1276);
nor U4281 (N_4281,In_1355,In_1128);
nand U4282 (N_4282,In_1836,In_1786);
or U4283 (N_4283,In_281,In_867);
nor U4284 (N_4284,In_1240,In_1700);
and U4285 (N_4285,In_256,In_1889);
and U4286 (N_4286,In_1981,In_13);
or U4287 (N_4287,In_869,In_1918);
nand U4288 (N_4288,In_875,In_109);
and U4289 (N_4289,In_1970,In_1472);
or U4290 (N_4290,In_1789,In_1631);
nor U4291 (N_4291,In_441,In_1379);
nor U4292 (N_4292,In_380,In_272);
nor U4293 (N_4293,In_199,In_1695);
nor U4294 (N_4294,In_143,In_119);
nand U4295 (N_4295,In_1908,In_854);
nand U4296 (N_4296,In_1139,In_992);
nor U4297 (N_4297,In_65,In_415);
and U4298 (N_4298,In_769,In_1927);
nor U4299 (N_4299,In_267,In_1622);
or U4300 (N_4300,In_508,In_1270);
nand U4301 (N_4301,In_228,In_1224);
nand U4302 (N_4302,In_1505,In_1034);
nand U4303 (N_4303,In_1920,In_1912);
nand U4304 (N_4304,In_1672,In_1009);
nor U4305 (N_4305,In_1410,In_443);
nor U4306 (N_4306,In_445,In_139);
or U4307 (N_4307,In_252,In_1742);
or U4308 (N_4308,In_628,In_1886);
nand U4309 (N_4309,In_1277,In_965);
nand U4310 (N_4310,In_1984,In_1287);
nand U4311 (N_4311,In_1549,In_873);
nand U4312 (N_4312,In_481,In_393);
nor U4313 (N_4313,In_1671,In_453);
or U4314 (N_4314,In_1513,In_66);
nor U4315 (N_4315,In_1551,In_1167);
nor U4316 (N_4316,In_1256,In_1610);
and U4317 (N_4317,In_357,In_936);
nor U4318 (N_4318,In_508,In_561);
or U4319 (N_4319,In_711,In_1592);
nand U4320 (N_4320,In_612,In_392);
and U4321 (N_4321,In_1196,In_1400);
nand U4322 (N_4322,In_1902,In_1741);
or U4323 (N_4323,In_1900,In_435);
nor U4324 (N_4324,In_1467,In_1726);
or U4325 (N_4325,In_815,In_163);
nor U4326 (N_4326,In_155,In_1604);
nor U4327 (N_4327,In_1057,In_1511);
or U4328 (N_4328,In_1686,In_1467);
nor U4329 (N_4329,In_652,In_635);
or U4330 (N_4330,In_1457,In_1587);
and U4331 (N_4331,In_1912,In_279);
xnor U4332 (N_4332,In_1215,In_755);
nand U4333 (N_4333,In_1158,In_1756);
nor U4334 (N_4334,In_298,In_240);
nor U4335 (N_4335,In_1120,In_193);
and U4336 (N_4336,In_377,In_292);
nor U4337 (N_4337,In_647,In_931);
or U4338 (N_4338,In_589,In_364);
and U4339 (N_4339,In_1971,In_1772);
nor U4340 (N_4340,In_1418,In_698);
nand U4341 (N_4341,In_1997,In_945);
nand U4342 (N_4342,In_989,In_345);
or U4343 (N_4343,In_534,In_1056);
nor U4344 (N_4344,In_1093,In_1292);
and U4345 (N_4345,In_1088,In_947);
and U4346 (N_4346,In_1683,In_1693);
or U4347 (N_4347,In_433,In_1712);
or U4348 (N_4348,In_304,In_153);
and U4349 (N_4349,In_797,In_1501);
and U4350 (N_4350,In_552,In_930);
or U4351 (N_4351,In_1737,In_1041);
or U4352 (N_4352,In_277,In_495);
xnor U4353 (N_4353,In_801,In_855);
nor U4354 (N_4354,In_1341,In_1802);
nand U4355 (N_4355,In_1080,In_998);
nand U4356 (N_4356,In_1282,In_5);
nor U4357 (N_4357,In_234,In_1589);
or U4358 (N_4358,In_1168,In_1589);
nand U4359 (N_4359,In_1870,In_657);
or U4360 (N_4360,In_170,In_1311);
and U4361 (N_4361,In_1694,In_1907);
and U4362 (N_4362,In_1513,In_321);
nor U4363 (N_4363,In_786,In_1563);
or U4364 (N_4364,In_1248,In_1525);
and U4365 (N_4365,In_912,In_645);
nand U4366 (N_4366,In_601,In_1264);
and U4367 (N_4367,In_1833,In_691);
and U4368 (N_4368,In_1325,In_802);
nand U4369 (N_4369,In_1069,In_1302);
nor U4370 (N_4370,In_1975,In_571);
or U4371 (N_4371,In_1101,In_1325);
nor U4372 (N_4372,In_608,In_1433);
nand U4373 (N_4373,In_124,In_716);
nor U4374 (N_4374,In_328,In_1602);
or U4375 (N_4375,In_1178,In_654);
nor U4376 (N_4376,In_1731,In_1744);
and U4377 (N_4377,In_1960,In_83);
nand U4378 (N_4378,In_1839,In_486);
or U4379 (N_4379,In_415,In_582);
nor U4380 (N_4380,In_948,In_1653);
nand U4381 (N_4381,In_632,In_1368);
nand U4382 (N_4382,In_345,In_1171);
and U4383 (N_4383,In_480,In_1486);
nor U4384 (N_4384,In_676,In_957);
and U4385 (N_4385,In_1758,In_1362);
or U4386 (N_4386,In_1275,In_1038);
and U4387 (N_4387,In_223,In_910);
nand U4388 (N_4388,In_523,In_60);
nor U4389 (N_4389,In_1422,In_277);
or U4390 (N_4390,In_501,In_1399);
nor U4391 (N_4391,In_526,In_1364);
nand U4392 (N_4392,In_305,In_1637);
nor U4393 (N_4393,In_174,In_1065);
nor U4394 (N_4394,In_1921,In_450);
and U4395 (N_4395,In_1670,In_571);
or U4396 (N_4396,In_291,In_652);
nor U4397 (N_4397,In_1273,In_1451);
nand U4398 (N_4398,In_799,In_1578);
and U4399 (N_4399,In_1510,In_1972);
nand U4400 (N_4400,In_1281,In_489);
or U4401 (N_4401,In_517,In_988);
nor U4402 (N_4402,In_1075,In_582);
and U4403 (N_4403,In_640,In_391);
xnor U4404 (N_4404,In_258,In_1219);
and U4405 (N_4405,In_1216,In_99);
nor U4406 (N_4406,In_1681,In_743);
nand U4407 (N_4407,In_1955,In_1229);
nand U4408 (N_4408,In_111,In_1961);
nand U4409 (N_4409,In_1255,In_993);
nand U4410 (N_4410,In_1876,In_192);
nand U4411 (N_4411,In_804,In_1563);
nor U4412 (N_4412,In_1466,In_852);
and U4413 (N_4413,In_878,In_784);
and U4414 (N_4414,In_1128,In_1413);
nand U4415 (N_4415,In_1128,In_885);
xnor U4416 (N_4416,In_608,In_916);
or U4417 (N_4417,In_1678,In_30);
nor U4418 (N_4418,In_999,In_1644);
nor U4419 (N_4419,In_1773,In_188);
and U4420 (N_4420,In_1127,In_1151);
nand U4421 (N_4421,In_1001,In_1743);
or U4422 (N_4422,In_251,In_1756);
or U4423 (N_4423,In_1939,In_900);
or U4424 (N_4424,In_740,In_1514);
or U4425 (N_4425,In_1407,In_1563);
or U4426 (N_4426,In_1109,In_549);
nor U4427 (N_4427,In_1555,In_1784);
nand U4428 (N_4428,In_22,In_819);
nand U4429 (N_4429,In_1317,In_257);
or U4430 (N_4430,In_1339,In_44);
nor U4431 (N_4431,In_162,In_134);
or U4432 (N_4432,In_1033,In_1215);
nand U4433 (N_4433,In_722,In_560);
or U4434 (N_4434,In_106,In_1810);
or U4435 (N_4435,In_262,In_1810);
nand U4436 (N_4436,In_87,In_204);
and U4437 (N_4437,In_1325,In_660);
nor U4438 (N_4438,In_1078,In_1771);
nor U4439 (N_4439,In_1933,In_1182);
and U4440 (N_4440,In_838,In_950);
nor U4441 (N_4441,In_617,In_1031);
or U4442 (N_4442,In_952,In_1035);
nand U4443 (N_4443,In_294,In_383);
or U4444 (N_4444,In_225,In_1446);
and U4445 (N_4445,In_1453,In_698);
nor U4446 (N_4446,In_618,In_688);
nand U4447 (N_4447,In_1909,In_985);
nor U4448 (N_4448,In_710,In_1586);
nor U4449 (N_4449,In_629,In_383);
xor U4450 (N_4450,In_1116,In_1613);
and U4451 (N_4451,In_140,In_646);
nand U4452 (N_4452,In_1206,In_1581);
nand U4453 (N_4453,In_1714,In_640);
nand U4454 (N_4454,In_317,In_1801);
or U4455 (N_4455,In_162,In_1397);
nand U4456 (N_4456,In_50,In_1052);
nand U4457 (N_4457,In_926,In_302);
and U4458 (N_4458,In_1170,In_1130);
or U4459 (N_4459,In_1517,In_264);
and U4460 (N_4460,In_1747,In_172);
nor U4461 (N_4461,In_1373,In_1557);
nor U4462 (N_4462,In_1881,In_566);
nor U4463 (N_4463,In_1978,In_1290);
nand U4464 (N_4464,In_1537,In_1249);
and U4465 (N_4465,In_329,In_811);
and U4466 (N_4466,In_13,In_1365);
nor U4467 (N_4467,In_105,In_1962);
nand U4468 (N_4468,In_1086,In_1838);
nand U4469 (N_4469,In_1989,In_1612);
and U4470 (N_4470,In_1842,In_1794);
nand U4471 (N_4471,In_1600,In_1399);
nor U4472 (N_4472,In_1629,In_798);
nor U4473 (N_4473,In_1690,In_19);
nand U4474 (N_4474,In_1025,In_1477);
nand U4475 (N_4475,In_254,In_1351);
nor U4476 (N_4476,In_1544,In_101);
nand U4477 (N_4477,In_1007,In_133);
nand U4478 (N_4478,In_201,In_600);
nor U4479 (N_4479,In_986,In_1793);
nor U4480 (N_4480,In_272,In_1864);
nand U4481 (N_4481,In_1386,In_1140);
or U4482 (N_4482,In_826,In_1316);
and U4483 (N_4483,In_1700,In_700);
nor U4484 (N_4484,In_186,In_1695);
and U4485 (N_4485,In_1589,In_177);
and U4486 (N_4486,In_270,In_289);
nand U4487 (N_4487,In_818,In_1509);
nor U4488 (N_4488,In_156,In_1050);
and U4489 (N_4489,In_703,In_1826);
nand U4490 (N_4490,In_1769,In_1510);
nor U4491 (N_4491,In_1061,In_603);
or U4492 (N_4492,In_1403,In_1395);
nand U4493 (N_4493,In_1307,In_205);
nor U4494 (N_4494,In_526,In_540);
nor U4495 (N_4495,In_1173,In_751);
or U4496 (N_4496,In_236,In_1909);
nor U4497 (N_4497,In_1439,In_346);
and U4498 (N_4498,In_903,In_840);
nand U4499 (N_4499,In_1454,In_816);
nor U4500 (N_4500,In_387,In_804);
or U4501 (N_4501,In_7,In_247);
xnor U4502 (N_4502,In_999,In_1801);
and U4503 (N_4503,In_913,In_1364);
nand U4504 (N_4504,In_1326,In_578);
and U4505 (N_4505,In_1167,In_1144);
nand U4506 (N_4506,In_720,In_377);
nand U4507 (N_4507,In_1050,In_72);
or U4508 (N_4508,In_1937,In_1633);
and U4509 (N_4509,In_915,In_1116);
nor U4510 (N_4510,In_817,In_149);
nand U4511 (N_4511,In_1321,In_1785);
nand U4512 (N_4512,In_341,In_386);
or U4513 (N_4513,In_100,In_741);
nor U4514 (N_4514,In_1434,In_1328);
nand U4515 (N_4515,In_1453,In_646);
nor U4516 (N_4516,In_537,In_1885);
and U4517 (N_4517,In_435,In_1927);
nor U4518 (N_4518,In_1082,In_915);
or U4519 (N_4519,In_1292,In_753);
or U4520 (N_4520,In_36,In_1708);
nor U4521 (N_4521,In_351,In_1054);
nor U4522 (N_4522,In_1818,In_998);
and U4523 (N_4523,In_376,In_403);
or U4524 (N_4524,In_1377,In_1095);
xor U4525 (N_4525,In_1384,In_64);
and U4526 (N_4526,In_1126,In_101);
nor U4527 (N_4527,In_673,In_1377);
and U4528 (N_4528,In_642,In_1095);
nor U4529 (N_4529,In_252,In_122);
nand U4530 (N_4530,In_732,In_751);
nor U4531 (N_4531,In_1511,In_305);
nor U4532 (N_4532,In_1554,In_781);
nand U4533 (N_4533,In_1164,In_548);
nand U4534 (N_4534,In_15,In_397);
nor U4535 (N_4535,In_1712,In_1916);
nor U4536 (N_4536,In_268,In_432);
and U4537 (N_4537,In_816,In_975);
and U4538 (N_4538,In_1357,In_1355);
nand U4539 (N_4539,In_1833,In_1057);
nand U4540 (N_4540,In_228,In_1183);
and U4541 (N_4541,In_816,In_1130);
and U4542 (N_4542,In_178,In_447);
nor U4543 (N_4543,In_1778,In_8);
and U4544 (N_4544,In_556,In_1217);
nand U4545 (N_4545,In_323,In_1640);
or U4546 (N_4546,In_1125,In_682);
nand U4547 (N_4547,In_931,In_935);
nand U4548 (N_4548,In_19,In_381);
and U4549 (N_4549,In_37,In_701);
and U4550 (N_4550,In_72,In_617);
and U4551 (N_4551,In_1361,In_269);
nand U4552 (N_4552,In_861,In_1141);
nand U4553 (N_4553,In_1259,In_492);
or U4554 (N_4554,In_1939,In_1837);
nand U4555 (N_4555,In_1736,In_637);
and U4556 (N_4556,In_1623,In_279);
or U4557 (N_4557,In_246,In_989);
and U4558 (N_4558,In_649,In_534);
nand U4559 (N_4559,In_1054,In_1559);
xnor U4560 (N_4560,In_1950,In_41);
nor U4561 (N_4561,In_1761,In_1456);
nor U4562 (N_4562,In_1207,In_501);
nand U4563 (N_4563,In_1352,In_1366);
nor U4564 (N_4564,In_156,In_1901);
xnor U4565 (N_4565,In_1507,In_883);
and U4566 (N_4566,In_525,In_79);
and U4567 (N_4567,In_1658,In_377);
nand U4568 (N_4568,In_1749,In_629);
nor U4569 (N_4569,In_1669,In_218);
or U4570 (N_4570,In_350,In_1361);
and U4571 (N_4571,In_724,In_277);
nand U4572 (N_4572,In_1128,In_1997);
nor U4573 (N_4573,In_49,In_1497);
nor U4574 (N_4574,In_864,In_370);
and U4575 (N_4575,In_1070,In_1274);
nor U4576 (N_4576,In_1862,In_685);
nand U4577 (N_4577,In_1092,In_1202);
nand U4578 (N_4578,In_1815,In_685);
and U4579 (N_4579,In_1320,In_40);
or U4580 (N_4580,In_909,In_449);
nor U4581 (N_4581,In_363,In_1662);
or U4582 (N_4582,In_59,In_1109);
nor U4583 (N_4583,In_1532,In_1711);
nand U4584 (N_4584,In_717,In_2);
and U4585 (N_4585,In_1302,In_812);
nor U4586 (N_4586,In_1723,In_405);
nor U4587 (N_4587,In_1375,In_931);
nor U4588 (N_4588,In_718,In_1517);
xnor U4589 (N_4589,In_1683,In_48);
or U4590 (N_4590,In_912,In_84);
or U4591 (N_4591,In_1887,In_1497);
nand U4592 (N_4592,In_885,In_969);
and U4593 (N_4593,In_1706,In_1368);
and U4594 (N_4594,In_319,In_385);
nand U4595 (N_4595,In_1521,In_902);
nor U4596 (N_4596,In_1593,In_1892);
nor U4597 (N_4597,In_1644,In_1690);
nand U4598 (N_4598,In_1563,In_1762);
nor U4599 (N_4599,In_522,In_96);
nand U4600 (N_4600,In_628,In_1305);
nor U4601 (N_4601,In_1446,In_1508);
and U4602 (N_4602,In_1037,In_1597);
nor U4603 (N_4603,In_1448,In_1847);
nor U4604 (N_4604,In_570,In_1135);
nand U4605 (N_4605,In_548,In_1702);
and U4606 (N_4606,In_336,In_1231);
or U4607 (N_4607,In_1981,In_979);
nand U4608 (N_4608,In_1771,In_1562);
nor U4609 (N_4609,In_746,In_919);
and U4610 (N_4610,In_439,In_665);
and U4611 (N_4611,In_636,In_1325);
and U4612 (N_4612,In_52,In_1173);
and U4613 (N_4613,In_507,In_1725);
or U4614 (N_4614,In_1540,In_743);
or U4615 (N_4615,In_1008,In_928);
or U4616 (N_4616,In_1122,In_1422);
nand U4617 (N_4617,In_980,In_1779);
or U4618 (N_4618,In_1786,In_987);
or U4619 (N_4619,In_1161,In_1927);
or U4620 (N_4620,In_1723,In_901);
nor U4621 (N_4621,In_210,In_672);
nor U4622 (N_4622,In_272,In_235);
and U4623 (N_4623,In_1198,In_852);
xnor U4624 (N_4624,In_931,In_1966);
nor U4625 (N_4625,In_898,In_1864);
or U4626 (N_4626,In_228,In_1528);
and U4627 (N_4627,In_152,In_1000);
nand U4628 (N_4628,In_435,In_857);
and U4629 (N_4629,In_1601,In_903);
nand U4630 (N_4630,In_613,In_1656);
or U4631 (N_4631,In_743,In_1805);
or U4632 (N_4632,In_528,In_1835);
nand U4633 (N_4633,In_1366,In_1019);
and U4634 (N_4634,In_1714,In_1604);
nor U4635 (N_4635,In_648,In_1607);
nand U4636 (N_4636,In_1169,In_558);
nor U4637 (N_4637,In_1046,In_708);
or U4638 (N_4638,In_1937,In_1818);
nor U4639 (N_4639,In_899,In_597);
or U4640 (N_4640,In_85,In_1466);
nand U4641 (N_4641,In_1026,In_476);
nand U4642 (N_4642,In_21,In_215);
nand U4643 (N_4643,In_533,In_1904);
and U4644 (N_4644,In_431,In_478);
nand U4645 (N_4645,In_1460,In_1805);
nand U4646 (N_4646,In_40,In_1589);
nor U4647 (N_4647,In_940,In_1381);
or U4648 (N_4648,In_245,In_1161);
nor U4649 (N_4649,In_1340,In_211);
and U4650 (N_4650,In_1099,In_573);
or U4651 (N_4651,In_1313,In_1476);
nor U4652 (N_4652,In_399,In_424);
and U4653 (N_4653,In_1316,In_1261);
and U4654 (N_4654,In_1382,In_536);
or U4655 (N_4655,In_194,In_1692);
or U4656 (N_4656,In_1885,In_1528);
nand U4657 (N_4657,In_1595,In_1610);
nand U4658 (N_4658,In_1372,In_1696);
and U4659 (N_4659,In_114,In_593);
nand U4660 (N_4660,In_954,In_1103);
or U4661 (N_4661,In_1608,In_1133);
and U4662 (N_4662,In_647,In_314);
nor U4663 (N_4663,In_1183,In_737);
and U4664 (N_4664,In_1846,In_1106);
nor U4665 (N_4665,In_283,In_25);
and U4666 (N_4666,In_635,In_1984);
or U4667 (N_4667,In_358,In_80);
nor U4668 (N_4668,In_163,In_3);
nand U4669 (N_4669,In_1088,In_1014);
or U4670 (N_4670,In_507,In_1169);
nor U4671 (N_4671,In_1122,In_1007);
and U4672 (N_4672,In_493,In_549);
or U4673 (N_4673,In_936,In_1909);
and U4674 (N_4674,In_967,In_1405);
nor U4675 (N_4675,In_1697,In_1629);
nor U4676 (N_4676,In_545,In_1311);
nor U4677 (N_4677,In_1458,In_612);
or U4678 (N_4678,In_1325,In_1962);
nor U4679 (N_4679,In_1890,In_932);
and U4680 (N_4680,In_1374,In_1344);
nand U4681 (N_4681,In_1154,In_1208);
and U4682 (N_4682,In_1919,In_1041);
or U4683 (N_4683,In_52,In_166);
nand U4684 (N_4684,In_1529,In_872);
or U4685 (N_4685,In_1897,In_1437);
or U4686 (N_4686,In_1335,In_682);
and U4687 (N_4687,In_891,In_1992);
or U4688 (N_4688,In_715,In_1405);
nand U4689 (N_4689,In_865,In_1815);
nor U4690 (N_4690,In_762,In_1400);
and U4691 (N_4691,In_1279,In_545);
or U4692 (N_4692,In_189,In_1919);
nor U4693 (N_4693,In_1150,In_412);
and U4694 (N_4694,In_238,In_452);
and U4695 (N_4695,In_595,In_856);
nor U4696 (N_4696,In_153,In_723);
nand U4697 (N_4697,In_1988,In_1613);
nand U4698 (N_4698,In_864,In_940);
and U4699 (N_4699,In_141,In_1674);
and U4700 (N_4700,In_665,In_755);
and U4701 (N_4701,In_1322,In_1506);
nand U4702 (N_4702,In_353,In_1879);
and U4703 (N_4703,In_1909,In_1295);
and U4704 (N_4704,In_266,In_125);
nand U4705 (N_4705,In_154,In_1094);
nand U4706 (N_4706,In_1810,In_559);
nor U4707 (N_4707,In_1899,In_1562);
nand U4708 (N_4708,In_1743,In_420);
nand U4709 (N_4709,In_936,In_44);
nor U4710 (N_4710,In_923,In_1063);
or U4711 (N_4711,In_1374,In_1133);
nor U4712 (N_4712,In_168,In_241);
and U4713 (N_4713,In_998,In_196);
and U4714 (N_4714,In_1356,In_1793);
nand U4715 (N_4715,In_1562,In_939);
xnor U4716 (N_4716,In_1925,In_356);
and U4717 (N_4717,In_1727,In_1426);
nand U4718 (N_4718,In_817,In_70);
and U4719 (N_4719,In_117,In_898);
or U4720 (N_4720,In_1256,In_1975);
or U4721 (N_4721,In_224,In_590);
nor U4722 (N_4722,In_1696,In_1418);
or U4723 (N_4723,In_1018,In_1430);
nand U4724 (N_4724,In_1358,In_1542);
nor U4725 (N_4725,In_1721,In_1585);
nand U4726 (N_4726,In_1034,In_1852);
nand U4727 (N_4727,In_253,In_1161);
or U4728 (N_4728,In_879,In_1612);
or U4729 (N_4729,In_775,In_1009);
nand U4730 (N_4730,In_1643,In_64);
nand U4731 (N_4731,In_736,In_154);
or U4732 (N_4732,In_287,In_1081);
nor U4733 (N_4733,In_1406,In_777);
or U4734 (N_4734,In_766,In_1931);
or U4735 (N_4735,In_1489,In_15);
nor U4736 (N_4736,In_1622,In_50);
nand U4737 (N_4737,In_1424,In_975);
and U4738 (N_4738,In_1395,In_1378);
nor U4739 (N_4739,In_969,In_813);
nor U4740 (N_4740,In_938,In_121);
or U4741 (N_4741,In_1705,In_1184);
nand U4742 (N_4742,In_619,In_1970);
nand U4743 (N_4743,In_1997,In_1151);
or U4744 (N_4744,In_638,In_494);
or U4745 (N_4745,In_1492,In_1778);
nor U4746 (N_4746,In_1284,In_1796);
or U4747 (N_4747,In_48,In_1641);
nand U4748 (N_4748,In_102,In_479);
nand U4749 (N_4749,In_471,In_842);
and U4750 (N_4750,In_324,In_187);
and U4751 (N_4751,In_90,In_1009);
nor U4752 (N_4752,In_490,In_65);
nor U4753 (N_4753,In_877,In_956);
and U4754 (N_4754,In_1892,In_654);
and U4755 (N_4755,In_83,In_1524);
and U4756 (N_4756,In_1351,In_870);
xnor U4757 (N_4757,In_1851,In_53);
or U4758 (N_4758,In_144,In_925);
nand U4759 (N_4759,In_357,In_1773);
nand U4760 (N_4760,In_455,In_141);
nand U4761 (N_4761,In_1884,In_1989);
or U4762 (N_4762,In_991,In_1633);
nand U4763 (N_4763,In_1521,In_1611);
or U4764 (N_4764,In_1732,In_1312);
nor U4765 (N_4765,In_761,In_121);
nor U4766 (N_4766,In_1029,In_821);
or U4767 (N_4767,In_1544,In_123);
or U4768 (N_4768,In_669,In_1328);
and U4769 (N_4769,In_1306,In_1132);
or U4770 (N_4770,In_275,In_969);
nand U4771 (N_4771,In_348,In_1257);
nor U4772 (N_4772,In_157,In_1225);
nand U4773 (N_4773,In_94,In_740);
nand U4774 (N_4774,In_1320,In_1682);
and U4775 (N_4775,In_2,In_1962);
nand U4776 (N_4776,In_135,In_1680);
nand U4777 (N_4777,In_1381,In_1511);
nor U4778 (N_4778,In_1422,In_48);
nor U4779 (N_4779,In_915,In_210);
nor U4780 (N_4780,In_783,In_1008);
and U4781 (N_4781,In_344,In_1032);
nand U4782 (N_4782,In_1541,In_1757);
and U4783 (N_4783,In_662,In_1319);
xor U4784 (N_4784,In_1835,In_1851);
and U4785 (N_4785,In_1364,In_408);
or U4786 (N_4786,In_387,In_36);
or U4787 (N_4787,In_1050,In_1435);
nand U4788 (N_4788,In_1094,In_925);
nor U4789 (N_4789,In_1148,In_1921);
nor U4790 (N_4790,In_1465,In_1986);
nor U4791 (N_4791,In_924,In_1802);
nand U4792 (N_4792,In_1092,In_1680);
and U4793 (N_4793,In_1568,In_1866);
or U4794 (N_4794,In_575,In_554);
nor U4795 (N_4795,In_461,In_503);
nand U4796 (N_4796,In_670,In_393);
or U4797 (N_4797,In_519,In_751);
nand U4798 (N_4798,In_4,In_1069);
nor U4799 (N_4799,In_4,In_233);
or U4800 (N_4800,In_965,In_839);
or U4801 (N_4801,In_790,In_753);
nor U4802 (N_4802,In_1640,In_580);
and U4803 (N_4803,In_1962,In_1968);
nand U4804 (N_4804,In_747,In_456);
or U4805 (N_4805,In_1236,In_242);
nor U4806 (N_4806,In_1662,In_1542);
and U4807 (N_4807,In_420,In_428);
or U4808 (N_4808,In_1941,In_821);
nand U4809 (N_4809,In_1348,In_1261);
nor U4810 (N_4810,In_1863,In_1143);
or U4811 (N_4811,In_131,In_1948);
nand U4812 (N_4812,In_1158,In_97);
or U4813 (N_4813,In_1773,In_1048);
nor U4814 (N_4814,In_376,In_1154);
or U4815 (N_4815,In_980,In_61);
and U4816 (N_4816,In_497,In_1695);
and U4817 (N_4817,In_1308,In_405);
nor U4818 (N_4818,In_257,In_974);
nand U4819 (N_4819,In_1288,In_410);
and U4820 (N_4820,In_264,In_47);
or U4821 (N_4821,In_44,In_366);
nor U4822 (N_4822,In_1994,In_496);
xor U4823 (N_4823,In_1186,In_316);
and U4824 (N_4824,In_572,In_141);
nand U4825 (N_4825,In_1366,In_1591);
nor U4826 (N_4826,In_619,In_1471);
nand U4827 (N_4827,In_1963,In_93);
or U4828 (N_4828,In_344,In_1022);
nand U4829 (N_4829,In_1324,In_1096);
xnor U4830 (N_4830,In_1925,In_900);
nand U4831 (N_4831,In_1090,In_1371);
nor U4832 (N_4832,In_1844,In_1296);
or U4833 (N_4833,In_1411,In_1918);
nor U4834 (N_4834,In_1248,In_156);
nor U4835 (N_4835,In_442,In_1140);
and U4836 (N_4836,In_90,In_604);
nor U4837 (N_4837,In_1263,In_52);
nor U4838 (N_4838,In_1704,In_466);
nor U4839 (N_4839,In_38,In_1847);
or U4840 (N_4840,In_101,In_1078);
nand U4841 (N_4841,In_989,In_1247);
nand U4842 (N_4842,In_1910,In_1859);
nor U4843 (N_4843,In_1802,In_1909);
nand U4844 (N_4844,In_1643,In_1480);
nor U4845 (N_4845,In_425,In_1003);
or U4846 (N_4846,In_1530,In_459);
nor U4847 (N_4847,In_1303,In_72);
nand U4848 (N_4848,In_375,In_1734);
nor U4849 (N_4849,In_1632,In_874);
or U4850 (N_4850,In_1681,In_1796);
nand U4851 (N_4851,In_295,In_822);
and U4852 (N_4852,In_460,In_1071);
and U4853 (N_4853,In_443,In_847);
nand U4854 (N_4854,In_1106,In_1747);
and U4855 (N_4855,In_1907,In_535);
or U4856 (N_4856,In_1022,In_260);
nor U4857 (N_4857,In_347,In_1888);
nor U4858 (N_4858,In_141,In_1363);
and U4859 (N_4859,In_862,In_1094);
or U4860 (N_4860,In_108,In_425);
or U4861 (N_4861,In_820,In_1020);
or U4862 (N_4862,In_1391,In_1129);
or U4863 (N_4863,In_1528,In_225);
nand U4864 (N_4864,In_292,In_533);
nand U4865 (N_4865,In_117,In_753);
and U4866 (N_4866,In_1172,In_463);
nand U4867 (N_4867,In_1033,In_501);
or U4868 (N_4868,In_1835,In_1745);
nor U4869 (N_4869,In_316,In_464);
or U4870 (N_4870,In_1033,In_476);
nor U4871 (N_4871,In_1443,In_1409);
nand U4872 (N_4872,In_460,In_761);
nor U4873 (N_4873,In_1894,In_73);
nor U4874 (N_4874,In_368,In_270);
or U4875 (N_4875,In_1863,In_1927);
nand U4876 (N_4876,In_1386,In_1499);
nand U4877 (N_4877,In_452,In_993);
or U4878 (N_4878,In_745,In_608);
nand U4879 (N_4879,In_1342,In_1360);
or U4880 (N_4880,In_145,In_40);
and U4881 (N_4881,In_1023,In_1260);
nand U4882 (N_4882,In_514,In_868);
or U4883 (N_4883,In_806,In_245);
xor U4884 (N_4884,In_1877,In_805);
nand U4885 (N_4885,In_1524,In_779);
nand U4886 (N_4886,In_1874,In_870);
and U4887 (N_4887,In_1104,In_1239);
or U4888 (N_4888,In_1467,In_176);
or U4889 (N_4889,In_924,In_1948);
xor U4890 (N_4890,In_690,In_486);
and U4891 (N_4891,In_782,In_130);
nand U4892 (N_4892,In_938,In_724);
or U4893 (N_4893,In_1480,In_1306);
or U4894 (N_4894,In_1346,In_1463);
and U4895 (N_4895,In_105,In_940);
nand U4896 (N_4896,In_1156,In_718);
nand U4897 (N_4897,In_1660,In_946);
or U4898 (N_4898,In_1272,In_1009);
and U4899 (N_4899,In_973,In_594);
nor U4900 (N_4900,In_1076,In_1936);
nor U4901 (N_4901,In_885,In_1711);
and U4902 (N_4902,In_1849,In_7);
nand U4903 (N_4903,In_122,In_683);
nand U4904 (N_4904,In_1299,In_1519);
or U4905 (N_4905,In_1012,In_848);
or U4906 (N_4906,In_1567,In_98);
nand U4907 (N_4907,In_325,In_214);
nor U4908 (N_4908,In_1184,In_170);
nor U4909 (N_4909,In_362,In_1189);
nand U4910 (N_4910,In_275,In_1496);
and U4911 (N_4911,In_1114,In_784);
and U4912 (N_4912,In_349,In_416);
nand U4913 (N_4913,In_400,In_1074);
and U4914 (N_4914,In_1817,In_1213);
and U4915 (N_4915,In_801,In_1772);
nor U4916 (N_4916,In_1149,In_1699);
nand U4917 (N_4917,In_643,In_1044);
nor U4918 (N_4918,In_1866,In_608);
nand U4919 (N_4919,In_1130,In_356);
nor U4920 (N_4920,In_1005,In_1063);
or U4921 (N_4921,In_1662,In_36);
or U4922 (N_4922,In_407,In_635);
and U4923 (N_4923,In_1835,In_1161);
and U4924 (N_4924,In_205,In_426);
or U4925 (N_4925,In_1959,In_423);
or U4926 (N_4926,In_618,In_1552);
nand U4927 (N_4927,In_549,In_913);
nor U4928 (N_4928,In_1062,In_1724);
or U4929 (N_4929,In_185,In_1928);
nor U4930 (N_4930,In_1908,In_1855);
nor U4931 (N_4931,In_331,In_1338);
or U4932 (N_4932,In_1858,In_97);
nand U4933 (N_4933,In_367,In_1);
and U4934 (N_4934,In_422,In_1724);
nand U4935 (N_4935,In_990,In_1712);
nand U4936 (N_4936,In_515,In_1956);
xor U4937 (N_4937,In_258,In_1088);
nand U4938 (N_4938,In_1413,In_1022);
nand U4939 (N_4939,In_325,In_516);
or U4940 (N_4940,In_312,In_1757);
nor U4941 (N_4941,In_1399,In_837);
or U4942 (N_4942,In_1506,In_1087);
or U4943 (N_4943,In_513,In_688);
nand U4944 (N_4944,In_591,In_600);
or U4945 (N_4945,In_1873,In_1751);
nand U4946 (N_4946,In_1216,In_1522);
or U4947 (N_4947,In_1656,In_604);
nor U4948 (N_4948,In_1267,In_4);
nand U4949 (N_4949,In_388,In_537);
or U4950 (N_4950,In_120,In_450);
or U4951 (N_4951,In_248,In_1950);
and U4952 (N_4952,In_1770,In_1267);
nor U4953 (N_4953,In_1295,In_1151);
and U4954 (N_4954,In_815,In_449);
nand U4955 (N_4955,In_756,In_1449);
nand U4956 (N_4956,In_1977,In_628);
and U4957 (N_4957,In_1488,In_1293);
nand U4958 (N_4958,In_809,In_121);
and U4959 (N_4959,In_81,In_1279);
and U4960 (N_4960,In_590,In_319);
and U4961 (N_4961,In_284,In_67);
or U4962 (N_4962,In_1852,In_1323);
nand U4963 (N_4963,In_1498,In_1772);
and U4964 (N_4964,In_835,In_719);
xnor U4965 (N_4965,In_480,In_1305);
nand U4966 (N_4966,In_1887,In_907);
nand U4967 (N_4967,In_1522,In_1371);
and U4968 (N_4968,In_142,In_1966);
nor U4969 (N_4969,In_1754,In_964);
and U4970 (N_4970,In_1546,In_1397);
or U4971 (N_4971,In_360,In_149);
nand U4972 (N_4972,In_1102,In_438);
or U4973 (N_4973,In_351,In_1822);
and U4974 (N_4974,In_835,In_659);
and U4975 (N_4975,In_1898,In_1213);
or U4976 (N_4976,In_211,In_736);
nand U4977 (N_4977,In_872,In_1764);
nand U4978 (N_4978,In_264,In_933);
and U4979 (N_4979,In_479,In_1594);
or U4980 (N_4980,In_1499,In_1756);
and U4981 (N_4981,In_1678,In_1024);
nor U4982 (N_4982,In_454,In_371);
nand U4983 (N_4983,In_1016,In_305);
or U4984 (N_4984,In_125,In_1148);
and U4985 (N_4985,In_143,In_392);
nand U4986 (N_4986,In_1435,In_1018);
and U4987 (N_4987,In_1292,In_592);
nand U4988 (N_4988,In_825,In_1898);
or U4989 (N_4989,In_798,In_307);
and U4990 (N_4990,In_1800,In_942);
nand U4991 (N_4991,In_1914,In_423);
nor U4992 (N_4992,In_866,In_1307);
nor U4993 (N_4993,In_134,In_17);
nand U4994 (N_4994,In_1883,In_337);
or U4995 (N_4995,In_216,In_1661);
and U4996 (N_4996,In_1896,In_1992);
nand U4997 (N_4997,In_759,In_1310);
nand U4998 (N_4998,In_1248,In_1377);
and U4999 (N_4999,In_1541,In_195);
or U5000 (N_5000,N_2858,N_2685);
nor U5001 (N_5001,N_897,N_911);
nor U5002 (N_5002,N_4400,N_4805);
nand U5003 (N_5003,N_2125,N_1972);
nand U5004 (N_5004,N_137,N_2051);
and U5005 (N_5005,N_3302,N_1369);
or U5006 (N_5006,N_1412,N_622);
and U5007 (N_5007,N_4962,N_4316);
nor U5008 (N_5008,N_3178,N_1415);
or U5009 (N_5009,N_4835,N_712);
nand U5010 (N_5010,N_2162,N_853);
xnor U5011 (N_5011,N_733,N_1480);
nor U5012 (N_5012,N_2460,N_2718);
or U5013 (N_5013,N_3914,N_1327);
nand U5014 (N_5014,N_1657,N_2534);
nor U5015 (N_5015,N_3964,N_2152);
and U5016 (N_5016,N_1940,N_4601);
nor U5017 (N_5017,N_2937,N_1650);
and U5018 (N_5018,N_486,N_820);
or U5019 (N_5019,N_2184,N_402);
and U5020 (N_5020,N_2489,N_3069);
nor U5021 (N_5021,N_1803,N_1547);
nand U5022 (N_5022,N_1594,N_2900);
or U5023 (N_5023,N_3037,N_4153);
or U5024 (N_5024,N_3473,N_1132);
and U5025 (N_5025,N_2958,N_2969);
nor U5026 (N_5026,N_3440,N_210);
nor U5027 (N_5027,N_2077,N_4480);
or U5028 (N_5028,N_1147,N_3714);
nor U5029 (N_5029,N_2486,N_1507);
nor U5030 (N_5030,N_89,N_1346);
nand U5031 (N_5031,N_2786,N_2113);
nand U5032 (N_5032,N_3033,N_4483);
and U5033 (N_5033,N_4969,N_3472);
nor U5034 (N_5034,N_3906,N_47);
nor U5035 (N_5035,N_3375,N_334);
nand U5036 (N_5036,N_1521,N_381);
nand U5037 (N_5037,N_4172,N_466);
and U5038 (N_5038,N_817,N_2879);
nand U5039 (N_5039,N_1334,N_4113);
and U5040 (N_5040,N_2740,N_2285);
nand U5041 (N_5041,N_3333,N_2748);
nand U5042 (N_5042,N_3727,N_3471);
or U5043 (N_5043,N_2003,N_3595);
and U5044 (N_5044,N_1637,N_3656);
or U5045 (N_5045,N_3229,N_2765);
nor U5046 (N_5046,N_2790,N_35);
nor U5047 (N_5047,N_2211,N_452);
nand U5048 (N_5048,N_2716,N_3636);
or U5049 (N_5049,N_3266,N_1220);
xnor U5050 (N_5050,N_2216,N_1638);
nand U5051 (N_5051,N_4277,N_326);
and U5052 (N_5052,N_4292,N_575);
and U5053 (N_5053,N_2672,N_131);
or U5054 (N_5054,N_1506,N_3316);
nor U5055 (N_5055,N_2278,N_3516);
nor U5056 (N_5056,N_501,N_2274);
or U5057 (N_5057,N_3548,N_4629);
or U5058 (N_5058,N_4798,N_4789);
and U5059 (N_5059,N_2381,N_1783);
nand U5060 (N_5060,N_147,N_3131);
or U5061 (N_5061,N_678,N_2139);
and U5062 (N_5062,N_2866,N_2940);
or U5063 (N_5063,N_2532,N_2126);
nand U5064 (N_5064,N_4406,N_4708);
and U5065 (N_5065,N_2608,N_1781);
and U5066 (N_5066,N_4306,N_4010);
nand U5067 (N_5067,N_3115,N_3317);
or U5068 (N_5068,N_1873,N_73);
or U5069 (N_5069,N_1761,N_2140);
nor U5070 (N_5070,N_2804,N_4122);
nand U5071 (N_5071,N_2794,N_976);
and U5072 (N_5072,N_2288,N_3557);
nor U5073 (N_5073,N_959,N_4848);
or U5074 (N_5074,N_3759,N_1678);
or U5075 (N_5075,N_367,N_256);
and U5076 (N_5076,N_311,N_99);
nand U5077 (N_5077,N_2237,N_2040);
nor U5078 (N_5078,N_2757,N_4164);
and U5079 (N_5079,N_1896,N_3721);
nand U5080 (N_5080,N_2268,N_4834);
nand U5081 (N_5081,N_1510,N_1798);
or U5082 (N_5082,N_1936,N_2731);
or U5083 (N_5083,N_142,N_3612);
and U5084 (N_5084,N_384,N_3735);
and U5085 (N_5085,N_961,N_3629);
or U5086 (N_5086,N_996,N_1171);
nor U5087 (N_5087,N_1123,N_2895);
nand U5088 (N_5088,N_4575,N_3467);
nand U5089 (N_5089,N_1977,N_3364);
nand U5090 (N_5090,N_282,N_3796);
nand U5091 (N_5091,N_2719,N_615);
nor U5092 (N_5092,N_1116,N_1205);
or U5093 (N_5093,N_139,N_2433);
xor U5094 (N_5094,N_3801,N_4822);
or U5095 (N_5095,N_4856,N_1701);
or U5096 (N_5096,N_4026,N_1540);
and U5097 (N_5097,N_2807,N_4654);
xnor U5098 (N_5098,N_3954,N_163);
nand U5099 (N_5099,N_3483,N_2362);
and U5100 (N_5100,N_3263,N_4594);
or U5101 (N_5101,N_4377,N_986);
or U5102 (N_5102,N_4180,N_444);
and U5103 (N_5103,N_1963,N_1582);
and U5104 (N_5104,N_4154,N_3663);
nand U5105 (N_5105,N_1859,N_3855);
nand U5106 (N_5106,N_2739,N_1418);
nand U5107 (N_5107,N_4426,N_473);
and U5108 (N_5108,N_859,N_4478);
nand U5109 (N_5109,N_4661,N_2800);
and U5110 (N_5110,N_4497,N_1734);
nor U5111 (N_5111,N_3840,N_3336);
nand U5112 (N_5112,N_4887,N_2842);
nor U5113 (N_5113,N_2476,N_1067);
and U5114 (N_5114,N_3904,N_4281);
nand U5115 (N_5115,N_574,N_3705);
nand U5116 (N_5116,N_4726,N_4949);
nand U5117 (N_5117,N_2621,N_644);
nor U5118 (N_5118,N_3039,N_492);
and U5119 (N_5119,N_1693,N_1219);
nor U5120 (N_5120,N_924,N_2744);
or U5121 (N_5121,N_2981,N_1679);
or U5122 (N_5122,N_3099,N_4626);
or U5123 (N_5123,N_5,N_3508);
nand U5124 (N_5124,N_3081,N_4101);
and U5125 (N_5125,N_2217,N_2523);
nor U5126 (N_5126,N_3752,N_1771);
and U5127 (N_5127,N_2029,N_2324);
or U5128 (N_5128,N_3746,N_3551);
xor U5129 (N_5129,N_18,N_2674);
and U5130 (N_5130,N_2049,N_2267);
nand U5131 (N_5131,N_1293,N_3095);
and U5132 (N_5132,N_4937,N_1494);
nand U5133 (N_5133,N_2984,N_389);
nand U5134 (N_5134,N_1773,N_667);
nor U5135 (N_5135,N_4695,N_2552);
or U5136 (N_5136,N_4772,N_2463);
and U5137 (N_5137,N_3560,N_1643);
nor U5138 (N_5138,N_3292,N_1986);
or U5139 (N_5139,N_705,N_4442);
or U5140 (N_5140,N_4673,N_2458);
and U5141 (N_5141,N_3521,N_1230);
nor U5142 (N_5142,N_23,N_320);
nor U5143 (N_5143,N_2510,N_446);
nor U5144 (N_5144,N_2776,N_3432);
and U5145 (N_5145,N_4585,N_86);
and U5146 (N_5146,N_3005,N_790);
nand U5147 (N_5147,N_1862,N_539);
or U5148 (N_5148,N_4552,N_3831);
nor U5149 (N_5149,N_222,N_4947);
nand U5150 (N_5150,N_225,N_2974);
and U5151 (N_5151,N_3638,N_3146);
and U5152 (N_5152,N_2747,N_1534);
nand U5153 (N_5153,N_2105,N_1910);
nand U5154 (N_5154,N_406,N_1146);
or U5155 (N_5155,N_2714,N_3662);
nand U5156 (N_5156,N_4034,N_4779);
nand U5157 (N_5157,N_2814,N_3541);
nand U5158 (N_5158,N_1424,N_1367);
xor U5159 (N_5159,N_844,N_2189);
or U5160 (N_5160,N_3041,N_3997);
nor U5161 (N_5161,N_2686,N_260);
and U5162 (N_5162,N_115,N_4989);
or U5163 (N_5163,N_3108,N_1307);
or U5164 (N_5164,N_1348,N_4469);
or U5165 (N_5165,N_3715,N_3057);
or U5166 (N_5166,N_1635,N_2212);
or U5167 (N_5167,N_723,N_4749);
or U5168 (N_5168,N_2064,N_4495);
or U5169 (N_5169,N_360,N_2684);
xnor U5170 (N_5170,N_2665,N_520);
and U5171 (N_5171,N_1530,N_3635);
or U5172 (N_5172,N_4405,N_4028);
and U5173 (N_5173,N_827,N_4500);
nand U5174 (N_5174,N_743,N_93);
nor U5175 (N_5175,N_631,N_4268);
nor U5176 (N_5176,N_2408,N_3280);
nor U5177 (N_5177,N_3815,N_3777);
and U5178 (N_5178,N_487,N_1462);
or U5179 (N_5179,N_1057,N_3382);
or U5180 (N_5180,N_1273,N_1713);
nand U5181 (N_5181,N_3968,N_2559);
or U5182 (N_5182,N_2202,N_209);
and U5183 (N_5183,N_2293,N_1448);
nor U5184 (N_5184,N_2963,N_1772);
or U5185 (N_5185,N_3224,N_3117);
nor U5186 (N_5186,N_2312,N_217);
nor U5187 (N_5187,N_3052,N_2956);
or U5188 (N_5188,N_786,N_1290);
or U5189 (N_5189,N_2075,N_3460);
nor U5190 (N_5190,N_1471,N_1013);
and U5191 (N_5191,N_842,N_3545);
and U5192 (N_5192,N_4525,N_4985);
and U5193 (N_5193,N_4819,N_938);
and U5194 (N_5194,N_268,N_788);
or U5195 (N_5195,N_3434,N_4423);
nand U5196 (N_5196,N_2543,N_259);
xnor U5197 (N_5197,N_1899,N_981);
xor U5198 (N_5198,N_3335,N_1680);
and U5199 (N_5199,N_410,N_3667);
nor U5200 (N_5200,N_1019,N_2473);
xor U5201 (N_5201,N_2390,N_4678);
and U5202 (N_5202,N_2972,N_3343);
and U5203 (N_5203,N_2085,N_253);
and U5204 (N_5204,N_1355,N_1129);
xor U5205 (N_5205,N_3799,N_4724);
nor U5206 (N_5206,N_2167,N_877);
nand U5207 (N_5207,N_3781,N_3249);
and U5208 (N_5208,N_2385,N_4986);
or U5209 (N_5209,N_2478,N_2525);
and U5210 (N_5210,N_4355,N_3067);
nor U5211 (N_5211,N_674,N_2999);
nor U5212 (N_5212,N_1338,N_577);
nor U5213 (N_5213,N_4078,N_799);
nand U5214 (N_5214,N_508,N_1074);
nand U5215 (N_5215,N_2834,N_3744);
or U5216 (N_5216,N_2986,N_2041);
and U5217 (N_5217,N_2816,N_1632);
nor U5218 (N_5218,N_3451,N_4606);
or U5219 (N_5219,N_887,N_2774);
and U5220 (N_5220,N_3643,N_3911);
nor U5221 (N_5221,N_2613,N_2423);
nand U5222 (N_5222,N_4057,N_557);
or U5223 (N_5223,N_1554,N_3262);
xnor U5224 (N_5224,N_2181,N_3969);
nand U5225 (N_5225,N_822,N_2634);
and U5226 (N_5226,N_72,N_4275);
or U5227 (N_5227,N_2912,N_3826);
and U5228 (N_5228,N_413,N_1105);
nor U5229 (N_5229,N_971,N_2676);
nor U5230 (N_5230,N_67,N_2018);
xnor U5231 (N_5231,N_1216,N_4462);
nand U5232 (N_5232,N_3361,N_4156);
nand U5233 (N_5233,N_3481,N_1989);
nand U5234 (N_5234,N_4252,N_105);
nand U5235 (N_5235,N_2365,N_927);
nand U5236 (N_5236,N_3524,N_4928);
and U5237 (N_5237,N_3120,N_4501);
nand U5238 (N_5238,N_1177,N_541);
and U5239 (N_5239,N_4251,N_4563);
nand U5240 (N_5240,N_4553,N_4639);
xor U5241 (N_5241,N_2661,N_368);
nand U5242 (N_5242,N_3258,N_2507);
nor U5243 (N_5243,N_2277,N_1141);
nor U5244 (N_5244,N_3967,N_1770);
and U5245 (N_5245,N_3765,N_547);
nor U5246 (N_5246,N_4382,N_3942);
nand U5247 (N_5247,N_3998,N_3231);
nor U5248 (N_5248,N_3975,N_1890);
or U5249 (N_5249,N_1204,N_2841);
and U5250 (N_5250,N_3561,N_3384);
xor U5251 (N_5251,N_2705,N_1207);
nand U5252 (N_5252,N_3431,N_1006);
nor U5253 (N_5253,N_1416,N_1302);
or U5254 (N_5254,N_1201,N_169);
nand U5255 (N_5255,N_3737,N_2763);
or U5256 (N_5256,N_4123,N_2080);
nand U5257 (N_5257,N_1702,N_4735);
nand U5258 (N_5258,N_1505,N_1523);
nand U5259 (N_5259,N_1549,N_2646);
nand U5260 (N_5260,N_1401,N_1258);
or U5261 (N_5261,N_4351,N_4301);
or U5262 (N_5262,N_4318,N_3490);
nor U5263 (N_5263,N_629,N_1064);
and U5264 (N_5264,N_1945,N_4412);
xor U5265 (N_5265,N_2086,N_2625);
nor U5266 (N_5266,N_1345,N_665);
nor U5267 (N_5267,N_4846,N_862);
nor U5268 (N_5268,N_3778,N_4658);
nand U5269 (N_5269,N_2222,N_4033);
nand U5270 (N_5270,N_1848,N_2773);
or U5271 (N_5271,N_4430,N_2449);
nor U5272 (N_5272,N_400,N_1498);
nor U5273 (N_5273,N_1502,N_2944);
nand U5274 (N_5274,N_4266,N_3747);
and U5275 (N_5275,N_2750,N_4983);
or U5276 (N_5276,N_3695,N_2038);
or U5277 (N_5277,N_4754,N_4234);
and U5278 (N_5278,N_4904,N_735);
nand U5279 (N_5279,N_2901,N_2770);
nand U5280 (N_5280,N_2553,N_694);
nand U5281 (N_5281,N_1911,N_1280);
and U5282 (N_5282,N_3182,N_526);
nand U5283 (N_5283,N_4721,N_3456);
nand U5284 (N_5284,N_3754,N_478);
nand U5285 (N_5285,N_3710,N_946);
or U5286 (N_5286,N_4013,N_2659);
and U5287 (N_5287,N_3520,N_4918);
and U5288 (N_5288,N_2624,N_1532);
and U5289 (N_5289,N_1585,N_3062);
and U5290 (N_5290,N_3716,N_2562);
or U5291 (N_5291,N_2154,N_4143);
nand U5292 (N_5292,N_1755,N_3502);
nor U5293 (N_5293,N_4433,N_2952);
nand U5294 (N_5294,N_2451,N_3681);
or U5295 (N_5295,N_3809,N_4702);
or U5296 (N_5296,N_3122,N_2567);
nand U5297 (N_5297,N_2376,N_4207);
and U5298 (N_5298,N_1126,N_4372);
nor U5299 (N_5299,N_4560,N_1186);
nor U5300 (N_5300,N_900,N_1908);
and U5301 (N_5301,N_1829,N_2782);
and U5302 (N_5302,N_2078,N_2788);
nor U5303 (N_5303,N_3406,N_2370);
and U5304 (N_5304,N_757,N_593);
nand U5305 (N_5305,N_4006,N_2355);
and U5306 (N_5306,N_669,N_995);
nand U5307 (N_5307,N_1144,N_695);
nand U5308 (N_5308,N_2467,N_417);
nor U5309 (N_5309,N_4631,N_1703);
or U5310 (N_5310,N_1932,N_1659);
nor U5311 (N_5311,N_278,N_1618);
or U5312 (N_5312,N_947,N_1305);
nand U5313 (N_5313,N_4079,N_3386);
or U5314 (N_5314,N_2880,N_1974);
nand U5315 (N_5315,N_4707,N_4539);
nor U5316 (N_5316,N_3301,N_1551);
nand U5317 (N_5317,N_453,N_3620);
nand U5318 (N_5318,N_2039,N_218);
or U5319 (N_5319,N_2910,N_39);
xnor U5320 (N_5320,N_34,N_1634);
and U5321 (N_5321,N_2928,N_2276);
nand U5322 (N_5322,N_3112,N_2128);
or U5323 (N_5323,N_1891,N_1166);
and U5324 (N_5324,N_1970,N_162);
nand U5325 (N_5325,N_3870,N_3366);
xor U5326 (N_5326,N_4841,N_3800);
nand U5327 (N_5327,N_4692,N_1208);
or U5328 (N_5328,N_3953,N_2334);
nor U5329 (N_5329,N_2652,N_1744);
nand U5330 (N_5330,N_3443,N_4868);
nor U5331 (N_5331,N_3402,N_4948);
nand U5332 (N_5332,N_2230,N_302);
or U5333 (N_5333,N_4617,N_2208);
nand U5334 (N_5334,N_4700,N_3334);
nor U5335 (N_5335,N_3246,N_3797);
or U5336 (N_5336,N_3938,N_1259);
or U5337 (N_5337,N_1452,N_3477);
nand U5338 (N_5338,N_2374,N_2005);
nor U5339 (N_5339,N_1094,N_2469);
nand U5340 (N_5340,N_1020,N_3532);
or U5341 (N_5341,N_4460,N_2261);
nand U5342 (N_5342,N_2030,N_4806);
or U5343 (N_5343,N_4977,N_2045);
and U5344 (N_5344,N_860,N_1636);
xnor U5345 (N_5345,N_2443,N_1825);
nor U5346 (N_5346,N_237,N_327);
nor U5347 (N_5347,N_425,N_488);
and U5348 (N_5348,N_1847,N_823);
nand U5349 (N_5349,N_1410,N_3875);
nor U5350 (N_5350,N_4745,N_1886);
and U5351 (N_5351,N_3369,N_412);
nand U5352 (N_5352,N_934,N_1603);
nand U5353 (N_5353,N_907,N_4035);
nand U5354 (N_5354,N_298,N_4104);
nand U5355 (N_5355,N_397,N_2820);
and U5356 (N_5356,N_4857,N_4581);
nand U5357 (N_5357,N_506,N_3771);
nand U5358 (N_5358,N_286,N_1919);
nand U5359 (N_5359,N_1090,N_1271);
or U5360 (N_5360,N_2915,N_3485);
and U5361 (N_5361,N_3841,N_3603);
nor U5362 (N_5362,N_831,N_2417);
nor U5363 (N_5363,N_4727,N_3926);
nor U5364 (N_5364,N_829,N_1739);
nor U5365 (N_5365,N_4227,N_528);
and U5366 (N_5366,N_305,N_1159);
nand U5367 (N_5367,N_4701,N_1255);
nand U5368 (N_5368,N_2123,N_2456);
nand U5369 (N_5369,N_3675,N_2190);
nand U5370 (N_5370,N_1654,N_977);
and U5371 (N_5371,N_2514,N_1473);
nand U5372 (N_5372,N_3090,N_2074);
nand U5373 (N_5373,N_3785,N_3252);
nor U5374 (N_5374,N_1430,N_52);
and U5375 (N_5375,N_4386,N_1902);
nand U5376 (N_5376,N_4213,N_3021);
nor U5377 (N_5377,N_888,N_10);
nor U5378 (N_5378,N_4816,N_2207);
nor U5379 (N_5379,N_1962,N_990);
or U5380 (N_5380,N_1938,N_3355);
and U5381 (N_5381,N_3750,N_4349);
and U5382 (N_5382,N_1628,N_3708);
xnor U5383 (N_5383,N_180,N_2031);
and U5384 (N_5384,N_3275,N_879);
nor U5385 (N_5385,N_2752,N_3559);
or U5386 (N_5386,N_81,N_3614);
and U5387 (N_5387,N_1438,N_161);
or U5388 (N_5388,N_857,N_4087);
nand U5389 (N_5389,N_4394,N_2540);
nand U5390 (N_5390,N_1252,N_457);
or U5391 (N_5391,N_1782,N_3948);
nor U5392 (N_5392,N_2699,N_1368);
and U5393 (N_5393,N_2819,N_1969);
nand U5394 (N_5394,N_3944,N_3528);
nand U5395 (N_5395,N_689,N_2439);
nand U5396 (N_5396,N_1880,N_3136);
nand U5397 (N_5397,N_1573,N_4981);
and U5398 (N_5398,N_2822,N_725);
and U5399 (N_5399,N_2353,N_2294);
and U5400 (N_5400,N_3396,N_4831);
xor U5401 (N_5401,N_1061,N_3839);
and U5402 (N_5402,N_2890,N_1040);
and U5403 (N_5403,N_3915,N_1762);
nor U5404 (N_5404,N_3522,N_471);
or U5405 (N_5405,N_4162,N_4170);
and U5406 (N_5406,N_594,N_4350);
or U5407 (N_5407,N_1719,N_1037);
or U5408 (N_5408,N_848,N_1027);
and U5409 (N_5409,N_3293,N_3408);
or U5410 (N_5410,N_2083,N_178);
nand U5411 (N_5411,N_2985,N_4328);
nand U5412 (N_5412,N_2250,N_884);
nor U5413 (N_5413,N_1232,N_3223);
nand U5414 (N_5414,N_4690,N_891);
or U5415 (N_5415,N_2000,N_2612);
nand U5416 (N_5416,N_409,N_4637);
nor U5417 (N_5417,N_585,N_3946);
nand U5418 (N_5418,N_3177,N_2011);
or U5419 (N_5419,N_2251,N_96);
nand U5420 (N_5420,N_342,N_1254);
nor U5421 (N_5421,N_727,N_3659);
nor U5422 (N_5422,N_138,N_4840);
nor U5423 (N_5423,N_3160,N_4693);
nand U5424 (N_5424,N_4456,N_3327);
nand U5425 (N_5425,N_1564,N_2993);
and U5426 (N_5426,N_3306,N_3836);
and U5427 (N_5427,N_785,N_2709);
nor U5428 (N_5428,N_2130,N_3218);
nand U5429 (N_5429,N_3325,N_1543);
nand U5430 (N_5430,N_3457,N_345);
nand U5431 (N_5431,N_261,N_3417);
or U5432 (N_5432,N_691,N_3454);
or U5433 (N_5433,N_4890,N_558);
xor U5434 (N_5434,N_4267,N_2533);
nand U5435 (N_5435,N_4402,N_172);
nand U5436 (N_5436,N_1720,N_1802);
and U5437 (N_5437,N_188,N_4398);
nand U5438 (N_5438,N_3399,N_2499);
and U5439 (N_5439,N_460,N_926);
or U5440 (N_5440,N_4375,N_3513);
nor U5441 (N_5441,N_1934,N_780);
nor U5442 (N_5442,N_4076,N_2528);
or U5443 (N_5443,N_4557,N_3027);
and U5444 (N_5444,N_4176,N_4112);
or U5445 (N_5445,N_50,N_1373);
or U5446 (N_5446,N_3853,N_2441);
and U5447 (N_5447,N_2155,N_4345);
nor U5448 (N_5448,N_4600,N_1672);
nor U5449 (N_5449,N_3758,N_133);
nor U5450 (N_5450,N_978,N_673);
or U5451 (N_5451,N_532,N_2341);
nor U5452 (N_5452,N_1269,N_3203);
nor U5453 (N_5453,N_4570,N_620);
and U5454 (N_5454,N_4605,N_3963);
or U5455 (N_5455,N_49,N_1125);
nor U5456 (N_5456,N_4524,N_3931);
nor U5457 (N_5457,N_1351,N_117);
or U5458 (N_5458,N_3862,N_522);
nor U5459 (N_5459,N_315,N_4408);
nand U5460 (N_5460,N_4723,N_143);
or U5461 (N_5461,N_1794,N_2257);
nor U5462 (N_5462,N_1222,N_3554);
nor U5463 (N_5463,N_1428,N_2766);
nor U5464 (N_5464,N_4031,N_3891);
and U5465 (N_5465,N_3547,N_3588);
nor U5466 (N_5466,N_4713,N_297);
and U5467 (N_5467,N_1362,N_4625);
and U5468 (N_5468,N_6,N_2796);
or U5469 (N_5469,N_2389,N_4820);
and U5470 (N_5470,N_2445,N_1777);
and U5471 (N_5471,N_3933,N_3889);
and U5472 (N_5472,N_2163,N_1646);
and U5473 (N_5473,N_2799,N_430);
and U5474 (N_5474,N_1000,N_2255);
nor U5475 (N_5475,N_4136,N_401);
nor U5476 (N_5476,N_2679,N_1690);
and U5477 (N_5477,N_4541,N_1343);
and U5478 (N_5478,N_685,N_3173);
nand U5479 (N_5479,N_3181,N_2670);
or U5480 (N_5480,N_4615,N_1839);
or U5481 (N_5481,N_1820,N_2239);
nor U5482 (N_5482,N_1842,N_556);
or U5483 (N_5483,N_193,N_2537);
or U5484 (N_5484,N_3215,N_3276);
nand U5485 (N_5485,N_2304,N_3354);
and U5486 (N_5486,N_1806,N_607);
nand U5487 (N_5487,N_3199,N_1641);
xnor U5488 (N_5488,N_3265,N_2863);
and U5489 (N_5489,N_4307,N_2065);
nor U5490 (N_5490,N_4029,N_3388);
nor U5491 (N_5491,N_1846,N_4638);
nor U5492 (N_5492,N_3717,N_4926);
nand U5493 (N_5493,N_2234,N_1192);
and U5494 (N_5494,N_1298,N_3118);
and U5495 (N_5495,N_2639,N_3049);
nor U5496 (N_5496,N_1931,N_2572);
nor U5497 (N_5497,N_2792,N_1799);
nand U5498 (N_5498,N_4662,N_4125);
and U5499 (N_5499,N_51,N_3051);
nand U5500 (N_5500,N_2953,N_2736);
nand U5501 (N_5501,N_2839,N_1566);
or U5502 (N_5502,N_4340,N_551);
nand U5503 (N_5503,N_1535,N_4990);
and U5504 (N_5504,N_943,N_496);
and U5505 (N_5505,N_3808,N_4748);
nor U5506 (N_5506,N_2253,N_3390);
and U5507 (N_5507,N_4616,N_4751);
or U5508 (N_5508,N_1256,N_4413);
and U5509 (N_5509,N_114,N_2371);
or U5510 (N_5510,N_1472,N_2368);
and U5511 (N_5511,N_2104,N_4959);
or U5512 (N_5512,N_3932,N_4320);
and U5513 (N_5513,N_572,N_4150);
nor U5514 (N_5514,N_4151,N_46);
or U5515 (N_5515,N_421,N_580);
and U5516 (N_5516,N_2348,N_1303);
nor U5517 (N_5517,N_1073,N_4036);
and U5518 (N_5518,N_4777,N_3464);
nor U5519 (N_5519,N_2743,N_3330);
nand U5520 (N_5520,N_4011,N_1914);
and U5521 (N_5521,N_3092,N_4738);
or U5522 (N_5522,N_1101,N_4517);
nand U5523 (N_5523,N_254,N_1590);
or U5524 (N_5524,N_3999,N_2050);
and U5525 (N_5525,N_333,N_2808);
or U5526 (N_5526,N_4080,N_763);
nor U5527 (N_5527,N_3920,N_1737);
nand U5528 (N_5528,N_2767,N_3574);
or U5529 (N_5529,N_2124,N_1644);
nor U5530 (N_5530,N_732,N_1958);
nand U5531 (N_5531,N_2047,N_2934);
or U5532 (N_5532,N_1152,N_1861);
or U5533 (N_5533,N_251,N_4177);
or U5534 (N_5534,N_1286,N_2144);
nand U5535 (N_5535,N_3972,N_127);
or U5536 (N_5536,N_1695,N_3167);
nand U5537 (N_5537,N_3138,N_1451);
nor U5538 (N_5538,N_796,N_653);
nand U5539 (N_5539,N_4567,N_4212);
nor U5540 (N_5540,N_1454,N_2061);
xor U5541 (N_5541,N_1952,N_2580);
xor U5542 (N_5542,N_3593,N_688);
and U5543 (N_5543,N_4163,N_2861);
nor U5544 (N_5544,N_1706,N_2415);
nand U5545 (N_5545,N_3405,N_1470);
or U5546 (N_5546,N_4124,N_2785);
nor U5547 (N_5547,N_1612,N_2330);
or U5548 (N_5548,N_2233,N_66);
nand U5549 (N_5549,N_776,N_4741);
or U5550 (N_5550,N_3449,N_2611);
or U5551 (N_5551,N_3535,N_4934);
nor U5552 (N_5552,N_3079,N_3674);
nand U5553 (N_5553,N_3517,N_2758);
or U5554 (N_5554,N_1170,N_923);
and U5555 (N_5555,N_281,N_819);
nor U5556 (N_5556,N_4786,N_3846);
and U5557 (N_5557,N_3843,N_3227);
nand U5558 (N_5558,N_4547,N_1774);
or U5559 (N_5559,N_2185,N_16);
and U5560 (N_5560,N_4363,N_627);
nor U5561 (N_5561,N_1278,N_239);
or U5562 (N_5562,N_3236,N_1526);
and U5563 (N_5563,N_45,N_4368);
and U5564 (N_5564,N_2325,N_2284);
and U5565 (N_5565,N_830,N_930);
and U5566 (N_5566,N_4037,N_813);
nor U5567 (N_5567,N_4602,N_3803);
nor U5568 (N_5568,N_4470,N_1411);
nor U5569 (N_5569,N_155,N_338);
nand U5570 (N_5570,N_1553,N_1017);
nand U5571 (N_5571,N_2328,N_2016);
and U5572 (N_5572,N_270,N_2220);
or U5573 (N_5573,N_4305,N_519);
nand U5574 (N_5574,N_868,N_4710);
and U5575 (N_5575,N_3995,N_1808);
nand U5576 (N_5576,N_3437,N_2931);
nand U5577 (N_5577,N_874,N_1217);
and U5578 (N_5578,N_748,N_166);
nand U5579 (N_5579,N_2723,N_1050);
or U5580 (N_5580,N_999,N_4105);
nand U5581 (N_5581,N_4696,N_1209);
nor U5582 (N_5582,N_608,N_4687);
xnor U5583 (N_5583,N_3546,N_4110);
or U5584 (N_5584,N_1926,N_2508);
nor U5585 (N_5585,N_4071,N_3219);
nor U5586 (N_5586,N_4595,N_1676);
or U5587 (N_5587,N_4416,N_2690);
nand U5588 (N_5588,N_1753,N_2957);
and U5589 (N_5589,N_3212,N_2198);
nor U5590 (N_5590,N_596,N_1583);
nor U5591 (N_5591,N_568,N_395);
and U5592 (N_5592,N_1289,N_3491);
and U5593 (N_5593,N_3341,N_3702);
or U5594 (N_5594,N_3232,N_1115);
nor U5595 (N_5595,N_1785,N_2602);
or U5596 (N_5596,N_1980,N_692);
nor U5597 (N_5597,N_3577,N_175);
nand U5598 (N_5598,N_1887,N_351);
nand U5599 (N_5599,N_1512,N_1999);
and U5600 (N_5600,N_3882,N_3056);
nand U5601 (N_5601,N_3880,N_3459);
nor U5602 (N_5602,N_4128,N_4424);
nand U5603 (N_5603,N_2735,N_2491);
nand U5604 (N_5604,N_2280,N_4537);
nor U5605 (N_5605,N_59,N_3934);
nand U5606 (N_5606,N_3194,N_1358);
nor U5607 (N_5607,N_4828,N_4330);
and U5608 (N_5608,N_681,N_4608);
and U5609 (N_5609,N_1961,N_3610);
and U5610 (N_5610,N_4326,N_675);
or U5611 (N_5611,N_1893,N_2465);
nand U5612 (N_5612,N_1225,N_3505);
nand U5613 (N_5613,N_3989,N_325);
and U5614 (N_5614,N_2843,N_4670);
nor U5615 (N_5615,N_1649,N_145);
or U5616 (N_5616,N_4717,N_1993);
nand U5617 (N_5617,N_1950,N_4643);
nor U5618 (N_5618,N_3712,N_3697);
nand U5619 (N_5619,N_4698,N_2698);
or U5620 (N_5620,N_2446,N_2687);
nand U5621 (N_5621,N_894,N_2529);
or U5622 (N_5622,N_3654,N_3901);
or U5623 (N_5623,N_2983,N_1464);
nor U5624 (N_5624,N_1021,N_1684);
nand U5625 (N_5625,N_2094,N_2935);
nor U5626 (N_5626,N_525,N_4287);
nor U5627 (N_5627,N_2967,N_3581);
nor U5628 (N_5628,N_4987,N_3297);
or U5629 (N_5629,N_1218,N_1237);
nor U5630 (N_5630,N_3303,N_2158);
nor U5631 (N_5631,N_1811,N_1432);
or U5632 (N_5632,N_3802,N_1112);
and U5633 (N_5633,N_2724,N_3930);
nand U5634 (N_5634,N_4366,N_773);
or U5635 (N_5635,N_1817,N_3608);
or U5636 (N_5636,N_814,N_4861);
nand U5637 (N_5637,N_4053,N_700);
and U5638 (N_5638,N_265,N_4535);
nor U5639 (N_5639,N_20,N_841);
and U5640 (N_5640,N_1018,N_1578);
nor U5641 (N_5641,N_3871,N_3003);
nand U5642 (N_5642,N_283,N_2172);
nor U5643 (N_5643,N_639,N_2333);
nand U5644 (N_5644,N_2166,N_1747);
nand U5645 (N_5645,N_2058,N_3496);
and U5646 (N_5646,N_4569,N_523);
and U5647 (N_5647,N_3628,N_62);
or U5648 (N_5648,N_4097,N_4199);
nand U5649 (N_5649,N_3171,N_2903);
nor U5650 (N_5650,N_2619,N_4451);
nor U5651 (N_5651,N_3234,N_1202);
or U5652 (N_5652,N_4905,N_3525);
and U5653 (N_5653,N_4682,N_1163);
and U5654 (N_5654,N_2345,N_106);
and U5655 (N_5655,N_869,N_191);
and U5656 (N_5656,N_4783,N_2420);
and U5657 (N_5657,N_1663,N_1648);
or U5658 (N_5658,N_1760,N_1079);
nor U5659 (N_5659,N_2650,N_1339);
nand U5660 (N_5660,N_1251,N_411);
nand U5661 (N_5661,N_3866,N_3818);
nor U5662 (N_5662,N_909,N_2290);
nor U5663 (N_5663,N_718,N_1183);
or U5664 (N_5664,N_2302,N_3631);
or U5665 (N_5665,N_3272,N_4597);
nor U5666 (N_5666,N_2784,N_4931);
nor U5667 (N_5667,N_4774,N_3287);
nor U5668 (N_5668,N_3271,N_1742);
or U5669 (N_5669,N_2635,N_628);
or U5670 (N_5670,N_3976,N_1407);
nor U5671 (N_5671,N_3085,N_1569);
or U5672 (N_5672,N_3349,N_55);
nor U5673 (N_5673,N_4360,N_4362);
nor U5674 (N_5674,N_369,N_687);
nand U5675 (N_5675,N_1484,N_294);
nor U5676 (N_5676,N_3617,N_238);
or U5677 (N_5677,N_3632,N_838);
xnor U5678 (N_5678,N_3865,N_3020);
nor U5679 (N_5679,N_716,N_4640);
xnor U5680 (N_5680,N_1740,N_4334);
or U5681 (N_5681,N_762,N_1609);
and U5682 (N_5682,N_717,N_4801);
or U5683 (N_5683,N_2096,N_2941);
or U5684 (N_5684,N_4485,N_1022);
and U5685 (N_5685,N_3387,N_3751);
or U5686 (N_5686,N_683,N_985);
nand U5687 (N_5687,N_811,N_4272);
nor U5688 (N_5688,N_2361,N_3176);
nor U5689 (N_5689,N_3217,N_2300);
or U5690 (N_5690,N_901,N_4651);
xor U5691 (N_5691,N_3533,N_4930);
nand U5692 (N_5692,N_4787,N_2296);
nand U5693 (N_5693,N_4095,N_1640);
nand U5694 (N_5694,N_1426,N_1750);
or U5695 (N_5695,N_2979,N_3291);
nand U5696 (N_5696,N_3211,N_1499);
xor U5697 (N_5697,N_1458,N_3650);
and U5698 (N_5698,N_2405,N_3668);
nor U5699 (N_5699,N_4414,N_4791);
nand U5700 (N_5700,N_356,N_2823);
or U5701 (N_5701,N_1957,N_2159);
nand U5702 (N_5702,N_4908,N_2098);
or U5703 (N_5703,N_420,N_416);
or U5704 (N_5704,N_3110,N_2087);
nor U5705 (N_5705,N_590,N_2471);
nor U5706 (N_5706,N_834,N_2996);
and U5707 (N_5707,N_1881,N_1892);
and U5708 (N_5708,N_2173,N_4231);
or U5709 (N_5709,N_4487,N_2846);
nor U5710 (N_5710,N_3127,N_4722);
or U5711 (N_5711,N_4577,N_3665);
and U5712 (N_5712,N_3607,N_3286);
nand U5713 (N_5713,N_1544,N_1924);
and U5714 (N_5714,N_2591,N_1492);
or U5715 (N_5715,N_1692,N_292);
and U5716 (N_5716,N_3134,N_1832);
nand U5717 (N_5717,N_2103,N_1009);
xnor U5718 (N_5718,N_4126,N_2459);
and U5719 (N_5719,N_104,N_2654);
nand U5720 (N_5720,N_1386,N_2976);
nand U5721 (N_5721,N_3277,N_2675);
and U5722 (N_5722,N_2357,N_4490);
and U5723 (N_5723,N_738,N_1075);
or U5724 (N_5724,N_3004,N_546);
and U5725 (N_5725,N_1705,N_967);
and U5726 (N_5726,N_1223,N_2379);
or U5727 (N_5727,N_423,N_3766);
or U5728 (N_5728,N_1460,N_4491);
and U5729 (N_5729,N_3804,N_1403);
or U5730 (N_5730,N_1682,N_1459);
nand U5731 (N_5731,N_676,N_3377);
and U5732 (N_5732,N_4038,N_1599);
and U5733 (N_5733,N_125,N_3530);
nand U5734 (N_5734,N_4395,N_1597);
nand U5735 (N_5735,N_4810,N_11);
and U5736 (N_5736,N_2316,N_386);
and U5737 (N_5737,N_2945,N_2954);
xnor U5738 (N_5738,N_70,N_2084);
nor U5739 (N_5739,N_3633,N_1190);
nor U5740 (N_5740,N_4496,N_2885);
or U5741 (N_5741,N_309,N_3314);
nor U5742 (N_5742,N_2313,N_1389);
nor U5743 (N_5743,N_870,N_3929);
nand U5744 (N_5744,N_4254,N_29);
nand U5745 (N_5745,N_1212,N_672);
or U5746 (N_5746,N_4860,N_28);
xnor U5747 (N_5747,N_1605,N_613);
or U5748 (N_5748,N_1983,N_3619);
or U5749 (N_5749,N_76,N_257);
xnor U5750 (N_5750,N_3391,N_329);
nand U5751 (N_5751,N_2218,N_2043);
nand U5752 (N_5752,N_174,N_3660);
and U5753 (N_5753,N_2637,N_2165);
nor U5754 (N_5754,N_4186,N_3974);
xnor U5755 (N_5755,N_3596,N_921);
and U5756 (N_5756,N_2893,N_2610);
or U5757 (N_5757,N_1724,N_1408);
nor U5758 (N_5758,N_3331,N_1158);
or U5759 (N_5759,N_965,N_1184);
and U5760 (N_5760,N_4335,N_1107);
or U5761 (N_5761,N_1272,N_1002);
nand U5762 (N_5762,N_4808,N_57);
or U5763 (N_5763,N_2965,N_1195);
nand U5764 (N_5764,N_1784,N_3309);
nor U5765 (N_5765,N_3337,N_3907);
or U5766 (N_5766,N_2223,N_4131);
or U5767 (N_5767,N_1966,N_3019);
and U5768 (N_5768,N_680,N_4171);
or U5769 (N_5769,N_1546,N_236);
nor U5770 (N_5770,N_3616,N_3410);
and U5771 (N_5771,N_1359,N_2141);
or U5772 (N_5772,N_299,N_3956);
xor U5773 (N_5773,N_266,N_3365);
nand U5774 (N_5774,N_2497,N_4476);
or U5775 (N_5775,N_1294,N_407);
nor U5776 (N_5776,N_4106,N_3861);
nand U5777 (N_5777,N_1897,N_3157);
nor U5778 (N_5778,N_3200,N_4902);
or U5779 (N_5779,N_255,N_398);
and U5780 (N_5780,N_3921,N_1148);
nand U5781 (N_5781,N_2247,N_3694);
nor U5782 (N_5782,N_2490,N_153);
or U5783 (N_5783,N_3097,N_3007);
nor U5784 (N_5784,N_3151,N_4331);
or U5785 (N_5785,N_3814,N_4778);
nor U5786 (N_5786,N_128,N_68);
or U5787 (N_5787,N_310,N_3655);
nor U5788 (N_5788,N_3304,N_3450);
and U5789 (N_5789,N_4782,N_1145);
nor U5790 (N_5790,N_1670,N_872);
nor U5791 (N_5791,N_349,N_141);
and U5792 (N_5792,N_4944,N_3868);
nor U5793 (N_5793,N_1399,N_4803);
nor U5794 (N_5794,N_1137,N_4716);
or U5795 (N_5795,N_3584,N_4198);
nand U5796 (N_5796,N_4457,N_1756);
and U5797 (N_5797,N_4603,N_4498);
and U5798 (N_5798,N_122,N_2106);
nor U5799 (N_5799,N_1933,N_4796);
and U5800 (N_5800,N_1405,N_3640);
nand U5801 (N_5801,N_4921,N_3763);
and U5802 (N_5802,N_4488,N_3571);
and U5803 (N_5803,N_2806,N_1736);
nor U5804 (N_5804,N_2430,N_586);
and U5805 (N_5805,N_982,N_3196);
nand U5806 (N_5806,N_4099,N_2575);
nor U5807 (N_5807,N_1951,N_1363);
nor U5808 (N_5808,N_455,N_1841);
nand U5809 (N_5809,N_3476,N_954);
nor U5810 (N_5810,N_3074,N_4845);
or U5811 (N_5811,N_3973,N_1550);
or U5812 (N_5812,N_4192,N_2034);
nor U5813 (N_5813,N_4542,N_1084);
nand U5814 (N_5814,N_4436,N_1572);
or U5815 (N_5815,N_1639,N_4967);
and U5816 (N_5816,N_4428,N_4359);
nand U5817 (N_5817,N_3507,N_3435);
xnor U5818 (N_5818,N_1032,N_1033);
nand U5819 (N_5819,N_3339,N_2947);
xnor U5820 (N_5820,N_4083,N_1035);
or U5821 (N_5821,N_549,N_4431);
and U5822 (N_5822,N_4242,N_3602);
nor U5823 (N_5823,N_1948,N_632);
or U5824 (N_5824,N_4094,N_3677);
and U5825 (N_5825,N_4680,N_1360);
nor U5826 (N_5826,N_792,N_1069);
nor U5827 (N_5827,N_1949,N_2840);
and U5828 (N_5828,N_2265,N_4761);
and U5829 (N_5829,N_2872,N_4103);
nor U5830 (N_5830,N_4957,N_1985);
nand U5831 (N_5831,N_3198,N_228);
nor U5832 (N_5832,N_3475,N_3939);
and U5833 (N_5833,N_3542,N_4996);
nand U5834 (N_5834,N_4239,N_437);
nor U5835 (N_5835,N_2753,N_2745);
nand U5836 (N_5836,N_3701,N_2662);
or U5837 (N_5837,N_3149,N_2092);
nand U5838 (N_5838,N_2052,N_2232);
and U5839 (N_5839,N_664,N_1392);
and U5840 (N_5840,N_2955,N_295);
or U5841 (N_5841,N_752,N_3486);
nand U5842 (N_5842,N_4587,N_2521);
nand U5843 (N_5843,N_2048,N_958);
and U5844 (N_5844,N_1689,N_603);
or U5845 (N_5845,N_194,N_3703);
nand U5846 (N_5846,N_2209,N_307);
nor U5847 (N_5847,N_2444,N_4086);
and U5848 (N_5848,N_616,N_359);
or U5849 (N_5849,N_4219,N_1552);
xnor U5850 (N_5850,N_1091,N_612);
nor U5851 (N_5851,N_2535,N_4437);
and U5852 (N_5852,N_3690,N_2134);
nor U5853 (N_5853,N_1189,N_4014);
and U5854 (N_5854,N_697,N_2664);
nor U5855 (N_5855,N_75,N_2044);
and U5856 (N_5856,N_4672,N_4566);
nand U5857 (N_5857,N_2256,N_3468);
nor U5858 (N_5858,N_4197,N_3404);
and U5859 (N_5859,N_1093,N_442);
and U5860 (N_5860,N_3586,N_165);
and U5861 (N_5861,N_1733,N_3374);
nand U5862 (N_5862,N_650,N_1160);
or U5863 (N_5863,N_4676,N_3226);
or U5864 (N_5864,N_2364,N_1879);
and U5865 (N_5865,N_2169,N_3237);
nor U5866 (N_5866,N_4285,N_1133);
nor U5867 (N_5867,N_249,N_1296);
nor U5868 (N_5868,N_3319,N_2352);
or U5869 (N_5869,N_641,N_2899);
nor U5870 (N_5870,N_392,N_2582);
nand U5871 (N_5871,N_4303,N_509);
nor U5872 (N_5872,N_2273,N_0);
and U5873 (N_5873,N_2622,N_3222);
nor U5874 (N_5874,N_882,N_196);
nor U5875 (N_5875,N_659,N_4472);
and U5876 (N_5876,N_719,N_4253);
or U5877 (N_5877,N_3014,N_3984);
and U5878 (N_5878,N_840,N_3943);
nor U5879 (N_5879,N_451,N_3842);
nor U5880 (N_5880,N_4020,N_316);
nor U5881 (N_5881,N_4200,N_4503);
and U5882 (N_5882,N_3795,N_2609);
nor U5883 (N_5883,N_726,N_3065);
nor U5884 (N_5884,N_1463,N_1909);
nor U5885 (N_5885,N_4127,N_2633);
and U5886 (N_5886,N_3242,N_2642);
and U5887 (N_5887,N_1263,N_212);
and U5888 (N_5888,N_1700,N_740);
and U5889 (N_5889,N_2697,N_4019);
nand U5890 (N_5890,N_2168,N_44);
nand U5891 (N_5891,N_1855,N_4407);
or U5892 (N_5892,N_4897,N_536);
and U5893 (N_5893,N_4747,N_109);
or U5894 (N_5894,N_301,N_4232);
nor U5895 (N_5895,N_3031,N_2925);
nand U5896 (N_5896,N_4753,N_4461);
and U5897 (N_5897,N_1387,N_2111);
or U5898 (N_5898,N_1349,N_779);
and U5899 (N_5899,N_3087,N_113);
or U5900 (N_5900,N_3941,N_837);
or U5901 (N_5901,N_4137,N_3578);
nand U5902 (N_5902,N_1826,N_2298);
and U5903 (N_5903,N_3488,N_231);
and U5904 (N_5904,N_3844,N_3106);
and U5905 (N_5905,N_1108,N_2225);
or U5906 (N_5906,N_4286,N_1900);
nor U5907 (N_5907,N_772,N_2715);
nand U5908 (N_5908,N_1686,N_4323);
or U5909 (N_5909,N_4465,N_3083);
nand U5910 (N_5910,N_149,N_2411);
and U5911 (N_5911,N_4108,N_3063);
and U5912 (N_5912,N_1130,N_4576);
nor U5913 (N_5913,N_4068,N_2161);
nor U5914 (N_5914,N_1699,N_531);
nor U5915 (N_5915,N_1981,N_4012);
or U5916 (N_5916,N_3392,N_248);
nand U5917 (N_5917,N_1623,N_4052);
or U5918 (N_5918,N_3109,N_3924);
or U5919 (N_5919,N_2797,N_2502);
and U5920 (N_5920,N_2079,N_4953);
nand U5921 (N_5921,N_1688,N_2701);
nand U5922 (N_5922,N_1815,N_4574);
and U5923 (N_5923,N_3088,N_2558);
nor U5924 (N_5924,N_2214,N_4914);
and U5925 (N_5925,N_4925,N_377);
and U5926 (N_5926,N_2127,N_4737);
nand U5927 (N_5927,N_4224,N_502);
nand U5928 (N_5928,N_2360,N_376);
nand U5929 (N_5929,N_2235,N_4964);
nor U5930 (N_5930,N_1943,N_2645);
nor U5931 (N_5931,N_1175,N_3183);
or U5932 (N_5932,N_1083,N_1097);
or U5933 (N_5933,N_195,N_4118);
nand U5934 (N_5934,N_2195,N_1082);
and U5935 (N_5935,N_206,N_3624);
nand U5936 (N_5936,N_2204,N_4299);
or U5937 (N_5937,N_4780,N_4998);
and U5938 (N_5938,N_462,N_4054);
or U5939 (N_5939,N_4869,N_1814);
nand U5940 (N_5940,N_2488,N_3310);
nand U5941 (N_5941,N_78,N_3753);
nand U5942 (N_5942,N_3270,N_3892);
or U5943 (N_5943,N_1257,N_4149);
nand U5944 (N_5944,N_662,N_883);
or U5945 (N_5945,N_1396,N_1517);
xor U5946 (N_5946,N_1624,N_4644);
or U5947 (N_5947,N_1987,N_2373);
and U5948 (N_5948,N_2781,N_322);
nor U5949 (N_5949,N_3427,N_4976);
nor U5950 (N_5950,N_1575,N_475);
or U5951 (N_5951,N_2164,N_391);
nor U5952 (N_5952,N_2068,N_2351);
and U5953 (N_5953,N_668,N_1292);
or U5954 (N_5954,N_3724,N_1457);
and U5955 (N_5955,N_373,N_198);
nor U5956 (N_5956,N_375,N_1656);
or U5957 (N_5957,N_2803,N_3154);
nor U5958 (N_5958,N_1078,N_2722);
or U5959 (N_5959,N_2737,N_4769);
and U5960 (N_5960,N_4800,N_1642);
nand U5961 (N_5961,N_4811,N_3145);
or U5962 (N_5962,N_4849,N_2626);
and U5963 (N_5963,N_1336,N_919);
or U5964 (N_5964,N_759,N_121);
nand U5965 (N_5965,N_1178,N_1587);
and U5966 (N_5966,N_4088,N_1162);
nand U5967 (N_5967,N_2531,N_637);
nand U5968 (N_5968,N_3641,N_3452);
nor U5969 (N_5969,N_3935,N_2911);
or U5970 (N_5970,N_3462,N_1812);
nor U5971 (N_5971,N_4278,N_3509);
or U5972 (N_5972,N_2651,N_1913);
and U5973 (N_5973,N_2171,N_2655);
or U5974 (N_5974,N_1317,N_1406);
nand U5975 (N_5975,N_635,N_3600);
nand U5976 (N_5976,N_3845,N_3282);
or U5977 (N_5977,N_2203,N_88);
nand U5978 (N_5978,N_4657,N_2066);
or U5979 (N_5979,N_998,N_3418);
xor U5980 (N_5980,N_48,N_2588);
or U5981 (N_5981,N_3637,N_2587);
nor U5982 (N_5982,N_1118,N_1319);
or U5983 (N_5983,N_1673,N_4938);
or U5984 (N_5984,N_2756,N_3664);
nor U5985 (N_5985,N_638,N_4240);
or U5986 (N_5986,N_328,N_2182);
or U5987 (N_5987,N_207,N_4183);
nor U5988 (N_5988,N_1751,N_4440);
or U5989 (N_5989,N_1791,N_190);
or U5990 (N_5990,N_433,N_1625);
and U5991 (N_5991,N_144,N_4579);
xnor U5992 (N_5992,N_4527,N_871);
and U5993 (N_5993,N_4622,N_350);
nor U5994 (N_5994,N_510,N_3728);
and U5995 (N_5995,N_3500,N_390);
nor U5996 (N_5996,N_2617,N_234);
nand U5997 (N_5997,N_3849,N_3368);
xor U5998 (N_5998,N_2805,N_240);
or U5999 (N_5999,N_3143,N_2320);
and U6000 (N_6000,N_521,N_2498);
nand U6001 (N_6001,N_176,N_2817);
and U6002 (N_6002,N_2309,N_79);
nand U6003 (N_6003,N_4767,N_2998);
nand U6004 (N_6004,N_4130,N_524);
nand U6005 (N_6005,N_1340,N_3426);
nand U6006 (N_6006,N_2746,N_1787);
and U6007 (N_6007,N_3372,N_361);
or U6008 (N_6008,N_624,N_803);
nor U6009 (N_6009,N_2271,N_3447);
nor U6010 (N_6010,N_1722,N_4321);
and U6011 (N_6011,N_3121,N_3740);
and U6012 (N_6012,N_1347,N_3768);
nor U6013 (N_6013,N_4671,N_22);
and U6014 (N_6014,N_3806,N_1151);
or U6015 (N_6015,N_4588,N_4);
nand U6016 (N_6016,N_2755,N_1801);
nor U6017 (N_6017,N_184,N_3902);
or U6018 (N_6018,N_4258,N_3105);
and U6019 (N_6019,N_2137,N_3254);
nand U6020 (N_6020,N_1172,N_4384);
nand U6021 (N_6021,N_1046,N_3592);
or U6022 (N_6022,N_1921,N_2397);
nor U6023 (N_6023,N_3864,N_3050);
nor U6024 (N_6024,N_3338,N_4619);
nor U6025 (N_6025,N_3983,N_1604);
and U6026 (N_6026,N_3979,N_1589);
or U6027 (N_6027,N_348,N_2815);
or U6028 (N_6028,N_2643,N_2666);
and U6029 (N_6029,N_36,N_4047);
nand U6030 (N_6030,N_4614,N_2754);
nand U6031 (N_6031,N_1490,N_4338);
or U6032 (N_6032,N_2384,N_3527);
or U6033 (N_6033,N_4582,N_744);
and U6034 (N_6034,N_4314,N_815);
and U6035 (N_6035,N_3130,N_2852);
nand U6036 (N_6036,N_2378,N_1904);
and U6037 (N_6037,N_1198,N_2706);
or U6038 (N_6038,N_2053,N_3326);
and U6039 (N_6039,N_4847,N_91);
and U6040 (N_6040,N_3204,N_863);
nor U6041 (N_6041,N_2778,N_988);
nor U6042 (N_6042,N_4590,N_3982);
or U6043 (N_6043,N_997,N_1824);
or U6044 (N_6044,N_3245,N_2242);
nor U6045 (N_6045,N_3350,N_4514);
nor U6046 (N_6046,N_1486,N_2673);
nand U6047 (N_6047,N_1853,N_1203);
nor U6048 (N_6048,N_3422,N_1850);
or U6049 (N_6049,N_3539,N_2939);
or U6050 (N_6050,N_4851,N_1167);
or U6051 (N_6051,N_4248,N_4115);
and U6052 (N_6052,N_670,N_289);
nand U6053 (N_6053,N_3133,N_2076);
or U6054 (N_6054,N_2851,N_858);
nor U6055 (N_6055,N_2894,N_2303);
or U6056 (N_6056,N_474,N_4309);
and U6057 (N_6057,N_1350,N_736);
nand U6058 (N_6058,N_2669,N_1041);
or U6059 (N_6059,N_2281,N_83);
and U6060 (N_6060,N_341,N_1056);
and U6061 (N_6061,N_2414,N_4548);
nor U6062 (N_6062,N_1052,N_1889);
or U6063 (N_6063,N_1315,N_1998);
and U6064 (N_6064,N_3949,N_2272);
nor U6065 (N_6065,N_4941,N_1038);
and U6066 (N_6066,N_602,N_2317);
or U6067 (N_6067,N_1795,N_3278);
xor U6068 (N_6068,N_1710,N_2429);
and U6069 (N_6069,N_808,N_4439);
or U6070 (N_6070,N_3784,N_1528);
or U6071 (N_6071,N_107,N_2227);
or U6072 (N_6072,N_1281,N_1391);
or U6073 (N_6073,N_3783,N_3453);
or U6074 (N_6074,N_787,N_3811);
or U6075 (N_6075,N_1616,N_3064);
and U6076 (N_6076,N_3340,N_2477);
or U6077 (N_6077,N_2015,N_1089);
or U6078 (N_6078,N_1849,N_3821);
nor U6079 (N_6079,N_3478,N_4261);
nor U6080 (N_6080,N_3479,N_2452);
and U6081 (N_6081,N_1978,N_630);
nor U6082 (N_6082,N_3591,N_671);
and U6083 (N_6083,N_4565,N_949);
nand U6084 (N_6084,N_4235,N_3318);
nand U6085 (N_6085,N_2989,N_2007);
nor U6086 (N_6086,N_1935,N_979);
nor U6087 (N_6087,N_3678,N_2107);
nor U6088 (N_6088,N_4821,N_3298);
xnor U6089 (N_6089,N_477,N_4445);
or U6090 (N_6090,N_4888,N_2628);
nand U6091 (N_6091,N_2777,N_4444);
and U6092 (N_6092,N_3268,N_724);
nor U6093 (N_6093,N_2421,N_713);
nor U6094 (N_6094,N_3782,N_3625);
and U6095 (N_6095,N_38,N_2010);
and U6096 (N_6096,N_4139,N_3166);
nor U6097 (N_6097,N_571,N_904);
and U6098 (N_6098,N_4066,N_4265);
and U6099 (N_6099,N_1888,N_1300);
nor U6100 (N_6100,N_151,N_3244);
and U6101 (N_6101,N_1843,N_1885);
nand U6102 (N_6102,N_2980,N_2629);
nand U6103 (N_6103,N_4188,N_1804);
nand U6104 (N_6104,N_1299,N_2870);
and U6105 (N_6105,N_1282,N_1869);
nand U6106 (N_6106,N_435,N_476);
nor U6107 (N_6107,N_4211,N_1851);
and U6108 (N_6108,N_3825,N_589);
or U6109 (N_6109,N_4409,N_387);
nor U6110 (N_6110,N_3072,N_1752);
or U6111 (N_6111,N_1711,N_1601);
or U6112 (N_6112,N_2436,N_518);
nor U6113 (N_6113,N_4070,N_4952);
or U6114 (N_6114,N_4473,N_1942);
nor U6115 (N_6115,N_1611,N_4369);
nand U6116 (N_6116,N_3580,N_1511);
xnor U6117 (N_6117,N_4705,N_1054);
nor U6118 (N_6118,N_721,N_2907);
and U6119 (N_6119,N_503,N_1567);
nand U6120 (N_6120,N_3013,N_633);
and U6121 (N_6121,N_2199,N_4510);
or U6122 (N_6122,N_1620,N_2908);
and U6123 (N_6123,N_4584,N_3729);
nand U6124 (N_6124,N_4443,N_157);
and U6125 (N_6125,N_3107,N_2783);
nor U6126 (N_6126,N_709,N_2323);
nor U6127 (N_6127,N_4269,N_2056);
and U6128 (N_6128,N_937,N_781);
nor U6129 (N_6129,N_2299,N_1522);
nand U6130 (N_6130,N_4746,N_1185);
nor U6131 (N_6131,N_569,N_783);
or U6132 (N_6132,N_3622,N_3739);
nand U6133 (N_6133,N_1982,N_2975);
nor U6134 (N_6134,N_3730,N_2121);
nor U6135 (N_6135,N_2122,N_1247);
and U6136 (N_6136,N_3923,N_4874);
or U6137 (N_6137,N_3952,N_1557);
or U6138 (N_6138,N_989,N_3235);
and U6139 (N_6139,N_183,N_4315);
and U6140 (N_6140,N_1221,N_2326);
nor U6141 (N_6141,N_4332,N_2991);
or U6142 (N_6142,N_258,N_4950);
and U6143 (N_6143,N_4304,N_3470);
or U6144 (N_6144,N_3260,N_211);
nor U6145 (N_6145,N_821,N_2369);
and U6146 (N_6146,N_2779,N_2279);
and U6147 (N_6147,N_2791,N_185);
nor U6148 (N_6148,N_4295,N_3493);
and U6149 (N_6149,N_2683,N_1095);
or U6150 (N_6150,N_3775,N_4920);
and U6151 (N_6151,N_4100,N_2667);
nor U6152 (N_6152,N_498,N_4159);
and U6153 (N_6153,N_4243,N_4193);
and U6154 (N_6154,N_4980,N_810);
xnor U6155 (N_6155,N_4233,N_2394);
or U6156 (N_6156,N_1045,N_3047);
nand U6157 (N_6157,N_1179,N_3380);
nand U6158 (N_6158,N_739,N_2725);
nor U6159 (N_6159,N_4771,N_3514);
or U6160 (N_6160,N_1366,N_4393);
nand U6161 (N_6161,N_1503,N_1939);
and U6162 (N_6162,N_382,N_120);
or U6163 (N_6163,N_7,N_3446);
and U6164 (N_6164,N_578,N_3011);
or U6165 (N_6165,N_4650,N_454);
and U6166 (N_6166,N_2245,N_805);
nor U6167 (N_6167,N_1384,N_4632);
and U6168 (N_6168,N_4788,N_2968);
or U6169 (N_6169,N_2729,N_2437);
nor U6170 (N_6170,N_4449,N_4280);
or U6171 (N_6171,N_4203,N_554);
nand U6172 (N_6172,N_3538,N_4161);
nor U6173 (N_6173,N_1725,N_3816);
and U6174 (N_6174,N_4895,N_794);
nor U6175 (N_6175,N_2501,N_1447);
nor U6176 (N_6176,N_3207,N_3356);
or U6177 (N_6177,N_895,N_1245);
nand U6178 (N_6178,N_2359,N_2494);
nand U6179 (N_6179,N_123,N_2896);
nand U6180 (N_6180,N_1574,N_108);
nand U6181 (N_6181,N_4852,N_1708);
and U6182 (N_6182,N_4991,N_2618);
and U6183 (N_6183,N_2109,N_4002);
or U6184 (N_6184,N_1157,N_4358);
and U6185 (N_6185,N_3965,N_21);
and U6186 (N_6186,N_2308,N_3187);
or U6187 (N_6187,N_2019,N_553);
nor U6188 (N_6188,N_1588,N_2001);
nand U6189 (N_6189,N_4114,N_816);
and U6190 (N_6190,N_4390,N_2761);
or U6191 (N_6191,N_3394,N_1548);
nor U6192 (N_6192,N_2033,N_2927);
nor U6193 (N_6193,N_408,N_1816);
and U6194 (N_6194,N_4781,N_2603);
nor U6195 (N_6195,N_339,N_2142);
and U6196 (N_6196,N_229,N_1874);
nor U6197 (N_6197,N_2102,N_737);
or U6198 (N_6198,N_80,N_2539);
nand U6199 (N_6199,N_767,N_2700);
nand U6200 (N_6200,N_4441,N_3059);
or U6201 (N_6201,N_3351,N_2905);
nand U6202 (N_6202,N_2112,N_1493);
or U6203 (N_6203,N_1778,N_527);
or U6204 (N_6204,N_3076,N_3830);
or U6205 (N_6205,N_4583,N_2170);
or U6206 (N_6206,N_973,N_1518);
and U6207 (N_6207,N_2620,N_1867);
nor U6208 (N_6208,N_3344,N_1211);
and U6209 (N_6209,N_1905,N_1556);
and U6210 (N_6210,N_1104,N_3001);
or U6211 (N_6211,N_1417,N_1788);
and U6212 (N_6212,N_1884,N_1353);
or U6213 (N_6213,N_2720,N_201);
nand U6214 (N_6214,N_1732,N_1235);
nor U6215 (N_6215,N_1529,N_1227);
or U6216 (N_6216,N_4842,N_722);
nor U6217 (N_6217,N_2406,N_4665);
and U6218 (N_6218,N_4166,N_3412);
and U6219 (N_6219,N_778,N_567);
or U6220 (N_6220,N_626,N_3503);
nand U6221 (N_6221,N_3764,N_4872);
nor U6222 (N_6222,N_1823,N_3205);
and U6223 (N_6223,N_3794,N_90);
nor U6224 (N_6224,N_2848,N_434);
nor U6225 (N_6225,N_1792,N_4817);
nor U6226 (N_6226,N_4311,N_1617);
and U6227 (N_6227,N_4051,N_4468);
and U6228 (N_6228,N_94,N_4418);
nor U6229 (N_6229,N_4628,N_1310);
nand U6230 (N_6230,N_1568,N_4669);
or U6231 (N_6231,N_2475,N_2466);
nand U6232 (N_6232,N_2566,N_4489);
and U6233 (N_6233,N_1857,N_2921);
or U6234 (N_6234,N_3583,N_3359);
or U6235 (N_6235,N_4836,N_699);
and U6236 (N_6236,N_2244,N_354);
and U6237 (N_6237,N_1131,N_4818);
or U6238 (N_6238,N_124,N_4182);
and U6239 (N_6239,N_1029,N_1922);
or U6240 (N_6240,N_2824,N_3732);
or U6241 (N_6241,N_1048,N_3537);
nor U6242 (N_6242,N_1371,N_1124);
and U6243 (N_6243,N_1443,N_4568);
and U6244 (N_6244,N_2691,N_1249);
and U6245 (N_6245,N_3102,N_1577);
and U6246 (N_6246,N_152,N_2088);
and U6247 (N_6247,N_4484,N_3718);
and U6248 (N_6248,N_4205,N_974);
nor U6249 (N_6249,N_1250,N_461);
and U6250 (N_6250,N_1425,N_1514);
nand U6251 (N_6251,N_3767,N_3397);
or U6252 (N_6252,N_4477,N_708);
or U6253 (N_6253,N_4784,N_1615);
or U6254 (N_6254,N_4361,N_2923);
nand U6255 (N_6255,N_3142,N_4916);
nand U6256 (N_6256,N_4009,N_4129);
and U6257 (N_6257,N_4940,N_4289);
nor U6258 (N_6258,N_2889,N_1984);
nand U6259 (N_6259,N_214,N_1694);
or U6260 (N_6260,N_3755,N_1483);
and U6261 (N_6261,N_2009,N_4220);
or U6262 (N_6262,N_4141,N_529);
or U6263 (N_6263,N_3358,N_2516);
xor U6264 (N_6264,N_4901,N_3627);
xor U6265 (N_6265,N_1729,N_4322);
and U6266 (N_6266,N_2789,N_4144);
and U6267 (N_6267,N_3779,N_1119);
and U6268 (N_6268,N_2728,N_4337);
nor U6269 (N_6269,N_4178,N_4256);
and U6270 (N_6270,N_1100,N_2349);
nor U6271 (N_6271,N_4121,N_4530);
nor U6272 (N_6272,N_1236,N_4829);
or U6273 (N_6273,N_950,N_4453);
nor U6274 (N_6274,N_4562,N_2407);
and U6275 (N_6275,N_1513,N_2228);
or U6276 (N_6276,N_4720,N_1238);
nand U6277 (N_6277,N_250,N_2243);
or U6278 (N_6278,N_1378,N_4627);
and U6279 (N_6279,N_3269,N_3489);
and U6280 (N_6280,N_3856,N_2145);
and U6281 (N_6281,N_3756,N_4221);
nor U6282 (N_6282,N_731,N_126);
nor U6283 (N_6283,N_135,N_3009);
nand U6284 (N_6284,N_484,N_87);
nor U6285 (N_6285,N_2229,N_2727);
nand U6286 (N_6286,N_2696,N_3273);
or U6287 (N_6287,N_3086,N_3444);
or U6288 (N_6288,N_1324,N_756);
and U6289 (N_6289,N_3433,N_3113);
or U6290 (N_6290,N_4458,N_610);
or U6291 (N_6291,N_1631,N_548);
and U6292 (N_6292,N_2545,N_33);
nand U6293 (N_6293,N_512,N_1633);
and U6294 (N_6294,N_922,N_619);
nor U6295 (N_6295,N_3925,N_917);
and U6296 (N_6296,N_2422,N_4966);
and U6297 (N_6297,N_4257,N_3415);
or U6298 (N_6298,N_306,N_1697);
or U6299 (N_6299,N_3558,N_646);
or U6300 (N_6300,N_1034,N_1608);
nand U6301 (N_6301,N_2592,N_1153);
nor U6302 (N_6302,N_4325,N_4554);
nor U6303 (N_6303,N_849,N_4018);
nand U6304 (N_6304,N_4045,N_287);
xnor U6305 (N_6305,N_1929,N_2193);
or U6306 (N_6306,N_12,N_4797);
or U6307 (N_6307,N_3575,N_1036);
or U6308 (N_6308,N_4513,N_4403);
or U6309 (N_6309,N_4237,N_2055);
and U6310 (N_6310,N_4191,N_1818);
or U6311 (N_6311,N_372,N_1579);
nand U6312 (N_6312,N_3893,N_714);
nand U6313 (N_6313,N_1085,N_4319);
nor U6314 (N_6314,N_378,N_3940);
nor U6315 (N_6315,N_491,N_2409);
nor U6316 (N_6316,N_4728,N_1423);
nand U6317 (N_6317,N_4873,N_4247);
and U6318 (N_6318,N_933,N_3461);
or U6319 (N_6319,N_399,N_3045);
or U6320 (N_6320,N_1866,N_2809);
and U6321 (N_6321,N_3566,N_4893);
nor U6322 (N_6322,N_71,N_4743);
and U6323 (N_6323,N_1745,N_4718);
and U6324 (N_6324,N_2616,N_4048);
or U6325 (N_6325,N_3054,N_647);
and U6326 (N_6326,N_2093,N_3058);
nand U6327 (N_6327,N_544,N_4173);
nand U6328 (N_6328,N_374,N_134);
nor U6329 (N_6329,N_2689,N_3970);
nor U6330 (N_6330,N_775,N_1004);
and U6331 (N_6331,N_4312,N_1012);
nand U6332 (N_6332,N_2156,N_766);
nand U6333 (N_6333,N_1111,N_3370);
nor U6334 (N_6334,N_3124,N_4978);
or U6335 (N_6335,N_839,N_4809);
nor U6336 (N_6336,N_963,N_3773);
and U6337 (N_6337,N_1647,N_4853);
or U6338 (N_6338,N_3188,N_2071);
nand U6339 (N_6339,N_2382,N_1856);
or U6340 (N_6340,N_2319,N_4142);
and U6341 (N_6341,N_2978,N_2704);
nor U6342 (N_6342,N_1592,N_4598);
nand U6343 (N_6343,N_1780,N_4664);
nor U6344 (N_6344,N_3295,N_4731);
or U6345 (N_6345,N_4175,N_2213);
or U6346 (N_6346,N_2875,N_4032);
nor U6347 (N_6347,N_4734,N_2248);
or U6348 (N_6348,N_4960,N_944);
and U6349 (N_6349,N_3689,N_3912);
nand U6350 (N_6350,N_741,N_835);
nand U6351 (N_6351,N_4555,N_747);
nand U6352 (N_6352,N_1354,N_3651);
nor U6353 (N_6353,N_1790,N_3055);
nand U6354 (N_6354,N_3676,N_599);
or U6355 (N_6355,N_4586,N_1645);
nand U6356 (N_6356,N_3025,N_3238);
nor U6357 (N_6357,N_1525,N_4357);
xnor U6358 (N_6358,N_3279,N_600);
and U6359 (N_6359,N_4512,N_2401);
nand U6360 (N_6360,N_4046,N_4591);
or U6361 (N_6361,N_750,N_782);
nand U6362 (N_6362,N_962,N_4041);
xor U6363 (N_6363,N_2002,N_4336);
or U6364 (N_6364,N_1053,N_2069);
or U6365 (N_6365,N_4730,N_4984);
and U6366 (N_6366,N_771,N_3713);
or U6367 (N_6367,N_1822,N_4624);
or U6368 (N_6368,N_2527,N_4912);
nor U6369 (N_6369,N_3916,N_605);
nor U6370 (N_6370,N_3299,N_4534);
nor U6371 (N_6371,N_4757,N_179);
and U6372 (N_6372,N_3790,N_1357);
xor U6373 (N_6373,N_2522,N_1173);
and U6374 (N_6374,N_1614,N_2867);
nor U6375 (N_6375,N_1967,N_2177);
and U6376 (N_6376,N_2143,N_3798);
nor U6377 (N_6377,N_3672,N_2874);
and U6378 (N_6378,N_2346,N_1287);
or U6379 (N_6379,N_3034,N_4017);
and U6380 (N_6380,N_1081,N_1010);
nand U6381 (N_6381,N_4520,N_598);
and U6382 (N_6382,N_4238,N_15);
nand U6383 (N_6383,N_2149,N_4230);
or U6384 (N_6384,N_2836,N_1845);
nand U6385 (N_6385,N_219,N_728);
and U6386 (N_6386,N_3860,N_1453);
nand U6387 (N_6387,N_3376,N_4903);
xnor U6388 (N_6388,N_1437,N_1828);
or U6389 (N_6389,N_1206,N_2636);
xnor U6390 (N_6390,N_4740,N_2375);
or U6391 (N_6391,N_2004,N_1667);
and U6392 (N_6392,N_2653,N_1382);
nor U6393 (N_6393,N_243,N_2830);
nor U6394 (N_6394,N_886,N_1871);
nor U6395 (N_6395,N_2606,N_1135);
or U6396 (N_6396,N_3501,N_2054);
nor U6397 (N_6397,N_4526,N_3421);
nor U6398 (N_6398,N_230,N_2020);
nor U6399 (N_6399,N_3652,N_2589);
nand U6400 (N_6400,N_4668,N_3693);
or U6401 (N_6401,N_276,N_267);
or U6402 (N_6402,N_1668,N_684);
nor U6403 (N_6403,N_4982,N_3428);
or U6404 (N_6404,N_3180,N_4120);
nor U6405 (N_6405,N_2462,N_102);
or U6406 (N_6406,N_252,N_4260);
or U6407 (N_6407,N_3834,N_1288);
nor U6408 (N_6408,N_666,N_383);
nor U6409 (N_6409,N_1110,N_3032);
or U6410 (N_6410,N_4882,N_4370);
nand U6411 (N_6411,N_154,N_2640);
nor U6412 (N_6412,N_17,N_3741);
xnor U6413 (N_6413,N_4850,N_4823);
and U6414 (N_6414,N_1992,N_939);
and U6415 (N_6415,N_2563,N_2240);
nor U6416 (N_6416,N_2219,N_3618);
or U6417 (N_6417,N_4686,N_505);
and U6418 (N_6418,N_3089,N_3572);
nand U6419 (N_6419,N_2868,N_2615);
and U6420 (N_6420,N_414,N_3529);
nand U6421 (N_6421,N_3950,N_4799);
nor U6422 (N_6422,N_3857,N_204);
nor U6423 (N_6423,N_2344,N_2292);
nor U6424 (N_6424,N_2827,N_1024);
and U6425 (N_6425,N_4954,N_1766);
nor U6426 (N_6426,N_690,N_3630);
nor U6427 (N_6427,N_2657,N_507);
nor U6428 (N_6428,N_3255,N_2483);
nor U6429 (N_6429,N_2897,N_3858);
or U6430 (N_6430,N_3357,N_1169);
nor U6431 (N_6431,N_2264,N_4729);
xnor U6432 (N_6432,N_2095,N_2434);
nand U6433 (N_6433,N_916,N_3769);
and U6434 (N_6434,N_4208,N_1142);
nand U6435 (N_6435,N_3206,N_2964);
or U6436 (N_6436,N_2847,N_1342);
and U6437 (N_6437,N_3407,N_2568);
nor U6438 (N_6438,N_1906,N_9);
nor U6439 (N_6439,N_4815,N_2495);
nand U6440 (N_6440,N_2254,N_2035);
nor U6441 (N_6441,N_570,N_2266);
or U6442 (N_6442,N_4179,N_2108);
nor U6443 (N_6443,N_215,N_3311);
nor U6444 (N_6444,N_3829,N_2623);
or U6445 (N_6445,N_2668,N_1442);
nor U6446 (N_6446,N_2855,N_3371);
or U6447 (N_6447,N_170,N_2100);
and U6448 (N_6448,N_1769,N_2188);
or U6449 (N_6449,N_4401,N_4310);
xor U6450 (N_6450,N_4528,N_1593);
and U6451 (N_6451,N_2913,N_1055);
nor U6452 (N_6452,N_1721,N_197);
nor U6453 (N_6453,N_4206,N_4474);
and U6454 (N_6454,N_56,N_1267);
or U6455 (N_6455,N_4900,N_1727);
or U6456 (N_6456,N_4194,N_3576);
or U6457 (N_6457,N_1176,N_1797);
nand U6458 (N_6458,N_1714,N_905);
nand U6459 (N_6459,N_3913,N_4225);
nand U6460 (N_6460,N_4050,N_428);
xnor U6461 (N_6461,N_918,N_2835);
nor U6462 (N_6462,N_890,N_2549);
nand U6463 (N_6463,N_1284,N_734);
nand U6464 (N_6464,N_824,N_177);
nand U6465 (N_6465,N_4392,N_3704);
nand U6466 (N_6466,N_2920,N_899);
nand U6467 (N_6467,N_3749,N_2574);
nand U6468 (N_6468,N_4025,N_1268);
and U6469 (N_6469,N_625,N_1374);
or U6470 (N_6470,N_2259,N_1383);
and U6471 (N_6471,N_3562,N_101);
and U6472 (N_6472,N_4063,N_3024);
and U6473 (N_6473,N_2681,N_2082);
nor U6474 (N_6474,N_760,N_4342);
nor U6475 (N_6475,N_679,N_1776);
nand U6476 (N_6476,N_4864,N_1677);
nor U6477 (N_6477,N_3645,N_3381);
or U6478 (N_6478,N_3230,N_3696);
nand U6479 (N_6479,N_1059,N_192);
and U6480 (N_6480,N_2933,N_2457);
and U6481 (N_6481,N_1555,N_1231);
nor U6482 (N_6482,N_4935,N_3565);
xor U6483 (N_6483,N_2342,N_2366);
nand U6484 (N_6484,N_1106,N_2270);
and U6485 (N_6485,N_393,N_4015);
nor U6486 (N_6486,N_2310,N_1565);
or U6487 (N_6487,N_4580,N_3772);
nor U6488 (N_6488,N_4229,N_4502);
and U6489 (N_6489,N_1875,N_40);
and U6490 (N_6490,N_1927,N_199);
nand U6491 (N_6491,N_3859,N_449);
nand U6492 (N_6492,N_1103,N_1602);
or U6493 (N_6493,N_3193,N_4691);
nor U6494 (N_6494,N_2598,N_3253);
or U6495 (N_6495,N_37,N_4082);
nor U6496 (N_6496,N_4434,N_2764);
and U6497 (N_6497,N_991,N_4589);
and U6498 (N_6498,N_4347,N_4463);
nand U6499 (N_6499,N_2336,N_1096);
and U6500 (N_6500,N_707,N_2557);
or U6501 (N_6501,N_3793,N_2942);
and U6502 (N_6502,N_171,N_1456);
nor U6503 (N_6503,N_903,N_4365);
and U6504 (N_6504,N_2632,N_913);
nand U6505 (N_6505,N_1915,N_4521);
and U6506 (N_6506,N_4218,N_2768);
nor U6507 (N_6507,N_2395,N_1793);
or U6508 (N_6508,N_429,N_436);
nor U6509 (N_6509,N_4899,N_1030);
nor U6510 (N_6510,N_1092,N_1304);
nand U6511 (N_6511,N_1134,N_1870);
nand U6512 (N_6512,N_3043,N_2829);
nor U6513 (N_6513,N_3519,N_1139);
nand U6514 (N_6514,N_2627,N_2426);
nor U6515 (N_6515,N_3742,N_2513);
and U6516 (N_6516,N_931,N_3734);
nor U6517 (N_6517,N_472,N_3908);
or U6518 (N_6518,N_2614,N_1835);
nand U6519 (N_6519,N_4965,N_2073);
or U6520 (N_6520,N_3315,N_4561);
nand U6521 (N_6521,N_1901,N_4870);
nor U6522 (N_6522,N_2129,N_945);
and U6523 (N_6523,N_4464,N_4069);
and U6524 (N_6524,N_3308,N_4195);
nand U6525 (N_6525,N_4504,N_2110);
nand U6526 (N_6526,N_2419,N_4324);
nand U6527 (N_6527,N_910,N_2032);
or U6528 (N_6528,N_1988,N_1077);
xor U6529 (N_6529,N_1121,N_1584);
and U6530 (N_6530,N_2605,N_2196);
or U6531 (N_6531,N_3597,N_1414);
nand U6532 (N_6532,N_4824,N_2221);
and U6533 (N_6533,N_4621,N_4979);
nor U6534 (N_6534,N_2343,N_3480);
and U6535 (N_6535,N_3240,N_2215);
nor U6536 (N_6536,N_2854,N_1065);
nor U6537 (N_6537,N_4992,N_4196);
nand U6538 (N_6538,N_2372,N_3324);
nand U6539 (N_6539,N_418,N_2862);
nor U6540 (N_6540,N_1956,N_4648);
nand U6541 (N_6541,N_1076,N_1197);
nor U6542 (N_6542,N_3322,N_3220);
and U6543 (N_6543,N_4770,N_1500);
nor U6544 (N_6544,N_1831,N_3609);
nand U6545 (N_6545,N_1323,N_1434);
nor U6546 (N_6546,N_2649,N_4830);
and U6547 (N_6547,N_1291,N_64);
nand U6548 (N_6548,N_2063,N_1515);
nand U6549 (N_6549,N_1025,N_4043);
or U6550 (N_6550,N_1509,N_2226);
or U6551 (N_6551,N_856,N_3161);
nor U6552 (N_6552,N_82,N_561);
or U6553 (N_6553,N_3140,N_1469);
xor U6554 (N_6554,N_1496,N_4858);
nand U6555 (N_6555,N_63,N_4146);
and U6556 (N_6556,N_652,N_1049);
and U6557 (N_6557,N_2971,N_2484);
and U6558 (N_6558,N_4479,N_2837);
and U6559 (N_6559,N_1671,N_4725);
nand U6560 (N_6560,N_3762,N_1402);
xnor U6561 (N_6561,N_303,N_3626);
and U6562 (N_6562,N_1964,N_4084);
or U6563 (N_6563,N_2881,N_3874);
and U6564 (N_6564,N_2579,N_4396);
and U6565 (N_6565,N_2402,N_618);
nand U6566 (N_6566,N_1226,N_1903);
xor U6567 (N_6567,N_4838,N_3835);
nand U6568 (N_6568,N_1066,N_3887);
and U6569 (N_6569,N_3883,N_3848);
nor U6570 (N_6570,N_2425,N_2849);
or U6571 (N_6571,N_4884,N_2772);
nand U6572 (N_6572,N_4647,N_4371);
and U6573 (N_6573,N_908,N_4410);
nor U6574 (N_6574,N_2569,N_4641);
or U6575 (N_6575,N_1375,N_836);
or U6576 (N_6576,N_2338,N_1419);
or U6577 (N_6577,N_4573,N_2601);
or U6578 (N_6578,N_4263,N_1007);
or U6579 (N_6579,N_3685,N_3373);
xnor U6580 (N_6580,N_1928,N_3137);
and U6581 (N_6581,N_394,N_4329);
nor U6582 (N_6582,N_4997,N_2946);
nand U6583 (N_6583,N_3986,N_2269);
and U6584 (N_6584,N_3094,N_745);
or U6585 (N_6585,N_2350,N_1306);
and U6586 (N_6586,N_1975,N_1031);
nand U6587 (N_6587,N_3409,N_1800);
or U6588 (N_6588,N_4999,N_552);
nor U6589 (N_6589,N_3959,N_25);
or U6590 (N_6590,N_3680,N_3869);
and U6591 (N_6591,N_4971,N_4333);
nand U6592 (N_6592,N_1390,N_227);
and U6593 (N_6593,N_1436,N_246);
nor U6594 (N_6594,N_873,N_1008);
nor U6595 (N_6595,N_318,N_3463);
nand U6596 (N_6596,N_4446,N_4762);
or U6597 (N_6597,N_3534,N_1253);
nor U6598 (N_6598,N_3910,N_1128);
nand U6599 (N_6599,N_4564,N_3996);
and U6600 (N_6600,N_1833,N_164);
nor U6601 (N_6601,N_3060,N_4367);
nor U6602 (N_6602,N_617,N_160);
or U6603 (N_6603,N_4759,N_4760);
xor U6604 (N_6604,N_3898,N_2464);
or U6605 (N_6605,N_4003,N_4276);
nor U6606 (N_6606,N_3812,N_2197);
nand U6607 (N_6607,N_2306,N_1421);
or U6608 (N_6608,N_3378,N_4951);
nand U6609 (N_6609,N_3482,N_2114);
and U6610 (N_6610,N_4259,N_3172);
and U6611 (N_6611,N_1449,N_1838);
nand U6612 (N_6612,N_482,N_4373);
nand U6613 (N_6613,N_4450,N_534);
nor U6614 (N_6614,N_4135,N_953);
xnor U6615 (N_6615,N_3002,N_2787);
or U6616 (N_6616,N_1626,N_4507);
or U6617 (N_6617,N_1325,N_648);
nor U6618 (N_6618,N_2194,N_1337);
or U6619 (N_6619,N_4859,N_4630);
nand U6620 (N_6620,N_2472,N_3156);
nor U6621 (N_6621,N_1996,N_4339);
xnor U6622 (N_6622,N_634,N_4245);
or U6623 (N_6623,N_2059,N_1215);
or U6624 (N_6624,N_1234,N_4226);
nor U6625 (N_6625,N_330,N_279);
or U6626 (N_6626,N_4538,N_465);
or U6627 (N_6627,N_1380,N_4519);
or U6628 (N_6628,N_1537,N_4343);
and U6629 (N_6629,N_4675,N_533);
nor U6630 (N_6630,N_3347,N_1596);
or U6631 (N_6631,N_1662,N_331);
or U6632 (N_6632,N_1827,N_4578);
nand U6633 (N_6633,N_2717,N_4293);
and U6634 (N_6634,N_4642,N_3684);
or U6635 (N_6635,N_2206,N_2546);
or U6636 (N_6636,N_2179,N_4714);
nor U6637 (N_6637,N_2238,N_1352);
nor U6638 (N_6638,N_881,N_1433);
or U6639 (N_6639,N_1191,N_1309);
or U6640 (N_6640,N_915,N_504);
nor U6641 (N_6641,N_3820,N_970);
and U6642 (N_6642,N_1877,N_563);
and U6643 (N_6643,N_2377,N_4298);
or U6644 (N_6644,N_4736,N_4004);
nor U6645 (N_6645,N_300,N_2877);
nor U6646 (N_6646,N_1786,N_2291);
nand U6647 (N_6647,N_1539,N_867);
nand U6648 (N_6648,N_969,N_362);
or U6649 (N_6649,N_4755,N_1807);
nand U6650 (N_6650,N_2555,N_4685);
and U6651 (N_6651,N_4448,N_1270);
or U6652 (N_6652,N_4119,N_4607);
and U6653 (N_6653,N_1431,N_657);
nor U6654 (N_6654,N_4109,N_1295);
and U6655 (N_6655,N_4827,N_784);
or U6656 (N_6656,N_4758,N_2386);
nor U6657 (N_6657,N_2734,N_3264);
xnor U6658 (N_6658,N_4896,N_1427);
nor U6659 (N_6659,N_371,N_3398);
and U6660 (N_6660,N_4711,N_912);
nor U6661 (N_6661,N_4214,N_1332);
nor U6662 (N_6662,N_2526,N_441);
or U6663 (N_6663,N_4007,N_1837);
and U6664 (N_6664,N_4096,N_3261);
nor U6665 (N_6665,N_3168,N_2118);
or U6666 (N_6666,N_4187,N_3029);
and U6667 (N_6667,N_951,N_1990);
nand U6668 (N_6668,N_495,N_3169);
and U6669 (N_6669,N_2960,N_1730);
nor U6670 (N_6670,N_693,N_61);
nand U6671 (N_6671,N_216,N_1283);
nor U6672 (N_6672,N_1995,N_2638);
or U6673 (N_6673,N_4889,N_642);
or U6674 (N_6674,N_2882,N_1907);
nor U6675 (N_6675,N_1086,N_3123);
nand U6676 (N_6676,N_3474,N_878);
nor U6677 (N_6677,N_2151,N_701);
or U6678 (N_6678,N_4056,N_3015);
and U6679 (N_6679,N_4892,N_4447);
and U6680 (N_6680,N_424,N_4545);
nor U6681 (N_6681,N_702,N_2481);
nor U6682 (N_6682,N_3307,N_2262);
or U6683 (N_6683,N_3854,N_1937);
and U6684 (N_6684,N_3683,N_2448);
nand U6685 (N_6685,N_321,N_2703);
nor U6686 (N_6686,N_3540,N_2081);
nand U6687 (N_6687,N_1898,N_3511);
and U6688 (N_6688,N_2046,N_4877);
nor U6689 (N_6689,N_2115,N_1023);
nand U6690 (N_6690,N_273,N_1276);
and U6691 (N_6691,N_3290,N_1979);
or U6692 (N_6692,N_1365,N_304);
nand U6693 (N_6693,N_4744,N_2515);
nor U6694 (N_6694,N_3699,N_4518);
and U6695 (N_6695,N_3040,N_2828);
or U6696 (N_6696,N_621,N_499);
and U6697 (N_6697,N_4885,N_3186);
or U6698 (N_6698,N_396,N_2607);
or U6699 (N_6699,N_1420,N_1576);
xor U6700 (N_6700,N_1653,N_583);
nand U6701 (N_6701,N_2331,N_2884);
nor U6702 (N_6702,N_450,N_861);
or U6703 (N_6703,N_3987,N_1497);
xnor U6704 (N_6704,N_2924,N_2593);
nand U6705 (N_6705,N_2600,N_1014);
and U6706 (N_6706,N_2542,N_1520);
nor U6707 (N_6707,N_1854,N_2644);
nor U6708 (N_6708,N_1813,N_855);
nand U6709 (N_6709,N_1731,N_2090);
nand U6710 (N_6710,N_4475,N_419);
or U6711 (N_6711,N_3621,N_4623);
nand U6712 (N_6712,N_4061,N_2630);
and U6713 (N_6713,N_3465,N_3492);
or U6714 (N_6714,N_41,N_3329);
nand U6715 (N_6715,N_60,N_1333);
xnor U6716 (N_6716,N_2022,N_3884);
or U6717 (N_6717,N_2192,N_1852);
and U6718 (N_6718,N_3810,N_4022);
nor U6719 (N_6719,N_4679,N_4482);
or U6720 (N_6720,N_3195,N_4550);
nor U6721 (N_6721,N_264,N_4044);
nand U6722 (N_6722,N_843,N_187);
nand U6723 (N_6723,N_703,N_4509);
nand U6724 (N_6724,N_4913,N_4794);
nor U6725 (N_6725,N_4190,N_2656);
and U6726 (N_6726,N_4246,N_3634);
or U6727 (N_6727,N_2450,N_3362);
nand U6728 (N_6728,N_1044,N_1261);
nor U6729 (N_6729,N_4494,N_2988);
nor U6730 (N_6730,N_4493,N_4839);
nand U6731 (N_6731,N_3881,N_3247);
nor U6732 (N_6732,N_3780,N_4592);
nor U6733 (N_6733,N_955,N_3896);
and U6734 (N_6734,N_1759,N_2671);
nand U6735 (N_6735,N_1665,N_3994);
nand U6736 (N_6736,N_3682,N_4098);
and U6737 (N_6737,N_1376,N_3851);
and U6738 (N_6738,N_3679,N_3776);
nor U6739 (N_6739,N_1717,N_4024);
and U6740 (N_6740,N_1765,N_2762);
nand U6741 (N_6741,N_3736,N_1240);
nand U6742 (N_6742,N_655,N_706);
nand U6743 (N_6743,N_3053,N_1422);
xnor U6744 (N_6744,N_4956,N_2153);
or U6745 (N_6745,N_698,N_388);
nor U6746 (N_6746,N_1916,N_1666);
nor U6747 (N_6747,N_288,N_4290);
or U6748 (N_6748,N_715,N_186);
nor U6749 (N_6749,N_3723,N_2871);
and U6750 (N_6750,N_3543,N_4522);
nand U6751 (N_6751,N_404,N_4348);
or U6752 (N_6752,N_4223,N_579);
or U6753 (N_6753,N_3243,N_1476);
nand U6754 (N_6754,N_4346,N_146);
nor U6755 (N_6755,N_366,N_3209);
or U6756 (N_6756,N_3028,N_2712);
nand U6757 (N_6757,N_845,N_1508);
or U6758 (N_6758,N_3671,N_3201);
nor U6759 (N_6759,N_4855,N_2301);
nor U6760 (N_6760,N_1199,N_4467);
or U6761 (N_6761,N_308,N_774);
or U6762 (N_6762,N_4646,N_4911);
and U6763 (N_6763,N_4922,N_3978);
nor U6764 (N_6764,N_2519,N_150);
and U6765 (N_6765,N_3424,N_645);
nor U6766 (N_6766,N_3900,N_3688);
nor U6767 (N_6767,N_3141,N_1698);
nor U6768 (N_6768,N_3328,N_1467);
nor U6769 (N_6769,N_1767,N_758);
nor U6770 (N_6770,N_4894,N_1439);
or U6771 (N_6771,N_4092,N_2057);
nor U6772 (N_6772,N_4709,N_609);
nand U6773 (N_6773,N_3284,N_3993);
nand U6774 (N_6774,N_2902,N_4689);
and U6775 (N_6775,N_1501,N_1768);
nand U6776 (N_6776,N_275,N_235);
nor U6777 (N_6777,N_1941,N_3152);
and U6778 (N_6778,N_2730,N_2037);
nand U6779 (N_6779,N_1619,N_3917);
or U6780 (N_6780,N_809,N_3774);
and U6781 (N_6781,N_3082,N_3615);
and U6782 (N_6782,N_941,N_565);
or U6783 (N_6783,N_2175,N_4558);
nand U6784 (N_6784,N_3613,N_3174);
or U6785 (N_6785,N_2771,N_1266);
nor U6786 (N_6786,N_2688,N_4147);
and U6787 (N_6787,N_4875,N_2493);
nand U6788 (N_6788,N_3981,N_2832);
or U6789 (N_6789,N_1994,N_4210);
nor U6790 (N_6790,N_847,N_4907);
or U6791 (N_6791,N_2886,N_3312);
and U6792 (N_6792,N_226,N_1541);
or U6793 (N_6793,N_2210,N_2550);
nor U6794 (N_6794,N_932,N_2482);
nand U6795 (N_6795,N_1477,N_2811);
nand U6796 (N_6796,N_205,N_224);
and U6797 (N_6797,N_2586,N_606);
or U6798 (N_6798,N_3250,N_3162);
nand U6799 (N_6799,N_4341,N_3563);
nand U6800 (N_6800,N_2695,N_132);
or U6801 (N_6801,N_3213,N_555);
or U6802 (N_6802,N_352,N_3568);
nand U6803 (N_6803,N_3420,N_182);
or U6804 (N_6804,N_2930,N_3553);
and U6805 (N_6805,N_1563,N_852);
or U6806 (N_6806,N_4667,N_801);
nor U6807 (N_6807,N_323,N_4389);
or U6808 (N_6808,N_3544,N_4432);
nor U6809 (N_6809,N_422,N_3175);
and U6810 (N_6810,N_4093,N_1136);
or U6811 (N_6811,N_4531,N_1570);
and U6812 (N_6812,N_4865,N_4795);
nor U6813 (N_6813,N_1331,N_806);
nor U6814 (N_6814,N_1959,N_2380);
nand U6815 (N_6815,N_1161,N_3267);
nand U6816 (N_6816,N_3918,N_3832);
nand U6817 (N_6817,N_3100,N_4813);
and U6818 (N_6818,N_3283,N_2150);
nand U6819 (N_6819,N_3601,N_4883);
or U6820 (N_6820,N_2072,N_3743);
and U6821 (N_6821,N_1758,N_3342);
nand U6822 (N_6822,N_4064,N_2);
nand U6823 (N_6823,N_3,N_3202);
nor U6824 (N_6824,N_1674,N_4975);
and U6825 (N_6825,N_3922,N_4620);
or U6826 (N_6826,N_3163,N_3745);
nand U6827 (N_6827,N_1400,N_2801);
nand U6828 (N_6828,N_4697,N_4021);
nand U6829 (N_6829,N_1479,N_3395);
nand U6830 (N_6830,N_262,N_4215);
or U6831 (N_6831,N_3587,N_4313);
nand U6832 (N_6832,N_4995,N_826);
and U6833 (N_6833,N_95,N_854);
nor U6834 (N_6834,N_4906,N_3506);
and U6835 (N_6835,N_1109,N_3611);
and U6836 (N_6836,N_1675,N_4107);
and U6837 (N_6837,N_4506,N_3214);
nand U6838 (N_6838,N_3257,N_69);
nand U6839 (N_6839,N_4968,N_2966);
or U6840 (N_6840,N_3827,N_4804);
xnor U6841 (N_6841,N_1865,N_3445);
nor U6842 (N_6842,N_1953,N_511);
or U6843 (N_6843,N_793,N_4189);
nor U6844 (N_6844,N_3556,N_3691);
or U6845 (N_6845,N_4544,N_1446);
nand U6846 (N_6846,N_4515,N_4077);
and U6847 (N_6847,N_4209,N_380);
and U6848 (N_6848,N_458,N_1444);
or U6849 (N_6849,N_935,N_3425);
nand U6850 (N_6850,N_3383,N_440);
and U6851 (N_6851,N_980,N_2547);
xnor U6852 (N_6852,N_140,N_1621);
xnor U6853 (N_6853,N_221,N_640);
nor U6854 (N_6854,N_1213,N_4060);
and U6855 (N_6855,N_3971,N_730);
or U6856 (N_6856,N_2091,N_1917);
and U6857 (N_6857,N_470,N_812);
or U6858 (N_6858,N_2741,N_3788);
nor U6859 (N_6859,N_661,N_1465);
nand U6860 (N_6860,N_3098,N_3905);
nand U6861 (N_6861,N_4001,N_1685);
nand U6862 (N_6862,N_3073,N_1749);
xor U6863 (N_6863,N_445,N_3838);
nand U6864 (N_6864,N_3036,N_4158);
nor U6865 (N_6865,N_3947,N_514);
and U6866 (N_6866,N_4262,N_3103);
nor U6867 (N_6867,N_3919,N_3128);
and U6868 (N_6868,N_1704,N_1156);
and U6869 (N_6869,N_3585,N_4942);
and U6870 (N_6870,N_4140,N_833);
and U6871 (N_6871,N_4715,N_54);
nand U6872 (N_6872,N_1878,N_1775);
nand U6873 (N_6873,N_2231,N_4145);
or U6874 (N_6874,N_24,N_1920);
and U6875 (N_6875,N_1821,N_3879);
or U6876 (N_6876,N_3564,N_3469);
and U6877 (N_6877,N_3061,N_2398);
and U6878 (N_6878,N_2116,N_2951);
or U6879 (N_6879,N_755,N_3786);
and U6880 (N_6880,N_4636,N_4356);
nor U6881 (N_6881,N_241,N_481);
or U6882 (N_6882,N_3139,N_92);
and U6883 (N_6883,N_4927,N_65);
or U6884 (N_6884,N_2692,N_464);
or U6885 (N_6885,N_4270,N_1664);
nor U6886 (N_6886,N_906,N_4533);
nor U6887 (N_6887,N_3044,N_851);
nand U6888 (N_6888,N_3828,N_469);
nor U6889 (N_6889,N_1001,N_2707);
nor U6890 (N_6890,N_4429,N_3569);
nor U6891 (N_6891,N_1810,N_2844);
nand U6892 (N_6892,N_4826,N_3878);
nand U6893 (N_6893,N_1882,N_1474);
or U6894 (N_6894,N_3401,N_1595);
or U6895 (N_6895,N_1393,N_1149);
nand U6896 (N_6896,N_77,N_3961);
xor U6897 (N_6897,N_651,N_3129);
or U6898 (N_6898,N_2136,N_1894);
nand U6899 (N_6899,N_4454,N_4091);
or U6900 (N_6900,N_2067,N_3579);
and U6901 (N_6901,N_4866,N_1876);
nor U6902 (N_6902,N_1011,N_2873);
nand U6903 (N_6903,N_1441,N_3536);
nand U6904 (N_6904,N_4415,N_4536);
or U6905 (N_6905,N_3552,N_129);
or U6906 (N_6906,N_3992,N_4540);
nand U6907 (N_6907,N_2438,N_4065);
nand U6908 (N_6908,N_2876,N_3419);
nand U6909 (N_6909,N_4435,N_3353);
or U6910 (N_6910,N_3761,N_4604);
nor U6911 (N_6911,N_2943,N_2258);
and U6912 (N_6912,N_1181,N_4633);
nand U6913 (N_6913,N_1622,N_2990);
and U6914 (N_6914,N_4891,N_3000);
and U6915 (N_6915,N_448,N_2354);
or U6916 (N_6916,N_611,N_4148);
xnor U6917 (N_6917,N_1533,N_1723);
nand U6918 (N_6918,N_1930,N_2201);
or U6919 (N_6919,N_3042,N_4297);
nor U6920 (N_6920,N_314,N_4283);
or U6921 (N_6921,N_1180,N_2399);
nor U6922 (N_6922,N_573,N_2702);
nand U6923 (N_6923,N_3046,N_720);
nor U6924 (N_6924,N_136,N_1);
nor U6925 (N_6925,N_994,N_3605);
and U6926 (N_6926,N_3448,N_972);
nor U6927 (N_6927,N_2565,N_1661);
nand U6928 (N_6928,N_1003,N_4862);
and U6929 (N_6929,N_3241,N_3360);
nor U6930 (N_6930,N_2160,N_479);
and U6931 (N_6931,N_682,N_530);
and U6932 (N_6932,N_4492,N_467);
or U6933 (N_6933,N_4102,N_1043);
nor U6934 (N_6934,N_952,N_2479);
or U6935 (N_6935,N_2793,N_3813);
or U6936 (N_6936,N_2660,N_623);
and U6937 (N_6937,N_3008,N_1200);
and U6938 (N_6938,N_4023,N_1516);
nand U6939 (N_6939,N_1187,N_2023);
and U6940 (N_6940,N_4936,N_4222);
or U6941 (N_6941,N_208,N_2008);
and U6942 (N_6942,N_2997,N_1120);
nand U6943 (N_6943,N_3084,N_1265);
nand U6944 (N_6944,N_4532,N_8);
or U6945 (N_6945,N_2099,N_2585);
nor U6946 (N_6946,N_291,N_1482);
or U6947 (N_6947,N_966,N_1954);
and U6948 (N_6948,N_3125,N_1140);
nor U6949 (N_6949,N_2751,N_4364);
and U6950 (N_6950,N_1098,N_3822);
and U6951 (N_6951,N_1613,N_4790);
nor U6952 (N_6952,N_517,N_4871);
or U6953 (N_6953,N_560,N_1329);
or U6954 (N_6954,N_343,N_1344);
and U6955 (N_6955,N_4972,N_3296);
and U6956 (N_6956,N_2424,N_4411);
and U6957 (N_6957,N_2388,N_4775);
nor U6958 (N_6958,N_1322,N_2982);
and U6959 (N_6959,N_431,N_2025);
nor U6960 (N_6960,N_1757,N_2888);
xnor U6961 (N_6961,N_3648,N_2573);
and U6962 (N_6962,N_2485,N_1260);
and U6963 (N_6963,N_4438,N_1955);
or U6964 (N_6964,N_58,N_3135);
nand U6965 (N_6965,N_2391,N_2187);
nand U6966 (N_6966,N_3294,N_1560);
nor U6967 (N_6967,N_3192,N_3233);
nand U6968 (N_6968,N_2641,N_2097);
and U6969 (N_6969,N_1377,N_2287);
xnor U6970 (N_6970,N_576,N_4279);
and U6971 (N_6971,N_2089,N_746);
nor U6972 (N_6972,N_807,N_1912);
nand U6973 (N_6973,N_4397,N_1944);
nor U6974 (N_6974,N_677,N_4344);
nor U6975 (N_6975,N_3760,N_3731);
nand U6976 (N_6976,N_2013,N_3012);
and U6977 (N_6977,N_1051,N_3673);
or U6978 (N_6978,N_3006,N_2544);
or U6979 (N_6979,N_2812,N_2387);
nor U6980 (N_6980,N_1741,N_4016);
and U6981 (N_6981,N_2138,N_3852);
or U6982 (N_6982,N_3770,N_3890);
nand U6983 (N_6983,N_4958,N_4074);
nand U6984 (N_6984,N_2959,N_232);
or U6985 (N_6985,N_1895,N_4634);
and U6986 (N_6986,N_3977,N_2693);
and U6987 (N_6987,N_542,N_3594);
nand U6988 (N_6988,N_2135,N_4499);
and U6989 (N_6989,N_3707,N_3873);
nor U6990 (N_6990,N_480,N_791);
or U6991 (N_6991,N_4963,N_4505);
and U6992 (N_6992,N_1071,N_1748);
nand U6993 (N_6993,N_1478,N_1718);
nor U6994 (N_6994,N_663,N_898);
or U6995 (N_6995,N_4352,N_4165);
or U6996 (N_6996,N_1164,N_3184);
and U6997 (N_6997,N_4073,N_2186);
nor U6998 (N_6998,N_1461,N_765);
and U6999 (N_6999,N_2403,N_902);
or U7000 (N_7000,N_1379,N_158);
nor U7001 (N_7001,N_3590,N_4924);
or U7002 (N_7002,N_4027,N_4814);
nor U7003 (N_7003,N_4455,N_3863);
and U7004 (N_7004,N_658,N_3179);
or U7005 (N_7005,N_4385,N_4773);
nand U7006 (N_7006,N_1918,N_2305);
nand U7007 (N_7007,N_2860,N_3026);
nand U7008 (N_7008,N_1763,N_920);
and U7009 (N_7009,N_3413,N_4174);
nor U7010 (N_7010,N_1099,N_3111);
and U7011 (N_7011,N_4138,N_4988);
and U7012 (N_7012,N_3888,N_3126);
or U7013 (N_7013,N_358,N_3990);
and U7014 (N_7014,N_3091,N_2878);
nor U7015 (N_7015,N_3711,N_379);
and U7016 (N_7016,N_896,N_3748);
nor U7017 (N_7017,N_3239,N_2631);
or U7018 (N_7018,N_3116,N_2909);
or U7019 (N_7019,N_2780,N_2826);
nor U7020 (N_7020,N_3016,N_516);
nor U7021 (N_7021,N_3604,N_223);
nor U7022 (N_7022,N_795,N_4072);
nand U7023 (N_7023,N_2314,N_3567);
or U7024 (N_7024,N_3256,N_3757);
or U7025 (N_7025,N_32,N_4766);
or U7026 (N_7026,N_2311,N_2898);
nor U7027 (N_7027,N_4085,N_111);
nor U7028 (N_7028,N_4719,N_1155);
or U7029 (N_7029,N_1558,N_2455);
and U7030 (N_7030,N_4167,N_2246);
or U7031 (N_7031,N_4380,N_3439);
nor U7032 (N_7032,N_3071,N_1538);
xnor U7033 (N_7033,N_2530,N_880);
nand U7034 (N_7034,N_3725,N_1531);
or U7035 (N_7035,N_4217,N_1726);
and U7036 (N_7036,N_4216,N_2183);
nor U7037 (N_7037,N_1016,N_1976);
or U7038 (N_7038,N_4452,N_2337);
nand U7039 (N_7039,N_2500,N_2891);
or U7040 (N_7040,N_4703,N_2356);
and U7041 (N_7041,N_4792,N_1562);
nand U7042 (N_7042,N_925,N_3606);
or U7043 (N_7043,N_4683,N_2474);
or U7044 (N_7044,N_485,N_30);
nor U7045 (N_7045,N_4250,N_993);
and U7046 (N_7046,N_914,N_385);
and U7047 (N_7047,N_4739,N_1356);
xnor U7048 (N_7048,N_1241,N_2760);
or U7049 (N_7049,N_4420,N_2282);
and U7050 (N_7050,N_489,N_3706);
or U7051 (N_7051,N_3666,N_202);
nor U7052 (N_7052,N_3647,N_4807);
and U7053 (N_7053,N_749,N_564);
and U7054 (N_7054,N_2561,N_74);
nand U7055 (N_7055,N_1182,N_1715);
or U7056 (N_7056,N_2710,N_2932);
nor U7057 (N_7057,N_1630,N_4466);
and U7058 (N_7058,N_2404,N_1026);
and U7059 (N_7059,N_497,N_271);
nor U7060 (N_7060,N_2694,N_4684);
or U7061 (N_7061,N_2289,N_3164);
and U7062 (N_7062,N_447,N_370);
and U7063 (N_7063,N_543,N_2026);
nand U7064 (N_7064,N_1070,N_3639);
nand U7065 (N_7065,N_1364,N_2551);
and U7066 (N_7066,N_769,N_335);
and U7067 (N_7067,N_2813,N_2864);
nand U7068 (N_7068,N_1973,N_4427);
and U7069 (N_7069,N_1946,N_2859);
or U7070 (N_7070,N_584,N_2973);
and U7071 (N_7071,N_285,N_189);
nand U7072 (N_7072,N_4837,N_1117);
nand U7073 (N_7073,N_1102,N_4886);
and U7074 (N_7074,N_3148,N_2865);
and U7075 (N_7075,N_865,N_4880);
nor U7076 (N_7076,N_3928,N_3191);
nor U7077 (N_7077,N_4549,N_768);
nor U7078 (N_7078,N_1127,N_2260);
and U7079 (N_7079,N_2570,N_2845);
and U7080 (N_7080,N_2180,N_3216);
and U7081 (N_7081,N_3022,N_4706);
and U7082 (N_7082,N_363,N_3649);
nand U7083 (N_7083,N_4202,N_4919);
and U7084 (N_7084,N_1743,N_2838);
nor U7085 (N_7085,N_2749,N_1651);
nor U7086 (N_7086,N_2315,N_3093);
nand U7087 (N_7087,N_97,N_2883);
nand U7088 (N_7088,N_2461,N_649);
and U7089 (N_7089,N_4354,N_3722);
nand U7090 (N_7090,N_116,N_3068);
nor U7091 (N_7091,N_1062,N_4075);
nand U7092 (N_7092,N_984,N_2120);
nand U7093 (N_7093,N_968,N_4618);
nand U7094 (N_7094,N_3899,N_3510);
or U7095 (N_7095,N_804,N_3466);
xnor U7096 (N_7096,N_4752,N_3114);
or U7097 (N_7097,N_4005,N_4040);
nor U7098 (N_7098,N_4611,N_1194);
or U7099 (N_7099,N_2992,N_3789);
nor U7100 (N_7100,N_3363,N_540);
nand U7101 (N_7101,N_1779,N_1301);
or U7102 (N_7102,N_3518,N_4291);
and U7103 (N_7103,N_2340,N_1150);
or U7104 (N_7104,N_2367,N_1488);
and U7105 (N_7105,N_1519,N_3498);
nor U7106 (N_7106,N_1683,N_1114);
and U7107 (N_7107,N_4655,N_355);
and U7108 (N_7108,N_2517,N_4610);
or U7109 (N_7109,N_1313,N_2682);
or U7110 (N_7110,N_2191,N_4111);
nand U7111 (N_7111,N_3687,N_1860);
nor U7112 (N_7112,N_26,N_27);
nor U7113 (N_7113,N_2564,N_2648);
and U7114 (N_7114,N_2595,N_159);
and U7115 (N_7115,N_4381,N_3937);
nor U7116 (N_7116,N_1335,N_4609);
and U7117 (N_7117,N_686,N_1536);
or U7118 (N_7118,N_1087,N_1716);
and U7119 (N_7119,N_2393,N_4802);
nor U7120 (N_7120,N_1559,N_4284);
nor U7121 (N_7121,N_940,N_4379);
nand U7122 (N_7122,N_4970,N_3787);
or U7123 (N_7123,N_1960,N_2133);
nand U7124 (N_7124,N_1264,N_2249);
or U7125 (N_7125,N_2857,N_2442);
or U7126 (N_7126,N_3442,N_2036);
and U7127 (N_7127,N_2962,N_244);
or U7128 (N_7128,N_3077,N_2658);
and U7129 (N_7129,N_2252,N_3847);
and U7130 (N_7130,N_1233,N_2412);
nor U7131 (N_7131,N_1796,N_2892);
and U7132 (N_7132,N_3499,N_957);
and U7133 (N_7133,N_3165,N_3531);
nor U7134 (N_7134,N_4300,N_4055);
nor U7135 (N_7135,N_4058,N_284);
nor U7136 (N_7136,N_4244,N_3709);
nor U7137 (N_7137,N_3980,N_4832);
and U7138 (N_7138,N_992,N_112);
nand U7139 (N_7139,N_3599,N_3885);
nand U7140 (N_7140,N_4049,N_2286);
nand U7141 (N_7141,N_3320,N_2948);
nor U7142 (N_7142,N_1154,N_1591);
nand U7143 (N_7143,N_742,N_2321);
or U7144 (N_7144,N_2307,N_4681);
nand U7145 (N_7145,N_4274,N_233);
nor U7146 (N_7146,N_654,N_353);
nor U7147 (N_7147,N_2825,N_4481);
or U7148 (N_7148,N_3850,N_200);
or U7149 (N_7149,N_1248,N_2802);
and U7150 (N_7150,N_2101,N_3210);
or U7151 (N_7151,N_319,N_3153);
nand U7152 (N_7152,N_3646,N_3288);
or U7153 (N_7153,N_2432,N_3352);
and U7154 (N_7154,N_2157,N_3158);
nor U7155 (N_7155,N_797,N_3738);
and U7156 (N_7156,N_3289,N_2726);
xor U7157 (N_7157,N_3429,N_4973);
or U7158 (N_7158,N_3323,N_1923);
or U7159 (N_7159,N_3414,N_4271);
or U7160 (N_7160,N_277,N_4551);
nor U7161 (N_7161,N_636,N_53);
nand U7162 (N_7162,N_3285,N_4168);
and U7163 (N_7163,N_4785,N_2936);
and U7164 (N_7164,N_2524,N_1691);
or U7165 (N_7165,N_2678,N_588);
or U7166 (N_7166,N_4353,N_3030);
nor U7167 (N_7167,N_1707,N_1789);
nor U7168 (N_7168,N_2416,N_4867);
nand U7169 (N_7169,N_3274,N_2440);
nand U7170 (N_7170,N_4419,N_274);
xor U7171 (N_7171,N_770,N_4282);
nand U7172 (N_7172,N_3903,N_1607);
nor U7173 (N_7173,N_4543,N_4571);
nor U7174 (N_7174,N_2132,N_2577);
xnor U7175 (N_7175,N_764,N_4733);
or U7176 (N_7176,N_3792,N_3494);
nand U7177 (N_7177,N_2511,N_4556);
and U7178 (N_7178,N_1858,N_3960);
and U7179 (N_7179,N_1122,N_3484);
and U7180 (N_7180,N_1606,N_2995);
nand U7181 (N_7181,N_4241,N_3070);
nor U7182 (N_7182,N_84,N_4663);
nor U7183 (N_7183,N_1277,N_4160);
nor U7184 (N_7184,N_3833,N_3403);
and U7185 (N_7185,N_2599,N_2518);
nor U7186 (N_7186,N_4656,N_4201);
and U7187 (N_7187,N_2590,N_4062);
nand U7188 (N_7188,N_1388,N_103);
nor U7189 (N_7189,N_4660,N_3248);
or U7190 (N_7190,N_1440,N_42);
and U7191 (N_7191,N_2869,N_2335);
nand U7192 (N_7192,N_2918,N_2970);
and U7193 (N_7193,N_1229,N_443);
and U7194 (N_7194,N_2413,N_4089);
nor U7195 (N_7195,N_562,N_1318);
nand U7196 (N_7196,N_1489,N_3582);
nand U7197 (N_7197,N_2512,N_956);
nand U7198 (N_7198,N_1485,N_3686);
nor U7199 (N_7199,N_4117,N_4712);
nor U7200 (N_7200,N_4296,N_1738);
nor U7201 (N_7201,N_4067,N_4878);
nand U7202 (N_7202,N_3720,N_3119);
nor U7203 (N_7203,N_4915,N_337);
nor U7204 (N_7204,N_4635,N_4236);
nand U7205 (N_7205,N_4511,N_3096);
and U7206 (N_7206,N_1397,N_332);
nor U7207 (N_7207,N_2295,N_864);
nor U7208 (N_7208,N_2146,N_1481);
nor U7209 (N_7209,N_13,N_2818);
nand U7210 (N_7210,N_3570,N_4833);
nand U7211 (N_7211,N_1308,N_2977);
nor U7212 (N_7212,N_1320,N_4750);
nor U7213 (N_7213,N_643,N_459);
nand U7214 (N_7214,N_456,N_4264);
or U7215 (N_7215,N_3048,N_4812);
nor U7216 (N_7216,N_1262,N_1545);
or U7217 (N_7217,N_3367,N_3991);
or U7218 (N_7218,N_3807,N_1138);
or U7219 (N_7219,N_3190,N_4288);
or U7220 (N_7220,N_3867,N_4929);
nand U7221 (N_7221,N_1450,N_1404);
and U7222 (N_7222,N_2680,N_3951);
xnor U7223 (N_7223,N_3670,N_4612);
nand U7224 (N_7224,N_2410,N_3221);
nor U7225 (N_7225,N_3385,N_4945);
or U7226 (N_7226,N_2504,N_1527);
nor U7227 (N_7227,N_2914,N_1068);
nand U7228 (N_7228,N_2711,N_4388);
or U7229 (N_7229,N_3170,N_1487);
or U7230 (N_7230,N_2200,N_4421);
or U7231 (N_7231,N_710,N_1728);
or U7232 (N_7232,N_4674,N_3877);
nor U7233 (N_7233,N_711,N_4294);
or U7234 (N_7234,N_3346,N_3305);
nand U7235 (N_7235,N_846,N_340);
and U7236 (N_7236,N_2810,N_3497);
nor U7237 (N_7237,N_1475,N_2759);
nand U7238 (N_7238,N_4688,N_1328);
or U7239 (N_7239,N_247,N_3487);
and U7240 (N_7240,N_513,N_2006);
nor U7241 (N_7241,N_2447,N_364);
xor U7242 (N_7242,N_2480,N_2024);
or U7243 (N_7243,N_3332,N_1971);
nor U7244 (N_7244,N_4879,N_3985);
or U7245 (N_7245,N_4933,N_2383);
or U7246 (N_7246,N_538,N_1580);
and U7247 (N_7247,N_798,N_3228);
or U7248 (N_7248,N_2428,N_1466);
or U7249 (N_7249,N_4249,N_4694);
nor U7250 (N_7250,N_2926,N_4994);
nand U7251 (N_7251,N_1658,N_4572);
nand U7252 (N_7252,N_1819,N_1242);
or U7253 (N_7253,N_2117,N_2496);
or U7254 (N_7254,N_1341,N_2505);
nand U7255 (N_7255,N_31,N_2798);
nand U7256 (N_7256,N_2297,N_1709);
nor U7257 (N_7257,N_3824,N_591);
and U7258 (N_7258,N_3147,N_1491);
nand U7259 (N_7259,N_3101,N_3726);
and U7260 (N_7260,N_4659,N_312);
or U7261 (N_7261,N_582,N_789);
and U7262 (N_7262,N_4704,N_1840);
nor U7263 (N_7263,N_4486,N_3017);
or U7264 (N_7264,N_1188,N_181);
nor U7265 (N_7265,N_130,N_2554);
and U7266 (N_7266,N_2339,N_4993);
or U7267 (N_7267,N_1246,N_1435);
or U7268 (N_7268,N_936,N_1228);
xnor U7269 (N_7269,N_3598,N_4081);
and U7270 (N_7270,N_4854,N_1370);
or U7271 (N_7271,N_148,N_1868);
nand U7272 (N_7272,N_4613,N_4763);
or U7273 (N_7273,N_3927,N_2732);
and U7274 (N_7274,N_3791,N_4157);
nand U7275 (N_7275,N_3495,N_4255);
nand U7276 (N_7276,N_1311,N_2708);
nor U7277 (N_7277,N_3259,N_3208);
nor U7278 (N_7278,N_3075,N_203);
and U7279 (N_7279,N_4649,N_1165);
nand U7280 (N_7280,N_3423,N_2594);
or U7281 (N_7281,N_948,N_1385);
and U7282 (N_7282,N_1239,N_432);
or U7283 (N_7283,N_696,N_601);
and U7284 (N_7284,N_3653,N_4399);
or U7285 (N_7285,N_269,N_494);
and U7286 (N_7286,N_4923,N_2916);
nor U7287 (N_7287,N_3988,N_876);
and U7288 (N_7288,N_3348,N_592);
and U7289 (N_7289,N_1581,N_4843);
nand U7290 (N_7290,N_4425,N_4378);
nand U7291 (N_7291,N_1372,N_483);
nor U7292 (N_7292,N_828,N_2795);
and U7293 (N_7293,N_1947,N_4273);
or U7294 (N_7294,N_1060,N_3010);
nor U7295 (N_7295,N_1314,N_3155);
nand U7296 (N_7296,N_3197,N_4943);
nand U7297 (N_7297,N_1805,N_3159);
or U7298 (N_7298,N_2906,N_4593);
nor U7299 (N_7299,N_4939,N_4039);
nor U7300 (N_7300,N_4876,N_118);
or U7301 (N_7301,N_2470,N_3698);
nor U7302 (N_7302,N_3504,N_2453);
and U7303 (N_7303,N_2327,N_4422);
and U7304 (N_7304,N_3512,N_3936);
nor U7305 (N_7305,N_595,N_2014);
or U7306 (N_7306,N_3644,N_2506);
and U7307 (N_7307,N_2427,N_3515);
or U7308 (N_7308,N_2769,N_2541);
nor U7309 (N_7309,N_110,N_4417);
nand U7310 (N_7310,N_3909,N_4863);
or U7311 (N_7311,N_1005,N_587);
nand U7312 (N_7312,N_2961,N_3379);
nand U7313 (N_7313,N_3623,N_4756);
nor U7314 (N_7314,N_761,N_2454);
nor U7315 (N_7315,N_3080,N_4152);
nand U7316 (N_7316,N_3819,N_889);
nand U7317 (N_7317,N_3078,N_2435);
nand U7318 (N_7318,N_293,N_975);
nor U7319 (N_7319,N_167,N_426);
or U7320 (N_7320,N_3189,N_2174);
nor U7321 (N_7321,N_777,N_1746);
and U7322 (N_7322,N_2775,N_1058);
nand U7323 (N_7323,N_2332,N_280);
or U7324 (N_7324,N_3455,N_3035);
and U7325 (N_7325,N_1143,N_1015);
or U7326 (N_7326,N_1997,N_405);
nor U7327 (N_7327,N_336,N_2738);
nor U7328 (N_7328,N_1965,N_4652);
and U7329 (N_7329,N_929,N_1735);
nor U7330 (N_7330,N_2604,N_2042);
and U7331 (N_7331,N_2418,N_2236);
nand U7332 (N_7332,N_3555,N_960);
and U7333 (N_7333,N_3958,N_1196);
nand U7334 (N_7334,N_3132,N_2178);
or U7335 (N_7335,N_3251,N_1598);
or U7336 (N_7336,N_100,N_4946);
and U7337 (N_7337,N_3400,N_1321);
nor U7338 (N_7338,N_604,N_1113);
or U7339 (N_7339,N_4042,N_2318);
nor U7340 (N_7340,N_2224,N_4974);
nor U7341 (N_7341,N_1627,N_2922);
and U7342 (N_7342,N_4516,N_4881);
xnor U7343 (N_7343,N_2322,N_2950);
and U7344 (N_7344,N_2021,N_2578);
and U7345 (N_7345,N_3700,N_1429);
nor U7346 (N_7346,N_1445,N_3669);
nor U7347 (N_7347,N_2062,N_4459);
and U7348 (N_7348,N_1836,N_2358);
nor U7349 (N_7349,N_1279,N_2400);
or U7350 (N_7350,N_1214,N_4765);
nor U7351 (N_7351,N_3150,N_4181);
nor U7352 (N_7352,N_2027,N_3895);
nor U7353 (N_7353,N_535,N_4529);
or U7354 (N_7354,N_1274,N_1042);
and U7355 (N_7355,N_1652,N_2263);
or U7356 (N_7356,N_3657,N_3823);
and U7357 (N_7357,N_2283,N_344);
xor U7358 (N_7358,N_4169,N_4546);
nor U7359 (N_7359,N_3345,N_3550);
or U7360 (N_7360,N_3692,N_1168);
or U7361 (N_7361,N_3023,N_2850);
nand U7362 (N_7362,N_4910,N_4844);
and U7363 (N_7363,N_4204,N_3104);
and U7364 (N_7364,N_4961,N_1413);
or U7365 (N_7365,N_4184,N_4000);
nand U7366 (N_7366,N_3661,N_2468);
or U7367 (N_7367,N_892,N_1660);
nor U7368 (N_7368,N_4825,N_614);
and U7369 (N_7369,N_4508,N_2994);
or U7370 (N_7370,N_4030,N_1872);
nor U7371 (N_7371,N_2713,N_43);
nor U7372 (N_7372,N_559,N_1655);
and U7373 (N_7373,N_3018,N_3438);
or U7374 (N_7374,N_1193,N_4133);
nand U7375 (N_7375,N_3549,N_4677);
nor U7376 (N_7376,N_85,N_220);
nor U7377 (N_7377,N_403,N_2487);
nor U7378 (N_7378,N_515,N_500);
and U7379 (N_7379,N_2831,N_2596);
or U7380 (N_7380,N_4374,N_2275);
and U7381 (N_7381,N_3441,N_4793);
nor U7382 (N_7382,N_825,N_1326);
nor U7383 (N_7383,N_3837,N_4471);
nand U7384 (N_7384,N_3389,N_4391);
nand U7385 (N_7385,N_4308,N_2347);
nand U7386 (N_7386,N_1610,N_3817);
or U7387 (N_7387,N_2548,N_2987);
nand U7388 (N_7388,N_3038,N_263);
nand U7389 (N_7389,N_4764,N_2742);
nor U7390 (N_7390,N_983,N_317);
nor U7391 (N_7391,N_19,N_597);
or U7392 (N_7392,N_4599,N_1696);
nand U7393 (N_7393,N_1863,N_1495);
nand U7394 (N_7394,N_415,N_4302);
and U7395 (N_7395,N_173,N_3589);
nor U7396 (N_7396,N_1968,N_3066);
xnor U7397 (N_7397,N_3886,N_2028);
nor U7398 (N_7398,N_2904,N_1244);
nor U7399 (N_7399,N_818,N_1809);
or U7400 (N_7400,N_213,N_2721);
or U7401 (N_7401,N_850,N_324);
or U7402 (N_7402,N_2856,N_347);
and U7403 (N_7403,N_2131,N_3458);
and U7404 (N_7404,N_2241,N_2070);
and U7405 (N_7405,N_1028,N_4732);
or U7406 (N_7406,N_4559,N_365);
or U7407 (N_7407,N_2536,N_885);
or U7408 (N_7408,N_463,N_4909);
nor U7409 (N_7409,N_2148,N_3281);
or U7410 (N_7410,N_1174,N_987);
or U7411 (N_7411,N_3321,N_1330);
nor U7412 (N_7412,N_1312,N_2329);
or U7413 (N_7413,N_2576,N_2492);
xnor U7414 (N_7414,N_4768,N_2919);
and U7415 (N_7415,N_1088,N_2396);
nor U7416 (N_7416,N_1381,N_866);
nor U7417 (N_7417,N_4317,N_1047);
nand U7418 (N_7418,N_964,N_272);
and U7419 (N_7419,N_2176,N_4596);
or U7420 (N_7420,N_3523,N_3876);
and U7421 (N_7421,N_1764,N_439);
or U7422 (N_7422,N_1455,N_2119);
nand U7423 (N_7423,N_4917,N_296);
and U7424 (N_7424,N_2571,N_1571);
and U7425 (N_7425,N_1883,N_1504);
nor U7426 (N_7426,N_1925,N_3436);
and U7427 (N_7427,N_1394,N_1830);
nor U7428 (N_7428,N_4653,N_3225);
nor U7429 (N_7429,N_1687,N_550);
nand U7430 (N_7430,N_4645,N_290);
or U7431 (N_7431,N_4776,N_493);
nand U7432 (N_7432,N_98,N_942);
nand U7433 (N_7433,N_1600,N_2012);
or U7434 (N_7434,N_4376,N_581);
nor U7435 (N_7435,N_3573,N_168);
or U7436 (N_7436,N_2833,N_119);
or U7437 (N_7437,N_4008,N_3416);
or U7438 (N_7438,N_3658,N_753);
nor U7439 (N_7439,N_2853,N_1834);
or U7440 (N_7440,N_2556,N_3185);
nand U7441 (N_7441,N_704,N_2733);
nor U7442 (N_7442,N_566,N_754);
nand U7443 (N_7443,N_4404,N_1524);
or U7444 (N_7444,N_2538,N_4955);
nand U7445 (N_7445,N_1395,N_1063);
and U7446 (N_7446,N_2917,N_2392);
and U7447 (N_7447,N_438,N_2597);
or U7448 (N_7448,N_3393,N_4059);
nor U7449 (N_7449,N_1669,N_3430);
nand U7450 (N_7450,N_1409,N_4699);
or U7451 (N_7451,N_490,N_1561);
nand U7452 (N_7452,N_14,N_3733);
nand U7453 (N_7453,N_2017,N_800);
nor U7454 (N_7454,N_1586,N_3945);
nor U7455 (N_7455,N_1224,N_3719);
or U7456 (N_7456,N_4387,N_2363);
and U7457 (N_7457,N_4134,N_3805);
nor U7458 (N_7458,N_4383,N_1712);
nor U7459 (N_7459,N_1991,N_245);
nand U7460 (N_7460,N_2929,N_3411);
and U7461 (N_7461,N_346,N_3897);
and U7462 (N_7462,N_545,N_427);
nand U7463 (N_7463,N_3966,N_3872);
or U7464 (N_7464,N_2677,N_1316);
nand U7465 (N_7465,N_3313,N_4327);
nand U7466 (N_7466,N_2584,N_4185);
xnor U7467 (N_7467,N_1072,N_1864);
nand U7468 (N_7468,N_2503,N_729);
nor U7469 (N_7469,N_2060,N_3955);
nor U7470 (N_7470,N_357,N_1629);
or U7471 (N_7471,N_3526,N_1039);
and U7472 (N_7472,N_660,N_4932);
xor U7473 (N_7473,N_2821,N_875);
and U7474 (N_7474,N_2949,N_4666);
or U7475 (N_7475,N_2583,N_3144);
nor U7476 (N_7476,N_1681,N_1468);
and U7477 (N_7477,N_1243,N_928);
nor U7478 (N_7478,N_2663,N_1297);
nand U7479 (N_7479,N_313,N_2581);
nand U7480 (N_7480,N_893,N_1542);
and U7481 (N_7481,N_156,N_4228);
nand U7482 (N_7482,N_2887,N_3894);
or U7483 (N_7483,N_3957,N_1210);
and U7484 (N_7484,N_2938,N_1080);
nand U7485 (N_7485,N_1275,N_1398);
and U7486 (N_7486,N_4742,N_3962);
nand U7487 (N_7487,N_2431,N_2520);
nand U7488 (N_7488,N_4523,N_2147);
nor U7489 (N_7489,N_4132,N_1844);
nand U7490 (N_7490,N_4155,N_1361);
nand U7491 (N_7491,N_1285,N_2560);
and U7492 (N_7492,N_2205,N_656);
and U7493 (N_7493,N_2647,N_802);
and U7494 (N_7494,N_3300,N_3642);
nor U7495 (N_7495,N_468,N_4116);
xnor U7496 (N_7496,N_1754,N_4898);
and U7497 (N_7497,N_751,N_242);
nor U7498 (N_7498,N_2509,N_537);
nor U7499 (N_7499,N_832,N_4090);
nor U7500 (N_7500,N_1692,N_2795);
and U7501 (N_7501,N_3474,N_2338);
nand U7502 (N_7502,N_2225,N_2355);
nand U7503 (N_7503,N_913,N_3294);
or U7504 (N_7504,N_2439,N_3273);
or U7505 (N_7505,N_4112,N_2675);
nor U7506 (N_7506,N_4883,N_1663);
and U7507 (N_7507,N_1519,N_409);
nor U7508 (N_7508,N_4792,N_3731);
nand U7509 (N_7509,N_2481,N_2729);
nor U7510 (N_7510,N_3860,N_3277);
and U7511 (N_7511,N_4441,N_1950);
and U7512 (N_7512,N_3808,N_1389);
and U7513 (N_7513,N_3627,N_3311);
nand U7514 (N_7514,N_4220,N_4321);
and U7515 (N_7515,N_3680,N_2270);
nand U7516 (N_7516,N_2425,N_1972);
or U7517 (N_7517,N_4366,N_3539);
and U7518 (N_7518,N_4683,N_1539);
nand U7519 (N_7519,N_4847,N_4884);
nor U7520 (N_7520,N_3570,N_1349);
and U7521 (N_7521,N_4093,N_3555);
nand U7522 (N_7522,N_3474,N_1078);
nand U7523 (N_7523,N_2371,N_2252);
nand U7524 (N_7524,N_996,N_4242);
or U7525 (N_7525,N_534,N_3251);
nor U7526 (N_7526,N_2430,N_4697);
or U7527 (N_7527,N_2043,N_883);
and U7528 (N_7528,N_4029,N_2885);
and U7529 (N_7529,N_1718,N_3261);
nor U7530 (N_7530,N_1698,N_217);
or U7531 (N_7531,N_1069,N_1206);
and U7532 (N_7532,N_1300,N_4550);
and U7533 (N_7533,N_2815,N_2626);
or U7534 (N_7534,N_3745,N_502);
nand U7535 (N_7535,N_581,N_3170);
xnor U7536 (N_7536,N_2417,N_1340);
or U7537 (N_7537,N_2947,N_2307);
nand U7538 (N_7538,N_4007,N_3600);
xnor U7539 (N_7539,N_3943,N_4004);
and U7540 (N_7540,N_1829,N_4301);
xnor U7541 (N_7541,N_959,N_2473);
nand U7542 (N_7542,N_3261,N_2686);
nor U7543 (N_7543,N_4614,N_413);
nor U7544 (N_7544,N_1058,N_1908);
and U7545 (N_7545,N_2828,N_4893);
or U7546 (N_7546,N_1932,N_566);
or U7547 (N_7547,N_2089,N_3755);
or U7548 (N_7548,N_104,N_2618);
or U7549 (N_7549,N_4412,N_3374);
or U7550 (N_7550,N_2400,N_701);
nand U7551 (N_7551,N_2468,N_3258);
and U7552 (N_7552,N_1650,N_1590);
and U7553 (N_7553,N_1266,N_1885);
and U7554 (N_7554,N_3631,N_3357);
nor U7555 (N_7555,N_1228,N_810);
or U7556 (N_7556,N_4270,N_3252);
or U7557 (N_7557,N_3323,N_4633);
nand U7558 (N_7558,N_1292,N_4425);
or U7559 (N_7559,N_1471,N_2355);
or U7560 (N_7560,N_2935,N_477);
and U7561 (N_7561,N_1695,N_1916);
nand U7562 (N_7562,N_4155,N_3326);
or U7563 (N_7563,N_3414,N_1596);
or U7564 (N_7564,N_127,N_3943);
and U7565 (N_7565,N_2471,N_4142);
nand U7566 (N_7566,N_2536,N_3837);
nand U7567 (N_7567,N_852,N_1232);
nand U7568 (N_7568,N_4022,N_1646);
and U7569 (N_7569,N_3367,N_4008);
and U7570 (N_7570,N_2099,N_4357);
nor U7571 (N_7571,N_3636,N_4810);
xnor U7572 (N_7572,N_64,N_3028);
nor U7573 (N_7573,N_741,N_1983);
nor U7574 (N_7574,N_3368,N_1787);
nand U7575 (N_7575,N_188,N_1184);
or U7576 (N_7576,N_4743,N_1736);
nand U7577 (N_7577,N_3053,N_933);
and U7578 (N_7578,N_80,N_4814);
or U7579 (N_7579,N_584,N_142);
or U7580 (N_7580,N_4111,N_4820);
and U7581 (N_7581,N_3749,N_151);
nand U7582 (N_7582,N_2161,N_4547);
xor U7583 (N_7583,N_1076,N_347);
and U7584 (N_7584,N_1005,N_3659);
nand U7585 (N_7585,N_1877,N_2186);
or U7586 (N_7586,N_4429,N_728);
nand U7587 (N_7587,N_308,N_1661);
nor U7588 (N_7588,N_4983,N_2962);
and U7589 (N_7589,N_2030,N_2630);
or U7590 (N_7590,N_193,N_3522);
and U7591 (N_7591,N_2538,N_3422);
or U7592 (N_7592,N_1817,N_2439);
and U7593 (N_7593,N_3721,N_238);
nand U7594 (N_7594,N_4972,N_3668);
and U7595 (N_7595,N_2013,N_4292);
nand U7596 (N_7596,N_3739,N_626);
nand U7597 (N_7597,N_2739,N_946);
nor U7598 (N_7598,N_1561,N_1052);
and U7599 (N_7599,N_1602,N_1511);
and U7600 (N_7600,N_3643,N_4607);
nand U7601 (N_7601,N_1823,N_4246);
and U7602 (N_7602,N_4215,N_1482);
nand U7603 (N_7603,N_4768,N_3727);
or U7604 (N_7604,N_3578,N_2361);
nand U7605 (N_7605,N_2682,N_2164);
nand U7606 (N_7606,N_1596,N_1831);
nand U7607 (N_7607,N_4179,N_4555);
nand U7608 (N_7608,N_4198,N_1093);
nor U7609 (N_7609,N_4167,N_2568);
or U7610 (N_7610,N_1173,N_3291);
nand U7611 (N_7611,N_725,N_3664);
nand U7612 (N_7612,N_2936,N_3706);
nand U7613 (N_7613,N_1080,N_1561);
and U7614 (N_7614,N_4636,N_519);
and U7615 (N_7615,N_4775,N_3621);
or U7616 (N_7616,N_1748,N_4075);
or U7617 (N_7617,N_4847,N_360);
nor U7618 (N_7618,N_2894,N_1857);
or U7619 (N_7619,N_3750,N_884);
nand U7620 (N_7620,N_4160,N_1577);
or U7621 (N_7621,N_311,N_3167);
or U7622 (N_7622,N_4499,N_518);
nor U7623 (N_7623,N_1764,N_342);
and U7624 (N_7624,N_696,N_2419);
nor U7625 (N_7625,N_4503,N_4672);
or U7626 (N_7626,N_4384,N_227);
nand U7627 (N_7627,N_3153,N_863);
nor U7628 (N_7628,N_3816,N_99);
and U7629 (N_7629,N_4445,N_4141);
or U7630 (N_7630,N_3443,N_3086);
nor U7631 (N_7631,N_1457,N_4601);
nand U7632 (N_7632,N_4983,N_3415);
nor U7633 (N_7633,N_1264,N_844);
nand U7634 (N_7634,N_3856,N_4161);
xor U7635 (N_7635,N_3657,N_1717);
xnor U7636 (N_7636,N_792,N_1259);
xor U7637 (N_7637,N_2740,N_1972);
xnor U7638 (N_7638,N_4861,N_2136);
nand U7639 (N_7639,N_3774,N_1540);
xor U7640 (N_7640,N_1425,N_328);
nand U7641 (N_7641,N_3244,N_810);
or U7642 (N_7642,N_2694,N_2984);
or U7643 (N_7643,N_3634,N_1537);
nor U7644 (N_7644,N_681,N_4708);
nor U7645 (N_7645,N_271,N_2514);
and U7646 (N_7646,N_4380,N_2981);
nand U7647 (N_7647,N_4374,N_350);
nand U7648 (N_7648,N_3364,N_4630);
and U7649 (N_7649,N_363,N_430);
or U7650 (N_7650,N_3185,N_4339);
nand U7651 (N_7651,N_1364,N_1959);
nor U7652 (N_7652,N_2473,N_3085);
nand U7653 (N_7653,N_2571,N_2051);
nand U7654 (N_7654,N_1056,N_2584);
nor U7655 (N_7655,N_205,N_662);
or U7656 (N_7656,N_1300,N_1574);
and U7657 (N_7657,N_1116,N_907);
nor U7658 (N_7658,N_3795,N_493);
nor U7659 (N_7659,N_2963,N_3642);
xor U7660 (N_7660,N_113,N_3691);
and U7661 (N_7661,N_1566,N_2942);
or U7662 (N_7662,N_3691,N_2922);
nand U7663 (N_7663,N_2071,N_2909);
or U7664 (N_7664,N_426,N_1776);
nor U7665 (N_7665,N_1741,N_2122);
nand U7666 (N_7666,N_3170,N_935);
or U7667 (N_7667,N_2299,N_22);
nand U7668 (N_7668,N_682,N_3026);
nor U7669 (N_7669,N_4974,N_4401);
and U7670 (N_7670,N_2504,N_1272);
or U7671 (N_7671,N_4658,N_193);
nor U7672 (N_7672,N_2132,N_3116);
or U7673 (N_7673,N_3416,N_3131);
nor U7674 (N_7674,N_2921,N_3701);
or U7675 (N_7675,N_2277,N_1850);
and U7676 (N_7676,N_2848,N_3274);
xnor U7677 (N_7677,N_1774,N_2708);
and U7678 (N_7678,N_3018,N_1668);
nor U7679 (N_7679,N_3572,N_4793);
nand U7680 (N_7680,N_4677,N_1443);
nor U7681 (N_7681,N_2067,N_1827);
nand U7682 (N_7682,N_20,N_4974);
nand U7683 (N_7683,N_959,N_1316);
and U7684 (N_7684,N_1683,N_4444);
nand U7685 (N_7685,N_1988,N_4802);
nand U7686 (N_7686,N_1576,N_2045);
or U7687 (N_7687,N_3007,N_4518);
and U7688 (N_7688,N_3393,N_3579);
and U7689 (N_7689,N_1114,N_945);
nand U7690 (N_7690,N_109,N_3112);
nor U7691 (N_7691,N_4319,N_735);
nor U7692 (N_7692,N_1607,N_3798);
nor U7693 (N_7693,N_4016,N_13);
nor U7694 (N_7694,N_4890,N_504);
nor U7695 (N_7695,N_2168,N_4666);
nand U7696 (N_7696,N_4203,N_203);
nor U7697 (N_7697,N_4497,N_958);
nor U7698 (N_7698,N_2763,N_2092);
nor U7699 (N_7699,N_4939,N_2008);
nor U7700 (N_7700,N_4361,N_4433);
nor U7701 (N_7701,N_4324,N_2218);
or U7702 (N_7702,N_3094,N_940);
nand U7703 (N_7703,N_1273,N_406);
nor U7704 (N_7704,N_788,N_4594);
or U7705 (N_7705,N_3385,N_4458);
xor U7706 (N_7706,N_2612,N_534);
nand U7707 (N_7707,N_2984,N_1970);
or U7708 (N_7708,N_2190,N_4158);
nor U7709 (N_7709,N_1803,N_2359);
nand U7710 (N_7710,N_66,N_3399);
nand U7711 (N_7711,N_4636,N_4538);
nand U7712 (N_7712,N_3319,N_2787);
nand U7713 (N_7713,N_3334,N_2053);
or U7714 (N_7714,N_423,N_4961);
and U7715 (N_7715,N_1692,N_4052);
nor U7716 (N_7716,N_4945,N_1674);
or U7717 (N_7717,N_4455,N_3922);
or U7718 (N_7718,N_2648,N_1234);
or U7719 (N_7719,N_1921,N_1290);
nor U7720 (N_7720,N_675,N_3526);
or U7721 (N_7721,N_884,N_4275);
nand U7722 (N_7722,N_272,N_653);
xor U7723 (N_7723,N_648,N_3252);
and U7724 (N_7724,N_1346,N_417);
or U7725 (N_7725,N_3325,N_991);
or U7726 (N_7726,N_1970,N_2030);
nand U7727 (N_7727,N_3211,N_3257);
and U7728 (N_7728,N_4636,N_1249);
nor U7729 (N_7729,N_2960,N_915);
nor U7730 (N_7730,N_3763,N_4529);
nor U7731 (N_7731,N_2620,N_1759);
xor U7732 (N_7732,N_2322,N_917);
nor U7733 (N_7733,N_4431,N_492);
nand U7734 (N_7734,N_4424,N_498);
nor U7735 (N_7735,N_447,N_2548);
nand U7736 (N_7736,N_3454,N_4614);
and U7737 (N_7737,N_2408,N_3568);
nand U7738 (N_7738,N_1576,N_3146);
or U7739 (N_7739,N_1703,N_4549);
nand U7740 (N_7740,N_4246,N_1983);
or U7741 (N_7741,N_2012,N_4855);
or U7742 (N_7742,N_3833,N_4969);
or U7743 (N_7743,N_3882,N_4376);
or U7744 (N_7744,N_344,N_2798);
and U7745 (N_7745,N_4687,N_3238);
nor U7746 (N_7746,N_1876,N_1766);
nand U7747 (N_7747,N_355,N_4473);
or U7748 (N_7748,N_1468,N_1884);
nor U7749 (N_7749,N_2939,N_3177);
or U7750 (N_7750,N_1974,N_1317);
or U7751 (N_7751,N_3752,N_1280);
nand U7752 (N_7752,N_4491,N_3562);
nand U7753 (N_7753,N_4425,N_2821);
nor U7754 (N_7754,N_3845,N_2825);
or U7755 (N_7755,N_3591,N_1425);
nor U7756 (N_7756,N_852,N_1788);
nor U7757 (N_7757,N_4677,N_447);
nor U7758 (N_7758,N_1525,N_2650);
and U7759 (N_7759,N_4232,N_3108);
nor U7760 (N_7760,N_3114,N_3786);
and U7761 (N_7761,N_1676,N_2241);
and U7762 (N_7762,N_3488,N_1146);
nor U7763 (N_7763,N_327,N_4907);
and U7764 (N_7764,N_494,N_3279);
or U7765 (N_7765,N_1821,N_3736);
nand U7766 (N_7766,N_231,N_2328);
or U7767 (N_7767,N_844,N_1677);
nand U7768 (N_7768,N_1811,N_2636);
nand U7769 (N_7769,N_1974,N_1405);
nand U7770 (N_7770,N_2099,N_4429);
nand U7771 (N_7771,N_701,N_1627);
or U7772 (N_7772,N_664,N_2136);
nor U7773 (N_7773,N_3666,N_1132);
nand U7774 (N_7774,N_1475,N_4630);
nand U7775 (N_7775,N_3882,N_3166);
or U7776 (N_7776,N_2808,N_32);
nor U7777 (N_7777,N_2131,N_3093);
and U7778 (N_7778,N_2423,N_1771);
and U7779 (N_7779,N_3861,N_3007);
and U7780 (N_7780,N_3954,N_3563);
nand U7781 (N_7781,N_2556,N_4124);
and U7782 (N_7782,N_1377,N_205);
nand U7783 (N_7783,N_3033,N_3616);
and U7784 (N_7784,N_1810,N_4692);
or U7785 (N_7785,N_2771,N_4503);
or U7786 (N_7786,N_2512,N_758);
nor U7787 (N_7787,N_1851,N_2075);
xor U7788 (N_7788,N_4291,N_4228);
or U7789 (N_7789,N_4923,N_4687);
or U7790 (N_7790,N_978,N_4788);
or U7791 (N_7791,N_1269,N_374);
and U7792 (N_7792,N_4269,N_4422);
nand U7793 (N_7793,N_3531,N_4436);
or U7794 (N_7794,N_3277,N_1022);
and U7795 (N_7795,N_2674,N_97);
nor U7796 (N_7796,N_2823,N_2412);
nor U7797 (N_7797,N_2075,N_4455);
nand U7798 (N_7798,N_25,N_1546);
nor U7799 (N_7799,N_2414,N_3757);
and U7800 (N_7800,N_2880,N_2750);
or U7801 (N_7801,N_903,N_1220);
nor U7802 (N_7802,N_3307,N_2996);
and U7803 (N_7803,N_4516,N_3410);
nor U7804 (N_7804,N_1660,N_2403);
or U7805 (N_7805,N_3953,N_790);
and U7806 (N_7806,N_1707,N_3466);
and U7807 (N_7807,N_3813,N_4099);
nor U7808 (N_7808,N_46,N_1083);
or U7809 (N_7809,N_2431,N_4395);
or U7810 (N_7810,N_3180,N_4333);
and U7811 (N_7811,N_2026,N_457);
nor U7812 (N_7812,N_3776,N_3698);
nor U7813 (N_7813,N_1653,N_2195);
xnor U7814 (N_7814,N_2335,N_4129);
nand U7815 (N_7815,N_4512,N_2154);
and U7816 (N_7816,N_4941,N_3586);
nand U7817 (N_7817,N_4087,N_1232);
and U7818 (N_7818,N_1546,N_4094);
and U7819 (N_7819,N_2696,N_4553);
nor U7820 (N_7820,N_4190,N_1832);
nor U7821 (N_7821,N_1547,N_632);
and U7822 (N_7822,N_3773,N_2343);
nor U7823 (N_7823,N_1772,N_1110);
nand U7824 (N_7824,N_3226,N_999);
nand U7825 (N_7825,N_1551,N_4825);
nor U7826 (N_7826,N_231,N_1243);
nand U7827 (N_7827,N_1712,N_3144);
nand U7828 (N_7828,N_4842,N_2522);
or U7829 (N_7829,N_3211,N_2750);
nand U7830 (N_7830,N_17,N_2692);
nand U7831 (N_7831,N_184,N_3564);
and U7832 (N_7832,N_1378,N_4648);
or U7833 (N_7833,N_1598,N_3055);
nand U7834 (N_7834,N_3182,N_3073);
nor U7835 (N_7835,N_2360,N_1058);
or U7836 (N_7836,N_1805,N_4590);
or U7837 (N_7837,N_4798,N_2696);
nor U7838 (N_7838,N_372,N_3116);
nand U7839 (N_7839,N_1721,N_1577);
nor U7840 (N_7840,N_4729,N_3976);
and U7841 (N_7841,N_1152,N_913);
and U7842 (N_7842,N_1040,N_3963);
or U7843 (N_7843,N_2030,N_1227);
and U7844 (N_7844,N_215,N_3434);
and U7845 (N_7845,N_408,N_3195);
or U7846 (N_7846,N_2414,N_1928);
xnor U7847 (N_7847,N_3955,N_2046);
nand U7848 (N_7848,N_4212,N_740);
nor U7849 (N_7849,N_989,N_4030);
or U7850 (N_7850,N_3505,N_413);
or U7851 (N_7851,N_4354,N_572);
nand U7852 (N_7852,N_1608,N_4969);
nand U7853 (N_7853,N_2311,N_1675);
nor U7854 (N_7854,N_1593,N_1235);
nand U7855 (N_7855,N_2845,N_4944);
nor U7856 (N_7856,N_4595,N_1408);
nor U7857 (N_7857,N_2256,N_1677);
nand U7858 (N_7858,N_2383,N_3798);
and U7859 (N_7859,N_1667,N_3023);
xnor U7860 (N_7860,N_4167,N_3436);
nand U7861 (N_7861,N_4852,N_441);
nand U7862 (N_7862,N_4648,N_3819);
and U7863 (N_7863,N_1364,N_1107);
or U7864 (N_7864,N_609,N_3376);
or U7865 (N_7865,N_2951,N_3819);
nor U7866 (N_7866,N_4359,N_4099);
and U7867 (N_7867,N_1417,N_2850);
or U7868 (N_7868,N_225,N_1012);
or U7869 (N_7869,N_896,N_4248);
nor U7870 (N_7870,N_3344,N_4726);
and U7871 (N_7871,N_1982,N_4223);
nand U7872 (N_7872,N_2653,N_3437);
or U7873 (N_7873,N_86,N_826);
and U7874 (N_7874,N_3788,N_4062);
nand U7875 (N_7875,N_1664,N_2072);
nand U7876 (N_7876,N_1556,N_3551);
and U7877 (N_7877,N_4010,N_2229);
nand U7878 (N_7878,N_1185,N_228);
and U7879 (N_7879,N_107,N_3138);
xnor U7880 (N_7880,N_2948,N_2838);
nor U7881 (N_7881,N_2634,N_3628);
or U7882 (N_7882,N_815,N_3279);
nand U7883 (N_7883,N_2273,N_332);
and U7884 (N_7884,N_1941,N_2354);
nor U7885 (N_7885,N_740,N_1211);
and U7886 (N_7886,N_1891,N_2145);
xnor U7887 (N_7887,N_4685,N_3814);
or U7888 (N_7888,N_583,N_3272);
nand U7889 (N_7889,N_3471,N_1710);
or U7890 (N_7890,N_4314,N_2948);
and U7891 (N_7891,N_2229,N_1593);
nand U7892 (N_7892,N_1797,N_2778);
and U7893 (N_7893,N_3495,N_1711);
nand U7894 (N_7894,N_2430,N_4183);
and U7895 (N_7895,N_2525,N_909);
nor U7896 (N_7896,N_1710,N_2159);
nor U7897 (N_7897,N_2827,N_3615);
or U7898 (N_7898,N_4571,N_4547);
or U7899 (N_7899,N_1094,N_650);
and U7900 (N_7900,N_4246,N_2887);
and U7901 (N_7901,N_4787,N_3083);
or U7902 (N_7902,N_4173,N_3368);
nand U7903 (N_7903,N_4444,N_2075);
nor U7904 (N_7904,N_4860,N_2419);
and U7905 (N_7905,N_194,N_2133);
nor U7906 (N_7906,N_973,N_4588);
and U7907 (N_7907,N_4112,N_1027);
nor U7908 (N_7908,N_2396,N_3876);
and U7909 (N_7909,N_3811,N_3590);
nand U7910 (N_7910,N_2370,N_806);
nor U7911 (N_7911,N_2316,N_2200);
nand U7912 (N_7912,N_971,N_1636);
or U7913 (N_7913,N_4169,N_4137);
and U7914 (N_7914,N_2837,N_1397);
nand U7915 (N_7915,N_2405,N_1086);
nor U7916 (N_7916,N_4094,N_514);
nand U7917 (N_7917,N_722,N_4562);
nor U7918 (N_7918,N_35,N_293);
nor U7919 (N_7919,N_560,N_4831);
and U7920 (N_7920,N_2786,N_4553);
nand U7921 (N_7921,N_4101,N_4450);
or U7922 (N_7922,N_1362,N_984);
nor U7923 (N_7923,N_860,N_2538);
nand U7924 (N_7924,N_3185,N_3108);
xor U7925 (N_7925,N_4660,N_4177);
nand U7926 (N_7926,N_3317,N_4538);
nor U7927 (N_7927,N_1974,N_4415);
or U7928 (N_7928,N_64,N_631);
or U7929 (N_7929,N_4808,N_1506);
nor U7930 (N_7930,N_1288,N_2888);
nand U7931 (N_7931,N_3536,N_2960);
nor U7932 (N_7932,N_1390,N_1621);
and U7933 (N_7933,N_3324,N_2924);
nand U7934 (N_7934,N_1187,N_4312);
nand U7935 (N_7935,N_1458,N_4664);
nand U7936 (N_7936,N_3831,N_2407);
or U7937 (N_7937,N_2533,N_17);
or U7938 (N_7938,N_3003,N_1547);
and U7939 (N_7939,N_1516,N_2726);
nor U7940 (N_7940,N_4793,N_4163);
and U7941 (N_7941,N_18,N_1061);
and U7942 (N_7942,N_3550,N_1816);
and U7943 (N_7943,N_154,N_1312);
xor U7944 (N_7944,N_1375,N_4710);
nor U7945 (N_7945,N_1034,N_436);
nor U7946 (N_7946,N_3661,N_639);
or U7947 (N_7947,N_2721,N_2042);
or U7948 (N_7948,N_4835,N_3976);
or U7949 (N_7949,N_2132,N_735);
and U7950 (N_7950,N_1709,N_1612);
and U7951 (N_7951,N_3216,N_4063);
or U7952 (N_7952,N_4449,N_342);
and U7953 (N_7953,N_651,N_2929);
or U7954 (N_7954,N_2406,N_4194);
nor U7955 (N_7955,N_811,N_3957);
or U7956 (N_7956,N_1736,N_4381);
nand U7957 (N_7957,N_1847,N_4013);
and U7958 (N_7958,N_1551,N_4982);
nor U7959 (N_7959,N_787,N_2151);
nor U7960 (N_7960,N_4019,N_3919);
nand U7961 (N_7961,N_4186,N_1716);
and U7962 (N_7962,N_3398,N_1284);
nor U7963 (N_7963,N_2568,N_1297);
or U7964 (N_7964,N_3637,N_2774);
xnor U7965 (N_7965,N_1767,N_280);
nor U7966 (N_7966,N_2777,N_4931);
nor U7967 (N_7967,N_251,N_2900);
or U7968 (N_7968,N_1226,N_1261);
nand U7969 (N_7969,N_3693,N_40);
and U7970 (N_7970,N_1963,N_4910);
and U7971 (N_7971,N_567,N_3507);
nor U7972 (N_7972,N_105,N_4746);
or U7973 (N_7973,N_1283,N_1508);
or U7974 (N_7974,N_4840,N_456);
xor U7975 (N_7975,N_1655,N_4168);
nand U7976 (N_7976,N_3708,N_367);
nor U7977 (N_7977,N_3685,N_473);
and U7978 (N_7978,N_3113,N_246);
or U7979 (N_7979,N_1237,N_1247);
nor U7980 (N_7980,N_989,N_1797);
nand U7981 (N_7981,N_1857,N_3704);
and U7982 (N_7982,N_1622,N_2699);
nand U7983 (N_7983,N_3870,N_1557);
and U7984 (N_7984,N_3115,N_3169);
nand U7985 (N_7985,N_14,N_3728);
and U7986 (N_7986,N_3197,N_4634);
or U7987 (N_7987,N_3504,N_3032);
nand U7988 (N_7988,N_2715,N_4771);
and U7989 (N_7989,N_1947,N_4397);
nand U7990 (N_7990,N_4683,N_35);
nor U7991 (N_7991,N_1135,N_4353);
xor U7992 (N_7992,N_2773,N_1859);
and U7993 (N_7993,N_1352,N_1676);
or U7994 (N_7994,N_1507,N_3110);
or U7995 (N_7995,N_2351,N_728);
xor U7996 (N_7996,N_2860,N_3034);
nor U7997 (N_7997,N_1332,N_1614);
or U7998 (N_7998,N_3874,N_3051);
or U7999 (N_7999,N_3535,N_1169);
nand U8000 (N_8000,N_2703,N_3172);
nand U8001 (N_8001,N_3320,N_878);
and U8002 (N_8002,N_3437,N_4801);
and U8003 (N_8003,N_113,N_4715);
xor U8004 (N_8004,N_689,N_4126);
nor U8005 (N_8005,N_1101,N_1973);
and U8006 (N_8006,N_3693,N_1610);
nor U8007 (N_8007,N_39,N_1597);
nor U8008 (N_8008,N_270,N_1775);
nor U8009 (N_8009,N_2298,N_3892);
or U8010 (N_8010,N_2027,N_95);
and U8011 (N_8011,N_3941,N_4843);
nand U8012 (N_8012,N_882,N_2444);
or U8013 (N_8013,N_3806,N_2129);
nand U8014 (N_8014,N_64,N_3675);
nor U8015 (N_8015,N_4451,N_2579);
and U8016 (N_8016,N_2221,N_1936);
or U8017 (N_8017,N_4392,N_1291);
and U8018 (N_8018,N_2219,N_1500);
or U8019 (N_8019,N_1079,N_2128);
xor U8020 (N_8020,N_3660,N_2105);
or U8021 (N_8021,N_1151,N_278);
xor U8022 (N_8022,N_2125,N_2170);
and U8023 (N_8023,N_3403,N_617);
nand U8024 (N_8024,N_264,N_1449);
nor U8025 (N_8025,N_2840,N_291);
nand U8026 (N_8026,N_1974,N_283);
nor U8027 (N_8027,N_147,N_23);
nand U8028 (N_8028,N_1210,N_3695);
xor U8029 (N_8029,N_3881,N_3609);
nor U8030 (N_8030,N_2264,N_2610);
or U8031 (N_8031,N_3298,N_1094);
nand U8032 (N_8032,N_700,N_4669);
and U8033 (N_8033,N_3983,N_4860);
nor U8034 (N_8034,N_898,N_2870);
nand U8035 (N_8035,N_4063,N_3717);
and U8036 (N_8036,N_2672,N_3478);
and U8037 (N_8037,N_449,N_1424);
nand U8038 (N_8038,N_4428,N_2744);
nand U8039 (N_8039,N_89,N_4947);
nand U8040 (N_8040,N_1889,N_1359);
and U8041 (N_8041,N_2505,N_3324);
nand U8042 (N_8042,N_3835,N_4600);
nor U8043 (N_8043,N_1104,N_1859);
nand U8044 (N_8044,N_913,N_3225);
nor U8045 (N_8045,N_3425,N_4204);
nor U8046 (N_8046,N_4819,N_2697);
nor U8047 (N_8047,N_3982,N_2780);
nand U8048 (N_8048,N_1095,N_4767);
nor U8049 (N_8049,N_2882,N_422);
nor U8050 (N_8050,N_2043,N_4224);
and U8051 (N_8051,N_4843,N_77);
and U8052 (N_8052,N_2943,N_54);
nand U8053 (N_8053,N_3197,N_941);
and U8054 (N_8054,N_1215,N_1705);
or U8055 (N_8055,N_228,N_834);
and U8056 (N_8056,N_138,N_3393);
or U8057 (N_8057,N_2234,N_1687);
or U8058 (N_8058,N_3068,N_920);
nand U8059 (N_8059,N_3356,N_330);
and U8060 (N_8060,N_2198,N_4443);
nor U8061 (N_8061,N_4789,N_414);
or U8062 (N_8062,N_3230,N_1320);
nand U8063 (N_8063,N_4441,N_1536);
and U8064 (N_8064,N_3114,N_2520);
nand U8065 (N_8065,N_2662,N_2704);
or U8066 (N_8066,N_1369,N_4577);
nand U8067 (N_8067,N_3021,N_4767);
or U8068 (N_8068,N_3319,N_2028);
nand U8069 (N_8069,N_2260,N_1450);
or U8070 (N_8070,N_2294,N_4039);
and U8071 (N_8071,N_2954,N_2265);
or U8072 (N_8072,N_4822,N_4200);
and U8073 (N_8073,N_2956,N_4434);
nor U8074 (N_8074,N_4616,N_2173);
and U8075 (N_8075,N_4954,N_3649);
and U8076 (N_8076,N_229,N_1857);
nand U8077 (N_8077,N_4007,N_555);
or U8078 (N_8078,N_3734,N_1226);
nand U8079 (N_8079,N_3853,N_4596);
nor U8080 (N_8080,N_4019,N_4897);
nor U8081 (N_8081,N_746,N_3087);
xnor U8082 (N_8082,N_987,N_3699);
and U8083 (N_8083,N_1617,N_2806);
nor U8084 (N_8084,N_954,N_4070);
and U8085 (N_8085,N_1490,N_4357);
nor U8086 (N_8086,N_4520,N_4127);
nor U8087 (N_8087,N_4048,N_3422);
and U8088 (N_8088,N_1474,N_354);
xor U8089 (N_8089,N_657,N_4379);
nor U8090 (N_8090,N_2276,N_4080);
nor U8091 (N_8091,N_2273,N_3367);
nand U8092 (N_8092,N_1262,N_2789);
and U8093 (N_8093,N_4291,N_1744);
and U8094 (N_8094,N_574,N_3404);
nor U8095 (N_8095,N_3775,N_3251);
or U8096 (N_8096,N_4396,N_2715);
nand U8097 (N_8097,N_194,N_3425);
nand U8098 (N_8098,N_2845,N_3061);
nand U8099 (N_8099,N_4679,N_1472);
xor U8100 (N_8100,N_426,N_4720);
or U8101 (N_8101,N_1267,N_297);
and U8102 (N_8102,N_219,N_911);
and U8103 (N_8103,N_1451,N_1359);
or U8104 (N_8104,N_819,N_3687);
or U8105 (N_8105,N_4754,N_1364);
nand U8106 (N_8106,N_4018,N_2207);
nand U8107 (N_8107,N_1647,N_1674);
and U8108 (N_8108,N_2612,N_3470);
nor U8109 (N_8109,N_943,N_698);
nand U8110 (N_8110,N_3785,N_1849);
or U8111 (N_8111,N_1333,N_3174);
and U8112 (N_8112,N_914,N_850);
or U8113 (N_8113,N_3195,N_3550);
nand U8114 (N_8114,N_1506,N_2651);
and U8115 (N_8115,N_4946,N_1973);
and U8116 (N_8116,N_3947,N_2133);
or U8117 (N_8117,N_4020,N_1019);
nor U8118 (N_8118,N_1881,N_3369);
nor U8119 (N_8119,N_4608,N_2634);
nand U8120 (N_8120,N_1182,N_305);
and U8121 (N_8121,N_153,N_3340);
or U8122 (N_8122,N_3918,N_709);
nor U8123 (N_8123,N_4374,N_2);
nand U8124 (N_8124,N_2743,N_2579);
and U8125 (N_8125,N_3811,N_2986);
nor U8126 (N_8126,N_1494,N_1167);
nand U8127 (N_8127,N_1107,N_2814);
and U8128 (N_8128,N_1520,N_296);
nor U8129 (N_8129,N_625,N_4518);
nand U8130 (N_8130,N_1231,N_1483);
and U8131 (N_8131,N_3927,N_509);
nor U8132 (N_8132,N_1301,N_2266);
nand U8133 (N_8133,N_166,N_2848);
and U8134 (N_8134,N_3451,N_2426);
or U8135 (N_8135,N_1245,N_4706);
and U8136 (N_8136,N_2544,N_2957);
or U8137 (N_8137,N_337,N_2798);
nor U8138 (N_8138,N_1832,N_4211);
and U8139 (N_8139,N_4945,N_1153);
nand U8140 (N_8140,N_2289,N_1972);
nand U8141 (N_8141,N_2031,N_3532);
nor U8142 (N_8142,N_3424,N_1414);
or U8143 (N_8143,N_4900,N_4607);
or U8144 (N_8144,N_68,N_204);
nand U8145 (N_8145,N_2511,N_1628);
and U8146 (N_8146,N_1882,N_3074);
or U8147 (N_8147,N_3992,N_1522);
and U8148 (N_8148,N_3440,N_2454);
nor U8149 (N_8149,N_197,N_1301);
nor U8150 (N_8150,N_4265,N_391);
and U8151 (N_8151,N_1454,N_3859);
or U8152 (N_8152,N_2063,N_1040);
nand U8153 (N_8153,N_3613,N_227);
nand U8154 (N_8154,N_721,N_4678);
or U8155 (N_8155,N_3671,N_4507);
or U8156 (N_8156,N_932,N_1467);
or U8157 (N_8157,N_1271,N_807);
nand U8158 (N_8158,N_2850,N_2468);
nand U8159 (N_8159,N_2100,N_4027);
nand U8160 (N_8160,N_4444,N_3012);
or U8161 (N_8161,N_599,N_646);
or U8162 (N_8162,N_4309,N_3783);
nor U8163 (N_8163,N_2745,N_1580);
nand U8164 (N_8164,N_1885,N_4374);
nand U8165 (N_8165,N_2674,N_87);
nor U8166 (N_8166,N_634,N_2542);
or U8167 (N_8167,N_1134,N_3662);
and U8168 (N_8168,N_4062,N_433);
and U8169 (N_8169,N_1143,N_2381);
and U8170 (N_8170,N_124,N_614);
or U8171 (N_8171,N_3312,N_2873);
and U8172 (N_8172,N_669,N_4677);
nand U8173 (N_8173,N_4584,N_4160);
nor U8174 (N_8174,N_2677,N_947);
nand U8175 (N_8175,N_415,N_1387);
nand U8176 (N_8176,N_612,N_3297);
or U8177 (N_8177,N_389,N_4899);
nand U8178 (N_8178,N_819,N_1739);
or U8179 (N_8179,N_2375,N_1232);
or U8180 (N_8180,N_365,N_4326);
or U8181 (N_8181,N_4903,N_1974);
nand U8182 (N_8182,N_3047,N_1273);
and U8183 (N_8183,N_1409,N_2599);
nand U8184 (N_8184,N_3654,N_7);
nor U8185 (N_8185,N_3578,N_41);
xor U8186 (N_8186,N_641,N_2347);
and U8187 (N_8187,N_2985,N_2428);
and U8188 (N_8188,N_2116,N_4278);
or U8189 (N_8189,N_4554,N_3385);
nand U8190 (N_8190,N_4657,N_2495);
and U8191 (N_8191,N_4410,N_4773);
nor U8192 (N_8192,N_1190,N_3491);
and U8193 (N_8193,N_3648,N_4994);
and U8194 (N_8194,N_2761,N_1727);
nand U8195 (N_8195,N_3029,N_1482);
or U8196 (N_8196,N_539,N_1117);
nor U8197 (N_8197,N_1095,N_1277);
or U8198 (N_8198,N_549,N_295);
or U8199 (N_8199,N_856,N_438);
nor U8200 (N_8200,N_1800,N_4400);
nand U8201 (N_8201,N_4374,N_926);
and U8202 (N_8202,N_2184,N_481);
or U8203 (N_8203,N_4503,N_1979);
and U8204 (N_8204,N_3292,N_4680);
and U8205 (N_8205,N_4420,N_4073);
nor U8206 (N_8206,N_3894,N_3012);
nor U8207 (N_8207,N_775,N_4334);
xnor U8208 (N_8208,N_1828,N_3055);
and U8209 (N_8209,N_1162,N_1294);
or U8210 (N_8210,N_216,N_2606);
and U8211 (N_8211,N_3852,N_3627);
nor U8212 (N_8212,N_1347,N_3362);
xor U8213 (N_8213,N_1724,N_2909);
and U8214 (N_8214,N_3336,N_4506);
nand U8215 (N_8215,N_770,N_196);
or U8216 (N_8216,N_3580,N_1810);
nand U8217 (N_8217,N_1418,N_2870);
nand U8218 (N_8218,N_4934,N_3266);
or U8219 (N_8219,N_848,N_2508);
nand U8220 (N_8220,N_492,N_2664);
nor U8221 (N_8221,N_237,N_738);
or U8222 (N_8222,N_842,N_2333);
nor U8223 (N_8223,N_2901,N_3300);
nand U8224 (N_8224,N_2297,N_170);
nand U8225 (N_8225,N_2689,N_2790);
or U8226 (N_8226,N_4971,N_761);
nand U8227 (N_8227,N_506,N_3784);
nor U8228 (N_8228,N_721,N_1466);
nand U8229 (N_8229,N_1717,N_273);
nor U8230 (N_8230,N_4786,N_2416);
nor U8231 (N_8231,N_2964,N_2626);
or U8232 (N_8232,N_3596,N_548);
nand U8233 (N_8233,N_1543,N_1507);
or U8234 (N_8234,N_4882,N_3285);
nor U8235 (N_8235,N_1913,N_2955);
nand U8236 (N_8236,N_1758,N_3742);
nand U8237 (N_8237,N_3581,N_1921);
nor U8238 (N_8238,N_1641,N_1918);
and U8239 (N_8239,N_2489,N_3779);
and U8240 (N_8240,N_1186,N_1461);
and U8241 (N_8241,N_494,N_52);
or U8242 (N_8242,N_2155,N_3453);
nor U8243 (N_8243,N_336,N_1384);
nor U8244 (N_8244,N_2729,N_1826);
nor U8245 (N_8245,N_1321,N_4388);
or U8246 (N_8246,N_1573,N_2203);
and U8247 (N_8247,N_3572,N_822);
nand U8248 (N_8248,N_3798,N_2846);
nor U8249 (N_8249,N_2790,N_4512);
or U8250 (N_8250,N_3549,N_4212);
and U8251 (N_8251,N_1101,N_2952);
nand U8252 (N_8252,N_2034,N_1562);
or U8253 (N_8253,N_2437,N_3420);
and U8254 (N_8254,N_572,N_2153);
or U8255 (N_8255,N_577,N_760);
nand U8256 (N_8256,N_2331,N_3438);
and U8257 (N_8257,N_2083,N_4874);
or U8258 (N_8258,N_89,N_1649);
nor U8259 (N_8259,N_4005,N_3311);
or U8260 (N_8260,N_4351,N_1936);
and U8261 (N_8261,N_1298,N_44);
nand U8262 (N_8262,N_1883,N_3357);
nand U8263 (N_8263,N_1542,N_1169);
or U8264 (N_8264,N_1311,N_2722);
and U8265 (N_8265,N_1581,N_624);
nand U8266 (N_8266,N_2522,N_3615);
and U8267 (N_8267,N_4859,N_3215);
nand U8268 (N_8268,N_2937,N_867);
nor U8269 (N_8269,N_2096,N_167);
and U8270 (N_8270,N_2921,N_2200);
nor U8271 (N_8271,N_1753,N_2147);
nand U8272 (N_8272,N_1996,N_3796);
nor U8273 (N_8273,N_1808,N_4744);
or U8274 (N_8274,N_3720,N_115);
or U8275 (N_8275,N_1393,N_124);
nor U8276 (N_8276,N_2124,N_4724);
and U8277 (N_8277,N_4099,N_4952);
nand U8278 (N_8278,N_3449,N_1957);
or U8279 (N_8279,N_286,N_4933);
nand U8280 (N_8280,N_3172,N_2098);
or U8281 (N_8281,N_1145,N_4493);
nor U8282 (N_8282,N_3817,N_4926);
nand U8283 (N_8283,N_1487,N_2262);
nand U8284 (N_8284,N_341,N_1914);
nand U8285 (N_8285,N_958,N_1915);
nand U8286 (N_8286,N_1278,N_3741);
and U8287 (N_8287,N_432,N_4838);
nand U8288 (N_8288,N_702,N_992);
and U8289 (N_8289,N_1849,N_4988);
nor U8290 (N_8290,N_292,N_1944);
nor U8291 (N_8291,N_3441,N_599);
nand U8292 (N_8292,N_3497,N_2353);
nand U8293 (N_8293,N_2175,N_4811);
or U8294 (N_8294,N_925,N_1056);
nor U8295 (N_8295,N_3490,N_2041);
nand U8296 (N_8296,N_2698,N_3781);
and U8297 (N_8297,N_4817,N_2367);
nand U8298 (N_8298,N_953,N_4506);
or U8299 (N_8299,N_4741,N_4580);
and U8300 (N_8300,N_3421,N_2002);
nand U8301 (N_8301,N_168,N_336);
nand U8302 (N_8302,N_3689,N_1859);
or U8303 (N_8303,N_1990,N_4465);
or U8304 (N_8304,N_2436,N_3308);
nor U8305 (N_8305,N_1451,N_3781);
nor U8306 (N_8306,N_381,N_730);
nor U8307 (N_8307,N_1140,N_1930);
nand U8308 (N_8308,N_2096,N_1304);
nand U8309 (N_8309,N_4900,N_3991);
and U8310 (N_8310,N_1202,N_518);
or U8311 (N_8311,N_1507,N_3900);
nand U8312 (N_8312,N_1434,N_3539);
or U8313 (N_8313,N_4094,N_786);
nand U8314 (N_8314,N_4460,N_3540);
nand U8315 (N_8315,N_87,N_4740);
nor U8316 (N_8316,N_1669,N_2084);
nor U8317 (N_8317,N_4190,N_4807);
nand U8318 (N_8318,N_3084,N_2281);
nor U8319 (N_8319,N_1552,N_2554);
or U8320 (N_8320,N_2573,N_2625);
or U8321 (N_8321,N_4735,N_3232);
or U8322 (N_8322,N_2856,N_727);
and U8323 (N_8323,N_3615,N_1955);
and U8324 (N_8324,N_2630,N_4192);
nand U8325 (N_8325,N_676,N_1409);
nor U8326 (N_8326,N_1413,N_4835);
or U8327 (N_8327,N_241,N_4318);
nor U8328 (N_8328,N_597,N_1565);
and U8329 (N_8329,N_2063,N_94);
and U8330 (N_8330,N_3346,N_4302);
nand U8331 (N_8331,N_4499,N_4618);
nor U8332 (N_8332,N_700,N_2648);
nand U8333 (N_8333,N_982,N_1901);
and U8334 (N_8334,N_726,N_605);
nor U8335 (N_8335,N_3963,N_4476);
nor U8336 (N_8336,N_3458,N_3201);
nor U8337 (N_8337,N_4667,N_1412);
nand U8338 (N_8338,N_1980,N_4928);
nand U8339 (N_8339,N_1614,N_4247);
nor U8340 (N_8340,N_222,N_281);
or U8341 (N_8341,N_4511,N_2405);
nand U8342 (N_8342,N_4940,N_1321);
nand U8343 (N_8343,N_4411,N_114);
or U8344 (N_8344,N_2314,N_981);
and U8345 (N_8345,N_504,N_3391);
nand U8346 (N_8346,N_1826,N_3933);
or U8347 (N_8347,N_534,N_4264);
nand U8348 (N_8348,N_2557,N_4546);
nor U8349 (N_8349,N_910,N_2942);
and U8350 (N_8350,N_2506,N_2837);
and U8351 (N_8351,N_90,N_4338);
nor U8352 (N_8352,N_2786,N_233);
nand U8353 (N_8353,N_1929,N_1007);
and U8354 (N_8354,N_1040,N_2524);
nand U8355 (N_8355,N_2910,N_1745);
nand U8356 (N_8356,N_1835,N_2634);
or U8357 (N_8357,N_3717,N_2671);
nand U8358 (N_8358,N_4917,N_2636);
and U8359 (N_8359,N_933,N_799);
nand U8360 (N_8360,N_640,N_4458);
and U8361 (N_8361,N_778,N_2817);
and U8362 (N_8362,N_1436,N_1265);
or U8363 (N_8363,N_2059,N_562);
and U8364 (N_8364,N_2665,N_4899);
nor U8365 (N_8365,N_4498,N_2532);
or U8366 (N_8366,N_2119,N_3084);
nand U8367 (N_8367,N_2296,N_1457);
or U8368 (N_8368,N_4800,N_295);
nor U8369 (N_8369,N_2324,N_1515);
or U8370 (N_8370,N_4307,N_822);
xnor U8371 (N_8371,N_2588,N_3737);
nor U8372 (N_8372,N_4020,N_3444);
nor U8373 (N_8373,N_2183,N_2982);
or U8374 (N_8374,N_110,N_1060);
or U8375 (N_8375,N_4111,N_67);
or U8376 (N_8376,N_2690,N_2106);
nor U8377 (N_8377,N_797,N_4213);
or U8378 (N_8378,N_1452,N_167);
or U8379 (N_8379,N_2780,N_4871);
nand U8380 (N_8380,N_2804,N_3152);
nand U8381 (N_8381,N_2979,N_251);
or U8382 (N_8382,N_2929,N_3935);
or U8383 (N_8383,N_1264,N_4229);
nand U8384 (N_8384,N_4107,N_3294);
and U8385 (N_8385,N_3632,N_1493);
xnor U8386 (N_8386,N_276,N_2572);
or U8387 (N_8387,N_168,N_2755);
nor U8388 (N_8388,N_4380,N_4030);
or U8389 (N_8389,N_2823,N_3077);
or U8390 (N_8390,N_766,N_4165);
nor U8391 (N_8391,N_2463,N_4404);
nor U8392 (N_8392,N_3870,N_1270);
or U8393 (N_8393,N_4684,N_3993);
or U8394 (N_8394,N_2407,N_3460);
or U8395 (N_8395,N_230,N_677);
or U8396 (N_8396,N_1636,N_335);
and U8397 (N_8397,N_2178,N_411);
and U8398 (N_8398,N_255,N_1900);
or U8399 (N_8399,N_2242,N_4979);
nand U8400 (N_8400,N_213,N_727);
or U8401 (N_8401,N_2200,N_2905);
nor U8402 (N_8402,N_2493,N_1746);
nand U8403 (N_8403,N_1296,N_230);
and U8404 (N_8404,N_398,N_479);
or U8405 (N_8405,N_826,N_1823);
nand U8406 (N_8406,N_1416,N_3554);
nand U8407 (N_8407,N_1754,N_267);
nand U8408 (N_8408,N_176,N_94);
or U8409 (N_8409,N_2350,N_4006);
and U8410 (N_8410,N_3922,N_4007);
or U8411 (N_8411,N_2452,N_4050);
nor U8412 (N_8412,N_3792,N_1907);
and U8413 (N_8413,N_43,N_4011);
or U8414 (N_8414,N_714,N_688);
xnor U8415 (N_8415,N_3463,N_4954);
nand U8416 (N_8416,N_2838,N_2071);
xnor U8417 (N_8417,N_3429,N_4142);
and U8418 (N_8418,N_2777,N_3235);
nor U8419 (N_8419,N_993,N_2104);
nand U8420 (N_8420,N_3861,N_34);
and U8421 (N_8421,N_2029,N_4325);
or U8422 (N_8422,N_4342,N_4219);
or U8423 (N_8423,N_4113,N_1649);
nor U8424 (N_8424,N_3463,N_1437);
nand U8425 (N_8425,N_1614,N_2966);
and U8426 (N_8426,N_4646,N_1794);
nand U8427 (N_8427,N_2682,N_1642);
nand U8428 (N_8428,N_2516,N_3158);
nand U8429 (N_8429,N_4948,N_3292);
or U8430 (N_8430,N_4033,N_2976);
or U8431 (N_8431,N_4327,N_826);
nor U8432 (N_8432,N_893,N_87);
xnor U8433 (N_8433,N_3170,N_1144);
nor U8434 (N_8434,N_4821,N_1828);
nand U8435 (N_8435,N_3371,N_4841);
nand U8436 (N_8436,N_3107,N_212);
or U8437 (N_8437,N_4600,N_3821);
nor U8438 (N_8438,N_4356,N_4866);
and U8439 (N_8439,N_1962,N_3073);
nor U8440 (N_8440,N_2958,N_3339);
nand U8441 (N_8441,N_304,N_3834);
nor U8442 (N_8442,N_3365,N_2225);
nor U8443 (N_8443,N_3275,N_4429);
xnor U8444 (N_8444,N_1551,N_1762);
and U8445 (N_8445,N_4237,N_1084);
and U8446 (N_8446,N_1936,N_4584);
nand U8447 (N_8447,N_372,N_3394);
or U8448 (N_8448,N_4725,N_4629);
nor U8449 (N_8449,N_3692,N_1708);
and U8450 (N_8450,N_4500,N_3820);
nor U8451 (N_8451,N_3082,N_2001);
and U8452 (N_8452,N_3948,N_3610);
nand U8453 (N_8453,N_1593,N_381);
and U8454 (N_8454,N_3548,N_2731);
nand U8455 (N_8455,N_1769,N_88);
nand U8456 (N_8456,N_1170,N_3444);
nor U8457 (N_8457,N_1615,N_718);
and U8458 (N_8458,N_841,N_3277);
and U8459 (N_8459,N_4198,N_3798);
nor U8460 (N_8460,N_2009,N_213);
and U8461 (N_8461,N_1124,N_2882);
nand U8462 (N_8462,N_781,N_3724);
and U8463 (N_8463,N_2298,N_1102);
nor U8464 (N_8464,N_4563,N_368);
nand U8465 (N_8465,N_1448,N_4151);
or U8466 (N_8466,N_3891,N_2095);
nor U8467 (N_8467,N_1698,N_2629);
nand U8468 (N_8468,N_1687,N_698);
and U8469 (N_8469,N_296,N_1489);
and U8470 (N_8470,N_3840,N_4767);
and U8471 (N_8471,N_3146,N_3116);
nor U8472 (N_8472,N_832,N_1429);
or U8473 (N_8473,N_3499,N_2455);
or U8474 (N_8474,N_4448,N_2582);
or U8475 (N_8475,N_4933,N_2830);
and U8476 (N_8476,N_4693,N_2957);
nand U8477 (N_8477,N_4749,N_705);
or U8478 (N_8478,N_3033,N_1546);
nand U8479 (N_8479,N_1066,N_1397);
nor U8480 (N_8480,N_3418,N_3891);
xor U8481 (N_8481,N_3439,N_3092);
and U8482 (N_8482,N_1583,N_615);
nand U8483 (N_8483,N_4000,N_3160);
and U8484 (N_8484,N_1264,N_1064);
nand U8485 (N_8485,N_3265,N_3361);
nand U8486 (N_8486,N_3714,N_2104);
nor U8487 (N_8487,N_4061,N_3285);
nand U8488 (N_8488,N_1886,N_4889);
and U8489 (N_8489,N_592,N_2484);
and U8490 (N_8490,N_4529,N_3478);
nand U8491 (N_8491,N_2068,N_69);
nor U8492 (N_8492,N_2890,N_3382);
or U8493 (N_8493,N_4019,N_4793);
and U8494 (N_8494,N_1468,N_4755);
nand U8495 (N_8495,N_4439,N_3762);
xnor U8496 (N_8496,N_2047,N_3055);
nand U8497 (N_8497,N_256,N_618);
nor U8498 (N_8498,N_3272,N_703);
or U8499 (N_8499,N_557,N_3937);
and U8500 (N_8500,N_2764,N_4276);
nand U8501 (N_8501,N_3498,N_3699);
or U8502 (N_8502,N_1704,N_2008);
and U8503 (N_8503,N_87,N_2017);
and U8504 (N_8504,N_1545,N_1134);
nand U8505 (N_8505,N_2261,N_3354);
and U8506 (N_8506,N_4978,N_585);
or U8507 (N_8507,N_2084,N_2081);
or U8508 (N_8508,N_1905,N_423);
nand U8509 (N_8509,N_4246,N_450);
or U8510 (N_8510,N_3105,N_4214);
or U8511 (N_8511,N_3834,N_2959);
and U8512 (N_8512,N_4730,N_3767);
nor U8513 (N_8513,N_4807,N_422);
and U8514 (N_8514,N_3296,N_620);
xnor U8515 (N_8515,N_3241,N_4908);
xor U8516 (N_8516,N_3390,N_4592);
and U8517 (N_8517,N_4524,N_524);
or U8518 (N_8518,N_397,N_1343);
and U8519 (N_8519,N_940,N_1319);
or U8520 (N_8520,N_3539,N_2732);
or U8521 (N_8521,N_4972,N_138);
or U8522 (N_8522,N_1981,N_2047);
and U8523 (N_8523,N_1109,N_397);
or U8524 (N_8524,N_1653,N_2145);
nor U8525 (N_8525,N_3553,N_989);
and U8526 (N_8526,N_4914,N_3097);
nor U8527 (N_8527,N_4897,N_797);
and U8528 (N_8528,N_4324,N_608);
nand U8529 (N_8529,N_3891,N_3215);
nor U8530 (N_8530,N_2482,N_35);
or U8531 (N_8531,N_3408,N_4227);
or U8532 (N_8532,N_570,N_4659);
nor U8533 (N_8533,N_2870,N_3334);
nor U8534 (N_8534,N_1959,N_1502);
or U8535 (N_8535,N_1543,N_25);
nor U8536 (N_8536,N_2150,N_2895);
nor U8537 (N_8537,N_4231,N_1669);
nand U8538 (N_8538,N_1669,N_2549);
nand U8539 (N_8539,N_3506,N_1757);
nor U8540 (N_8540,N_2676,N_3349);
and U8541 (N_8541,N_1091,N_2465);
nor U8542 (N_8542,N_3339,N_848);
nand U8543 (N_8543,N_3255,N_2944);
nand U8544 (N_8544,N_2737,N_4208);
nand U8545 (N_8545,N_236,N_3998);
and U8546 (N_8546,N_3235,N_2920);
nor U8547 (N_8547,N_3305,N_3284);
nand U8548 (N_8548,N_4921,N_2943);
and U8549 (N_8549,N_739,N_1055);
nor U8550 (N_8550,N_3558,N_167);
nand U8551 (N_8551,N_149,N_1837);
nor U8552 (N_8552,N_3711,N_2943);
and U8553 (N_8553,N_1582,N_3265);
or U8554 (N_8554,N_1312,N_412);
or U8555 (N_8555,N_2410,N_3149);
and U8556 (N_8556,N_1174,N_1083);
or U8557 (N_8557,N_1388,N_1036);
and U8558 (N_8558,N_2647,N_2609);
nand U8559 (N_8559,N_2439,N_2613);
and U8560 (N_8560,N_2869,N_1166);
nand U8561 (N_8561,N_778,N_981);
and U8562 (N_8562,N_102,N_1450);
and U8563 (N_8563,N_3778,N_278);
and U8564 (N_8564,N_4772,N_1398);
nand U8565 (N_8565,N_391,N_4115);
and U8566 (N_8566,N_4884,N_2034);
nor U8567 (N_8567,N_3108,N_2556);
xor U8568 (N_8568,N_19,N_806);
nand U8569 (N_8569,N_4164,N_2423);
nor U8570 (N_8570,N_4410,N_3258);
nor U8571 (N_8571,N_2456,N_1392);
or U8572 (N_8572,N_857,N_305);
or U8573 (N_8573,N_4838,N_537);
and U8574 (N_8574,N_2181,N_3907);
or U8575 (N_8575,N_1783,N_2233);
nand U8576 (N_8576,N_369,N_1033);
and U8577 (N_8577,N_3228,N_1126);
and U8578 (N_8578,N_4721,N_1144);
and U8579 (N_8579,N_1022,N_678);
nor U8580 (N_8580,N_1347,N_2913);
and U8581 (N_8581,N_2001,N_3316);
and U8582 (N_8582,N_1569,N_2942);
nor U8583 (N_8583,N_4394,N_315);
or U8584 (N_8584,N_3195,N_1097);
nand U8585 (N_8585,N_4998,N_4422);
nand U8586 (N_8586,N_336,N_2157);
or U8587 (N_8587,N_2426,N_1336);
or U8588 (N_8588,N_4712,N_42);
nand U8589 (N_8589,N_4469,N_4658);
nand U8590 (N_8590,N_465,N_4586);
xor U8591 (N_8591,N_1275,N_2044);
and U8592 (N_8592,N_4452,N_3944);
nor U8593 (N_8593,N_471,N_3856);
or U8594 (N_8594,N_2976,N_3517);
or U8595 (N_8595,N_4477,N_3388);
and U8596 (N_8596,N_4522,N_1500);
and U8597 (N_8597,N_173,N_2262);
nor U8598 (N_8598,N_3908,N_2047);
and U8599 (N_8599,N_2936,N_4716);
xnor U8600 (N_8600,N_997,N_3426);
and U8601 (N_8601,N_4575,N_35);
and U8602 (N_8602,N_4801,N_1487);
nand U8603 (N_8603,N_3089,N_1);
and U8604 (N_8604,N_1520,N_3957);
and U8605 (N_8605,N_3120,N_838);
and U8606 (N_8606,N_4299,N_751);
or U8607 (N_8607,N_1751,N_4596);
nor U8608 (N_8608,N_3586,N_3218);
nand U8609 (N_8609,N_4142,N_804);
nor U8610 (N_8610,N_1254,N_3530);
or U8611 (N_8611,N_3562,N_1231);
and U8612 (N_8612,N_1241,N_904);
nor U8613 (N_8613,N_2916,N_1042);
or U8614 (N_8614,N_710,N_3958);
nor U8615 (N_8615,N_4482,N_2829);
nand U8616 (N_8616,N_2091,N_1369);
or U8617 (N_8617,N_3702,N_4184);
and U8618 (N_8618,N_3670,N_3275);
or U8619 (N_8619,N_52,N_3916);
and U8620 (N_8620,N_44,N_3502);
and U8621 (N_8621,N_1671,N_867);
and U8622 (N_8622,N_3107,N_3044);
or U8623 (N_8623,N_2009,N_4861);
nor U8624 (N_8624,N_668,N_2532);
nor U8625 (N_8625,N_3387,N_2431);
or U8626 (N_8626,N_1251,N_3860);
and U8627 (N_8627,N_3874,N_28);
nand U8628 (N_8628,N_3524,N_4620);
nand U8629 (N_8629,N_1529,N_948);
nor U8630 (N_8630,N_1454,N_4300);
nand U8631 (N_8631,N_1541,N_1701);
nor U8632 (N_8632,N_4284,N_2900);
nor U8633 (N_8633,N_4734,N_882);
nor U8634 (N_8634,N_1791,N_193);
nor U8635 (N_8635,N_1877,N_3736);
nand U8636 (N_8636,N_2435,N_1638);
or U8637 (N_8637,N_1061,N_3587);
nand U8638 (N_8638,N_1904,N_910);
or U8639 (N_8639,N_4072,N_3008);
nor U8640 (N_8640,N_2358,N_4510);
nand U8641 (N_8641,N_492,N_1839);
and U8642 (N_8642,N_1578,N_1691);
nand U8643 (N_8643,N_1583,N_1795);
nand U8644 (N_8644,N_535,N_2404);
and U8645 (N_8645,N_1879,N_4029);
and U8646 (N_8646,N_626,N_3924);
and U8647 (N_8647,N_4211,N_398);
and U8648 (N_8648,N_974,N_4172);
nand U8649 (N_8649,N_4100,N_907);
or U8650 (N_8650,N_4412,N_4809);
or U8651 (N_8651,N_4309,N_3010);
nand U8652 (N_8652,N_509,N_1910);
and U8653 (N_8653,N_6,N_2869);
nand U8654 (N_8654,N_4293,N_1796);
and U8655 (N_8655,N_3041,N_4767);
nand U8656 (N_8656,N_155,N_1365);
nand U8657 (N_8657,N_4518,N_886);
and U8658 (N_8658,N_4983,N_2181);
nor U8659 (N_8659,N_4992,N_4190);
nor U8660 (N_8660,N_2503,N_3273);
nor U8661 (N_8661,N_104,N_3639);
or U8662 (N_8662,N_2045,N_446);
nand U8663 (N_8663,N_3238,N_3179);
nor U8664 (N_8664,N_2033,N_2708);
nand U8665 (N_8665,N_703,N_337);
or U8666 (N_8666,N_3681,N_1081);
and U8667 (N_8667,N_3180,N_2015);
xor U8668 (N_8668,N_3370,N_1512);
or U8669 (N_8669,N_3174,N_4205);
nor U8670 (N_8670,N_968,N_3954);
nand U8671 (N_8671,N_1511,N_4781);
or U8672 (N_8672,N_1287,N_2050);
nor U8673 (N_8673,N_937,N_4377);
nand U8674 (N_8674,N_4439,N_1730);
nor U8675 (N_8675,N_1214,N_4255);
and U8676 (N_8676,N_3211,N_3283);
nand U8677 (N_8677,N_2338,N_898);
or U8678 (N_8678,N_1957,N_2777);
nand U8679 (N_8679,N_766,N_646);
nand U8680 (N_8680,N_3146,N_1198);
or U8681 (N_8681,N_841,N_3268);
nand U8682 (N_8682,N_660,N_411);
or U8683 (N_8683,N_481,N_4297);
nand U8684 (N_8684,N_2221,N_3617);
nor U8685 (N_8685,N_4616,N_2451);
nand U8686 (N_8686,N_3402,N_1489);
or U8687 (N_8687,N_3809,N_539);
and U8688 (N_8688,N_729,N_4927);
and U8689 (N_8689,N_1794,N_4395);
nand U8690 (N_8690,N_1498,N_3592);
and U8691 (N_8691,N_1057,N_1146);
nand U8692 (N_8692,N_2538,N_3703);
and U8693 (N_8693,N_166,N_1953);
nor U8694 (N_8694,N_1600,N_156);
or U8695 (N_8695,N_577,N_1858);
or U8696 (N_8696,N_3205,N_280);
and U8697 (N_8697,N_3164,N_1344);
nand U8698 (N_8698,N_254,N_1758);
nor U8699 (N_8699,N_1374,N_2957);
nor U8700 (N_8700,N_1723,N_3414);
nor U8701 (N_8701,N_2440,N_283);
or U8702 (N_8702,N_270,N_1675);
nand U8703 (N_8703,N_3712,N_52);
xnor U8704 (N_8704,N_3867,N_1140);
nand U8705 (N_8705,N_2430,N_2241);
nand U8706 (N_8706,N_1153,N_2287);
or U8707 (N_8707,N_4109,N_473);
nand U8708 (N_8708,N_3684,N_3354);
or U8709 (N_8709,N_2275,N_1478);
or U8710 (N_8710,N_4342,N_3932);
or U8711 (N_8711,N_1187,N_955);
nor U8712 (N_8712,N_202,N_1473);
or U8713 (N_8713,N_668,N_1073);
nand U8714 (N_8714,N_1237,N_2759);
or U8715 (N_8715,N_613,N_4607);
nor U8716 (N_8716,N_2848,N_4219);
nor U8717 (N_8717,N_1698,N_1672);
nor U8718 (N_8718,N_4633,N_2868);
nor U8719 (N_8719,N_251,N_2698);
nand U8720 (N_8720,N_4201,N_4702);
and U8721 (N_8721,N_1842,N_712);
nand U8722 (N_8722,N_2752,N_991);
nor U8723 (N_8723,N_2988,N_3499);
nand U8724 (N_8724,N_1780,N_283);
or U8725 (N_8725,N_4304,N_3254);
nor U8726 (N_8726,N_2637,N_4983);
nor U8727 (N_8727,N_1261,N_2639);
or U8728 (N_8728,N_1145,N_4963);
nand U8729 (N_8729,N_3120,N_699);
and U8730 (N_8730,N_3690,N_4270);
nor U8731 (N_8731,N_917,N_3965);
or U8732 (N_8732,N_3399,N_1449);
and U8733 (N_8733,N_1208,N_3661);
nand U8734 (N_8734,N_3284,N_3785);
or U8735 (N_8735,N_2916,N_2421);
nand U8736 (N_8736,N_4943,N_2522);
nand U8737 (N_8737,N_811,N_1864);
nor U8738 (N_8738,N_430,N_2053);
or U8739 (N_8739,N_890,N_4617);
nand U8740 (N_8740,N_1731,N_3025);
or U8741 (N_8741,N_1375,N_3227);
nand U8742 (N_8742,N_2729,N_1383);
nor U8743 (N_8743,N_3123,N_2146);
nand U8744 (N_8744,N_1234,N_1352);
nand U8745 (N_8745,N_2975,N_63);
and U8746 (N_8746,N_1256,N_554);
and U8747 (N_8747,N_4586,N_4500);
or U8748 (N_8748,N_1312,N_4186);
nand U8749 (N_8749,N_372,N_4901);
nand U8750 (N_8750,N_190,N_2088);
nand U8751 (N_8751,N_2133,N_353);
and U8752 (N_8752,N_3607,N_2118);
nor U8753 (N_8753,N_3205,N_4981);
nand U8754 (N_8754,N_4258,N_758);
nor U8755 (N_8755,N_1061,N_3672);
nand U8756 (N_8756,N_1123,N_498);
nand U8757 (N_8757,N_4601,N_3061);
nand U8758 (N_8758,N_1659,N_4668);
nand U8759 (N_8759,N_139,N_4293);
or U8760 (N_8760,N_3901,N_1347);
and U8761 (N_8761,N_3135,N_3409);
and U8762 (N_8762,N_1363,N_439);
nand U8763 (N_8763,N_4689,N_1706);
nand U8764 (N_8764,N_1528,N_3547);
nor U8765 (N_8765,N_1942,N_4326);
nor U8766 (N_8766,N_975,N_2988);
or U8767 (N_8767,N_1084,N_4656);
and U8768 (N_8768,N_242,N_981);
nor U8769 (N_8769,N_3102,N_1745);
nor U8770 (N_8770,N_1146,N_520);
or U8771 (N_8771,N_4350,N_531);
and U8772 (N_8772,N_1927,N_3214);
nand U8773 (N_8773,N_3472,N_4062);
nor U8774 (N_8774,N_2902,N_2004);
xnor U8775 (N_8775,N_3647,N_228);
and U8776 (N_8776,N_2887,N_364);
nand U8777 (N_8777,N_2256,N_1067);
or U8778 (N_8778,N_507,N_1371);
nor U8779 (N_8779,N_4817,N_1586);
nand U8780 (N_8780,N_1557,N_4413);
and U8781 (N_8781,N_3815,N_4357);
and U8782 (N_8782,N_3861,N_3138);
or U8783 (N_8783,N_1365,N_4543);
nor U8784 (N_8784,N_3046,N_4162);
and U8785 (N_8785,N_2895,N_380);
and U8786 (N_8786,N_4485,N_925);
and U8787 (N_8787,N_4782,N_43);
and U8788 (N_8788,N_1033,N_3575);
nor U8789 (N_8789,N_1525,N_3677);
nand U8790 (N_8790,N_3959,N_4238);
nand U8791 (N_8791,N_2832,N_3613);
or U8792 (N_8792,N_1581,N_2859);
or U8793 (N_8793,N_1560,N_4995);
and U8794 (N_8794,N_749,N_4114);
nand U8795 (N_8795,N_3022,N_1234);
nand U8796 (N_8796,N_759,N_1907);
and U8797 (N_8797,N_3971,N_2204);
nor U8798 (N_8798,N_26,N_1082);
xnor U8799 (N_8799,N_4104,N_2402);
or U8800 (N_8800,N_4761,N_441);
nor U8801 (N_8801,N_3279,N_2930);
and U8802 (N_8802,N_4982,N_3450);
xor U8803 (N_8803,N_2224,N_2012);
or U8804 (N_8804,N_755,N_1498);
nor U8805 (N_8805,N_2127,N_3906);
nor U8806 (N_8806,N_3734,N_450);
nor U8807 (N_8807,N_2138,N_1126);
nand U8808 (N_8808,N_680,N_2896);
or U8809 (N_8809,N_2493,N_3322);
nand U8810 (N_8810,N_4949,N_4833);
and U8811 (N_8811,N_4363,N_2738);
nor U8812 (N_8812,N_782,N_4192);
and U8813 (N_8813,N_4732,N_4115);
and U8814 (N_8814,N_3237,N_2562);
or U8815 (N_8815,N_4234,N_2108);
and U8816 (N_8816,N_4763,N_1726);
or U8817 (N_8817,N_1063,N_3918);
nor U8818 (N_8818,N_4368,N_3082);
and U8819 (N_8819,N_2597,N_2408);
nor U8820 (N_8820,N_333,N_1296);
or U8821 (N_8821,N_2050,N_4442);
nor U8822 (N_8822,N_2128,N_2426);
nor U8823 (N_8823,N_4404,N_4319);
or U8824 (N_8824,N_740,N_2450);
nand U8825 (N_8825,N_1370,N_3821);
nor U8826 (N_8826,N_711,N_4355);
or U8827 (N_8827,N_783,N_2600);
and U8828 (N_8828,N_1717,N_4568);
or U8829 (N_8829,N_1952,N_4153);
nor U8830 (N_8830,N_2275,N_1174);
nand U8831 (N_8831,N_2264,N_2054);
and U8832 (N_8832,N_4869,N_2972);
and U8833 (N_8833,N_4666,N_711);
nor U8834 (N_8834,N_2227,N_350);
nand U8835 (N_8835,N_3704,N_3737);
or U8836 (N_8836,N_2918,N_2125);
nand U8837 (N_8837,N_473,N_115);
and U8838 (N_8838,N_1425,N_3843);
or U8839 (N_8839,N_547,N_303);
and U8840 (N_8840,N_4929,N_740);
nand U8841 (N_8841,N_736,N_2561);
and U8842 (N_8842,N_4899,N_4931);
nor U8843 (N_8843,N_2920,N_3806);
nor U8844 (N_8844,N_2106,N_4749);
or U8845 (N_8845,N_3489,N_2141);
nand U8846 (N_8846,N_3602,N_3924);
or U8847 (N_8847,N_1171,N_1211);
nand U8848 (N_8848,N_2233,N_2368);
nand U8849 (N_8849,N_3152,N_3184);
nand U8850 (N_8850,N_4488,N_4606);
nor U8851 (N_8851,N_3840,N_3850);
nand U8852 (N_8852,N_526,N_344);
and U8853 (N_8853,N_2792,N_268);
or U8854 (N_8854,N_1112,N_3313);
and U8855 (N_8855,N_540,N_382);
or U8856 (N_8856,N_1925,N_743);
nor U8857 (N_8857,N_198,N_3883);
nand U8858 (N_8858,N_3966,N_2079);
and U8859 (N_8859,N_830,N_3982);
nor U8860 (N_8860,N_2945,N_4691);
and U8861 (N_8861,N_1039,N_3416);
nand U8862 (N_8862,N_2414,N_4939);
nor U8863 (N_8863,N_4825,N_3780);
nand U8864 (N_8864,N_521,N_3976);
or U8865 (N_8865,N_1554,N_698);
nor U8866 (N_8866,N_2251,N_226);
and U8867 (N_8867,N_3695,N_754);
and U8868 (N_8868,N_427,N_898);
nor U8869 (N_8869,N_939,N_3626);
nand U8870 (N_8870,N_37,N_586);
nand U8871 (N_8871,N_4084,N_2814);
nor U8872 (N_8872,N_4383,N_2497);
or U8873 (N_8873,N_221,N_1267);
or U8874 (N_8874,N_1876,N_1288);
nor U8875 (N_8875,N_2137,N_4344);
and U8876 (N_8876,N_3044,N_3439);
and U8877 (N_8877,N_4867,N_3144);
or U8878 (N_8878,N_1349,N_469);
nand U8879 (N_8879,N_1963,N_2224);
nor U8880 (N_8880,N_3237,N_3848);
and U8881 (N_8881,N_419,N_4816);
nor U8882 (N_8882,N_4352,N_226);
nand U8883 (N_8883,N_3401,N_2920);
nand U8884 (N_8884,N_1360,N_1613);
nand U8885 (N_8885,N_644,N_1087);
xnor U8886 (N_8886,N_1017,N_2256);
and U8887 (N_8887,N_4000,N_3806);
or U8888 (N_8888,N_51,N_1006);
nor U8889 (N_8889,N_2938,N_4016);
nor U8890 (N_8890,N_2405,N_3700);
nand U8891 (N_8891,N_1591,N_3175);
nor U8892 (N_8892,N_4533,N_3943);
nor U8893 (N_8893,N_2616,N_4499);
xnor U8894 (N_8894,N_379,N_2009);
nor U8895 (N_8895,N_4409,N_3273);
and U8896 (N_8896,N_1369,N_858);
or U8897 (N_8897,N_668,N_4902);
and U8898 (N_8898,N_4642,N_2574);
nor U8899 (N_8899,N_2747,N_1589);
nand U8900 (N_8900,N_1716,N_4649);
and U8901 (N_8901,N_3890,N_814);
nand U8902 (N_8902,N_2149,N_1580);
nor U8903 (N_8903,N_4039,N_4746);
nand U8904 (N_8904,N_4495,N_3364);
or U8905 (N_8905,N_3650,N_1890);
or U8906 (N_8906,N_1387,N_140);
or U8907 (N_8907,N_233,N_3710);
nor U8908 (N_8908,N_97,N_1464);
nor U8909 (N_8909,N_2851,N_96);
and U8910 (N_8910,N_2367,N_3996);
or U8911 (N_8911,N_2676,N_3106);
and U8912 (N_8912,N_2124,N_1858);
nor U8913 (N_8913,N_3972,N_2304);
nand U8914 (N_8914,N_3464,N_2687);
or U8915 (N_8915,N_1872,N_4269);
or U8916 (N_8916,N_4244,N_295);
xor U8917 (N_8917,N_750,N_2361);
nor U8918 (N_8918,N_4628,N_3797);
or U8919 (N_8919,N_101,N_4627);
nor U8920 (N_8920,N_73,N_4534);
and U8921 (N_8921,N_3064,N_224);
and U8922 (N_8922,N_4595,N_1399);
nand U8923 (N_8923,N_2369,N_2257);
nand U8924 (N_8924,N_2736,N_669);
nor U8925 (N_8925,N_3540,N_1857);
nor U8926 (N_8926,N_1597,N_1013);
nand U8927 (N_8927,N_228,N_1996);
nand U8928 (N_8928,N_253,N_2807);
nand U8929 (N_8929,N_2180,N_1105);
nand U8930 (N_8930,N_3320,N_1177);
nand U8931 (N_8931,N_1586,N_3997);
nor U8932 (N_8932,N_678,N_2488);
and U8933 (N_8933,N_2747,N_4834);
nor U8934 (N_8934,N_459,N_4382);
and U8935 (N_8935,N_1049,N_850);
or U8936 (N_8936,N_1759,N_1749);
or U8937 (N_8937,N_4518,N_2747);
xnor U8938 (N_8938,N_3710,N_2183);
nor U8939 (N_8939,N_274,N_958);
nand U8940 (N_8940,N_3320,N_1408);
or U8941 (N_8941,N_228,N_4796);
nand U8942 (N_8942,N_4770,N_2634);
and U8943 (N_8943,N_3637,N_351);
or U8944 (N_8944,N_195,N_3001);
nand U8945 (N_8945,N_4673,N_1803);
nand U8946 (N_8946,N_1460,N_4400);
nand U8947 (N_8947,N_2264,N_1374);
nor U8948 (N_8948,N_2196,N_898);
nand U8949 (N_8949,N_1856,N_1653);
or U8950 (N_8950,N_2092,N_4929);
nor U8951 (N_8951,N_954,N_2185);
nand U8952 (N_8952,N_1911,N_314);
nor U8953 (N_8953,N_3578,N_1403);
nand U8954 (N_8954,N_1850,N_1558);
or U8955 (N_8955,N_650,N_3939);
and U8956 (N_8956,N_2027,N_3594);
nor U8957 (N_8957,N_4560,N_177);
or U8958 (N_8958,N_3555,N_4924);
and U8959 (N_8959,N_4395,N_4545);
and U8960 (N_8960,N_375,N_1588);
nor U8961 (N_8961,N_4731,N_1283);
or U8962 (N_8962,N_2376,N_1859);
or U8963 (N_8963,N_4880,N_3751);
or U8964 (N_8964,N_2574,N_800);
nand U8965 (N_8965,N_4608,N_1646);
nor U8966 (N_8966,N_2841,N_805);
and U8967 (N_8967,N_4466,N_2628);
nand U8968 (N_8968,N_2901,N_4744);
nor U8969 (N_8969,N_2536,N_114);
and U8970 (N_8970,N_1601,N_904);
and U8971 (N_8971,N_1272,N_2292);
nand U8972 (N_8972,N_4932,N_4606);
nand U8973 (N_8973,N_2168,N_1153);
or U8974 (N_8974,N_2230,N_1105);
nand U8975 (N_8975,N_1472,N_3012);
and U8976 (N_8976,N_1462,N_2056);
nor U8977 (N_8977,N_4300,N_3775);
and U8978 (N_8978,N_903,N_4188);
nand U8979 (N_8979,N_4385,N_1204);
or U8980 (N_8980,N_418,N_3970);
and U8981 (N_8981,N_3336,N_4267);
and U8982 (N_8982,N_4622,N_2899);
nor U8983 (N_8983,N_4720,N_3748);
or U8984 (N_8984,N_2811,N_373);
nand U8985 (N_8985,N_3394,N_4702);
nand U8986 (N_8986,N_249,N_1153);
or U8987 (N_8987,N_3071,N_3733);
xor U8988 (N_8988,N_4364,N_2699);
or U8989 (N_8989,N_4478,N_3751);
nand U8990 (N_8990,N_1469,N_3396);
and U8991 (N_8991,N_1227,N_2583);
nand U8992 (N_8992,N_3336,N_2338);
or U8993 (N_8993,N_3424,N_4288);
or U8994 (N_8994,N_4323,N_3547);
nor U8995 (N_8995,N_3002,N_1962);
nand U8996 (N_8996,N_1504,N_3775);
nor U8997 (N_8997,N_1432,N_4700);
or U8998 (N_8998,N_2616,N_1924);
nand U8999 (N_8999,N_3339,N_4408);
nor U9000 (N_9000,N_4760,N_3258);
or U9001 (N_9001,N_2149,N_3627);
and U9002 (N_9002,N_2641,N_2575);
nand U9003 (N_9003,N_1912,N_1334);
or U9004 (N_9004,N_794,N_1063);
nand U9005 (N_9005,N_4377,N_1577);
nor U9006 (N_9006,N_980,N_2305);
nand U9007 (N_9007,N_4898,N_2727);
nor U9008 (N_9008,N_1882,N_3245);
or U9009 (N_9009,N_326,N_3527);
or U9010 (N_9010,N_3986,N_316);
and U9011 (N_9011,N_840,N_4950);
nand U9012 (N_9012,N_2434,N_2444);
nand U9013 (N_9013,N_1293,N_1379);
nor U9014 (N_9014,N_3654,N_562);
nor U9015 (N_9015,N_377,N_4723);
and U9016 (N_9016,N_4834,N_3807);
nor U9017 (N_9017,N_973,N_1749);
nand U9018 (N_9018,N_723,N_1175);
or U9019 (N_9019,N_3611,N_503);
nand U9020 (N_9020,N_4472,N_802);
and U9021 (N_9021,N_4613,N_3014);
or U9022 (N_9022,N_1913,N_1138);
nor U9023 (N_9023,N_410,N_3333);
nand U9024 (N_9024,N_998,N_2040);
nor U9025 (N_9025,N_4786,N_2250);
and U9026 (N_9026,N_4361,N_4017);
or U9027 (N_9027,N_2416,N_39);
nand U9028 (N_9028,N_3802,N_3771);
and U9029 (N_9029,N_2372,N_1152);
nor U9030 (N_9030,N_157,N_4260);
xnor U9031 (N_9031,N_1447,N_3598);
and U9032 (N_9032,N_4693,N_2963);
nand U9033 (N_9033,N_3672,N_2687);
nand U9034 (N_9034,N_1750,N_3692);
nor U9035 (N_9035,N_1213,N_4055);
nand U9036 (N_9036,N_262,N_2887);
or U9037 (N_9037,N_2911,N_4150);
nand U9038 (N_9038,N_1978,N_4184);
nor U9039 (N_9039,N_4585,N_3842);
nand U9040 (N_9040,N_2304,N_1303);
nor U9041 (N_9041,N_1910,N_3167);
nand U9042 (N_9042,N_3436,N_3636);
nand U9043 (N_9043,N_1260,N_4984);
and U9044 (N_9044,N_2177,N_4185);
nand U9045 (N_9045,N_765,N_2667);
and U9046 (N_9046,N_3550,N_1560);
nand U9047 (N_9047,N_974,N_1261);
nor U9048 (N_9048,N_1546,N_431);
and U9049 (N_9049,N_2268,N_41);
nor U9050 (N_9050,N_77,N_3399);
and U9051 (N_9051,N_4382,N_1471);
or U9052 (N_9052,N_787,N_4563);
nor U9053 (N_9053,N_698,N_1912);
nor U9054 (N_9054,N_4840,N_3679);
nor U9055 (N_9055,N_3005,N_3116);
nand U9056 (N_9056,N_1696,N_5);
nor U9057 (N_9057,N_4958,N_2484);
nor U9058 (N_9058,N_1520,N_1409);
nor U9059 (N_9059,N_3363,N_479);
nand U9060 (N_9060,N_2655,N_3623);
nand U9061 (N_9061,N_2976,N_1892);
and U9062 (N_9062,N_2293,N_1097);
and U9063 (N_9063,N_1610,N_300);
or U9064 (N_9064,N_1137,N_1126);
or U9065 (N_9065,N_3770,N_995);
nor U9066 (N_9066,N_236,N_2297);
nor U9067 (N_9067,N_4333,N_3999);
or U9068 (N_9068,N_1819,N_2671);
nor U9069 (N_9069,N_2118,N_1682);
or U9070 (N_9070,N_1809,N_1418);
nand U9071 (N_9071,N_2263,N_486);
nor U9072 (N_9072,N_3152,N_3246);
nor U9073 (N_9073,N_677,N_1294);
nor U9074 (N_9074,N_975,N_2876);
and U9075 (N_9075,N_576,N_3321);
and U9076 (N_9076,N_84,N_3894);
nand U9077 (N_9077,N_3494,N_4992);
nand U9078 (N_9078,N_2203,N_4164);
and U9079 (N_9079,N_4517,N_1208);
or U9080 (N_9080,N_2639,N_1220);
nand U9081 (N_9081,N_1455,N_3698);
and U9082 (N_9082,N_1554,N_3492);
nor U9083 (N_9083,N_116,N_1987);
nor U9084 (N_9084,N_3805,N_2155);
or U9085 (N_9085,N_3967,N_1003);
nor U9086 (N_9086,N_4321,N_3896);
nand U9087 (N_9087,N_2101,N_2861);
and U9088 (N_9088,N_3522,N_794);
or U9089 (N_9089,N_3178,N_2089);
and U9090 (N_9090,N_1487,N_530);
xor U9091 (N_9091,N_809,N_3888);
nand U9092 (N_9092,N_910,N_797);
or U9093 (N_9093,N_34,N_4173);
or U9094 (N_9094,N_4507,N_944);
and U9095 (N_9095,N_4123,N_4168);
nor U9096 (N_9096,N_3416,N_4275);
nor U9097 (N_9097,N_2768,N_1138);
xnor U9098 (N_9098,N_4723,N_2581);
xor U9099 (N_9099,N_4046,N_3250);
or U9100 (N_9100,N_3006,N_4752);
or U9101 (N_9101,N_3731,N_4850);
nand U9102 (N_9102,N_3030,N_3733);
nand U9103 (N_9103,N_1213,N_4792);
or U9104 (N_9104,N_3646,N_3815);
and U9105 (N_9105,N_1550,N_103);
or U9106 (N_9106,N_2315,N_3443);
and U9107 (N_9107,N_3212,N_107);
nand U9108 (N_9108,N_4767,N_2491);
and U9109 (N_9109,N_4126,N_159);
nor U9110 (N_9110,N_3114,N_2507);
nor U9111 (N_9111,N_1495,N_3235);
and U9112 (N_9112,N_3946,N_1170);
nor U9113 (N_9113,N_3547,N_1255);
nor U9114 (N_9114,N_4781,N_2472);
or U9115 (N_9115,N_2687,N_1822);
or U9116 (N_9116,N_4061,N_4125);
nor U9117 (N_9117,N_801,N_3823);
nand U9118 (N_9118,N_4814,N_3721);
nand U9119 (N_9119,N_878,N_2424);
nand U9120 (N_9120,N_560,N_2744);
nor U9121 (N_9121,N_4030,N_3023);
nand U9122 (N_9122,N_8,N_3941);
nand U9123 (N_9123,N_508,N_2206);
and U9124 (N_9124,N_4772,N_945);
nor U9125 (N_9125,N_167,N_1208);
nand U9126 (N_9126,N_3728,N_1746);
nand U9127 (N_9127,N_2925,N_1400);
or U9128 (N_9128,N_935,N_1010);
nand U9129 (N_9129,N_3103,N_394);
nand U9130 (N_9130,N_3492,N_4583);
and U9131 (N_9131,N_3716,N_2015);
and U9132 (N_9132,N_2034,N_3132);
nand U9133 (N_9133,N_3073,N_654);
and U9134 (N_9134,N_4411,N_4958);
and U9135 (N_9135,N_2315,N_2660);
nor U9136 (N_9136,N_4092,N_3349);
nor U9137 (N_9137,N_932,N_1144);
nand U9138 (N_9138,N_4008,N_4642);
or U9139 (N_9139,N_3763,N_2428);
nand U9140 (N_9140,N_4572,N_2473);
nor U9141 (N_9141,N_592,N_1967);
nand U9142 (N_9142,N_2934,N_4314);
and U9143 (N_9143,N_1146,N_231);
nand U9144 (N_9144,N_4767,N_576);
or U9145 (N_9145,N_867,N_1584);
and U9146 (N_9146,N_2865,N_2964);
or U9147 (N_9147,N_2464,N_674);
nor U9148 (N_9148,N_765,N_912);
nand U9149 (N_9149,N_3327,N_128);
or U9150 (N_9150,N_766,N_3009);
nor U9151 (N_9151,N_3387,N_781);
nor U9152 (N_9152,N_3734,N_3358);
nor U9153 (N_9153,N_1013,N_1449);
nand U9154 (N_9154,N_4580,N_961);
nor U9155 (N_9155,N_1588,N_130);
nand U9156 (N_9156,N_2910,N_3305);
and U9157 (N_9157,N_2230,N_2936);
nor U9158 (N_9158,N_1200,N_1375);
nor U9159 (N_9159,N_206,N_993);
or U9160 (N_9160,N_1285,N_784);
and U9161 (N_9161,N_4899,N_2755);
nor U9162 (N_9162,N_838,N_2735);
nor U9163 (N_9163,N_4314,N_2028);
and U9164 (N_9164,N_508,N_202);
nor U9165 (N_9165,N_1722,N_3418);
xor U9166 (N_9166,N_139,N_4688);
nand U9167 (N_9167,N_3267,N_1105);
nand U9168 (N_9168,N_700,N_3596);
or U9169 (N_9169,N_1251,N_4905);
nor U9170 (N_9170,N_1411,N_3316);
and U9171 (N_9171,N_3548,N_555);
nand U9172 (N_9172,N_3431,N_2480);
nor U9173 (N_9173,N_2832,N_4235);
or U9174 (N_9174,N_581,N_2709);
nor U9175 (N_9175,N_2704,N_4984);
and U9176 (N_9176,N_4313,N_4626);
nor U9177 (N_9177,N_47,N_4541);
nor U9178 (N_9178,N_1167,N_2364);
nand U9179 (N_9179,N_557,N_1241);
nor U9180 (N_9180,N_3590,N_3327);
nand U9181 (N_9181,N_2690,N_3931);
and U9182 (N_9182,N_2473,N_203);
nand U9183 (N_9183,N_2682,N_3322);
nand U9184 (N_9184,N_2369,N_2186);
or U9185 (N_9185,N_3487,N_961);
and U9186 (N_9186,N_771,N_4);
nand U9187 (N_9187,N_2709,N_4983);
nor U9188 (N_9188,N_3864,N_1274);
and U9189 (N_9189,N_1305,N_934);
or U9190 (N_9190,N_2542,N_1332);
nor U9191 (N_9191,N_679,N_670);
and U9192 (N_9192,N_811,N_2591);
or U9193 (N_9193,N_4719,N_3443);
or U9194 (N_9194,N_3070,N_4935);
and U9195 (N_9195,N_2207,N_4388);
nor U9196 (N_9196,N_1313,N_4700);
nor U9197 (N_9197,N_4489,N_1071);
and U9198 (N_9198,N_901,N_143);
nand U9199 (N_9199,N_1752,N_2608);
or U9200 (N_9200,N_3545,N_2251);
and U9201 (N_9201,N_3300,N_1447);
and U9202 (N_9202,N_597,N_748);
nor U9203 (N_9203,N_3393,N_3339);
or U9204 (N_9204,N_4530,N_1757);
nor U9205 (N_9205,N_1336,N_2786);
nand U9206 (N_9206,N_654,N_1448);
nor U9207 (N_9207,N_1413,N_2331);
and U9208 (N_9208,N_536,N_3316);
and U9209 (N_9209,N_4629,N_4524);
nor U9210 (N_9210,N_3778,N_4950);
nor U9211 (N_9211,N_2840,N_4864);
or U9212 (N_9212,N_1346,N_2769);
and U9213 (N_9213,N_4964,N_3791);
nand U9214 (N_9214,N_2410,N_2798);
xor U9215 (N_9215,N_4014,N_683);
or U9216 (N_9216,N_10,N_3825);
and U9217 (N_9217,N_4198,N_2127);
or U9218 (N_9218,N_3996,N_2389);
or U9219 (N_9219,N_67,N_2579);
nand U9220 (N_9220,N_3028,N_1957);
and U9221 (N_9221,N_2886,N_1816);
and U9222 (N_9222,N_2613,N_597);
xor U9223 (N_9223,N_1514,N_2999);
nor U9224 (N_9224,N_4671,N_3351);
or U9225 (N_9225,N_3982,N_2548);
nor U9226 (N_9226,N_502,N_3535);
nor U9227 (N_9227,N_372,N_2123);
nand U9228 (N_9228,N_2660,N_2729);
and U9229 (N_9229,N_731,N_4928);
nand U9230 (N_9230,N_87,N_1514);
and U9231 (N_9231,N_1150,N_3504);
or U9232 (N_9232,N_401,N_4601);
and U9233 (N_9233,N_1195,N_2390);
or U9234 (N_9234,N_685,N_860);
nand U9235 (N_9235,N_3845,N_660);
nand U9236 (N_9236,N_4047,N_4199);
nor U9237 (N_9237,N_4484,N_4181);
nand U9238 (N_9238,N_3665,N_3307);
and U9239 (N_9239,N_1646,N_3547);
nor U9240 (N_9240,N_2779,N_341);
nand U9241 (N_9241,N_3231,N_1624);
nand U9242 (N_9242,N_380,N_1354);
xor U9243 (N_9243,N_2857,N_2252);
nand U9244 (N_9244,N_449,N_4602);
or U9245 (N_9245,N_4747,N_3675);
and U9246 (N_9246,N_4808,N_3591);
xor U9247 (N_9247,N_4803,N_1922);
nand U9248 (N_9248,N_186,N_2272);
nor U9249 (N_9249,N_3521,N_1099);
nand U9250 (N_9250,N_4830,N_3436);
xor U9251 (N_9251,N_2277,N_746);
nand U9252 (N_9252,N_1052,N_1550);
nand U9253 (N_9253,N_596,N_348);
nand U9254 (N_9254,N_4985,N_3205);
nor U9255 (N_9255,N_661,N_2271);
or U9256 (N_9256,N_2321,N_3381);
nand U9257 (N_9257,N_2994,N_2160);
or U9258 (N_9258,N_337,N_127);
nand U9259 (N_9259,N_3227,N_3887);
xor U9260 (N_9260,N_15,N_2814);
or U9261 (N_9261,N_2433,N_3382);
nor U9262 (N_9262,N_1075,N_3659);
and U9263 (N_9263,N_3765,N_1383);
and U9264 (N_9264,N_2945,N_4891);
and U9265 (N_9265,N_1555,N_2761);
nand U9266 (N_9266,N_4209,N_4980);
and U9267 (N_9267,N_1754,N_2285);
or U9268 (N_9268,N_3162,N_1077);
nand U9269 (N_9269,N_13,N_2696);
or U9270 (N_9270,N_2915,N_1684);
xnor U9271 (N_9271,N_3804,N_4579);
or U9272 (N_9272,N_1985,N_4858);
nor U9273 (N_9273,N_4154,N_2461);
or U9274 (N_9274,N_1718,N_3930);
and U9275 (N_9275,N_507,N_54);
and U9276 (N_9276,N_4416,N_4850);
and U9277 (N_9277,N_2501,N_1009);
nor U9278 (N_9278,N_271,N_2946);
or U9279 (N_9279,N_2097,N_3049);
or U9280 (N_9280,N_123,N_1347);
and U9281 (N_9281,N_2893,N_1394);
nor U9282 (N_9282,N_1532,N_828);
nand U9283 (N_9283,N_710,N_2913);
and U9284 (N_9284,N_823,N_3246);
or U9285 (N_9285,N_4523,N_4302);
nand U9286 (N_9286,N_2394,N_632);
or U9287 (N_9287,N_4643,N_3947);
and U9288 (N_9288,N_6,N_2408);
nor U9289 (N_9289,N_4943,N_4321);
nand U9290 (N_9290,N_4630,N_3047);
and U9291 (N_9291,N_860,N_2870);
nor U9292 (N_9292,N_411,N_4110);
or U9293 (N_9293,N_381,N_3676);
and U9294 (N_9294,N_4058,N_906);
nor U9295 (N_9295,N_3017,N_1943);
xor U9296 (N_9296,N_2628,N_3495);
nand U9297 (N_9297,N_441,N_2547);
or U9298 (N_9298,N_1441,N_729);
or U9299 (N_9299,N_762,N_773);
nor U9300 (N_9300,N_3792,N_3883);
nand U9301 (N_9301,N_1211,N_3106);
and U9302 (N_9302,N_3856,N_3248);
and U9303 (N_9303,N_83,N_2208);
nor U9304 (N_9304,N_4889,N_1223);
nand U9305 (N_9305,N_2497,N_678);
nand U9306 (N_9306,N_1474,N_2222);
xor U9307 (N_9307,N_3286,N_3457);
or U9308 (N_9308,N_2372,N_1794);
nor U9309 (N_9309,N_3718,N_4558);
nor U9310 (N_9310,N_3576,N_565);
or U9311 (N_9311,N_3306,N_4412);
nand U9312 (N_9312,N_1136,N_4343);
nand U9313 (N_9313,N_753,N_3582);
and U9314 (N_9314,N_2399,N_854);
and U9315 (N_9315,N_1227,N_891);
nand U9316 (N_9316,N_3122,N_3615);
and U9317 (N_9317,N_1069,N_2227);
or U9318 (N_9318,N_1518,N_1320);
or U9319 (N_9319,N_4528,N_3715);
and U9320 (N_9320,N_2913,N_3788);
or U9321 (N_9321,N_1032,N_1262);
and U9322 (N_9322,N_648,N_570);
nand U9323 (N_9323,N_2641,N_3753);
nor U9324 (N_9324,N_345,N_830);
nand U9325 (N_9325,N_3069,N_1249);
or U9326 (N_9326,N_692,N_3763);
and U9327 (N_9327,N_3467,N_516);
nor U9328 (N_9328,N_1959,N_3501);
or U9329 (N_9329,N_4616,N_693);
nand U9330 (N_9330,N_2978,N_3056);
nand U9331 (N_9331,N_1129,N_735);
xor U9332 (N_9332,N_2600,N_2598);
or U9333 (N_9333,N_170,N_909);
nand U9334 (N_9334,N_2079,N_3666);
or U9335 (N_9335,N_4672,N_2022);
and U9336 (N_9336,N_3211,N_2426);
and U9337 (N_9337,N_3441,N_4607);
or U9338 (N_9338,N_1102,N_1267);
or U9339 (N_9339,N_1465,N_4790);
nor U9340 (N_9340,N_1631,N_2594);
or U9341 (N_9341,N_1391,N_4603);
nand U9342 (N_9342,N_1664,N_3202);
or U9343 (N_9343,N_4922,N_3429);
nand U9344 (N_9344,N_928,N_3688);
or U9345 (N_9345,N_4798,N_2077);
or U9346 (N_9346,N_1780,N_2011);
nand U9347 (N_9347,N_4527,N_1406);
nor U9348 (N_9348,N_4937,N_3282);
and U9349 (N_9349,N_2003,N_872);
nand U9350 (N_9350,N_3792,N_2585);
nand U9351 (N_9351,N_3564,N_4249);
or U9352 (N_9352,N_750,N_2830);
and U9353 (N_9353,N_4955,N_3887);
and U9354 (N_9354,N_4522,N_2537);
or U9355 (N_9355,N_2896,N_3213);
nor U9356 (N_9356,N_2231,N_4702);
nor U9357 (N_9357,N_290,N_4520);
nand U9358 (N_9358,N_2570,N_2085);
nor U9359 (N_9359,N_4242,N_4745);
nand U9360 (N_9360,N_4770,N_4354);
and U9361 (N_9361,N_559,N_931);
and U9362 (N_9362,N_352,N_3008);
nor U9363 (N_9363,N_3173,N_144);
and U9364 (N_9364,N_788,N_5);
nand U9365 (N_9365,N_4659,N_183);
and U9366 (N_9366,N_3287,N_3594);
nand U9367 (N_9367,N_3793,N_2835);
and U9368 (N_9368,N_739,N_718);
and U9369 (N_9369,N_3924,N_2870);
nor U9370 (N_9370,N_3802,N_1693);
nor U9371 (N_9371,N_2415,N_113);
and U9372 (N_9372,N_857,N_3856);
nor U9373 (N_9373,N_3118,N_817);
or U9374 (N_9374,N_696,N_2253);
nor U9375 (N_9375,N_4607,N_907);
nor U9376 (N_9376,N_2604,N_3026);
or U9377 (N_9377,N_682,N_2825);
or U9378 (N_9378,N_3304,N_1083);
nand U9379 (N_9379,N_283,N_478);
and U9380 (N_9380,N_1005,N_4425);
and U9381 (N_9381,N_2794,N_4970);
or U9382 (N_9382,N_2631,N_2238);
or U9383 (N_9383,N_4125,N_4513);
and U9384 (N_9384,N_2397,N_3061);
or U9385 (N_9385,N_4044,N_1637);
and U9386 (N_9386,N_3597,N_3768);
nand U9387 (N_9387,N_2920,N_3111);
or U9388 (N_9388,N_1238,N_1184);
nor U9389 (N_9389,N_1511,N_834);
nand U9390 (N_9390,N_4170,N_1794);
and U9391 (N_9391,N_4700,N_4154);
nand U9392 (N_9392,N_1587,N_4376);
or U9393 (N_9393,N_2065,N_973);
or U9394 (N_9394,N_2136,N_1224);
or U9395 (N_9395,N_263,N_2259);
or U9396 (N_9396,N_3458,N_3188);
or U9397 (N_9397,N_2814,N_4743);
nor U9398 (N_9398,N_2839,N_2334);
nand U9399 (N_9399,N_2056,N_2058);
nor U9400 (N_9400,N_1385,N_3195);
nand U9401 (N_9401,N_3320,N_2474);
and U9402 (N_9402,N_233,N_670);
nand U9403 (N_9403,N_4418,N_521);
nand U9404 (N_9404,N_733,N_572);
nand U9405 (N_9405,N_2547,N_127);
xnor U9406 (N_9406,N_182,N_644);
nand U9407 (N_9407,N_3412,N_3071);
and U9408 (N_9408,N_2419,N_1562);
nand U9409 (N_9409,N_1890,N_3852);
nand U9410 (N_9410,N_1271,N_1969);
and U9411 (N_9411,N_4102,N_2449);
nor U9412 (N_9412,N_2312,N_3335);
nand U9413 (N_9413,N_4872,N_3398);
nand U9414 (N_9414,N_4867,N_4697);
nand U9415 (N_9415,N_2455,N_1293);
or U9416 (N_9416,N_1042,N_499);
and U9417 (N_9417,N_1763,N_4179);
and U9418 (N_9418,N_1286,N_4706);
nand U9419 (N_9419,N_3018,N_4785);
xnor U9420 (N_9420,N_183,N_355);
nor U9421 (N_9421,N_337,N_2435);
nand U9422 (N_9422,N_1156,N_3869);
and U9423 (N_9423,N_492,N_1157);
xor U9424 (N_9424,N_4936,N_4199);
and U9425 (N_9425,N_3797,N_460);
or U9426 (N_9426,N_757,N_1310);
nand U9427 (N_9427,N_3819,N_64);
nor U9428 (N_9428,N_3330,N_1271);
nand U9429 (N_9429,N_4140,N_4110);
and U9430 (N_9430,N_1017,N_748);
nor U9431 (N_9431,N_548,N_2104);
nor U9432 (N_9432,N_3204,N_2245);
or U9433 (N_9433,N_1685,N_3395);
nor U9434 (N_9434,N_2693,N_3667);
or U9435 (N_9435,N_4600,N_3907);
and U9436 (N_9436,N_3621,N_4277);
and U9437 (N_9437,N_1499,N_4232);
and U9438 (N_9438,N_3352,N_4555);
nor U9439 (N_9439,N_1648,N_1353);
and U9440 (N_9440,N_107,N_1880);
nand U9441 (N_9441,N_1360,N_2012);
or U9442 (N_9442,N_1988,N_601);
or U9443 (N_9443,N_4271,N_1198);
and U9444 (N_9444,N_3893,N_2770);
or U9445 (N_9445,N_4327,N_3427);
nand U9446 (N_9446,N_1719,N_3418);
nor U9447 (N_9447,N_3627,N_1660);
nor U9448 (N_9448,N_2643,N_3289);
or U9449 (N_9449,N_1562,N_1194);
nand U9450 (N_9450,N_4111,N_4708);
nand U9451 (N_9451,N_4652,N_2941);
or U9452 (N_9452,N_3131,N_3563);
nor U9453 (N_9453,N_2608,N_2627);
or U9454 (N_9454,N_2308,N_1845);
nor U9455 (N_9455,N_178,N_1225);
or U9456 (N_9456,N_2735,N_1972);
nand U9457 (N_9457,N_3814,N_4112);
or U9458 (N_9458,N_4493,N_207);
and U9459 (N_9459,N_24,N_2992);
or U9460 (N_9460,N_3126,N_1188);
and U9461 (N_9461,N_3283,N_403);
nand U9462 (N_9462,N_3140,N_365);
nand U9463 (N_9463,N_896,N_4562);
nor U9464 (N_9464,N_3408,N_1445);
and U9465 (N_9465,N_4432,N_3333);
and U9466 (N_9466,N_3971,N_4999);
nor U9467 (N_9467,N_1403,N_15);
and U9468 (N_9468,N_1452,N_467);
nor U9469 (N_9469,N_2568,N_582);
nor U9470 (N_9470,N_1124,N_3151);
or U9471 (N_9471,N_1712,N_1329);
or U9472 (N_9472,N_760,N_2768);
nand U9473 (N_9473,N_1995,N_2154);
nand U9474 (N_9474,N_4087,N_3762);
and U9475 (N_9475,N_2878,N_4488);
nor U9476 (N_9476,N_1031,N_3734);
and U9477 (N_9477,N_1707,N_3010);
nor U9478 (N_9478,N_958,N_4401);
or U9479 (N_9479,N_2702,N_4954);
nand U9480 (N_9480,N_3448,N_3441);
and U9481 (N_9481,N_19,N_4404);
nand U9482 (N_9482,N_3775,N_149);
nand U9483 (N_9483,N_4874,N_3106);
and U9484 (N_9484,N_4405,N_1378);
and U9485 (N_9485,N_704,N_860);
nor U9486 (N_9486,N_1669,N_2307);
and U9487 (N_9487,N_554,N_3117);
and U9488 (N_9488,N_4865,N_738);
nand U9489 (N_9489,N_4199,N_4140);
and U9490 (N_9490,N_3886,N_3557);
nor U9491 (N_9491,N_1572,N_3233);
or U9492 (N_9492,N_3719,N_4141);
nor U9493 (N_9493,N_4531,N_1282);
nor U9494 (N_9494,N_4840,N_4326);
and U9495 (N_9495,N_4319,N_2094);
and U9496 (N_9496,N_4589,N_523);
or U9497 (N_9497,N_2272,N_2433);
nand U9498 (N_9498,N_2966,N_2795);
and U9499 (N_9499,N_419,N_1340);
and U9500 (N_9500,N_785,N_1691);
or U9501 (N_9501,N_3079,N_888);
and U9502 (N_9502,N_663,N_552);
or U9503 (N_9503,N_696,N_196);
xor U9504 (N_9504,N_265,N_1345);
and U9505 (N_9505,N_2974,N_1970);
nand U9506 (N_9506,N_2352,N_1937);
nand U9507 (N_9507,N_4883,N_1250);
nor U9508 (N_9508,N_581,N_4890);
and U9509 (N_9509,N_546,N_1120);
or U9510 (N_9510,N_2710,N_676);
nor U9511 (N_9511,N_3244,N_588);
and U9512 (N_9512,N_4287,N_2795);
nor U9513 (N_9513,N_2278,N_674);
and U9514 (N_9514,N_1898,N_2420);
or U9515 (N_9515,N_3716,N_1671);
nor U9516 (N_9516,N_1321,N_2595);
and U9517 (N_9517,N_4984,N_3967);
or U9518 (N_9518,N_498,N_1534);
nand U9519 (N_9519,N_1817,N_3556);
or U9520 (N_9520,N_4914,N_2790);
nand U9521 (N_9521,N_4575,N_3480);
nand U9522 (N_9522,N_4266,N_2065);
or U9523 (N_9523,N_2801,N_513);
nand U9524 (N_9524,N_1283,N_1150);
or U9525 (N_9525,N_4500,N_4753);
nand U9526 (N_9526,N_476,N_4419);
nand U9527 (N_9527,N_4672,N_994);
xnor U9528 (N_9528,N_2598,N_3015);
nand U9529 (N_9529,N_1888,N_2744);
and U9530 (N_9530,N_1303,N_3630);
nor U9531 (N_9531,N_2856,N_471);
xor U9532 (N_9532,N_758,N_3977);
and U9533 (N_9533,N_1351,N_4480);
or U9534 (N_9534,N_4790,N_1080);
and U9535 (N_9535,N_3966,N_1255);
and U9536 (N_9536,N_3930,N_4331);
or U9537 (N_9537,N_4412,N_4187);
nand U9538 (N_9538,N_732,N_1684);
nor U9539 (N_9539,N_3919,N_1025);
or U9540 (N_9540,N_2373,N_1259);
or U9541 (N_9541,N_1526,N_479);
nand U9542 (N_9542,N_4832,N_1078);
nand U9543 (N_9543,N_2722,N_647);
nand U9544 (N_9544,N_710,N_4204);
or U9545 (N_9545,N_1545,N_2418);
and U9546 (N_9546,N_4036,N_899);
or U9547 (N_9547,N_3920,N_4642);
or U9548 (N_9548,N_4424,N_93);
or U9549 (N_9549,N_467,N_2598);
and U9550 (N_9550,N_2082,N_18);
or U9551 (N_9551,N_2618,N_2656);
and U9552 (N_9552,N_2453,N_4197);
and U9553 (N_9553,N_4632,N_4441);
and U9554 (N_9554,N_4383,N_3177);
nor U9555 (N_9555,N_2314,N_4575);
and U9556 (N_9556,N_1555,N_474);
and U9557 (N_9557,N_1962,N_277);
and U9558 (N_9558,N_1976,N_1344);
or U9559 (N_9559,N_4207,N_3405);
and U9560 (N_9560,N_2454,N_1464);
nor U9561 (N_9561,N_931,N_2252);
nand U9562 (N_9562,N_2716,N_1754);
nor U9563 (N_9563,N_2429,N_3712);
or U9564 (N_9564,N_3979,N_3717);
or U9565 (N_9565,N_1387,N_141);
or U9566 (N_9566,N_375,N_178);
and U9567 (N_9567,N_867,N_398);
xor U9568 (N_9568,N_3362,N_2562);
and U9569 (N_9569,N_10,N_215);
nand U9570 (N_9570,N_3248,N_2176);
nand U9571 (N_9571,N_3632,N_4233);
nor U9572 (N_9572,N_4299,N_1679);
nand U9573 (N_9573,N_2142,N_4196);
or U9574 (N_9574,N_1882,N_900);
or U9575 (N_9575,N_2034,N_1997);
and U9576 (N_9576,N_2414,N_300);
or U9577 (N_9577,N_2843,N_4901);
and U9578 (N_9578,N_4392,N_1803);
or U9579 (N_9579,N_1098,N_1871);
and U9580 (N_9580,N_2448,N_4063);
nor U9581 (N_9581,N_1115,N_3285);
nor U9582 (N_9582,N_1935,N_1762);
and U9583 (N_9583,N_4029,N_2307);
or U9584 (N_9584,N_3615,N_730);
and U9585 (N_9585,N_3338,N_357);
nor U9586 (N_9586,N_3283,N_699);
xnor U9587 (N_9587,N_124,N_3102);
xor U9588 (N_9588,N_530,N_3839);
nand U9589 (N_9589,N_4340,N_243);
or U9590 (N_9590,N_637,N_1516);
nor U9591 (N_9591,N_2038,N_2384);
and U9592 (N_9592,N_4,N_4650);
nand U9593 (N_9593,N_4024,N_750);
and U9594 (N_9594,N_28,N_4714);
nor U9595 (N_9595,N_1765,N_2792);
nor U9596 (N_9596,N_4397,N_1731);
xnor U9597 (N_9597,N_1515,N_4833);
xor U9598 (N_9598,N_2388,N_817);
or U9599 (N_9599,N_2745,N_2956);
nor U9600 (N_9600,N_1579,N_2738);
or U9601 (N_9601,N_4258,N_2009);
nor U9602 (N_9602,N_514,N_4811);
nor U9603 (N_9603,N_1698,N_1000);
nand U9604 (N_9604,N_2055,N_2615);
or U9605 (N_9605,N_1160,N_616);
nand U9606 (N_9606,N_1978,N_4586);
and U9607 (N_9607,N_2173,N_2698);
or U9608 (N_9608,N_1851,N_1317);
or U9609 (N_9609,N_3509,N_2459);
nand U9610 (N_9610,N_3657,N_1591);
and U9611 (N_9611,N_29,N_744);
nand U9612 (N_9612,N_3642,N_1327);
or U9613 (N_9613,N_3771,N_4243);
nand U9614 (N_9614,N_4039,N_982);
nor U9615 (N_9615,N_1278,N_4475);
or U9616 (N_9616,N_582,N_529);
or U9617 (N_9617,N_1739,N_3153);
nand U9618 (N_9618,N_1659,N_4246);
or U9619 (N_9619,N_905,N_4199);
or U9620 (N_9620,N_3029,N_3314);
nor U9621 (N_9621,N_3995,N_1139);
nor U9622 (N_9622,N_4062,N_3547);
nand U9623 (N_9623,N_2737,N_3726);
or U9624 (N_9624,N_4238,N_443);
nand U9625 (N_9625,N_3199,N_1739);
nor U9626 (N_9626,N_1562,N_2212);
nand U9627 (N_9627,N_3801,N_1634);
and U9628 (N_9628,N_4642,N_4026);
nand U9629 (N_9629,N_4577,N_3752);
nand U9630 (N_9630,N_2387,N_812);
and U9631 (N_9631,N_1868,N_214);
and U9632 (N_9632,N_3969,N_160);
or U9633 (N_9633,N_3943,N_2236);
nand U9634 (N_9634,N_3500,N_1855);
or U9635 (N_9635,N_2214,N_1294);
nor U9636 (N_9636,N_3048,N_1163);
nor U9637 (N_9637,N_4652,N_4697);
nor U9638 (N_9638,N_4469,N_4395);
or U9639 (N_9639,N_3311,N_2875);
and U9640 (N_9640,N_724,N_356);
nand U9641 (N_9641,N_1932,N_704);
and U9642 (N_9642,N_2066,N_390);
or U9643 (N_9643,N_1828,N_3478);
nor U9644 (N_9644,N_4128,N_308);
nor U9645 (N_9645,N_3007,N_516);
nor U9646 (N_9646,N_4313,N_1004);
or U9647 (N_9647,N_2636,N_1433);
nand U9648 (N_9648,N_2802,N_4993);
nand U9649 (N_9649,N_878,N_1330);
nor U9650 (N_9650,N_950,N_4905);
nand U9651 (N_9651,N_3434,N_3341);
nor U9652 (N_9652,N_4661,N_3956);
nand U9653 (N_9653,N_168,N_1601);
nor U9654 (N_9654,N_4237,N_4671);
and U9655 (N_9655,N_323,N_3423);
nor U9656 (N_9656,N_369,N_2841);
nand U9657 (N_9657,N_4605,N_872);
or U9658 (N_9658,N_2932,N_1421);
or U9659 (N_9659,N_4767,N_1220);
nand U9660 (N_9660,N_4372,N_1759);
or U9661 (N_9661,N_4886,N_1209);
or U9662 (N_9662,N_452,N_4998);
and U9663 (N_9663,N_4541,N_943);
and U9664 (N_9664,N_82,N_3869);
and U9665 (N_9665,N_3682,N_2816);
nand U9666 (N_9666,N_3190,N_3675);
and U9667 (N_9667,N_4998,N_3151);
nor U9668 (N_9668,N_890,N_2427);
nand U9669 (N_9669,N_532,N_3454);
or U9670 (N_9670,N_1950,N_1220);
nor U9671 (N_9671,N_880,N_761);
nand U9672 (N_9672,N_2019,N_1534);
nor U9673 (N_9673,N_561,N_4857);
or U9674 (N_9674,N_709,N_1946);
nand U9675 (N_9675,N_3150,N_564);
or U9676 (N_9676,N_938,N_4063);
and U9677 (N_9677,N_655,N_4363);
or U9678 (N_9678,N_209,N_4181);
nor U9679 (N_9679,N_1999,N_4708);
nand U9680 (N_9680,N_4730,N_1994);
nor U9681 (N_9681,N_3341,N_4980);
xor U9682 (N_9682,N_4176,N_4968);
nor U9683 (N_9683,N_2105,N_3352);
or U9684 (N_9684,N_370,N_1328);
and U9685 (N_9685,N_3076,N_1805);
and U9686 (N_9686,N_4020,N_2968);
nand U9687 (N_9687,N_481,N_4716);
nor U9688 (N_9688,N_12,N_2756);
nand U9689 (N_9689,N_2504,N_2033);
or U9690 (N_9690,N_1091,N_4366);
and U9691 (N_9691,N_1324,N_3597);
and U9692 (N_9692,N_4007,N_2516);
nand U9693 (N_9693,N_524,N_2004);
nor U9694 (N_9694,N_3128,N_2860);
nand U9695 (N_9695,N_994,N_727);
and U9696 (N_9696,N_4945,N_1498);
and U9697 (N_9697,N_4395,N_762);
or U9698 (N_9698,N_2286,N_3092);
or U9699 (N_9699,N_172,N_1536);
nor U9700 (N_9700,N_357,N_83);
or U9701 (N_9701,N_4073,N_2247);
or U9702 (N_9702,N_1745,N_1403);
or U9703 (N_9703,N_1053,N_2585);
or U9704 (N_9704,N_3043,N_4914);
nand U9705 (N_9705,N_4278,N_1828);
or U9706 (N_9706,N_4808,N_474);
nand U9707 (N_9707,N_4626,N_4083);
nor U9708 (N_9708,N_314,N_1276);
nand U9709 (N_9709,N_268,N_2969);
and U9710 (N_9710,N_4116,N_4010);
nand U9711 (N_9711,N_1316,N_2007);
nand U9712 (N_9712,N_4001,N_2566);
nand U9713 (N_9713,N_448,N_2451);
or U9714 (N_9714,N_1747,N_4485);
nand U9715 (N_9715,N_3247,N_2765);
and U9716 (N_9716,N_1538,N_1124);
nand U9717 (N_9717,N_4621,N_2633);
or U9718 (N_9718,N_134,N_408);
and U9719 (N_9719,N_1948,N_4698);
nor U9720 (N_9720,N_4053,N_749);
nor U9721 (N_9721,N_4397,N_2543);
and U9722 (N_9722,N_4931,N_2830);
and U9723 (N_9723,N_681,N_2600);
and U9724 (N_9724,N_3587,N_2831);
nor U9725 (N_9725,N_2738,N_4682);
or U9726 (N_9726,N_1528,N_528);
and U9727 (N_9727,N_3116,N_2600);
nor U9728 (N_9728,N_4382,N_1128);
nor U9729 (N_9729,N_1960,N_1357);
or U9730 (N_9730,N_4538,N_219);
and U9731 (N_9731,N_3239,N_4900);
and U9732 (N_9732,N_4591,N_60);
nor U9733 (N_9733,N_2878,N_1960);
and U9734 (N_9734,N_4573,N_3323);
nor U9735 (N_9735,N_4584,N_1105);
or U9736 (N_9736,N_923,N_1559);
nor U9737 (N_9737,N_3060,N_3868);
and U9738 (N_9738,N_3075,N_2394);
and U9739 (N_9739,N_2357,N_1493);
nor U9740 (N_9740,N_1673,N_4453);
and U9741 (N_9741,N_1582,N_2578);
nand U9742 (N_9742,N_1272,N_2995);
nor U9743 (N_9743,N_1059,N_4907);
or U9744 (N_9744,N_3344,N_678);
and U9745 (N_9745,N_3200,N_235);
or U9746 (N_9746,N_1146,N_4492);
and U9747 (N_9747,N_2527,N_2364);
nand U9748 (N_9748,N_4893,N_3021);
or U9749 (N_9749,N_2175,N_3570);
nor U9750 (N_9750,N_3967,N_2018);
or U9751 (N_9751,N_2998,N_3465);
or U9752 (N_9752,N_4181,N_2675);
or U9753 (N_9753,N_1408,N_1104);
xnor U9754 (N_9754,N_1846,N_4875);
or U9755 (N_9755,N_2846,N_4678);
or U9756 (N_9756,N_4598,N_3578);
and U9757 (N_9757,N_52,N_1905);
nor U9758 (N_9758,N_2685,N_3824);
nor U9759 (N_9759,N_2313,N_2145);
and U9760 (N_9760,N_4491,N_3500);
and U9761 (N_9761,N_1832,N_1226);
nand U9762 (N_9762,N_1504,N_4491);
nor U9763 (N_9763,N_3574,N_1265);
nand U9764 (N_9764,N_753,N_998);
and U9765 (N_9765,N_3603,N_739);
nand U9766 (N_9766,N_4846,N_1778);
and U9767 (N_9767,N_4093,N_1191);
and U9768 (N_9768,N_1879,N_4566);
and U9769 (N_9769,N_4658,N_685);
and U9770 (N_9770,N_1085,N_4678);
and U9771 (N_9771,N_3231,N_2038);
xnor U9772 (N_9772,N_2362,N_1011);
or U9773 (N_9773,N_4352,N_4017);
nor U9774 (N_9774,N_2643,N_2572);
and U9775 (N_9775,N_3663,N_4725);
nand U9776 (N_9776,N_4486,N_769);
nor U9777 (N_9777,N_348,N_150);
nor U9778 (N_9778,N_3936,N_2456);
or U9779 (N_9779,N_3117,N_3475);
and U9780 (N_9780,N_2722,N_2671);
or U9781 (N_9781,N_631,N_205);
and U9782 (N_9782,N_968,N_2413);
and U9783 (N_9783,N_3275,N_224);
or U9784 (N_9784,N_228,N_997);
nor U9785 (N_9785,N_1472,N_371);
nor U9786 (N_9786,N_4017,N_636);
and U9787 (N_9787,N_4501,N_2565);
or U9788 (N_9788,N_2516,N_3669);
and U9789 (N_9789,N_1211,N_1221);
nand U9790 (N_9790,N_4599,N_3985);
nor U9791 (N_9791,N_2946,N_3386);
nor U9792 (N_9792,N_1813,N_4816);
and U9793 (N_9793,N_4675,N_2823);
nand U9794 (N_9794,N_2666,N_490);
and U9795 (N_9795,N_3749,N_2802);
nand U9796 (N_9796,N_484,N_1561);
and U9797 (N_9797,N_4077,N_4142);
nand U9798 (N_9798,N_3144,N_419);
or U9799 (N_9799,N_452,N_3702);
and U9800 (N_9800,N_3887,N_3935);
nor U9801 (N_9801,N_746,N_3314);
or U9802 (N_9802,N_1063,N_4081);
nor U9803 (N_9803,N_535,N_4565);
and U9804 (N_9804,N_420,N_2027);
or U9805 (N_9805,N_3390,N_2502);
nor U9806 (N_9806,N_3633,N_1521);
or U9807 (N_9807,N_3895,N_3464);
nor U9808 (N_9808,N_2963,N_2488);
or U9809 (N_9809,N_4507,N_1389);
nor U9810 (N_9810,N_4003,N_1588);
nand U9811 (N_9811,N_2891,N_3716);
and U9812 (N_9812,N_3600,N_1995);
nor U9813 (N_9813,N_2633,N_234);
nor U9814 (N_9814,N_3984,N_4622);
nor U9815 (N_9815,N_1756,N_388);
nand U9816 (N_9816,N_1101,N_1462);
or U9817 (N_9817,N_1082,N_901);
or U9818 (N_9818,N_4915,N_3405);
or U9819 (N_9819,N_4464,N_4888);
or U9820 (N_9820,N_595,N_3519);
nand U9821 (N_9821,N_4237,N_1977);
and U9822 (N_9822,N_2014,N_633);
or U9823 (N_9823,N_3017,N_701);
nor U9824 (N_9824,N_1592,N_4738);
nor U9825 (N_9825,N_3143,N_3284);
xor U9826 (N_9826,N_4651,N_1229);
and U9827 (N_9827,N_1700,N_1200);
or U9828 (N_9828,N_185,N_247);
and U9829 (N_9829,N_24,N_1259);
nand U9830 (N_9830,N_113,N_2096);
and U9831 (N_9831,N_3949,N_2189);
and U9832 (N_9832,N_2525,N_1325);
or U9833 (N_9833,N_1685,N_2978);
and U9834 (N_9834,N_2721,N_3627);
nor U9835 (N_9835,N_3008,N_2949);
nor U9836 (N_9836,N_2143,N_530);
and U9837 (N_9837,N_4403,N_1301);
nor U9838 (N_9838,N_4758,N_4457);
or U9839 (N_9839,N_2314,N_3188);
or U9840 (N_9840,N_3825,N_4863);
and U9841 (N_9841,N_612,N_1761);
or U9842 (N_9842,N_4923,N_830);
or U9843 (N_9843,N_4940,N_4444);
and U9844 (N_9844,N_4669,N_1135);
and U9845 (N_9845,N_3300,N_643);
or U9846 (N_9846,N_800,N_79);
or U9847 (N_9847,N_1342,N_1729);
nand U9848 (N_9848,N_2479,N_3774);
nand U9849 (N_9849,N_389,N_882);
nand U9850 (N_9850,N_4400,N_4155);
nand U9851 (N_9851,N_1781,N_2916);
nand U9852 (N_9852,N_4446,N_4863);
and U9853 (N_9853,N_2684,N_4263);
or U9854 (N_9854,N_120,N_2509);
nand U9855 (N_9855,N_4861,N_1996);
nand U9856 (N_9856,N_2513,N_815);
nand U9857 (N_9857,N_4901,N_1863);
nand U9858 (N_9858,N_2687,N_4954);
or U9859 (N_9859,N_4584,N_1816);
nor U9860 (N_9860,N_1208,N_130);
nand U9861 (N_9861,N_351,N_2579);
nand U9862 (N_9862,N_4921,N_4990);
nor U9863 (N_9863,N_1645,N_2907);
or U9864 (N_9864,N_3008,N_4639);
nor U9865 (N_9865,N_831,N_1269);
nand U9866 (N_9866,N_3485,N_1006);
or U9867 (N_9867,N_3852,N_645);
nand U9868 (N_9868,N_1977,N_4242);
nand U9869 (N_9869,N_4373,N_1802);
nand U9870 (N_9870,N_4395,N_4655);
or U9871 (N_9871,N_2354,N_4907);
nand U9872 (N_9872,N_2576,N_4030);
nand U9873 (N_9873,N_1421,N_4261);
or U9874 (N_9874,N_578,N_4115);
nand U9875 (N_9875,N_1079,N_935);
and U9876 (N_9876,N_342,N_3536);
or U9877 (N_9877,N_2618,N_4848);
nor U9878 (N_9878,N_1583,N_3375);
xor U9879 (N_9879,N_1654,N_3464);
or U9880 (N_9880,N_4906,N_823);
and U9881 (N_9881,N_2571,N_1835);
or U9882 (N_9882,N_3595,N_3290);
or U9883 (N_9883,N_2025,N_1013);
and U9884 (N_9884,N_443,N_2484);
xnor U9885 (N_9885,N_2933,N_2043);
and U9886 (N_9886,N_340,N_1704);
nand U9887 (N_9887,N_2876,N_981);
nand U9888 (N_9888,N_699,N_3799);
nor U9889 (N_9889,N_624,N_3966);
nor U9890 (N_9890,N_4045,N_4388);
xnor U9891 (N_9891,N_2685,N_4633);
nor U9892 (N_9892,N_4343,N_1906);
and U9893 (N_9893,N_235,N_246);
nor U9894 (N_9894,N_1009,N_3303);
and U9895 (N_9895,N_3651,N_1370);
or U9896 (N_9896,N_891,N_3969);
nor U9897 (N_9897,N_1936,N_1832);
and U9898 (N_9898,N_4838,N_2649);
and U9899 (N_9899,N_2244,N_3710);
or U9900 (N_9900,N_2829,N_4890);
and U9901 (N_9901,N_1957,N_1963);
nand U9902 (N_9902,N_56,N_3477);
or U9903 (N_9903,N_4411,N_2528);
or U9904 (N_9904,N_393,N_4652);
nor U9905 (N_9905,N_1510,N_1459);
nor U9906 (N_9906,N_4119,N_4463);
and U9907 (N_9907,N_3181,N_1178);
nand U9908 (N_9908,N_3933,N_2060);
xnor U9909 (N_9909,N_511,N_509);
or U9910 (N_9910,N_3151,N_2886);
and U9911 (N_9911,N_936,N_646);
nor U9912 (N_9912,N_3139,N_1117);
nor U9913 (N_9913,N_1173,N_248);
nor U9914 (N_9914,N_4432,N_460);
nor U9915 (N_9915,N_1145,N_4754);
nor U9916 (N_9916,N_1224,N_1482);
or U9917 (N_9917,N_3474,N_4848);
and U9918 (N_9918,N_3433,N_3377);
and U9919 (N_9919,N_3187,N_4381);
nor U9920 (N_9920,N_2919,N_2938);
and U9921 (N_9921,N_2372,N_2200);
nand U9922 (N_9922,N_2534,N_1208);
nor U9923 (N_9923,N_593,N_421);
or U9924 (N_9924,N_4281,N_2514);
or U9925 (N_9925,N_4205,N_4084);
or U9926 (N_9926,N_3606,N_1652);
nand U9927 (N_9927,N_551,N_3961);
and U9928 (N_9928,N_2004,N_4731);
nor U9929 (N_9929,N_4752,N_1913);
or U9930 (N_9930,N_3166,N_11);
nand U9931 (N_9931,N_443,N_2671);
nor U9932 (N_9932,N_4929,N_4353);
nand U9933 (N_9933,N_708,N_4295);
nand U9934 (N_9934,N_1719,N_374);
and U9935 (N_9935,N_3698,N_122);
or U9936 (N_9936,N_3755,N_164);
or U9937 (N_9937,N_304,N_955);
or U9938 (N_9938,N_1114,N_4212);
or U9939 (N_9939,N_4904,N_309);
or U9940 (N_9940,N_553,N_4751);
and U9941 (N_9941,N_1981,N_1797);
nand U9942 (N_9942,N_3476,N_924);
nand U9943 (N_9943,N_4329,N_3253);
and U9944 (N_9944,N_1057,N_2290);
nand U9945 (N_9945,N_4996,N_3071);
nor U9946 (N_9946,N_3108,N_4891);
nor U9947 (N_9947,N_2107,N_4608);
nand U9948 (N_9948,N_716,N_3884);
xnor U9949 (N_9949,N_3655,N_1190);
xor U9950 (N_9950,N_376,N_2640);
and U9951 (N_9951,N_859,N_3131);
nor U9952 (N_9952,N_2926,N_863);
and U9953 (N_9953,N_599,N_4602);
nor U9954 (N_9954,N_2351,N_488);
nor U9955 (N_9955,N_1478,N_802);
xnor U9956 (N_9956,N_3748,N_502);
nor U9957 (N_9957,N_88,N_4960);
or U9958 (N_9958,N_189,N_1471);
or U9959 (N_9959,N_3251,N_740);
or U9960 (N_9960,N_1372,N_694);
nor U9961 (N_9961,N_2671,N_3796);
nand U9962 (N_9962,N_2689,N_1710);
nor U9963 (N_9963,N_4393,N_510);
nor U9964 (N_9964,N_970,N_1801);
nor U9965 (N_9965,N_4081,N_1784);
nand U9966 (N_9966,N_4653,N_4523);
xnor U9967 (N_9967,N_3181,N_3327);
xor U9968 (N_9968,N_531,N_2128);
and U9969 (N_9969,N_4805,N_722);
and U9970 (N_9970,N_356,N_3210);
nor U9971 (N_9971,N_424,N_1215);
nand U9972 (N_9972,N_1196,N_443);
nor U9973 (N_9973,N_4395,N_4095);
or U9974 (N_9974,N_1983,N_3850);
nand U9975 (N_9975,N_1015,N_2997);
and U9976 (N_9976,N_1633,N_2814);
and U9977 (N_9977,N_4779,N_1808);
nand U9978 (N_9978,N_3091,N_264);
or U9979 (N_9979,N_4517,N_4330);
or U9980 (N_9980,N_513,N_1232);
and U9981 (N_9981,N_4690,N_28);
nand U9982 (N_9982,N_559,N_1826);
and U9983 (N_9983,N_4933,N_4552);
nand U9984 (N_9984,N_3991,N_476);
or U9985 (N_9985,N_3166,N_4675);
and U9986 (N_9986,N_254,N_2121);
and U9987 (N_9987,N_1898,N_2019);
or U9988 (N_9988,N_3151,N_4983);
and U9989 (N_9989,N_3733,N_309);
nand U9990 (N_9990,N_1067,N_3795);
nor U9991 (N_9991,N_4930,N_1324);
nor U9992 (N_9992,N_4209,N_3935);
or U9993 (N_9993,N_4341,N_2303);
nor U9994 (N_9994,N_3668,N_4279);
nand U9995 (N_9995,N_799,N_4790);
nand U9996 (N_9996,N_4062,N_4669);
and U9997 (N_9997,N_2702,N_1349);
nand U9998 (N_9998,N_4276,N_2720);
or U9999 (N_9999,N_3525,N_3350);
nand U10000 (N_10000,N_9906,N_5401);
or U10001 (N_10001,N_9622,N_5736);
nor U10002 (N_10002,N_9818,N_9964);
and U10003 (N_10003,N_8354,N_8270);
or U10004 (N_10004,N_9394,N_7492);
or U10005 (N_10005,N_6759,N_9276);
nand U10006 (N_10006,N_6315,N_8802);
and U10007 (N_10007,N_6629,N_7062);
xor U10008 (N_10008,N_7385,N_9686);
or U10009 (N_10009,N_9192,N_5290);
or U10010 (N_10010,N_5999,N_5744);
and U10011 (N_10011,N_5682,N_9855);
and U10012 (N_10012,N_8001,N_6439);
and U10013 (N_10013,N_5314,N_6991);
or U10014 (N_10014,N_5877,N_9318);
nand U10015 (N_10015,N_7513,N_6911);
nor U10016 (N_10016,N_6066,N_5034);
and U10017 (N_10017,N_5924,N_9474);
nor U10018 (N_10018,N_9213,N_8220);
nand U10019 (N_10019,N_6146,N_5408);
nor U10020 (N_10020,N_6669,N_6976);
nor U10021 (N_10021,N_6494,N_5753);
nor U10022 (N_10022,N_6938,N_7920);
nand U10023 (N_10023,N_6215,N_7774);
and U10024 (N_10024,N_7945,N_9031);
or U10025 (N_10025,N_9901,N_9999);
nand U10026 (N_10026,N_5449,N_9458);
or U10027 (N_10027,N_6865,N_5621);
or U10028 (N_10028,N_6607,N_7688);
nand U10029 (N_10029,N_8797,N_9446);
or U10030 (N_10030,N_8574,N_8915);
and U10031 (N_10031,N_9732,N_5973);
or U10032 (N_10032,N_7532,N_7816);
or U10033 (N_10033,N_7488,N_6412);
nor U10034 (N_10034,N_9698,N_8312);
or U10035 (N_10035,N_6294,N_7763);
nor U10036 (N_10036,N_7271,N_8558);
nor U10037 (N_10037,N_5029,N_6372);
nor U10038 (N_10038,N_6906,N_6462);
nand U10039 (N_10039,N_8218,N_5939);
and U10040 (N_10040,N_9969,N_8686);
nor U10041 (N_10041,N_9072,N_8066);
and U10042 (N_10042,N_8019,N_9646);
and U10043 (N_10043,N_5895,N_5176);
nor U10044 (N_10044,N_6077,N_5522);
nand U10045 (N_10045,N_7058,N_5321);
nand U10046 (N_10046,N_9106,N_5425);
nand U10047 (N_10047,N_6919,N_8688);
or U10048 (N_10048,N_5198,N_7667);
nand U10049 (N_10049,N_7915,N_7470);
or U10050 (N_10050,N_7857,N_9239);
or U10051 (N_10051,N_6529,N_5389);
nand U10052 (N_10052,N_9699,N_6133);
and U10053 (N_10053,N_6762,N_5247);
or U10054 (N_10054,N_9330,N_9028);
or U10055 (N_10055,N_9862,N_8930);
and U10056 (N_10056,N_7267,N_9603);
and U10057 (N_10057,N_9570,N_7429);
and U10058 (N_10058,N_5043,N_8828);
nor U10059 (N_10059,N_5160,N_7115);
or U10060 (N_10060,N_8496,N_7328);
or U10061 (N_10061,N_6861,N_6791);
or U10062 (N_10062,N_7051,N_7472);
or U10063 (N_10063,N_5732,N_6994);
nand U10064 (N_10064,N_7600,N_6450);
and U10065 (N_10065,N_6880,N_5243);
nand U10066 (N_10066,N_9724,N_9558);
or U10067 (N_10067,N_5880,N_7041);
and U10068 (N_10068,N_5585,N_6005);
nand U10069 (N_10069,N_9094,N_9015);
nand U10070 (N_10070,N_9151,N_5801);
nand U10071 (N_10071,N_7085,N_8091);
and U10072 (N_10072,N_8861,N_8808);
nand U10073 (N_10073,N_9842,N_9697);
xor U10074 (N_10074,N_6178,N_6986);
or U10075 (N_10075,N_8081,N_9451);
or U10076 (N_10076,N_6828,N_9419);
or U10077 (N_10077,N_6770,N_7476);
nor U10078 (N_10078,N_5493,N_9748);
or U10079 (N_10079,N_6645,N_8581);
and U10080 (N_10080,N_5051,N_7593);
or U10081 (N_10081,N_5267,N_8801);
nand U10082 (N_10082,N_7338,N_9073);
nor U10083 (N_10083,N_5604,N_6139);
or U10084 (N_10084,N_9742,N_6259);
nor U10085 (N_10085,N_9866,N_7790);
and U10086 (N_10086,N_5322,N_9963);
or U10087 (N_10087,N_8219,N_8903);
nor U10088 (N_10088,N_7639,N_7680);
nand U10089 (N_10089,N_9684,N_8414);
nor U10090 (N_10090,N_5009,N_6422);
xor U10091 (N_10091,N_9762,N_5205);
or U10092 (N_10092,N_9362,N_9783);
nand U10093 (N_10093,N_7377,N_6147);
nor U10094 (N_10094,N_8022,N_8487);
and U10095 (N_10095,N_5110,N_5157);
or U10096 (N_10096,N_6163,N_6881);
and U10097 (N_10097,N_8046,N_9281);
and U10098 (N_10098,N_5560,N_6324);
and U10099 (N_10099,N_8604,N_8642);
or U10100 (N_10100,N_6948,N_5388);
or U10101 (N_10101,N_9562,N_5628);
nor U10102 (N_10102,N_5847,N_5074);
nand U10103 (N_10103,N_7992,N_7000);
nand U10104 (N_10104,N_5437,N_9214);
or U10105 (N_10105,N_9477,N_5533);
nor U10106 (N_10106,N_6845,N_5250);
or U10107 (N_10107,N_7113,N_6067);
xor U10108 (N_10108,N_8386,N_7164);
nor U10109 (N_10109,N_9756,N_7989);
or U10110 (N_10110,N_8174,N_7918);
nor U10111 (N_10111,N_7794,N_7868);
and U10112 (N_10112,N_6300,N_7055);
or U10113 (N_10113,N_7906,N_7908);
xor U10114 (N_10114,N_8234,N_9011);
nor U10115 (N_10115,N_5768,N_9879);
or U10116 (N_10116,N_7169,N_6411);
nor U10117 (N_10117,N_5954,N_8902);
nand U10118 (N_10118,N_9676,N_9173);
nand U10119 (N_10119,N_5120,N_9545);
and U10120 (N_10120,N_5173,N_7626);
nor U10121 (N_10121,N_5625,N_7151);
or U10122 (N_10122,N_7033,N_9508);
xor U10123 (N_10123,N_6103,N_7694);
and U10124 (N_10124,N_5891,N_6522);
nand U10125 (N_10125,N_5126,N_9821);
or U10126 (N_10126,N_6849,N_8334);
or U10127 (N_10127,N_6024,N_7421);
nand U10128 (N_10128,N_7026,N_9655);
nor U10129 (N_10129,N_7150,N_5724);
nand U10130 (N_10130,N_6662,N_9802);
nand U10131 (N_10131,N_5101,N_8189);
or U10132 (N_10132,N_9645,N_9060);
or U10133 (N_10133,N_7437,N_7562);
nand U10134 (N_10134,N_8914,N_6457);
or U10135 (N_10135,N_5980,N_8578);
nand U10136 (N_10136,N_6748,N_9472);
or U10137 (N_10137,N_8768,N_9129);
nand U10138 (N_10138,N_8564,N_9255);
or U10139 (N_10139,N_5300,N_9457);
and U10140 (N_10140,N_9062,N_9672);
nor U10141 (N_10141,N_9246,N_7685);
nor U10142 (N_10142,N_7661,N_5192);
or U10143 (N_10143,N_6839,N_9071);
and U10144 (N_10144,N_5244,N_6942);
nor U10145 (N_10145,N_8593,N_6757);
nand U10146 (N_10146,N_7324,N_5215);
and U10147 (N_10147,N_7962,N_7783);
nand U10148 (N_10148,N_5197,N_7076);
or U10149 (N_10149,N_8853,N_9585);
or U10150 (N_10150,N_8908,N_7690);
or U10151 (N_10151,N_7795,N_5874);
nand U10152 (N_10152,N_9825,N_7960);
or U10153 (N_10153,N_6953,N_7642);
and U10154 (N_10154,N_8211,N_8423);
or U10155 (N_10155,N_8199,N_9306);
or U10156 (N_10156,N_6696,N_9565);
xor U10157 (N_10157,N_6446,N_5918);
or U10158 (N_10158,N_8568,N_9487);
and U10159 (N_10159,N_8494,N_9867);
and U10160 (N_10160,N_8783,N_6175);
and U10161 (N_10161,N_9381,N_7280);
nand U10162 (N_10162,N_6594,N_9393);
nor U10163 (N_10163,N_5607,N_8567);
nand U10164 (N_10164,N_8116,N_5210);
or U10165 (N_10165,N_5920,N_8843);
or U10166 (N_10166,N_8000,N_7102);
nand U10167 (N_10167,N_7522,N_6417);
nor U10168 (N_10168,N_7198,N_6341);
and U10169 (N_10169,N_7994,N_7602);
nand U10170 (N_10170,N_8086,N_8790);
or U10171 (N_10171,N_8398,N_5399);
and U10172 (N_10172,N_7482,N_8160);
nand U10173 (N_10173,N_8241,N_5123);
and U10174 (N_10174,N_9627,N_6838);
and U10175 (N_10175,N_8878,N_6719);
nor U10176 (N_10176,N_6779,N_9261);
nor U10177 (N_10177,N_6473,N_7106);
or U10178 (N_10178,N_9510,N_8426);
or U10179 (N_10179,N_6290,N_9341);
nand U10180 (N_10180,N_9061,N_5330);
nand U10181 (N_10181,N_7349,N_5155);
or U10182 (N_10182,N_6304,N_6380);
nand U10183 (N_10183,N_5571,N_6519);
and U10184 (N_10184,N_9104,N_8480);
nand U10185 (N_10185,N_7497,N_9186);
nor U10186 (N_10186,N_6384,N_6079);
xnor U10187 (N_10187,N_6499,N_9916);
nor U10188 (N_10188,N_9909,N_8532);
nand U10189 (N_10189,N_6279,N_9338);
or U10190 (N_10190,N_6898,N_8984);
or U10191 (N_10191,N_7676,N_6233);
nor U10192 (N_10192,N_7656,N_8089);
nor U10193 (N_10193,N_6443,N_9848);
and U10194 (N_10194,N_6071,N_7067);
and U10195 (N_10195,N_5605,N_6227);
and U10196 (N_10196,N_9004,N_9943);
nor U10197 (N_10197,N_5953,N_6007);
nand U10198 (N_10198,N_5730,N_5985);
nand U10199 (N_10199,N_8483,N_5667);
and U10200 (N_10200,N_6463,N_8047);
nor U10201 (N_10201,N_5125,N_6799);
nand U10202 (N_10202,N_5767,N_6878);
xnor U10203 (N_10203,N_7884,N_9179);
or U10204 (N_10204,N_8159,N_9251);
or U10205 (N_10205,N_6542,N_6467);
and U10206 (N_10206,N_6735,N_5906);
and U10207 (N_10207,N_9103,N_9122);
or U10208 (N_10208,N_6366,N_6676);
nand U10209 (N_10209,N_9088,N_5282);
or U10210 (N_10210,N_5579,N_7941);
nand U10211 (N_10211,N_6404,N_5093);
nand U10212 (N_10212,N_6927,N_7397);
nor U10213 (N_10213,N_5111,N_7448);
nor U10214 (N_10214,N_5837,N_9337);
and U10215 (N_10215,N_9860,N_7954);
xnor U10216 (N_10216,N_8320,N_9165);
and U10217 (N_10217,N_5228,N_9953);
or U10218 (N_10218,N_7742,N_8084);
nand U10219 (N_10219,N_9735,N_7930);
nor U10220 (N_10220,N_9668,N_5103);
nand U10221 (N_10221,N_8064,N_5580);
or U10222 (N_10222,N_7615,N_7436);
nor U10223 (N_10223,N_8836,N_7108);
nand U10224 (N_10224,N_5776,N_6954);
nand U10225 (N_10225,N_8834,N_5639);
and U10226 (N_10226,N_9206,N_6670);
nand U10227 (N_10227,N_8944,N_5256);
nor U10228 (N_10228,N_7321,N_8978);
nand U10229 (N_10229,N_5075,N_7802);
nor U10230 (N_10230,N_6243,N_7266);
nor U10231 (N_10231,N_6508,N_5731);
and U10232 (N_10232,N_8599,N_8013);
or U10233 (N_10233,N_8940,N_9811);
and U10234 (N_10234,N_5128,N_7809);
and U10235 (N_10235,N_7381,N_6060);
and U10236 (N_10236,N_5398,N_9237);
and U10237 (N_10237,N_9870,N_9934);
xor U10238 (N_10238,N_6479,N_6338);
or U10239 (N_10239,N_7326,N_9852);
and U10240 (N_10240,N_8052,N_5411);
nor U10241 (N_10241,N_6438,N_5692);
and U10242 (N_10242,N_9947,N_9736);
nand U10243 (N_10243,N_9121,N_7773);
and U10244 (N_10244,N_9583,N_8246);
nand U10245 (N_10245,N_7242,N_7314);
or U10246 (N_10246,N_7786,N_7713);
nor U10247 (N_10247,N_8233,N_6964);
and U10248 (N_10248,N_9659,N_6336);
and U10249 (N_10249,N_5104,N_6397);
nand U10250 (N_10250,N_7308,N_9409);
nand U10251 (N_10251,N_9701,N_5709);
nand U10252 (N_10252,N_6726,N_6245);
nand U10253 (N_10253,N_5270,N_8315);
and U10254 (N_10254,N_9951,N_8909);
and U10255 (N_10255,N_6042,N_5905);
xnor U10256 (N_10256,N_5316,N_9141);
and U10257 (N_10257,N_5631,N_7705);
nor U10258 (N_10258,N_9405,N_5262);
or U10259 (N_10259,N_7898,N_6254);
nand U10260 (N_10260,N_9689,N_5440);
xnor U10261 (N_10261,N_6855,N_9635);
nor U10262 (N_10262,N_9722,N_5152);
nand U10263 (N_10263,N_5718,N_7717);
and U10264 (N_10264,N_6317,N_5934);
nand U10265 (N_10265,N_7817,N_9492);
or U10266 (N_10266,N_5911,N_5167);
nor U10267 (N_10267,N_6608,N_6430);
nor U10268 (N_10268,N_8666,N_9392);
nand U10269 (N_10269,N_5531,N_6612);
and U10270 (N_10270,N_9054,N_7651);
or U10271 (N_10271,N_9924,N_9354);
and U10272 (N_10272,N_7233,N_6753);
and U10273 (N_10273,N_9021,N_9481);
or U10274 (N_10274,N_9534,N_6741);
nor U10275 (N_10275,N_6742,N_5028);
nand U10276 (N_10276,N_5457,N_6699);
or U10277 (N_10277,N_5748,N_5416);
nand U10278 (N_10278,N_7515,N_8586);
and U10279 (N_10279,N_5410,N_8101);
and U10280 (N_10280,N_7226,N_6088);
nor U10281 (N_10281,N_5749,N_7673);
nor U10282 (N_10282,N_8209,N_8530);
or U10283 (N_10283,N_9417,N_5964);
and U10284 (N_10284,N_5626,N_7101);
and U10285 (N_10285,N_5808,N_5142);
and U10286 (N_10286,N_9703,N_7380);
and U10287 (N_10287,N_8849,N_6378);
and U10288 (N_10288,N_9796,N_7252);
or U10289 (N_10289,N_5651,N_6917);
or U10290 (N_10290,N_6221,N_9713);
nor U10291 (N_10291,N_5060,N_6248);
nand U10292 (N_10292,N_8736,N_8042);
and U10293 (N_10293,N_6729,N_9435);
nor U10294 (N_10294,N_8297,N_5986);
and U10295 (N_10295,N_6774,N_7619);
or U10296 (N_10296,N_8695,N_5670);
nor U10297 (N_10297,N_7311,N_5283);
and U10298 (N_10298,N_9172,N_5432);
nand U10299 (N_10299,N_7096,N_9024);
or U10300 (N_10300,N_8791,N_7531);
and U10301 (N_10301,N_5082,N_5599);
xor U10302 (N_10302,N_8602,N_9163);
nand U10303 (N_10303,N_7956,N_9928);
nand U10304 (N_10304,N_5171,N_5785);
or U10305 (N_10305,N_9184,N_9984);
or U10306 (N_10306,N_6034,N_6541);
nor U10307 (N_10307,N_7319,N_9897);
nor U10308 (N_10308,N_5168,N_6203);
and U10309 (N_10309,N_6143,N_7373);
nand U10310 (N_10310,N_8493,N_8507);
nand U10311 (N_10311,N_5042,N_8479);
nor U10312 (N_10312,N_6061,N_9826);
or U10313 (N_10313,N_9930,N_7216);
and U10314 (N_10314,N_8088,N_8007);
nand U10315 (N_10315,N_9720,N_6135);
nor U10316 (N_10316,N_5400,N_8138);
and U10317 (N_10317,N_9158,N_9939);
and U10318 (N_10318,N_8239,N_9356);
or U10319 (N_10319,N_5269,N_5616);
and U10320 (N_10320,N_7479,N_9611);
nand U10321 (N_10321,N_8035,N_8287);
nor U10322 (N_10322,N_9065,N_9706);
nor U10323 (N_10323,N_6613,N_6540);
and U10324 (N_10324,N_8440,N_9333);
nand U10325 (N_10325,N_8855,N_5045);
and U10326 (N_10326,N_7306,N_7057);
or U10327 (N_10327,N_9990,N_5258);
or U10328 (N_10328,N_8387,N_7674);
and U10329 (N_10329,N_8690,N_7894);
xnor U10330 (N_10330,N_6514,N_9447);
nand U10331 (N_10331,N_5273,N_6068);
nand U10332 (N_10332,N_7175,N_5078);
and U10333 (N_10333,N_9480,N_8729);
nor U10334 (N_10334,N_6533,N_8971);
or U10335 (N_10335,N_7391,N_6744);
and U10336 (N_10336,N_7166,N_5841);
nand U10337 (N_10337,N_9966,N_9566);
or U10338 (N_10338,N_9167,N_8309);
and U10339 (N_10339,N_8215,N_9473);
and U10340 (N_10340,N_5040,N_5097);
and U10341 (N_10341,N_5673,N_5129);
and U10342 (N_10342,N_6251,N_9751);
and U10343 (N_10343,N_7978,N_8513);
and U10344 (N_10344,N_5712,N_6513);
nand U10345 (N_10345,N_9584,N_9958);
xor U10346 (N_10346,N_9295,N_7430);
or U10347 (N_10347,N_9280,N_5955);
or U10348 (N_10348,N_5342,N_7103);
xor U10349 (N_10349,N_9055,N_6225);
nor U10350 (N_10350,N_7720,N_5348);
nor U10351 (N_10351,N_5429,N_5644);
nor U10352 (N_10352,N_9576,N_8226);
or U10353 (N_10353,N_7741,N_5726);
or U10354 (N_10354,N_8640,N_5116);
nand U10355 (N_10355,N_6381,N_6206);
nor U10356 (N_10356,N_8165,N_9787);
and U10357 (N_10357,N_9828,N_7521);
and U10358 (N_10358,N_7776,N_8896);
and U10359 (N_10359,N_8306,N_9497);
and U10360 (N_10360,N_6761,N_5902);
or U10361 (N_10361,N_6382,N_9387);
nor U10362 (N_10362,N_5313,N_8812);
and U10363 (N_10363,N_9675,N_8924);
or U10364 (N_10364,N_5794,N_9131);
nand U10365 (N_10365,N_5061,N_7177);
and U10366 (N_10366,N_8929,N_9965);
or U10367 (N_10367,N_9652,N_7820);
nor U10368 (N_10368,N_5004,N_8938);
or U10369 (N_10369,N_9944,N_7703);
nor U10370 (N_10370,N_5144,N_6451);
nor U10371 (N_10371,N_8054,N_9115);
nand U10372 (N_10372,N_7432,N_8117);
nand U10373 (N_10373,N_7872,N_6686);
nand U10374 (N_10374,N_6489,N_9669);
xnor U10375 (N_10375,N_5175,N_9514);
nor U10376 (N_10376,N_5222,N_9283);
nor U10377 (N_10377,N_7416,N_7581);
and U10378 (N_10378,N_9962,N_6781);
nand U10379 (N_10379,N_8845,N_8910);
and U10380 (N_10380,N_9768,N_6349);
nand U10381 (N_10381,N_9066,N_5583);
or U10382 (N_10382,N_7109,N_6918);
or U10383 (N_10383,N_8850,N_6958);
and U10384 (N_10384,N_5907,N_6485);
nand U10385 (N_10385,N_5271,N_6063);
or U10386 (N_10386,N_7065,N_6978);
nor U10387 (N_10387,N_7854,N_8254);
nor U10388 (N_10388,N_8527,N_6287);
nand U10389 (N_10389,N_9486,N_8027);
nand U10390 (N_10390,N_7384,N_9034);
nor U10391 (N_10391,N_6692,N_5005);
and U10392 (N_10392,N_7539,N_5892);
nand U10393 (N_10393,N_8373,N_5434);
or U10394 (N_10394,N_6016,N_7253);
or U10395 (N_10395,N_9279,N_9342);
nor U10396 (N_10396,N_7003,N_7236);
nor U10397 (N_10397,N_5665,N_9026);
nand U10398 (N_10398,N_7912,N_5421);
and U10399 (N_10399,N_7625,N_9705);
nand U10400 (N_10400,N_7212,N_7796);
nor U10401 (N_10401,N_5239,N_8073);
or U10402 (N_10402,N_5134,N_6162);
and U10403 (N_10403,N_7826,N_9196);
nand U10404 (N_10404,N_9006,N_6140);
and U10405 (N_10405,N_7707,N_6172);
nand U10406 (N_10406,N_8016,N_7935);
and U10407 (N_10407,N_5046,N_9216);
nor U10408 (N_10408,N_7823,N_5196);
and U10409 (N_10409,N_9621,N_8988);
nor U10410 (N_10410,N_6159,N_9022);
nor U10411 (N_10411,N_9120,N_7158);
and U10412 (N_10412,N_8360,N_6655);
or U10413 (N_10413,N_5600,N_9444);
xor U10414 (N_10414,N_5693,N_6894);
and U10415 (N_10415,N_8789,N_7045);
and U10416 (N_10416,N_5526,N_9126);
and U10417 (N_10417,N_6588,N_8539);
nor U10418 (N_10418,N_6641,N_6258);
nand U10419 (N_10419,N_8363,N_8181);
or U10420 (N_10420,N_6039,N_8272);
nand U10421 (N_10421,N_6501,N_9555);
nand U10422 (N_10422,N_9027,N_5280);
xor U10423 (N_10423,N_8974,N_5535);
nor U10424 (N_10424,N_6926,N_8382);
or U10425 (N_10425,N_8708,N_7985);
nor U10426 (N_10426,N_7803,N_6712);
and U10427 (N_10427,N_9604,N_7740);
or U10428 (N_10428,N_8153,N_6385);
nand U10429 (N_10429,N_9128,N_6623);
nand U10430 (N_10430,N_6435,N_6905);
and U10431 (N_10431,N_7426,N_9553);
or U10432 (N_10432,N_6511,N_6065);
nand U10433 (N_10433,N_8502,N_8105);
or U10434 (N_10434,N_6076,N_6295);
and U10435 (N_10435,N_8252,N_7133);
nor U10436 (N_10436,N_6424,N_9225);
nor U10437 (N_10437,N_6325,N_5113);
and U10438 (N_10438,N_7679,N_8684);
nor U10439 (N_10439,N_8609,N_7142);
nand U10440 (N_10440,N_6937,N_7555);
and U10441 (N_10441,N_7630,N_5520);
nand U10442 (N_10442,N_8776,N_5377);
and U10443 (N_10443,N_5848,N_6142);
or U10444 (N_10444,N_8848,N_5549);
and U10445 (N_10445,N_5541,N_6493);
nor U10446 (N_10446,N_9302,N_5771);
nand U10447 (N_10447,N_5236,N_5011);
nor U10448 (N_10448,N_5648,N_6057);
nor U10449 (N_10449,N_9308,N_6805);
nor U10450 (N_10450,N_8351,N_5761);
xnor U10451 (N_10451,N_8628,N_8847);
or U10452 (N_10452,N_5336,N_5772);
nand U10453 (N_10453,N_9479,N_9526);
and U10454 (N_10454,N_8190,N_9992);
nor U10455 (N_10455,N_9933,N_8777);
and U10456 (N_10456,N_9873,N_8550);
or U10457 (N_10457,N_6086,N_7913);
and U10458 (N_10458,N_8150,N_7905);
nor U10459 (N_10459,N_8919,N_5624);
or U10460 (N_10460,N_8113,N_6817);
nand U10461 (N_10461,N_5340,N_5494);
and U10462 (N_10462,N_5386,N_9695);
and U10463 (N_10463,N_9851,N_6503);
or U10464 (N_10464,N_7583,N_7578);
nor U10465 (N_10465,N_8420,N_7862);
nand U10466 (N_10466,N_9009,N_6337);
nand U10467 (N_10467,N_8969,N_5983);
nor U10468 (N_10468,N_8650,N_7764);
nor U10469 (N_10469,N_9369,N_6752);
xor U10470 (N_10470,N_5627,N_9436);
nand U10471 (N_10471,N_9426,N_5255);
nor U10472 (N_10472,N_7654,N_5289);
nand U10473 (N_10473,N_8024,N_5309);
and U10474 (N_10474,N_7502,N_9579);
or U10475 (N_10475,N_8279,N_7163);
nor U10476 (N_10476,N_7700,N_8547);
nand U10477 (N_10477,N_6822,N_9876);
or U10478 (N_10478,N_9687,N_9997);
and U10479 (N_10479,N_6740,N_5504);
xnor U10480 (N_10480,N_8157,N_5414);
nor U10481 (N_10481,N_6399,N_7087);
and U10482 (N_10482,N_7274,N_8689);
nand U10483 (N_10483,N_5067,N_8566);
nor U10484 (N_10484,N_9157,N_9657);
or U10485 (N_10485,N_6318,N_5527);
nor U10486 (N_10486,N_7964,N_5559);
or U10487 (N_10487,N_6923,N_7459);
nand U10488 (N_10488,N_8478,N_5395);
nor U10489 (N_10489,N_7971,N_6156);
and U10490 (N_10490,N_5048,N_9390);
or U10491 (N_10491,N_9693,N_9463);
and U10492 (N_10492,N_8166,N_7801);
and U10493 (N_10493,N_6532,N_9005);
nor U10494 (N_10494,N_6483,N_6054);
or U10495 (N_10495,N_7383,N_8362);
nor U10496 (N_10496,N_5402,N_9312);
nand U10497 (N_10497,N_5789,N_9532);
nor U10498 (N_10498,N_5591,N_8374);
and U10499 (N_10499,N_7849,N_9607);
nor U10500 (N_10500,N_6628,N_7440);
and U10501 (N_10501,N_6598,N_9140);
or U10502 (N_10502,N_9113,N_7950);
nor U10503 (N_10503,N_7839,N_6475);
or U10504 (N_10504,N_5720,N_7732);
or U10505 (N_10505,N_5420,N_5332);
and U10506 (N_10506,N_9240,N_5413);
nand U10507 (N_10507,N_7039,N_5385);
or U10508 (N_10508,N_9344,N_6889);
nor U10509 (N_10509,N_9183,N_8963);
or U10510 (N_10510,N_9755,N_7767);
nor U10511 (N_10511,N_5084,N_5752);
and U10512 (N_10512,N_8589,N_7881);
or U10513 (N_10513,N_9226,N_6272);
nor U10514 (N_10514,N_7154,N_9968);
nor U10515 (N_10515,N_7167,N_7998);
nand U10516 (N_10516,N_8734,N_5746);
nand U10517 (N_10517,N_6468,N_7004);
and U10518 (N_10518,N_6092,N_9494);
and U10519 (N_10519,N_7406,N_5092);
or U10520 (N_10520,N_5513,N_9111);
nand U10521 (N_10521,N_7535,N_8034);
nand U10522 (N_10522,N_5643,N_7494);
nor U10523 (N_10523,N_5925,N_6646);
nor U10524 (N_10524,N_6796,N_5131);
nor U10525 (N_10525,N_7305,N_7709);
and U10526 (N_10526,N_7877,N_5929);
and U10527 (N_10527,N_6314,N_9247);
and U10528 (N_10528,N_8546,N_8477);
and U10529 (N_10529,N_7238,N_8787);
nor U10530 (N_10530,N_8009,N_7018);
xnor U10531 (N_10531,N_7341,N_7910);
nor U10532 (N_10532,N_7892,N_8085);
nor U10533 (N_10533,N_8506,N_8225);
or U10534 (N_10534,N_6126,N_8470);
and U10535 (N_10535,N_9895,N_7100);
nor U10536 (N_10536,N_5186,N_5130);
and U10537 (N_10537,N_9665,N_8661);
or U10538 (N_10538,N_7159,N_6996);
or U10539 (N_10539,N_9413,N_6981);
nor U10540 (N_10540,N_7901,N_5371);
nor U10541 (N_10541,N_9039,N_8879);
or U10542 (N_10542,N_9259,N_6802);
nor U10543 (N_10543,N_6939,N_8949);
nand U10544 (N_10544,N_7889,N_5355);
or U10545 (N_10545,N_6844,N_7805);
or U10546 (N_10546,N_9277,N_8749);
or U10547 (N_10547,N_9149,N_9937);
and U10548 (N_10548,N_7135,N_9979);
and U10549 (N_10549,N_5486,N_6804);
nor U10550 (N_10550,N_6704,N_8617);
nand U10551 (N_10551,N_8605,N_7541);
or U10552 (N_10552,N_5066,N_9452);
or U10553 (N_10553,N_5710,N_6566);
and U10554 (N_10554,N_8028,N_7608);
nand U10555 (N_10555,N_8031,N_9294);
and U10556 (N_10556,N_5164,N_8488);
or U10557 (N_10557,N_8560,N_9644);
nor U10558 (N_10558,N_9483,N_7678);
and U10559 (N_10559,N_6104,N_6323);
and U10560 (N_10560,N_5868,N_5584);
nand U10561 (N_10561,N_6736,N_7197);
nand U10562 (N_10562,N_8983,N_5502);
and U10563 (N_10563,N_7368,N_8316);
nand U10564 (N_10564,N_9936,N_6659);
or U10565 (N_10565,N_5124,N_5013);
nand U10566 (N_10566,N_9769,N_6618);
nand U10567 (N_10567,N_8645,N_6136);
or U10568 (N_10568,N_7850,N_6261);
and U10569 (N_10569,N_8169,N_5363);
xor U10570 (N_10570,N_6552,N_7746);
nor U10571 (N_10571,N_9696,N_9445);
or U10572 (N_10572,N_8203,N_7457);
nor U10573 (N_10573,N_6120,N_9778);
or U10574 (N_10574,N_6702,N_9109);
and U10575 (N_10575,N_7592,N_7507);
and U10576 (N_10576,N_6959,N_7194);
nand U10577 (N_10577,N_7529,N_8486);
or U10578 (N_10578,N_5814,N_7708);
nor U10579 (N_10579,N_8207,N_5885);
or U10580 (N_10580,N_9135,N_9591);
and U10581 (N_10581,N_9462,N_5334);
nand U10582 (N_10582,N_7543,N_5207);
and U10583 (N_10583,N_7070,N_5650);
and U10584 (N_10584,N_9014,N_8145);
nor U10585 (N_10585,N_6112,N_7921);
xor U10586 (N_10586,N_8582,N_6041);
and U10587 (N_10587,N_5966,N_8410);
and U10588 (N_10588,N_7360,N_9367);
and U10589 (N_10589,N_8076,N_6745);
nor U10590 (N_10590,N_9047,N_6535);
or U10591 (N_10591,N_8408,N_8837);
nand U10592 (N_10592,N_7320,N_8806);
or U10593 (N_10593,N_8238,N_7633);
nand U10594 (N_10594,N_6925,N_8458);
or U10595 (N_10595,N_6070,N_8725);
nand U10596 (N_10596,N_9456,N_6733);
nor U10597 (N_10597,N_9900,N_5077);
and U10598 (N_10598,N_8534,N_8573);
xnor U10599 (N_10599,N_6567,N_6600);
nand U10600 (N_10600,N_8464,N_5380);
nor U10601 (N_10601,N_8627,N_6565);
and U10602 (N_10602,N_8223,N_7968);
and U10603 (N_10603,N_7394,N_9412);
nor U10604 (N_10604,N_9515,N_5817);
and U10605 (N_10605,N_5284,N_8931);
and U10606 (N_10606,N_9721,N_5151);
or U10607 (N_10607,N_7168,N_6396);
or U10608 (N_10608,N_7174,N_8361);
or U10609 (N_10609,N_9980,N_6963);
and U10610 (N_10610,N_6377,N_8888);
and U10611 (N_10611,N_8319,N_8434);
nand U10612 (N_10612,N_7528,N_7833);
and U10613 (N_10613,N_7079,N_5447);
and U10614 (N_10614,N_5539,N_6524);
and U10615 (N_10615,N_6228,N_8119);
nor U10616 (N_10616,N_6731,N_7512);
nor U10617 (N_10617,N_6436,N_9967);
and U10618 (N_10618,N_9894,N_5422);
nand U10619 (N_10619,N_7582,N_5614);
or U10620 (N_10620,N_7006,N_8669);
or U10621 (N_10621,N_6447,N_5366);
nor U10622 (N_10622,N_8103,N_8445);
and U10623 (N_10623,N_6102,N_5136);
nand U10624 (N_10624,N_8402,N_7789);
nand U10625 (N_10625,N_6051,N_6903);
or U10626 (N_10626,N_6816,N_9488);
or U10627 (N_10627,N_9210,N_5094);
xor U10628 (N_10628,N_6862,N_6346);
nand U10629 (N_10629,N_7455,N_8664);
nand U10630 (N_10630,N_6149,N_6573);
nand U10631 (N_10631,N_8820,N_5178);
and U10632 (N_10632,N_8583,N_7655);
and U10633 (N_10633,N_6576,N_9609);
or U10634 (N_10634,N_9288,N_9133);
nand U10635 (N_10635,N_9854,N_7304);
nand U10636 (N_10636,N_8817,N_7420);
nand U10637 (N_10637,N_9287,N_6118);
nor U10638 (N_10638,N_5390,N_6809);
nor U10639 (N_10639,N_6453,N_5834);
nor U10640 (N_10640,N_6474,N_8953);
or U10641 (N_10641,N_7333,N_6012);
nand U10642 (N_10642,N_8428,N_5546);
and U10643 (N_10643,N_8475,N_6006);
or U10644 (N_10644,N_6247,N_6370);
nand U10645 (N_10645,N_9972,N_9679);
nand U10646 (N_10646,N_8647,N_8061);
and U10647 (N_10647,N_7276,N_6653);
and U10648 (N_10648,N_8618,N_6609);
or U10649 (N_10649,N_7022,N_5510);
nand U10650 (N_10650,N_5081,N_9000);
nand U10651 (N_10651,N_6984,N_8401);
or U10652 (N_10652,N_9921,N_5276);
and U10653 (N_10653,N_5932,N_5495);
nor U10654 (N_10654,N_8796,N_8718);
nor U10655 (N_10655,N_6466,N_5260);
or U10656 (N_10656,N_6311,N_5729);
or U10657 (N_10657,N_8770,N_6459);
xor U10658 (N_10658,N_8308,N_6182);
and U10659 (N_10659,N_8325,N_9298);
and U10660 (N_10660,N_6128,N_5292);
and U10661 (N_10661,N_8142,N_7880);
or U10662 (N_10662,N_6482,N_8122);
nor U10663 (N_10663,N_8449,N_6028);
and U10664 (N_10664,N_5357,N_8839);
nand U10665 (N_10665,N_8925,N_9708);
nand U10666 (N_10666,N_7111,N_5523);
nand U10667 (N_10667,N_8750,N_7490);
or U10668 (N_10668,N_9938,N_8713);
nand U10669 (N_10669,N_8333,N_7411);
nor U10670 (N_10670,N_6402,N_8163);
or U10671 (N_10671,N_9322,N_8522);
nor U10672 (N_10672,N_8115,N_8439);
and U10673 (N_10673,N_6936,N_8455);
nor U10674 (N_10674,N_6615,N_5378);
nor U10675 (N_10675,N_5943,N_8512);
nor U10676 (N_10676,N_7363,N_8679);
or U10677 (N_10677,N_6831,N_6201);
and U10678 (N_10678,N_7465,N_6718);
and U10679 (N_10679,N_9228,N_6944);
and U10680 (N_10680,N_8018,N_5503);
xor U10681 (N_10681,N_5242,N_7162);
and U10682 (N_10682,N_8979,N_8883);
nor U10683 (N_10683,N_7542,N_8017);
and U10684 (N_10684,N_9327,N_7038);
and U10685 (N_10685,N_7050,N_7695);
xor U10686 (N_10686,N_7359,N_6167);
and U10687 (N_10687,N_6749,N_8130);
nor U10688 (N_10688,N_5636,N_9215);
and U10689 (N_10689,N_6687,N_8851);
and U10690 (N_10690,N_8485,N_6302);
nor U10691 (N_10691,N_6000,N_7725);
and U10692 (N_10692,N_5870,N_5717);
xor U10693 (N_10693,N_8656,N_9428);
nor U10694 (N_10694,N_9431,N_7043);
and U10695 (N_10695,N_8247,N_8212);
and U10696 (N_10696,N_7422,N_6291);
nand U10697 (N_10697,N_9733,N_7389);
nor U10698 (N_10698,N_5146,N_8032);
nand U10699 (N_10699,N_6059,N_6445);
nand U10700 (N_10700,N_5014,N_7566);
and U10701 (N_10701,N_5166,N_9805);
and U10702 (N_10702,N_9263,N_5989);
and U10703 (N_10703,N_7735,N_6620);
or U10704 (N_10704,N_5212,N_5470);
nor U10705 (N_10705,N_9045,N_5335);
or U10706 (N_10706,N_7590,N_6358);
and U10707 (N_10707,N_7290,N_7259);
or U10708 (N_10708,N_6408,N_5846);
or U10709 (N_10709,N_5049,N_5900);
nor U10710 (N_10710,N_7780,N_9998);
nor U10711 (N_10711,N_9470,N_8624);
and U10712 (N_10712,N_5908,N_7092);
nand U10713 (N_10713,N_8704,N_7013);
or U10714 (N_10714,N_9749,N_8870);
nor U10715 (N_10715,N_8767,N_9162);
and U10716 (N_10716,N_5177,N_7375);
or U10717 (N_10717,N_7757,N_8549);
nor U10718 (N_10718,N_9630,N_7646);
nor U10719 (N_10719,N_6764,N_7640);
nor U10720 (N_10720,N_5468,N_8692);
and U10721 (N_10721,N_6709,N_5909);
nor U10722 (N_10722,N_5678,N_7584);
nor U10723 (N_10723,N_9002,N_9092);
nand U10724 (N_10724,N_9893,N_8995);
or U10725 (N_10725,N_7565,N_6593);
and U10726 (N_10726,N_7972,N_6058);
or U10727 (N_10727,N_7885,N_9587);
or U10728 (N_10728,N_9319,N_5039);
and U10729 (N_10729,N_7315,N_7228);
and U10730 (N_10730,N_6893,N_5676);
or U10731 (N_10731,N_6425,N_7404);
or U10732 (N_10732,N_5824,N_7231);
or U10733 (N_10733,N_7307,N_6452);
nor U10734 (N_10734,N_6101,N_5536);
and U10735 (N_10735,N_7957,N_5705);
nor U10736 (N_10736,N_9236,N_7224);
or U10737 (N_10737,N_9053,N_9830);
or U10738 (N_10738,N_6776,N_9789);
nor U10739 (N_10739,N_9846,N_9971);
and U10740 (N_10740,N_5716,N_5068);
nand U10741 (N_10741,N_8266,N_5406);
nand U10742 (N_10742,N_9529,N_8409);
and U10743 (N_10743,N_5947,N_6972);
nor U10744 (N_10744,N_9174,N_8662);
nand U10745 (N_10745,N_7083,N_5945);
nand U10746 (N_10746,N_6660,N_5596);
nor U10747 (N_10747,N_9915,N_5086);
nand U10748 (N_10748,N_6650,N_7869);
or U10749 (N_10749,N_9955,N_5156);
nand U10750 (N_10750,N_7128,N_9651);
or U10751 (N_10751,N_9459,N_6990);
and U10752 (N_10752,N_9782,N_7234);
and U10753 (N_10753,N_9535,N_6498);
or U10754 (N_10754,N_6940,N_5442);
nor U10755 (N_10755,N_8687,N_5024);
nor U10756 (N_10756,N_9123,N_7926);
nand U10757 (N_10757,N_9482,N_8660);
nor U10758 (N_10758,N_8262,N_6597);
nand U10759 (N_10759,N_7506,N_9037);
or U10760 (N_10760,N_7505,N_8731);
nor U10761 (N_10761,N_7053,N_6890);
nand U10762 (N_10762,N_5512,N_9430);
nand U10763 (N_10763,N_8170,N_9058);
nor U10764 (N_10764,N_7628,N_9248);
and U10765 (N_10765,N_8592,N_8463);
nor U10766 (N_10766,N_9256,N_5783);
and U10767 (N_10767,N_5225,N_5773);
or U10768 (N_10768,N_5364,N_6583);
nor U10769 (N_10769,N_7843,N_9907);
nor U10770 (N_10770,N_9827,N_6014);
xor U10771 (N_10771,N_8058,N_8961);
nand U10772 (N_10772,N_7286,N_5708);
nand U10773 (N_10773,N_9682,N_5542);
and U10774 (N_10774,N_8611,N_7556);
nand U10775 (N_10775,N_5352,N_5170);
nor U10776 (N_10776,N_9485,N_6860);
or U10777 (N_10777,N_5697,N_6643);
nor U10778 (N_10778,N_8087,N_6684);
nand U10779 (N_10779,N_6138,N_9757);
or U10780 (N_10780,N_6352,N_7414);
xor U10781 (N_10781,N_5672,N_5564);
nor U10782 (N_10782,N_6196,N_9520);
or U10783 (N_10783,N_9269,N_9878);
nor U10784 (N_10784,N_5937,N_8899);
or U10785 (N_10785,N_7951,N_6357);
nor U10786 (N_10786,N_8381,N_9561);
and U10787 (N_10787,N_6852,N_6048);
or U10788 (N_10788,N_6563,N_6153);
and U10789 (N_10789,N_7828,N_6721);
nand U10790 (N_10790,N_8379,N_6539);
nand U10791 (N_10791,N_9977,N_6544);
nand U10792 (N_10792,N_9478,N_9305);
nor U10793 (N_10793,N_9046,N_8610);
and U10794 (N_10794,N_9550,N_8785);
or U10795 (N_10795,N_6571,N_8964);
nand U10796 (N_10796,N_6191,N_5427);
xor U10797 (N_10797,N_5702,N_6663);
nand U10798 (N_10798,N_5287,N_6031);
nor U10799 (N_10799,N_6454,N_9754);
nor U10800 (N_10800,N_6569,N_5311);
or U10801 (N_10801,N_5594,N_7875);
or U10802 (N_10802,N_7609,N_5635);
nor U10803 (N_10803,N_7469,N_8741);
nand U10804 (N_10804,N_9597,N_7976);
nor U10805 (N_10805,N_9365,N_9525);
and U10806 (N_10806,N_5102,N_7382);
and U10807 (N_10807,N_6818,N_6853);
nor U10808 (N_10808,N_6536,N_9704);
nor U10809 (N_10809,N_9819,N_9043);
and U10810 (N_10810,N_5797,N_5430);
or U10811 (N_10811,N_5563,N_6943);
nand U10812 (N_10812,N_7331,N_5691);
and U10813 (N_10813,N_6364,N_7132);
or U10814 (N_10814,N_5884,N_6379);
and U10815 (N_10815,N_5959,N_5795);
nand U10816 (N_10816,N_7215,N_9575);
and U10817 (N_10817,N_9085,N_8129);
and U10818 (N_10818,N_8260,N_6309);
nand U10819 (N_10819,N_9727,N_6798);
nand U10820 (N_10820,N_8168,N_9030);
nor U10821 (N_10821,N_5608,N_6183);
xor U10822 (N_10822,N_5471,N_9408);
nor U10823 (N_10823,N_5358,N_5524);
or U10824 (N_10824,N_5463,N_6293);
nor U10825 (N_10825,N_7023,N_8951);
or U10826 (N_10826,N_5277,N_9124);
or U10827 (N_10827,N_5589,N_6409);
nor U10828 (N_10828,N_6461,N_7379);
and U10829 (N_10829,N_5065,N_8608);
nor U10830 (N_10830,N_5516,N_7220);
xnor U10831 (N_10831,N_9032,N_9872);
or U10832 (N_10832,N_7475,N_8231);
and U10833 (N_10833,N_7126,N_5926);
or U10834 (N_10834,N_7374,N_8305);
nand U10835 (N_10835,N_9709,N_6851);
nor U10836 (N_10836,N_6928,N_5232);
nand U10837 (N_10837,N_5760,N_5181);
nor U10838 (N_10838,N_9772,N_7412);
or U10839 (N_10839,N_9820,N_5933);
and U10840 (N_10840,N_5278,N_9610);
and U10841 (N_10841,N_7579,N_9293);
or U10842 (N_10842,N_7417,N_7352);
and U10843 (N_10843,N_7681,N_8634);
nor U10844 (N_10844,N_6044,N_5409);
nor U10845 (N_10845,N_6197,N_6465);
and U10846 (N_10846,N_8562,N_9148);
nor U10847 (N_10847,N_6433,N_5577);
nor U10848 (N_10848,N_6292,N_9068);
nand U10849 (N_10849,N_8338,N_7317);
nor U10850 (N_10850,N_8191,N_5441);
and U10851 (N_10851,N_6638,N_6035);
or U10852 (N_10852,N_9493,N_8482);
nor U10853 (N_10853,N_6160,N_7078);
nor U10854 (N_10854,N_6614,N_9386);
or U10855 (N_10855,N_5960,N_6017);
nor U10856 (N_10856,N_9150,N_7295);
nor U10857 (N_10857,N_8495,N_7134);
or U10858 (N_10858,N_6002,N_5387);
or U10859 (N_10859,N_8552,N_7318);
and U10860 (N_10860,N_8193,N_5558);
or U10861 (N_10861,N_6040,N_9637);
and U10862 (N_10862,N_5855,N_5310);
or U10863 (N_10863,N_8921,N_6560);
nor U10864 (N_10864,N_7895,N_5339);
and U10865 (N_10865,N_8754,N_7060);
and U10866 (N_10866,N_7537,N_9539);
nand U10867 (N_10867,N_6207,N_5108);
or U10868 (N_10868,N_9325,N_7759);
and U10869 (N_10869,N_5894,N_9258);
nand U10870 (N_10870,N_6835,N_7035);
nand U10871 (N_10871,N_7660,N_8738);
and U10872 (N_10872,N_5806,N_5297);
xnor U10873 (N_10873,N_7914,N_5344);
nand U10874 (N_10874,N_7196,N_6363);
nand U10875 (N_10875,N_6455,N_5132);
nand U10876 (N_10876,N_8389,N_5403);
or U10877 (N_10877,N_7888,N_8942);
nor U10878 (N_10878,N_7595,N_8372);
nand U10879 (N_10879,N_7099,N_6368);
nand U10880 (N_10880,N_5659,N_9618);
and U10881 (N_10881,N_5597,N_8818);
xnor U10882 (N_10882,N_7210,N_5143);
and U10883 (N_10883,N_6255,N_8358);
nand U10884 (N_10884,N_7471,N_5453);
nor U10885 (N_10885,N_8991,N_6870);
nor U10886 (N_10886,N_7086,N_8356);
or U10887 (N_10887,N_6899,N_9227);
nand U10888 (N_10888,N_5219,N_5598);
xor U10889 (N_10889,N_8698,N_8281);
or U10890 (N_10890,N_9193,N_7925);
or U10891 (N_10891,N_6094,N_8598);
nand U10892 (N_10892,N_7818,N_5613);
nor U10893 (N_10893,N_7567,N_6758);
and U10894 (N_10894,N_7395,N_8779);
and U10895 (N_10895,N_6879,N_9108);
nand U10896 (N_10896,N_9764,N_6520);
nor U10897 (N_10897,N_9407,N_6577);
nand U10898 (N_10898,N_8867,N_5353);
nand U10899 (N_10899,N_6800,N_9217);
or U10900 (N_10900,N_7649,N_9523);
and U10901 (N_10901,N_7544,N_7330);
and U10902 (N_10902,N_9832,N_8816);
nand U10903 (N_10903,N_8341,N_7346);
xor U10904 (N_10904,N_9301,N_7069);
nand U10905 (N_10905,N_6929,N_6589);
nor U10906 (N_10906,N_6231,N_8996);
nor U10907 (N_10907,N_7093,N_9309);
and U10908 (N_10908,N_8575,N_6130);
and U10909 (N_10909,N_9840,N_7643);
nand U10910 (N_10910,N_5456,N_9244);
nand U10911 (N_10911,N_5368,N_9945);
or U10912 (N_10912,N_6648,N_7545);
or U10913 (N_10913,N_5006,N_6369);
xnor U10914 (N_10914,N_8336,N_5713);
nor U10915 (N_10915,N_9593,N_5252);
xnor U10916 (N_10916,N_9865,N_8451);
and U10917 (N_10917,N_9010,N_7714);
nor U10918 (N_10918,N_8441,N_8282);
or U10919 (N_10919,N_9070,N_8700);
nor U10920 (N_10920,N_6768,N_6946);
xnor U10921 (N_10921,N_9634,N_8570);
nor U10922 (N_10922,N_5461,N_6406);
and U10923 (N_10923,N_6916,N_9049);
nor U10924 (N_10924,N_9718,N_8433);
or U10925 (N_10925,N_9540,N_8538);
and U10926 (N_10926,N_5565,N_9898);
nand U10927 (N_10927,N_5784,N_8852);
nand U10928 (N_10928,N_8049,N_5876);
nand U10929 (N_10929,N_8473,N_9926);
nand U10930 (N_10930,N_7137,N_5703);
and U10931 (N_10931,N_9357,N_5443);
nand U10932 (N_10932,N_9917,N_5557);
or U10933 (N_10933,N_9181,N_8544);
nor U10934 (N_10934,N_8503,N_8882);
xor U10935 (N_10935,N_9323,N_7370);
and U10936 (N_10936,N_8886,N_8758);
nor U10937 (N_10937,N_5064,N_9781);
nand U10938 (N_10938,N_6808,N_5254);
nand U10939 (N_10939,N_6842,N_5230);
nand U10940 (N_10940,N_6176,N_6367);
nand U10941 (N_10941,N_6515,N_8436);
nand U10942 (N_10942,N_6192,N_7511);
or U10943 (N_10943,N_9991,N_5862);
nor U10944 (N_10944,N_6989,N_5865);
nor U10945 (N_10945,N_6825,N_8588);
or U10946 (N_10946,N_7296,N_6164);
and U10947 (N_10947,N_7762,N_5978);
and U10948 (N_10948,N_5799,N_7601);
or U10949 (N_10949,N_5245,N_9615);
nor U10950 (N_10950,N_8472,N_9427);
nand U10951 (N_10951,N_8620,N_6543);
nor U10952 (N_10952,N_7540,N_6260);
nor U10953 (N_10953,N_6434,N_5003);
nor U10954 (N_10954,N_8437,N_8809);
and U10955 (N_10955,N_7265,N_7657);
or U10956 (N_10956,N_7675,N_8565);
or U10957 (N_10957,N_7400,N_7325);
or U10958 (N_10958,N_5619,N_8328);
nor U10959 (N_10959,N_5912,N_6875);
nand U10960 (N_10960,N_9267,N_7364);
nor U10961 (N_10961,N_6230,N_6784);
nand U10962 (N_10962,N_9588,N_9516);
or U10963 (N_10963,N_9201,N_9512);
xor U10964 (N_10964,N_5903,N_5741);
nand U10965 (N_10965,N_8601,N_9329);
or U10966 (N_10966,N_8124,N_7036);
nand U10967 (N_10967,N_8154,N_7855);
nand U10968 (N_10968,N_9041,N_6547);
or U10969 (N_10969,N_8213,N_5037);
and U10970 (N_10970,N_6312,N_5786);
nor U10971 (N_10971,N_8603,N_5990);
and U10972 (N_10972,N_6194,N_7255);
nand U10973 (N_10973,N_8340,N_8771);
nand U10974 (N_10974,N_9132,N_7922);
xor U10975 (N_10975,N_9311,N_5031);
nand U10976 (N_10976,N_6658,N_7523);
nor U10977 (N_10977,N_7909,N_6833);
nor U10978 (N_10978,N_8525,N_5373);
nand U10979 (N_10979,N_9680,N_5091);
or U10980 (N_10980,N_8317,N_5574);
nand U10981 (N_10981,N_8990,N_6158);
nor U10982 (N_10982,N_7393,N_9717);
nor U10983 (N_10983,N_5238,N_8541);
or U10984 (N_10984,N_9450,N_5263);
or U10985 (N_10985,N_6606,N_9856);
nor U10986 (N_10986,N_8029,N_5053);
or U10987 (N_10987,N_7907,N_9836);
and U10988 (N_10988,N_6239,N_7949);
or U10989 (N_10989,N_8854,N_9844);
nand U10990 (N_10990,N_5948,N_9650);
and U10991 (N_10991,N_9775,N_7345);
nand U10992 (N_10992,N_6974,N_8710);
nand U10993 (N_10993,N_5822,N_9956);
and U10994 (N_10994,N_6891,N_9808);
and U10995 (N_10995,N_7353,N_6407);
and U10996 (N_10996,N_8236,N_7650);
nand U10997 (N_10997,N_5030,N_5838);
or U10998 (N_10998,N_7848,N_7146);
nor U10999 (N_10999,N_8202,N_5100);
nor U11000 (N_11000,N_9642,N_9803);
and U11001 (N_11001,N_6812,N_7279);
nor U11002 (N_11002,N_6073,N_5165);
or U11003 (N_11003,N_8553,N_7934);
nor U11004 (N_11004,N_8222,N_6630);
nand U11005 (N_11005,N_7719,N_6777);
nand U11006 (N_11006,N_8533,N_5154);
and U11007 (N_11007,N_8863,N_6846);
xnor U11008 (N_11008,N_8600,N_9433);
nand U11009 (N_11009,N_8947,N_7270);
or U11010 (N_11010,N_7284,N_9541);
or U11011 (N_11011,N_8784,N_7048);
or U11012 (N_11012,N_5180,N_7618);
nor U11013 (N_11013,N_7696,N_5548);
and U11014 (N_11014,N_7002,N_6640);
and U11015 (N_11015,N_5467,N_5391);
or U11016 (N_11016,N_6273,N_5790);
xnor U11017 (N_11017,N_6559,N_5997);
nor U11018 (N_11018,N_8293,N_8460);
nor U11019 (N_11019,N_9388,N_9671);
or U11020 (N_11020,N_7335,N_7677);
nand U11021 (N_11021,N_5382,N_5759);
and U11022 (N_11022,N_5898,N_7011);
or U11023 (N_11023,N_6344,N_5419);
or U11024 (N_11024,N_6262,N_9880);
nor U11025 (N_11025,N_8342,N_8591);
and U11026 (N_11026,N_8778,N_7339);
and U11027 (N_11027,N_5172,N_7007);
nor U11028 (N_11028,N_6610,N_5988);
or U11029 (N_11029,N_8466,N_8310);
nor U11030 (N_11030,N_5609,N_6403);
nor U11031 (N_11031,N_7323,N_7495);
nand U11032 (N_11032,N_7249,N_6241);
and U11033 (N_11033,N_6965,N_9766);
nor U11034 (N_11034,N_8404,N_9981);
or U11035 (N_11035,N_9970,N_8162);
nor U11036 (N_11036,N_5889,N_5472);
and U11037 (N_11037,N_8136,N_8435);
and U11038 (N_11038,N_7860,N_8301);
and U11039 (N_11039,N_5474,N_6097);
xor U11040 (N_11040,N_7726,N_7611);
nand U11041 (N_11041,N_8010,N_8090);
nor U11042 (N_11042,N_6018,N_9794);
and U11043 (N_11043,N_6557,N_5079);
and U11044 (N_11044,N_9320,N_9841);
or U11045 (N_11045,N_6739,N_9882);
nand U11046 (N_11046,N_9986,N_8594);
nor U11047 (N_11047,N_7546,N_8149);
or U11048 (N_11048,N_8430,N_9993);
nand U11049 (N_11049,N_6973,N_8606);
nor U11050 (N_11050,N_6730,N_6632);
and U11051 (N_11051,N_6360,N_9340);
nor U11052 (N_11052,N_8523,N_6672);
nand U11053 (N_11053,N_5318,N_7724);
nor U11054 (N_11054,N_7081,N_6401);
or U11055 (N_11055,N_5547,N_9728);
nand U11056 (N_11056,N_7890,N_5458);
nor U11057 (N_11057,N_7485,N_7481);
nand U11058 (N_11058,N_5308,N_9469);
nor U11059 (N_11059,N_7403,N_8590);
nor U11060 (N_11060,N_6429,N_7147);
nand U11061 (N_11061,N_9702,N_9595);
nand U11062 (N_11062,N_9460,N_5294);
nand U11063 (N_11063,N_9960,N_9044);
nor U11064 (N_11064,N_5423,N_6581);
or U11065 (N_11065,N_9185,N_5404);
nand U11066 (N_11066,N_5998,N_6788);
nor U11067 (N_11067,N_8484,N_8810);
nand U11068 (N_11068,N_8905,N_8045);
or U11069 (N_11069,N_9877,N_5951);
nor U11070 (N_11070,N_7009,N_9519);
nor U11071 (N_11071,N_6661,N_9683);
nor U11072 (N_11072,N_9719,N_5849);
nand U11073 (N_11073,N_6003,N_8025);
nand U11074 (N_11074,N_7016,N_8936);
nand U11075 (N_11075,N_6320,N_5888);
nand U11076 (N_11076,N_9743,N_6590);
nand U11077 (N_11077,N_5852,N_6208);
or U11078 (N_11078,N_9443,N_8352);
or U11079 (N_11079,N_9404,N_5038);
or U11080 (N_11080,N_6242,N_6331);
nand U11081 (N_11081,N_6204,N_6824);
nor U11082 (N_11082,N_9219,N_5582);
nor U11083 (N_11083,N_9291,N_8760);
nand U11084 (N_11084,N_7029,N_7449);
and U11085 (N_11085,N_7825,N_5910);
nand U11086 (N_11086,N_9326,N_9352);
xor U11087 (N_11087,N_7899,N_9360);
or U11088 (N_11088,N_7256,N_7165);
nand U11089 (N_11089,N_5105,N_6935);
nor U11090 (N_11090,N_9596,N_8192);
or U11091 (N_11091,N_8442,N_6480);
or U11092 (N_11092,N_5617,N_8210);
nand U11093 (N_11093,N_6021,N_9798);
nand U11094 (N_11094,N_7232,N_9816);
nand U11095 (N_11095,N_8075,N_8037);
and U11096 (N_11096,N_5251,N_8327);
or U11097 (N_11097,N_8505,N_9667);
and U11098 (N_11098,N_9199,N_9531);
nand U11099 (N_11099,N_7748,N_6780);
nor U11100 (N_11100,N_7670,N_8461);
or U11101 (N_11101,N_7613,N_9397);
nand U11102 (N_11102,N_8545,N_5027);
and U11103 (N_11103,N_9069,N_9268);
or U11104 (N_11104,N_5688,N_7001);
nand U11105 (N_11105,N_8376,N_8977);
or U11106 (N_11106,N_7456,N_6674);
and U11107 (N_11107,N_6885,N_8900);
nand U11108 (N_11108,N_5098,N_8476);
and U11109 (N_11109,N_7230,N_7807);
nor U11110 (N_11110,N_5982,N_7221);
and U11111 (N_11111,N_9674,N_8295);
or U11112 (N_11112,N_9569,N_8151);
nand U11113 (N_11113,N_7066,N_6356);
or U11114 (N_11114,N_5832,N_7399);
or U11115 (N_11115,N_6166,N_5861);
nor U11116 (N_11116,N_8876,N_8249);
nor U11117 (N_11117,N_5687,N_6093);
or U11118 (N_11118,N_9350,N_5685);
and U11119 (N_11119,N_5793,N_5087);
and U11120 (N_11120,N_5917,N_8637);
and U11121 (N_11121,N_9208,N_6200);
nor U11122 (N_11122,N_7754,N_7310);
nand U11123 (N_11123,N_6055,N_6096);
and U11124 (N_11124,N_7692,N_8137);
and U11125 (N_11125,N_8672,N_8871);
and U11126 (N_11126,N_8508,N_5424);
nand U11127 (N_11127,N_6627,N_5117);
and U11128 (N_11128,N_7815,N_8511);
nand U11129 (N_11129,N_9336,N_5121);
and U11130 (N_11130,N_5323,N_9307);
or U11131 (N_11131,N_9159,N_7648);
and U11132 (N_11132,N_6275,N_7261);
or U11133 (N_11133,N_8639,N_8649);
or U11134 (N_11134,N_9812,N_6856);
and U11135 (N_11135,N_9912,N_6472);
nand U11136 (N_11136,N_7965,N_8244);
nand U11137 (N_11137,N_9594,N_9249);
and U11138 (N_11138,N_7771,N_5690);
nor U11139 (N_11139,N_8276,N_6554);
nand U11140 (N_11140,N_7859,N_9589);
nor U11141 (N_11141,N_9499,N_8872);
nand U11142 (N_11142,N_5505,N_5873);
or U11143 (N_11143,N_9284,N_8383);
nand U11144 (N_11144,N_8406,N_7017);
nand U11145 (N_11145,N_8814,N_7610);
or U11146 (N_11146,N_7206,N_6967);
nor U11147 (N_11147,N_5774,N_6724);
nor U11148 (N_11148,N_6591,N_6148);
or U11149 (N_11149,N_6326,N_6289);
nor U11150 (N_11150,N_5015,N_6282);
or U11151 (N_11151,N_9617,N_6339);
nand U11152 (N_11152,N_8556,N_7452);
and U11153 (N_11153,N_8892,N_6516);
and U11154 (N_11154,N_8127,N_7684);
nor U11155 (N_11155,N_8519,N_8958);
or U11156 (N_11156,N_8006,N_5499);
or U11157 (N_11157,N_7733,N_5804);
nor U11158 (N_11158,N_8499,N_5106);
nand U11159 (N_11159,N_9093,N_7961);
nand U11160 (N_11160,N_9685,N_6604);
or U11161 (N_11161,N_8623,N_5952);
and U11162 (N_11162,N_9194,N_8965);
nor U11163 (N_11163,N_8557,N_6701);
and U11164 (N_11164,N_8630,N_8250);
nor U11165 (N_11165,N_6680,N_8307);
nor U11166 (N_11166,N_9620,N_7973);
xor U11167 (N_11167,N_5706,N_6960);
xnor U11168 (N_11168,N_8391,N_9950);
nor U11169 (N_11169,N_7728,N_6694);
nand U11170 (N_11170,N_5813,N_7564);
and U11171 (N_11171,N_6697,N_8955);
nor U11172 (N_11172,N_7721,N_7904);
and U11173 (N_11173,N_8543,N_5554);
nand U11174 (N_11174,N_5875,N_6491);
and U11175 (N_11175,N_6274,N_8330);
and U11176 (N_11176,N_6226,N_9983);
and U11177 (N_11177,N_8107,N_9461);
or U11178 (N_11178,N_8268,N_9884);
nor U11179 (N_11179,N_9209,N_8015);
nor U11180 (N_11180,N_5528,N_6526);
nor U11181 (N_11181,N_8677,N_6423);
and U11182 (N_11182,N_5274,N_9467);
or U11183 (N_11183,N_8786,N_5568);
nand U11184 (N_11184,N_7827,N_8982);
and U11185 (N_11185,N_5532,N_9304);
nand U11186 (N_11186,N_7886,N_6155);
and U11187 (N_11187,N_9164,N_7863);
nand U11188 (N_11188,N_5211,N_6168);
or U11189 (N_11189,N_7037,N_5199);
and U11190 (N_11190,N_5249,N_7329);
or U11191 (N_11191,N_5668,N_9765);
and U11192 (N_11192,N_9625,N_9358);
and U11193 (N_11193,N_5728,N_5803);
nor U11194 (N_11194,N_6601,N_9638);
or U11195 (N_11195,N_5551,N_9101);
or U11196 (N_11196,N_5115,N_7524);
nand U11197 (N_11197,N_7073,N_7477);
xor U11198 (N_11198,N_5750,N_7585);
nor U11199 (N_11199,N_9626,N_7982);
or U11200 (N_11200,N_5587,N_7765);
and U11201 (N_11201,N_7237,N_7362);
and U11202 (N_11202,N_6100,N_9019);
and U11203 (N_11203,N_7813,N_5921);
or U11204 (N_11204,N_5867,N_5899);
and U11205 (N_11205,N_7837,N_5922);
and U11206 (N_11206,N_6765,N_8245);
nand U11207 (N_11207,N_8976,N_8962);
or U11208 (N_11208,N_6909,N_9504);
nor U11209 (N_11209,N_7144,N_7919);
nand U11210 (N_11210,N_6654,N_5842);
or U11211 (N_11211,N_6922,N_8835);
nand U11212 (N_11212,N_8743,N_9745);
and U11213 (N_11213,N_5476,N_5623);
or U11214 (N_11214,N_8471,N_6656);
nand U11215 (N_11215,N_8827,N_8651);
and U11216 (N_11216,N_7084,N_6421);
or U11217 (N_11217,N_6108,N_8367);
nand U11218 (N_11218,N_8273,N_8446);
nor U11219 (N_11219,N_8671,N_9759);
nor U11220 (N_11220,N_7990,N_5214);
and U11221 (N_11221,N_6713,N_8407);
or U11222 (N_11222,N_8106,N_9590);
nor U11223 (N_11223,N_9361,N_8587);
and U11224 (N_11224,N_6151,N_7181);
nand U11225 (N_11225,N_6224,N_9220);
nor U11226 (N_11226,N_6476,N_5714);
nand U11227 (N_11227,N_6621,N_7172);
nand U11228 (N_11228,N_9339,N_8569);
nor U11229 (N_11229,N_8673,N_7760);
and U11230 (N_11230,N_6912,N_6043);
and U11231 (N_11231,N_8819,N_7077);
nor U11232 (N_11232,N_5233,N_5666);
or U11233 (N_11233,N_7313,N_9503);
nand U11234 (N_11234,N_9859,N_5059);
and U11235 (N_11235,N_8759,N_6448);
and U11236 (N_11236,N_5872,N_5747);
nand U11237 (N_11237,N_8044,N_8283);
and U11238 (N_11238,N_5840,N_9785);
and U11239 (N_11239,N_7701,N_5695);
and U11240 (N_11240,N_5141,N_6026);
nand U11241 (N_11241,N_8148,N_9712);
nor U11242 (N_11242,N_8186,N_7299);
and U11243 (N_11243,N_7580,N_8318);
nor U11244 (N_11244,N_6931,N_7064);
and U11245 (N_11245,N_8681,N_6022);
nand U11246 (N_11246,N_9035,N_6993);
and U11247 (N_11247,N_7788,N_7327);
nand U11248 (N_11248,N_7110,N_9649);
nor U11249 (N_11249,N_5991,N_8748);
nand U11250 (N_11250,N_5622,N_8937);
nor U11251 (N_11251,N_5916,N_9632);
nand U11252 (N_11252,N_9048,N_8071);
nand U11253 (N_11253,N_9203,N_8701);
nand U11254 (N_11254,N_7263,N_8842);
and U11255 (N_11255,N_5970,N_5976);
nor U11256 (N_11256,N_7182,N_6234);
or U11257 (N_11257,N_8884,N_7179);
nor U11258 (N_11258,N_7450,N_5365);
or U11259 (N_11259,N_6217,N_7900);
or U11260 (N_11260,N_8348,N_9598);
or U11261 (N_11261,N_9730,N_7205);
nand U11262 (N_11262,N_6854,N_5479);
and U11263 (N_11263,N_9257,N_7878);
nand U11264 (N_11264,N_9299,N_8343);
nand U11265 (N_11265,N_8265,N_5303);
and U11266 (N_11266,N_8187,N_9752);
nor U11267 (N_11267,N_6933,N_8739);
and U11268 (N_11268,N_7711,N_9142);
nand U11269 (N_11269,N_7865,N_5054);
or U11270 (N_11270,N_5780,N_7021);
or U11271 (N_11271,N_8359,N_9211);
nor U11272 (N_11272,N_8693,N_6956);
xor U11273 (N_11273,N_9090,N_6010);
nor U11274 (N_11274,N_6582,N_7797);
and U11275 (N_11275,N_8537,N_5007);
and U11276 (N_11276,N_8135,N_9270);
or U11277 (N_11277,N_6488,N_6947);
and U11278 (N_11278,N_8014,N_5392);
and U11279 (N_11279,N_7729,N_6471);
and U11280 (N_11280,N_8392,N_8504);
nor U11281 (N_11281,N_5041,N_8638);
and U11282 (N_11282,N_8769,N_6580);
and U11283 (N_11283,N_8735,N_5935);
nand U11284 (N_11284,N_5018,N_8683);
nand U11285 (N_11285,N_5073,N_8548);
nand U11286 (N_11286,N_7487,N_6125);
nor U11287 (N_11287,N_6920,N_8957);
and U11288 (N_11288,N_6518,N_9166);
and U11289 (N_11289,N_5811,N_8011);
nand U11290 (N_11290,N_5969,N_5514);
or U11291 (N_11291,N_9903,N_5220);
and U11292 (N_11292,N_6306,N_5519);
nor U11293 (N_11293,N_9224,N_7879);
or U11294 (N_11294,N_9552,N_9564);
or U11295 (N_11295,N_8826,N_9229);
nor U11296 (N_11296,N_9154,N_8322);
or U11297 (N_11297,N_5057,N_9465);
nand U11298 (N_11298,N_9506,N_9139);
nand U11299 (N_11299,N_6850,N_6229);
nand U11300 (N_11300,N_6198,N_5213);
nand U11301 (N_11301,N_8946,N_6827);
nor U11302 (N_11302,N_5044,N_7525);
nor U11303 (N_11303,N_7768,N_9377);
nor U11304 (N_11304,N_7219,N_7519);
and U11305 (N_11305,N_7882,N_6847);
and U11306 (N_11306,N_6276,N_5630);
nor U11307 (N_11307,N_6393,N_8294);
nor U11308 (N_11308,N_9624,N_5237);
and U11309 (N_11309,N_5656,N_7120);
nand U11310 (N_11310,N_9574,N_6075);
or U11311 (N_11311,N_8906,N_7291);
nor U11312 (N_11312,N_5552,N_6313);
nor U11313 (N_11313,N_8987,N_9266);
nor U11314 (N_11314,N_5491,N_8821);
nor U11315 (N_11315,N_5492,N_5661);
or U11316 (N_11316,N_9692,N_7489);
nor U11317 (N_11317,N_8204,N_8146);
or U11318 (N_11318,N_5634,N_7631);
nor U11319 (N_11319,N_6790,N_9038);
nand U11320 (N_11320,N_8048,N_6080);
nor U11321 (N_11321,N_7464,N_8706);
or U11322 (N_11322,N_5566,N_6914);
nand U11323 (N_11323,N_7257,N_7247);
and U11324 (N_11324,N_7445,N_9847);
nand U11325 (N_11325,N_7442,N_8128);
or U11326 (N_11326,N_5231,N_6706);
and U11327 (N_11327,N_9726,N_6820);
and U11328 (N_11328,N_5393,N_7075);
or U11329 (N_11329,N_8069,N_8928);
or U11330 (N_11330,N_9599,N_7702);
or U11331 (N_11331,N_7342,N_5019);
nand U11332 (N_11332,N_6400,N_9289);
nor U11333 (N_11333,N_6913,N_9885);
nor U11334 (N_11334,N_9188,N_8514);
nor U11335 (N_11335,N_5394,N_5229);
and U11336 (N_11336,N_7095,N_5349);
nand U11337 (N_11337,N_8346,N_6637);
nor U11338 (N_11338,N_9946,N_7647);
nor U11339 (N_11339,N_5950,N_5700);
or U11340 (N_11340,N_6213,N_7461);
and U11341 (N_11341,N_8917,N_7852);
or U11342 (N_11342,N_8125,N_5281);
or U11343 (N_11343,N_7756,N_5987);
nand U11344 (N_11344,N_9155,N_9853);
or U11345 (N_11345,N_9834,N_8585);
and U11346 (N_11346,N_5721,N_8577);
and U11347 (N_11347,N_5979,N_7570);
or U11348 (N_11348,N_8092,N_8912);
nand U11349 (N_11349,N_5792,N_9817);
nor U11350 (N_11350,N_7088,N_8644);
or U11351 (N_11351,N_5831,N_9670);
nand U11352 (N_11352,N_7371,N_8396);
nand U11353 (N_11353,N_5191,N_9863);
or U11354 (N_11354,N_8528,N_9511);
nand U11355 (N_11355,N_5961,N_6284);
nor U11356 (N_11356,N_8813,N_9799);
and U11357 (N_11357,N_6374,N_7082);
nand U11358 (N_11358,N_6746,N_8877);
nor U11359 (N_11359,N_7853,N_8703);
and U11360 (N_11360,N_8761,N_7446);
nor U11361 (N_11361,N_8970,N_9118);
nor U11362 (N_11362,N_6371,N_7435);
nand U11363 (N_11363,N_6308,N_6826);
nor U11364 (N_11364,N_5017,N_7727);
nand U11365 (N_11365,N_5020,N_6105);
nand U11366 (N_11366,N_5329,N_6264);
nor U11367 (N_11367,N_6690,N_9232);
nor U11368 (N_11368,N_7254,N_8986);
and U11369 (N_11369,N_7572,N_7312);
and U11370 (N_11370,N_9737,N_6330);
or U11371 (N_11371,N_5525,N_6592);
and U11372 (N_11372,N_8985,N_7822);
or U11373 (N_11373,N_8654,N_7503);
or U11374 (N_11374,N_7686,N_7887);
or U11375 (N_11375,N_5965,N_7672);
nand U11376 (N_11376,N_8763,N_9833);
and U11377 (N_11377,N_6819,N_9978);
nor U11378 (N_11378,N_9399,N_6185);
nand U11379 (N_11379,N_8916,N_8467);
nand U11380 (N_11380,N_8967,N_5302);
nand U11381 (N_11381,N_7246,N_7218);
nand U11382 (N_11382,N_7439,N_9952);
or U11383 (N_11383,N_9791,N_5854);
nor U11384 (N_11384,N_6930,N_9948);
nor U11385 (N_11385,N_9064,N_5938);
and U11386 (N_11386,N_7376,N_7140);
nor U11387 (N_11387,N_6867,N_8321);
or U11388 (N_11388,N_6419,N_9389);
nor U11389 (N_11389,N_7473,N_6383);
or U11390 (N_11390,N_5901,N_6157);
and U11391 (N_11391,N_9838,N_8291);
and U11392 (N_11392,N_9082,N_6211);
nand U11393 (N_11393,N_5138,N_6622);
nand U11394 (N_11394,N_8429,N_9278);
and U11395 (N_11395,N_7258,N_9631);
and U11396 (N_11396,N_7997,N_5850);
nand U11397 (N_11397,N_6530,N_6811);
nand U11398 (N_11398,N_6886,N_8456);
nand U11399 (N_11399,N_8765,N_7378);
nand U11400 (N_11400,N_5610,N_9471);
and U11401 (N_11401,N_5016,N_8992);
nor U11402 (N_11402,N_8781,N_8070);
or U11403 (N_11403,N_5464,N_7980);
nor U11404 (N_11404,N_5679,N_8468);
nor U11405 (N_11405,N_8004,N_8078);
nand U11406 (N_11406,N_8728,N_8551);
or U11407 (N_11407,N_9509,N_9501);
and U11408 (N_11408,N_6932,N_6728);
nand U11409 (N_11409,N_7520,N_7157);
and U11410 (N_11410,N_9195,N_6416);
or U11411 (N_11411,N_8285,N_6652);
nor U11412 (N_11412,N_8762,N_8176);
or U11413 (N_11413,N_7358,N_5487);
and U11414 (N_11414,N_5829,N_9453);
nor U11415 (N_11415,N_8074,N_5663);
nor U11416 (N_11416,N_9557,N_8002);
nand U11417 (N_11417,N_6117,N_9522);
or U11418 (N_11418,N_7125,N_8773);
nor U11419 (N_11419,N_9690,N_5620);
nor U11420 (N_11420,N_7658,N_7616);
nor U11421 (N_11421,N_7576,N_5507);
nand U11422 (N_11422,N_6236,N_5347);
and U11423 (N_11423,N_8531,N_7217);
nand U11424 (N_11424,N_8932,N_7829);
and U11425 (N_11425,N_5538,N_7948);
nand U11426 (N_11426,N_7824,N_6050);
or U11427 (N_11427,N_7864,N_5974);
xnor U11428 (N_11428,N_9810,N_6992);
and U11429 (N_11429,N_5830,N_7942);
nor U11430 (N_11430,N_6004,N_9942);
nand U11431 (N_11431,N_5185,N_7614);
or U11432 (N_11432,N_9628,N_6975);
or U11433 (N_11433,N_6477,N_8555);
or U11434 (N_11434,N_7975,N_6442);
nor U11435 (N_11435,N_9559,N_5417);
nand U11436 (N_11436,N_5362,N_5556);
nand U11437 (N_11437,N_5291,N_6333);
and U11438 (N_11438,N_8431,N_5805);
nor U11439 (N_11439,N_7669,N_6553);
and U11440 (N_11440,N_9374,N_7928);
and U11441 (N_11441,N_8263,N_7223);
nor U11442 (N_11442,N_9779,N_9423);
and U11443 (N_11443,N_6388,N_6141);
nor U11444 (N_11444,N_6205,N_8721);
and U11445 (N_11445,N_7836,N_8418);
or U11446 (N_11446,N_7782,N_7354);
nand U11447 (N_11447,N_9177,N_6815);
and U11448 (N_11448,N_7423,N_7213);
nor U11449 (N_11449,N_6470,N_9454);
nand U11450 (N_11450,N_6773,N_7138);
nand U11451 (N_11451,N_7974,N_8621);
nor U11452 (N_11452,N_6813,N_5070);
or U11453 (N_11453,N_5821,N_9464);
or U11454 (N_11454,N_8300,N_5361);
nor U11455 (N_11455,N_6265,N_9440);
or U11456 (N_11456,N_5286,N_6256);
nor U11457 (N_11457,N_9551,N_7204);
nor U11458 (N_11458,N_6145,N_9056);
and U11459 (N_11459,N_9187,N_6353);
nor U11460 (N_11460,N_9253,N_9112);
nand U11461 (N_11461,N_6555,N_5863);
and U11462 (N_11462,N_7665,N_5595);
or U11463 (N_11463,N_6700,N_6072);
nand U11464 (N_11464,N_7644,N_7431);
nand U11465 (N_11465,N_9363,N_6481);
and U11466 (N_11466,N_7235,N_6970);
nand U11467 (N_11467,N_5193,N_5208);
and U11468 (N_11468,N_6249,N_6152);
nor U11469 (N_11469,N_5076,N_9776);
nor U11470 (N_11470,N_8038,N_7480);
or U11471 (N_11471,N_6299,N_9400);
or U11472 (N_11472,N_9372,N_6209);
nor U11473 (N_11473,N_9581,N_8082);
and U11474 (N_11474,N_6506,N_7028);
or U11475 (N_11475,N_5967,N_8715);
nor U11476 (N_11476,N_5845,N_5469);
or U11477 (N_11477,N_5743,N_8873);
and U11478 (N_11478,N_9807,N_5629);
or U11479 (N_11479,N_9161,N_6180);
nor U11480 (N_11480,N_8208,N_6955);
or U11481 (N_11481,N_7214,N_6548);
nor U11482 (N_11482,N_6214,N_9544);
and U11483 (N_11483,N_8051,N_9774);
or U11484 (N_11484,N_9171,N_5163);
and U11485 (N_11485,N_5866,N_8290);
nor U11486 (N_11486,N_9114,N_7699);
and U11487 (N_11487,N_8927,N_6415);
and U11488 (N_11488,N_7272,N_8994);
nand U11489 (N_11489,N_9218,N_7068);
or U11490 (N_11490,N_7059,N_5489);
nand U11491 (N_11491,N_9572,N_5632);
xnor U11492 (N_11492,N_5674,N_6252);
and U11493 (N_11493,N_7830,N_5734);
nand U11494 (N_11494,N_5268,N_6165);
xor U11495 (N_11495,N_9592,N_7268);
nand U11496 (N_11496,N_6551,N_8633);
or U11497 (N_11497,N_6271,N_7663);
or U11498 (N_11498,N_6755,N_6375);
and U11499 (N_11499,N_7867,N_7861);
nor U11500 (N_11500,N_5127,N_8752);
or U11501 (N_11501,N_7145,N_8950);
nand U11502 (N_11502,N_8711,N_9896);
nand U11503 (N_11503,N_7846,N_8100);
xnor U11504 (N_11504,N_8913,N_8155);
nor U11505 (N_11505,N_7091,N_8240);
nor U11506 (N_11506,N_5488,N_5010);
nand U11507 (N_11507,N_5701,N_9029);
or U11508 (N_11508,N_7834,N_6549);
and U11509 (N_11509,N_6872,N_8298);
nor U11510 (N_11510,N_9605,N_7603);
and U11511 (N_11511,N_6492,N_9422);
or U11512 (N_11512,N_7056,N_8368);
nor U11513 (N_11513,N_5883,N_6297);
xor U11514 (N_11514,N_8457,N_6267);
or U11515 (N_11515,N_7736,N_6715);
nor U11516 (N_11516,N_9091,N_6711);
or U11517 (N_11517,N_8057,N_9042);
xor U11518 (N_11518,N_7527,N_7396);
or U11519 (N_11519,N_7574,N_8095);
and U11520 (N_11520,N_8740,N_5881);
nor U11521 (N_11521,N_5763,N_6394);
nand U11522 (N_11522,N_5496,N_6998);
nor U11523 (N_11523,N_6089,N_7207);
and U11524 (N_11524,N_5756,N_6570);
or U11525 (N_11525,N_6437,N_9949);
or U11526 (N_11526,N_9640,N_6074);
or U11527 (N_11527,N_9647,N_9147);
xnor U11528 (N_11528,N_9548,N_5993);
nand U11529 (N_11529,N_9353,N_7499);
or U11530 (N_11530,N_6432,N_8999);
or U11531 (N_11531,N_5052,N_7977);
or U11532 (N_11532,N_9262,N_7478);
nand U11533 (N_11533,N_6985,N_9252);
or U11534 (N_11534,N_7203,N_5914);
or U11535 (N_11535,N_7493,N_6743);
nor U11536 (N_11536,N_8257,N_7597);
or U11537 (N_11537,N_9809,N_9376);
nand U11538 (N_11538,N_8235,N_6283);
and U11539 (N_11539,N_8271,N_7264);
nand U11540 (N_11540,N_9076,N_7999);
or U11541 (N_11541,N_5968,N_6395);
nor U11542 (N_11542,N_5025,N_6703);
nor U11543 (N_11543,N_7668,N_9795);
or U11544 (N_11544,N_9316,N_9084);
nand U11545 (N_11545,N_7730,N_6897);
or U11546 (N_11546,N_9688,N_6095);
or U11547 (N_11547,N_5055,N_6199);
nand U11548 (N_11548,N_5930,N_5050);
nand U11549 (N_11549,N_8171,N_9119);
and U11550 (N_11550,N_6843,N_6263);
nor U11551 (N_11551,N_5397,N_7498);
nand U11552 (N_11552,N_8008,N_7787);
and U11553 (N_11553,N_5162,N_5501);
or U11554 (N_11554,N_6868,N_7344);
nand U11555 (N_11555,N_6969,N_7876);
or U11556 (N_11556,N_9403,N_7821);
and U11557 (N_11557,N_8898,N_9793);
xnor U11558 (N_11558,N_9750,N_5913);
nand U11559 (N_11559,N_7959,N_7874);
or U11560 (N_11560,N_5647,N_7737);
nand U11561 (N_11561,N_7316,N_7180);
xnor U11562 (N_11562,N_5782,N_6154);
nand U11563 (N_11563,N_8375,N_7534);
and U11564 (N_11564,N_8400,N_6009);
or U11565 (N_11565,N_6714,N_8622);
nand U11566 (N_11566,N_7710,N_7682);
or U11567 (N_11567,N_5586,N_8377);
nor U11568 (N_11568,N_8397,N_8616);
or U11569 (N_11569,N_8200,N_8459);
nor U11570 (N_11570,N_5819,N_5085);
nand U11571 (N_11571,N_7199,N_6486);
nand U11572 (N_11572,N_6509,N_6531);
or U11573 (N_11573,N_6027,N_5462);
nand U11574 (N_11574,N_7866,N_8516);
and U11575 (N_11575,N_6328,N_6238);
nor U11576 (N_11576,N_8629,N_5246);
nor U11577 (N_11577,N_8026,N_9869);
nor U11578 (N_11578,N_5444,N_5775);
or U11579 (N_11579,N_8489,N_7747);
or U11580 (N_11580,N_6137,N_7870);
nor U11581 (N_11581,N_6848,N_8665);
and U11582 (N_11582,N_6750,N_5498);
nor U11583 (N_11583,N_9710,N_7873);
nand U11584 (N_11584,N_9887,N_6685);
and U11585 (N_11585,N_7847,N_6578);
nor U11586 (N_11586,N_5203,N_9379);
or U11587 (N_11587,N_8079,N_7243);
or U11588 (N_11588,N_9396,N_9910);
nand U11589 (N_11589,N_9767,N_8742);
and U11590 (N_11590,N_5853,N_7561);
or U11591 (N_11591,N_6307,N_8907);
or U11592 (N_11592,N_9438,N_8632);
and U11593 (N_11593,N_6887,N_7192);
nor U11594 (N_11594,N_6237,N_8939);
nand U11595 (N_11595,N_9636,N_5080);
nand U11596 (N_11596,N_8173,N_7697);
nand U11597 (N_11597,N_9608,N_8126);
and U11598 (N_11598,N_7538,N_5815);
and U11599 (N_11599,N_8846,N_6521);
nand U11600 (N_11600,N_8869,N_5588);
nor U11601 (N_11601,N_6098,N_8667);
nor U11602 (N_11602,N_7387,N_8993);
and U11603 (N_11603,N_9758,N_7653);
nor U11604 (N_11604,N_5107,N_8954);
or U11605 (N_11605,N_5766,N_8584);
nand U11606 (N_11606,N_8380,N_7559);
or U11607 (N_11607,N_8055,N_6354);
or U11608 (N_11608,N_6864,N_8278);
nor U11609 (N_11609,N_8920,N_9919);
and U11610 (N_11610,N_6836,N_6301);
or U11611 (N_11611,N_7637,N_7453);
or U11612 (N_11612,N_7769,N_9373);
nand U11613 (N_11613,N_8895,N_9290);
or U11614 (N_11614,N_7491,N_6787);
and U11615 (N_11615,N_7923,N_6001);
nand U11616 (N_11616,N_9234,N_7798);
or U11617 (N_11617,N_6771,N_8680);
or U11618 (N_11618,N_9875,N_7275);
or U11619 (N_11619,N_6038,N_6725);
and U11620 (N_11620,N_9102,N_9098);
nor U11621 (N_11621,N_7671,N_5217);
nand U11622 (N_11622,N_9382,N_9395);
and U11623 (N_11623,N_7129,N_7987);
nand U11624 (N_11624,N_7044,N_6793);
nor U11625 (N_11625,N_8104,N_9418);
nand U11626 (N_11626,N_6502,N_9714);
nor U11627 (N_11627,N_8782,N_5787);
nand U11628 (N_11628,N_5275,N_5265);
or U11629 (N_11629,N_9272,N_8065);
nand U11630 (N_11630,N_7739,N_8258);
or U11631 (N_11631,N_6069,N_6988);
nor U11632 (N_11632,N_6717,N_6083);
nor U11633 (N_11633,N_8184,N_9017);
or U11634 (N_11634,N_9573,N_7530);
xnor U11635 (N_11635,N_7577,N_7390);
nor U11636 (N_11636,N_5174,N_5664);
nor U11637 (N_11637,N_6390,N_6223);
xor U11638 (N_11638,N_7594,N_9913);
nor U11639 (N_11639,N_5816,N_9739);
nor U11640 (N_11640,N_8510,N_8960);
nor U11641 (N_11641,N_8275,N_7288);
nor U11642 (N_11642,N_7931,N_9923);
or U11643 (N_11643,N_7273,N_9410);
or U11644 (N_11644,N_6202,N_6184);
and U11645 (N_11645,N_7425,N_6348);
and U11646 (N_11646,N_8120,N_7840);
nand U11647 (N_11647,N_5194,N_6823);
and U11648 (N_11648,N_6968,N_5448);
and U11649 (N_11649,N_9770,N_9437);
nand U11650 (N_11650,N_9079,N_9334);
nor U11651 (N_11651,N_7598,N_5707);
nand U11652 (N_11652,N_6596,N_7510);
or U11653 (N_11653,N_8774,N_6871);
nor U11654 (N_11654,N_5326,N_8292);
nor U11655 (N_11655,N_7173,N_9521);
nor U11656 (N_11656,N_8830,N_8648);
or U11657 (N_11657,N_5521,N_8535);
xnor U11658 (N_11658,N_9273,N_9420);
or U11659 (N_11659,N_6980,N_8005);
or U11660 (N_11660,N_8438,N_6169);
or U11661 (N_11661,N_5611,N_7483);
or U11662 (N_11662,N_9271,N_7031);
and U11663 (N_11663,N_7842,N_5537);
or U11664 (N_11664,N_9441,N_5684);
nor U11665 (N_11665,N_7766,N_9134);
and U11666 (N_11666,N_8339,N_8299);
and U11667 (N_11667,N_8795,N_8385);
nand U11668 (N_11668,N_8469,N_8636);
and U11669 (N_11669,N_8335,N_5757);
nand U11670 (N_11670,N_7835,N_7916);
and U11671 (N_11671,N_7054,N_9753);
xor U11672 (N_11672,N_8403,N_8772);
nand U11673 (N_11673,N_6298,N_9429);
or U11674 (N_11674,N_5545,N_9892);
and U11675 (N_11675,N_7123,N_9911);
and U11676 (N_11676,N_6642,N_8793);
or U11677 (N_11677,N_5654,N_6691);
nand U11678 (N_11678,N_9518,N_5257);
and U11679 (N_11679,N_6444,N_9664);
nand U11680 (N_11680,N_9007,N_6281);
nand U11681 (N_11681,N_9052,N_9348);
and U11682 (N_11682,N_5770,N_9406);
nor U11683 (N_11683,N_6782,N_8419);
nand U11684 (N_11684,N_9666,N_5956);
or U11685 (N_11685,N_5135,N_5293);
nor U11686 (N_11686,N_7814,N_7105);
nand U11687 (N_11687,N_8179,N_9858);
xor U11688 (N_11688,N_9835,N_8536);
nor U11689 (N_11689,N_7761,N_7800);
xor U11690 (N_11690,N_8968,N_9959);
nand U11691 (N_11691,N_7558,N_7447);
nand U11692 (N_11692,N_7127,N_5161);
nor U11693 (N_11693,N_7551,N_7178);
nor U11694 (N_11694,N_9763,N_7458);
and U11695 (N_11695,N_8369,N_8237);
nand U11696 (N_11696,N_8072,N_5745);
nand U11697 (N_11697,N_9489,N_8096);
or U11698 (N_11698,N_6062,N_5511);
or U11699 (N_11699,N_9995,N_8753);
nor U11700 (N_11700,N_5835,N_9571);
nor U11701 (N_11701,N_6049,N_6863);
nand U11702 (N_11702,N_6666,N_8685);
nand U11703 (N_11703,N_5446,N_8935);
or U11704 (N_11704,N_7466,N_8966);
or U11705 (N_11705,N_8860,N_8973);
nand U11706 (N_11706,N_5058,N_9012);
nand U11707 (N_11707,N_5518,N_7589);
nor U11708 (N_11708,N_9074,N_6081);
nor U11709 (N_11709,N_6797,N_6689);
or U11710 (N_11710,N_9931,N_7080);
and U11711 (N_11711,N_9839,N_8823);
nand U11712 (N_11712,N_9922,N_5227);
or U11713 (N_11713,N_7337,N_9994);
xor U11714 (N_11714,N_6961,N_5919);
nor U11715 (N_11715,N_9100,N_7282);
nor U11716 (N_11716,N_8831,N_8705);
and U11717 (N_11717,N_7351,N_5490);
nand U11718 (N_11718,N_8614,N_5356);
nand U11719 (N_11719,N_5426,N_7758);
nand U11720 (N_11720,N_7121,N_5601);
nor U11721 (N_11721,N_6500,N_5618);
nand U11722 (N_11722,N_9107,N_9138);
nand U11723 (N_11723,N_9988,N_7278);
and U11724 (N_11724,N_5285,N_9495);
nand U11725 (N_11725,N_8180,N_6428);
nand U11726 (N_11726,N_8448,N_8745);
and U11727 (N_11727,N_9105,N_9616);
or U11728 (N_11728,N_8780,N_5360);
and U11729 (N_11729,N_7392,N_6756);
or U11730 (N_11730,N_7460,N_7191);
nor U11731 (N_11731,N_7136,N_8794);
nand U11732 (N_11732,N_8253,N_6874);
nand U11733 (N_11733,N_6647,N_7300);
nor U11734 (N_11734,N_9095,N_7634);
nor U11735 (N_11735,N_7176,N_7209);
and U11736 (N_11736,N_9018,N_9500);
nand U11737 (N_11737,N_6668,N_7841);
and U11738 (N_11738,N_5879,N_7187);
nor U11739 (N_11739,N_7114,N_6277);
or U11740 (N_11740,N_6504,N_9366);
or U11741 (N_11741,N_8615,N_9254);
and U11742 (N_11742,N_9554,N_9814);
nand U11743 (N_11743,N_8893,N_9606);
nand U11744 (N_11744,N_9886,N_5981);
or U11745 (N_11745,N_8707,N_8347);
nor U11746 (N_11746,N_7752,N_8227);
nor U11747 (N_11747,N_8554,N_8719);
nor U11748 (N_11748,N_9641,N_6795);
nand U11749 (N_11749,N_5658,N_9110);
nor U11750 (N_11750,N_7413,N_8844);
nand U11751 (N_11751,N_5158,N_6345);
nand U11752 (N_11752,N_7939,N_9491);
or U11753 (N_11753,N_6945,N_6525);
nand U11754 (N_11754,N_5095,N_9198);
and U11755 (N_11755,N_7687,N_5871);
nor U11756 (N_11756,N_5369,N_8112);
and U11757 (N_11757,N_5032,N_7683);
or U11758 (N_11758,N_5791,N_6469);
and U11759 (N_11759,N_5936,N_6321);
nand U11760 (N_11760,N_9623,N_8923);
nor U11761 (N_11761,N_8500,N_8003);
nor U11762 (N_11762,N_5089,N_9700);
nor U11763 (N_11763,N_6639,N_7285);
nor U11764 (N_11764,N_9542,N_6413);
and U11765 (N_11765,N_7063,N_5769);
and U11766 (N_11766,N_9260,N_8757);
and U11767 (N_11767,N_6305,N_6545);
and U11768 (N_11768,N_9345,N_5450);
xnor U11769 (N_11769,N_9222,N_8798);
or U11770 (N_11770,N_6528,N_9282);
nor U11771 (N_11771,N_7356,N_8998);
and U11772 (N_11772,N_8303,N_9662);
nand U11773 (N_11773,N_6456,N_7778);
and U11774 (N_11774,N_5200,N_6391);
nand U11775 (N_11775,N_6087,N_9822);
nor U11776 (N_11776,N_7560,N_9792);
nor U11777 (N_11777,N_9250,N_6319);
nor U11778 (N_11778,N_5299,N_9899);
xnor U11779 (N_11779,N_8133,N_9448);
nand U11780 (N_11780,N_6737,N_8068);
nor U11781 (N_11781,N_7185,N_8518);
nor U11782 (N_11782,N_7292,N_8756);
or U11783 (N_11783,N_9169,N_6599);
and U11784 (N_11784,N_9200,N_7119);
nand U11785 (N_11785,N_9036,N_9050);
or U11786 (N_11786,N_6631,N_8702);
or U11787 (N_11787,N_6999,N_7744);
nor U11788 (N_11788,N_6997,N_5482);
nand U11789 (N_11789,N_5949,N_7995);
and U11790 (N_11790,N_8746,N_8668);
and U11791 (N_11791,N_9099,N_9125);
or U11792 (N_11792,N_7027,N_6505);
and U11793 (N_11793,N_7793,N_5940);
nand U11794 (N_11794,N_8324,N_5384);
or U11795 (N_11795,N_6873,N_8080);
nor U11796 (N_11796,N_8394,N_5405);
and U11797 (N_11797,N_6310,N_8641);
nor U11798 (N_11798,N_6801,N_5603);
or U11799 (N_11799,N_6240,N_6052);
nand U11800 (N_11800,N_8111,N_8972);
nand U11801 (N_11801,N_8156,N_7010);
and U11802 (N_11802,N_8841,N_8345);
nor U11803 (N_11803,N_6619,N_6053);
nor U11804 (N_11804,N_9297,N_7988);
or U11805 (N_11805,N_6602,N_6420);
or U11806 (N_11806,N_6460,N_5445);
nand U11807 (N_11807,N_8675,N_8311);
and U11808 (N_11808,N_5671,N_8355);
nand U11809 (N_11809,N_5338,N_9466);
or U11810 (N_11810,N_7072,N_6332);
nor U11811 (N_11811,N_8904,N_7124);
and U11812 (N_11812,N_5928,N_6830);
nand U11813 (N_11813,N_9890,N_6924);
or U11814 (N_11814,N_8804,N_8110);
nand U11815 (N_11815,N_8228,N_5715);
nand U11816 (N_11816,N_6747,N_7573);
nor U11817 (N_11817,N_9658,N_5109);
or U11818 (N_11818,N_5305,N_8349);
nand U11819 (N_11819,N_7716,N_5810);
and U11820 (N_11820,N_9586,N_8811);
nand U11821 (N_11821,N_6008,N_8114);
or U11822 (N_11822,N_5465,N_7418);
or U11823 (N_11823,N_5755,N_7664);
and U11824 (N_11824,N_7750,N_7160);
nor U11825 (N_11825,N_8399,N_9904);
and U11826 (N_11826,N_8658,N_5572);
nand U11827 (N_11827,N_7775,N_7240);
or U11828 (N_11828,N_8788,N_9315);
and U11829 (N_11829,N_9941,N_5012);
or U11830 (N_11830,N_8041,N_9117);
or U11831 (N_11831,N_9850,N_9191);
nor U11832 (N_11832,N_6334,N_7294);
nor U11833 (N_11833,N_7933,N_5500);
nor U11834 (N_11834,N_5139,N_9694);
and U11835 (N_11835,N_5543,N_5023);
or U11836 (N_11836,N_7605,N_9286);
nor U11837 (N_11837,N_9080,N_5567);
and U11838 (N_11838,N_5026,N_9023);
nand U11839 (N_11839,N_7552,N_8326);
or U11840 (N_11840,N_5887,N_9801);
nand U11841 (N_11841,N_6114,N_8529);
nand U11842 (N_11842,N_5615,N_7303);
and U11843 (N_11843,N_7666,N_9543);
nand U11844 (N_11844,N_5301,N_6810);
xnor U11845 (N_11845,N_9130,N_6716);
nand U11846 (N_11846,N_6170,N_9368);
or U11847 (N_11847,N_5540,N_7936);
and U11848 (N_11848,N_7332,N_7896);
or U11849 (N_11849,N_5860,N_6624);
nor U11850 (N_11850,N_5047,N_5459);
nand U11851 (N_11851,N_7770,N_6587);
and U11852 (N_11852,N_9600,N_6244);
nor U11853 (N_11853,N_7388,N_9619);
or U11854 (N_11854,N_9414,N_9168);
and U11855 (N_11855,N_9905,N_5765);
or U11856 (N_11856,N_6011,N_7586);
nor U11857 (N_11857,N_8158,N_8097);
nand U11858 (N_11858,N_6857,N_5056);
and U11859 (N_11859,N_5653,N_8036);
nor U11860 (N_11860,N_9813,N_7693);
and U11861 (N_11861,N_7074,N_8559);
nand U11862 (N_11862,N_9439,N_7569);
nor U11863 (N_11863,N_9961,N_5145);
nand U11864 (N_11864,N_6115,N_8424);
or U11865 (N_11865,N_8751,N_6722);
nand U11866 (N_11866,N_6020,N_5436);
nand U11867 (N_11867,N_6030,N_8020);
nand U11868 (N_11868,N_5994,N_7428);
or U11869 (N_11869,N_6512,N_9449);
nand U11870 (N_11870,N_8185,N_5477);
or U11871 (N_11871,N_8824,N_7831);
and U11872 (N_11872,N_9274,N_5826);
or U11873 (N_11873,N_6617,N_7405);
xor U11874 (N_11874,N_7632,N_9182);
nor U11875 (N_11875,N_5370,N_9223);
nand U11876 (N_11876,N_5864,N_5751);
nor U11877 (N_11877,N_5641,N_7924);
or U11878 (N_11878,N_6484,N_5240);
nand U11879 (N_11879,N_6888,N_6440);
and U11880 (N_11880,N_7302,N_6033);
nor U11881 (N_11881,N_6904,N_9402);
xor U11882 (N_11882,N_8452,N_6732);
nor U11883 (N_11883,N_6124,N_9929);
xor U11884 (N_11884,N_8329,N_8412);
nand U11885 (N_11885,N_8866,N_5367);
or U11886 (N_11886,N_9265,N_9746);
or U11887 (N_11887,N_5331,N_5735);
nor U11888 (N_11888,N_9391,N_8277);
nand U11889 (N_11889,N_8314,N_6934);
nor U11890 (N_11890,N_7444,N_6901);
nor U11891 (N_11891,N_5189,N_9849);
nor U11892 (N_11892,N_5298,N_5719);
nand U11893 (N_11893,N_5963,N_9476);
xnor U11894 (N_11894,N_8229,N_8595);
nor U11895 (N_11895,N_9546,N_6786);
and U11896 (N_11896,N_6387,N_8323);
or U11897 (N_11897,N_6150,N_5351);
and U11898 (N_11898,N_6667,N_9383);
and U11899 (N_11899,N_8894,N_7260);
nand U11900 (N_11900,N_8945,N_6688);
and U11901 (N_11901,N_9932,N_6921);
or U11902 (N_11902,N_5640,N_5857);
xor U11903 (N_11903,N_6523,N_7623);
and U11904 (N_11904,N_5375,N_6595);
nand U11905 (N_11905,N_5374,N_8653);
nand U11906 (N_11906,N_5677,N_9484);
and U11907 (N_11907,N_9908,N_6884);
and U11908 (N_11908,N_7468,N_7153);
nor U11909 (N_11909,N_5346,N_6723);
xor U11910 (N_11910,N_5530,N_6603);
nor U11911 (N_11911,N_8161,N_5485);
nand U11912 (N_11912,N_9442,N_8118);
nand U11913 (N_11913,N_8868,N_6537);
and U11914 (N_11914,N_5415,N_7504);
or U11915 (N_11915,N_6389,N_7858);
nor U11916 (N_11916,N_6373,N_5593);
nand U11917 (N_11917,N_8050,N_7222);
and U11918 (N_11918,N_6876,N_7772);
and U11919 (N_11919,N_7496,N_9178);
or U11920 (N_11920,N_9040,N_5699);
and U11921 (N_11921,N_6190,N_5226);
and U11922 (N_11922,N_5555,N_6085);
nor U11923 (N_11923,N_7433,N_6783);
nor U11924 (N_11924,N_5333,N_8194);
and U11925 (N_11925,N_5454,N_7832);
or U11926 (N_11926,N_7201,N_7952);
nand U11927 (N_11927,N_7097,N_7514);
nor U11928 (N_11928,N_6099,N_8255);
or U11929 (N_11929,N_9567,N_7427);
nand U11930 (N_11930,N_7025,N_7200);
nand U11931 (N_11931,N_6129,N_5962);
and U11932 (N_11932,N_5035,N_6355);
xnor U11933 (N_11933,N_9067,N_6829);
and U11934 (N_11934,N_9957,N_7098);
or U11935 (N_11935,N_6376,N_9691);
xor U11936 (N_11936,N_9556,N_8217);
and U11937 (N_11937,N_8799,N_6649);
or U11938 (N_11938,N_6803,N_6019);
nand U11939 (N_11939,N_6181,N_5069);
nor U11940 (N_11940,N_7208,N_6144);
or U11941 (N_11941,N_6605,N_7283);
or U11942 (N_11942,N_5858,N_9292);
and U11943 (N_11943,N_7917,N_5878);
nand U11944 (N_11944,N_9189,N_9536);
or U11945 (N_11945,N_7718,N_7141);
or U11946 (N_11946,N_6106,N_7691);
nand U11947 (N_11947,N_5984,N_5942);
or U11948 (N_11948,N_9180,N_7893);
and U11949 (N_11949,N_6907,N_5327);
nand U11950 (N_11950,N_6707,N_7575);
or U11951 (N_11951,N_7940,N_6837);
nor U11952 (N_11952,N_5694,N_7367);
nand U11953 (N_11953,N_7443,N_8887);
or U11954 (N_11954,N_5633,N_7195);
nor U11955 (N_11955,N_6987,N_8131);
and U11956 (N_11956,N_8059,N_9241);
nand U11957 (N_11957,N_8132,N_5481);
nand U11958 (N_11958,N_9744,N_8365);
and U11959 (N_11959,N_6111,N_5828);
and U11960 (N_11960,N_9317,N_8911);
and U11961 (N_11961,N_8491,N_5869);
or U11962 (N_11962,N_5612,N_7516);
nor U11963 (N_11963,N_7946,N_6286);
nor U11964 (N_11964,N_6966,N_6859);
nor U11965 (N_11965,N_5777,N_8302);
and U11966 (N_11966,N_7365,N_8094);
or U11967 (N_11967,N_6586,N_9359);
nor U11968 (N_11968,N_8093,N_5033);
nor U11969 (N_11969,N_6883,N_5550);
nand U11970 (N_11970,N_5337,N_6754);
or U11971 (N_11971,N_9127,N_8980);
nand U11972 (N_11972,N_6635,N_5544);
nand U11973 (N_11973,N_8563,N_8596);
nor U11974 (N_11974,N_7903,N_6585);
or U11975 (N_11975,N_8183,N_8123);
or U11976 (N_11976,N_7484,N_5812);
or U11977 (N_11977,N_5977,N_9296);
nand U11978 (N_11978,N_6695,N_7704);
nor U11979 (N_11979,N_9144,N_7955);
or U11980 (N_11980,N_8775,N_9806);
nor U11981 (N_11981,N_7911,N_7547);
nor U11982 (N_11982,N_8221,N_8631);
nor U11983 (N_11983,N_6900,N_9914);
nor U11984 (N_11984,N_6268,N_5675);
or U11985 (N_11985,N_9891,N_8880);
or U11986 (N_11986,N_6023,N_8261);
nand U11987 (N_11987,N_9788,N_5431);
nor U11988 (N_11988,N_7130,N_9230);
or U11989 (N_11989,N_7811,N_6751);
nor U11990 (N_11990,N_9078,N_8607);
or U11991 (N_11991,N_8726,N_6029);
nor U11992 (N_11992,N_6832,N_7844);
nor U11993 (N_11993,N_7089,N_8053);
and U11994 (N_11994,N_8652,N_7550);
and U11995 (N_11995,N_5383,N_8744);
nand U11996 (N_11996,N_5071,N_8444);
nor U11997 (N_11997,N_6657,N_9560);
and U11998 (N_11998,N_9496,N_9001);
nor U11999 (N_11999,N_5923,N_9385);
nor U12000 (N_12000,N_5376,N_6882);
and U12001 (N_12001,N_8121,N_8926);
or U12002 (N_12002,N_5133,N_9498);
or U12003 (N_12003,N_5778,N_6303);
nand U12004 (N_12004,N_8296,N_6633);
xnor U12005 (N_12005,N_7251,N_9725);
nor U12006 (N_12006,N_6834,N_5169);
nor U12007 (N_12007,N_5324,N_5649);
nor U12008 (N_12008,N_9145,N_5460);
or U12009 (N_12009,N_9824,N_6510);
and U12010 (N_12010,N_9375,N_5099);
nor U12011 (N_12011,N_6186,N_7851);
nand U12012 (N_12012,N_8447,N_6681);
and U12013 (N_12013,N_8175,N_5083);
nor U12014 (N_12014,N_8682,N_5581);
nand U12015 (N_12015,N_8077,N_7553);
nor U12016 (N_12016,N_7467,N_6179);
nand U12017 (N_12017,N_9175,N_8747);
and U12018 (N_12018,N_7734,N_5345);
nor U12019 (N_12019,N_8259,N_7662);
or U12020 (N_12020,N_6032,N_7155);
or U12021 (N_12021,N_6410,N_6625);
nand U12022 (N_12022,N_9003,N_5602);
nand U12023 (N_12023,N_5696,N_7871);
nand U12024 (N_12024,N_9761,N_8989);
nand U12025 (N_12025,N_5638,N_8021);
nor U12026 (N_12026,N_5307,N_5224);
nand U12027 (N_12027,N_5118,N_7245);
nor U12028 (N_12028,N_6250,N_9823);
nand U12029 (N_12029,N_5209,N_5480);
or U12030 (N_12030,N_5833,N_9987);
nand U12031 (N_12031,N_6220,N_8699);
nand U12032 (N_12032,N_7112,N_6679);
or U12033 (N_12033,N_8952,N_9883);
xor U12034 (N_12034,N_9673,N_9264);
and U12035 (N_12035,N_5036,N_8807);
nand U12036 (N_12036,N_9502,N_9137);
or U12037 (N_12037,N_9245,N_7617);
or U12038 (N_12038,N_8540,N_7804);
nor U12039 (N_12039,N_5372,N_8694);
and U12040 (N_12040,N_6109,N_5206);
or U12041 (N_12041,N_7269,N_6426);
nor U12042 (N_12042,N_7969,N_7441);
and U12043 (N_12043,N_8384,N_5683);
and U12044 (N_12044,N_6575,N_8858);
nor U12045 (N_12045,N_8415,N_9613);
nor U12046 (N_12046,N_7309,N_6671);
or U12047 (N_12047,N_5187,N_8232);
nand U12048 (N_12048,N_9156,N_9974);
and U12049 (N_12049,N_8197,N_8109);
and U12050 (N_12050,N_8515,N_6350);
nor U12051 (N_12051,N_9275,N_8625);
or U12052 (N_12052,N_9212,N_8709);
nor U12053 (N_12053,N_6343,N_7731);
or U12054 (N_12054,N_9355,N_9221);
and U12055 (N_12055,N_7984,N_6340);
and U12056 (N_12056,N_8388,N_8890);
nor U12057 (N_12057,N_8413,N_8370);
nor U12058 (N_12058,N_7799,N_8840);
nand U12059 (N_12059,N_7953,N_8501);
or U12060 (N_12060,N_9771,N_8579);
nor U12061 (N_12061,N_5886,N_8230);
nor U12062 (N_12062,N_8182,N_5882);
and U12063 (N_12063,N_9864,N_8524);
or U12064 (N_12064,N_7262,N_5662);
nand U12065 (N_12065,N_6982,N_8243);
or U12066 (N_12066,N_6673,N_7568);
nand U12067 (N_12067,N_5578,N_6132);
or U12068 (N_12068,N_6025,N_8829);
nor U12069 (N_12069,N_8164,N_9086);
and U12070 (N_12070,N_5646,N_6789);
nand U12071 (N_12071,N_9136,N_7554);
and U12072 (N_12072,N_8815,N_9313);
nand U12073 (N_12073,N_9738,N_8274);
or U12074 (N_12074,N_7241,N_8196);
or U12075 (N_12075,N_6449,N_6127);
nand U12076 (N_12076,N_8332,N_7563);
or U12077 (N_12077,N_9434,N_8733);
and U12078 (N_12078,N_8108,N_5090);
nand U12079 (N_12079,N_5764,N_7606);
or U12080 (N_12080,N_9831,N_6892);
nor U12081 (N_12081,N_6495,N_8214);
and U12082 (N_12082,N_6090,N_7347);
nor U12083 (N_12083,N_8766,N_8803);
nor U12084 (N_12084,N_9777,N_8030);
or U12085 (N_12085,N_9790,N_7227);
nand U12086 (N_12086,N_9780,N_6458);
or U12087 (N_12087,N_6778,N_7117);
or U12088 (N_12088,N_8833,N_7967);
or U12089 (N_12089,N_9346,N_5669);
or U12090 (N_12090,N_5253,N_8856);
or U12091 (N_12091,N_9537,N_9332);
or U12092 (N_12092,N_9678,N_9063);
nor U12093 (N_12093,N_9380,N_6296);
and U12094 (N_12094,N_6329,N_5455);
or U12095 (N_12095,N_8450,N_6113);
and U12096 (N_12096,N_8805,N_6538);
and U12097 (N_12097,N_6738,N_8498);
or U12098 (N_12098,N_9829,N_9328);
or U12099 (N_12099,N_6110,N_7636);
nand U12100 (N_12100,N_9364,N_6497);
nor U12101 (N_12101,N_8357,N_6362);
nand U12102 (N_12102,N_8364,N_7350);
nor U12103 (N_12103,N_6950,N_9888);
xnor U12104 (N_12104,N_9143,N_7293);
and U12105 (N_12105,N_5201,N_9973);
nand U12106 (N_12106,N_8635,N_7034);
or U12107 (N_12107,N_7745,N_5652);
and U12108 (N_12108,N_7474,N_9347);
or U12109 (N_12109,N_8542,N_8948);
and U12110 (N_12110,N_9773,N_7792);
nand U12111 (N_12111,N_9424,N_9843);
or U12112 (N_12112,N_9527,N_5657);
and U12113 (N_12113,N_7751,N_6174);
and U12114 (N_12114,N_7225,N_7607);
or U12115 (N_12115,N_7612,N_6134);
and U12116 (N_12116,N_9152,N_8619);
nand U12117 (N_12117,N_7408,N_5153);
or U12118 (N_12118,N_6951,N_7808);
and U12119 (N_12119,N_8580,N_6698);
nand U12120 (N_12120,N_8881,N_8492);
nand U12121 (N_12121,N_6767,N_5844);
nand U12122 (N_12122,N_7991,N_9051);
or U12123 (N_12123,N_9059,N_7042);
nand U12124 (N_12124,N_6414,N_6616);
and U12125 (N_12125,N_7943,N_8177);
and U12126 (N_12126,N_9416,N_6398);
nor U12127 (N_12127,N_9025,N_8304);
nor U12128 (N_12128,N_8862,N_7944);
and U12129 (N_12129,N_5515,N_7348);
nand U12130 (N_12130,N_6807,N_6634);
and U12131 (N_12131,N_7622,N_5235);
nor U12132 (N_12132,N_7749,N_6568);
nand U12133 (N_12133,N_9517,N_9716);
nand U12134 (N_12134,N_7557,N_6327);
nand U12135 (N_12135,N_8147,N_6036);
and U12136 (N_12136,N_8286,N_6122);
or U12137 (N_12137,N_5325,N_5957);
and U12138 (N_12138,N_6675,N_5159);
or U12139 (N_12139,N_6840,N_5008);
nor U12140 (N_12140,N_5754,N_6792);
and U12141 (N_12141,N_9602,N_8067);
nand U12142 (N_12142,N_7500,N_7143);
or U12143 (N_12143,N_7297,N_8509);
xor U12144 (N_12144,N_8737,N_5435);
and U12145 (N_12145,N_5739,N_7755);
nor U12146 (N_12146,N_8453,N_7986);
nor U12147 (N_12147,N_7738,N_5742);
or U12148 (N_12148,N_7604,N_7689);
nand U12149 (N_12149,N_8178,N_8678);
or U12150 (N_12150,N_5592,N_7190);
nor U12151 (N_12151,N_5740,N_6047);
nand U12152 (N_12152,N_7152,N_6013);
nand U12153 (N_12153,N_8755,N_9233);
nand U12154 (N_12154,N_6734,N_9370);
and U12155 (N_12155,N_6056,N_9881);
nor U12156 (N_12156,N_6841,N_5122);
xor U12157 (N_12157,N_7047,N_6257);
nor U12158 (N_12158,N_5645,N_6269);
or U12159 (N_12159,N_5529,N_5896);
nor U12160 (N_12160,N_5483,N_8167);
or U12161 (N_12161,N_5261,N_7277);
nand U12162 (N_12162,N_5971,N_5809);
or U12163 (N_12163,N_6177,N_8289);
or U12164 (N_12164,N_7019,N_8981);
nor U12165 (N_12165,N_9920,N_7409);
or U12166 (N_12166,N_5534,N_9331);
nand U12167 (N_12167,N_9401,N_8857);
nor U12168 (N_12168,N_7438,N_5836);
or U12169 (N_12169,N_9020,N_8421);
and U12170 (N_12170,N_7963,N_8350);
and U12171 (N_12171,N_6116,N_6351);
or U12172 (N_12172,N_5328,N_9077);
and U12173 (N_12173,N_5359,N_6550);
nand U12174 (N_12174,N_8941,N_5354);
nor U12175 (N_12175,N_5711,N_7810);
or U12176 (N_12176,N_9954,N_6046);
and U12177 (N_12177,N_8526,N_9160);
or U12178 (N_12178,N_8454,N_6187);
nor U12179 (N_12179,N_6107,N_8897);
nand U12180 (N_12180,N_5241,N_8353);
or U12181 (N_12181,N_7361,N_8891);
nand U12182 (N_12182,N_8663,N_7526);
and U12183 (N_12183,N_5451,N_8724);
nand U12184 (N_12184,N_7812,N_5975);
nand U12185 (N_12185,N_9371,N_7587);
nand U12186 (N_12186,N_5698,N_9577);
or U12187 (N_12187,N_5851,N_7289);
nand U12188 (N_12188,N_9711,N_7131);
or U12189 (N_12189,N_9349,N_9081);
xor U12190 (N_12190,N_7629,N_5221);
nand U12191 (N_12191,N_8676,N_5820);
or U12192 (N_12192,N_8313,N_7463);
or U12193 (N_12193,N_9677,N_9861);
and U12194 (N_12194,N_7599,N_8427);
nand U12195 (N_12195,N_7883,N_9918);
or U12196 (N_12196,N_9568,N_9784);
or U12197 (N_12197,N_6210,N_6941);
nor U12198 (N_12198,N_5341,N_8481);
nor U12199 (N_12199,N_7652,N_6161);
nand U12200 (N_12200,N_6546,N_7624);
or U12201 (N_12201,N_8874,N_7090);
or U12202 (N_12202,N_5248,N_9190);
nor U12203 (N_12203,N_7336,N_8098);
nor U12204 (N_12204,N_9303,N_5904);
and U12205 (N_12205,N_9153,N_8943);
nor U12206 (N_12206,N_8691,N_8571);
nand U12207 (N_12207,N_6562,N_9455);
or U12208 (N_12208,N_9205,N_7402);
or U12209 (N_12209,N_5779,N_7334);
nand U12210 (N_12210,N_9513,N_5856);
nand U12211 (N_12211,N_8832,N_5996);
or U12212 (N_12212,N_7706,N_9800);
and U12213 (N_12213,N_9707,N_9601);
xnor U12214 (N_12214,N_6285,N_7030);
or U12215 (N_12215,N_8720,N_9538);
nor U12216 (N_12216,N_8288,N_8251);
and U12217 (N_12217,N_5606,N_5517);
nor U12218 (N_12218,N_5183,N_5350);
and U12219 (N_12219,N_8140,N_8918);
nand U12220 (N_12220,N_8462,N_9582);
nand U12221 (N_12221,N_9033,N_8416);
nor U12222 (N_12222,N_7743,N_6487);
or U12223 (N_12223,N_6235,N_8670);
nor U12224 (N_12224,N_8172,N_7845);
nand U12225 (N_12225,N_7723,N_9889);
nor U12226 (N_12226,N_7897,N_7434);
or U12227 (N_12227,N_6869,N_8378);
nor U12228 (N_12228,N_6078,N_5317);
or U12229 (N_12229,N_9384,N_7020);
nor U12230 (N_12230,N_6895,N_9797);
or U12231 (N_12231,N_7104,N_6995);
and U12232 (N_12232,N_5680,N_5553);
and U12233 (N_12233,N_8060,N_8395);
and U12234 (N_12234,N_8730,N_6361);
nand U12235 (N_12235,N_6335,N_9653);
nand U12236 (N_12236,N_8646,N_8023);
or U12237 (N_12237,N_7966,N_8901);
nor U12238 (N_12238,N_8825,N_9415);
or U12239 (N_12239,N_6769,N_8405);
or U12240 (N_12240,N_9238,N_7806);
nor U12241 (N_12241,N_7188,N_6232);
and U12242 (N_12242,N_5800,N_8922);
nand U12243 (N_12243,N_5195,N_9940);
or U12244 (N_12244,N_5062,N_7094);
or U12245 (N_12245,N_9731,N_9231);
or U12246 (N_12246,N_6693,N_5150);
or U12247 (N_12247,N_7071,N_8152);
nand U12248 (N_12248,N_8188,N_7932);
nor U12249 (N_12249,N_8613,N_9378);
nor U12250 (N_12250,N_6189,N_6644);
or U12251 (N_12251,N_7149,N_8934);
nor U12252 (N_12252,N_7454,N_6814);
nand U12253 (N_12253,N_6785,N_6866);
nor U12254 (N_12254,N_9533,N_7838);
nand U12255 (N_12255,N_5995,N_7993);
or U12256 (N_12256,N_9982,N_5897);
and U12257 (N_12257,N_5000,N_8997);
and U12258 (N_12258,N_6427,N_8280);
nand U12259 (N_12259,N_5823,N_9857);
nand U12260 (N_12260,N_9815,N_8674);
nor U12261 (N_12261,N_5484,N_6121);
or U12262 (N_12262,N_9475,N_7937);
and U12263 (N_12263,N_8264,N_5001);
xor U12264 (N_12264,N_9243,N_6678);
and U12265 (N_12265,N_7501,N_5473);
and U12266 (N_12266,N_5590,N_9530);
or U12267 (N_12267,N_7588,N_5306);
nor U12268 (N_12268,N_6431,N_6253);
and U12269 (N_12269,N_9976,N_6794);
nand U12270 (N_12270,N_8033,N_5072);
nand U12271 (N_12271,N_9300,N_5843);
nand U12272 (N_12272,N_7698,N_6971);
nand U12273 (N_12273,N_6359,N_6902);
nand U12274 (N_12274,N_8717,N_5723);
nor U12275 (N_12275,N_6131,N_5418);
and U12276 (N_12276,N_6979,N_5573);
and U12277 (N_12277,N_6664,N_5762);
nor U12278 (N_12278,N_5788,N_9528);
nor U12279 (N_12279,N_7024,N_9008);
nand U12280 (N_12280,N_5140,N_9505);
nand U12281 (N_12281,N_8822,N_9013);
nor U12282 (N_12282,N_5946,N_7620);
nor U12283 (N_12283,N_5478,N_5506);
or U12284 (N_12284,N_8012,N_7366);
and U12285 (N_12285,N_7645,N_8056);
nor U12286 (N_12286,N_9170,N_6682);
and U12287 (N_12287,N_7785,N_6775);
nor U12288 (N_12288,N_8256,N_5704);
or U12289 (N_12289,N_5264,N_5637);
or U12290 (N_12290,N_8134,N_7996);
and U12291 (N_12291,N_9321,N_7486);
nor U12292 (N_12292,N_6266,N_5114);
or U12293 (N_12293,N_9845,N_8659);
or U12294 (N_12294,N_5295,N_6216);
or U12295 (N_12295,N_6915,N_8865);
or U12296 (N_12296,N_7032,N_5428);
nor U12297 (N_12297,N_9547,N_6651);
nand U12298 (N_12298,N_8083,N_5733);
nand U12299 (N_12299,N_7929,N_9996);
nand U12300 (N_12300,N_9868,N_5725);
nand U12301 (N_12301,N_7641,N_7049);
and U12302 (N_12302,N_7791,N_5758);
or U12303 (N_12303,N_6064,N_8102);
or U12304 (N_12304,N_6858,N_9563);
nand U12305 (N_12305,N_7239,N_9421);
nand U12306 (N_12306,N_9314,N_9927);
nand U12307 (N_12307,N_8723,N_6665);
and U12308 (N_12308,N_6123,N_8201);
nand U12309 (N_12309,N_6316,N_7419);
nor U12310 (N_12310,N_5063,N_7229);
and U12311 (N_12311,N_8474,N_9146);
nand U12312 (N_12312,N_6278,N_6574);
and U12313 (N_12313,N_7509,N_5944);
or U12314 (N_12314,N_7281,N_5992);
or U12315 (N_12315,N_8267,N_5958);
or U12316 (N_12316,N_6212,N_9580);
or U12317 (N_12317,N_8561,N_7186);
nor U12318 (N_12318,N_8885,N_8764);
and U12319 (N_12319,N_7322,N_6119);
nand U12320 (N_12320,N_9176,N_9661);
nand U12321 (N_12321,N_5266,N_7372);
and U12322 (N_12322,N_6760,N_5320);
or U12323 (N_12323,N_8465,N_6365);
nor U12324 (N_12324,N_8696,N_6677);
or U12325 (N_12325,N_5575,N_7548);
nor U12326 (N_12326,N_9975,N_5149);
or U12327 (N_12327,N_8269,N_9837);
or U12328 (N_12328,N_6084,N_7549);
nand U12329 (N_12329,N_9734,N_6910);
nor U12330 (N_12330,N_9723,N_5296);
or U12331 (N_12331,N_7596,N_8643);
nand U12332 (N_12332,N_5439,N_5204);
xnor U12333 (N_12333,N_9760,N_5655);
and U12334 (N_12334,N_9197,N_7014);
and U12335 (N_12335,N_8205,N_8040);
or U12336 (N_12336,N_7621,N_6270);
nor U12337 (N_12337,N_9786,N_6534);
and U12338 (N_12338,N_6464,N_7248);
or U12339 (N_12339,N_5569,N_9874);
nand U12340 (N_12340,N_5466,N_7040);
nand U12341 (N_12341,N_8716,N_6558);
or U12342 (N_12342,N_8432,N_5218);
nand U12343 (N_12343,N_9741,N_6517);
and U12344 (N_12344,N_6218,N_7508);
and U12345 (N_12345,N_9524,N_5796);
and U12346 (N_12346,N_8417,N_5119);
nand U12347 (N_12347,N_6705,N_9242);
nor U12348 (N_12348,N_9335,N_6908);
nor U12349 (N_12349,N_5576,N_6418);
nand U12350 (N_12350,N_7779,N_8520);
nand U12351 (N_12351,N_7244,N_7015);
nor U12352 (N_12352,N_7970,N_9097);
nand U12353 (N_12353,N_8875,N_5148);
nand U12354 (N_12354,N_5223,N_7979);
nand U12355 (N_12355,N_8933,N_8422);
nor U12356 (N_12356,N_9985,N_6952);
or U12357 (N_12357,N_7638,N_5319);
nor U12358 (N_12358,N_6556,N_9549);
or U12359 (N_12359,N_8411,N_6392);
and U12360 (N_12360,N_8712,N_9075);
and U12361 (N_12361,N_7784,N_8099);
and U12362 (N_12362,N_9411,N_7161);
or U12363 (N_12363,N_6636,N_6584);
and U12364 (N_12364,N_6572,N_7517);
and U12365 (N_12365,N_6949,N_5931);
nand U12366 (N_12366,N_6983,N_7202);
or U12367 (N_12367,N_9057,N_7938);
nor U12368 (N_12368,N_6710,N_5781);
nor U12369 (N_12369,N_7343,N_7156);
nand U12370 (N_12370,N_8732,N_9096);
or U12371 (N_12371,N_5202,N_5562);
or U12372 (N_12372,N_5279,N_6478);
or U12373 (N_12373,N_9432,N_6173);
nand U12374 (N_12374,N_9681,N_7635);
nand U12375 (N_12375,N_6280,N_5002);
and U12376 (N_12376,N_8141,N_5727);
and U12377 (N_12377,N_5915,N_8975);
and U12378 (N_12378,N_8521,N_6564);
and U12379 (N_12379,N_8144,N_5839);
nor U12380 (N_12380,N_8657,N_6496);
nand U12381 (N_12381,N_9871,N_7107);
nor U12382 (N_12382,N_5343,N_7781);
nand U12383 (N_12383,N_5798,N_9235);
or U12384 (N_12384,N_5315,N_8337);
nor U12385 (N_12385,N_5412,N_7061);
and U12386 (N_12386,N_8576,N_7902);
nand U12387 (N_12387,N_7386,N_8390);
nand U12388 (N_12388,N_7983,N_8206);
and U12389 (N_12389,N_9656,N_9925);
nand U12390 (N_12390,N_6441,N_8063);
nand U12391 (N_12391,N_5147,N_9715);
nand U12392 (N_12392,N_7533,N_8956);
nor U12393 (N_12393,N_6763,N_9654);
or U12394 (N_12394,N_6490,N_6037);
or U12395 (N_12395,N_6386,N_5190);
and U12396 (N_12396,N_8889,N_7250);
or U12397 (N_12397,N_8864,N_5642);
nand U12398 (N_12398,N_5288,N_6766);
and U12399 (N_12399,N_9083,N_9116);
nand U12400 (N_12400,N_5807,N_8959);
nand U12401 (N_12401,N_8490,N_8722);
nand U12402 (N_12402,N_7410,N_5188);
nor U12403 (N_12403,N_5738,N_8284);
nor U12404 (N_12404,N_6171,N_5381);
nor U12405 (N_12405,N_8612,N_6405);
xor U12406 (N_12406,N_9639,N_7722);
nor U12407 (N_12407,N_6342,N_5686);
nand U12408 (N_12408,N_9398,N_7052);
or U12409 (N_12409,N_5509,N_9902);
nand U12410 (N_12410,N_5433,N_9629);
nand U12411 (N_12411,N_7407,N_7536);
nor U12412 (N_12412,N_7369,N_7189);
nor U12413 (N_12413,N_7927,N_9310);
or U12414 (N_12414,N_7424,N_7856);
and U12415 (N_12415,N_8626,N_5021);
nand U12416 (N_12416,N_5312,N_7398);
nor U12417 (N_12417,N_5475,N_6347);
nand U12418 (N_12418,N_5508,N_6045);
or U12419 (N_12419,N_7116,N_7193);
nand U12420 (N_12420,N_6962,N_6877);
and U12421 (N_12421,N_5182,N_5737);
nor U12422 (N_12422,N_6561,N_8655);
or U12423 (N_12423,N_9425,N_9016);
or U12424 (N_12424,N_6322,N_6288);
nor U12425 (N_12425,N_6626,N_5184);
or U12426 (N_12426,N_8062,N_8344);
and U12427 (N_12427,N_8366,N_9324);
or U12428 (N_12428,N_8139,N_5818);
or U12429 (N_12429,N_5438,N_9663);
nor U12430 (N_12430,N_5802,N_9468);
or U12431 (N_12431,N_5272,N_7170);
nor U12432 (N_12432,N_5660,N_8198);
and U12433 (N_12433,N_9351,N_5681);
nand U12434 (N_12434,N_6222,N_9747);
and U12435 (N_12435,N_7301,N_5407);
nand U12436 (N_12436,N_7401,N_5304);
nand U12437 (N_12437,N_5379,N_7357);
nor U12438 (N_12438,N_8697,N_9285);
nor U12439 (N_12439,N_9089,N_7005);
or U12440 (N_12440,N_9740,N_8838);
or U12441 (N_12441,N_6683,N_5022);
nor U12442 (N_12442,N_6219,N_5179);
nor U12443 (N_12443,N_9578,N_5096);
nor U12444 (N_12444,N_9204,N_6611);
or U12445 (N_12445,N_5452,N_7355);
nand U12446 (N_12446,N_5497,N_8242);
or U12447 (N_12447,N_6527,N_7122);
nand U12448 (N_12448,N_9989,N_6091);
nand U12449 (N_12449,N_6188,N_6246);
and U12450 (N_12450,N_9660,N_8043);
or U12451 (N_12451,N_5827,N_5396);
or U12452 (N_12452,N_7287,N_8195);
and U12453 (N_12453,N_9729,N_7627);
and U12454 (N_12454,N_7819,N_7715);
nand U12455 (N_12455,N_5941,N_7211);
nor U12456 (N_12456,N_9202,N_7958);
nor U12457 (N_12457,N_5570,N_6579);
or U12458 (N_12458,N_5088,N_8572);
and U12459 (N_12459,N_8331,N_8224);
nand U12460 (N_12460,N_7947,N_8425);
nand U12461 (N_12461,N_7777,N_7148);
or U12462 (N_12462,N_9804,N_7518);
nor U12463 (N_12463,N_5216,N_8517);
or U12464 (N_12464,N_8714,N_7981);
nor U12465 (N_12465,N_7012,N_8248);
nand U12466 (N_12466,N_7415,N_7659);
or U12467 (N_12467,N_9614,N_7184);
or U12468 (N_12468,N_8597,N_5825);
nor U12469 (N_12469,N_6193,N_7183);
nand U12470 (N_12470,N_6507,N_7891);
or U12471 (N_12471,N_9087,N_7171);
nand U12472 (N_12472,N_5259,N_7340);
nand U12473 (N_12473,N_7046,N_9935);
nand U12474 (N_12474,N_8393,N_7753);
and U12475 (N_12475,N_5859,N_6720);
nor U12476 (N_12476,N_6806,N_6082);
and U12477 (N_12477,N_6977,N_8143);
nor U12478 (N_12478,N_7451,N_9633);
nor U12479 (N_12479,N_8497,N_8443);
nand U12480 (N_12480,N_9343,N_5927);
and U12481 (N_12481,N_7712,N_7462);
and U12482 (N_12482,N_9643,N_9507);
nand U12483 (N_12483,N_7591,N_8792);
nand U12484 (N_12484,N_6195,N_8216);
nand U12485 (N_12485,N_8859,N_6015);
nor U12486 (N_12486,N_7139,N_5972);
nand U12487 (N_12487,N_5112,N_5137);
and U12488 (N_12488,N_8800,N_8039);
or U12489 (N_12489,N_6821,N_8371);
or U12490 (N_12490,N_9612,N_9490);
and U12491 (N_12491,N_6896,N_7571);
nor U12492 (N_12492,N_6727,N_7118);
and U12493 (N_12493,N_5722,N_9207);
nor U12494 (N_12494,N_6708,N_9648);
nor U12495 (N_12495,N_6772,N_6957);
nand U12496 (N_12496,N_5561,N_5893);
or U12497 (N_12497,N_7008,N_5689);
nand U12498 (N_12498,N_7298,N_5234);
and U12499 (N_12499,N_5890,N_8727);
nor U12500 (N_12500,N_5058,N_9428);
nand U12501 (N_12501,N_8078,N_6270);
and U12502 (N_12502,N_5904,N_7333);
nor U12503 (N_12503,N_8904,N_7514);
nor U12504 (N_12504,N_7978,N_8234);
and U12505 (N_12505,N_6235,N_9013);
nor U12506 (N_12506,N_8504,N_8768);
or U12507 (N_12507,N_8243,N_5360);
nand U12508 (N_12508,N_9094,N_9463);
nand U12509 (N_12509,N_6617,N_6713);
or U12510 (N_12510,N_7630,N_8816);
nor U12511 (N_12511,N_5529,N_5605);
and U12512 (N_12512,N_5153,N_6296);
nor U12513 (N_12513,N_6168,N_5906);
nor U12514 (N_12514,N_9352,N_5788);
or U12515 (N_12515,N_8570,N_6925);
and U12516 (N_12516,N_6124,N_5155);
nand U12517 (N_12517,N_9363,N_7458);
and U12518 (N_12518,N_5245,N_7291);
nand U12519 (N_12519,N_5356,N_6526);
or U12520 (N_12520,N_5857,N_6726);
nand U12521 (N_12521,N_6514,N_6755);
nor U12522 (N_12522,N_9786,N_6911);
nand U12523 (N_12523,N_7059,N_9823);
nand U12524 (N_12524,N_6861,N_9583);
nor U12525 (N_12525,N_8749,N_8775);
nor U12526 (N_12526,N_6670,N_9236);
and U12527 (N_12527,N_6327,N_7712);
and U12528 (N_12528,N_9723,N_6648);
or U12529 (N_12529,N_9170,N_9619);
and U12530 (N_12530,N_6208,N_8993);
nand U12531 (N_12531,N_6064,N_9525);
nor U12532 (N_12532,N_8430,N_9634);
nand U12533 (N_12533,N_7709,N_6030);
or U12534 (N_12534,N_6177,N_9786);
and U12535 (N_12535,N_6827,N_8621);
nor U12536 (N_12536,N_6913,N_5022);
nor U12537 (N_12537,N_7659,N_5053);
and U12538 (N_12538,N_9506,N_5293);
nand U12539 (N_12539,N_9532,N_5046);
and U12540 (N_12540,N_5054,N_5329);
and U12541 (N_12541,N_8286,N_9282);
nand U12542 (N_12542,N_7404,N_6029);
and U12543 (N_12543,N_9457,N_9127);
or U12544 (N_12544,N_8923,N_6982);
nor U12545 (N_12545,N_9385,N_8668);
nor U12546 (N_12546,N_9331,N_6916);
or U12547 (N_12547,N_6857,N_7988);
and U12548 (N_12548,N_9681,N_5327);
xnor U12549 (N_12549,N_8700,N_5941);
nor U12550 (N_12550,N_8895,N_6896);
and U12551 (N_12551,N_8179,N_5534);
nand U12552 (N_12552,N_9368,N_5716);
and U12553 (N_12553,N_7770,N_8102);
or U12554 (N_12554,N_7491,N_5671);
nand U12555 (N_12555,N_8944,N_5872);
nand U12556 (N_12556,N_7279,N_6677);
or U12557 (N_12557,N_8815,N_9203);
nor U12558 (N_12558,N_7521,N_7600);
and U12559 (N_12559,N_9431,N_9550);
nor U12560 (N_12560,N_8371,N_7326);
or U12561 (N_12561,N_6170,N_6680);
nand U12562 (N_12562,N_5480,N_8038);
or U12563 (N_12563,N_5667,N_8940);
nand U12564 (N_12564,N_7913,N_5847);
or U12565 (N_12565,N_5457,N_9474);
nand U12566 (N_12566,N_7426,N_9683);
or U12567 (N_12567,N_7730,N_9856);
and U12568 (N_12568,N_7599,N_7413);
and U12569 (N_12569,N_8589,N_5483);
nand U12570 (N_12570,N_5313,N_8005);
nand U12571 (N_12571,N_6498,N_6646);
and U12572 (N_12572,N_8346,N_5032);
or U12573 (N_12573,N_7311,N_9944);
nor U12574 (N_12574,N_5068,N_7328);
and U12575 (N_12575,N_5049,N_7692);
and U12576 (N_12576,N_8739,N_8371);
and U12577 (N_12577,N_6894,N_9153);
nand U12578 (N_12578,N_9923,N_5456);
or U12579 (N_12579,N_7472,N_9259);
nand U12580 (N_12580,N_5363,N_7776);
or U12581 (N_12581,N_8282,N_9237);
or U12582 (N_12582,N_5029,N_8438);
nand U12583 (N_12583,N_8764,N_9738);
or U12584 (N_12584,N_9286,N_6917);
nor U12585 (N_12585,N_7251,N_5920);
nand U12586 (N_12586,N_8476,N_7801);
and U12587 (N_12587,N_8048,N_8537);
nor U12588 (N_12588,N_6798,N_8674);
and U12589 (N_12589,N_7722,N_6218);
nand U12590 (N_12590,N_7233,N_6726);
nor U12591 (N_12591,N_8389,N_6083);
nor U12592 (N_12592,N_6325,N_5767);
nor U12593 (N_12593,N_9800,N_8200);
nand U12594 (N_12594,N_9618,N_8983);
and U12595 (N_12595,N_7928,N_7615);
or U12596 (N_12596,N_5685,N_9749);
and U12597 (N_12597,N_8692,N_6276);
and U12598 (N_12598,N_7395,N_5399);
nand U12599 (N_12599,N_5479,N_8884);
nand U12600 (N_12600,N_9188,N_8224);
nand U12601 (N_12601,N_8997,N_7256);
nor U12602 (N_12602,N_6252,N_7582);
nor U12603 (N_12603,N_7114,N_7810);
nand U12604 (N_12604,N_5246,N_5446);
xor U12605 (N_12605,N_7964,N_7479);
or U12606 (N_12606,N_5730,N_8475);
nor U12607 (N_12607,N_8876,N_6997);
nand U12608 (N_12608,N_5324,N_8369);
nand U12609 (N_12609,N_7987,N_5762);
xnor U12610 (N_12610,N_7323,N_6186);
xnor U12611 (N_12611,N_9662,N_9021);
and U12612 (N_12612,N_8420,N_9974);
xnor U12613 (N_12613,N_6180,N_6386);
or U12614 (N_12614,N_6650,N_6426);
nand U12615 (N_12615,N_7874,N_7599);
and U12616 (N_12616,N_5951,N_9125);
nand U12617 (N_12617,N_7928,N_8296);
and U12618 (N_12618,N_7733,N_8023);
nor U12619 (N_12619,N_8361,N_5156);
or U12620 (N_12620,N_7169,N_6075);
xnor U12621 (N_12621,N_9380,N_7171);
or U12622 (N_12622,N_6885,N_7206);
and U12623 (N_12623,N_5241,N_6949);
nand U12624 (N_12624,N_8051,N_6059);
or U12625 (N_12625,N_5366,N_5142);
and U12626 (N_12626,N_9740,N_6188);
and U12627 (N_12627,N_7856,N_8590);
and U12628 (N_12628,N_9819,N_9947);
or U12629 (N_12629,N_6648,N_6854);
and U12630 (N_12630,N_5443,N_7205);
and U12631 (N_12631,N_5063,N_6376);
nand U12632 (N_12632,N_7742,N_8315);
nand U12633 (N_12633,N_6833,N_6161);
nand U12634 (N_12634,N_6245,N_8181);
nor U12635 (N_12635,N_7561,N_7019);
nor U12636 (N_12636,N_8124,N_7046);
and U12637 (N_12637,N_6945,N_5627);
nand U12638 (N_12638,N_7012,N_9880);
and U12639 (N_12639,N_8915,N_6680);
or U12640 (N_12640,N_9973,N_5027);
nor U12641 (N_12641,N_5577,N_6112);
and U12642 (N_12642,N_8714,N_8782);
nor U12643 (N_12643,N_9478,N_9715);
or U12644 (N_12644,N_9082,N_5756);
xnor U12645 (N_12645,N_7714,N_9897);
nor U12646 (N_12646,N_8443,N_5834);
nand U12647 (N_12647,N_7572,N_9631);
or U12648 (N_12648,N_8347,N_5789);
and U12649 (N_12649,N_6110,N_7038);
nor U12650 (N_12650,N_9643,N_7505);
nor U12651 (N_12651,N_8486,N_5811);
and U12652 (N_12652,N_9231,N_7470);
and U12653 (N_12653,N_8355,N_5280);
and U12654 (N_12654,N_6866,N_5347);
nand U12655 (N_12655,N_9389,N_9152);
or U12656 (N_12656,N_8186,N_9333);
or U12657 (N_12657,N_8191,N_7836);
nand U12658 (N_12658,N_9489,N_9840);
nand U12659 (N_12659,N_6103,N_9170);
or U12660 (N_12660,N_6223,N_8295);
and U12661 (N_12661,N_7658,N_6682);
nor U12662 (N_12662,N_8928,N_7279);
or U12663 (N_12663,N_6970,N_9662);
nand U12664 (N_12664,N_8197,N_5849);
and U12665 (N_12665,N_9961,N_8932);
or U12666 (N_12666,N_7985,N_6470);
nor U12667 (N_12667,N_8210,N_7880);
nand U12668 (N_12668,N_9528,N_6671);
and U12669 (N_12669,N_8684,N_8775);
nand U12670 (N_12670,N_8180,N_7115);
nand U12671 (N_12671,N_9913,N_5893);
or U12672 (N_12672,N_5427,N_5718);
nand U12673 (N_12673,N_6282,N_5818);
and U12674 (N_12674,N_5892,N_5895);
or U12675 (N_12675,N_5687,N_9529);
and U12676 (N_12676,N_5009,N_6506);
and U12677 (N_12677,N_5516,N_9066);
nor U12678 (N_12678,N_5552,N_5274);
or U12679 (N_12679,N_6138,N_7656);
and U12680 (N_12680,N_6644,N_7089);
nand U12681 (N_12681,N_6834,N_8630);
nor U12682 (N_12682,N_8751,N_7866);
and U12683 (N_12683,N_9635,N_5478);
nor U12684 (N_12684,N_5737,N_7034);
and U12685 (N_12685,N_8843,N_6914);
nand U12686 (N_12686,N_7847,N_6484);
nor U12687 (N_12687,N_5884,N_9645);
nor U12688 (N_12688,N_6792,N_9844);
or U12689 (N_12689,N_5438,N_8729);
nor U12690 (N_12690,N_6542,N_5088);
nand U12691 (N_12691,N_5153,N_9883);
and U12692 (N_12692,N_5089,N_8183);
and U12693 (N_12693,N_7895,N_7168);
and U12694 (N_12694,N_6766,N_6030);
nand U12695 (N_12695,N_9059,N_9216);
nand U12696 (N_12696,N_6657,N_7654);
and U12697 (N_12697,N_9450,N_6931);
or U12698 (N_12698,N_7882,N_6317);
and U12699 (N_12699,N_9193,N_9779);
and U12700 (N_12700,N_5889,N_8762);
nor U12701 (N_12701,N_9236,N_9816);
nand U12702 (N_12702,N_8511,N_9766);
and U12703 (N_12703,N_9822,N_5601);
nor U12704 (N_12704,N_5920,N_8142);
xnor U12705 (N_12705,N_9075,N_5025);
nand U12706 (N_12706,N_7706,N_7472);
nor U12707 (N_12707,N_8400,N_9971);
nand U12708 (N_12708,N_6579,N_5410);
nor U12709 (N_12709,N_7373,N_8469);
and U12710 (N_12710,N_6654,N_7782);
or U12711 (N_12711,N_5877,N_8070);
xor U12712 (N_12712,N_5739,N_9415);
nand U12713 (N_12713,N_9681,N_6969);
or U12714 (N_12714,N_9091,N_5446);
nand U12715 (N_12715,N_8239,N_8322);
or U12716 (N_12716,N_6788,N_7039);
nor U12717 (N_12717,N_6293,N_9171);
and U12718 (N_12718,N_5478,N_5647);
nor U12719 (N_12719,N_7662,N_9427);
nand U12720 (N_12720,N_8955,N_5392);
and U12721 (N_12721,N_8980,N_9976);
and U12722 (N_12722,N_6798,N_6686);
nor U12723 (N_12723,N_8636,N_5799);
nor U12724 (N_12724,N_7434,N_9695);
nor U12725 (N_12725,N_5273,N_7713);
and U12726 (N_12726,N_8803,N_8437);
or U12727 (N_12727,N_6557,N_6896);
or U12728 (N_12728,N_8789,N_7846);
nor U12729 (N_12729,N_8922,N_8354);
xnor U12730 (N_12730,N_6513,N_7426);
nand U12731 (N_12731,N_8265,N_6435);
or U12732 (N_12732,N_8173,N_9213);
and U12733 (N_12733,N_6816,N_7861);
nand U12734 (N_12734,N_6297,N_5851);
and U12735 (N_12735,N_5132,N_9068);
nand U12736 (N_12736,N_8080,N_6017);
nor U12737 (N_12737,N_8914,N_9881);
xor U12738 (N_12738,N_6018,N_9438);
nor U12739 (N_12739,N_9958,N_5924);
nand U12740 (N_12740,N_7036,N_9631);
and U12741 (N_12741,N_8067,N_6057);
and U12742 (N_12742,N_8510,N_8938);
and U12743 (N_12743,N_5963,N_5329);
or U12744 (N_12744,N_6877,N_9046);
nor U12745 (N_12745,N_9644,N_5911);
or U12746 (N_12746,N_6757,N_8105);
nor U12747 (N_12747,N_9723,N_9452);
or U12748 (N_12748,N_6818,N_8681);
nand U12749 (N_12749,N_8490,N_7042);
nand U12750 (N_12750,N_6221,N_9174);
and U12751 (N_12751,N_5932,N_8466);
and U12752 (N_12752,N_6347,N_7277);
xnor U12753 (N_12753,N_6845,N_5131);
nor U12754 (N_12754,N_9182,N_9137);
and U12755 (N_12755,N_5021,N_8889);
xnor U12756 (N_12756,N_7714,N_6298);
or U12757 (N_12757,N_9203,N_7634);
nor U12758 (N_12758,N_5563,N_7943);
nor U12759 (N_12759,N_9806,N_6420);
nor U12760 (N_12760,N_7967,N_7902);
or U12761 (N_12761,N_9714,N_7599);
nand U12762 (N_12762,N_7139,N_6960);
nand U12763 (N_12763,N_9308,N_6511);
nor U12764 (N_12764,N_9894,N_7387);
and U12765 (N_12765,N_9187,N_5819);
nor U12766 (N_12766,N_5511,N_9601);
nand U12767 (N_12767,N_5158,N_8704);
and U12768 (N_12768,N_7910,N_6454);
nor U12769 (N_12769,N_9830,N_7214);
nand U12770 (N_12770,N_5866,N_7017);
nand U12771 (N_12771,N_7208,N_8436);
nor U12772 (N_12772,N_9269,N_7224);
nor U12773 (N_12773,N_8873,N_7403);
nor U12774 (N_12774,N_6023,N_6297);
and U12775 (N_12775,N_7091,N_9639);
nand U12776 (N_12776,N_9512,N_9471);
or U12777 (N_12777,N_9322,N_5997);
or U12778 (N_12778,N_5430,N_8807);
nand U12779 (N_12779,N_5172,N_8135);
nand U12780 (N_12780,N_5206,N_5673);
nand U12781 (N_12781,N_6637,N_9335);
nor U12782 (N_12782,N_5315,N_5208);
xnor U12783 (N_12783,N_5630,N_9367);
and U12784 (N_12784,N_5132,N_8482);
nor U12785 (N_12785,N_7601,N_8778);
nand U12786 (N_12786,N_8093,N_6385);
nor U12787 (N_12787,N_6735,N_7249);
nor U12788 (N_12788,N_8790,N_6718);
and U12789 (N_12789,N_6677,N_6579);
nor U12790 (N_12790,N_9149,N_9174);
or U12791 (N_12791,N_6275,N_9955);
nor U12792 (N_12792,N_6473,N_9368);
nor U12793 (N_12793,N_6332,N_7750);
or U12794 (N_12794,N_8772,N_9196);
nand U12795 (N_12795,N_7332,N_6819);
nor U12796 (N_12796,N_8502,N_5383);
nand U12797 (N_12797,N_8803,N_8120);
nand U12798 (N_12798,N_8562,N_9049);
nor U12799 (N_12799,N_8806,N_6350);
nand U12800 (N_12800,N_6047,N_7614);
nand U12801 (N_12801,N_5860,N_9790);
or U12802 (N_12802,N_7567,N_6922);
or U12803 (N_12803,N_7223,N_7364);
and U12804 (N_12804,N_7635,N_9822);
and U12805 (N_12805,N_8346,N_9941);
nor U12806 (N_12806,N_9370,N_6816);
and U12807 (N_12807,N_8176,N_8942);
nor U12808 (N_12808,N_8040,N_6379);
nor U12809 (N_12809,N_8289,N_7337);
and U12810 (N_12810,N_5818,N_6107);
nor U12811 (N_12811,N_7798,N_8527);
nor U12812 (N_12812,N_8375,N_8736);
or U12813 (N_12813,N_7401,N_7646);
and U12814 (N_12814,N_7393,N_7100);
and U12815 (N_12815,N_7146,N_5912);
nand U12816 (N_12816,N_5515,N_8500);
nor U12817 (N_12817,N_8920,N_5454);
nand U12818 (N_12818,N_6420,N_7158);
or U12819 (N_12819,N_7540,N_5989);
xnor U12820 (N_12820,N_7313,N_9633);
and U12821 (N_12821,N_9890,N_5139);
nand U12822 (N_12822,N_7761,N_5724);
nor U12823 (N_12823,N_6473,N_9936);
or U12824 (N_12824,N_9020,N_5896);
nor U12825 (N_12825,N_5280,N_6489);
or U12826 (N_12826,N_9441,N_8653);
and U12827 (N_12827,N_8786,N_6781);
nor U12828 (N_12828,N_9264,N_7974);
nor U12829 (N_12829,N_8025,N_5923);
nand U12830 (N_12830,N_8237,N_9637);
nor U12831 (N_12831,N_9314,N_7175);
nor U12832 (N_12832,N_5255,N_7738);
or U12833 (N_12833,N_7108,N_5346);
or U12834 (N_12834,N_6333,N_5117);
nor U12835 (N_12835,N_5845,N_6087);
nor U12836 (N_12836,N_8691,N_6772);
or U12837 (N_12837,N_5251,N_5847);
or U12838 (N_12838,N_6200,N_9814);
nand U12839 (N_12839,N_7066,N_5117);
nor U12840 (N_12840,N_9123,N_9711);
and U12841 (N_12841,N_7987,N_8500);
nand U12842 (N_12842,N_7754,N_7668);
or U12843 (N_12843,N_7379,N_6442);
nor U12844 (N_12844,N_6979,N_5632);
xor U12845 (N_12845,N_5194,N_6559);
or U12846 (N_12846,N_9529,N_5454);
nand U12847 (N_12847,N_6295,N_6686);
or U12848 (N_12848,N_7416,N_5253);
or U12849 (N_12849,N_7042,N_8006);
or U12850 (N_12850,N_5680,N_5649);
nor U12851 (N_12851,N_6350,N_5182);
nand U12852 (N_12852,N_5148,N_8880);
nor U12853 (N_12853,N_5981,N_5834);
or U12854 (N_12854,N_9847,N_5777);
or U12855 (N_12855,N_9323,N_9507);
nand U12856 (N_12856,N_5304,N_5394);
nor U12857 (N_12857,N_9486,N_5822);
nor U12858 (N_12858,N_8177,N_7259);
and U12859 (N_12859,N_6304,N_5749);
and U12860 (N_12860,N_9201,N_7512);
nor U12861 (N_12861,N_9499,N_8550);
nand U12862 (N_12862,N_9961,N_8387);
nor U12863 (N_12863,N_7140,N_5512);
nand U12864 (N_12864,N_7563,N_6410);
and U12865 (N_12865,N_5434,N_7691);
nand U12866 (N_12866,N_9078,N_6879);
or U12867 (N_12867,N_6047,N_8332);
and U12868 (N_12868,N_9358,N_5284);
nor U12869 (N_12869,N_7475,N_8870);
nand U12870 (N_12870,N_8217,N_5452);
and U12871 (N_12871,N_7210,N_8059);
or U12872 (N_12872,N_9000,N_8927);
or U12873 (N_12873,N_7321,N_9430);
nand U12874 (N_12874,N_5887,N_7047);
xnor U12875 (N_12875,N_8565,N_6854);
nand U12876 (N_12876,N_6155,N_8949);
and U12877 (N_12877,N_7966,N_5650);
nand U12878 (N_12878,N_5882,N_7913);
nor U12879 (N_12879,N_9066,N_6783);
nor U12880 (N_12880,N_6809,N_7513);
nand U12881 (N_12881,N_8501,N_7595);
and U12882 (N_12882,N_9825,N_9998);
nand U12883 (N_12883,N_5136,N_9343);
and U12884 (N_12884,N_6517,N_6264);
nor U12885 (N_12885,N_5468,N_6171);
or U12886 (N_12886,N_8692,N_8975);
and U12887 (N_12887,N_8126,N_9986);
nand U12888 (N_12888,N_6294,N_8817);
nor U12889 (N_12889,N_8134,N_5855);
nand U12890 (N_12890,N_8802,N_8720);
or U12891 (N_12891,N_6693,N_6722);
nor U12892 (N_12892,N_9302,N_8965);
or U12893 (N_12893,N_9892,N_9714);
nand U12894 (N_12894,N_6955,N_6935);
nand U12895 (N_12895,N_6121,N_6682);
nor U12896 (N_12896,N_6837,N_6431);
nor U12897 (N_12897,N_9763,N_6578);
and U12898 (N_12898,N_6802,N_9925);
or U12899 (N_12899,N_5558,N_9070);
or U12900 (N_12900,N_9265,N_5867);
nor U12901 (N_12901,N_7616,N_7302);
nand U12902 (N_12902,N_6184,N_7399);
or U12903 (N_12903,N_8791,N_6088);
nand U12904 (N_12904,N_6280,N_7848);
xnor U12905 (N_12905,N_6373,N_9007);
and U12906 (N_12906,N_6051,N_8720);
nand U12907 (N_12907,N_9160,N_5138);
nand U12908 (N_12908,N_6183,N_5589);
and U12909 (N_12909,N_8391,N_9560);
nor U12910 (N_12910,N_7564,N_8825);
nor U12911 (N_12911,N_9091,N_9824);
nand U12912 (N_12912,N_7998,N_8242);
and U12913 (N_12913,N_8648,N_9908);
nand U12914 (N_12914,N_6369,N_6064);
or U12915 (N_12915,N_5710,N_7156);
and U12916 (N_12916,N_9450,N_7899);
nor U12917 (N_12917,N_5156,N_9896);
nor U12918 (N_12918,N_8869,N_6760);
nor U12919 (N_12919,N_6730,N_8391);
nor U12920 (N_12920,N_9477,N_5325);
nand U12921 (N_12921,N_5388,N_8076);
and U12922 (N_12922,N_6797,N_6086);
or U12923 (N_12923,N_8229,N_7750);
and U12924 (N_12924,N_6654,N_6983);
nand U12925 (N_12925,N_5375,N_7227);
nor U12926 (N_12926,N_7801,N_6971);
nor U12927 (N_12927,N_6478,N_8826);
nor U12928 (N_12928,N_5414,N_5889);
or U12929 (N_12929,N_8820,N_5184);
or U12930 (N_12930,N_9292,N_7587);
nor U12931 (N_12931,N_6600,N_8662);
nor U12932 (N_12932,N_8604,N_7420);
nand U12933 (N_12933,N_8626,N_5942);
and U12934 (N_12934,N_7447,N_6041);
nor U12935 (N_12935,N_9841,N_5236);
and U12936 (N_12936,N_9054,N_5528);
or U12937 (N_12937,N_5409,N_8231);
nand U12938 (N_12938,N_6828,N_8665);
and U12939 (N_12939,N_6682,N_5375);
nor U12940 (N_12940,N_6036,N_7990);
and U12941 (N_12941,N_5777,N_5548);
and U12942 (N_12942,N_6481,N_6923);
nor U12943 (N_12943,N_5623,N_8828);
and U12944 (N_12944,N_8762,N_8138);
nor U12945 (N_12945,N_9138,N_8333);
nand U12946 (N_12946,N_7744,N_5236);
and U12947 (N_12947,N_7049,N_7857);
nand U12948 (N_12948,N_5576,N_7971);
nand U12949 (N_12949,N_8404,N_6270);
or U12950 (N_12950,N_9185,N_6965);
and U12951 (N_12951,N_5481,N_7102);
and U12952 (N_12952,N_9733,N_9287);
and U12953 (N_12953,N_9759,N_7978);
and U12954 (N_12954,N_6233,N_7666);
or U12955 (N_12955,N_7242,N_9339);
nor U12956 (N_12956,N_5163,N_5443);
nand U12957 (N_12957,N_7299,N_9369);
nor U12958 (N_12958,N_5806,N_9271);
nor U12959 (N_12959,N_9073,N_8040);
nor U12960 (N_12960,N_6398,N_8257);
and U12961 (N_12961,N_8819,N_6248);
nand U12962 (N_12962,N_6239,N_5018);
nand U12963 (N_12963,N_7059,N_9749);
xor U12964 (N_12964,N_8502,N_6406);
nand U12965 (N_12965,N_9039,N_6319);
or U12966 (N_12966,N_5539,N_5722);
or U12967 (N_12967,N_5354,N_6565);
nand U12968 (N_12968,N_7864,N_8332);
and U12969 (N_12969,N_9542,N_7611);
xnor U12970 (N_12970,N_7171,N_8683);
nand U12971 (N_12971,N_9337,N_5126);
or U12972 (N_12972,N_6838,N_8319);
or U12973 (N_12973,N_8768,N_5905);
and U12974 (N_12974,N_9043,N_6555);
or U12975 (N_12975,N_7562,N_9943);
and U12976 (N_12976,N_7962,N_5179);
nand U12977 (N_12977,N_6394,N_9123);
nor U12978 (N_12978,N_7591,N_8179);
and U12979 (N_12979,N_5621,N_9585);
and U12980 (N_12980,N_6773,N_7018);
or U12981 (N_12981,N_6308,N_6595);
nor U12982 (N_12982,N_9596,N_6247);
or U12983 (N_12983,N_5392,N_9069);
or U12984 (N_12984,N_7280,N_8876);
and U12985 (N_12985,N_7733,N_9501);
nand U12986 (N_12986,N_8468,N_8172);
or U12987 (N_12987,N_6164,N_9522);
xor U12988 (N_12988,N_9619,N_6518);
nand U12989 (N_12989,N_9302,N_9917);
and U12990 (N_12990,N_9485,N_5461);
xnor U12991 (N_12991,N_8423,N_8863);
and U12992 (N_12992,N_8105,N_7638);
and U12993 (N_12993,N_9763,N_5535);
or U12994 (N_12994,N_5956,N_8468);
or U12995 (N_12995,N_7559,N_8854);
nand U12996 (N_12996,N_6316,N_8015);
and U12997 (N_12997,N_8109,N_9211);
nand U12998 (N_12998,N_7923,N_5441);
and U12999 (N_12999,N_5818,N_6479);
and U13000 (N_13000,N_7911,N_6389);
xor U13001 (N_13001,N_8813,N_5185);
or U13002 (N_13002,N_7390,N_8948);
nand U13003 (N_13003,N_5822,N_7531);
nand U13004 (N_13004,N_9966,N_9854);
nand U13005 (N_13005,N_8826,N_6328);
or U13006 (N_13006,N_6062,N_9542);
nand U13007 (N_13007,N_7033,N_5674);
and U13008 (N_13008,N_6773,N_8332);
or U13009 (N_13009,N_7075,N_6892);
and U13010 (N_13010,N_5491,N_6802);
nor U13011 (N_13011,N_6033,N_9247);
nand U13012 (N_13012,N_6632,N_5182);
or U13013 (N_13013,N_6940,N_5935);
nand U13014 (N_13014,N_9549,N_6617);
nand U13015 (N_13015,N_6491,N_6370);
nand U13016 (N_13016,N_6273,N_9897);
and U13017 (N_13017,N_9484,N_7087);
or U13018 (N_13018,N_9850,N_6419);
and U13019 (N_13019,N_5191,N_6988);
and U13020 (N_13020,N_8731,N_6853);
and U13021 (N_13021,N_6781,N_7989);
or U13022 (N_13022,N_5201,N_6525);
nand U13023 (N_13023,N_5294,N_5545);
nand U13024 (N_13024,N_7052,N_7908);
nand U13025 (N_13025,N_5399,N_5997);
and U13026 (N_13026,N_9182,N_6323);
and U13027 (N_13027,N_7856,N_6731);
nor U13028 (N_13028,N_9068,N_6934);
and U13029 (N_13029,N_5385,N_6761);
and U13030 (N_13030,N_9906,N_9289);
nand U13031 (N_13031,N_5321,N_9988);
or U13032 (N_13032,N_6375,N_6626);
and U13033 (N_13033,N_5130,N_8246);
and U13034 (N_13034,N_7926,N_9766);
nor U13035 (N_13035,N_6616,N_7321);
or U13036 (N_13036,N_7478,N_8476);
or U13037 (N_13037,N_6820,N_8689);
nor U13038 (N_13038,N_7921,N_5321);
and U13039 (N_13039,N_9573,N_6897);
nand U13040 (N_13040,N_6679,N_9841);
or U13041 (N_13041,N_5677,N_6211);
and U13042 (N_13042,N_7840,N_7132);
nor U13043 (N_13043,N_8256,N_7846);
and U13044 (N_13044,N_9995,N_7989);
and U13045 (N_13045,N_7006,N_9739);
or U13046 (N_13046,N_8216,N_5327);
or U13047 (N_13047,N_7935,N_9566);
nor U13048 (N_13048,N_8966,N_7237);
or U13049 (N_13049,N_9694,N_9256);
nor U13050 (N_13050,N_6646,N_6881);
or U13051 (N_13051,N_7534,N_6132);
or U13052 (N_13052,N_9931,N_5514);
or U13053 (N_13053,N_5837,N_6935);
nand U13054 (N_13054,N_7396,N_6196);
nor U13055 (N_13055,N_6016,N_8345);
and U13056 (N_13056,N_7769,N_6488);
and U13057 (N_13057,N_8348,N_6656);
nor U13058 (N_13058,N_8289,N_9110);
and U13059 (N_13059,N_7642,N_7720);
nand U13060 (N_13060,N_9510,N_6082);
or U13061 (N_13061,N_8224,N_8845);
nor U13062 (N_13062,N_8222,N_6277);
nand U13063 (N_13063,N_5475,N_5723);
and U13064 (N_13064,N_5386,N_5392);
nand U13065 (N_13065,N_9256,N_5724);
nand U13066 (N_13066,N_5753,N_5200);
nand U13067 (N_13067,N_7595,N_6647);
or U13068 (N_13068,N_5751,N_9805);
and U13069 (N_13069,N_7259,N_6815);
nand U13070 (N_13070,N_6037,N_9700);
or U13071 (N_13071,N_6650,N_5170);
or U13072 (N_13072,N_7229,N_5149);
nor U13073 (N_13073,N_7120,N_7613);
and U13074 (N_13074,N_5055,N_7827);
nand U13075 (N_13075,N_7773,N_7191);
nor U13076 (N_13076,N_9237,N_9686);
nor U13077 (N_13077,N_8211,N_9057);
nand U13078 (N_13078,N_9247,N_5727);
or U13079 (N_13079,N_5419,N_6749);
or U13080 (N_13080,N_5923,N_9909);
nor U13081 (N_13081,N_7262,N_5525);
or U13082 (N_13082,N_7529,N_7178);
and U13083 (N_13083,N_7517,N_9292);
nor U13084 (N_13084,N_9806,N_9342);
and U13085 (N_13085,N_6063,N_9400);
or U13086 (N_13086,N_8126,N_7756);
xor U13087 (N_13087,N_9997,N_8762);
nand U13088 (N_13088,N_7336,N_8542);
nand U13089 (N_13089,N_7548,N_5397);
and U13090 (N_13090,N_6334,N_8208);
nor U13091 (N_13091,N_7168,N_6250);
nand U13092 (N_13092,N_7216,N_7673);
and U13093 (N_13093,N_5189,N_9917);
and U13094 (N_13094,N_8590,N_5907);
nand U13095 (N_13095,N_5026,N_7339);
or U13096 (N_13096,N_9522,N_5121);
nor U13097 (N_13097,N_7150,N_8691);
or U13098 (N_13098,N_5121,N_9128);
xnor U13099 (N_13099,N_7103,N_5429);
xor U13100 (N_13100,N_7296,N_8755);
and U13101 (N_13101,N_7194,N_9379);
nor U13102 (N_13102,N_5012,N_8726);
nand U13103 (N_13103,N_8484,N_8700);
nand U13104 (N_13104,N_7056,N_9980);
nor U13105 (N_13105,N_6567,N_8227);
nand U13106 (N_13106,N_6625,N_7081);
nor U13107 (N_13107,N_8844,N_8267);
nor U13108 (N_13108,N_5348,N_8952);
and U13109 (N_13109,N_7364,N_7302);
nand U13110 (N_13110,N_6846,N_8150);
nor U13111 (N_13111,N_5267,N_7546);
and U13112 (N_13112,N_9042,N_5322);
nor U13113 (N_13113,N_7982,N_7992);
and U13114 (N_13114,N_8311,N_6994);
nand U13115 (N_13115,N_5928,N_9501);
or U13116 (N_13116,N_5622,N_9758);
nand U13117 (N_13117,N_7118,N_9759);
and U13118 (N_13118,N_8350,N_6179);
nor U13119 (N_13119,N_6606,N_9858);
or U13120 (N_13120,N_9591,N_8849);
nand U13121 (N_13121,N_7558,N_6825);
nand U13122 (N_13122,N_6778,N_5910);
nor U13123 (N_13123,N_8433,N_8736);
and U13124 (N_13124,N_6992,N_5215);
xor U13125 (N_13125,N_8354,N_6682);
nor U13126 (N_13126,N_7540,N_7297);
nor U13127 (N_13127,N_6080,N_5334);
and U13128 (N_13128,N_7818,N_6496);
nand U13129 (N_13129,N_7254,N_6521);
and U13130 (N_13130,N_6777,N_7171);
nand U13131 (N_13131,N_6667,N_5579);
nand U13132 (N_13132,N_5130,N_7194);
and U13133 (N_13133,N_8481,N_8243);
nand U13134 (N_13134,N_7895,N_6822);
nor U13135 (N_13135,N_6753,N_5776);
and U13136 (N_13136,N_8454,N_7387);
and U13137 (N_13137,N_5161,N_5016);
and U13138 (N_13138,N_8175,N_7214);
or U13139 (N_13139,N_8957,N_8111);
nand U13140 (N_13140,N_7559,N_7755);
or U13141 (N_13141,N_7002,N_6274);
and U13142 (N_13142,N_7643,N_8585);
and U13143 (N_13143,N_8988,N_7558);
or U13144 (N_13144,N_8916,N_7222);
nand U13145 (N_13145,N_7163,N_5698);
and U13146 (N_13146,N_9257,N_6793);
nor U13147 (N_13147,N_7179,N_8759);
nor U13148 (N_13148,N_9626,N_6759);
nor U13149 (N_13149,N_7967,N_5322);
xor U13150 (N_13150,N_8053,N_5544);
and U13151 (N_13151,N_7701,N_7931);
nand U13152 (N_13152,N_7082,N_7863);
or U13153 (N_13153,N_8288,N_8294);
or U13154 (N_13154,N_7667,N_8976);
or U13155 (N_13155,N_5368,N_8474);
and U13156 (N_13156,N_5574,N_8044);
nand U13157 (N_13157,N_5015,N_5204);
or U13158 (N_13158,N_9778,N_5375);
nor U13159 (N_13159,N_8791,N_5324);
and U13160 (N_13160,N_6978,N_7311);
or U13161 (N_13161,N_9324,N_9494);
nor U13162 (N_13162,N_8148,N_5649);
nor U13163 (N_13163,N_7577,N_6871);
nor U13164 (N_13164,N_7675,N_5515);
and U13165 (N_13165,N_9928,N_9698);
nand U13166 (N_13166,N_9442,N_6949);
and U13167 (N_13167,N_8946,N_9514);
or U13168 (N_13168,N_5899,N_7303);
or U13169 (N_13169,N_8420,N_7978);
nor U13170 (N_13170,N_7492,N_8658);
xor U13171 (N_13171,N_8266,N_6203);
and U13172 (N_13172,N_9689,N_6770);
or U13173 (N_13173,N_9977,N_6702);
or U13174 (N_13174,N_5574,N_5798);
nand U13175 (N_13175,N_6755,N_7799);
or U13176 (N_13176,N_8767,N_8978);
nand U13177 (N_13177,N_6232,N_7273);
or U13178 (N_13178,N_9340,N_8803);
or U13179 (N_13179,N_5408,N_7056);
nand U13180 (N_13180,N_8906,N_9249);
nand U13181 (N_13181,N_7998,N_5315);
nand U13182 (N_13182,N_8762,N_6769);
or U13183 (N_13183,N_6774,N_7781);
or U13184 (N_13184,N_5127,N_9745);
nor U13185 (N_13185,N_7261,N_9486);
nor U13186 (N_13186,N_7938,N_9699);
nand U13187 (N_13187,N_8688,N_7667);
nand U13188 (N_13188,N_9614,N_9343);
and U13189 (N_13189,N_9402,N_7623);
and U13190 (N_13190,N_7467,N_5185);
xnor U13191 (N_13191,N_5518,N_7822);
nand U13192 (N_13192,N_6193,N_5882);
nand U13193 (N_13193,N_8986,N_6227);
and U13194 (N_13194,N_7413,N_5174);
and U13195 (N_13195,N_8126,N_6260);
nand U13196 (N_13196,N_9044,N_5411);
or U13197 (N_13197,N_5976,N_6062);
or U13198 (N_13198,N_5214,N_8662);
and U13199 (N_13199,N_6434,N_9505);
nand U13200 (N_13200,N_7680,N_8101);
or U13201 (N_13201,N_9416,N_9451);
or U13202 (N_13202,N_5417,N_8566);
nand U13203 (N_13203,N_8557,N_6937);
nand U13204 (N_13204,N_7116,N_6869);
and U13205 (N_13205,N_7153,N_6377);
nor U13206 (N_13206,N_7356,N_5437);
or U13207 (N_13207,N_9165,N_9920);
nand U13208 (N_13208,N_6532,N_7238);
or U13209 (N_13209,N_9468,N_7563);
and U13210 (N_13210,N_8412,N_7573);
nor U13211 (N_13211,N_5390,N_6373);
nand U13212 (N_13212,N_6608,N_5752);
and U13213 (N_13213,N_6021,N_7492);
or U13214 (N_13214,N_8369,N_7088);
nand U13215 (N_13215,N_5563,N_6899);
xnor U13216 (N_13216,N_9627,N_5139);
and U13217 (N_13217,N_6220,N_9679);
nor U13218 (N_13218,N_6255,N_6300);
and U13219 (N_13219,N_7321,N_5993);
xor U13220 (N_13220,N_8001,N_9278);
or U13221 (N_13221,N_6004,N_9236);
and U13222 (N_13222,N_7795,N_8047);
nor U13223 (N_13223,N_6875,N_9740);
nor U13224 (N_13224,N_9277,N_6650);
nor U13225 (N_13225,N_8078,N_9700);
nor U13226 (N_13226,N_5298,N_7163);
or U13227 (N_13227,N_5923,N_8378);
and U13228 (N_13228,N_6194,N_7183);
nand U13229 (N_13229,N_6453,N_8447);
and U13230 (N_13230,N_9258,N_5403);
and U13231 (N_13231,N_5351,N_6353);
or U13232 (N_13232,N_6971,N_7958);
and U13233 (N_13233,N_9369,N_9914);
nor U13234 (N_13234,N_8196,N_8213);
and U13235 (N_13235,N_5798,N_9888);
or U13236 (N_13236,N_7365,N_9565);
nor U13237 (N_13237,N_9654,N_6512);
nor U13238 (N_13238,N_6542,N_5677);
nand U13239 (N_13239,N_7962,N_6315);
or U13240 (N_13240,N_7523,N_7764);
and U13241 (N_13241,N_7666,N_6120);
and U13242 (N_13242,N_5868,N_5410);
or U13243 (N_13243,N_5287,N_8295);
nand U13244 (N_13244,N_6648,N_5425);
nor U13245 (N_13245,N_5199,N_6959);
nor U13246 (N_13246,N_5023,N_6519);
nand U13247 (N_13247,N_9081,N_9483);
nor U13248 (N_13248,N_5170,N_5387);
or U13249 (N_13249,N_5635,N_5539);
or U13250 (N_13250,N_8775,N_6904);
or U13251 (N_13251,N_7366,N_7761);
and U13252 (N_13252,N_7734,N_8995);
and U13253 (N_13253,N_5052,N_8277);
or U13254 (N_13254,N_6608,N_6219);
or U13255 (N_13255,N_5928,N_8684);
nand U13256 (N_13256,N_7317,N_8412);
nor U13257 (N_13257,N_9594,N_6088);
or U13258 (N_13258,N_7271,N_7967);
and U13259 (N_13259,N_5841,N_6732);
nor U13260 (N_13260,N_8593,N_7117);
nand U13261 (N_13261,N_9231,N_5445);
nand U13262 (N_13262,N_9391,N_8384);
xor U13263 (N_13263,N_7621,N_6828);
or U13264 (N_13264,N_8616,N_6771);
nand U13265 (N_13265,N_9915,N_5525);
or U13266 (N_13266,N_9460,N_5972);
or U13267 (N_13267,N_8118,N_8137);
nor U13268 (N_13268,N_6982,N_9527);
or U13269 (N_13269,N_6174,N_5612);
nand U13270 (N_13270,N_7134,N_9766);
or U13271 (N_13271,N_5810,N_8956);
and U13272 (N_13272,N_5154,N_9803);
or U13273 (N_13273,N_7000,N_8235);
nor U13274 (N_13274,N_6828,N_5987);
or U13275 (N_13275,N_6663,N_8351);
nor U13276 (N_13276,N_7092,N_8510);
and U13277 (N_13277,N_5547,N_9400);
and U13278 (N_13278,N_5825,N_7959);
nor U13279 (N_13279,N_9408,N_7412);
nor U13280 (N_13280,N_7963,N_7356);
nor U13281 (N_13281,N_5583,N_9632);
or U13282 (N_13282,N_6091,N_9065);
nor U13283 (N_13283,N_8314,N_7490);
and U13284 (N_13284,N_9925,N_7570);
nand U13285 (N_13285,N_8753,N_9929);
or U13286 (N_13286,N_9083,N_6146);
and U13287 (N_13287,N_7643,N_5981);
nand U13288 (N_13288,N_5354,N_8051);
or U13289 (N_13289,N_6823,N_9942);
or U13290 (N_13290,N_6950,N_8930);
nand U13291 (N_13291,N_7796,N_6926);
or U13292 (N_13292,N_7586,N_8612);
nor U13293 (N_13293,N_8985,N_8924);
and U13294 (N_13294,N_9090,N_7328);
nor U13295 (N_13295,N_6069,N_5230);
and U13296 (N_13296,N_6105,N_8511);
nor U13297 (N_13297,N_9126,N_9735);
nor U13298 (N_13298,N_9117,N_8575);
nand U13299 (N_13299,N_5192,N_5383);
or U13300 (N_13300,N_9860,N_9357);
nand U13301 (N_13301,N_6819,N_5271);
or U13302 (N_13302,N_9076,N_5596);
and U13303 (N_13303,N_7700,N_8343);
nand U13304 (N_13304,N_9875,N_6021);
nor U13305 (N_13305,N_9664,N_7017);
nor U13306 (N_13306,N_9148,N_6079);
nor U13307 (N_13307,N_7413,N_9237);
nand U13308 (N_13308,N_5768,N_6831);
nand U13309 (N_13309,N_8320,N_7163);
nor U13310 (N_13310,N_6249,N_6748);
nand U13311 (N_13311,N_8806,N_7697);
nor U13312 (N_13312,N_8967,N_6863);
or U13313 (N_13313,N_7377,N_6672);
nor U13314 (N_13314,N_7401,N_7084);
or U13315 (N_13315,N_8094,N_6276);
and U13316 (N_13316,N_7017,N_7335);
or U13317 (N_13317,N_8990,N_7900);
nor U13318 (N_13318,N_8924,N_5327);
and U13319 (N_13319,N_6406,N_9167);
or U13320 (N_13320,N_6177,N_9569);
nor U13321 (N_13321,N_5970,N_9335);
and U13322 (N_13322,N_7156,N_9720);
nor U13323 (N_13323,N_9264,N_7881);
nand U13324 (N_13324,N_7461,N_8128);
nor U13325 (N_13325,N_5875,N_8063);
and U13326 (N_13326,N_9194,N_8014);
or U13327 (N_13327,N_9773,N_9401);
nand U13328 (N_13328,N_7833,N_6593);
and U13329 (N_13329,N_7212,N_9810);
or U13330 (N_13330,N_8760,N_9354);
nor U13331 (N_13331,N_7655,N_5889);
and U13332 (N_13332,N_9685,N_6395);
nor U13333 (N_13333,N_9431,N_7932);
or U13334 (N_13334,N_5221,N_7264);
nand U13335 (N_13335,N_6827,N_6251);
nand U13336 (N_13336,N_6586,N_7448);
nand U13337 (N_13337,N_5971,N_5545);
nor U13338 (N_13338,N_7122,N_5735);
or U13339 (N_13339,N_7161,N_6220);
nor U13340 (N_13340,N_5807,N_9859);
nand U13341 (N_13341,N_6963,N_5612);
or U13342 (N_13342,N_5985,N_8267);
nor U13343 (N_13343,N_9430,N_9055);
and U13344 (N_13344,N_6777,N_5671);
and U13345 (N_13345,N_6744,N_7335);
or U13346 (N_13346,N_5727,N_5929);
and U13347 (N_13347,N_6201,N_9656);
or U13348 (N_13348,N_7041,N_8639);
nor U13349 (N_13349,N_6582,N_5863);
and U13350 (N_13350,N_7914,N_8626);
and U13351 (N_13351,N_6221,N_5785);
xor U13352 (N_13352,N_9952,N_5111);
nand U13353 (N_13353,N_8178,N_7095);
nor U13354 (N_13354,N_7922,N_6779);
nand U13355 (N_13355,N_6231,N_7863);
nor U13356 (N_13356,N_6638,N_7008);
nor U13357 (N_13357,N_8786,N_7153);
and U13358 (N_13358,N_5408,N_7964);
or U13359 (N_13359,N_5433,N_7140);
nand U13360 (N_13360,N_6683,N_8658);
and U13361 (N_13361,N_6102,N_5235);
nor U13362 (N_13362,N_8994,N_5846);
nand U13363 (N_13363,N_8843,N_9765);
nand U13364 (N_13364,N_5338,N_6830);
nor U13365 (N_13365,N_7935,N_5902);
or U13366 (N_13366,N_9772,N_9905);
nand U13367 (N_13367,N_9184,N_5881);
nand U13368 (N_13368,N_6759,N_6054);
and U13369 (N_13369,N_8113,N_6753);
nor U13370 (N_13370,N_6840,N_8284);
and U13371 (N_13371,N_9752,N_6746);
or U13372 (N_13372,N_5892,N_9310);
nand U13373 (N_13373,N_9702,N_9781);
or U13374 (N_13374,N_7604,N_5904);
and U13375 (N_13375,N_5070,N_8465);
and U13376 (N_13376,N_6141,N_7777);
nand U13377 (N_13377,N_9834,N_6285);
xor U13378 (N_13378,N_7364,N_6078);
and U13379 (N_13379,N_9811,N_9797);
nor U13380 (N_13380,N_5128,N_5738);
or U13381 (N_13381,N_7002,N_5018);
nand U13382 (N_13382,N_8449,N_6600);
and U13383 (N_13383,N_8676,N_7266);
nand U13384 (N_13384,N_5484,N_7240);
or U13385 (N_13385,N_6466,N_8145);
or U13386 (N_13386,N_7331,N_8179);
and U13387 (N_13387,N_6654,N_8919);
or U13388 (N_13388,N_7740,N_9363);
nor U13389 (N_13389,N_7426,N_8047);
and U13390 (N_13390,N_5652,N_5571);
nor U13391 (N_13391,N_9962,N_8903);
nor U13392 (N_13392,N_9353,N_9596);
nand U13393 (N_13393,N_7438,N_5341);
or U13394 (N_13394,N_8518,N_7534);
nor U13395 (N_13395,N_5216,N_5505);
or U13396 (N_13396,N_7428,N_5722);
nand U13397 (N_13397,N_9461,N_6536);
or U13398 (N_13398,N_9752,N_8564);
or U13399 (N_13399,N_5143,N_8868);
and U13400 (N_13400,N_6898,N_6251);
nor U13401 (N_13401,N_7995,N_9609);
nor U13402 (N_13402,N_7636,N_5090);
nor U13403 (N_13403,N_5003,N_6729);
nor U13404 (N_13404,N_7393,N_6841);
or U13405 (N_13405,N_7591,N_6417);
nand U13406 (N_13406,N_6719,N_7173);
and U13407 (N_13407,N_5176,N_8164);
nand U13408 (N_13408,N_6047,N_5840);
nor U13409 (N_13409,N_5899,N_6356);
nor U13410 (N_13410,N_9012,N_8151);
nand U13411 (N_13411,N_5225,N_9178);
and U13412 (N_13412,N_6940,N_9573);
nor U13413 (N_13413,N_7163,N_6567);
and U13414 (N_13414,N_5796,N_9212);
and U13415 (N_13415,N_6554,N_6941);
xor U13416 (N_13416,N_7925,N_5596);
or U13417 (N_13417,N_9784,N_8963);
xor U13418 (N_13418,N_7160,N_9044);
or U13419 (N_13419,N_9867,N_8038);
nand U13420 (N_13420,N_7082,N_9370);
nand U13421 (N_13421,N_8920,N_5058);
xor U13422 (N_13422,N_7157,N_5886);
and U13423 (N_13423,N_5689,N_8836);
nand U13424 (N_13424,N_8792,N_7565);
and U13425 (N_13425,N_9822,N_6544);
and U13426 (N_13426,N_7222,N_8748);
nand U13427 (N_13427,N_6478,N_5668);
and U13428 (N_13428,N_5479,N_8866);
and U13429 (N_13429,N_9576,N_8778);
nor U13430 (N_13430,N_9050,N_6673);
nand U13431 (N_13431,N_6965,N_8889);
or U13432 (N_13432,N_5602,N_6025);
nand U13433 (N_13433,N_9372,N_5082);
and U13434 (N_13434,N_5426,N_6083);
nor U13435 (N_13435,N_9864,N_5084);
or U13436 (N_13436,N_9583,N_6494);
and U13437 (N_13437,N_8863,N_6330);
or U13438 (N_13438,N_8801,N_6625);
or U13439 (N_13439,N_7079,N_7980);
and U13440 (N_13440,N_7287,N_7247);
nand U13441 (N_13441,N_7873,N_9664);
nand U13442 (N_13442,N_7529,N_7758);
nor U13443 (N_13443,N_5204,N_9553);
nor U13444 (N_13444,N_7315,N_7733);
nor U13445 (N_13445,N_6587,N_6383);
or U13446 (N_13446,N_9190,N_7854);
nand U13447 (N_13447,N_9582,N_8413);
nor U13448 (N_13448,N_5694,N_8497);
nor U13449 (N_13449,N_9551,N_8769);
nand U13450 (N_13450,N_7308,N_8373);
nand U13451 (N_13451,N_7756,N_8984);
and U13452 (N_13452,N_7588,N_5434);
and U13453 (N_13453,N_8371,N_8053);
nand U13454 (N_13454,N_6508,N_6360);
xnor U13455 (N_13455,N_5694,N_6637);
nor U13456 (N_13456,N_8490,N_6284);
nor U13457 (N_13457,N_8727,N_9257);
nor U13458 (N_13458,N_8617,N_6585);
nor U13459 (N_13459,N_7535,N_7904);
and U13460 (N_13460,N_6396,N_5392);
nand U13461 (N_13461,N_6988,N_9393);
nand U13462 (N_13462,N_8792,N_5410);
nand U13463 (N_13463,N_5563,N_8777);
nand U13464 (N_13464,N_9122,N_5330);
or U13465 (N_13465,N_8660,N_8989);
xnor U13466 (N_13466,N_7097,N_7032);
nand U13467 (N_13467,N_8806,N_6372);
nand U13468 (N_13468,N_5704,N_5887);
nor U13469 (N_13469,N_5690,N_9178);
nor U13470 (N_13470,N_9110,N_7929);
xor U13471 (N_13471,N_8583,N_5084);
and U13472 (N_13472,N_8197,N_7044);
nand U13473 (N_13473,N_6952,N_7635);
and U13474 (N_13474,N_7041,N_8560);
nand U13475 (N_13475,N_5732,N_9189);
nor U13476 (N_13476,N_8770,N_6431);
and U13477 (N_13477,N_7466,N_6047);
nor U13478 (N_13478,N_6616,N_9344);
nor U13479 (N_13479,N_6489,N_8944);
nand U13480 (N_13480,N_5795,N_5642);
nor U13481 (N_13481,N_9030,N_6460);
nand U13482 (N_13482,N_9236,N_7532);
xnor U13483 (N_13483,N_7514,N_7653);
and U13484 (N_13484,N_9694,N_8698);
nor U13485 (N_13485,N_7459,N_8987);
and U13486 (N_13486,N_6418,N_9213);
nand U13487 (N_13487,N_8750,N_5634);
nand U13488 (N_13488,N_5946,N_6921);
and U13489 (N_13489,N_9822,N_7356);
nor U13490 (N_13490,N_9740,N_9583);
or U13491 (N_13491,N_7375,N_5674);
and U13492 (N_13492,N_7834,N_7936);
xor U13493 (N_13493,N_6101,N_9595);
nor U13494 (N_13494,N_6003,N_7881);
and U13495 (N_13495,N_8641,N_7018);
nor U13496 (N_13496,N_6003,N_9053);
or U13497 (N_13497,N_6809,N_6985);
nand U13498 (N_13498,N_8332,N_7700);
nand U13499 (N_13499,N_5693,N_9723);
nand U13500 (N_13500,N_6480,N_8036);
or U13501 (N_13501,N_8205,N_5078);
or U13502 (N_13502,N_7432,N_8085);
and U13503 (N_13503,N_9263,N_8657);
nor U13504 (N_13504,N_5614,N_7765);
and U13505 (N_13505,N_8245,N_7123);
nor U13506 (N_13506,N_9865,N_6321);
nor U13507 (N_13507,N_9408,N_7603);
nand U13508 (N_13508,N_6050,N_8153);
nand U13509 (N_13509,N_5516,N_9220);
or U13510 (N_13510,N_8307,N_9997);
nand U13511 (N_13511,N_5260,N_5529);
and U13512 (N_13512,N_8868,N_8196);
nand U13513 (N_13513,N_6492,N_9766);
and U13514 (N_13514,N_9247,N_8082);
and U13515 (N_13515,N_9363,N_9887);
or U13516 (N_13516,N_6064,N_5033);
or U13517 (N_13517,N_6268,N_6745);
or U13518 (N_13518,N_7376,N_6938);
or U13519 (N_13519,N_8369,N_9058);
and U13520 (N_13520,N_8843,N_8799);
or U13521 (N_13521,N_6592,N_9465);
and U13522 (N_13522,N_9573,N_6466);
or U13523 (N_13523,N_6847,N_8848);
or U13524 (N_13524,N_9090,N_6272);
and U13525 (N_13525,N_5938,N_6799);
nor U13526 (N_13526,N_7167,N_5823);
nor U13527 (N_13527,N_5352,N_8641);
or U13528 (N_13528,N_6391,N_6868);
and U13529 (N_13529,N_7351,N_7305);
nor U13530 (N_13530,N_7199,N_7964);
nor U13531 (N_13531,N_6529,N_8897);
nand U13532 (N_13532,N_6771,N_6983);
nor U13533 (N_13533,N_5277,N_5044);
nand U13534 (N_13534,N_8601,N_9649);
or U13535 (N_13535,N_8126,N_7935);
nand U13536 (N_13536,N_6801,N_5412);
and U13537 (N_13537,N_7186,N_6445);
nand U13538 (N_13538,N_5778,N_6042);
and U13539 (N_13539,N_9038,N_8025);
nor U13540 (N_13540,N_6584,N_6480);
and U13541 (N_13541,N_7426,N_5377);
nor U13542 (N_13542,N_8687,N_7176);
xor U13543 (N_13543,N_6186,N_5877);
or U13544 (N_13544,N_8640,N_7593);
nor U13545 (N_13545,N_5126,N_8803);
nor U13546 (N_13546,N_7345,N_9562);
or U13547 (N_13547,N_6190,N_6892);
and U13548 (N_13548,N_5568,N_5649);
or U13549 (N_13549,N_7392,N_9598);
nor U13550 (N_13550,N_7797,N_9557);
nor U13551 (N_13551,N_5360,N_6543);
and U13552 (N_13552,N_9258,N_5480);
nor U13553 (N_13553,N_8064,N_7727);
nor U13554 (N_13554,N_8027,N_5709);
and U13555 (N_13555,N_9364,N_7382);
nand U13556 (N_13556,N_5054,N_6279);
xnor U13557 (N_13557,N_6917,N_9181);
nand U13558 (N_13558,N_8946,N_9321);
or U13559 (N_13559,N_7077,N_6904);
and U13560 (N_13560,N_5057,N_7273);
nand U13561 (N_13561,N_6293,N_9347);
and U13562 (N_13562,N_5349,N_8802);
or U13563 (N_13563,N_8632,N_5771);
or U13564 (N_13564,N_7585,N_6450);
nor U13565 (N_13565,N_6868,N_6136);
and U13566 (N_13566,N_6871,N_9215);
or U13567 (N_13567,N_5789,N_7021);
and U13568 (N_13568,N_6746,N_9045);
or U13569 (N_13569,N_9394,N_9637);
or U13570 (N_13570,N_7460,N_8554);
nand U13571 (N_13571,N_8520,N_6856);
nand U13572 (N_13572,N_5616,N_7302);
or U13573 (N_13573,N_7020,N_5900);
nand U13574 (N_13574,N_5212,N_8100);
or U13575 (N_13575,N_6583,N_8456);
nor U13576 (N_13576,N_7494,N_8158);
nand U13577 (N_13577,N_8338,N_6295);
or U13578 (N_13578,N_8822,N_9706);
nor U13579 (N_13579,N_9013,N_7377);
nor U13580 (N_13580,N_9799,N_7330);
nand U13581 (N_13581,N_5334,N_5786);
and U13582 (N_13582,N_9335,N_5246);
or U13583 (N_13583,N_5141,N_7034);
and U13584 (N_13584,N_5415,N_9190);
and U13585 (N_13585,N_7546,N_8980);
or U13586 (N_13586,N_8133,N_5986);
nor U13587 (N_13587,N_9509,N_6069);
nor U13588 (N_13588,N_8979,N_5894);
nand U13589 (N_13589,N_9101,N_7255);
and U13590 (N_13590,N_6320,N_5612);
xor U13591 (N_13591,N_7243,N_6489);
nand U13592 (N_13592,N_8968,N_7126);
and U13593 (N_13593,N_9728,N_7657);
or U13594 (N_13594,N_7883,N_6483);
or U13595 (N_13595,N_8265,N_5223);
nand U13596 (N_13596,N_7542,N_8648);
nand U13597 (N_13597,N_7837,N_8635);
nor U13598 (N_13598,N_9185,N_6516);
or U13599 (N_13599,N_8107,N_5240);
and U13600 (N_13600,N_9581,N_8290);
nor U13601 (N_13601,N_5809,N_7460);
nor U13602 (N_13602,N_8139,N_7362);
nor U13603 (N_13603,N_6997,N_6153);
or U13604 (N_13604,N_6960,N_5453);
or U13605 (N_13605,N_5092,N_6845);
nor U13606 (N_13606,N_7205,N_9629);
nand U13607 (N_13607,N_6184,N_8798);
nor U13608 (N_13608,N_7546,N_8735);
and U13609 (N_13609,N_6459,N_8238);
nand U13610 (N_13610,N_7292,N_7607);
or U13611 (N_13611,N_5506,N_8844);
or U13612 (N_13612,N_8980,N_8352);
nand U13613 (N_13613,N_8824,N_5342);
and U13614 (N_13614,N_6745,N_7623);
or U13615 (N_13615,N_7875,N_6291);
and U13616 (N_13616,N_6765,N_5120);
nand U13617 (N_13617,N_7730,N_7610);
nand U13618 (N_13618,N_6213,N_6266);
and U13619 (N_13619,N_5556,N_5682);
or U13620 (N_13620,N_7227,N_5452);
nor U13621 (N_13621,N_9718,N_8343);
or U13622 (N_13622,N_6564,N_8223);
or U13623 (N_13623,N_6844,N_6575);
nand U13624 (N_13624,N_5451,N_6448);
nor U13625 (N_13625,N_8256,N_9579);
nor U13626 (N_13626,N_9002,N_5016);
or U13627 (N_13627,N_6428,N_8459);
and U13628 (N_13628,N_5555,N_5638);
or U13629 (N_13629,N_7769,N_5419);
nand U13630 (N_13630,N_6917,N_9780);
and U13631 (N_13631,N_9506,N_6237);
or U13632 (N_13632,N_6086,N_6326);
and U13633 (N_13633,N_6216,N_6288);
nand U13634 (N_13634,N_6378,N_9997);
nor U13635 (N_13635,N_8880,N_6856);
nand U13636 (N_13636,N_5099,N_5176);
or U13637 (N_13637,N_9434,N_6578);
and U13638 (N_13638,N_8469,N_6831);
or U13639 (N_13639,N_8524,N_7047);
or U13640 (N_13640,N_8608,N_6527);
or U13641 (N_13641,N_6955,N_6580);
and U13642 (N_13642,N_6439,N_9595);
nor U13643 (N_13643,N_6656,N_9335);
or U13644 (N_13644,N_7152,N_8799);
nand U13645 (N_13645,N_9297,N_7697);
or U13646 (N_13646,N_8405,N_8765);
and U13647 (N_13647,N_5146,N_7065);
and U13648 (N_13648,N_8803,N_7601);
nand U13649 (N_13649,N_9467,N_9678);
nor U13650 (N_13650,N_9672,N_8089);
or U13651 (N_13651,N_7331,N_6589);
and U13652 (N_13652,N_9187,N_5917);
nand U13653 (N_13653,N_8527,N_9590);
and U13654 (N_13654,N_8481,N_8277);
or U13655 (N_13655,N_6385,N_5169);
or U13656 (N_13656,N_8756,N_6499);
nand U13657 (N_13657,N_9453,N_5750);
nand U13658 (N_13658,N_5512,N_5457);
nor U13659 (N_13659,N_6328,N_6576);
or U13660 (N_13660,N_5217,N_5120);
nor U13661 (N_13661,N_7795,N_7842);
or U13662 (N_13662,N_5387,N_5050);
nor U13663 (N_13663,N_7755,N_5038);
and U13664 (N_13664,N_9877,N_5049);
and U13665 (N_13665,N_8403,N_7798);
and U13666 (N_13666,N_6104,N_9357);
nand U13667 (N_13667,N_8013,N_6373);
nand U13668 (N_13668,N_7029,N_7455);
nor U13669 (N_13669,N_8474,N_8043);
nand U13670 (N_13670,N_7679,N_7199);
nor U13671 (N_13671,N_6227,N_6360);
and U13672 (N_13672,N_8704,N_8795);
nor U13673 (N_13673,N_8810,N_8791);
nor U13674 (N_13674,N_5830,N_8236);
and U13675 (N_13675,N_9206,N_9879);
and U13676 (N_13676,N_8605,N_6397);
or U13677 (N_13677,N_5059,N_7287);
nand U13678 (N_13678,N_7699,N_7503);
nor U13679 (N_13679,N_8812,N_6737);
and U13680 (N_13680,N_9064,N_5683);
or U13681 (N_13681,N_9565,N_5451);
and U13682 (N_13682,N_8896,N_8638);
or U13683 (N_13683,N_8393,N_5159);
or U13684 (N_13684,N_5582,N_9201);
and U13685 (N_13685,N_5010,N_9694);
nand U13686 (N_13686,N_8119,N_5656);
nand U13687 (N_13687,N_8806,N_9169);
nand U13688 (N_13688,N_8210,N_5410);
or U13689 (N_13689,N_6701,N_5825);
nor U13690 (N_13690,N_7925,N_7628);
or U13691 (N_13691,N_9637,N_9908);
nor U13692 (N_13692,N_7443,N_8301);
nor U13693 (N_13693,N_8501,N_7797);
or U13694 (N_13694,N_9007,N_8558);
and U13695 (N_13695,N_5218,N_5972);
and U13696 (N_13696,N_6952,N_5314);
and U13697 (N_13697,N_8226,N_9440);
and U13698 (N_13698,N_6204,N_7227);
or U13699 (N_13699,N_6467,N_7602);
and U13700 (N_13700,N_9285,N_8261);
nor U13701 (N_13701,N_7982,N_5158);
or U13702 (N_13702,N_8951,N_5070);
and U13703 (N_13703,N_6174,N_9833);
nor U13704 (N_13704,N_9914,N_6195);
or U13705 (N_13705,N_6633,N_5768);
or U13706 (N_13706,N_7848,N_5426);
or U13707 (N_13707,N_5576,N_7041);
or U13708 (N_13708,N_8614,N_8339);
nor U13709 (N_13709,N_7123,N_5367);
or U13710 (N_13710,N_9208,N_6594);
or U13711 (N_13711,N_6421,N_5432);
nand U13712 (N_13712,N_8172,N_9323);
nor U13713 (N_13713,N_6797,N_9960);
nand U13714 (N_13714,N_7266,N_8996);
or U13715 (N_13715,N_5466,N_9418);
nand U13716 (N_13716,N_7248,N_5272);
and U13717 (N_13717,N_5229,N_8072);
nor U13718 (N_13718,N_5151,N_9455);
or U13719 (N_13719,N_9335,N_8423);
and U13720 (N_13720,N_7071,N_9199);
nand U13721 (N_13721,N_7196,N_5743);
nor U13722 (N_13722,N_5725,N_9756);
or U13723 (N_13723,N_9070,N_9709);
and U13724 (N_13724,N_9852,N_7388);
and U13725 (N_13725,N_9737,N_6110);
nor U13726 (N_13726,N_5679,N_5438);
nand U13727 (N_13727,N_5653,N_5169);
and U13728 (N_13728,N_6579,N_9240);
and U13729 (N_13729,N_6650,N_5639);
nor U13730 (N_13730,N_8172,N_6664);
and U13731 (N_13731,N_8085,N_9369);
or U13732 (N_13732,N_7584,N_8135);
nor U13733 (N_13733,N_8706,N_8199);
and U13734 (N_13734,N_9255,N_9495);
and U13735 (N_13735,N_6199,N_9887);
or U13736 (N_13736,N_7350,N_8365);
nor U13737 (N_13737,N_6649,N_7102);
nand U13738 (N_13738,N_6525,N_6381);
or U13739 (N_13739,N_5436,N_6048);
nor U13740 (N_13740,N_9823,N_6184);
nand U13741 (N_13741,N_9922,N_6371);
nand U13742 (N_13742,N_9706,N_7420);
nand U13743 (N_13743,N_6058,N_6896);
nand U13744 (N_13744,N_7444,N_6101);
nor U13745 (N_13745,N_6048,N_6435);
or U13746 (N_13746,N_8626,N_8953);
or U13747 (N_13747,N_5040,N_6398);
or U13748 (N_13748,N_8815,N_8060);
nor U13749 (N_13749,N_7750,N_5799);
nand U13750 (N_13750,N_9083,N_6843);
nand U13751 (N_13751,N_6074,N_8693);
and U13752 (N_13752,N_7324,N_9001);
or U13753 (N_13753,N_5453,N_9231);
xnor U13754 (N_13754,N_9904,N_5469);
or U13755 (N_13755,N_6109,N_8038);
nand U13756 (N_13756,N_8507,N_5084);
nor U13757 (N_13757,N_6471,N_5427);
nand U13758 (N_13758,N_6412,N_9266);
nor U13759 (N_13759,N_5607,N_8096);
or U13760 (N_13760,N_6913,N_5433);
nand U13761 (N_13761,N_8394,N_7692);
nor U13762 (N_13762,N_7583,N_6227);
and U13763 (N_13763,N_6502,N_6532);
nand U13764 (N_13764,N_5125,N_7483);
nor U13765 (N_13765,N_5902,N_6997);
and U13766 (N_13766,N_5681,N_9301);
nand U13767 (N_13767,N_7441,N_7767);
nor U13768 (N_13768,N_9002,N_5509);
nor U13769 (N_13769,N_9885,N_5838);
or U13770 (N_13770,N_5567,N_8156);
nor U13771 (N_13771,N_8333,N_5134);
and U13772 (N_13772,N_6311,N_5768);
nand U13773 (N_13773,N_7758,N_5094);
nand U13774 (N_13774,N_7382,N_9816);
and U13775 (N_13775,N_6825,N_7272);
nor U13776 (N_13776,N_7819,N_5474);
nor U13777 (N_13777,N_5266,N_9073);
nor U13778 (N_13778,N_9770,N_8724);
or U13779 (N_13779,N_5021,N_9660);
or U13780 (N_13780,N_7998,N_7620);
nand U13781 (N_13781,N_5357,N_8966);
or U13782 (N_13782,N_9221,N_5401);
nand U13783 (N_13783,N_6275,N_7745);
and U13784 (N_13784,N_8910,N_5074);
or U13785 (N_13785,N_6214,N_6786);
or U13786 (N_13786,N_7598,N_5294);
or U13787 (N_13787,N_8966,N_7086);
and U13788 (N_13788,N_9461,N_7588);
nor U13789 (N_13789,N_8764,N_9837);
and U13790 (N_13790,N_7832,N_5287);
nand U13791 (N_13791,N_5620,N_6639);
and U13792 (N_13792,N_9211,N_5026);
nor U13793 (N_13793,N_9517,N_8066);
or U13794 (N_13794,N_6834,N_7376);
nor U13795 (N_13795,N_9806,N_9810);
nor U13796 (N_13796,N_5929,N_8494);
or U13797 (N_13797,N_7993,N_6935);
and U13798 (N_13798,N_8834,N_5565);
or U13799 (N_13799,N_5042,N_9393);
nand U13800 (N_13800,N_8865,N_8382);
or U13801 (N_13801,N_9214,N_6673);
or U13802 (N_13802,N_6772,N_6992);
and U13803 (N_13803,N_5472,N_8734);
nand U13804 (N_13804,N_8515,N_7215);
and U13805 (N_13805,N_5056,N_6843);
or U13806 (N_13806,N_7750,N_6330);
or U13807 (N_13807,N_7491,N_9566);
nor U13808 (N_13808,N_9435,N_8596);
or U13809 (N_13809,N_9486,N_6643);
and U13810 (N_13810,N_6140,N_9400);
or U13811 (N_13811,N_8372,N_6855);
or U13812 (N_13812,N_6104,N_8951);
or U13813 (N_13813,N_5371,N_5149);
or U13814 (N_13814,N_6384,N_7637);
or U13815 (N_13815,N_7834,N_7197);
nor U13816 (N_13816,N_6351,N_8668);
nor U13817 (N_13817,N_8432,N_6149);
xnor U13818 (N_13818,N_5381,N_5597);
or U13819 (N_13819,N_9755,N_7149);
nor U13820 (N_13820,N_9165,N_7144);
nor U13821 (N_13821,N_5591,N_6166);
or U13822 (N_13822,N_9533,N_6808);
nand U13823 (N_13823,N_8374,N_7296);
xnor U13824 (N_13824,N_9617,N_7287);
nor U13825 (N_13825,N_6422,N_6787);
and U13826 (N_13826,N_7350,N_9711);
and U13827 (N_13827,N_8493,N_6184);
and U13828 (N_13828,N_5812,N_5745);
or U13829 (N_13829,N_7594,N_7275);
nor U13830 (N_13830,N_7555,N_5059);
nor U13831 (N_13831,N_6368,N_5464);
nand U13832 (N_13832,N_5325,N_9185);
xnor U13833 (N_13833,N_8612,N_7456);
nor U13834 (N_13834,N_8750,N_8517);
and U13835 (N_13835,N_8236,N_8998);
nor U13836 (N_13836,N_6764,N_9772);
or U13837 (N_13837,N_6710,N_7097);
or U13838 (N_13838,N_9254,N_7200);
or U13839 (N_13839,N_8071,N_5437);
or U13840 (N_13840,N_8795,N_6353);
nand U13841 (N_13841,N_7132,N_5499);
nand U13842 (N_13842,N_7557,N_5529);
and U13843 (N_13843,N_7448,N_7997);
and U13844 (N_13844,N_8668,N_9102);
and U13845 (N_13845,N_7354,N_8295);
and U13846 (N_13846,N_8928,N_6667);
and U13847 (N_13847,N_8718,N_7369);
nand U13848 (N_13848,N_5589,N_9495);
nand U13849 (N_13849,N_9103,N_5056);
and U13850 (N_13850,N_8225,N_6355);
and U13851 (N_13851,N_8643,N_6333);
and U13852 (N_13852,N_7501,N_7923);
or U13853 (N_13853,N_6995,N_6973);
xnor U13854 (N_13854,N_9962,N_7842);
or U13855 (N_13855,N_8784,N_9444);
nand U13856 (N_13856,N_7648,N_8931);
nand U13857 (N_13857,N_9489,N_6178);
and U13858 (N_13858,N_6679,N_8251);
or U13859 (N_13859,N_6603,N_7280);
or U13860 (N_13860,N_9474,N_6730);
and U13861 (N_13861,N_5893,N_7879);
nand U13862 (N_13862,N_7528,N_8124);
or U13863 (N_13863,N_6763,N_5875);
or U13864 (N_13864,N_8828,N_9781);
or U13865 (N_13865,N_6858,N_7302);
and U13866 (N_13866,N_7162,N_8047);
nor U13867 (N_13867,N_7934,N_9416);
and U13868 (N_13868,N_5695,N_8194);
and U13869 (N_13869,N_6737,N_7326);
or U13870 (N_13870,N_9127,N_7247);
nand U13871 (N_13871,N_9851,N_6265);
or U13872 (N_13872,N_7173,N_5583);
nand U13873 (N_13873,N_9974,N_7535);
xnor U13874 (N_13874,N_5333,N_5582);
nand U13875 (N_13875,N_9178,N_5550);
or U13876 (N_13876,N_5844,N_9217);
nand U13877 (N_13877,N_9719,N_7787);
or U13878 (N_13878,N_9045,N_5365);
and U13879 (N_13879,N_6373,N_9047);
nand U13880 (N_13880,N_6552,N_6882);
nor U13881 (N_13881,N_9277,N_7047);
nand U13882 (N_13882,N_5793,N_5509);
or U13883 (N_13883,N_5371,N_8473);
or U13884 (N_13884,N_5237,N_5041);
nand U13885 (N_13885,N_9864,N_6888);
or U13886 (N_13886,N_5351,N_7042);
or U13887 (N_13887,N_9157,N_6930);
nand U13888 (N_13888,N_9746,N_8938);
or U13889 (N_13889,N_9117,N_9221);
nor U13890 (N_13890,N_6845,N_5903);
or U13891 (N_13891,N_7545,N_6575);
or U13892 (N_13892,N_5650,N_6481);
nand U13893 (N_13893,N_9354,N_8994);
nand U13894 (N_13894,N_9190,N_5249);
nand U13895 (N_13895,N_8106,N_5907);
or U13896 (N_13896,N_6611,N_7020);
nor U13897 (N_13897,N_7956,N_7720);
nor U13898 (N_13898,N_5997,N_8352);
or U13899 (N_13899,N_9484,N_5030);
nand U13900 (N_13900,N_8079,N_9965);
xor U13901 (N_13901,N_7970,N_5603);
nand U13902 (N_13902,N_7755,N_9453);
or U13903 (N_13903,N_7219,N_7231);
or U13904 (N_13904,N_6335,N_5401);
and U13905 (N_13905,N_7631,N_8950);
or U13906 (N_13906,N_7998,N_5212);
or U13907 (N_13907,N_7617,N_5259);
nor U13908 (N_13908,N_6811,N_8628);
nor U13909 (N_13909,N_6241,N_6981);
or U13910 (N_13910,N_6753,N_6804);
or U13911 (N_13911,N_9275,N_5134);
nor U13912 (N_13912,N_8179,N_5903);
or U13913 (N_13913,N_9240,N_9363);
nor U13914 (N_13914,N_5627,N_8502);
nor U13915 (N_13915,N_7567,N_5662);
nor U13916 (N_13916,N_7660,N_5053);
nand U13917 (N_13917,N_8558,N_6362);
or U13918 (N_13918,N_6552,N_6453);
nand U13919 (N_13919,N_9621,N_9401);
nand U13920 (N_13920,N_6375,N_5286);
nand U13921 (N_13921,N_8360,N_7857);
and U13922 (N_13922,N_7610,N_5837);
or U13923 (N_13923,N_7840,N_5586);
or U13924 (N_13924,N_9815,N_5374);
nand U13925 (N_13925,N_6500,N_5726);
nand U13926 (N_13926,N_9217,N_9171);
nand U13927 (N_13927,N_5846,N_9854);
or U13928 (N_13928,N_9660,N_5985);
and U13929 (N_13929,N_5146,N_9021);
nor U13930 (N_13930,N_8860,N_6955);
and U13931 (N_13931,N_7172,N_6049);
nand U13932 (N_13932,N_7270,N_6653);
and U13933 (N_13933,N_6610,N_8936);
nor U13934 (N_13934,N_6943,N_5973);
nor U13935 (N_13935,N_5395,N_7021);
nand U13936 (N_13936,N_7283,N_5242);
nor U13937 (N_13937,N_7667,N_8081);
or U13938 (N_13938,N_6642,N_7488);
xnor U13939 (N_13939,N_7872,N_5554);
or U13940 (N_13940,N_7615,N_5435);
or U13941 (N_13941,N_5436,N_5024);
or U13942 (N_13942,N_6419,N_9783);
nand U13943 (N_13943,N_5418,N_5364);
nor U13944 (N_13944,N_5085,N_6638);
and U13945 (N_13945,N_7174,N_8354);
and U13946 (N_13946,N_9208,N_8152);
or U13947 (N_13947,N_9680,N_8734);
nand U13948 (N_13948,N_7218,N_7167);
nor U13949 (N_13949,N_7706,N_6486);
xor U13950 (N_13950,N_6406,N_9893);
nor U13951 (N_13951,N_8707,N_9341);
nand U13952 (N_13952,N_6221,N_8426);
nand U13953 (N_13953,N_6333,N_9444);
nor U13954 (N_13954,N_8420,N_9661);
nor U13955 (N_13955,N_6490,N_7225);
or U13956 (N_13956,N_8523,N_7590);
nor U13957 (N_13957,N_5919,N_7466);
nor U13958 (N_13958,N_9747,N_7922);
nor U13959 (N_13959,N_8837,N_5798);
nand U13960 (N_13960,N_5837,N_7093);
or U13961 (N_13961,N_8061,N_9224);
or U13962 (N_13962,N_6706,N_8811);
and U13963 (N_13963,N_8243,N_6469);
nor U13964 (N_13964,N_7112,N_8591);
nor U13965 (N_13965,N_7683,N_8591);
and U13966 (N_13966,N_6952,N_6676);
nor U13967 (N_13967,N_6774,N_7747);
nand U13968 (N_13968,N_7096,N_9297);
or U13969 (N_13969,N_7400,N_8469);
or U13970 (N_13970,N_9205,N_7287);
nor U13971 (N_13971,N_6253,N_6306);
nor U13972 (N_13972,N_9130,N_6787);
and U13973 (N_13973,N_5188,N_9708);
nand U13974 (N_13974,N_8193,N_5028);
nor U13975 (N_13975,N_5018,N_5246);
or U13976 (N_13976,N_9032,N_6429);
and U13977 (N_13977,N_6147,N_6566);
or U13978 (N_13978,N_8924,N_8525);
nor U13979 (N_13979,N_8833,N_9164);
or U13980 (N_13980,N_8526,N_6103);
nand U13981 (N_13981,N_7706,N_8120);
nor U13982 (N_13982,N_5660,N_8827);
nand U13983 (N_13983,N_7771,N_9800);
nor U13984 (N_13984,N_9720,N_8586);
nor U13985 (N_13985,N_6132,N_9109);
nand U13986 (N_13986,N_8288,N_9405);
nor U13987 (N_13987,N_6195,N_7815);
nand U13988 (N_13988,N_7355,N_7715);
nor U13989 (N_13989,N_8621,N_5032);
nor U13990 (N_13990,N_7984,N_6192);
and U13991 (N_13991,N_8361,N_7336);
nor U13992 (N_13992,N_7162,N_6682);
nor U13993 (N_13993,N_8046,N_7035);
and U13994 (N_13994,N_6211,N_7650);
or U13995 (N_13995,N_6491,N_5702);
nand U13996 (N_13996,N_8656,N_9345);
xnor U13997 (N_13997,N_6139,N_6588);
nor U13998 (N_13998,N_5898,N_6389);
or U13999 (N_13999,N_9011,N_6180);
nor U14000 (N_14000,N_9494,N_7342);
nand U14001 (N_14001,N_9545,N_7935);
nand U14002 (N_14002,N_6123,N_6658);
or U14003 (N_14003,N_8734,N_7495);
or U14004 (N_14004,N_6021,N_9270);
nor U14005 (N_14005,N_6042,N_9833);
or U14006 (N_14006,N_6124,N_9572);
nand U14007 (N_14007,N_8034,N_9469);
and U14008 (N_14008,N_8219,N_6358);
or U14009 (N_14009,N_6583,N_8030);
and U14010 (N_14010,N_9081,N_9149);
and U14011 (N_14011,N_5092,N_9695);
and U14012 (N_14012,N_7768,N_5517);
and U14013 (N_14013,N_5752,N_9129);
nor U14014 (N_14014,N_8920,N_8420);
or U14015 (N_14015,N_7120,N_6278);
or U14016 (N_14016,N_8121,N_6430);
or U14017 (N_14017,N_6326,N_7616);
or U14018 (N_14018,N_5580,N_6622);
and U14019 (N_14019,N_8050,N_6440);
nand U14020 (N_14020,N_8851,N_7740);
nand U14021 (N_14021,N_7606,N_9441);
nor U14022 (N_14022,N_6684,N_8319);
and U14023 (N_14023,N_7987,N_5558);
and U14024 (N_14024,N_8893,N_7097);
and U14025 (N_14025,N_9199,N_9593);
and U14026 (N_14026,N_9954,N_7200);
nand U14027 (N_14027,N_6025,N_5047);
and U14028 (N_14028,N_7483,N_6482);
nand U14029 (N_14029,N_6563,N_7964);
nand U14030 (N_14030,N_7521,N_6631);
or U14031 (N_14031,N_7198,N_5982);
and U14032 (N_14032,N_8916,N_6062);
or U14033 (N_14033,N_6284,N_9162);
nand U14034 (N_14034,N_7315,N_6925);
and U14035 (N_14035,N_7902,N_7582);
nor U14036 (N_14036,N_6473,N_8338);
or U14037 (N_14037,N_8114,N_5746);
or U14038 (N_14038,N_8188,N_9569);
nor U14039 (N_14039,N_9366,N_9000);
nand U14040 (N_14040,N_8385,N_6966);
or U14041 (N_14041,N_7163,N_9452);
and U14042 (N_14042,N_5573,N_8816);
nand U14043 (N_14043,N_9895,N_7930);
nor U14044 (N_14044,N_8062,N_7076);
nand U14045 (N_14045,N_7677,N_6804);
nand U14046 (N_14046,N_9597,N_6358);
and U14047 (N_14047,N_8694,N_5019);
nor U14048 (N_14048,N_6914,N_6274);
and U14049 (N_14049,N_5113,N_9106);
nor U14050 (N_14050,N_9279,N_9192);
and U14051 (N_14051,N_8644,N_9200);
and U14052 (N_14052,N_9555,N_9631);
and U14053 (N_14053,N_8452,N_8188);
or U14054 (N_14054,N_9502,N_5144);
and U14055 (N_14055,N_7515,N_5398);
nand U14056 (N_14056,N_6659,N_7538);
and U14057 (N_14057,N_5604,N_7301);
or U14058 (N_14058,N_7499,N_8707);
or U14059 (N_14059,N_7266,N_8659);
or U14060 (N_14060,N_6427,N_5751);
nand U14061 (N_14061,N_5046,N_9801);
nand U14062 (N_14062,N_6357,N_9336);
and U14063 (N_14063,N_8784,N_9182);
nor U14064 (N_14064,N_5892,N_8597);
or U14065 (N_14065,N_8543,N_6968);
nand U14066 (N_14066,N_7469,N_7680);
nand U14067 (N_14067,N_8203,N_9938);
nand U14068 (N_14068,N_7671,N_9112);
or U14069 (N_14069,N_6106,N_6936);
and U14070 (N_14070,N_9335,N_5268);
nor U14071 (N_14071,N_9133,N_9132);
or U14072 (N_14072,N_6641,N_6445);
or U14073 (N_14073,N_8032,N_6931);
and U14074 (N_14074,N_8354,N_7879);
nand U14075 (N_14075,N_8725,N_6474);
nor U14076 (N_14076,N_7285,N_7177);
nor U14077 (N_14077,N_7821,N_5022);
or U14078 (N_14078,N_7704,N_8836);
or U14079 (N_14079,N_7586,N_8452);
or U14080 (N_14080,N_8731,N_7303);
nand U14081 (N_14081,N_9532,N_5337);
and U14082 (N_14082,N_9320,N_7072);
and U14083 (N_14083,N_8893,N_8079);
and U14084 (N_14084,N_9211,N_6607);
and U14085 (N_14085,N_5388,N_7347);
and U14086 (N_14086,N_9940,N_6888);
nand U14087 (N_14087,N_9446,N_6396);
nor U14088 (N_14088,N_9464,N_5449);
and U14089 (N_14089,N_7324,N_9120);
and U14090 (N_14090,N_6845,N_5087);
nor U14091 (N_14091,N_8778,N_7137);
and U14092 (N_14092,N_9167,N_8436);
nor U14093 (N_14093,N_7417,N_7927);
nor U14094 (N_14094,N_9314,N_8928);
nor U14095 (N_14095,N_9360,N_9353);
and U14096 (N_14096,N_5670,N_7770);
and U14097 (N_14097,N_6559,N_5562);
or U14098 (N_14098,N_5898,N_8479);
and U14099 (N_14099,N_8399,N_9837);
nand U14100 (N_14100,N_8185,N_8058);
nand U14101 (N_14101,N_9135,N_7094);
nor U14102 (N_14102,N_5783,N_8588);
or U14103 (N_14103,N_6730,N_7607);
and U14104 (N_14104,N_9663,N_7885);
or U14105 (N_14105,N_5784,N_9042);
and U14106 (N_14106,N_7831,N_6988);
nor U14107 (N_14107,N_5050,N_5344);
nor U14108 (N_14108,N_6259,N_5405);
and U14109 (N_14109,N_7077,N_8814);
nand U14110 (N_14110,N_7283,N_5929);
nand U14111 (N_14111,N_8169,N_5325);
nand U14112 (N_14112,N_6475,N_7665);
nand U14113 (N_14113,N_8295,N_6336);
nand U14114 (N_14114,N_8930,N_6209);
and U14115 (N_14115,N_6684,N_7069);
and U14116 (N_14116,N_6467,N_5836);
nand U14117 (N_14117,N_6484,N_6650);
nand U14118 (N_14118,N_5394,N_9708);
or U14119 (N_14119,N_7925,N_9728);
nand U14120 (N_14120,N_9530,N_8888);
or U14121 (N_14121,N_9378,N_7181);
nand U14122 (N_14122,N_7451,N_9987);
nand U14123 (N_14123,N_5770,N_6113);
or U14124 (N_14124,N_5958,N_9069);
and U14125 (N_14125,N_6314,N_8440);
and U14126 (N_14126,N_7471,N_8290);
xor U14127 (N_14127,N_6592,N_5280);
nand U14128 (N_14128,N_8114,N_8451);
and U14129 (N_14129,N_8457,N_7469);
nor U14130 (N_14130,N_6472,N_8073);
xor U14131 (N_14131,N_9552,N_9188);
nor U14132 (N_14132,N_8604,N_6410);
nand U14133 (N_14133,N_8599,N_5481);
nand U14134 (N_14134,N_7830,N_7339);
or U14135 (N_14135,N_7171,N_9134);
or U14136 (N_14136,N_8447,N_8673);
nand U14137 (N_14137,N_6722,N_5619);
and U14138 (N_14138,N_7576,N_6040);
or U14139 (N_14139,N_8478,N_8504);
nor U14140 (N_14140,N_9937,N_7132);
or U14141 (N_14141,N_6210,N_7100);
nor U14142 (N_14142,N_8616,N_7067);
nand U14143 (N_14143,N_6650,N_6906);
and U14144 (N_14144,N_9536,N_9700);
nand U14145 (N_14145,N_5065,N_6047);
nand U14146 (N_14146,N_7702,N_7488);
nand U14147 (N_14147,N_5223,N_8734);
or U14148 (N_14148,N_5885,N_9890);
and U14149 (N_14149,N_9519,N_7634);
nor U14150 (N_14150,N_6004,N_7888);
nor U14151 (N_14151,N_5141,N_8060);
nand U14152 (N_14152,N_7140,N_9516);
nand U14153 (N_14153,N_6892,N_9640);
or U14154 (N_14154,N_7418,N_8780);
nand U14155 (N_14155,N_5215,N_6316);
or U14156 (N_14156,N_7273,N_8496);
nand U14157 (N_14157,N_6126,N_7710);
and U14158 (N_14158,N_9604,N_7831);
nor U14159 (N_14159,N_7902,N_5135);
nand U14160 (N_14160,N_5969,N_9563);
nor U14161 (N_14161,N_7730,N_9563);
xor U14162 (N_14162,N_8036,N_5858);
and U14163 (N_14163,N_7457,N_7669);
xor U14164 (N_14164,N_5881,N_8251);
nand U14165 (N_14165,N_7429,N_8449);
or U14166 (N_14166,N_7541,N_6355);
and U14167 (N_14167,N_5282,N_5827);
xor U14168 (N_14168,N_8644,N_8632);
nand U14169 (N_14169,N_8895,N_5754);
nor U14170 (N_14170,N_7963,N_8373);
nor U14171 (N_14171,N_7804,N_9471);
nand U14172 (N_14172,N_7930,N_9908);
or U14173 (N_14173,N_8441,N_9957);
and U14174 (N_14174,N_7858,N_7841);
or U14175 (N_14175,N_5676,N_6788);
and U14176 (N_14176,N_8287,N_6196);
nand U14177 (N_14177,N_5525,N_9060);
nor U14178 (N_14178,N_7489,N_6673);
nor U14179 (N_14179,N_8997,N_6198);
xnor U14180 (N_14180,N_5953,N_7557);
and U14181 (N_14181,N_6081,N_6460);
or U14182 (N_14182,N_8539,N_7096);
nor U14183 (N_14183,N_6524,N_5545);
or U14184 (N_14184,N_7305,N_7057);
and U14185 (N_14185,N_9639,N_5621);
and U14186 (N_14186,N_7937,N_5164);
and U14187 (N_14187,N_6781,N_7665);
nand U14188 (N_14188,N_6047,N_5711);
nand U14189 (N_14189,N_7312,N_9164);
nor U14190 (N_14190,N_5725,N_7177);
and U14191 (N_14191,N_5320,N_5248);
nand U14192 (N_14192,N_8062,N_7840);
nand U14193 (N_14193,N_6722,N_6314);
nand U14194 (N_14194,N_6817,N_8240);
nor U14195 (N_14195,N_7070,N_6894);
and U14196 (N_14196,N_7004,N_5976);
nor U14197 (N_14197,N_5977,N_7507);
nor U14198 (N_14198,N_5682,N_5699);
nand U14199 (N_14199,N_5198,N_7793);
or U14200 (N_14200,N_5143,N_5185);
nand U14201 (N_14201,N_5163,N_6054);
nand U14202 (N_14202,N_6930,N_9877);
or U14203 (N_14203,N_7579,N_9510);
and U14204 (N_14204,N_5623,N_6097);
or U14205 (N_14205,N_7150,N_5782);
or U14206 (N_14206,N_8747,N_7058);
nor U14207 (N_14207,N_7986,N_6243);
nand U14208 (N_14208,N_5421,N_8286);
nor U14209 (N_14209,N_8236,N_5691);
nand U14210 (N_14210,N_6728,N_9287);
or U14211 (N_14211,N_5077,N_6086);
nand U14212 (N_14212,N_7476,N_6147);
or U14213 (N_14213,N_5552,N_9992);
nand U14214 (N_14214,N_6223,N_7631);
nor U14215 (N_14215,N_6819,N_9784);
or U14216 (N_14216,N_5009,N_7336);
xor U14217 (N_14217,N_9900,N_9895);
and U14218 (N_14218,N_5780,N_9018);
nand U14219 (N_14219,N_9803,N_9064);
nand U14220 (N_14220,N_5206,N_5056);
nor U14221 (N_14221,N_9951,N_6162);
or U14222 (N_14222,N_9872,N_7220);
and U14223 (N_14223,N_5139,N_5574);
and U14224 (N_14224,N_5339,N_8935);
nor U14225 (N_14225,N_9082,N_5044);
nor U14226 (N_14226,N_8318,N_6355);
and U14227 (N_14227,N_9758,N_8551);
and U14228 (N_14228,N_8564,N_6384);
or U14229 (N_14229,N_5965,N_7806);
nand U14230 (N_14230,N_8380,N_8755);
nor U14231 (N_14231,N_8543,N_5688);
nand U14232 (N_14232,N_7183,N_8861);
nand U14233 (N_14233,N_9498,N_7508);
nor U14234 (N_14234,N_9553,N_9698);
and U14235 (N_14235,N_8715,N_7952);
or U14236 (N_14236,N_5694,N_9818);
or U14237 (N_14237,N_6093,N_7099);
nand U14238 (N_14238,N_5296,N_7611);
nor U14239 (N_14239,N_6305,N_6484);
nor U14240 (N_14240,N_9965,N_6394);
and U14241 (N_14241,N_9113,N_6660);
or U14242 (N_14242,N_6788,N_6176);
or U14243 (N_14243,N_7768,N_5047);
nor U14244 (N_14244,N_7725,N_5500);
and U14245 (N_14245,N_5005,N_8193);
nand U14246 (N_14246,N_8614,N_9223);
or U14247 (N_14247,N_9722,N_8032);
nor U14248 (N_14248,N_5664,N_5106);
and U14249 (N_14249,N_7812,N_9549);
nand U14250 (N_14250,N_9137,N_6744);
nand U14251 (N_14251,N_5815,N_9681);
or U14252 (N_14252,N_9477,N_9282);
or U14253 (N_14253,N_5182,N_6629);
or U14254 (N_14254,N_9132,N_7113);
nand U14255 (N_14255,N_6895,N_8401);
nand U14256 (N_14256,N_7536,N_8180);
nor U14257 (N_14257,N_5255,N_7959);
nor U14258 (N_14258,N_7664,N_5557);
and U14259 (N_14259,N_8673,N_8179);
nor U14260 (N_14260,N_7802,N_9617);
nand U14261 (N_14261,N_6399,N_8550);
nor U14262 (N_14262,N_5260,N_6167);
nor U14263 (N_14263,N_9490,N_7279);
nor U14264 (N_14264,N_9452,N_6465);
or U14265 (N_14265,N_7720,N_5448);
nand U14266 (N_14266,N_8316,N_6641);
and U14267 (N_14267,N_9057,N_7521);
nor U14268 (N_14268,N_6807,N_5000);
and U14269 (N_14269,N_7749,N_5259);
or U14270 (N_14270,N_9492,N_5058);
nand U14271 (N_14271,N_5769,N_5921);
nor U14272 (N_14272,N_8288,N_5021);
nand U14273 (N_14273,N_7580,N_6428);
nand U14274 (N_14274,N_9988,N_7099);
or U14275 (N_14275,N_5639,N_5001);
and U14276 (N_14276,N_6603,N_8090);
and U14277 (N_14277,N_9811,N_8747);
and U14278 (N_14278,N_8065,N_8950);
nor U14279 (N_14279,N_8689,N_7410);
or U14280 (N_14280,N_9163,N_9637);
nor U14281 (N_14281,N_6843,N_5849);
and U14282 (N_14282,N_5676,N_9061);
nor U14283 (N_14283,N_6715,N_7334);
and U14284 (N_14284,N_8415,N_7074);
and U14285 (N_14285,N_7569,N_7043);
and U14286 (N_14286,N_8795,N_9915);
or U14287 (N_14287,N_7499,N_9990);
nand U14288 (N_14288,N_9555,N_5339);
and U14289 (N_14289,N_8359,N_8920);
xnor U14290 (N_14290,N_6216,N_7955);
nor U14291 (N_14291,N_7984,N_7514);
or U14292 (N_14292,N_6043,N_6431);
nor U14293 (N_14293,N_8873,N_5387);
nor U14294 (N_14294,N_6620,N_9602);
or U14295 (N_14295,N_5777,N_9466);
and U14296 (N_14296,N_7361,N_9610);
nor U14297 (N_14297,N_7058,N_6254);
or U14298 (N_14298,N_6970,N_6404);
nand U14299 (N_14299,N_5224,N_5375);
and U14300 (N_14300,N_6257,N_9348);
nor U14301 (N_14301,N_5977,N_6285);
nor U14302 (N_14302,N_7614,N_5714);
and U14303 (N_14303,N_9642,N_5883);
and U14304 (N_14304,N_8756,N_6010);
nor U14305 (N_14305,N_5279,N_6944);
nor U14306 (N_14306,N_6227,N_9540);
nor U14307 (N_14307,N_8823,N_9422);
and U14308 (N_14308,N_8239,N_5221);
nor U14309 (N_14309,N_8004,N_6836);
or U14310 (N_14310,N_6407,N_9453);
nor U14311 (N_14311,N_8170,N_5061);
or U14312 (N_14312,N_8265,N_7322);
and U14313 (N_14313,N_7252,N_9884);
or U14314 (N_14314,N_5391,N_5491);
nand U14315 (N_14315,N_5093,N_8843);
nor U14316 (N_14316,N_6437,N_8885);
or U14317 (N_14317,N_6870,N_5231);
nand U14318 (N_14318,N_8504,N_7072);
nand U14319 (N_14319,N_8898,N_9762);
nor U14320 (N_14320,N_8946,N_8428);
or U14321 (N_14321,N_8081,N_9705);
nor U14322 (N_14322,N_9553,N_8738);
or U14323 (N_14323,N_6810,N_9486);
nand U14324 (N_14324,N_7902,N_5562);
nor U14325 (N_14325,N_8908,N_9085);
nor U14326 (N_14326,N_9062,N_8639);
nor U14327 (N_14327,N_8982,N_7267);
nand U14328 (N_14328,N_5637,N_7511);
nand U14329 (N_14329,N_9105,N_6361);
and U14330 (N_14330,N_9855,N_6887);
nand U14331 (N_14331,N_9272,N_9084);
xnor U14332 (N_14332,N_9081,N_5957);
and U14333 (N_14333,N_9320,N_5182);
or U14334 (N_14334,N_7781,N_9014);
or U14335 (N_14335,N_6933,N_6755);
or U14336 (N_14336,N_5758,N_8865);
and U14337 (N_14337,N_6534,N_7813);
or U14338 (N_14338,N_9115,N_7250);
nor U14339 (N_14339,N_6379,N_7704);
or U14340 (N_14340,N_7470,N_8456);
xor U14341 (N_14341,N_7470,N_7987);
and U14342 (N_14342,N_6917,N_6270);
nor U14343 (N_14343,N_6864,N_5950);
or U14344 (N_14344,N_6632,N_9159);
and U14345 (N_14345,N_8241,N_9829);
or U14346 (N_14346,N_5020,N_9803);
nand U14347 (N_14347,N_6344,N_9267);
and U14348 (N_14348,N_5001,N_5041);
or U14349 (N_14349,N_5097,N_5186);
nand U14350 (N_14350,N_6048,N_7422);
or U14351 (N_14351,N_5196,N_7768);
and U14352 (N_14352,N_5962,N_6970);
and U14353 (N_14353,N_5123,N_6600);
nand U14354 (N_14354,N_5219,N_7897);
nand U14355 (N_14355,N_8414,N_8337);
and U14356 (N_14356,N_5100,N_5052);
nand U14357 (N_14357,N_8761,N_7595);
nand U14358 (N_14358,N_6754,N_6258);
or U14359 (N_14359,N_8773,N_9567);
xor U14360 (N_14360,N_7621,N_6829);
or U14361 (N_14361,N_8084,N_9640);
nand U14362 (N_14362,N_5033,N_5842);
nand U14363 (N_14363,N_5230,N_8090);
nand U14364 (N_14364,N_6970,N_9231);
and U14365 (N_14365,N_7506,N_6197);
nand U14366 (N_14366,N_8933,N_7285);
nor U14367 (N_14367,N_7449,N_7576);
nand U14368 (N_14368,N_5553,N_8874);
or U14369 (N_14369,N_6474,N_5469);
nor U14370 (N_14370,N_8199,N_6853);
nor U14371 (N_14371,N_5148,N_6204);
nor U14372 (N_14372,N_8816,N_6717);
and U14373 (N_14373,N_9633,N_8257);
and U14374 (N_14374,N_7446,N_7399);
and U14375 (N_14375,N_8684,N_5990);
nand U14376 (N_14376,N_7872,N_7376);
nor U14377 (N_14377,N_5464,N_5490);
nand U14378 (N_14378,N_9971,N_8092);
or U14379 (N_14379,N_9921,N_5863);
or U14380 (N_14380,N_5384,N_7617);
and U14381 (N_14381,N_5163,N_8819);
nand U14382 (N_14382,N_6052,N_7066);
nor U14383 (N_14383,N_7046,N_8555);
nand U14384 (N_14384,N_8168,N_5743);
xnor U14385 (N_14385,N_5505,N_8546);
nand U14386 (N_14386,N_6005,N_6828);
and U14387 (N_14387,N_5864,N_9354);
and U14388 (N_14388,N_7581,N_5183);
nor U14389 (N_14389,N_7139,N_8010);
or U14390 (N_14390,N_7329,N_6064);
or U14391 (N_14391,N_7603,N_9810);
and U14392 (N_14392,N_8923,N_8479);
nand U14393 (N_14393,N_6377,N_8695);
nand U14394 (N_14394,N_9787,N_5707);
nand U14395 (N_14395,N_6544,N_9942);
nand U14396 (N_14396,N_7764,N_9917);
nand U14397 (N_14397,N_9074,N_5244);
nor U14398 (N_14398,N_5697,N_5252);
or U14399 (N_14399,N_5638,N_8804);
or U14400 (N_14400,N_6838,N_8551);
or U14401 (N_14401,N_5618,N_5886);
and U14402 (N_14402,N_7633,N_8732);
nor U14403 (N_14403,N_5202,N_7119);
and U14404 (N_14404,N_5492,N_5015);
or U14405 (N_14405,N_9420,N_8620);
and U14406 (N_14406,N_9391,N_6625);
nor U14407 (N_14407,N_7255,N_8043);
nor U14408 (N_14408,N_7550,N_8004);
nor U14409 (N_14409,N_5632,N_5865);
and U14410 (N_14410,N_6368,N_6299);
nand U14411 (N_14411,N_7714,N_8116);
nand U14412 (N_14412,N_8654,N_9374);
and U14413 (N_14413,N_6788,N_7094);
nor U14414 (N_14414,N_5338,N_7384);
xnor U14415 (N_14415,N_7402,N_6697);
xor U14416 (N_14416,N_5419,N_7693);
or U14417 (N_14417,N_5181,N_5975);
or U14418 (N_14418,N_5242,N_8421);
or U14419 (N_14419,N_6653,N_6149);
or U14420 (N_14420,N_9080,N_8803);
nor U14421 (N_14421,N_6146,N_8154);
and U14422 (N_14422,N_8160,N_9435);
nor U14423 (N_14423,N_5826,N_7293);
or U14424 (N_14424,N_8036,N_5710);
and U14425 (N_14425,N_5475,N_8916);
nand U14426 (N_14426,N_5648,N_6531);
or U14427 (N_14427,N_9336,N_8048);
nor U14428 (N_14428,N_7195,N_9327);
nor U14429 (N_14429,N_8976,N_9359);
and U14430 (N_14430,N_7923,N_9904);
nand U14431 (N_14431,N_5545,N_6224);
or U14432 (N_14432,N_7995,N_8451);
xnor U14433 (N_14433,N_7899,N_8161);
nor U14434 (N_14434,N_6580,N_5083);
nor U14435 (N_14435,N_8806,N_6697);
nand U14436 (N_14436,N_8814,N_7548);
nor U14437 (N_14437,N_7470,N_7721);
or U14438 (N_14438,N_7935,N_7287);
nor U14439 (N_14439,N_6458,N_8387);
or U14440 (N_14440,N_9925,N_8937);
and U14441 (N_14441,N_7091,N_5499);
and U14442 (N_14442,N_8013,N_6032);
nand U14443 (N_14443,N_9474,N_8468);
nor U14444 (N_14444,N_7681,N_9657);
or U14445 (N_14445,N_9016,N_9917);
and U14446 (N_14446,N_7531,N_5743);
nor U14447 (N_14447,N_9608,N_7278);
nor U14448 (N_14448,N_8734,N_6802);
nor U14449 (N_14449,N_7079,N_7868);
nor U14450 (N_14450,N_6689,N_5705);
nor U14451 (N_14451,N_7715,N_6955);
and U14452 (N_14452,N_6551,N_6060);
and U14453 (N_14453,N_6802,N_6551);
nand U14454 (N_14454,N_6815,N_9206);
or U14455 (N_14455,N_5838,N_9772);
or U14456 (N_14456,N_9477,N_8038);
or U14457 (N_14457,N_7264,N_9181);
nand U14458 (N_14458,N_7871,N_8660);
or U14459 (N_14459,N_8660,N_9592);
or U14460 (N_14460,N_6939,N_9383);
and U14461 (N_14461,N_7591,N_6797);
nand U14462 (N_14462,N_7760,N_7872);
nand U14463 (N_14463,N_6371,N_5547);
and U14464 (N_14464,N_8232,N_5461);
or U14465 (N_14465,N_5658,N_7486);
nor U14466 (N_14466,N_8110,N_7504);
and U14467 (N_14467,N_9851,N_6093);
or U14468 (N_14468,N_9003,N_6230);
nand U14469 (N_14469,N_5444,N_7294);
and U14470 (N_14470,N_7866,N_6133);
or U14471 (N_14471,N_8578,N_9493);
nor U14472 (N_14472,N_6690,N_8150);
or U14473 (N_14473,N_8906,N_8258);
nor U14474 (N_14474,N_5727,N_8397);
or U14475 (N_14475,N_7339,N_9709);
and U14476 (N_14476,N_5657,N_5214);
and U14477 (N_14477,N_6991,N_6221);
nor U14478 (N_14478,N_6345,N_7919);
nor U14479 (N_14479,N_5098,N_9857);
and U14480 (N_14480,N_9769,N_8320);
and U14481 (N_14481,N_7205,N_9953);
or U14482 (N_14482,N_8285,N_8307);
nand U14483 (N_14483,N_9932,N_8772);
nand U14484 (N_14484,N_9919,N_7682);
nand U14485 (N_14485,N_7434,N_5263);
xor U14486 (N_14486,N_5145,N_9793);
or U14487 (N_14487,N_8808,N_6899);
nand U14488 (N_14488,N_9017,N_9695);
nor U14489 (N_14489,N_6386,N_8806);
or U14490 (N_14490,N_6569,N_7822);
or U14491 (N_14491,N_5467,N_6744);
nand U14492 (N_14492,N_9751,N_8059);
nor U14493 (N_14493,N_9596,N_5975);
nand U14494 (N_14494,N_7996,N_7905);
or U14495 (N_14495,N_6164,N_7776);
nand U14496 (N_14496,N_5415,N_6750);
xor U14497 (N_14497,N_6912,N_7746);
or U14498 (N_14498,N_7583,N_5170);
and U14499 (N_14499,N_7613,N_7556);
nand U14500 (N_14500,N_9299,N_9209);
nor U14501 (N_14501,N_8734,N_7925);
or U14502 (N_14502,N_5457,N_9856);
or U14503 (N_14503,N_9355,N_5965);
nor U14504 (N_14504,N_8710,N_6313);
or U14505 (N_14505,N_7911,N_7335);
and U14506 (N_14506,N_8367,N_8376);
nand U14507 (N_14507,N_8594,N_5104);
or U14508 (N_14508,N_8513,N_6393);
xor U14509 (N_14509,N_7603,N_8205);
or U14510 (N_14510,N_6442,N_9708);
or U14511 (N_14511,N_9701,N_5641);
or U14512 (N_14512,N_6063,N_8725);
and U14513 (N_14513,N_6068,N_5417);
nand U14514 (N_14514,N_9104,N_7087);
or U14515 (N_14515,N_8184,N_5171);
or U14516 (N_14516,N_8894,N_9180);
and U14517 (N_14517,N_6088,N_8039);
nand U14518 (N_14518,N_8362,N_6986);
nand U14519 (N_14519,N_6606,N_9757);
nor U14520 (N_14520,N_8688,N_5812);
and U14521 (N_14521,N_7501,N_7215);
nor U14522 (N_14522,N_7190,N_6253);
and U14523 (N_14523,N_7972,N_6203);
or U14524 (N_14524,N_9457,N_9451);
and U14525 (N_14525,N_5688,N_5557);
and U14526 (N_14526,N_8178,N_8874);
nand U14527 (N_14527,N_7284,N_9603);
nand U14528 (N_14528,N_5274,N_6669);
or U14529 (N_14529,N_8054,N_9255);
and U14530 (N_14530,N_7645,N_7399);
or U14531 (N_14531,N_5930,N_6586);
nor U14532 (N_14532,N_7949,N_6347);
or U14533 (N_14533,N_7277,N_7824);
nor U14534 (N_14534,N_5889,N_8193);
or U14535 (N_14535,N_7173,N_8544);
xor U14536 (N_14536,N_9922,N_8025);
or U14537 (N_14537,N_9904,N_7034);
or U14538 (N_14538,N_7203,N_6930);
or U14539 (N_14539,N_7614,N_8755);
and U14540 (N_14540,N_5126,N_7421);
or U14541 (N_14541,N_8193,N_7611);
or U14542 (N_14542,N_9897,N_7037);
or U14543 (N_14543,N_8083,N_5106);
or U14544 (N_14544,N_7761,N_6653);
or U14545 (N_14545,N_7013,N_6642);
nand U14546 (N_14546,N_7135,N_7958);
or U14547 (N_14547,N_5730,N_7945);
and U14548 (N_14548,N_7766,N_5554);
and U14549 (N_14549,N_7046,N_8131);
nor U14550 (N_14550,N_9066,N_9805);
xor U14551 (N_14551,N_8555,N_7347);
nand U14552 (N_14552,N_6147,N_8785);
nand U14553 (N_14553,N_5637,N_7276);
xor U14554 (N_14554,N_7338,N_6360);
or U14555 (N_14555,N_8813,N_9251);
nor U14556 (N_14556,N_6326,N_5264);
nand U14557 (N_14557,N_9094,N_5502);
or U14558 (N_14558,N_7668,N_7925);
and U14559 (N_14559,N_7020,N_9232);
nand U14560 (N_14560,N_6245,N_7871);
or U14561 (N_14561,N_5181,N_5284);
nor U14562 (N_14562,N_6096,N_9019);
or U14563 (N_14563,N_7658,N_9975);
nand U14564 (N_14564,N_8071,N_9949);
and U14565 (N_14565,N_7020,N_8548);
and U14566 (N_14566,N_8663,N_5905);
nor U14567 (N_14567,N_9426,N_8692);
or U14568 (N_14568,N_5701,N_9178);
or U14569 (N_14569,N_9779,N_6079);
and U14570 (N_14570,N_7393,N_5551);
nor U14571 (N_14571,N_7782,N_8730);
nor U14572 (N_14572,N_5102,N_7779);
and U14573 (N_14573,N_9992,N_9131);
xor U14574 (N_14574,N_6530,N_9609);
and U14575 (N_14575,N_9306,N_8982);
xor U14576 (N_14576,N_9261,N_7631);
or U14577 (N_14577,N_7289,N_9053);
or U14578 (N_14578,N_6666,N_6194);
nand U14579 (N_14579,N_5363,N_5287);
and U14580 (N_14580,N_6110,N_9583);
or U14581 (N_14581,N_5631,N_8435);
nand U14582 (N_14582,N_8115,N_5636);
nand U14583 (N_14583,N_5841,N_9770);
nand U14584 (N_14584,N_6761,N_5295);
and U14585 (N_14585,N_5065,N_7095);
nand U14586 (N_14586,N_7937,N_7540);
and U14587 (N_14587,N_8578,N_8929);
nor U14588 (N_14588,N_5391,N_9847);
or U14589 (N_14589,N_9309,N_5548);
or U14590 (N_14590,N_6915,N_5878);
nand U14591 (N_14591,N_5132,N_9391);
or U14592 (N_14592,N_6258,N_5505);
xor U14593 (N_14593,N_5424,N_7519);
nor U14594 (N_14594,N_6586,N_7140);
nand U14595 (N_14595,N_6758,N_5542);
nor U14596 (N_14596,N_9096,N_7679);
or U14597 (N_14597,N_9002,N_8002);
and U14598 (N_14598,N_7399,N_9125);
nand U14599 (N_14599,N_6689,N_5734);
and U14600 (N_14600,N_6023,N_6686);
and U14601 (N_14601,N_5865,N_7534);
nand U14602 (N_14602,N_6906,N_9489);
or U14603 (N_14603,N_8740,N_8823);
nor U14604 (N_14604,N_9669,N_9602);
nor U14605 (N_14605,N_9378,N_6515);
or U14606 (N_14606,N_7622,N_7979);
or U14607 (N_14607,N_9318,N_8004);
or U14608 (N_14608,N_9742,N_8140);
nor U14609 (N_14609,N_6186,N_5662);
nand U14610 (N_14610,N_9972,N_6129);
and U14611 (N_14611,N_9063,N_6153);
or U14612 (N_14612,N_8019,N_7544);
or U14613 (N_14613,N_6820,N_8906);
nor U14614 (N_14614,N_8638,N_7400);
nand U14615 (N_14615,N_6652,N_7704);
nand U14616 (N_14616,N_9688,N_7197);
nand U14617 (N_14617,N_6802,N_5908);
or U14618 (N_14618,N_8468,N_8152);
xnor U14619 (N_14619,N_6865,N_6050);
or U14620 (N_14620,N_9782,N_7498);
or U14621 (N_14621,N_8158,N_7104);
nor U14622 (N_14622,N_5690,N_6202);
nand U14623 (N_14623,N_8818,N_8670);
or U14624 (N_14624,N_5723,N_5403);
and U14625 (N_14625,N_8887,N_5020);
nand U14626 (N_14626,N_8272,N_9069);
nor U14627 (N_14627,N_6880,N_6822);
or U14628 (N_14628,N_7778,N_7651);
and U14629 (N_14629,N_7541,N_9714);
nor U14630 (N_14630,N_5886,N_5912);
nand U14631 (N_14631,N_7179,N_7516);
or U14632 (N_14632,N_6014,N_9903);
nor U14633 (N_14633,N_8387,N_5916);
nor U14634 (N_14634,N_9333,N_5114);
or U14635 (N_14635,N_9897,N_9303);
nor U14636 (N_14636,N_8661,N_6737);
or U14637 (N_14637,N_5004,N_7110);
nand U14638 (N_14638,N_8631,N_9343);
or U14639 (N_14639,N_6272,N_8864);
nand U14640 (N_14640,N_6895,N_9447);
xnor U14641 (N_14641,N_9914,N_8954);
or U14642 (N_14642,N_5652,N_6628);
or U14643 (N_14643,N_7534,N_5498);
nand U14644 (N_14644,N_6848,N_9883);
nor U14645 (N_14645,N_7887,N_8497);
and U14646 (N_14646,N_6078,N_6895);
and U14647 (N_14647,N_8701,N_9040);
and U14648 (N_14648,N_7746,N_9088);
nor U14649 (N_14649,N_7216,N_9319);
nor U14650 (N_14650,N_8021,N_9647);
and U14651 (N_14651,N_7978,N_8490);
or U14652 (N_14652,N_7704,N_5496);
and U14653 (N_14653,N_6226,N_8576);
nor U14654 (N_14654,N_7726,N_5619);
or U14655 (N_14655,N_8742,N_9538);
nor U14656 (N_14656,N_9353,N_9804);
or U14657 (N_14657,N_6310,N_9667);
or U14658 (N_14658,N_7090,N_6623);
nor U14659 (N_14659,N_5512,N_5139);
or U14660 (N_14660,N_6133,N_5686);
nor U14661 (N_14661,N_6681,N_5647);
nor U14662 (N_14662,N_5204,N_5793);
and U14663 (N_14663,N_6102,N_9989);
or U14664 (N_14664,N_7483,N_9377);
and U14665 (N_14665,N_8533,N_9363);
xor U14666 (N_14666,N_7409,N_9216);
nand U14667 (N_14667,N_7721,N_6329);
nor U14668 (N_14668,N_5061,N_6270);
nor U14669 (N_14669,N_6694,N_7558);
nand U14670 (N_14670,N_5486,N_9483);
and U14671 (N_14671,N_6855,N_9338);
and U14672 (N_14672,N_5142,N_6300);
and U14673 (N_14673,N_5348,N_8362);
or U14674 (N_14674,N_7400,N_5692);
and U14675 (N_14675,N_5052,N_7251);
nand U14676 (N_14676,N_7250,N_5505);
or U14677 (N_14677,N_6780,N_7023);
nand U14678 (N_14678,N_5438,N_5227);
and U14679 (N_14679,N_5757,N_8680);
nor U14680 (N_14680,N_9214,N_8031);
or U14681 (N_14681,N_5191,N_8377);
and U14682 (N_14682,N_9428,N_7695);
xnor U14683 (N_14683,N_9838,N_8725);
and U14684 (N_14684,N_8327,N_5380);
or U14685 (N_14685,N_8101,N_9288);
or U14686 (N_14686,N_9901,N_7191);
nand U14687 (N_14687,N_6799,N_8000);
nor U14688 (N_14688,N_9000,N_5573);
nand U14689 (N_14689,N_5910,N_5869);
nor U14690 (N_14690,N_5203,N_7072);
or U14691 (N_14691,N_6674,N_5640);
nor U14692 (N_14692,N_5055,N_7213);
nor U14693 (N_14693,N_8899,N_7591);
nand U14694 (N_14694,N_6559,N_5466);
nand U14695 (N_14695,N_6139,N_8897);
and U14696 (N_14696,N_9197,N_7601);
nand U14697 (N_14697,N_6478,N_8627);
or U14698 (N_14698,N_8734,N_8432);
and U14699 (N_14699,N_6794,N_6483);
nor U14700 (N_14700,N_8429,N_5318);
or U14701 (N_14701,N_7788,N_9947);
or U14702 (N_14702,N_8117,N_9336);
and U14703 (N_14703,N_8829,N_5605);
and U14704 (N_14704,N_9990,N_6001);
nand U14705 (N_14705,N_7871,N_7715);
or U14706 (N_14706,N_9708,N_6767);
nor U14707 (N_14707,N_8716,N_9528);
nor U14708 (N_14708,N_8406,N_8723);
and U14709 (N_14709,N_8527,N_6634);
nor U14710 (N_14710,N_8774,N_6260);
and U14711 (N_14711,N_5597,N_6236);
or U14712 (N_14712,N_5814,N_7888);
and U14713 (N_14713,N_7687,N_5798);
nand U14714 (N_14714,N_9975,N_7249);
and U14715 (N_14715,N_6393,N_8750);
or U14716 (N_14716,N_6836,N_9068);
nor U14717 (N_14717,N_8281,N_5458);
nor U14718 (N_14718,N_6216,N_7018);
or U14719 (N_14719,N_6380,N_7384);
and U14720 (N_14720,N_8546,N_8820);
and U14721 (N_14721,N_8485,N_7834);
and U14722 (N_14722,N_6315,N_6741);
or U14723 (N_14723,N_8812,N_6184);
and U14724 (N_14724,N_8164,N_6876);
or U14725 (N_14725,N_9135,N_5034);
and U14726 (N_14726,N_8539,N_5101);
nand U14727 (N_14727,N_9661,N_6580);
and U14728 (N_14728,N_9754,N_9043);
nand U14729 (N_14729,N_7850,N_5660);
and U14730 (N_14730,N_7515,N_7506);
nand U14731 (N_14731,N_8153,N_7968);
and U14732 (N_14732,N_7114,N_9989);
or U14733 (N_14733,N_6918,N_9555);
and U14734 (N_14734,N_5124,N_8238);
or U14735 (N_14735,N_9639,N_5170);
nor U14736 (N_14736,N_7778,N_8045);
or U14737 (N_14737,N_9718,N_7099);
and U14738 (N_14738,N_5541,N_8942);
nor U14739 (N_14739,N_8544,N_8060);
nand U14740 (N_14740,N_5722,N_8873);
nand U14741 (N_14741,N_9869,N_5719);
nor U14742 (N_14742,N_9818,N_8807);
nand U14743 (N_14743,N_6918,N_7810);
and U14744 (N_14744,N_5191,N_8533);
nand U14745 (N_14745,N_6223,N_7447);
or U14746 (N_14746,N_6839,N_5452);
or U14747 (N_14747,N_7102,N_9699);
nand U14748 (N_14748,N_5490,N_7237);
nand U14749 (N_14749,N_5919,N_5442);
or U14750 (N_14750,N_8636,N_8486);
and U14751 (N_14751,N_8188,N_8547);
nor U14752 (N_14752,N_6655,N_6947);
or U14753 (N_14753,N_7763,N_8223);
nand U14754 (N_14754,N_6166,N_7412);
nor U14755 (N_14755,N_5016,N_5214);
xor U14756 (N_14756,N_6136,N_7995);
or U14757 (N_14757,N_9293,N_8094);
nor U14758 (N_14758,N_9542,N_8857);
xnor U14759 (N_14759,N_7906,N_6033);
nand U14760 (N_14760,N_8026,N_9992);
nand U14761 (N_14761,N_5704,N_9831);
nor U14762 (N_14762,N_5607,N_9353);
or U14763 (N_14763,N_5165,N_6662);
nand U14764 (N_14764,N_8251,N_5368);
xor U14765 (N_14765,N_6790,N_9478);
and U14766 (N_14766,N_8721,N_8362);
and U14767 (N_14767,N_6007,N_8207);
and U14768 (N_14768,N_7876,N_8237);
and U14769 (N_14769,N_6213,N_5966);
and U14770 (N_14770,N_9600,N_9665);
nand U14771 (N_14771,N_7113,N_9615);
nor U14772 (N_14772,N_9766,N_5093);
nor U14773 (N_14773,N_8555,N_5086);
or U14774 (N_14774,N_7479,N_6848);
and U14775 (N_14775,N_6299,N_9757);
and U14776 (N_14776,N_9676,N_7414);
and U14777 (N_14777,N_9775,N_7107);
nand U14778 (N_14778,N_7548,N_9866);
nor U14779 (N_14779,N_7014,N_9826);
or U14780 (N_14780,N_5167,N_9232);
nor U14781 (N_14781,N_7214,N_9216);
nand U14782 (N_14782,N_6998,N_7745);
nand U14783 (N_14783,N_6733,N_6591);
nand U14784 (N_14784,N_5568,N_9117);
or U14785 (N_14785,N_8913,N_8648);
and U14786 (N_14786,N_9850,N_7278);
or U14787 (N_14787,N_7082,N_7182);
nand U14788 (N_14788,N_9009,N_7872);
nand U14789 (N_14789,N_9118,N_6359);
nand U14790 (N_14790,N_6231,N_8474);
and U14791 (N_14791,N_5871,N_6056);
or U14792 (N_14792,N_7532,N_8793);
and U14793 (N_14793,N_5842,N_8807);
and U14794 (N_14794,N_7504,N_8507);
nand U14795 (N_14795,N_5474,N_7106);
and U14796 (N_14796,N_8754,N_9062);
nand U14797 (N_14797,N_7487,N_6268);
and U14798 (N_14798,N_9807,N_5402);
nor U14799 (N_14799,N_6835,N_9953);
or U14800 (N_14800,N_5097,N_7810);
or U14801 (N_14801,N_7422,N_6074);
nor U14802 (N_14802,N_9892,N_9876);
or U14803 (N_14803,N_9996,N_8152);
and U14804 (N_14804,N_7640,N_8811);
or U14805 (N_14805,N_9719,N_7542);
and U14806 (N_14806,N_5954,N_7122);
nor U14807 (N_14807,N_6946,N_7450);
nand U14808 (N_14808,N_8703,N_9416);
or U14809 (N_14809,N_8333,N_9101);
and U14810 (N_14810,N_6201,N_7125);
and U14811 (N_14811,N_8775,N_6059);
or U14812 (N_14812,N_5733,N_6036);
and U14813 (N_14813,N_8410,N_8939);
nand U14814 (N_14814,N_6741,N_5540);
nand U14815 (N_14815,N_5689,N_8761);
nand U14816 (N_14816,N_5540,N_6423);
nand U14817 (N_14817,N_5973,N_7717);
xor U14818 (N_14818,N_5159,N_6863);
or U14819 (N_14819,N_7050,N_9788);
and U14820 (N_14820,N_8728,N_9083);
nand U14821 (N_14821,N_9232,N_8286);
nand U14822 (N_14822,N_9439,N_9569);
nor U14823 (N_14823,N_9437,N_9531);
xor U14824 (N_14824,N_8992,N_6065);
nor U14825 (N_14825,N_8517,N_6439);
or U14826 (N_14826,N_8889,N_6094);
or U14827 (N_14827,N_8741,N_9996);
and U14828 (N_14828,N_5005,N_7024);
or U14829 (N_14829,N_8045,N_5519);
or U14830 (N_14830,N_9661,N_7436);
nor U14831 (N_14831,N_8102,N_5487);
or U14832 (N_14832,N_7256,N_6286);
nand U14833 (N_14833,N_6884,N_5371);
nor U14834 (N_14834,N_8851,N_5421);
nor U14835 (N_14835,N_8272,N_8959);
or U14836 (N_14836,N_7812,N_5915);
nand U14837 (N_14837,N_7146,N_8686);
and U14838 (N_14838,N_5620,N_9524);
or U14839 (N_14839,N_7083,N_8015);
and U14840 (N_14840,N_6886,N_8185);
and U14841 (N_14841,N_8057,N_7936);
or U14842 (N_14842,N_7730,N_5851);
or U14843 (N_14843,N_8107,N_8302);
nand U14844 (N_14844,N_7034,N_5916);
and U14845 (N_14845,N_8278,N_6802);
nor U14846 (N_14846,N_6518,N_6425);
xnor U14847 (N_14847,N_5842,N_7843);
or U14848 (N_14848,N_8039,N_6704);
or U14849 (N_14849,N_7563,N_6207);
nor U14850 (N_14850,N_5763,N_7236);
nand U14851 (N_14851,N_9474,N_9780);
nor U14852 (N_14852,N_9885,N_7496);
and U14853 (N_14853,N_7895,N_5887);
or U14854 (N_14854,N_6106,N_8239);
and U14855 (N_14855,N_7643,N_7163);
nand U14856 (N_14856,N_8953,N_7271);
nand U14857 (N_14857,N_7230,N_9131);
xor U14858 (N_14858,N_9249,N_9904);
nand U14859 (N_14859,N_9276,N_7557);
or U14860 (N_14860,N_5032,N_8717);
nand U14861 (N_14861,N_8967,N_6464);
or U14862 (N_14862,N_6031,N_9467);
or U14863 (N_14863,N_5451,N_9753);
and U14864 (N_14864,N_9694,N_9113);
and U14865 (N_14865,N_9886,N_9928);
or U14866 (N_14866,N_8517,N_8748);
nand U14867 (N_14867,N_7019,N_5681);
nand U14868 (N_14868,N_8977,N_6810);
and U14869 (N_14869,N_6937,N_7207);
or U14870 (N_14870,N_6020,N_9009);
and U14871 (N_14871,N_7981,N_8105);
or U14872 (N_14872,N_7491,N_7773);
or U14873 (N_14873,N_5836,N_8751);
and U14874 (N_14874,N_8649,N_7157);
nand U14875 (N_14875,N_7567,N_5115);
or U14876 (N_14876,N_6977,N_9406);
nor U14877 (N_14877,N_9120,N_8543);
or U14878 (N_14878,N_7347,N_7703);
or U14879 (N_14879,N_7604,N_9145);
nor U14880 (N_14880,N_8702,N_6740);
nor U14881 (N_14881,N_8774,N_8854);
or U14882 (N_14882,N_7882,N_7334);
and U14883 (N_14883,N_5058,N_7129);
xnor U14884 (N_14884,N_7806,N_9391);
nand U14885 (N_14885,N_9249,N_5374);
nand U14886 (N_14886,N_7455,N_7794);
nor U14887 (N_14887,N_9970,N_7719);
nor U14888 (N_14888,N_8296,N_6051);
nor U14889 (N_14889,N_8601,N_5426);
and U14890 (N_14890,N_7585,N_5271);
and U14891 (N_14891,N_7972,N_5650);
or U14892 (N_14892,N_8879,N_9162);
nor U14893 (N_14893,N_8182,N_6114);
nand U14894 (N_14894,N_9415,N_6681);
and U14895 (N_14895,N_8079,N_9985);
and U14896 (N_14896,N_6798,N_5666);
or U14897 (N_14897,N_6397,N_8800);
and U14898 (N_14898,N_5198,N_8290);
nand U14899 (N_14899,N_7432,N_7027);
nand U14900 (N_14900,N_8263,N_6867);
nand U14901 (N_14901,N_9065,N_8189);
or U14902 (N_14902,N_5601,N_7698);
nor U14903 (N_14903,N_8649,N_9761);
nor U14904 (N_14904,N_5143,N_6805);
and U14905 (N_14905,N_5606,N_5902);
or U14906 (N_14906,N_7200,N_8227);
or U14907 (N_14907,N_6905,N_7420);
and U14908 (N_14908,N_8394,N_7414);
nand U14909 (N_14909,N_8307,N_9816);
or U14910 (N_14910,N_8056,N_5352);
nand U14911 (N_14911,N_5761,N_8643);
and U14912 (N_14912,N_9583,N_6925);
and U14913 (N_14913,N_6193,N_6743);
or U14914 (N_14914,N_6387,N_5410);
nand U14915 (N_14915,N_6559,N_9408);
or U14916 (N_14916,N_5197,N_9678);
and U14917 (N_14917,N_6232,N_9529);
nand U14918 (N_14918,N_7194,N_9258);
and U14919 (N_14919,N_8611,N_9109);
nand U14920 (N_14920,N_9684,N_5663);
nor U14921 (N_14921,N_8908,N_6799);
or U14922 (N_14922,N_8484,N_8109);
nand U14923 (N_14923,N_9953,N_7864);
nand U14924 (N_14924,N_8142,N_7256);
and U14925 (N_14925,N_7260,N_6268);
xnor U14926 (N_14926,N_7340,N_8442);
nor U14927 (N_14927,N_6213,N_9188);
and U14928 (N_14928,N_8518,N_9800);
and U14929 (N_14929,N_8952,N_5132);
and U14930 (N_14930,N_6909,N_8659);
nor U14931 (N_14931,N_5579,N_7469);
nor U14932 (N_14932,N_5467,N_7497);
or U14933 (N_14933,N_8694,N_9798);
and U14934 (N_14934,N_6663,N_6556);
xnor U14935 (N_14935,N_6961,N_8800);
xor U14936 (N_14936,N_8707,N_8626);
or U14937 (N_14937,N_7943,N_8523);
or U14938 (N_14938,N_5463,N_5248);
nor U14939 (N_14939,N_6272,N_7544);
or U14940 (N_14940,N_8660,N_5516);
nand U14941 (N_14941,N_8291,N_8210);
and U14942 (N_14942,N_7454,N_5109);
and U14943 (N_14943,N_7811,N_5147);
nor U14944 (N_14944,N_7758,N_5247);
nor U14945 (N_14945,N_8900,N_7708);
or U14946 (N_14946,N_8902,N_7322);
nor U14947 (N_14947,N_8981,N_6188);
nor U14948 (N_14948,N_6998,N_8862);
nand U14949 (N_14949,N_6628,N_5271);
or U14950 (N_14950,N_6798,N_7048);
nand U14951 (N_14951,N_6751,N_6065);
nand U14952 (N_14952,N_9471,N_6072);
and U14953 (N_14953,N_9248,N_7285);
and U14954 (N_14954,N_5455,N_6199);
nor U14955 (N_14955,N_9418,N_5243);
nor U14956 (N_14956,N_8416,N_7305);
nand U14957 (N_14957,N_5089,N_6827);
nand U14958 (N_14958,N_8583,N_9468);
xor U14959 (N_14959,N_6411,N_9014);
nand U14960 (N_14960,N_5386,N_8304);
and U14961 (N_14961,N_9605,N_5967);
and U14962 (N_14962,N_6988,N_5255);
or U14963 (N_14963,N_8154,N_9780);
or U14964 (N_14964,N_6531,N_9891);
and U14965 (N_14965,N_7790,N_6972);
nor U14966 (N_14966,N_9080,N_6414);
and U14967 (N_14967,N_5768,N_6279);
nor U14968 (N_14968,N_6342,N_8483);
and U14969 (N_14969,N_5560,N_7932);
nand U14970 (N_14970,N_9441,N_6409);
nor U14971 (N_14971,N_9245,N_5823);
or U14972 (N_14972,N_6441,N_9814);
nand U14973 (N_14973,N_6530,N_6840);
xor U14974 (N_14974,N_7016,N_7785);
nand U14975 (N_14975,N_5601,N_9123);
nand U14976 (N_14976,N_6823,N_8729);
nand U14977 (N_14977,N_9735,N_9439);
nor U14978 (N_14978,N_9683,N_5680);
nor U14979 (N_14979,N_7644,N_6632);
and U14980 (N_14980,N_6646,N_7437);
nor U14981 (N_14981,N_5445,N_8042);
nand U14982 (N_14982,N_6140,N_6372);
and U14983 (N_14983,N_8519,N_7094);
nor U14984 (N_14984,N_6900,N_8681);
nor U14985 (N_14985,N_9070,N_5554);
or U14986 (N_14986,N_8103,N_9557);
nand U14987 (N_14987,N_9079,N_6495);
and U14988 (N_14988,N_8177,N_7514);
nand U14989 (N_14989,N_5783,N_8927);
nand U14990 (N_14990,N_5649,N_5827);
nor U14991 (N_14991,N_5784,N_7564);
or U14992 (N_14992,N_5624,N_8282);
and U14993 (N_14993,N_7368,N_7105);
nor U14994 (N_14994,N_6382,N_7570);
xnor U14995 (N_14995,N_9249,N_9049);
and U14996 (N_14996,N_6439,N_8459);
nand U14997 (N_14997,N_8697,N_9295);
and U14998 (N_14998,N_7208,N_8870);
nand U14999 (N_14999,N_5572,N_5209);
or U15000 (N_15000,N_12988,N_12130);
or U15001 (N_15001,N_12136,N_11176);
or U15002 (N_15002,N_11570,N_11479);
or U15003 (N_15003,N_11161,N_10686);
nand U15004 (N_15004,N_10380,N_11924);
and U15005 (N_15005,N_11228,N_13092);
nor U15006 (N_15006,N_12164,N_14957);
nand U15007 (N_15007,N_12784,N_14204);
nand U15008 (N_15008,N_11555,N_13679);
and U15009 (N_15009,N_14930,N_14787);
or U15010 (N_15010,N_12601,N_12915);
and U15011 (N_15011,N_12529,N_13081);
or U15012 (N_15012,N_12165,N_13082);
or U15013 (N_15013,N_13364,N_12934);
nor U15014 (N_15014,N_13657,N_14050);
and U15015 (N_15015,N_10951,N_14728);
or U15016 (N_15016,N_10364,N_11982);
and U15017 (N_15017,N_10041,N_11584);
nand U15018 (N_15018,N_12557,N_11026);
nor U15019 (N_15019,N_10851,N_14171);
nand U15020 (N_15020,N_14262,N_14547);
or U15021 (N_15021,N_11624,N_13483);
nand U15022 (N_15022,N_11623,N_14376);
and U15023 (N_15023,N_13410,N_10723);
nor U15024 (N_15024,N_11753,N_14384);
nor U15025 (N_15025,N_11090,N_13603);
nor U15026 (N_15026,N_14501,N_12450);
nor U15027 (N_15027,N_12480,N_13519);
and U15028 (N_15028,N_12242,N_11859);
nor U15029 (N_15029,N_11900,N_14567);
nand U15030 (N_15030,N_11170,N_13643);
nor U15031 (N_15031,N_14807,N_12019);
xor U15032 (N_15032,N_10334,N_10458);
and U15033 (N_15033,N_14583,N_13760);
or U15034 (N_15034,N_10983,N_12459);
and U15035 (N_15035,N_11270,N_10931);
nand U15036 (N_15036,N_11967,N_13016);
and U15037 (N_15037,N_10797,N_10978);
and U15038 (N_15038,N_14472,N_14990);
or U15039 (N_15039,N_13763,N_10308);
nor U15040 (N_15040,N_12455,N_11416);
and U15041 (N_15041,N_12024,N_13066);
and U15042 (N_15042,N_12674,N_13301);
or U15043 (N_15043,N_13709,N_14553);
nand U15044 (N_15044,N_12289,N_13246);
nor U15045 (N_15045,N_11512,N_14722);
nand U15046 (N_15046,N_11961,N_14349);
nor U15047 (N_15047,N_12399,N_11349);
or U15048 (N_15048,N_11181,N_10874);
or U15049 (N_15049,N_10321,N_10732);
nor U15050 (N_15050,N_12120,N_11152);
or U15051 (N_15051,N_14708,N_11607);
nor U15052 (N_15052,N_10633,N_13018);
and U15053 (N_15053,N_13486,N_13521);
or U15054 (N_15054,N_13038,N_12116);
nand U15055 (N_15055,N_11767,N_14261);
nand U15056 (N_15056,N_12448,N_13287);
and U15057 (N_15057,N_10876,N_11332);
and U15058 (N_15058,N_11507,N_12936);
nand U15059 (N_15059,N_12102,N_11188);
nor U15060 (N_15060,N_10117,N_14254);
or U15061 (N_15061,N_13089,N_14400);
and U15062 (N_15062,N_12226,N_14643);
nor U15063 (N_15063,N_10815,N_14983);
and U15064 (N_15064,N_14266,N_14962);
and U15065 (N_15065,N_10489,N_11149);
and U15066 (N_15066,N_11733,N_11817);
and U15067 (N_15067,N_14714,N_12265);
or U15068 (N_15068,N_13440,N_12214);
nor U15069 (N_15069,N_10840,N_12634);
nor U15070 (N_15070,N_10924,N_14710);
nor U15071 (N_15071,N_14445,N_14842);
and U15072 (N_15072,N_13153,N_12210);
nand U15073 (N_15073,N_14693,N_11340);
nor U15074 (N_15074,N_13737,N_12978);
nor U15075 (N_15075,N_12177,N_13094);
xor U15076 (N_15076,N_13717,N_11645);
or U15077 (N_15077,N_10599,N_11930);
nand U15078 (N_15078,N_11547,N_14464);
and U15079 (N_15079,N_11669,N_12990);
nand U15080 (N_15080,N_14759,N_14169);
nand U15081 (N_15081,N_13886,N_11429);
nand U15082 (N_15082,N_13481,N_10123);
and U15083 (N_15083,N_13857,N_13314);
nor U15084 (N_15084,N_10943,N_14903);
nor U15085 (N_15085,N_13101,N_10521);
nor U15086 (N_15086,N_13007,N_14928);
or U15087 (N_15087,N_10853,N_12447);
nand U15088 (N_15088,N_12572,N_14964);
or U15089 (N_15089,N_13658,N_13569);
and U15090 (N_15090,N_14539,N_11887);
or U15091 (N_15091,N_10381,N_14534);
or U15092 (N_15092,N_10543,N_10539);
or U15093 (N_15093,N_14176,N_12162);
and U15094 (N_15094,N_13666,N_14963);
nand U15095 (N_15095,N_13147,N_14460);
and U15096 (N_15096,N_13098,N_13839);
or U15097 (N_15097,N_13537,N_11463);
and U15098 (N_15098,N_14719,N_13680);
and U15099 (N_15099,N_11946,N_14636);
nor U15100 (N_15100,N_10766,N_13361);
and U15101 (N_15101,N_13581,N_14403);
and U15102 (N_15102,N_10469,N_14498);
nor U15103 (N_15103,N_12051,N_10059);
nor U15104 (N_15104,N_12734,N_12292);
nand U15105 (N_15105,N_11764,N_12350);
nor U15106 (N_15106,N_14530,N_12310);
nand U15107 (N_15107,N_10770,N_11067);
nor U15108 (N_15108,N_12538,N_11926);
and U15109 (N_15109,N_13404,N_12673);
nand U15110 (N_15110,N_14301,N_10249);
nand U15111 (N_15111,N_12706,N_10150);
or U15112 (N_15112,N_13422,N_14196);
and U15113 (N_15113,N_12542,N_13086);
nand U15114 (N_15114,N_14598,N_12754);
nand U15115 (N_15115,N_13131,N_11768);
nor U15116 (N_15116,N_10920,N_12908);
nor U15117 (N_15117,N_11711,N_11799);
or U15118 (N_15118,N_13302,N_14214);
xor U15119 (N_15119,N_10420,N_11263);
nor U15120 (N_15120,N_11418,N_14802);
or U15121 (N_15121,N_13023,N_11373);
nand U15122 (N_15122,N_14791,N_13326);
nor U15123 (N_15123,N_11486,N_12460);
or U15124 (N_15124,N_13753,N_11245);
nor U15125 (N_15125,N_10628,N_13973);
or U15126 (N_15126,N_13570,N_13381);
and U15127 (N_15127,N_11619,N_14136);
nand U15128 (N_15128,N_14825,N_13375);
nand U15129 (N_15129,N_10022,N_11941);
or U15130 (N_15130,N_13877,N_13645);
or U15131 (N_15131,N_10985,N_10804);
nand U15132 (N_15132,N_10970,N_14274);
nand U15133 (N_15133,N_10215,N_11268);
and U15134 (N_15134,N_13941,N_11474);
nand U15135 (N_15135,N_11943,N_12444);
nor U15136 (N_15136,N_10177,N_12345);
or U15137 (N_15137,N_13677,N_12597);
nand U15138 (N_15138,N_12021,N_10698);
nand U15139 (N_15139,N_12425,N_10522);
and U15140 (N_15140,N_11988,N_14372);
nor U15141 (N_15141,N_13727,N_10889);
and U15142 (N_15142,N_12294,N_13029);
and U15143 (N_15143,N_13074,N_14783);
xnor U15144 (N_15144,N_11398,N_14425);
nand U15145 (N_15145,N_13170,N_10456);
and U15146 (N_15146,N_14485,N_14006);
nor U15147 (N_15147,N_11459,N_10739);
or U15148 (N_15148,N_12325,N_14645);
nand U15149 (N_15149,N_12593,N_13851);
nor U15150 (N_15150,N_11363,N_11759);
xnor U15151 (N_15151,N_14788,N_12912);
nor U15152 (N_15152,N_10332,N_12385);
and U15153 (N_15153,N_12388,N_12604);
nand U15154 (N_15154,N_12243,N_12414);
and U15155 (N_15155,N_11047,N_11351);
or U15156 (N_15156,N_12745,N_13320);
and U15157 (N_15157,N_13437,N_10173);
nand U15158 (N_15158,N_14423,N_14115);
nor U15159 (N_15159,N_12917,N_10927);
nand U15160 (N_15160,N_14995,N_13718);
nand U15161 (N_15161,N_14480,N_13485);
or U15162 (N_15162,N_10894,N_12741);
nor U15163 (N_15163,N_13267,N_10486);
and U15164 (N_15164,N_13892,N_14684);
nand U15165 (N_15165,N_14489,N_14168);
or U15166 (N_15166,N_13154,N_10708);
or U15167 (N_15167,N_14926,N_14607);
nand U15168 (N_15168,N_10957,N_12326);
nor U15169 (N_15169,N_12690,N_13393);
nor U15170 (N_15170,N_14182,N_13487);
nor U15171 (N_15171,N_14904,N_14822);
nor U15172 (N_15172,N_10850,N_12771);
or U15173 (N_15173,N_14831,N_11060);
nor U15174 (N_15174,N_13704,N_10447);
nor U15175 (N_15175,N_11775,N_10141);
nand U15176 (N_15176,N_12454,N_14951);
nor U15177 (N_15177,N_13283,N_10484);
or U15178 (N_15178,N_13130,N_10276);
or U15179 (N_15179,N_10306,N_13420);
nand U15180 (N_15180,N_14860,N_11498);
nor U15181 (N_15181,N_10278,N_12622);
or U15182 (N_15182,N_14281,N_12232);
and U15183 (N_15183,N_12575,N_12500);
and U15184 (N_15184,N_13464,N_14560);
and U15185 (N_15185,N_11736,N_11940);
nor U15186 (N_15186,N_10438,N_12466);
xnor U15187 (N_15187,N_10568,N_14040);
xnor U15188 (N_15188,N_12303,N_14263);
or U15189 (N_15189,N_10771,N_10846);
and U15190 (N_15190,N_13212,N_11236);
and U15191 (N_15191,N_12481,N_14979);
nand U15192 (N_15192,N_10535,N_14541);
nor U15193 (N_15193,N_14624,N_12023);
nor U15194 (N_15194,N_13183,N_10558);
nand U15195 (N_15195,N_14733,N_14531);
nor U15196 (N_15196,N_13144,N_11034);
nor U15197 (N_15197,N_12327,N_14189);
nand U15198 (N_15198,N_11018,N_11960);
or U15199 (N_15199,N_14019,N_10922);
nor U15200 (N_15200,N_13938,N_13838);
and U15201 (N_15201,N_12660,N_12677);
nor U15202 (N_15202,N_14269,N_11849);
nand U15203 (N_15203,N_14556,N_11451);
and U15204 (N_15204,N_11954,N_13906);
or U15205 (N_15205,N_14276,N_12967);
nor U15206 (N_15206,N_10974,N_11288);
and U15207 (N_15207,N_14740,N_12037);
nor U15208 (N_15208,N_11316,N_12560);
nor U15209 (N_15209,N_14697,N_11395);
and U15210 (N_15210,N_14440,N_11882);
and U15211 (N_15211,N_14559,N_10800);
nand U15212 (N_15212,N_12011,N_13011);
and U15213 (N_15213,N_14187,N_11271);
nor U15214 (N_15214,N_11573,N_12358);
and U15215 (N_15215,N_12184,N_13005);
and U15216 (N_15216,N_13649,N_12403);
and U15217 (N_15217,N_13122,N_10742);
and U15218 (N_15218,N_14819,N_12919);
nand U15219 (N_15219,N_14601,N_12061);
nor U15220 (N_15220,N_11991,N_13057);
xor U15221 (N_15221,N_12486,N_10430);
and U15222 (N_15222,N_10361,N_13749);
nor U15223 (N_15223,N_13256,N_12647);
xor U15224 (N_15224,N_14426,N_13235);
and U15225 (N_15225,N_12651,N_12067);
nor U15226 (N_15226,N_13574,N_11706);
or U15227 (N_15227,N_10667,N_11850);
and U15228 (N_15228,N_13711,N_13405);
nor U15229 (N_15229,N_10477,N_10195);
nand U15230 (N_15230,N_13493,N_10485);
or U15231 (N_15231,N_10822,N_14153);
nor U15232 (N_15232,N_14396,N_10120);
or U15233 (N_15233,N_14148,N_11886);
nor U15234 (N_15234,N_14478,N_13530);
or U15235 (N_15235,N_10847,N_10488);
nor U15236 (N_15236,N_12257,N_14665);
and U15237 (N_15237,N_13242,N_10080);
or U15238 (N_15238,N_11990,N_11357);
and U15239 (N_15239,N_12779,N_11464);
or U15240 (N_15240,N_12318,N_14882);
or U15241 (N_15241,N_14449,N_14474);
nor U15242 (N_15242,N_10862,N_10424);
or U15243 (N_15243,N_12657,N_10998);
or U15244 (N_15244,N_12155,N_12810);
nand U15245 (N_15245,N_13697,N_14074);
and U15246 (N_15246,N_13380,N_11617);
and U15247 (N_15247,N_10119,N_11794);
xnor U15248 (N_15248,N_11339,N_13543);
and U15249 (N_15249,N_14484,N_12187);
or U15250 (N_15250,N_10689,N_12987);
nor U15251 (N_15251,N_14641,N_14760);
nand U15252 (N_15252,N_11232,N_13403);
and U15253 (N_15253,N_10452,N_11248);
and U15254 (N_15254,N_11216,N_11553);
nor U15255 (N_15255,N_14692,N_13049);
and U15256 (N_15256,N_12957,N_12473);
nand U15257 (N_15257,N_14758,N_13146);
or U15258 (N_15258,N_14273,N_10873);
nand U15259 (N_15259,N_13359,N_11899);
nor U15260 (N_15260,N_10218,N_10079);
and U15261 (N_15261,N_11262,N_11661);
nor U15262 (N_15262,N_10885,N_12293);
nor U15263 (N_15263,N_11806,N_13949);
or U15264 (N_15264,N_14139,N_12109);
or U15265 (N_15265,N_12646,N_13899);
or U15266 (N_15266,N_11590,N_12984);
nand U15267 (N_15267,N_12701,N_11894);
or U15268 (N_15268,N_14361,N_10167);
nand U15269 (N_15269,N_12629,N_10736);
nor U15270 (N_15270,N_12112,N_14119);
nand U15271 (N_15271,N_12360,N_10707);
nor U15272 (N_15272,N_12281,N_12369);
nand U15273 (N_15273,N_13477,N_14235);
and U15274 (N_15274,N_14065,N_12233);
or U15275 (N_15275,N_14395,N_12983);
nor U15276 (N_15276,N_11554,N_11680);
nor U15277 (N_15277,N_12737,N_11196);
nor U15278 (N_15278,N_12513,N_12705);
nor U15279 (N_15279,N_13424,N_12742);
or U15280 (N_15280,N_13732,N_10210);
nand U15281 (N_15281,N_13127,N_12456);
nand U15282 (N_15282,N_14496,N_13766);
or U15283 (N_15283,N_12556,N_11610);
nor U15284 (N_15284,N_11050,N_13823);
or U15285 (N_15285,N_12463,N_13844);
or U15286 (N_15286,N_12707,N_13588);
nor U15287 (N_15287,N_10097,N_14689);
nor U15288 (N_15288,N_11714,N_13332);
xnor U15289 (N_15289,N_11905,N_11042);
nor U15290 (N_15290,N_14775,N_11449);
and U15291 (N_15291,N_12838,N_11293);
and U15292 (N_15292,N_13745,N_13079);
nor U15293 (N_15293,N_11524,N_10919);
or U15294 (N_15294,N_11436,N_13455);
or U15295 (N_15295,N_10147,N_11186);
and U15296 (N_15296,N_13779,N_14035);
nand U15297 (N_15297,N_13444,N_14488);
and U15298 (N_15298,N_14118,N_11561);
nand U15299 (N_15299,N_12499,N_13670);
nor U15300 (N_15300,N_13612,N_14820);
nand U15301 (N_15301,N_12273,N_13847);
xnor U15302 (N_15302,N_14479,N_11783);
or U15303 (N_15303,N_10937,N_10038);
nand U15304 (N_15304,N_11121,N_11004);
nor U15305 (N_15305,N_11866,N_10396);
or U15306 (N_15306,N_11825,N_10001);
nand U15307 (N_15307,N_10179,N_14239);
nand U15308 (N_15308,N_13070,N_13635);
and U15309 (N_15309,N_11142,N_14854);
nor U15310 (N_15310,N_11198,N_10536);
nand U15311 (N_15311,N_12890,N_10949);
or U15312 (N_15312,N_12074,N_10880);
and U15313 (N_15313,N_11171,N_12491);
xnor U15314 (N_15314,N_10959,N_10004);
or U15315 (N_15315,N_14796,N_10342);
and U15316 (N_15316,N_14128,N_13004);
or U15317 (N_15317,N_10519,N_14918);
or U15318 (N_15318,N_12507,N_10542);
nor U15319 (N_15319,N_14014,N_12331);
nand U15320 (N_15320,N_13672,N_13565);
xor U15321 (N_15321,N_12946,N_13646);
or U15322 (N_15322,N_10440,N_13893);
or U15323 (N_15323,N_10273,N_14573);
xnor U15324 (N_15324,N_11548,N_11778);
nand U15325 (N_15325,N_10356,N_10216);
nor U15326 (N_15326,N_11038,N_10563);
or U15327 (N_15327,N_10325,N_13733);
or U15328 (N_15328,N_14342,N_10683);
and U15329 (N_15329,N_11519,N_10258);
and U15330 (N_15330,N_10121,N_14663);
nor U15331 (N_15331,N_13202,N_11699);
or U15332 (N_15332,N_12269,N_13830);
or U15333 (N_15333,N_10805,N_14314);
and U15334 (N_15334,N_13189,N_11546);
and U15335 (N_15335,N_10111,N_11355);
nor U15336 (N_15336,N_12221,N_12053);
or U15337 (N_15337,N_12259,N_11821);
nor U15338 (N_15338,N_12837,N_11322);
nand U15339 (N_15339,N_13193,N_13954);
xnor U15340 (N_15340,N_13648,N_13230);
and U15341 (N_15341,N_13063,N_12413);
nand U15342 (N_15342,N_13684,N_10403);
nor U15343 (N_15343,N_13213,N_10898);
and U15344 (N_15344,N_10901,N_13900);
nor U15345 (N_15345,N_12188,N_11781);
nor U15346 (N_15346,N_12899,N_10624);
nand U15347 (N_15347,N_13025,N_10500);
nor U15348 (N_15348,N_13250,N_14952);
nor U15349 (N_15349,N_12535,N_14510);
or U15350 (N_15350,N_12215,N_10413);
nand U15351 (N_15351,N_11409,N_10033);
nand U15352 (N_15352,N_10649,N_11743);
nand U15353 (N_15353,N_10789,N_13599);
or U15354 (N_15354,N_10255,N_13600);
or U15355 (N_15355,N_12445,N_13544);
or U15356 (N_15356,N_10421,N_12589);
and U15357 (N_15357,N_11311,N_14799);
or U15358 (N_15358,N_11278,N_10369);
nand U15359 (N_15359,N_11535,N_13036);
nor U15360 (N_15360,N_13308,N_11653);
nand U15361 (N_15361,N_13363,N_11480);
nor U15362 (N_15362,N_14463,N_11388);
and U15363 (N_15363,N_12260,N_10527);
nor U15364 (N_15364,N_12341,N_11013);
nor U15365 (N_15365,N_10827,N_11014);
nand U15366 (N_15366,N_11335,N_13654);
and U15367 (N_15367,N_13998,N_13972);
nor U15368 (N_15368,N_12173,N_14415);
nor U15369 (N_15369,N_12979,N_12346);
or U15370 (N_15370,N_10310,N_13429);
nor U15371 (N_15371,N_13741,N_10138);
nand U15372 (N_15372,N_14143,N_12351);
nand U15373 (N_15373,N_12235,N_13263);
nor U15374 (N_15374,N_10050,N_14847);
or U15375 (N_15375,N_11250,N_12541);
nor U15376 (N_15376,N_11620,N_11426);
and U15377 (N_15377,N_10836,N_11875);
or U15378 (N_15378,N_12678,N_10990);
or U15379 (N_15379,N_14275,N_11386);
or U15380 (N_15380,N_10618,N_13663);
xor U15381 (N_15381,N_14683,N_14348);
nor U15382 (N_15382,N_10231,N_14456);
or U15383 (N_15383,N_10843,N_11092);
nand U15384 (N_15384,N_13702,N_11745);
and U15385 (N_15385,N_11108,N_13416);
nand U15386 (N_15386,N_13328,N_12441);
xnor U15387 (N_15387,N_14878,N_13118);
and U15388 (N_15388,N_14914,N_12174);
nor U15389 (N_15389,N_12749,N_13333);
xnor U15390 (N_15390,N_12615,N_13143);
nand U15391 (N_15391,N_11998,N_13868);
nor U15392 (N_15392,N_11218,N_10900);
nand U15393 (N_15393,N_14121,N_14155);
and U15394 (N_15394,N_11174,N_14872);
and U15395 (N_15395,N_12344,N_10712);
or U15396 (N_15396,N_10912,N_14385);
and U15397 (N_15397,N_13536,N_13021);
and U15398 (N_15398,N_11410,N_14865);
nor U15399 (N_15399,N_14130,N_13223);
and U15400 (N_15400,N_14190,N_11717);
nor U15401 (N_15401,N_14768,N_11971);
nor U15402 (N_15402,N_10761,N_12623);
or U15403 (N_15403,N_14855,N_10436);
or U15404 (N_15404,N_10107,N_12090);
nand U15405 (N_15405,N_11118,N_12492);
or U15406 (N_15406,N_11842,N_10219);
or U15407 (N_15407,N_11190,N_13983);
and U15408 (N_15408,N_12758,N_14152);
nand U15409 (N_15409,N_14905,N_14521);
or U15410 (N_15410,N_13201,N_14292);
or U15411 (N_15411,N_10906,N_14499);
nor U15412 (N_15412,N_10475,N_12435);
nand U15413 (N_15413,N_11867,N_12044);
and U15414 (N_15414,N_10577,N_10463);
xnor U15415 (N_15415,N_11689,N_10935);
nand U15416 (N_15416,N_11734,N_10189);
nand U15417 (N_15417,N_12013,N_13052);
nand U15418 (N_15418,N_10832,N_10288);
nand U15419 (N_15419,N_14288,N_13699);
or U15420 (N_15420,N_13323,N_12652);
or U15421 (N_15421,N_14132,N_11615);
or U15422 (N_15422,N_13678,N_14828);
xor U15423 (N_15423,N_12016,N_10243);
or U15424 (N_15424,N_10584,N_10194);
nand U15425 (N_15425,N_14270,N_11932);
nand U15426 (N_15426,N_12603,N_11477);
and U15427 (N_15427,N_13650,N_14233);
or U15428 (N_15428,N_14563,N_12650);
nor U15429 (N_15429,N_10236,N_14402);
and U15430 (N_15430,N_13355,N_14699);
nand U15431 (N_15431,N_12725,N_14369);
nor U15432 (N_15432,N_10807,N_12471);
nand U15433 (N_15433,N_11044,N_14414);
and U15434 (N_15434,N_14451,N_14680);
nor U15435 (N_15435,N_11287,N_14388);
and U15436 (N_15436,N_14251,N_14336);
or U15437 (N_15437,N_12366,N_10213);
or U15438 (N_15438,N_14518,N_10106);
or U15439 (N_15439,N_12820,N_14294);
nand U15440 (N_15440,N_12052,N_10407);
or U15441 (N_15441,N_13069,N_10966);
and U15442 (N_15442,N_14900,N_11124);
and U15443 (N_15443,N_12371,N_10432);
or U15444 (N_15444,N_11165,N_11731);
or U15445 (N_15445,N_14315,N_14216);
and U15446 (N_15446,N_11175,N_14901);
nand U15447 (N_15447,N_13571,N_10710);
nor U15448 (N_15448,N_13494,N_12409);
and U15449 (N_15449,N_11679,N_14197);
nand U15450 (N_15450,N_10327,N_12852);
nand U15451 (N_15451,N_13706,N_10863);
nor U15452 (N_15452,N_13959,N_11888);
or U15453 (N_15453,N_12167,N_13808);
nand U15454 (N_15454,N_11267,N_13347);
or U15455 (N_15455,N_13577,N_11039);
nand U15456 (N_15456,N_11273,N_12079);
xnor U15457 (N_15457,N_12993,N_10755);
and U15458 (N_15458,N_14446,N_12540);
and U15459 (N_15459,N_12910,N_10303);
nor U15460 (N_15460,N_14891,N_12189);
or U15461 (N_15461,N_12947,N_12698);
nor U15462 (N_15462,N_11879,N_10392);
or U15463 (N_15463,N_12728,N_13948);
and U15464 (N_15464,N_14897,N_12223);
and U15465 (N_15465,N_12839,N_14554);
nor U15466 (N_15466,N_12075,N_11362);
or U15467 (N_15467,N_12977,N_11591);
nor U15468 (N_15468,N_12739,N_10299);
and U15469 (N_15469,N_13400,N_10277);
nand U15470 (N_15470,N_10507,N_10042);
nand U15471 (N_15471,N_10849,N_10331);
or U15472 (N_15472,N_14748,N_13383);
nor U15473 (N_15473,N_10196,N_14871);
or U15474 (N_15474,N_12914,N_12335);
or U15475 (N_15475,N_10478,N_13124);
nor U15476 (N_15476,N_14540,N_12710);
or U15477 (N_15477,N_12099,N_14508);
and U15478 (N_15478,N_11642,N_11139);
nor U15479 (N_15479,N_13724,N_10666);
nor U15480 (N_15480,N_14730,N_10802);
and U15481 (N_15481,N_11801,N_13020);
or U15482 (N_15482,N_11687,N_10127);
nand U15483 (N_15483,N_11021,N_10939);
or U15484 (N_15484,N_14422,N_10501);
or U15485 (N_15485,N_13630,N_14784);
nor U15486 (N_15486,N_13901,N_14550);
and U15487 (N_15487,N_10767,N_13575);
nand U15488 (N_15488,N_14178,N_11102);
and U15489 (N_15489,N_10910,N_12158);
nor U15490 (N_15490,N_14146,N_11189);
or U15491 (N_15491,N_12224,N_13239);
xnor U15492 (N_15492,N_10881,N_12815);
nand U15493 (N_15493,N_14492,N_13969);
and U15494 (N_15494,N_12082,N_13865);
or U15495 (N_15495,N_14394,N_11172);
or U15496 (N_15496,N_11350,N_11752);
nor U15497 (N_15497,N_10293,N_14971);
nor U15498 (N_15498,N_13156,N_14524);
or U15499 (N_15499,N_10244,N_12747);
nor U15500 (N_15500,N_10730,N_11500);
and U15501 (N_15501,N_14815,N_11608);
or U15502 (N_15502,N_12616,N_12217);
and U15503 (N_15503,N_10359,N_14310);
nor U15504 (N_15504,N_14711,N_13908);
or U15505 (N_15505,N_10201,N_10801);
nor U15506 (N_15506,N_12530,N_10465);
nor U15507 (N_15507,N_14803,N_11770);
nand U15508 (N_15508,N_12191,N_12125);
nor U15509 (N_15509,N_10634,N_10612);
nand U15510 (N_15510,N_14543,N_14106);
nor U15511 (N_15511,N_13631,N_12537);
and U15512 (N_15512,N_11542,N_10696);
or U15513 (N_15513,N_11810,N_11713);
and U15514 (N_15514,N_10096,N_12282);
and U15515 (N_15515,N_12431,N_10690);
or U15516 (N_15516,N_11098,N_10307);
nand U15517 (N_15517,N_10635,N_12380);
xnor U15518 (N_15518,N_10172,N_13339);
and U15519 (N_15519,N_10858,N_12778);
nor U15520 (N_15520,N_11581,N_13656);
and U15521 (N_15521,N_11545,N_14406);
nand U15522 (N_15522,N_13179,N_11670);
xor U15523 (N_15523,N_14381,N_13754);
xnor U15524 (N_15524,N_14193,N_10422);
or U15525 (N_15525,N_13059,N_12968);
nor U15526 (N_15526,N_13155,N_10598);
and U15527 (N_15527,N_14066,N_12665);
nor U15528 (N_15528,N_13854,N_12826);
nand U15529 (N_15529,N_12315,N_13623);
and U15530 (N_15530,N_11730,N_14244);
nand U15531 (N_15531,N_14911,N_10343);
nor U15532 (N_15532,N_11798,N_14353);
or U15533 (N_15533,N_11719,N_10098);
nand U15534 (N_15534,N_10125,N_13826);
and U15535 (N_15535,N_12662,N_14574);
or U15536 (N_15536,N_13317,N_10126);
and U15537 (N_15537,N_11688,N_13028);
nor U15538 (N_15538,N_13190,N_10679);
and U15539 (N_15539,N_14660,N_11086);
xor U15540 (N_15540,N_10192,N_12683);
or U15541 (N_15541,N_12057,N_10928);
or U15542 (N_15542,N_11747,N_10086);
nand U15543 (N_15543,N_10018,N_12692);
nor U15544 (N_15544,N_14927,N_11259);
nand U15545 (N_15545,N_13843,N_12585);
or U15546 (N_15546,N_13047,N_14629);
nand U15547 (N_15547,N_10318,N_11742);
nor U15548 (N_15548,N_14398,N_11465);
nand U15549 (N_15549,N_12343,N_11919);
nor U15550 (N_15550,N_14659,N_12036);
or U15551 (N_15551,N_13056,N_10282);
or U15552 (N_15552,N_14329,N_12525);
and U15553 (N_15553,N_13266,N_10729);
nor U15554 (N_15554,N_13158,N_11987);
or U15555 (N_15555,N_10035,N_14051);
nand U15556 (N_15556,N_12866,N_11240);
nor U15557 (N_15557,N_11716,N_10017);
or U15558 (N_15558,N_11433,N_10166);
nand U15559 (N_15559,N_14004,N_11802);
and U15560 (N_15560,N_11159,N_11404);
nor U15561 (N_15561,N_10207,N_13024);
nor U15562 (N_15562,N_14191,N_12251);
nor U15563 (N_15563,N_14652,N_14272);
nor U15564 (N_15564,N_11343,N_10721);
nor U15565 (N_15565,N_11291,N_10918);
nand U15566 (N_15566,N_10648,N_14477);
nor U15567 (N_15567,N_10235,N_10222);
nor U15568 (N_15568,N_14365,N_12744);
nand U15569 (N_15569,N_11931,N_12605);
nand U15570 (N_15570,N_12049,N_10416);
and U15571 (N_15571,N_13090,N_14507);
or U15572 (N_15572,N_10613,N_13946);
or U15573 (N_15573,N_13304,N_12107);
and U15574 (N_15574,N_13685,N_11312);
nand U15575 (N_15575,N_10028,N_10188);
and U15576 (N_15576,N_11402,N_12509);
or U15577 (N_15577,N_10794,N_11247);
and U15578 (N_15578,N_14053,N_14793);
xnor U15579 (N_15579,N_11660,N_12906);
nor U15580 (N_15580,N_10302,N_11379);
nand U15581 (N_15581,N_14305,N_10907);
nor U15582 (N_15582,N_11446,N_10434);
nor U15583 (N_15583,N_11975,N_14942);
or U15584 (N_15584,N_13927,N_13884);
and U15585 (N_15585,N_14590,N_11333);
nor U15586 (N_15586,N_10406,N_13840);
nand U15587 (N_15587,N_11099,N_11853);
and U15588 (N_15588,N_12421,N_11414);
or U15589 (N_15589,N_11365,N_11725);
or U15590 (N_15590,N_12782,N_12353);
nand U15591 (N_15591,N_11454,N_11577);
nand U15592 (N_15592,N_14649,N_13747);
nand U15593 (N_15593,N_10586,N_12986);
nor U15594 (N_15594,N_12594,N_13365);
nor U15595 (N_15595,N_11318,N_11130);
or U15596 (N_15596,N_13776,N_12299);
or U15597 (N_15597,N_10266,N_13182);
or U15598 (N_15598,N_12314,N_13296);
nor U15599 (N_15599,N_12196,N_11337);
or U15600 (N_15600,N_13064,N_10921);
and U15601 (N_15601,N_14709,N_14095);
nor U15602 (N_15602,N_13817,N_13407);
nor U15603 (N_15603,N_10466,N_13861);
and U15604 (N_15604,N_11983,N_12545);
or U15605 (N_15605,N_14713,N_10677);
or U15606 (N_15606,N_10694,N_13761);
nand U15607 (N_15607,N_14880,N_14206);
nor U15608 (N_15608,N_14974,N_10362);
and U15609 (N_15609,N_13115,N_11692);
nor U15610 (N_15610,N_13905,N_12270);
and U15611 (N_15611,N_11915,N_10205);
nand U15612 (N_15612,N_10220,N_10350);
nand U15613 (N_15613,N_13338,N_10021);
and U15614 (N_15614,N_13520,N_12971);
and U15615 (N_15615,N_14797,N_11569);
nand U15616 (N_15616,N_12997,N_10451);
nor U15617 (N_15617,N_12138,N_14925);
and U15618 (N_15618,N_14774,N_13376);
or U15619 (N_15619,N_14743,N_10152);
nand U15620 (N_15620,N_13428,N_10626);
and U15621 (N_15621,N_11836,N_13538);
nor U15622 (N_15622,N_11830,N_10768);
and U15623 (N_15623,N_14242,N_12790);
or U15624 (N_15624,N_10831,N_11834);
nand U15625 (N_15625,N_13693,N_14161);
nor U15626 (N_15626,N_11544,N_12482);
nor U15627 (N_15627,N_13999,N_12534);
or U15628 (N_15628,N_12803,N_10868);
nor U15629 (N_15629,N_13500,N_14399);
nor U15630 (N_15630,N_10214,N_13034);
nor U15631 (N_15631,N_14149,N_11659);
or U15632 (N_15632,N_11643,N_11153);
or U15633 (N_15633,N_11421,N_10941);
nor U15634 (N_15634,N_10629,N_11358);
or U15635 (N_15635,N_12774,N_13634);
nand U15636 (N_15636,N_10368,N_13356);
nand U15637 (N_15637,N_12667,N_10678);
and U15638 (N_15638,N_10074,N_14776);
and U15639 (N_15639,N_13984,N_10339);
or U15640 (N_15640,N_11822,N_11051);
or U15641 (N_15641,N_10980,N_10153);
or U15642 (N_15642,N_11633,N_12904);
and U15643 (N_15643,N_12252,N_14245);
nand U15644 (N_15644,N_11091,N_10161);
nor U15645 (N_15645,N_14890,N_14209);
and U15646 (N_15646,N_10744,N_11212);
or U15647 (N_15647,N_10981,N_10743);
xor U15648 (N_15648,N_11036,N_11505);
nand U15649 (N_15649,N_12641,N_14331);
nand U15650 (N_15650,N_10433,N_12408);
nand U15651 (N_15651,N_13318,N_10468);
nor U15652 (N_15652,N_10757,N_14284);
or U15653 (N_15653,N_13744,N_13837);
and U15654 (N_15654,N_13396,N_13807);
nand U15655 (N_15655,N_14098,N_13293);
or U15656 (N_15656,N_12970,N_10056);
nor U15657 (N_15657,N_14085,N_10140);
nand U15658 (N_15658,N_10204,N_10116);
or U15659 (N_15659,N_10639,N_10036);
nand U15660 (N_15660,N_13436,N_10971);
nand U15661 (N_15661,N_10006,N_12332);
and U15662 (N_15662,N_10292,N_14354);
nand U15663 (N_15663,N_10280,N_10829);
nor U15664 (N_15664,N_10144,N_12916);
nor U15665 (N_15665,N_14208,N_14142);
nand U15666 (N_15666,N_10168,N_14741);
or U15667 (N_15667,N_10841,N_11496);
or U15668 (N_15668,N_13087,N_14236);
nand U15669 (N_15669,N_14955,N_13695);
nor U15670 (N_15670,N_13819,N_10608);
nor U15671 (N_15671,N_12980,N_12928);
and U15672 (N_15672,N_11201,N_12100);
nor U15673 (N_15673,N_11101,N_12848);
or U15674 (N_15674,N_10367,N_12755);
nand U15675 (N_15675,N_10473,N_14046);
or U15676 (N_15676,N_11113,N_12080);
nor U15677 (N_15677,N_10217,N_13435);
nor U15678 (N_15678,N_10923,N_14669);
nor U15679 (N_15679,N_13665,N_14008);
nand U15680 (N_15680,N_11443,N_12822);
or U15681 (N_15681,N_10093,N_14028);
nor U15682 (N_15682,N_12874,N_10316);
nand U15683 (N_15683,N_11020,N_10848);
nand U15684 (N_15684,N_12546,N_11070);
nor U15685 (N_15685,N_11916,N_14993);
nor U15686 (N_15686,N_14677,N_14742);
nand U15687 (N_15687,N_14075,N_13379);
nor U15688 (N_15688,N_12329,N_13495);
nand U15689 (N_15689,N_12945,N_13965);
and U15690 (N_15690,N_14453,N_13238);
nand U15691 (N_15691,N_12935,N_13616);
nor U15692 (N_15692,N_11305,N_10039);
nand U15693 (N_15693,N_13810,N_13390);
xor U15694 (N_15694,N_10809,N_13871);
and U15695 (N_15695,N_13981,N_13466);
or U15696 (N_15696,N_12205,N_14009);
or U15697 (N_15697,N_11721,N_14250);
nand U15698 (N_15698,N_14468,N_10702);
nand U15699 (N_15699,N_10557,N_12769);
and U15700 (N_15700,N_13557,N_10043);
nor U15701 (N_15701,N_13205,N_11489);
nand U15702 (N_15702,N_12203,N_11635);
or U15703 (N_15703,N_13408,N_12618);
and U15704 (N_15704,N_14528,N_10287);
and U15705 (N_15705,N_12571,N_13518);
nand U15706 (N_15706,N_11727,N_10333);
nor U15707 (N_15707,N_10225,N_12239);
nor U15708 (N_15708,N_12859,N_11986);
nand U15709 (N_15709,N_14616,N_11984);
or U15710 (N_15710,N_11756,N_10899);
nand U15711 (N_15711,N_14447,N_13104);
nand U15712 (N_15712,N_12875,N_13698);
or U15713 (N_15713,N_12470,N_10516);
nand U15714 (N_15714,N_13457,N_14938);
or U15715 (N_15715,N_10005,N_13019);
and U15716 (N_15716,N_13012,N_10773);
or U15717 (N_15717,N_10082,N_14282);
nand U15718 (N_15718,N_11666,N_12956);
nor U15719 (N_15719,N_13818,N_12362);
or U15720 (N_15720,N_12268,N_11878);
or U15721 (N_15721,N_12168,N_12569);
nand U15722 (N_15722,N_11327,N_10174);
nor U15723 (N_15723,N_10186,N_11056);
and U15724 (N_15724,N_12216,N_13200);
or U15725 (N_15725,N_12145,N_11678);
or U15726 (N_15726,N_14055,N_14718);
nand U15727 (N_15727,N_12564,N_14473);
nor U15728 (N_15728,N_10015,N_11179);
nor U15729 (N_15729,N_14493,N_11406);
or U15730 (N_15730,N_11621,N_14587);
and U15731 (N_15731,N_10571,N_14727);
and U15732 (N_15732,N_14868,N_14077);
or U15733 (N_15733,N_10499,N_13736);
nand U15734 (N_15734,N_13515,N_10662);
nand U15735 (N_15735,N_13608,N_14920);
nand U15736 (N_15736,N_12248,N_13102);
or U15737 (N_15737,N_14939,N_12580);
nor U15738 (N_15738,N_14696,N_12279);
and U15739 (N_15739,N_12410,N_11787);
and U15740 (N_15740,N_10137,N_14124);
and U15741 (N_15741,N_12877,N_11583);
nor U15742 (N_15742,N_14902,N_11600);
or U15743 (N_15743,N_12206,N_13510);
nor U15744 (N_15744,N_10950,N_14611);
nand U15745 (N_15745,N_10428,N_13765);
nor U15746 (N_15746,N_14243,N_10779);
nor U15747 (N_15747,N_12584,N_12730);
nor U15748 (N_15748,N_10909,N_14744);
nor U15749 (N_15749,N_13957,N_14258);
nor U15750 (N_15750,N_11618,N_11482);
nor U15751 (N_15751,N_10719,N_11215);
and U15752 (N_15752,N_11007,N_11059);
and U15753 (N_15753,N_11658,N_10304);
or U15754 (N_15754,N_12813,N_12696);
nand U15755 (N_15755,N_14538,N_12098);
or U15756 (N_15756,N_14227,N_12583);
and U15757 (N_15757,N_11981,N_10897);
nand U15758 (N_15758,N_11490,N_12505);
nor U15759 (N_15759,N_12909,N_13929);
and U15760 (N_15760,N_10437,N_10425);
or U15761 (N_15761,N_10049,N_13522);
or U15762 (N_15762,N_10023,N_10241);
or U15763 (N_15763,N_13970,N_10312);
or U15764 (N_15764,N_10606,N_12108);
and U15765 (N_15765,N_13820,N_10999);
or U15766 (N_15766,N_11784,N_10833);
nor U15767 (N_15767,N_11413,N_12798);
nand U15768 (N_15768,N_12528,N_10600);
nor U15769 (N_15769,N_14110,N_10699);
nor U15770 (N_15770,N_11995,N_10940);
and U15771 (N_15771,N_12719,N_13735);
nor U15772 (N_15772,N_14482,N_11359);
nor U15773 (N_15773,N_13324,N_13506);
nor U15774 (N_15774,N_13958,N_11061);
nor U15775 (N_15775,N_10798,N_13805);
nor U15776 (N_15776,N_13027,N_12373);
xnor U15777 (N_15777,N_11673,N_12733);
nand U15778 (N_15778,N_14519,N_12181);
nand U15779 (N_15779,N_11602,N_10305);
nor U15780 (N_15780,N_10537,N_12923);
or U15781 (N_15781,N_10573,N_14411);
nand U15782 (N_15782,N_13335,N_10709);
or U15783 (N_15783,N_12645,N_10965);
nor U15784 (N_15784,N_11662,N_13053);
and U15785 (N_15785,N_10375,N_12402);
nand U15786 (N_15786,N_14432,N_13953);
and U15787 (N_15787,N_13438,N_14304);
nand U15788 (N_15788,N_13468,N_13345);
and U15789 (N_15789,N_12149,N_13584);
or U15790 (N_15790,N_13233,N_13633);
nand U15791 (N_15791,N_11740,N_10198);
nand U15792 (N_15792,N_14695,N_13401);
nor U15793 (N_15793,N_10553,N_13956);
and U15794 (N_15794,N_10726,N_10692);
or U15795 (N_15795,N_11475,N_14358);
and U15796 (N_15796,N_13231,N_12427);
or U15797 (N_15797,N_12762,N_11258);
or U15798 (N_15798,N_12284,N_10619);
or U15799 (N_15799,N_12802,N_11516);
or U15800 (N_15800,N_14870,N_10652);
nand U15801 (N_15801,N_12777,N_13382);
nand U15802 (N_15802,N_11985,N_13887);
nand U15803 (N_15803,N_14976,N_13831);
and U15804 (N_15804,N_10684,N_10377);
nand U15805 (N_15805,N_11163,N_10358);
nand U15806 (N_15806,N_14886,N_13642);
and U15807 (N_15807,N_11593,N_10787);
nor U15808 (N_15808,N_12590,N_13960);
and U15809 (N_15809,N_13639,N_13221);
or U15810 (N_15810,N_13395,N_12198);
or U15811 (N_15811,N_14097,N_13539);
and U15812 (N_15812,N_10092,N_12816);
nand U15813 (N_15813,N_10784,N_10704);
or U15814 (N_15814,N_12193,N_10984);
and U15815 (N_15815,N_12291,N_11272);
nand U15816 (N_15816,N_10068,N_11948);
or U15817 (N_15817,N_10884,N_11690);
or U15818 (N_15818,N_11024,N_13517);
nor U15819 (N_15819,N_10030,N_12743);
or U15820 (N_15820,N_14940,N_11114);
nand U15821 (N_15821,N_12628,N_12920);
and U15822 (N_15822,N_14751,N_14224);
or U15823 (N_15823,N_13815,N_11300);
nor U15824 (N_15824,N_11739,N_10602);
nand U15825 (N_15825,N_13249,N_10716);
nor U15826 (N_15826,N_10020,N_13045);
and U15827 (N_15827,N_14679,N_12829);
or U15828 (N_15828,N_14738,N_14612);
nand U15829 (N_15829,N_13367,N_11843);
or U15830 (N_15830,N_12220,N_13106);
or U15831 (N_15831,N_14861,N_13931);
and U15832 (N_15832,N_13352,N_12961);
nand U15833 (N_15833,N_14581,N_11045);
xnor U15834 (N_15834,N_12687,N_11686);
nor U15835 (N_15835,N_14184,N_14984);
nor U15836 (N_15836,N_10329,N_14810);
and U15837 (N_15837,N_14763,N_12748);
or U15838 (N_15838,N_11314,N_12262);
nor U15839 (N_15839,N_10655,N_11648);
nand U15840 (N_15840,N_13691,N_11950);
and U15841 (N_15841,N_12611,N_10130);
nor U15842 (N_15842,N_11969,N_10455);
nor U15843 (N_15843,N_12407,N_14851);
nor U15844 (N_15844,N_14017,N_11580);
or U15845 (N_15845,N_11700,N_11192);
or U15846 (N_15846,N_13513,N_13832);
nand U15847 (N_15847,N_12428,N_12863);
or U15848 (N_15848,N_14651,N_13525);
or U15849 (N_15849,N_13511,N_10774);
nor U15850 (N_15850,N_11494,N_14747);
nor U15851 (N_15851,N_12170,N_12422);
nor U15852 (N_15852,N_13441,N_10199);
or U15853 (N_15853,N_12805,N_10104);
or U15854 (N_15854,N_12896,N_14526);
and U15855 (N_15855,N_11632,N_11902);
or U15856 (N_15856,N_13060,N_14931);
and U15857 (N_15857,N_13195,N_14945);
xor U15858 (N_15858,N_10084,N_13874);
and U15859 (N_15859,N_11606,N_14211);
and U15860 (N_15860,N_13385,N_10374);
and U15861 (N_15861,N_11112,N_12256);
nor U15862 (N_15862,N_13586,N_12976);
and U15863 (N_15863,N_12998,N_13849);
and U15864 (N_15864,N_10552,N_12732);
or U15865 (N_15865,N_12411,N_13145);
nand U15866 (N_15866,N_12311,N_11741);
or U15867 (N_15867,N_12468,N_11910);
nand U15868 (N_15868,N_13850,N_14045);
nor U15869 (N_15869,N_13652,N_13336);
or U15870 (N_15870,N_11461,N_11906);
and U15871 (N_15871,N_13548,N_11481);
nand U15872 (N_15872,N_14427,N_10968);
and U15873 (N_15873,N_13940,N_11723);
nand U15874 (N_15874,N_14935,N_12412);
or U15875 (N_15875,N_13910,N_10311);
and U15876 (N_15876,N_13715,N_13191);
nor U15877 (N_15877,N_11261,N_12800);
nand U15878 (N_15878,N_10372,N_12553);
nand U15879 (N_15879,N_12617,N_10146);
nor U15880 (N_15880,N_11527,N_11214);
nand U15881 (N_15881,N_14832,N_14782);
nor U15882 (N_15882,N_13446,N_10270);
nand U15883 (N_15883,N_13909,N_13509);
or U15884 (N_15884,N_13095,N_13085);
nor U15885 (N_15885,N_13460,N_12612);
or U15886 (N_15886,N_10987,N_14162);
and U15887 (N_15887,N_11430,N_14549);
xor U15888 (N_15888,N_13606,N_11224);
nor U15889 (N_15889,N_13298,N_14458);
and U15890 (N_15890,N_14264,N_12999);
nor U15891 (N_15891,N_14600,N_14912);
nand U15892 (N_15892,N_10378,N_10247);
nand U15893 (N_15893,N_10100,N_11851);
nor U15894 (N_15894,N_10108,N_11876);
nor U15895 (N_15895,N_13590,N_13712);
and U15896 (N_15896,N_13458,N_13617);
nor U15897 (N_15897,N_14544,N_13700);
nand U15898 (N_15898,N_11411,N_14356);
nor U15899 (N_15899,N_13002,N_10674);
or U15900 (N_15900,N_13177,N_13554);
and U15901 (N_15901,N_11049,N_12426);
or U15902 (N_15902,N_14434,N_11484);
and U15903 (N_15903,N_13728,N_14757);
nor U15904 (N_15904,N_12451,N_12458);
and U15905 (N_15905,N_10482,N_10143);
and U15906 (N_15906,N_13876,N_11345);
and U15907 (N_15907,N_11031,N_11520);
nor U15908 (N_15908,N_14047,N_12166);
or U15909 (N_15909,N_13300,N_10349);
or U15910 (N_15910,N_13110,N_14769);
or U15911 (N_15911,N_11664,N_11353);
nand U15912 (N_15912,N_14992,N_12316);
nor U15913 (N_15913,N_10570,N_14011);
or U15914 (N_15914,N_13533,N_13255);
nor U15915 (N_15915,N_11965,N_10796);
and U15916 (N_15916,N_12078,N_12484);
and U15917 (N_15917,N_13930,N_11230);
and U15918 (N_15918,N_13987,N_10870);
or U15919 (N_15919,N_13853,N_10370);
nor U15920 (N_15920,N_11220,N_10226);
and U15921 (N_15921,N_12132,N_10803);
nor U15922 (N_15922,N_11522,N_13470);
and U15923 (N_15923,N_14150,N_11284);
and U15924 (N_15924,N_14407,N_11219);
xor U15925 (N_15925,N_12659,N_14170);
or U15926 (N_15926,N_12179,N_14630);
nor U15927 (N_15927,N_13542,N_11331);
or U15928 (N_15928,N_12213,N_12297);
nor U15929 (N_15929,N_11611,N_13535);
nor U15930 (N_15930,N_12656,N_13638);
nor U15931 (N_15931,N_11187,N_12072);
and U15932 (N_15932,N_11710,N_14091);
and U15933 (N_15933,N_11017,N_11495);
or U15934 (N_15934,N_13860,N_14707);
nand U15935 (N_15935,N_13080,N_13556);
nor U15936 (N_15936,N_13083,N_12069);
nand U15937 (N_15937,N_13508,N_10580);
and U15938 (N_15938,N_12364,N_12939);
or U15939 (N_15939,N_14205,N_13142);
nand U15940 (N_15940,N_10073,N_11627);
nor U15941 (N_15941,N_13421,N_12144);
nand U15942 (N_15942,N_10903,N_13353);
nor U15943 (N_15943,N_13568,N_11252);
nand U15944 (N_15944,N_13796,N_10286);
nand U15945 (N_15945,N_11435,N_11367);
nor U15946 (N_15946,N_13285,N_10623);
or U15947 (N_15947,N_10955,N_12415);
xor U15948 (N_15948,N_11302,N_12855);
or U15949 (N_15949,N_12485,N_12288);
and U15950 (N_15950,N_13236,N_11761);
or U15951 (N_15951,N_12868,N_13450);
nand U15952 (N_15952,N_13418,N_14134);
and U15953 (N_15953,N_10969,N_14946);
or U15954 (N_15954,N_10574,N_14805);
and U15955 (N_15955,N_11234,N_13253);
and U15956 (N_15956,N_10497,N_14202);
or U15957 (N_15957,N_13762,N_11264);
or U15958 (N_15958,N_10972,N_13835);
xnor U15959 (N_15959,N_12792,N_13614);
nand U15960 (N_15960,N_12740,N_12927);
nand U15961 (N_15961,N_13561,N_11306);
or U15962 (N_15962,N_10593,N_10389);
and U15963 (N_15963,N_14454,N_14307);
nor U15964 (N_15964,N_12510,N_10411);
and U15965 (N_15965,N_14430,N_13869);
or U15966 (N_15966,N_12119,N_13739);
or U15967 (N_15967,N_11929,N_14570);
and U15968 (N_15968,N_11466,N_13560);
nor U15969 (N_15969,N_13564,N_13541);
nor U15970 (N_15970,N_11035,N_13816);
xnor U15971 (N_15971,N_12237,N_11972);
nor U15972 (N_15972,N_13262,N_14715);
nand U15973 (N_15973,N_11456,N_13072);
nand U15974 (N_15974,N_10640,N_11579);
nor U15975 (N_15975,N_12858,N_10835);
nor U15976 (N_15976,N_10142,N_11483);
or U15977 (N_15977,N_14504,N_10942);
and U15978 (N_15978,N_14174,N_11251);
nand U15979 (N_15979,N_13578,N_12498);
nor U15980 (N_15980,N_13372,N_12359);
or U15981 (N_15981,N_11372,N_14109);
nor U15982 (N_15982,N_13748,N_11222);
and U15983 (N_15983,N_12076,N_10319);
and U15984 (N_15984,N_11082,N_10472);
or U15985 (N_15985,N_13188,N_11033);
nor U15986 (N_15986,N_11782,N_11766);
nand U15987 (N_15987,N_14048,N_12007);
xor U15988 (N_15988,N_11636,N_10933);
nor U15989 (N_15989,N_12394,N_14123);
nor U15990 (N_15990,N_14296,N_14924);
and U15991 (N_15991,N_11513,N_10886);
and U15992 (N_15992,N_13459,N_12347);
and U15993 (N_15993,N_10313,N_14404);
xor U15994 (N_15994,N_12825,N_14181);
nand U15995 (N_15995,N_12086,N_11737);
nand U15996 (N_15996,N_10638,N_14512);
or U15997 (N_15997,N_10676,N_12950);
nand U15998 (N_15998,N_11106,N_12009);
nor U15999 (N_15999,N_10842,N_13814);
nor U16000 (N_16000,N_10916,N_11568);
and U16001 (N_16001,N_12304,N_10099);
nand U16002 (N_16002,N_11510,N_12508);
or U16003 (N_16003,N_13022,N_10653);
xor U16004 (N_16004,N_14450,N_11909);
and U16005 (N_16005,N_10654,N_11675);
nand U16006 (N_16006,N_10529,N_10625);
and U16007 (N_16007,N_14079,N_10973);
and U16008 (N_16008,N_11760,N_10155);
or U16009 (N_16009,N_11707,N_13566);
nand U16010 (N_16010,N_13675,N_11777);
nor U16011 (N_16011,N_14967,N_10385);
or U16012 (N_16012,N_13821,N_10956);
xnor U16013 (N_16013,N_13427,N_13058);
and U16014 (N_16014,N_11156,N_12151);
nand U16015 (N_16015,N_10388,N_10470);
and U16016 (N_16016,N_14090,N_10069);
or U16017 (N_16017,N_14185,N_14666);
nand U16018 (N_16018,N_12888,N_10148);
nor U16019 (N_16019,N_13902,N_13259);
nand U16020 (N_16020,N_12148,N_14564);
and U16021 (N_16021,N_14969,N_12253);
nor U16022 (N_16022,N_12504,N_10695);
nor U16023 (N_16023,N_12142,N_14435);
nor U16024 (N_16024,N_14093,N_11835);
nor U16025 (N_16025,N_12381,N_13621);
nand U16026 (N_16026,N_11235,N_12309);
and U16027 (N_16027,N_10496,N_13312);
nand U16028 (N_16028,N_13474,N_11861);
nor U16029 (N_16029,N_13222,N_10769);
or U16030 (N_16030,N_10314,N_11622);
and U16031 (N_16031,N_10366,N_11281);
nand U16032 (N_16032,N_14018,N_12436);
or U16033 (N_16033,N_14505,N_12661);
or U16034 (N_16034,N_11285,N_12254);
and U16035 (N_16035,N_10133,N_12624);
nand U16036 (N_16036,N_10752,N_14879);
and U16037 (N_16037,N_14056,N_13674);
or U16038 (N_16038,N_13026,N_11229);
and U16039 (N_16039,N_10281,N_13215);
nor U16040 (N_16040,N_14194,N_13245);
and U16041 (N_16041,N_11790,N_13593);
nor U16042 (N_16042,N_11134,N_11989);
and U16043 (N_16043,N_11539,N_14885);
nand U16044 (N_16044,N_13690,N_10977);
nand U16045 (N_16045,N_12680,N_12654);
nand U16046 (N_16046,N_14007,N_11141);
nand U16047 (N_16047,N_12054,N_11195);
or U16048 (N_16048,N_12885,N_12750);
and U16049 (N_16049,N_10257,N_12377);
nand U16050 (N_16050,N_10819,N_13217);
or U16051 (N_16051,N_14306,N_12789);
nor U16052 (N_16052,N_10748,N_12882);
and U16053 (N_16053,N_14462,N_13227);
or U16054 (N_16054,N_11807,N_13842);
nor U16055 (N_16055,N_11143,N_13462);
or U16056 (N_16056,N_14864,N_14157);
nor U16057 (N_16057,N_10975,N_10051);
and U16058 (N_16058,N_12157,N_13883);
or U16059 (N_16059,N_11334,N_13756);
or U16060 (N_16060,N_14859,N_12897);
or U16061 (N_16061,N_10791,N_13995);
or U16062 (N_16062,N_10355,N_11392);
xnor U16063 (N_16063,N_13311,N_14915);
nand U16064 (N_16064,N_13540,N_11062);
nor U16065 (N_16065,N_12975,N_12878);
or U16066 (N_16066,N_13866,N_13346);
nand U16067 (N_16067,N_10518,N_11511);
or U16068 (N_16068,N_14922,N_14201);
nand U16069 (N_16069,N_12522,N_12958);
or U16070 (N_16070,N_12559,N_10435);
and U16071 (N_16071,N_13000,N_12948);
nor U16072 (N_16072,N_14830,N_11551);
nand U16073 (N_16073,N_11776,N_12686);
or U16074 (N_16074,N_13425,N_14588);
and U16075 (N_16075,N_12027,N_14688);
nand U16076 (N_16076,N_14192,N_13260);
or U16077 (N_16077,N_13882,N_12114);
and U16078 (N_16078,N_11376,N_11682);
or U16079 (N_16079,N_13100,N_11457);
and U16080 (N_16080,N_13945,N_12752);
nand U16081 (N_16081,N_12018,N_11726);
nor U16082 (N_16082,N_14240,N_11157);
nor U16083 (N_16083,N_13655,N_13919);
and U16084 (N_16084,N_10682,N_10193);
or U16085 (N_16085,N_12147,N_10245);
and U16086 (N_16086,N_13917,N_10668);
or U16087 (N_16087,N_12419,N_11518);
or U16088 (N_16088,N_13136,N_12695);
and U16089 (N_16089,N_12395,N_10524);
nor U16090 (N_16090,N_11368,N_13040);
and U16091 (N_16091,N_13725,N_12059);
and U16092 (N_16092,N_13192,N_11022);
or U16093 (N_16093,N_11244,N_14899);
nor U16094 (N_16094,N_11668,N_11944);
and U16095 (N_16095,N_12015,N_14705);
nor U16096 (N_16096,N_12123,N_10512);
xnor U16097 (N_16097,N_12760,N_14022);
nor U16098 (N_16098,N_12439,N_13030);
or U16099 (N_16099,N_10510,N_14137);
and U16100 (N_16100,N_14082,N_11378);
xor U16101 (N_16101,N_11384,N_13357);
nand U16102 (N_16102,N_11221,N_11309);
nor U16103 (N_16103,N_10261,N_14798);
or U16104 (N_16104,N_11815,N_10246);
nand U16105 (N_16105,N_12965,N_12201);
xor U16106 (N_16106,N_12186,N_14668);
and U16107 (N_16107,N_12083,N_11934);
and U16108 (N_16108,N_13392,N_10781);
nor U16109 (N_16109,N_11085,N_12751);
nor U16110 (N_16110,N_10765,N_14732);
or U16111 (N_16111,N_12862,N_12817);
and U16112 (N_16112,N_12093,N_12204);
nor U16113 (N_16113,N_13003,N_10952);
and U16114 (N_16114,N_13132,N_12763);
nand U16115 (N_16115,N_13067,N_14271);
nor U16116 (N_16116,N_10642,N_14502);
and U16117 (N_16117,N_11684,N_14070);
nor U16118 (N_16118,N_13181,N_10490);
or U16119 (N_16119,N_10260,N_13604);
nor U16120 (N_16120,N_10687,N_14323);
and U16121 (N_16121,N_11523,N_14491);
nor U16122 (N_16122,N_10081,N_14419);
nor U16123 (N_16123,N_12004,N_14771);
or U16124 (N_16124,N_10071,N_13813);
nor U16125 (N_16125,N_12836,N_13121);
nand U16126 (N_16126,N_12840,N_13148);
and U16127 (N_16127,N_13812,N_10754);
and U16128 (N_16128,N_10384,N_10379);
and U16129 (N_16129,N_10262,N_12348);
nor U16130 (N_16130,N_11329,N_10811);
nor U16131 (N_16131,N_10211,N_10651);
nor U16132 (N_16132,N_11407,N_12274);
nor U16133 (N_16133,N_14297,N_14778);
and U16134 (N_16134,N_14551,N_14234);
and U16135 (N_16135,N_13795,N_11501);
nor U16136 (N_16136,N_13017,N_12313);
nor U16137 (N_16137,N_14755,N_11374);
and U16138 (N_16138,N_11115,N_13746);
and U16139 (N_16139,N_14661,N_13068);
or U16140 (N_16140,N_14076,N_10163);
xnor U16141 (N_16141,N_12263,N_10614);
nor U16142 (N_16142,N_12514,N_13523);
and U16143 (N_16143,N_12032,N_14433);
nor U16144 (N_16144,N_11515,N_12610);
nor U16145 (N_16145,N_12574,N_13050);
xnor U16146 (N_16146,N_12989,N_10315);
nand U16147 (N_16147,N_12452,N_10135);
nand U16148 (N_16148,N_13789,N_10551);
nand U16149 (N_16149,N_10611,N_14965);
or U16150 (N_16150,N_10187,N_14023);
or U16151 (N_16151,N_13261,N_10783);
nor U16152 (N_16152,N_12639,N_10118);
or U16153 (N_16153,N_13097,N_10616);
or U16154 (N_16154,N_12001,N_10003);
or U16155 (N_16155,N_11832,N_11966);
or U16156 (N_16156,N_14876,N_14207);
nand U16157 (N_16157,N_14516,N_14687);
nor U16158 (N_16158,N_11586,N_13358);
and U16159 (N_16159,N_11437,N_14312);
nand U16160 (N_16160,N_13206,N_12898);
nor U16161 (N_16161,N_11604,N_14287);
nand U16162 (N_16162,N_13198,N_14476);
and U16163 (N_16163,N_11705,N_12511);
nand U16164 (N_16164,N_10620,N_13125);
nand U16165 (N_16165,N_14032,N_14344);
nor U16166 (N_16166,N_13247,N_11127);
nand U16167 (N_16167,N_13609,N_13912);
nor U16168 (N_16168,N_13426,N_11977);
or U16169 (N_16169,N_12275,N_13254);
nor U16170 (N_16170,N_13651,N_12638);
xnor U16171 (N_16171,N_11564,N_13785);
or U16172 (N_16172,N_11962,N_11103);
nand U16173 (N_16173,N_11823,N_11173);
nor U16174 (N_16174,N_12757,N_10637);
nand U16175 (N_16175,N_14700,N_11844);
nand U16176 (N_16176,N_14877,N_14063);
nor U16177 (N_16177,N_13726,N_11325);
or U16178 (N_16178,N_12097,N_14127);
nand U16179 (N_16179,N_12367,N_10564);
nand U16180 (N_16180,N_10491,N_14973);
nand U16181 (N_16181,N_14298,N_14203);
nor U16182 (N_16182,N_10945,N_10904);
or U16183 (N_16183,N_12429,N_12671);
nand U16184 (N_16184,N_13354,N_12324);
and U16185 (N_16185,N_11428,N_13514);
or U16186 (N_16186,N_14786,N_12799);
and U16187 (N_16187,N_13307,N_12003);
nor U16188 (N_16188,N_11858,N_14241);
nor U16189 (N_16189,N_12558,N_14513);
and U16190 (N_16190,N_11868,N_10075);
or U16191 (N_16191,N_12462,N_13913);
and U16192 (N_16192,N_10517,N_10572);
nand U16193 (N_16193,N_14767,N_11558);
nand U16194 (N_16194,N_11420,N_14812);
nand U16195 (N_16195,N_10178,N_11956);
nor U16196 (N_16196,N_11400,N_13664);
nand U16197 (N_16197,N_14373,N_10562);
and U16198 (N_16198,N_10929,N_11904);
nor U16199 (N_16199,N_11254,N_10269);
or U16200 (N_16200,N_13605,N_13224);
or U16201 (N_16201,N_14232,N_13313);
or U16202 (N_16202,N_11338,N_14163);
and U16203 (N_16203,N_13472,N_11533);
nand U16204 (N_16204,N_14334,N_10550);
and U16205 (N_16205,N_10065,N_14225);
and U16206 (N_16206,N_13950,N_10828);
and U16207 (N_16207,N_12781,N_10890);
or U16208 (N_16208,N_11280,N_13489);
and U16209 (N_16209,N_10158,N_13671);
or U16210 (N_16210,N_13982,N_12857);
or U16211 (N_16211,N_11126,N_13925);
and U16212 (N_16212,N_11506,N_13636);
nand U16213 (N_16213,N_10717,N_12354);
nand U16214 (N_16214,N_13109,N_10170);
nor U16215 (N_16215,N_14001,N_11169);
nand U16216 (N_16216,N_12131,N_12503);
or U16217 (N_16217,N_14621,N_12182);
nor U16218 (N_16218,N_11881,N_14105);
and U16219 (N_16219,N_11249,N_11896);
nand U16220 (N_16220,N_13562,N_14833);
nor U16221 (N_16221,N_10387,N_12921);
nand U16222 (N_16222,N_11712,N_10561);
nor U16223 (N_16223,N_14012,N_12356);
nor U16224 (N_16224,N_12709,N_10806);
nand U16225 (N_16225,N_11597,N_12026);
or U16226 (N_16226,N_12160,N_12047);
nand U16227 (N_16227,N_13681,N_11724);
or U16228 (N_16228,N_10483,N_11469);
and U16229 (N_16229,N_14745,N_12141);
nor U16230 (N_16230,N_13976,N_11129);
nand U16231 (N_16231,N_11027,N_14555);
nand U16232 (N_16232,N_10399,N_10511);
and U16233 (N_16233,N_11052,N_12400);
nor U16234 (N_16234,N_11609,N_13750);
and U16235 (N_16235,N_13708,N_14589);
or U16236 (N_16236,N_14503,N_14412);
nand U16237 (N_16237,N_11920,N_11088);
nand U16238 (N_16238,N_14228,N_11442);
nor U16239 (N_16239,N_14655,N_13175);
or U16240 (N_16240,N_12974,N_11709);
or U16241 (N_16241,N_13943,N_14857);
and U16242 (N_16242,N_11549,N_12714);
nor U16243 (N_16243,N_13234,N_11914);
or U16244 (N_16244,N_11780,N_10057);
and U16245 (N_16245,N_11029,N_12319);
or U16246 (N_16246,N_10808,N_11704);
nor U16247 (N_16247,N_14809,N_11953);
nor U16248 (N_16248,N_12688,N_13723);
nand U16249 (N_16249,N_12889,N_11774);
nand U16250 (N_16250,N_13516,N_14363);
nand U16251 (N_16251,N_12883,N_14625);
nor U16252 (N_16252,N_12870,N_13888);
nand U16253 (N_16253,N_10630,N_12962);
nor U16254 (N_16254,N_14691,N_10053);
and U16255 (N_16255,N_14067,N_13573);
nand U16256 (N_16256,N_11148,N_13926);
and U16257 (N_16257,N_12991,N_11685);
nand U16258 (N_16258,N_12649,N_12461);
nand U16259 (N_16259,N_10185,N_10504);
and U16260 (N_16260,N_12230,N_14827);
nor U16261 (N_16261,N_11182,N_14639);
and U16262 (N_16262,N_10066,N_10776);
nor U16263 (N_16263,N_10560,N_10383);
or U16264 (N_16264,N_11901,N_10348);
nor U16265 (N_16265,N_10888,N_11980);
and U16266 (N_16266,N_12808,N_10427);
xor U16267 (N_16267,N_10852,N_10232);
or U16268 (N_16268,N_10745,N_12301);
or U16269 (N_16269,N_14337,N_12853);
nor U16270 (N_16270,N_11855,N_14936);
nand U16271 (N_16271,N_14662,N_12391);
nand U16272 (N_16272,N_11958,N_11748);
nand U16273 (N_16273,N_11552,N_13980);
xor U16274 (N_16274,N_12372,N_14599);
nor U16275 (N_16275,N_10190,N_10265);
or U16276 (N_16276,N_11348,N_12434);
nand U16277 (N_16277,N_11380,N_14140);
nor U16278 (N_16278,N_10417,N_11063);
nor U16279 (N_16279,N_14068,N_11145);
and U16280 (N_16280,N_14933,N_11160);
or U16281 (N_16281,N_11470,N_12587);
or U16282 (N_16282,N_11105,N_11412);
or U16283 (N_16283,N_12081,N_10149);
or U16284 (N_16284,N_13252,N_14657);
nor U16285 (N_16285,N_13875,N_14319);
nand U16286 (N_16286,N_12070,N_13009);
nand U16287 (N_16287,N_14958,N_14638);
and U16288 (N_16288,N_14295,N_11274);
or U16289 (N_16289,N_14442,N_11556);
and U16290 (N_16290,N_13073,N_11755);
and U16291 (N_16291,N_10443,N_13989);
and U16292 (N_16292,N_13291,N_14133);
nor U16293 (N_16293,N_14988,N_10382);
nand U16294 (N_16294,N_12689,N_13478);
nand U16295 (N_16295,N_12488,N_14754);
or U16296 (N_16296,N_12937,N_10502);
nor U16297 (N_16297,N_13576,N_13934);
or U16298 (N_16298,N_14309,N_11800);
or U16299 (N_16299,N_12955,N_12518);
nand U16300 (N_16300,N_13445,N_10734);
nor U16301 (N_16301,N_10297,N_13661);
nor U16302 (N_16302,N_11942,N_11898);
nand U16303 (N_16303,N_14165,N_11694);
and U16304 (N_16304,N_12549,N_12850);
and U16305 (N_16305,N_11054,N_14511);
or U16306 (N_16306,N_12694,N_13033);
nor U16307 (N_16307,N_11877,N_13166);
nand U16308 (N_16308,N_14199,N_11538);
nor U16309 (N_16309,N_11936,N_14183);
or U16310 (N_16310,N_13918,N_12726);
or U16311 (N_16311,N_12720,N_13032);
and U16312 (N_16312,N_10444,N_12497);
nor U16313 (N_16313,N_10514,N_14409);
nor U16314 (N_16314,N_10253,N_10151);
and U16315 (N_16315,N_13889,N_11979);
nand U16316 (N_16316,N_12135,N_14752);
or U16317 (N_16317,N_13243,N_13001);
or U16318 (N_16318,N_11567,N_10954);
xor U16319 (N_16319,N_11213,N_13015);
or U16320 (N_16320,N_10636,N_14326);
nand U16321 (N_16321,N_12567,N_11344);
nand U16322 (N_16322,N_14231,N_12433);
or U16323 (N_16323,N_11095,N_12809);
and U16324 (N_16324,N_10725,N_14673);
or U16325 (N_16325,N_13743,N_12438);
or U16326 (N_16326,N_10239,N_10992);
nand U16327 (N_16327,N_11493,N_11326);
or U16328 (N_16328,N_14800,N_10991);
or U16329 (N_16329,N_13126,N_11812);
nor U16330 (N_16330,N_14355,N_10947);
nand U16331 (N_16331,N_12349,N_14117);
and U16332 (N_16332,N_10546,N_11241);
nand U16333 (N_16333,N_13161,N_12094);
nor U16334 (N_16334,N_14762,N_14058);
and U16335 (N_16335,N_12849,N_11702);
xnor U16336 (N_16336,N_10224,N_12644);
nand U16337 (N_16337,N_13279,N_14490);
nand U16338 (N_16338,N_13265,N_14849);
or U16339 (N_16339,N_14397,N_13769);
nor U16340 (N_16340,N_14811,N_13729);
nor U16341 (N_16341,N_14917,N_11792);
and U16342 (N_16342,N_10027,N_10722);
or U16343 (N_16343,N_12951,N_14389);
xor U16344 (N_16344,N_13168,N_10480);
or U16345 (N_16345,N_13878,N_13042);
and U16346 (N_16346,N_11164,N_14043);
or U16347 (N_16347,N_10124,N_14631);
or U16348 (N_16348,N_12185,N_11167);
nand U16349 (N_16349,N_11162,N_14853);
nor U16350 (N_16350,N_13078,N_14887);
nor U16351 (N_16351,N_11751,N_13203);
nor U16352 (N_16352,N_10229,N_12845);
nand U16353 (N_16353,N_13099,N_11037);
or U16354 (N_16354,N_14195,N_14002);
nand U16355 (N_16355,N_13475,N_12192);
or U16356 (N_16356,N_14527,N_12568);
and U16357 (N_16357,N_10445,N_11769);
nand U16358 (N_16358,N_13781,N_10337);
nand U16359 (N_16359,N_14253,N_11204);
xor U16360 (N_16360,N_11128,N_10129);
and U16361 (N_16361,N_13755,N_10938);
nor U16362 (N_16362,N_11217,N_11084);
nand U16363 (N_16363,N_10290,N_11845);
or U16364 (N_16364,N_13551,N_12417);
nor U16365 (N_16365,N_10180,N_10083);
nand U16366 (N_16366,N_11417,N_11693);
or U16367 (N_16367,N_14362,N_10016);
and U16368 (N_16368,N_14635,N_13610);
and U16369 (N_16369,N_11592,N_10905);
nand U16370 (N_16370,N_13272,N_10300);
nand U16371 (N_16371,N_12653,N_14721);
xor U16372 (N_16372,N_13862,N_13997);
and U16373 (N_16373,N_14532,N_10993);
nand U16374 (N_16374,N_13292,N_13240);
or U16375 (N_16375,N_11492,N_12851);
nand U16376 (N_16376,N_14795,N_11360);
and U16377 (N_16377,N_10391,N_12693);
and U16378 (N_16378,N_10996,N_14907);
xnor U16379 (N_16379,N_12930,N_12969);
nor U16380 (N_16380,N_11276,N_13640);
or U16381 (N_16381,N_13108,N_12321);
nand U16382 (N_16382,N_10883,N_14584);
nor U16383 (N_16383,N_14594,N_13703);
or U16384 (N_16384,N_12338,N_11447);
nand U16385 (N_16385,N_14602,N_13559);
or U16386 (N_16386,N_11448,N_12679);
nor U16387 (N_16387,N_13315,N_13615);
nor U16388 (N_16388,N_13904,N_14694);
nor U16389 (N_16389,N_12212,N_12476);
and U16390 (N_16390,N_12296,N_10830);
nor U16391 (N_16391,N_13991,N_11003);
nand U16392 (N_16392,N_13622,N_12077);
nor U16393 (N_16393,N_10181,N_11058);
or U16394 (N_16394,N_13151,N_10240);
and U16395 (N_16395,N_13449,N_10932);
and U16396 (N_16396,N_14154,N_14072);
or U16397 (N_16397,N_10837,N_14994);
nand U16398 (N_16398,N_13327,N_13864);
or U16399 (N_16399,N_13319,N_10627);
nor U16400 (N_16400,N_11282,N_12570);
nor U16401 (N_16401,N_14026,N_10110);
and U16402 (N_16402,N_10346,N_13442);
nand U16403 (N_16403,N_10982,N_12911);
and U16404 (N_16404,N_10409,N_10202);
or U16405 (N_16405,N_13492,N_14640);
nand U16406 (N_16406,N_10531,N_14062);
and U16407 (N_16407,N_13055,N_13330);
nand U16408 (N_16408,N_11001,N_10762);
and U16409 (N_16409,N_13476,N_13218);
nor U16410 (N_16410,N_14108,N_11885);
and U16411 (N_16411,N_14520,N_12765);
nand U16412 (N_16412,N_14044,N_12126);
nor U16413 (N_16413,N_12668,N_11471);
nand U16414 (N_16414,N_12180,N_10703);
and U16415 (N_16415,N_12533,N_10171);
nor U16416 (N_16416,N_13618,N_12020);
nor U16417 (N_16417,N_14577,N_11123);
nand U16418 (N_16418,N_11072,N_13567);
and U16419 (N_16419,N_10136,N_12776);
or U16420 (N_16420,N_13858,N_11077);
or U16421 (N_16421,N_10663,N_11462);
or U16422 (N_16422,N_11478,N_13759);
and U16423 (N_16423,N_13911,N_14781);
nor U16424 (N_16424,N_12600,N_14948);
or U16425 (N_16425,N_11892,N_10408);
nand U16426 (N_16426,N_11066,N_11838);
or U16427 (N_16427,N_12043,N_13244);
nand U16428 (N_16428,N_11949,N_12283);
nor U16429 (N_16429,N_13596,N_14617);
and U16430 (N_16430,N_11596,N_13277);
nand U16431 (N_16431,N_14934,N_12084);
and U16432 (N_16432,N_11432,N_12202);
and U16433 (N_16433,N_13978,N_13935);
nor U16434 (N_16434,N_12039,N_14308);
nor U16435 (N_16435,N_10223,N_13625);
nor U16436 (N_16436,N_13284,N_13117);
and U16437 (N_16437,N_11612,N_12128);
and U16438 (N_16438,N_12982,N_11816);
and U16439 (N_16439,N_11565,N_13394);
nor U16440 (N_16440,N_11223,N_12806);
and U16441 (N_16441,N_14024,N_13967);
nand U16442 (N_16442,N_14370,N_13975);
nand U16443 (N_16443,N_10024,N_14883);
or U16444 (N_16444,N_11729,N_14632);
nor U16445 (N_16445,N_14813,N_13454);
or U16446 (N_16446,N_12516,N_11672);
and U16447 (N_16447,N_11242,N_14034);
nand U16448 (N_16448,N_11576,N_12295);
or U16449 (N_16449,N_10089,N_11860);
nand U16450 (N_16450,N_12797,N_11387);
xor U16451 (N_16451,N_14374,N_12562);
nor U16452 (N_16452,N_11657,N_13722);
nor U16453 (N_16453,N_14726,N_12761);
nor U16454 (N_16454,N_10528,N_10701);
or U16455 (N_16455,N_11075,N_10589);
or U16456 (N_16456,N_14340,N_10877);
nor U16457 (N_16457,N_11064,N_14071);
nand U16458 (N_16458,N_14717,N_13163);
nand U16459 (N_16459,N_10031,N_13414);
and U16460 (N_16460,N_14226,N_14481);
nor U16461 (N_16461,N_10013,N_11869);
nor U16462 (N_16462,N_14277,N_13891);
nand U16463 (N_16463,N_14080,N_12333);
and U16464 (N_16464,N_14596,N_13257);
or U16465 (N_16465,N_13119,N_11589);
xor U16466 (N_16466,N_14390,N_10569);
nand U16467 (N_16467,N_13496,N_12565);
and U16468 (N_16468,N_13273,N_11955);
or U16469 (N_16469,N_11209,N_12681);
or U16470 (N_16470,N_12844,N_10448);
nor U16471 (N_16471,N_12010,N_10892);
nor U16472 (N_16472,N_14970,N_10660);
nand U16473 (N_16473,N_13992,N_11937);
or U16474 (N_16474,N_12966,N_14320);
and U16475 (N_16475,N_11342,N_11536);
or U16476 (N_16476,N_14648,N_13598);
nor U16477 (N_16477,N_12717,N_14382);
nor U16478 (N_16478,N_10869,N_10055);
nor U16479 (N_16479,N_11671,N_10441);
nor U16480 (N_16480,N_13362,N_12280);
and U16481 (N_16481,N_13463,N_14099);
xnor U16482 (N_16482,N_14318,N_10493);
and U16483 (N_16483,N_11588,N_13784);
and U16484 (N_16484,N_10714,N_12501);
and U16485 (N_16485,N_10492,N_11872);
nand U16486 (N_16486,N_14339,N_12110);
nand U16487 (N_16487,N_14138,N_14737);
nor U16488 (N_16488,N_10583,N_10559);
nand U16489 (N_16489,N_14675,N_13583);
or U16490 (N_16490,N_12901,N_11646);
nand U16491 (N_16491,N_11366,N_11562);
nor U16492 (N_16492,N_11993,N_11578);
and U16493 (N_16493,N_13286,N_11396);
nor U16494 (N_16494,N_13294,N_14506);
and U16495 (N_16495,N_14436,N_10212);
and U16496 (N_16496,N_11136,N_13932);
nor U16497 (N_16497,N_13668,N_13731);
nor U16498 (N_16498,N_13276,N_11297);
nand U16499 (N_16499,N_14837,N_12014);
or U16500 (N_16500,N_11434,N_11863);
or U16501 (N_16501,N_14280,N_13299);
and U16502 (N_16502,N_14084,N_12050);
nor U16503 (N_16503,N_14332,N_13653);
or U16504 (N_16504,N_13391,N_13114);
nor U16505 (N_16505,N_10738,N_10272);
or U16506 (N_16506,N_12702,N_13916);
and U16507 (N_16507,N_13281,N_14895);
nor U16508 (N_16508,N_10474,N_12382);
nor U16509 (N_16509,N_14223,N_10254);
xnor U16510 (N_16510,N_14135,N_13955);
nor U16511 (N_16511,N_14172,N_12404);
and U16512 (N_16512,N_10824,N_12941);
or U16513 (N_16513,N_13742,N_12795);
or U16514 (N_16514,N_13184,N_14420);
or U16515 (N_16515,N_10363,N_13811);
nor U16516 (N_16516,N_12118,N_14874);
and U16517 (N_16517,N_13229,N_13534);
or U16518 (N_16518,N_13529,N_10826);
xnor U16519 (N_16519,N_11487,N_12929);
nor U16520 (N_16520,N_14438,N_11012);
nor U16521 (N_16521,N_12127,N_10429);
nor U16522 (N_16522,N_11797,N_14620);
nand U16523 (N_16523,N_11788,N_14701);
and U16524 (N_16524,N_12117,N_11073);
and U16525 (N_16525,N_14772,N_14038);
nor U16526 (N_16526,N_13268,N_14317);
nand U16527 (N_16527,N_12708,N_14321);
nand U16528 (N_16528,N_10449,N_12387);
and U16529 (N_16529,N_10019,N_12715);
nand U16530 (N_16530,N_14368,N_13798);
nand U16531 (N_16531,N_10340,N_14923);
or U16532 (N_16532,N_11625,N_12115);
and U16533 (N_16533,N_10505,N_14557);
nor U16534 (N_16534,N_14200,N_11133);
or U16535 (N_16535,N_10197,N_10008);
nor U16536 (N_16536,N_10354,N_12796);
nand U16537 (N_16537,N_10454,N_12791);
nor U16538 (N_16538,N_10756,N_11884);
and U16539 (N_16539,N_14122,N_13386);
nor U16540 (N_16540,N_12942,N_13209);
nand U16541 (N_16541,N_14626,N_12153);
and U16542 (N_16542,N_11959,N_12894);
or U16543 (N_16543,N_11833,N_10285);
or U16544 (N_16544,N_10915,N_10911);
or U16545 (N_16545,N_12040,N_10341);
and U16546 (N_16546,N_11225,N_10631);
nand U16547 (N_16547,N_13803,N_13197);
and U16548 (N_16548,N_14761,N_11131);
or U16549 (N_16549,N_11637,N_13278);
and U16550 (N_16550,N_13187,N_11918);
and U16551 (N_16551,N_10404,N_12211);
nor U16552 (N_16552,N_14107,N_12682);
or U16553 (N_16553,N_13591,N_10617);
and U16554 (N_16554,N_10182,N_11703);
and U16555 (N_16555,N_11197,N_10294);
nor U16556 (N_16556,N_11100,N_13644);
nand U16557 (N_16557,N_12389,N_12457);
nor U16558 (N_16558,N_11847,N_14175);
nand U16559 (N_16559,N_10131,N_14856);
and U16560 (N_16560,N_14141,N_14597);
or U16561 (N_16561,N_10934,N_12169);
or U16562 (N_16562,N_12392,N_13799);
and U16563 (N_16563,N_13797,N_13974);
nand U16564 (N_16564,N_12386,N_11125);
nand U16565 (N_16565,N_13303,N_14566);
nor U16566 (N_16566,N_11572,N_11531);
and U16567 (N_16567,N_14015,N_12342);
and U16568 (N_16568,N_10298,N_13585);
nor U16569 (N_16569,N_11255,N_14448);
and U16570 (N_16570,N_10585,N_12264);
and U16571 (N_16571,N_11525,N_12625);
nand U16572 (N_16572,N_10113,N_11595);
nor U16573 (N_16573,N_12586,N_11019);
xnor U16574 (N_16574,N_13251,N_14030);
nand U16575 (N_16575,N_10534,N_14565);
nand U16576 (N_16576,N_11491,N_12536);
nor U16577 (N_16577,N_10063,N_12161);
nor U16578 (N_16578,N_10588,N_14568);
nor U16579 (N_16579,N_12490,N_10250);
and U16580 (N_16580,N_12626,N_14932);
and U16581 (N_16581,N_12159,N_11758);
and U16582 (N_16582,N_14892,N_12240);
and U16583 (N_16583,N_10670,N_13985);
nand U16584 (N_16584,N_13829,N_12423);
and U16585 (N_16585,N_12465,N_13683);
nor U16586 (N_16586,N_13076,N_14377);
nand U16587 (N_16587,N_14634,N_14954);
and U16588 (N_16588,N_10988,N_10782);
or U16589 (N_16589,N_11913,N_12124);
nand U16590 (N_16590,N_14112,N_11754);
or U16591 (N_16591,N_10032,N_12396);
or U16592 (N_16592,N_12532,N_14350);
nor U16593 (N_16593,N_13770,N_12952);
nor U16594 (N_16594,N_14145,N_14252);
and U16595 (N_16595,N_10944,N_11226);
or U16596 (N_16596,N_14217,N_12091);
nor U16597 (N_16597,N_11651,N_12842);
or U16598 (N_16598,N_14561,N_11796);
or U16599 (N_16599,N_10044,N_12902);
nand U16600 (N_16600,N_11194,N_12022);
and U16601 (N_16601,N_13366,N_11065);
or U16602 (N_16602,N_12502,N_13137);
nand U16603 (N_16603,N_14416,N_10301);
nor U16604 (N_16604,N_13043,N_13990);
nand U16605 (N_16605,N_14278,N_14552);
nor U16606 (N_16606,N_10724,N_11771);
or U16607 (N_16607,N_12841,N_12250);
nor U16608 (N_16608,N_12713,N_10259);
nor U16609 (N_16609,N_11628,N_13641);
or U16610 (N_16610,N_14401,N_10675);
nand U16611 (N_16611,N_12398,N_10605);
or U16612 (N_16612,N_13490,N_14977);
or U16613 (N_16613,N_11952,N_11336);
or U16614 (N_16614,N_13350,N_14441);
nand U16615 (N_16615,N_13772,N_14770);
nand U16616 (N_16616,N_11009,N_13196);
or U16617 (N_16617,N_13802,N_14016);
and U16618 (N_16618,N_14283,N_11191);
and U16619 (N_16619,N_14064,N_13778);
nor U16620 (N_16620,N_14247,N_14230);
and U16621 (N_16621,N_11346,N_11231);
and U16622 (N_16622,N_10864,N_14265);
and U16623 (N_16623,N_10581,N_12775);
nand U16624 (N_16624,N_11626,N_11652);
or U16625 (N_16625,N_14644,N_13116);
nor U16626 (N_16626,N_10162,N_10208);
xor U16627 (N_16627,N_14572,N_13977);
nand U16628 (N_16628,N_10582,N_10132);
nor U16629 (N_16629,N_13834,N_11499);
and U16630 (N_16630,N_11571,N_11151);
xor U16631 (N_16631,N_10659,N_13411);
and U16632 (N_16632,N_12271,N_14081);
or U16633 (N_16633,N_11808,N_10567);
nor U16634 (N_16634,N_12830,N_14392);
nor U16635 (N_16635,N_14846,N_14839);
nand U16636 (N_16636,N_13164,N_11401);
nor U16637 (N_16637,N_11865,N_14330);
nor U16638 (N_16638,N_12938,N_10014);
or U16639 (N_16639,N_13628,N_14483);
nand U16640 (N_16640,N_10790,N_10410);
nor U16641 (N_16641,N_12640,N_11811);
nor U16642 (N_16642,N_10948,N_14790);
or U16643 (N_16643,N_11116,N_12995);
and U16644 (N_16644,N_11364,N_10026);
and U16645 (N_16645,N_11978,N_14102);
and U16646 (N_16646,N_14347,N_10763);
nand U16647 (N_16647,N_11089,N_14215);
and U16648 (N_16648,N_11728,N_10860);
or U16649 (N_16649,N_14255,N_12731);
and U16650 (N_16650,N_14720,N_12913);
nor U16651 (N_16651,N_14909,N_10402);
or U16652 (N_16652,N_11994,N_11521);
and U16653 (N_16653,N_14328,N_10615);
or U16654 (N_16654,N_11405,N_14674);
and U16655 (N_16655,N_14465,N_10295);
and U16656 (N_16656,N_13936,N_13673);
and U16657 (N_16657,N_10401,N_10865);
nand U16658 (N_16658,N_10248,N_14676);
or U16659 (N_16659,N_12524,N_12046);
nor U16660 (N_16660,N_13105,N_10376);
or U16661 (N_16661,N_10917,N_11208);
and U16662 (N_16662,N_14985,N_12272);
or U16663 (N_16663,N_10459,N_14975);
nand U16664 (N_16664,N_10758,N_10645);
and U16665 (N_16665,N_11328,N_10390);
or U16666 (N_16666,N_13790,N_12588);
or U16667 (N_16667,N_13692,N_10227);
nor U16668 (N_16668,N_11791,N_12788);
nor U16669 (N_16669,N_13432,N_10508);
or U16670 (N_16670,N_12370,N_11559);
nor U16671 (N_16671,N_10184,N_14982);
nand U16672 (N_16672,N_13705,N_12609);
nor U16673 (N_16673,N_12469,N_11598);
and U16674 (N_16674,N_14667,N_14835);
and U16675 (N_16675,N_10554,N_11237);
and U16676 (N_16676,N_13374,N_11383);
or U16677 (N_16677,N_10532,N_13669);
nor U16678 (N_16678,N_13771,N_11650);
or U16679 (N_16679,N_10256,N_11354);
nor U16680 (N_16680,N_11321,N_11168);
and U16681 (N_16681,N_10457,N_14380);
nor U16682 (N_16682,N_13659,N_12416);
or U16683 (N_16683,N_13398,N_10323);
or U16684 (N_16684,N_13527,N_12140);
and U16685 (N_16685,N_10595,N_13417);
or U16686 (N_16686,N_11594,N_11277);
or U16687 (N_16687,N_14850,N_11938);
nand U16688 (N_16688,N_12931,N_13008);
or U16689 (N_16689,N_12477,N_12684);
or U16690 (N_16690,N_13075,N_13845);
or U16691 (N_16691,N_11968,N_12154);
or U16692 (N_16692,N_10650,N_11880);
or U16693 (N_16693,N_13872,N_14212);
and U16694 (N_16694,N_12636,N_11450);
or U16695 (N_16695,N_12697,N_14249);
nand U16696 (N_16696,N_10237,N_13595);
nor U16697 (N_16697,N_13933,N_14658);
and U16698 (N_16698,N_14322,N_13497);
nand U16699 (N_16699,N_10795,N_11292);
nor U16700 (N_16700,N_11999,N_11933);
nor U16701 (N_16701,N_13316,N_13903);
or U16702 (N_16702,N_12190,N_10820);
xnor U16703 (N_16703,N_12105,N_10338);
nor U16704 (N_16704,N_10357,N_12065);
or U16705 (N_16705,N_13046,N_10072);
nor U16706 (N_16706,N_10029,N_10058);
nand U16707 (N_16707,N_12375,N_14650);
and U16708 (N_16708,N_13264,N_12903);
or U16709 (N_16709,N_14575,N_13787);
nand U16710 (N_16710,N_14562,N_11352);
nor U16711 (N_16711,N_11485,N_13447);
or U16712 (N_16712,N_11473,N_10157);
and U16713 (N_16713,N_11681,N_12258);
nor U16714 (N_16714,N_13274,N_14542);
and U16715 (N_16715,N_10538,N_13275);
or U16716 (N_16716,N_11696,N_13174);
nor U16717 (N_16717,N_12566,N_14817);
nor U16718 (N_16718,N_11927,N_13310);
nand U16719 (N_16719,N_10094,N_14618);
and U16720 (N_16720,N_12048,N_12312);
xnor U16721 (N_16721,N_10159,N_10866);
or U16722 (N_16722,N_10967,N_12864);
nand U16723 (N_16723,N_11840,N_12964);
nor U16724 (N_16724,N_12255,N_14522);
or U16725 (N_16725,N_11947,N_12025);
xor U16726 (N_16726,N_13088,N_10844);
and U16727 (N_16727,N_10995,N_10271);
nand U16728 (N_16728,N_12630,N_14956);
nand U16729 (N_16729,N_14609,N_11603);
nor U16730 (N_16730,N_14580,N_11408);
or U16731 (N_16731,N_12871,N_13453);
and U16732 (N_16732,N_11508,N_13341);
or U16733 (N_16733,N_14739,N_12716);
and U16734 (N_16734,N_12137,N_13473);
nor U16735 (N_16735,N_10007,N_14841);
nor U16736 (N_16736,N_11560,N_13881);
or U16737 (N_16737,N_14000,N_10476);
and U16738 (N_16738,N_11415,N_11720);
nor U16739 (N_16739,N_10715,N_11117);
or U16740 (N_16740,N_10335,N_13589);
nand U16741 (N_16741,N_13792,N_11708);
nor U16742 (N_16742,N_11140,N_13186);
or U16743 (N_16743,N_11540,N_12614);
nand U16744 (N_16744,N_10867,N_14386);
and U16745 (N_16745,N_13526,N_11765);
or U16746 (N_16746,N_12176,N_12194);
or U16747 (N_16747,N_13103,N_13322);
and U16748 (N_16748,N_14052,N_10450);
and U16749 (N_16749,N_12627,N_10156);
and U16750 (N_16750,N_11537,N_12453);
or U16751 (N_16751,N_14804,N_12175);
or U16752 (N_16752,N_13093,N_11701);
nand U16753 (N_16753,N_12876,N_10034);
or U16754 (N_16754,N_11638,N_11298);
nand U16755 (N_16755,N_14608,N_11803);
nand U16756 (N_16756,N_14509,N_11069);
nand U16757 (N_16757,N_10176,N_13237);
nor U16758 (N_16758,N_11895,N_12060);
nand U16759 (N_16759,N_11698,N_14096);
nand U16760 (N_16760,N_13344,N_13767);
and U16761 (N_16761,N_13791,N_13479);
or U16762 (N_16762,N_13480,N_14908);
nand U16763 (N_16763,N_11997,N_13786);
nand U16764 (N_16764,N_14610,N_10925);
or U16765 (N_16765,N_14712,N_13924);
nor U16766 (N_16766,N_13793,N_13232);
and U16767 (N_16767,N_12756,N_12582);
or U16768 (N_16768,N_11005,N_12846);
nor U16769 (N_16769,N_11870,N_10994);
or U16770 (N_16770,N_11864,N_14487);
and U16771 (N_16771,N_11957,N_12475);
or U16772 (N_16772,N_10565,N_11370);
nand U16773 (N_16773,N_10556,N_12152);
nand U16774 (N_16774,N_10494,N_14585);
nand U16775 (N_16775,N_12517,N_13014);
or U16776 (N_16776,N_10506,N_13258);
nand U16777 (N_16777,N_13360,N_12563);
and U16778 (N_16778,N_10453,N_11534);
or U16779 (N_16779,N_11068,N_14537);
and U16780 (N_16780,N_13451,N_12801);
xnor U16781 (N_16781,N_13546,N_11613);
nand U16782 (N_16782,N_12994,N_11455);
nand U16783 (N_16783,N_14785,N_11025);
or U16784 (N_16784,N_13488,N_12121);
and U16785 (N_16785,N_14943,N_14366);
and U16786 (N_16786,N_13107,N_14779);
and U16787 (N_16787,N_13825,N_12322);
nand U16788 (N_16788,N_14335,N_13620);
nor U16789 (N_16789,N_10962,N_10090);
nor U16790 (N_16790,N_11440,N_12163);
or U16791 (N_16791,N_14533,N_12494);
or U16792 (N_16792,N_13873,N_11903);
or U16793 (N_16793,N_11178,N_14173);
nand U16794 (N_16794,N_10326,N_13563);
or U16795 (N_16795,N_14627,N_14120);
or U16796 (N_16796,N_11695,N_12246);
or U16797 (N_16797,N_10228,N_12607);
or U16798 (N_16798,N_11138,N_13719);
nand U16799 (N_16799,N_14529,N_13545);
nor U16800 (N_16800,N_10446,N_13607);
and U16801 (N_16801,N_11301,N_14966);
or U16802 (N_16802,N_11256,N_10764);
or U16803 (N_16803,N_11080,N_11391);
nand U16804 (N_16804,N_12843,N_11028);
nor U16805 (N_16805,N_14151,N_10685);
or U16806 (N_16806,N_14033,N_12101);
nand U16807 (N_16807,N_14723,N_14889);
and U16808 (N_16808,N_13306,N_13501);
or U16809 (N_16809,N_12330,N_13780);
nor U16810 (N_16810,N_13579,N_11912);
nor U16811 (N_16811,N_10101,N_10872);
nor U16812 (N_16812,N_14997,N_12241);
or U16813 (N_16813,N_14300,N_11296);
nor U16814 (N_16814,N_10078,N_12073);
nand U16815 (N_16815,N_13996,N_10700);
or U16816 (N_16816,N_13176,N_13667);
nor U16817 (N_16817,N_11476,N_11423);
or U16818 (N_16818,N_12531,N_14299);
nor U16819 (N_16819,N_11361,N_10834);
or U16820 (N_16820,N_11805,N_10891);
and U16821 (N_16821,N_14834,N_14656);
nor U16822 (N_16822,N_10845,N_12972);
nand U16823 (N_16823,N_14036,N_12467);
nand U16824 (N_16824,N_12089,N_13707);
nand U16825 (N_16825,N_11654,N_10085);
xor U16826 (N_16826,N_13140,N_12831);
and U16827 (N_16827,N_13282,N_10095);
nand U16828 (N_16828,N_11541,N_14248);
and U16829 (N_16829,N_14888,N_11422);
and U16830 (N_16830,N_14514,N_12608);
or U16831 (N_16831,N_12664,N_12886);
nand U16832 (N_16832,N_14571,N_11211);
nand U16833 (N_16833,N_13157,N_11078);
nand U16834 (N_16834,N_11184,N_12352);
or U16835 (N_16835,N_12727,N_12704);
xor U16836 (N_16836,N_10103,N_10964);
xnor U16837 (N_16837,N_13065,N_10540);
and U16838 (N_16838,N_11857,N_11016);
xnor U16839 (N_16839,N_14186,N_12735);
nand U16840 (N_16840,N_11917,N_11299);
nand U16841 (N_16841,N_12794,N_11543);
nand U16842 (N_16842,N_13433,N_10128);
nor U16843 (N_16843,N_12783,N_10464);
or U16844 (N_16844,N_12363,N_11614);
or U16845 (N_16845,N_12900,N_12592);
and U16846 (N_16846,N_10785,N_12483);
and U16847 (N_16847,N_11275,N_11772);
nor U16848 (N_16848,N_11893,N_11819);
nor U16849 (N_16849,N_11283,N_13051);
nor U16850 (N_16850,N_11002,N_12307);
nor U16851 (N_16851,N_13885,N_12405);
or U16852 (N_16852,N_11441,N_13248);
nor U16853 (N_16853,N_11202,N_12981);
and U16854 (N_16854,N_11243,N_13044);
nand U16855 (N_16855,N_12891,N_14246);
nor U16856 (N_16856,N_13775,N_10263);
or U16857 (N_16857,N_14177,N_14459);
nand U16858 (N_16858,N_11891,N_13800);
nand U16859 (N_16859,N_11757,N_14780);
nor U16860 (N_16860,N_11385,N_12208);
and U16861 (N_16861,N_14021,N_10936);
nand U16862 (N_16862,N_12195,N_13734);
nand U16863 (N_16863,N_13714,N_11107);
nand U16864 (N_16864,N_14703,N_14764);
xnor U16865 (N_16865,N_10760,N_14672);
nand U16866 (N_16866,N_12401,N_10545);
nand U16867 (N_16867,N_11144,N_14179);
and U16868 (N_16868,N_10009,N_14818);
and U16869 (N_16869,N_14595,N_10673);
xor U16870 (N_16870,N_10788,N_11856);
nor U16871 (N_16871,N_11634,N_13384);
nor U16872 (N_16872,N_14592,N_14352);
and U16873 (N_16873,N_13710,N_13343);
and U16874 (N_16874,N_12139,N_14311);
nor U16875 (N_16875,N_13378,N_13031);
and U16876 (N_16876,N_13951,N_11530);
or U16877 (N_16877,N_14260,N_14591);
nor U16878 (N_16878,N_10264,N_10825);
and U16879 (N_16879,N_14685,N_12854);
nand U16880 (N_16880,N_13920,N_14729);
nor U16881 (N_16881,N_14210,N_12736);
and U16882 (N_16882,N_11809,N_12339);
and U16883 (N_16883,N_11097,N_11973);
and U16884 (N_16884,N_10958,N_10267);
and U16885 (N_16885,N_12633,N_13922);
nor U16886 (N_16886,N_12552,N_10759);
or U16887 (N_16887,N_13676,N_12005);
and U16888 (N_16888,N_14794,N_13694);
and U16889 (N_16889,N_10596,N_11854);
or U16890 (N_16890,N_13531,N_13439);
or U16891 (N_16891,N_11655,N_10345);
and U16892 (N_16892,N_14999,N_11375);
and U16893 (N_16893,N_10115,N_14289);
or U16894 (N_16894,N_10664,N_13966);
or U16895 (N_16895,N_13730,N_12156);
and U16896 (N_16896,N_13895,N_14836);
or U16897 (N_16897,N_14147,N_11253);
xor U16898 (N_16898,N_10672,N_10462);
nor U16899 (N_16899,N_13452,N_11313);
nor U16900 (N_16900,N_13214,N_11928);
nor U16901 (N_16901,N_13305,N_14357);
nand U16902 (N_16902,N_13855,N_14159);
and U16903 (N_16903,N_14823,N_10322);
nor U16904 (N_16904,N_10737,N_10812);
and U16905 (N_16905,N_10405,N_12954);
nor U16906 (N_16906,N_13647,N_12521);
and U16907 (N_16907,N_11266,N_12178);
or U16908 (N_16908,N_12666,N_14753);
nor U16909 (N_16909,N_10091,N_11303);
nand U16910 (N_16910,N_11873,N_11503);
nand U16911 (N_16911,N_14749,N_11155);
nor U16912 (N_16912,N_14515,N_10238);
and U16913 (N_16913,N_12286,N_11789);
nor U16914 (N_16914,N_10746,N_10597);
or U16915 (N_16915,N_11502,N_12579);
nor U16916 (N_16916,N_12035,N_14777);
nand U16917 (N_16917,N_10643,N_10070);
nand U16918 (N_16918,N_13194,N_13128);
nand U16919 (N_16919,N_11566,N_13794);
nand U16920 (N_16920,N_13939,N_12430);
xnor U16921 (N_16921,N_10603,N_11132);
nor U16922 (N_16922,N_14237,N_12723);
and U16923 (N_16923,N_14005,N_10154);
nand U16924 (N_16924,N_11135,N_10048);
nand U16925 (N_16925,N_11310,N_12103);
and U16926 (N_16926,N_13269,N_12577);
nand U16927 (N_16927,N_12008,N_10691);
and U16928 (N_16928,N_12658,N_12884);
and U16929 (N_16929,N_10728,N_13409);
and U16930 (N_16930,N_10461,N_13896);
or U16931 (N_16931,N_13738,N_14010);
and U16932 (N_16932,N_10252,N_14972);
nand U16933 (N_16933,N_14256,N_14101);
nand U16934 (N_16934,N_10697,N_13597);
nand U16935 (N_16935,N_11096,N_11199);
and U16936 (N_16936,N_11587,N_14324);
nand U16937 (N_16937,N_12133,N_10859);
or U16938 (N_16938,N_11744,N_12440);
nand U16939 (N_16939,N_10460,N_14087);
or U16940 (N_16940,N_14910,N_12764);
nor U16941 (N_16941,N_10786,N_12278);
and U16942 (N_16942,N_12306,N_13828);
or U16943 (N_16943,N_14126,N_13035);
or U16944 (N_16944,N_14037,N_13524);
and U16945 (N_16945,N_13402,N_12996);
xor U16946 (N_16946,N_11286,N_10418);
nor U16947 (N_16947,N_11911,N_14647);
nand U16948 (N_16948,N_10590,N_12238);
and U16949 (N_16949,N_10902,N_14536);
and U16950 (N_16950,N_10592,N_11295);
and U16951 (N_16951,N_10487,N_10200);
or U16952 (N_16952,N_14756,N_13334);
and U16953 (N_16953,N_11677,N_10230);
and U16954 (N_16954,N_10365,N_13349);
or U16955 (N_16955,N_13804,N_13532);
or U16956 (N_16956,N_10509,N_14929);
or U16957 (N_16957,N_10646,N_14716);
and U16958 (N_16958,N_14736,N_12642);
nand U16959 (N_16959,N_11307,N_14569);
or U16960 (N_16960,N_12515,N_13039);
and U16961 (N_16961,N_12113,N_12368);
and U16962 (N_16962,N_12300,N_13491);
nand U16963 (N_16963,N_10953,N_10165);
and U16964 (N_16964,N_10693,N_10336);
or U16965 (N_16965,N_12247,N_12420);
nand U16966 (N_16966,N_12632,N_10060);
and U16967 (N_16967,N_12824,N_14220);
and U16968 (N_16968,N_12785,N_11908);
nor U16969 (N_16969,N_11445,N_12031);
nor U16970 (N_16970,N_13340,N_12340);
nor U16971 (N_16971,N_13112,N_11528);
and U16972 (N_16972,N_12648,N_13662);
or U16973 (N_16973,N_13859,N_12879);
or U16974 (N_16974,N_11083,N_13498);
nand U16975 (N_16975,N_10479,N_13288);
or U16976 (N_16976,N_13377,N_13971);
nand U16977 (N_16977,N_11239,N_13419);
or U16978 (N_16978,N_10665,N_13469);
nand U16979 (N_16979,N_11831,N_10324);
nand U16980 (N_16980,N_11674,N_10503);
and U16981 (N_16981,N_12245,N_14156);
nand U16982 (N_16982,N_14947,N_12122);
xor U16983 (N_16983,N_12066,N_10854);
nor U16984 (N_16984,N_13289,N_13348);
and U16985 (N_16985,N_14941,N_11032);
and U16986 (N_16986,N_11269,N_11497);
nor U16987 (N_16987,N_14302,N_12355);
or U16988 (N_16988,N_14375,N_11320);
nand U16989 (N_16989,N_12547,N_13993);
and U16990 (N_16990,N_10879,N_11294);
nor U16991 (N_16991,N_10780,N_14089);
and U16992 (N_16992,N_13448,N_14735);
or U16993 (N_16993,N_14125,N_13852);
nor U16994 (N_16994,N_11110,N_12539);
and U16995 (N_16995,N_12146,N_12062);
nand U16996 (N_16996,N_12940,N_11732);
or U16997 (N_16997,N_11779,N_10875);
or U16998 (N_16998,N_14622,N_14792);
nand U16999 (N_16999,N_14364,N_12085);
nand U17000 (N_17000,N_10134,N_11846);
nand U17001 (N_17001,N_14546,N_14838);
nand U17002 (N_17002,N_12002,N_10604);
nand U17003 (N_17003,N_13502,N_12963);
nand U17004 (N_17004,N_11601,N_12337);
nand U17005 (N_17005,N_13129,N_11631);
nand U17006 (N_17006,N_11015,N_12881);
nor U17007 (N_17007,N_13632,N_11053);
nand U17008 (N_17008,N_14906,N_10109);
nor U17009 (N_17009,N_11238,N_12038);
nand U17010 (N_17010,N_11427,N_11158);
nor U17011 (N_17011,N_12887,N_13923);
nor U17012 (N_17012,N_12277,N_14816);
nor U17013 (N_17013,N_13204,N_13111);
nand U17014 (N_17014,N_14603,N_14517);
nor U17015 (N_17015,N_12685,N_14867);
or U17016 (N_17016,N_14613,N_11488);
and U17017 (N_17017,N_12199,N_13185);
nand U17018 (N_17018,N_13550,N_12033);
nor U17019 (N_17019,N_14267,N_13159);
nor U17020 (N_17020,N_14486,N_14671);
and U17021 (N_17021,N_14164,N_10102);
nor U17022 (N_17022,N_11793,N_10533);
and U17023 (N_17023,N_14682,N_13431);
or U17024 (N_17024,N_11697,N_10997);
nor U17025 (N_17025,N_14027,N_10309);
nand U17026 (N_17026,N_11081,N_13783);
and U17027 (N_17027,N_13619,N_14092);
nor U17028 (N_17028,N_13580,N_10799);
or U17029 (N_17029,N_11691,N_14698);
or U17030 (N_17030,N_12602,N_13553);
nand U17031 (N_17031,N_13507,N_11382);
nand U17032 (N_17032,N_14898,N_13226);
nand U17033 (N_17033,N_12867,N_14604);
or U17034 (N_17034,N_13013,N_11233);
nand U17035 (N_17035,N_10274,N_11820);
or U17036 (N_17036,N_13048,N_13689);
nand U17037 (N_17037,N_12905,N_12183);
and U17038 (N_17038,N_10145,N_11639);
nor U17039 (N_17039,N_11074,N_13963);
xnor U17040 (N_17040,N_10415,N_11308);
or U17041 (N_17041,N_12092,N_13325);
nand U17042 (N_17042,N_13503,N_10658);
or U17043 (N_17043,N_14003,N_14558);
and U17044 (N_17044,N_14670,N_10855);
nand U17045 (N_17045,N_14343,N_14500);
or U17046 (N_17046,N_13295,N_12551);
nor U17047 (N_17047,N_12000,N_11057);
nor U17048 (N_17048,N_14166,N_11992);
or U17049 (N_17049,N_14042,N_11452);
or U17050 (N_17050,N_14706,N_14439);
or U17051 (N_17051,N_14160,N_12064);
and U17052 (N_17052,N_13863,N_14188);
or U17053 (N_17053,N_14766,N_11925);
or U17054 (N_17054,N_11111,N_12543);
nand U17055 (N_17055,N_12222,N_12724);
nor U17056 (N_17056,N_14968,N_11718);
nand U17057 (N_17057,N_14578,N_14346);
and U17058 (N_17058,N_14579,N_13721);
nand U17059 (N_17059,N_12298,N_10067);
nor U17060 (N_17060,N_13751,N_10913);
and U17061 (N_17061,N_14619,N_10669);
or U17062 (N_17062,N_14167,N_11315);
nor U17063 (N_17063,N_10045,N_12670);
and U17064 (N_17064,N_12823,N_12334);
nand U17065 (N_17065,N_14452,N_11030);
nor U17066 (N_17066,N_11504,N_10530);
or U17067 (N_17067,N_14333,N_11828);
and U17068 (N_17068,N_14824,N_14916);
nor U17069 (N_17069,N_13626,N_11193);
and U17070 (N_17070,N_11109,N_10105);
nor U17071 (N_17071,N_14387,N_12819);
xnor U17072 (N_17072,N_13962,N_13369);
xor U17073 (N_17073,N_14293,N_12925);
nor U17074 (N_17074,N_13321,N_10025);
nand U17075 (N_17075,N_11279,N_11071);
and U17076 (N_17076,N_11829,N_13207);
and U17077 (N_17077,N_11425,N_12150);
or U17078 (N_17078,N_13594,N_12672);
nand U17079 (N_17079,N_14418,N_13208);
nand U17080 (N_17080,N_13054,N_12219);
and U17081 (N_17081,N_14845,N_10289);
or U17082 (N_17082,N_13138,N_10139);
nor U17083 (N_17083,N_14424,N_12860);
nor U17084 (N_17084,N_10713,N_10037);
nand U17085 (N_17085,N_13688,N_12323);
and U17086 (N_17086,N_12519,N_11750);
nand U17087 (N_17087,N_12143,N_13370);
and U17088 (N_17088,N_13687,N_13123);
or U17089 (N_17089,N_11200,N_10268);
nand U17090 (N_17090,N_12171,N_11347);
and U17091 (N_17091,N_10088,N_13434);
and U17092 (N_17092,N_10838,N_13167);
and U17093 (N_17093,N_14987,N_11317);
and U17094 (N_17094,N_12718,N_14327);
nand U17095 (N_17095,N_13210,N_13133);
nand U17096 (N_17096,N_11210,N_12872);
or U17097 (N_17097,N_10061,N_12134);
or U17098 (N_17098,N_13456,N_13388);
nand U17099 (N_17099,N_14702,N_12770);
nor U17100 (N_17100,N_14961,N_13613);
nor U17101 (N_17101,N_14129,N_14025);
nand U17102 (N_17102,N_14843,N_14664);
and U17103 (N_17103,N_11574,N_14467);
and U17104 (N_17104,N_10395,N_12418);
or U17105 (N_17105,N_11804,N_12464);
and U17106 (N_17106,N_12700,N_10741);
or U17107 (N_17107,N_13592,N_14383);
and U17108 (N_17108,N_14313,N_12550);
or U17109 (N_17109,N_11862,N_14466);
and U17110 (N_17110,N_11377,N_11785);
and U17111 (N_17111,N_12487,N_10360);
nor U17112 (N_17112,N_11000,N_10426);
or U17113 (N_17113,N_13371,N_13041);
and U17114 (N_17114,N_11514,N_14525);
nand U17115 (N_17115,N_12437,N_13484);
and U17116 (N_17116,N_14351,N_11467);
or U17117 (N_17117,N_10718,N_14576);
and U17118 (N_17118,N_14114,N_13782);
nor U17119 (N_17119,N_11715,N_14286);
nor U17120 (N_17120,N_12266,N_10740);
nand U17121 (N_17121,N_12835,N_10661);
nor U17122 (N_17122,N_11616,N_12895);
nor U17123 (N_17123,N_12390,N_14937);
and U17124 (N_17124,N_12856,N_14268);
nor U17125 (N_17125,N_11180,N_10353);
or U17126 (N_17126,N_14475,N_11582);
nand U17127 (N_17127,N_12302,N_12056);
nand U17128 (N_17128,N_13331,N_11290);
nor U17129 (N_17129,N_14057,N_11257);
nor U17130 (N_17130,N_10961,N_14379);
nor U17131 (N_17131,N_13979,N_10747);
nor U17132 (N_17132,N_14690,N_11848);
or U17133 (N_17133,N_14221,N_13149);
and U17134 (N_17134,N_14020,N_13870);
or U17135 (N_17135,N_10352,N_13482);
or U17136 (N_17136,N_12753,N_13160);
nor U17137 (N_17137,N_12591,N_14894);
nor U17138 (N_17138,N_13096,N_12869);
and U17139 (N_17139,N_11319,N_11439);
nor U17140 (N_17140,N_13071,N_13552);
and U17141 (N_17141,N_11970,N_12576);
or U17142 (N_17142,N_14497,N_12229);
or U17143 (N_17143,N_13777,N_14408);
and U17144 (N_17144,N_10986,N_14991);
xor U17145 (N_17145,N_12446,N_11289);
nand U17146 (N_17146,N_10887,N_14884);
nand U17147 (N_17147,N_11599,N_14367);
or U17148 (N_17148,N_12267,N_11458);
or U17149 (N_17149,N_12924,N_11087);
nor U17150 (N_17150,N_11641,N_12012);
or U17151 (N_17151,N_13848,N_14290);
and U17152 (N_17152,N_12209,N_13757);
and U17153 (N_17153,N_10823,N_13555);
or U17154 (N_17154,N_14978,N_12236);
nand U17155 (N_17155,N_11575,N_10279);
nor U17156 (N_17156,N_11852,N_10792);
nand U17157 (N_17157,N_12880,N_13505);
and U17158 (N_17158,N_12231,N_13423);
nand U17159 (N_17159,N_10647,N_13682);
or U17160 (N_17160,N_11389,N_10054);
nor U17161 (N_17161,N_14131,N_14678);
and U17162 (N_17162,N_12029,N_11468);
nor U17163 (N_17163,N_11399,N_13601);
and U17164 (N_17164,N_12711,N_14378);
nor U17165 (N_17165,N_10621,N_11526);
and U17166 (N_17166,N_13219,N_12812);
and U17167 (N_17167,N_10393,N_14041);
and U17168 (N_17168,N_10431,N_11453);
nand U17169 (N_17169,N_12336,N_14049);
nand U17170 (N_17170,N_12712,N_12520);
nand U17171 (N_17171,N_12811,N_13342);
or U17172 (N_17172,N_14605,N_12773);
or U17173 (N_17173,N_10711,N_12225);
nor U17174 (N_17174,N_14615,N_11023);
nand U17175 (N_17175,N_11529,N_10160);
or U17176 (N_17176,N_10317,N_10878);
nor U17177 (N_17177,N_10423,N_10772);
and U17178 (N_17178,N_10575,N_12827);
nor U17179 (N_17179,N_12926,N_11786);
and U17180 (N_17180,N_12058,N_13841);
or U17181 (N_17181,N_10498,N_12959);
and U17182 (N_17182,N_14921,N_10328);
nand U17183 (N_17183,N_14073,N_10656);
or U17184 (N_17184,N_14863,N_10793);
or U17185 (N_17185,N_10419,N_13879);
nor U17186 (N_17186,N_11369,N_11824);
nand U17187 (N_17187,N_12218,N_13988);
or U17188 (N_17188,N_14614,N_12729);
or U17189 (N_17189,N_11818,N_14840);
or U17190 (N_17190,N_13660,N_13329);
and U17191 (N_17191,N_14431,N_13465);
nand U17192 (N_17192,N_10344,N_14405);
nand U17193 (N_17193,N_11683,N_10242);
and U17194 (N_17194,N_11166,N_10882);
nor U17195 (N_17195,N_13764,N_14345);
nand U17196 (N_17196,N_14950,N_12985);
xnor U17197 (N_17197,N_14980,N_13907);
and U17198 (N_17198,N_10818,N_14371);
nand U17199 (N_17199,N_14083,N_13430);
xnor U17200 (N_17200,N_11738,N_14285);
and U17201 (N_17201,N_10169,N_12766);
nand U17202 (N_17202,N_14848,N_11663);
and U17203 (N_17203,N_12620,N_11883);
nand U17204 (N_17204,N_11438,N_14443);
and U17205 (N_17205,N_14801,N_11964);
and U17206 (N_17206,N_13788,N_12772);
nor U17207 (N_17207,N_12320,N_11563);
xor U17208 (N_17208,N_12197,N_13809);
nor U17209 (N_17209,N_13836,N_13271);
nor U17210 (N_17210,N_13801,N_13942);
or U17211 (N_17211,N_12893,N_10751);
and U17212 (N_17212,N_12424,N_14494);
nand U17213 (N_17213,N_12675,N_13171);
and U17214 (N_17214,N_14858,N_10989);
nand U17215 (N_17215,N_14953,N_12544);
or U17216 (N_17216,N_13752,N_12207);
or U17217 (N_17217,N_10816,N_14104);
nor U17218 (N_17218,N_12290,N_10011);
nor U17219 (N_17219,N_11557,N_12818);
nor U17220 (N_17220,N_13010,N_11996);
nor U17221 (N_17221,N_12028,N_11094);
and U17222 (N_17222,N_12767,N_14686);
nor U17223 (N_17223,N_12489,N_10856);
or U17224 (N_17224,N_10221,N_11079);
xor U17225 (N_17225,N_14826,N_12613);
nand U17226 (N_17226,N_10002,N_12992);
or U17227 (N_17227,N_14421,N_12759);
nand U17228 (N_17228,N_11735,N_14646);
nor U17229 (N_17229,N_13225,N_10046);
and U17230 (N_17230,N_13880,N_13280);
nand U17231 (N_17231,N_11393,N_14461);
nor U17232 (N_17232,N_12523,N_14986);
nor U17233 (N_17233,N_11935,N_14029);
or U17234 (N_17234,N_10052,N_14746);
nor U17235 (N_17235,N_11183,N_11951);
and U17236 (N_17236,N_10010,N_11509);
nor U17237 (N_17237,N_11976,N_14291);
or U17238 (N_17238,N_14069,N_13914);
and U17239 (N_17239,N_13890,N_10283);
nand U17240 (N_17240,N_14359,N_11649);
and U17241 (N_17241,N_14844,N_10578);
and U17242 (N_17242,N_10926,N_11656);
nand U17243 (N_17243,N_12804,N_12828);
xor U17244 (N_17244,N_14455,N_13716);
nand U17245 (N_17245,N_12861,N_12526);
and U17246 (N_17246,N_13867,N_12305);
and U17247 (N_17247,N_11585,N_14654);
nand U17248 (N_17248,N_12095,N_11922);
and U17249 (N_17249,N_13309,N_12234);
nor U17250 (N_17250,N_13162,N_14873);
or U17251 (N_17251,N_12619,N_14428);
and U17252 (N_17252,N_12495,N_12907);
nor U17253 (N_17253,N_10164,N_14219);
nand U17254 (N_17254,N_11304,N_14229);
xor U17255 (N_17255,N_13558,N_11923);
and U17256 (N_17256,N_11762,N_10775);
nand U17257 (N_17257,N_11119,N_10587);
nor U17258 (N_17258,N_10576,N_13165);
nor U17259 (N_17259,N_14593,N_10481);
and U17260 (N_17260,N_12397,N_14341);
nor U17261 (N_17261,N_14681,N_14218);
nand U17262 (N_17262,N_11839,N_14088);
and U17263 (N_17263,N_12172,N_14548);
nand U17264 (N_17264,N_11444,N_11093);
or U17265 (N_17265,N_13113,N_13827);
or U17266 (N_17266,N_11043,N_11137);
nor U17267 (N_17267,N_13397,N_10681);
or U17268 (N_17268,N_10960,N_13406);
xnor U17269 (N_17269,N_10895,N_13091);
nand U17270 (N_17270,N_12055,N_11041);
nor U17271 (N_17271,N_14410,N_11813);
nor U17272 (N_17272,N_10893,N_12527);
or U17273 (N_17273,N_12493,N_12129);
nand U17274 (N_17274,N_11177,N_10296);
and U17275 (N_17275,N_12960,N_14086);
nand U17276 (N_17276,N_11897,N_12365);
nor U17277 (N_17277,N_13337,N_12663);
or U17278 (N_17278,N_11260,N_10813);
and U17279 (N_17279,N_11403,N_13415);
or U17280 (N_17280,N_11055,N_12034);
or U17281 (N_17281,N_14981,N_11227);
nand U17282 (N_17282,N_13758,N_12722);
or U17283 (N_17283,N_10735,N_10209);
or U17284 (N_17284,N_10914,N_11324);
or U17285 (N_17285,N_12378,N_13898);
nand U17286 (N_17286,N_14413,N_11550);
nor U17287 (N_17287,N_11150,N_14523);
nand U17288 (N_17288,N_13964,N_14059);
and U17289 (N_17289,N_11006,N_14949);
nand U17290 (N_17290,N_10976,N_10720);
and U17291 (N_17291,N_13986,N_14535);
or U17292 (N_17292,N_11008,N_10547);
or U17293 (N_17293,N_11665,N_12512);
and U17294 (N_17294,N_11841,N_12807);
nor U17295 (N_17295,N_10203,N_13937);
nand U17296 (N_17296,N_12285,N_12088);
nand U17297 (N_17297,N_12357,N_12472);
and U17298 (N_17298,N_13150,N_10400);
nand U17299 (N_17299,N_12361,N_13077);
and U17300 (N_17300,N_13961,N_13713);
nor U17301 (N_17301,N_13241,N_12768);
or U17302 (N_17302,N_14944,N_14113);
nor U17303 (N_17303,N_12087,N_13587);
xor U17304 (N_17304,N_13947,N_10979);
nand U17305 (N_17305,N_11040,N_11011);
and U17306 (N_17306,N_14862,N_13467);
and U17307 (N_17307,N_10857,N_10896);
or U17308 (N_17308,N_10706,N_13833);
and U17309 (N_17309,N_11431,N_14198);
and U17310 (N_17310,N_14829,N_13211);
nor U17311 (N_17311,N_13037,N_11330);
and U17312 (N_17312,N_14893,N_11419);
and U17313 (N_17313,N_13528,N_14789);
or U17314 (N_17314,N_13373,N_13504);
nor U17315 (N_17315,N_10513,N_14724);
nand U17316 (N_17316,N_14960,N_13846);
nand U17317 (N_17317,N_11722,N_11837);
nor U17318 (N_17318,N_12631,N_10077);
nor U17319 (N_17319,N_12834,N_10114);
nand U17320 (N_17320,N_12746,N_12786);
nor U17321 (N_17321,N_10064,N_10839);
nand U17322 (N_17322,N_12287,N_13120);
nand U17323 (N_17323,N_10750,N_14989);
nor U17324 (N_17324,N_11246,N_14773);
or U17325 (N_17325,N_10320,N_12393);
nand U17326 (N_17326,N_12045,N_10778);
or U17327 (N_17327,N_13806,N_14869);
or U17328 (N_17328,N_10610,N_14094);
or U17329 (N_17329,N_12249,N_13624);
or U17330 (N_17330,N_13134,N_10601);
nand U17331 (N_17331,N_12738,N_14469);
nor U17332 (N_17332,N_14725,N_13389);
or U17333 (N_17333,N_10000,N_14731);
nor U17334 (N_17334,N_10753,N_12635);
or U17335 (N_17335,N_14653,N_12561);
or U17336 (N_17336,N_10579,N_13773);
or U17337 (N_17337,N_13897,N_14429);
nor U17338 (N_17338,N_13549,N_14959);
nand U17339 (N_17339,N_12847,N_14545);
or U17340 (N_17340,N_10749,N_14222);
and U17341 (N_17341,N_10622,N_14996);
or U17342 (N_17342,N_13443,N_10330);
nand U17343 (N_17343,N_11630,N_13412);
nor U17344 (N_17344,N_11207,N_10047);
nor U17345 (N_17345,N_13637,N_12787);
or U17346 (N_17346,N_10566,N_14642);
nand U17347 (N_17347,N_13141,N_13180);
and U17348 (N_17348,N_11206,N_14704);
nor U17349 (N_17349,N_14111,N_10414);
nor U17350 (N_17350,N_10821,N_10040);
or U17351 (N_17351,N_14303,N_11323);
and U17352 (N_17352,N_12933,N_13413);
and U17353 (N_17353,N_10373,N_13178);
nand U17354 (N_17354,N_13471,N_11532);
nand U17355 (N_17355,N_12944,N_12317);
xor U17356 (N_17356,N_10523,N_13169);
and U17357 (N_17357,N_11203,N_13824);
nor U17358 (N_17358,N_10495,N_10871);
nor U17359 (N_17359,N_13915,N_10908);
nor U17360 (N_17360,N_14279,N_10861);
nor U17361 (N_17361,N_10705,N_12384);
and U17362 (N_17362,N_10777,N_14180);
xnor U17363 (N_17363,N_10609,N_10727);
and U17364 (N_17364,N_10733,N_14896);
xnor U17365 (N_17365,N_11667,N_12699);
and U17366 (N_17366,N_10520,N_12030);
nor U17367 (N_17367,N_13701,N_12276);
or U17368 (N_17368,N_11945,N_14393);
nand U17369 (N_17369,N_12244,N_11460);
nor U17370 (N_17370,N_14875,N_13152);
and U17371 (N_17371,N_13822,N_14061);
nor U17372 (N_17372,N_13139,N_12943);
or U17373 (N_17373,N_12669,N_14821);
and U17374 (N_17374,N_11795,N_11046);
or U17375 (N_17375,N_10351,N_12376);
and U17376 (N_17376,N_11763,N_10641);
and U17377 (N_17377,N_14582,N_13461);
nand U17378 (N_17378,N_10607,N_14471);
nand U17379 (N_17379,N_11205,N_10541);
or U17380 (N_17380,N_11076,N_11356);
nor U17381 (N_17381,N_12478,N_13572);
nor U17382 (N_17382,N_12703,N_13199);
or U17383 (N_17383,N_10814,N_12793);
or U17384 (N_17384,N_12496,N_13968);
or U17385 (N_17385,N_14213,N_12068);
or U17386 (N_17386,N_11120,N_12918);
nor U17387 (N_17387,N_14633,N_12780);
or U17388 (N_17388,N_11146,N_10206);
nor U17389 (N_17389,N_13547,N_10525);
nor U17390 (N_17390,N_10657,N_14457);
and U17391 (N_17391,N_14998,N_13368);
or U17392 (N_17392,N_11341,N_12691);
nand U17393 (N_17393,N_13921,N_10284);
nand U17394 (N_17394,N_12096,N_10817);
nand U17395 (N_17395,N_14417,N_10112);
nand U17396 (N_17396,N_10251,N_13216);
or U17397 (N_17397,N_13928,N_10291);
and U17398 (N_17398,N_13602,N_11381);
nor U17399 (N_17399,N_10062,N_11907);
nor U17400 (N_17400,N_14866,N_10076);
xnor U17401 (N_17401,N_14734,N_14637);
and U17402 (N_17402,N_11647,N_12578);
nand U17403 (N_17403,N_12442,N_11890);
nor U17404 (N_17404,N_14765,N_11963);
and U17405 (N_17405,N_12548,N_12833);
and U17406 (N_17406,N_11676,N_11746);
nor U17407 (N_17407,N_12581,N_12474);
or U17408 (N_17408,N_12973,N_10549);
nor U17409 (N_17409,N_10398,N_13062);
and U17410 (N_17410,N_12892,N_14060);
or U17411 (N_17411,N_11629,N_13512);
nor U17412 (N_17412,N_11826,N_11517);
or U17413 (N_17413,N_12873,N_11154);
nor U17414 (N_17414,N_14100,N_10632);
and U17415 (N_17415,N_12949,N_12228);
or U17416 (N_17416,N_14144,N_14495);
and U17417 (N_17417,N_12374,N_11939);
nor U17418 (N_17418,N_13627,N_10963);
or U17419 (N_17419,N_13399,N_14116);
or U17420 (N_17420,N_14360,N_10371);
and U17421 (N_17421,N_13270,N_13629);
nor U17422 (N_17422,N_10544,N_10087);
nor U17423 (N_17423,N_14623,N_14881);
nand U17424 (N_17424,N_13582,N_12637);
nand U17425 (N_17425,N_12383,N_12655);
and U17426 (N_17426,N_10644,N_11640);
and U17427 (N_17427,N_14158,N_10439);
and U17428 (N_17428,N_11749,N_11889);
nor U17429 (N_17429,N_12555,N_11605);
nand U17430 (N_17430,N_12443,N_10594);
nor U17431 (N_17431,N_11185,N_10930);
and U17432 (N_17432,N_14606,N_13220);
nor U17433 (N_17433,N_11773,N_11827);
or U17434 (N_17434,N_13774,N_13172);
and U17435 (N_17435,N_14750,N_12865);
and U17436 (N_17436,N_14013,N_12042);
nand U17437 (N_17437,N_12261,N_11010);
or U17438 (N_17438,N_12554,N_12479);
or U17439 (N_17439,N_13297,N_14257);
nor U17440 (N_17440,N_11390,N_10175);
nor U17441 (N_17441,N_14814,N_13952);
and U17442 (N_17442,N_11147,N_12111);
nand U17443 (N_17443,N_11644,N_13173);
and U17444 (N_17444,N_13135,N_12932);
or U17445 (N_17445,N_13686,N_12106);
nor U17446 (N_17446,N_12814,N_10688);
or U17447 (N_17447,N_11397,N_10591);
or U17448 (N_17448,N_11424,N_13290);
xor U17449 (N_17449,N_13740,N_12606);
nor U17450 (N_17450,N_10946,N_12449);
and U17451 (N_17451,N_14103,N_14391);
nor U17452 (N_17452,N_14628,N_14437);
nand U17453 (N_17453,N_14078,N_14316);
or U17454 (N_17454,N_10526,N_14338);
and U17455 (N_17455,N_11472,N_13084);
nor U17456 (N_17456,N_14031,N_10412);
nor U17457 (N_17457,N_14919,N_11265);
nor U17458 (N_17458,N_14039,N_13944);
or U17459 (N_17459,N_12406,N_13856);
nand U17460 (N_17460,N_12041,N_10548);
nor U17461 (N_17461,N_10680,N_12328);
nand U17462 (N_17462,N_13894,N_12432);
or U17463 (N_17463,N_10347,N_10234);
nor U17464 (N_17464,N_12063,N_10122);
nand U17465 (N_17465,N_14259,N_12379);
xor U17466 (N_17466,N_10442,N_10671);
and U17467 (N_17467,N_12676,N_14586);
or U17468 (N_17468,N_11371,N_10386);
nand U17469 (N_17469,N_13994,N_12599);
or U17470 (N_17470,N_14325,N_14852);
nand U17471 (N_17471,N_10467,N_12006);
and U17472 (N_17472,N_12643,N_10183);
nand U17473 (N_17473,N_12595,N_13387);
nor U17474 (N_17474,N_13006,N_14808);
or U17475 (N_17475,N_12200,N_13696);
nor U17476 (N_17476,N_13061,N_12573);
nor U17477 (N_17477,N_13499,N_12506);
and U17478 (N_17478,N_10515,N_14806);
nand U17479 (N_17479,N_11122,N_13351);
and U17480 (N_17480,N_12227,N_11871);
nand U17481 (N_17481,N_10810,N_11974);
nand U17482 (N_17482,N_10555,N_12953);
nor U17483 (N_17483,N_13228,N_10471);
nor U17484 (N_17484,N_10394,N_10397);
or U17485 (N_17485,N_12596,N_12832);
and U17486 (N_17486,N_11874,N_11921);
xor U17487 (N_17487,N_14913,N_12922);
or U17488 (N_17488,N_10233,N_13611);
nor U17489 (N_17489,N_13720,N_12017);
nand U17490 (N_17490,N_14054,N_14470);
nand U17491 (N_17491,N_12621,N_12308);
nor U17492 (N_17492,N_11104,N_14238);
or U17493 (N_17493,N_10012,N_11814);
nor U17494 (N_17494,N_12721,N_11048);
and U17495 (N_17495,N_14444,N_12104);
nand U17496 (N_17496,N_12598,N_11394);
nor U17497 (N_17497,N_12071,N_10275);
nor U17498 (N_17498,N_12821,N_10731);
nand U17499 (N_17499,N_10191,N_13768);
xnor U17500 (N_17500,N_12730,N_11403);
nand U17501 (N_17501,N_10312,N_12587);
or U17502 (N_17502,N_11728,N_11669);
nand U17503 (N_17503,N_13721,N_11611);
and U17504 (N_17504,N_10686,N_14112);
or U17505 (N_17505,N_10245,N_11161);
nand U17506 (N_17506,N_14433,N_13415);
nor U17507 (N_17507,N_11508,N_10212);
and U17508 (N_17508,N_12327,N_14005);
or U17509 (N_17509,N_10852,N_13746);
nand U17510 (N_17510,N_11060,N_11629);
or U17511 (N_17511,N_13046,N_13809);
nand U17512 (N_17512,N_14992,N_10333);
and U17513 (N_17513,N_11077,N_13155);
and U17514 (N_17514,N_13818,N_14062);
and U17515 (N_17515,N_11181,N_11915);
nor U17516 (N_17516,N_10467,N_12729);
nor U17517 (N_17517,N_14341,N_14939);
nor U17518 (N_17518,N_14532,N_12812);
nand U17519 (N_17519,N_12894,N_10458);
and U17520 (N_17520,N_11126,N_13397);
and U17521 (N_17521,N_12641,N_10362);
nand U17522 (N_17522,N_12778,N_10415);
or U17523 (N_17523,N_12244,N_11149);
and U17524 (N_17524,N_10112,N_12540);
and U17525 (N_17525,N_11206,N_13348);
nor U17526 (N_17526,N_12347,N_14465);
and U17527 (N_17527,N_14919,N_13272);
and U17528 (N_17528,N_11959,N_14425);
nor U17529 (N_17529,N_14960,N_13718);
nand U17530 (N_17530,N_11889,N_13390);
nand U17531 (N_17531,N_11677,N_10752);
and U17532 (N_17532,N_11735,N_14144);
or U17533 (N_17533,N_12252,N_14132);
nor U17534 (N_17534,N_10918,N_11588);
nor U17535 (N_17535,N_11366,N_12266);
xnor U17536 (N_17536,N_10337,N_12592);
and U17537 (N_17537,N_11364,N_14325);
and U17538 (N_17538,N_11718,N_12297);
and U17539 (N_17539,N_14982,N_10558);
and U17540 (N_17540,N_10256,N_14879);
xor U17541 (N_17541,N_10188,N_14581);
and U17542 (N_17542,N_10853,N_13783);
nand U17543 (N_17543,N_11798,N_11667);
or U17544 (N_17544,N_11024,N_11266);
nor U17545 (N_17545,N_12248,N_14711);
nor U17546 (N_17546,N_12551,N_11551);
and U17547 (N_17547,N_11733,N_14253);
or U17548 (N_17548,N_14926,N_12519);
or U17549 (N_17549,N_11171,N_10658);
and U17550 (N_17550,N_11056,N_12984);
xnor U17551 (N_17551,N_13701,N_10972);
nand U17552 (N_17552,N_12129,N_12321);
and U17553 (N_17553,N_13539,N_13168);
nor U17554 (N_17554,N_13897,N_11401);
and U17555 (N_17555,N_14487,N_14236);
nand U17556 (N_17556,N_14311,N_12719);
or U17557 (N_17557,N_10844,N_10963);
nor U17558 (N_17558,N_14296,N_13393);
nand U17559 (N_17559,N_10747,N_14366);
nand U17560 (N_17560,N_10494,N_11275);
or U17561 (N_17561,N_11244,N_14708);
and U17562 (N_17562,N_14656,N_14317);
nand U17563 (N_17563,N_14408,N_14447);
nand U17564 (N_17564,N_13791,N_10202);
or U17565 (N_17565,N_12895,N_12163);
nor U17566 (N_17566,N_13652,N_14113);
or U17567 (N_17567,N_14920,N_14095);
and U17568 (N_17568,N_12729,N_14057);
and U17569 (N_17569,N_10246,N_14035);
or U17570 (N_17570,N_14229,N_10434);
or U17571 (N_17571,N_13953,N_10782);
or U17572 (N_17572,N_12312,N_14764);
or U17573 (N_17573,N_10455,N_13112);
and U17574 (N_17574,N_12026,N_12524);
nor U17575 (N_17575,N_13671,N_13378);
nand U17576 (N_17576,N_10609,N_11692);
or U17577 (N_17577,N_14083,N_11389);
and U17578 (N_17578,N_11045,N_13565);
nor U17579 (N_17579,N_12226,N_12608);
and U17580 (N_17580,N_10532,N_13035);
and U17581 (N_17581,N_12018,N_14430);
or U17582 (N_17582,N_12205,N_11532);
or U17583 (N_17583,N_10512,N_12310);
or U17584 (N_17584,N_13759,N_12791);
nor U17585 (N_17585,N_10936,N_12500);
or U17586 (N_17586,N_11903,N_14155);
nand U17587 (N_17587,N_14800,N_11308);
and U17588 (N_17588,N_11035,N_12282);
or U17589 (N_17589,N_14837,N_13394);
or U17590 (N_17590,N_13540,N_12045);
and U17591 (N_17591,N_10732,N_12727);
or U17592 (N_17592,N_12244,N_12263);
or U17593 (N_17593,N_10193,N_14390);
or U17594 (N_17594,N_14154,N_10488);
and U17595 (N_17595,N_10522,N_13406);
or U17596 (N_17596,N_10086,N_13092);
xnor U17597 (N_17597,N_12058,N_10753);
nor U17598 (N_17598,N_13281,N_12673);
xnor U17599 (N_17599,N_13228,N_10776);
nand U17600 (N_17600,N_12793,N_12774);
or U17601 (N_17601,N_10913,N_10480);
nand U17602 (N_17602,N_12906,N_11860);
nor U17603 (N_17603,N_12539,N_11363);
nor U17604 (N_17604,N_13495,N_10930);
or U17605 (N_17605,N_13685,N_12398);
nand U17606 (N_17606,N_14085,N_12854);
nand U17607 (N_17607,N_14845,N_11151);
and U17608 (N_17608,N_14205,N_12750);
nand U17609 (N_17609,N_13990,N_12192);
or U17610 (N_17610,N_12324,N_11756);
or U17611 (N_17611,N_11639,N_13384);
and U17612 (N_17612,N_13051,N_12414);
and U17613 (N_17613,N_11243,N_12147);
or U17614 (N_17614,N_10639,N_14601);
nor U17615 (N_17615,N_13234,N_13579);
nand U17616 (N_17616,N_12316,N_10142);
or U17617 (N_17617,N_13920,N_11673);
and U17618 (N_17618,N_13997,N_10685);
nand U17619 (N_17619,N_13971,N_14619);
or U17620 (N_17620,N_13312,N_11279);
or U17621 (N_17621,N_13861,N_12718);
and U17622 (N_17622,N_13776,N_10489);
nor U17623 (N_17623,N_14741,N_11436);
nor U17624 (N_17624,N_14409,N_12760);
or U17625 (N_17625,N_10937,N_14058);
and U17626 (N_17626,N_13261,N_13410);
nand U17627 (N_17627,N_11129,N_10737);
nand U17628 (N_17628,N_10077,N_14242);
nand U17629 (N_17629,N_14254,N_12911);
nor U17630 (N_17630,N_14309,N_13021);
nand U17631 (N_17631,N_11354,N_10861);
nor U17632 (N_17632,N_13928,N_10634);
nand U17633 (N_17633,N_10074,N_14407);
or U17634 (N_17634,N_14997,N_11704);
nor U17635 (N_17635,N_14444,N_12358);
nor U17636 (N_17636,N_13317,N_11135);
or U17637 (N_17637,N_11339,N_14758);
nand U17638 (N_17638,N_14789,N_14295);
or U17639 (N_17639,N_11427,N_14048);
nor U17640 (N_17640,N_13487,N_13758);
and U17641 (N_17641,N_13464,N_10429);
or U17642 (N_17642,N_13131,N_13241);
or U17643 (N_17643,N_11706,N_14002);
nand U17644 (N_17644,N_14275,N_10177);
or U17645 (N_17645,N_11591,N_14910);
nor U17646 (N_17646,N_11254,N_12433);
and U17647 (N_17647,N_13287,N_11669);
and U17648 (N_17648,N_13448,N_11259);
nand U17649 (N_17649,N_13064,N_14616);
nor U17650 (N_17650,N_13098,N_10562);
and U17651 (N_17651,N_13385,N_11297);
nor U17652 (N_17652,N_10080,N_14869);
or U17653 (N_17653,N_14539,N_12110);
and U17654 (N_17654,N_13728,N_14071);
and U17655 (N_17655,N_12594,N_10774);
and U17656 (N_17656,N_11638,N_14243);
and U17657 (N_17657,N_13482,N_10323);
or U17658 (N_17658,N_11686,N_13324);
nor U17659 (N_17659,N_10170,N_10729);
nand U17660 (N_17660,N_10911,N_13362);
or U17661 (N_17661,N_10400,N_11469);
and U17662 (N_17662,N_12073,N_13487);
and U17663 (N_17663,N_11201,N_10400);
nor U17664 (N_17664,N_13823,N_11368);
and U17665 (N_17665,N_12565,N_10717);
nand U17666 (N_17666,N_14944,N_13590);
and U17667 (N_17667,N_13818,N_13925);
or U17668 (N_17668,N_12065,N_14542);
or U17669 (N_17669,N_10217,N_14182);
and U17670 (N_17670,N_10703,N_12893);
nor U17671 (N_17671,N_10206,N_13992);
and U17672 (N_17672,N_11663,N_13006);
and U17673 (N_17673,N_11276,N_14864);
or U17674 (N_17674,N_12107,N_11422);
or U17675 (N_17675,N_10204,N_10430);
or U17676 (N_17676,N_11048,N_10561);
nor U17677 (N_17677,N_10408,N_11648);
nor U17678 (N_17678,N_12318,N_12019);
or U17679 (N_17679,N_10451,N_14656);
nor U17680 (N_17680,N_14260,N_13545);
nand U17681 (N_17681,N_12522,N_13229);
nor U17682 (N_17682,N_10031,N_13626);
nor U17683 (N_17683,N_11857,N_11395);
nor U17684 (N_17684,N_12283,N_11284);
nor U17685 (N_17685,N_13656,N_14061);
or U17686 (N_17686,N_12360,N_10154);
nor U17687 (N_17687,N_13639,N_12492);
and U17688 (N_17688,N_14295,N_10408);
nand U17689 (N_17689,N_12748,N_13648);
or U17690 (N_17690,N_11238,N_14597);
nand U17691 (N_17691,N_14239,N_11616);
or U17692 (N_17692,N_13470,N_12587);
xor U17693 (N_17693,N_12399,N_14030);
and U17694 (N_17694,N_10273,N_10711);
and U17695 (N_17695,N_14344,N_10221);
nor U17696 (N_17696,N_10536,N_12475);
or U17697 (N_17697,N_14669,N_13551);
and U17698 (N_17698,N_12468,N_11945);
nor U17699 (N_17699,N_10592,N_12161);
or U17700 (N_17700,N_10850,N_12285);
nand U17701 (N_17701,N_11095,N_11858);
or U17702 (N_17702,N_14681,N_11687);
and U17703 (N_17703,N_13872,N_12305);
nor U17704 (N_17704,N_13983,N_14966);
nand U17705 (N_17705,N_10360,N_12131);
nand U17706 (N_17706,N_10033,N_11850);
and U17707 (N_17707,N_12165,N_11484);
or U17708 (N_17708,N_12160,N_13953);
nand U17709 (N_17709,N_11575,N_13145);
nand U17710 (N_17710,N_10586,N_14730);
and U17711 (N_17711,N_14042,N_13663);
and U17712 (N_17712,N_14606,N_13962);
nand U17713 (N_17713,N_11395,N_10996);
nor U17714 (N_17714,N_14901,N_13054);
or U17715 (N_17715,N_12654,N_13039);
nand U17716 (N_17716,N_11670,N_12485);
or U17717 (N_17717,N_10724,N_12148);
nand U17718 (N_17718,N_11082,N_10689);
or U17719 (N_17719,N_12162,N_12948);
nand U17720 (N_17720,N_11805,N_12357);
or U17721 (N_17721,N_12631,N_14564);
nand U17722 (N_17722,N_10237,N_11216);
nor U17723 (N_17723,N_13221,N_14672);
or U17724 (N_17724,N_12753,N_11988);
nand U17725 (N_17725,N_10187,N_11823);
or U17726 (N_17726,N_12620,N_10857);
nor U17727 (N_17727,N_13041,N_11047);
and U17728 (N_17728,N_14814,N_13349);
and U17729 (N_17729,N_10967,N_10229);
and U17730 (N_17730,N_14441,N_14610);
nor U17731 (N_17731,N_12035,N_13772);
and U17732 (N_17732,N_11724,N_12833);
nand U17733 (N_17733,N_14700,N_10669);
and U17734 (N_17734,N_11786,N_12726);
nand U17735 (N_17735,N_12356,N_14997);
nand U17736 (N_17736,N_12571,N_14660);
and U17737 (N_17737,N_10632,N_13147);
nor U17738 (N_17738,N_13636,N_13419);
nand U17739 (N_17739,N_11000,N_11387);
nand U17740 (N_17740,N_10172,N_13856);
and U17741 (N_17741,N_14555,N_14046);
or U17742 (N_17742,N_14701,N_13725);
or U17743 (N_17743,N_10307,N_12805);
nor U17744 (N_17744,N_10419,N_13612);
or U17745 (N_17745,N_12049,N_13179);
and U17746 (N_17746,N_11909,N_12374);
xnor U17747 (N_17747,N_13439,N_11110);
and U17748 (N_17748,N_11134,N_14023);
nor U17749 (N_17749,N_10514,N_10759);
nand U17750 (N_17750,N_12255,N_14463);
nor U17751 (N_17751,N_11020,N_10446);
nand U17752 (N_17752,N_14510,N_10975);
nand U17753 (N_17753,N_12620,N_13097);
nand U17754 (N_17754,N_14165,N_14310);
nor U17755 (N_17755,N_12725,N_10197);
or U17756 (N_17756,N_13057,N_14528);
or U17757 (N_17757,N_13755,N_10786);
nand U17758 (N_17758,N_14890,N_13754);
nor U17759 (N_17759,N_12933,N_11912);
or U17760 (N_17760,N_10786,N_10305);
nand U17761 (N_17761,N_10876,N_14125);
xnor U17762 (N_17762,N_11356,N_12823);
nor U17763 (N_17763,N_12702,N_12218);
nor U17764 (N_17764,N_12771,N_12734);
and U17765 (N_17765,N_13298,N_13863);
or U17766 (N_17766,N_13478,N_12411);
nor U17767 (N_17767,N_13440,N_11710);
nand U17768 (N_17768,N_14312,N_14548);
nor U17769 (N_17769,N_13564,N_10807);
and U17770 (N_17770,N_10412,N_10266);
nand U17771 (N_17771,N_12664,N_11529);
or U17772 (N_17772,N_12532,N_11888);
or U17773 (N_17773,N_11743,N_14055);
nor U17774 (N_17774,N_12360,N_13836);
and U17775 (N_17775,N_11755,N_10186);
and U17776 (N_17776,N_10705,N_11241);
xor U17777 (N_17777,N_12064,N_12659);
or U17778 (N_17778,N_10979,N_12396);
xor U17779 (N_17779,N_10737,N_12870);
nand U17780 (N_17780,N_12649,N_14724);
nand U17781 (N_17781,N_13546,N_14516);
and U17782 (N_17782,N_14165,N_12217);
or U17783 (N_17783,N_10348,N_10582);
and U17784 (N_17784,N_12613,N_13930);
nor U17785 (N_17785,N_13361,N_11374);
nor U17786 (N_17786,N_12794,N_10071);
nor U17787 (N_17787,N_10924,N_14033);
and U17788 (N_17788,N_14619,N_14572);
or U17789 (N_17789,N_13245,N_13348);
nor U17790 (N_17790,N_12779,N_10134);
nor U17791 (N_17791,N_14915,N_12331);
and U17792 (N_17792,N_14892,N_11284);
nand U17793 (N_17793,N_14074,N_14946);
and U17794 (N_17794,N_14103,N_13539);
or U17795 (N_17795,N_14996,N_14795);
nand U17796 (N_17796,N_14646,N_13925);
nand U17797 (N_17797,N_11651,N_11911);
nor U17798 (N_17798,N_13976,N_14043);
or U17799 (N_17799,N_13310,N_13018);
or U17800 (N_17800,N_13824,N_10326);
nand U17801 (N_17801,N_13716,N_10406);
nand U17802 (N_17802,N_11866,N_12504);
nand U17803 (N_17803,N_14754,N_14677);
nor U17804 (N_17804,N_11482,N_12139);
nor U17805 (N_17805,N_12620,N_11828);
and U17806 (N_17806,N_10719,N_13573);
nor U17807 (N_17807,N_14226,N_11433);
and U17808 (N_17808,N_12915,N_14396);
and U17809 (N_17809,N_14836,N_12819);
or U17810 (N_17810,N_11402,N_14334);
nand U17811 (N_17811,N_14807,N_13254);
nor U17812 (N_17812,N_14619,N_13544);
nor U17813 (N_17813,N_10913,N_11957);
or U17814 (N_17814,N_10322,N_11391);
nand U17815 (N_17815,N_10416,N_11858);
and U17816 (N_17816,N_10385,N_14684);
and U17817 (N_17817,N_12737,N_13258);
or U17818 (N_17818,N_11222,N_11350);
nor U17819 (N_17819,N_11155,N_13610);
or U17820 (N_17820,N_13367,N_11661);
nor U17821 (N_17821,N_10858,N_11917);
or U17822 (N_17822,N_10161,N_11941);
and U17823 (N_17823,N_11305,N_13038);
or U17824 (N_17824,N_11581,N_12713);
nand U17825 (N_17825,N_12721,N_11292);
nor U17826 (N_17826,N_14276,N_12527);
and U17827 (N_17827,N_10574,N_11496);
and U17828 (N_17828,N_14540,N_12692);
nand U17829 (N_17829,N_11555,N_11421);
xor U17830 (N_17830,N_13729,N_12054);
and U17831 (N_17831,N_10854,N_13393);
nor U17832 (N_17832,N_12461,N_11706);
nand U17833 (N_17833,N_14651,N_12118);
or U17834 (N_17834,N_11180,N_13146);
nand U17835 (N_17835,N_14218,N_12958);
nor U17836 (N_17836,N_10569,N_12348);
and U17837 (N_17837,N_11388,N_13580);
nor U17838 (N_17838,N_13395,N_14408);
and U17839 (N_17839,N_12262,N_13192);
nand U17840 (N_17840,N_12681,N_13421);
nor U17841 (N_17841,N_10256,N_12317);
or U17842 (N_17842,N_12788,N_10568);
nor U17843 (N_17843,N_10467,N_13853);
or U17844 (N_17844,N_10425,N_14166);
or U17845 (N_17845,N_10415,N_11750);
and U17846 (N_17846,N_12897,N_14941);
or U17847 (N_17847,N_11433,N_14775);
nor U17848 (N_17848,N_14178,N_11834);
nor U17849 (N_17849,N_10076,N_12212);
xor U17850 (N_17850,N_10669,N_11770);
nand U17851 (N_17851,N_11365,N_14849);
or U17852 (N_17852,N_14602,N_12884);
xnor U17853 (N_17853,N_12744,N_13533);
nand U17854 (N_17854,N_13864,N_14192);
nor U17855 (N_17855,N_10305,N_10196);
nor U17856 (N_17856,N_14175,N_13851);
or U17857 (N_17857,N_14899,N_12856);
and U17858 (N_17858,N_13437,N_11955);
nand U17859 (N_17859,N_14092,N_14194);
or U17860 (N_17860,N_14220,N_11589);
nor U17861 (N_17861,N_13091,N_14231);
nor U17862 (N_17862,N_11058,N_14676);
or U17863 (N_17863,N_13237,N_11415);
or U17864 (N_17864,N_13857,N_13620);
nor U17865 (N_17865,N_11835,N_12586);
nor U17866 (N_17866,N_11296,N_10448);
and U17867 (N_17867,N_12428,N_10841);
nand U17868 (N_17868,N_10248,N_10864);
and U17869 (N_17869,N_12697,N_10498);
nor U17870 (N_17870,N_11518,N_10441);
nor U17871 (N_17871,N_13916,N_13446);
and U17872 (N_17872,N_14645,N_11045);
nor U17873 (N_17873,N_11616,N_12996);
xnor U17874 (N_17874,N_14603,N_14826);
nor U17875 (N_17875,N_10999,N_14386);
nor U17876 (N_17876,N_11831,N_10622);
and U17877 (N_17877,N_10934,N_14145);
nor U17878 (N_17878,N_10230,N_12433);
nor U17879 (N_17879,N_10238,N_13313);
or U17880 (N_17880,N_12280,N_10396);
or U17881 (N_17881,N_10958,N_14925);
nor U17882 (N_17882,N_10816,N_14249);
nor U17883 (N_17883,N_11083,N_13042);
and U17884 (N_17884,N_10866,N_13753);
nor U17885 (N_17885,N_10378,N_10212);
nand U17886 (N_17886,N_10747,N_10413);
nand U17887 (N_17887,N_12816,N_12179);
and U17888 (N_17888,N_11897,N_12665);
nor U17889 (N_17889,N_13207,N_14176);
and U17890 (N_17890,N_14476,N_10445);
or U17891 (N_17891,N_13819,N_13138);
nor U17892 (N_17892,N_11666,N_11297);
nand U17893 (N_17893,N_11331,N_14324);
xnor U17894 (N_17894,N_13741,N_12015);
and U17895 (N_17895,N_10470,N_13070);
or U17896 (N_17896,N_12620,N_10955);
nand U17897 (N_17897,N_12212,N_13877);
nand U17898 (N_17898,N_12410,N_12661);
and U17899 (N_17899,N_11915,N_14165);
or U17900 (N_17900,N_10852,N_12924);
and U17901 (N_17901,N_13195,N_13466);
nand U17902 (N_17902,N_14329,N_10904);
nand U17903 (N_17903,N_14172,N_12748);
and U17904 (N_17904,N_13242,N_14856);
nor U17905 (N_17905,N_13974,N_10363);
or U17906 (N_17906,N_14749,N_10507);
nor U17907 (N_17907,N_14871,N_13844);
nand U17908 (N_17908,N_10365,N_13665);
and U17909 (N_17909,N_10632,N_12150);
nor U17910 (N_17910,N_14309,N_13251);
nor U17911 (N_17911,N_14895,N_12256);
nor U17912 (N_17912,N_14248,N_13923);
nor U17913 (N_17913,N_13293,N_10316);
nor U17914 (N_17914,N_10748,N_11298);
nand U17915 (N_17915,N_10996,N_11968);
nor U17916 (N_17916,N_13729,N_11430);
nor U17917 (N_17917,N_12947,N_13175);
and U17918 (N_17918,N_11888,N_13441);
nand U17919 (N_17919,N_14447,N_11236);
or U17920 (N_17920,N_10042,N_11583);
nor U17921 (N_17921,N_14288,N_14537);
nand U17922 (N_17922,N_14454,N_13798);
nand U17923 (N_17923,N_11781,N_14500);
nand U17924 (N_17924,N_14199,N_11226);
or U17925 (N_17925,N_13296,N_14999);
nand U17926 (N_17926,N_13763,N_13474);
or U17927 (N_17927,N_12401,N_11443);
or U17928 (N_17928,N_10296,N_14937);
nor U17929 (N_17929,N_14399,N_12055);
nor U17930 (N_17930,N_10510,N_12819);
and U17931 (N_17931,N_10635,N_10136);
nor U17932 (N_17932,N_14597,N_13468);
nor U17933 (N_17933,N_10415,N_13431);
nor U17934 (N_17934,N_14642,N_13919);
nand U17935 (N_17935,N_14301,N_13119);
or U17936 (N_17936,N_10088,N_11239);
or U17937 (N_17937,N_10454,N_11730);
or U17938 (N_17938,N_10622,N_13248);
or U17939 (N_17939,N_14457,N_12804);
xnor U17940 (N_17940,N_10776,N_13684);
nand U17941 (N_17941,N_11124,N_10975);
nand U17942 (N_17942,N_12084,N_11898);
nand U17943 (N_17943,N_12876,N_14484);
nand U17944 (N_17944,N_11779,N_10731);
and U17945 (N_17945,N_11742,N_10904);
xnor U17946 (N_17946,N_14688,N_10172);
or U17947 (N_17947,N_12897,N_14639);
nor U17948 (N_17948,N_14114,N_12245);
and U17949 (N_17949,N_13171,N_14183);
nor U17950 (N_17950,N_13936,N_13983);
and U17951 (N_17951,N_13470,N_11366);
nand U17952 (N_17952,N_11579,N_11483);
nand U17953 (N_17953,N_13974,N_13883);
nand U17954 (N_17954,N_10485,N_10680);
or U17955 (N_17955,N_10368,N_11094);
and U17956 (N_17956,N_10533,N_14634);
and U17957 (N_17957,N_13527,N_13358);
and U17958 (N_17958,N_11645,N_13151);
nand U17959 (N_17959,N_12297,N_11699);
and U17960 (N_17960,N_14160,N_14084);
or U17961 (N_17961,N_10406,N_14094);
or U17962 (N_17962,N_10906,N_12514);
or U17963 (N_17963,N_10861,N_14982);
nand U17964 (N_17964,N_11445,N_11218);
nor U17965 (N_17965,N_14306,N_11639);
or U17966 (N_17966,N_14489,N_10835);
and U17967 (N_17967,N_12301,N_13841);
and U17968 (N_17968,N_13370,N_14942);
or U17969 (N_17969,N_12106,N_10556);
or U17970 (N_17970,N_14706,N_13663);
and U17971 (N_17971,N_12270,N_14206);
or U17972 (N_17972,N_13624,N_12026);
and U17973 (N_17973,N_10927,N_12439);
nand U17974 (N_17974,N_10653,N_14090);
nand U17975 (N_17975,N_11797,N_12182);
nand U17976 (N_17976,N_12823,N_11874);
nand U17977 (N_17977,N_11482,N_13922);
nor U17978 (N_17978,N_10443,N_14504);
or U17979 (N_17979,N_10500,N_11625);
and U17980 (N_17980,N_11423,N_11648);
nor U17981 (N_17981,N_11655,N_13849);
and U17982 (N_17982,N_11380,N_11838);
nand U17983 (N_17983,N_14787,N_10832);
nor U17984 (N_17984,N_11533,N_13948);
nand U17985 (N_17985,N_13009,N_10025);
nor U17986 (N_17986,N_10785,N_11481);
and U17987 (N_17987,N_11226,N_14447);
nand U17988 (N_17988,N_12354,N_11052);
nand U17989 (N_17989,N_10125,N_11983);
nor U17990 (N_17990,N_11078,N_13245);
or U17991 (N_17991,N_13330,N_12277);
nor U17992 (N_17992,N_13413,N_14229);
xnor U17993 (N_17993,N_13469,N_12763);
nor U17994 (N_17994,N_11223,N_12232);
or U17995 (N_17995,N_14539,N_11767);
or U17996 (N_17996,N_11307,N_11658);
nand U17997 (N_17997,N_10646,N_13583);
nand U17998 (N_17998,N_10450,N_14922);
or U17999 (N_17999,N_12566,N_12416);
and U18000 (N_18000,N_11006,N_14056);
or U18001 (N_18001,N_11667,N_13841);
nand U18002 (N_18002,N_11793,N_13704);
xnor U18003 (N_18003,N_12695,N_12409);
nor U18004 (N_18004,N_14815,N_11567);
nor U18005 (N_18005,N_13061,N_14482);
nor U18006 (N_18006,N_12915,N_12234);
nor U18007 (N_18007,N_14878,N_14918);
nor U18008 (N_18008,N_10783,N_12879);
and U18009 (N_18009,N_11949,N_13556);
nor U18010 (N_18010,N_14361,N_14841);
nand U18011 (N_18011,N_13646,N_12322);
or U18012 (N_18012,N_11195,N_14015);
and U18013 (N_18013,N_11256,N_13851);
and U18014 (N_18014,N_14723,N_12771);
nor U18015 (N_18015,N_12981,N_12963);
and U18016 (N_18016,N_10223,N_13787);
and U18017 (N_18017,N_14221,N_11583);
or U18018 (N_18018,N_14794,N_11264);
nor U18019 (N_18019,N_11013,N_10390);
and U18020 (N_18020,N_13803,N_11461);
nor U18021 (N_18021,N_14017,N_13023);
nor U18022 (N_18022,N_12436,N_14859);
and U18023 (N_18023,N_12023,N_14323);
and U18024 (N_18024,N_11768,N_11780);
nand U18025 (N_18025,N_11366,N_10214);
xor U18026 (N_18026,N_10447,N_13965);
nand U18027 (N_18027,N_11629,N_14597);
nand U18028 (N_18028,N_14359,N_10159);
nand U18029 (N_18029,N_11064,N_10668);
xnor U18030 (N_18030,N_10429,N_11252);
and U18031 (N_18031,N_12933,N_12316);
nand U18032 (N_18032,N_12908,N_10273);
nor U18033 (N_18033,N_13747,N_10523);
nor U18034 (N_18034,N_11929,N_14297);
or U18035 (N_18035,N_11348,N_12127);
or U18036 (N_18036,N_11185,N_14096);
nand U18037 (N_18037,N_12489,N_11277);
nand U18038 (N_18038,N_12411,N_11956);
nand U18039 (N_18039,N_13692,N_10502);
nand U18040 (N_18040,N_10094,N_13151);
and U18041 (N_18041,N_14789,N_12192);
nand U18042 (N_18042,N_13848,N_10979);
nor U18043 (N_18043,N_11794,N_14532);
nor U18044 (N_18044,N_11123,N_12439);
or U18045 (N_18045,N_12512,N_12730);
or U18046 (N_18046,N_11216,N_14752);
nand U18047 (N_18047,N_12148,N_11893);
or U18048 (N_18048,N_14296,N_13605);
or U18049 (N_18049,N_10954,N_12979);
or U18050 (N_18050,N_10225,N_13170);
or U18051 (N_18051,N_13329,N_13019);
nor U18052 (N_18052,N_12976,N_11626);
and U18053 (N_18053,N_10157,N_10572);
or U18054 (N_18054,N_12258,N_10354);
nand U18055 (N_18055,N_11186,N_11182);
nor U18056 (N_18056,N_13157,N_11984);
nand U18057 (N_18057,N_14227,N_14543);
and U18058 (N_18058,N_13937,N_11858);
and U18059 (N_18059,N_14580,N_11218);
and U18060 (N_18060,N_10053,N_13022);
nand U18061 (N_18061,N_10361,N_14648);
and U18062 (N_18062,N_11549,N_10156);
and U18063 (N_18063,N_13746,N_12460);
nor U18064 (N_18064,N_13336,N_12037);
and U18065 (N_18065,N_11268,N_14243);
and U18066 (N_18066,N_10435,N_10731);
nand U18067 (N_18067,N_14642,N_14080);
or U18068 (N_18068,N_10594,N_14824);
or U18069 (N_18069,N_11517,N_11881);
nor U18070 (N_18070,N_12476,N_13028);
or U18071 (N_18071,N_14228,N_14285);
and U18072 (N_18072,N_13418,N_10004);
or U18073 (N_18073,N_11850,N_13109);
and U18074 (N_18074,N_13278,N_13869);
nor U18075 (N_18075,N_13187,N_11516);
nor U18076 (N_18076,N_10816,N_12119);
nand U18077 (N_18077,N_13992,N_13418);
nand U18078 (N_18078,N_13090,N_10661);
nand U18079 (N_18079,N_14599,N_12422);
nand U18080 (N_18080,N_13154,N_12694);
nor U18081 (N_18081,N_14896,N_13152);
and U18082 (N_18082,N_13453,N_10396);
nor U18083 (N_18083,N_14827,N_12657);
nor U18084 (N_18084,N_11700,N_11193);
or U18085 (N_18085,N_10143,N_13850);
nor U18086 (N_18086,N_10509,N_14549);
or U18087 (N_18087,N_14137,N_11035);
and U18088 (N_18088,N_10254,N_14813);
or U18089 (N_18089,N_13440,N_14608);
nand U18090 (N_18090,N_14578,N_13124);
nor U18091 (N_18091,N_10642,N_12671);
nand U18092 (N_18092,N_12325,N_12647);
nand U18093 (N_18093,N_11013,N_12169);
nand U18094 (N_18094,N_10961,N_12896);
nor U18095 (N_18095,N_14969,N_11332);
or U18096 (N_18096,N_10964,N_10052);
nand U18097 (N_18097,N_12364,N_13052);
or U18098 (N_18098,N_12146,N_11162);
nor U18099 (N_18099,N_14004,N_10155);
nor U18100 (N_18100,N_14395,N_13477);
nand U18101 (N_18101,N_10600,N_12892);
nand U18102 (N_18102,N_11316,N_13125);
nor U18103 (N_18103,N_11662,N_12440);
nand U18104 (N_18104,N_12748,N_13451);
or U18105 (N_18105,N_11299,N_10764);
nand U18106 (N_18106,N_10331,N_14959);
or U18107 (N_18107,N_11068,N_12789);
nor U18108 (N_18108,N_10889,N_11186);
nand U18109 (N_18109,N_13620,N_13700);
and U18110 (N_18110,N_14679,N_10306);
nand U18111 (N_18111,N_10818,N_10058);
and U18112 (N_18112,N_11632,N_13621);
xor U18113 (N_18113,N_11687,N_14632);
nor U18114 (N_18114,N_11922,N_13116);
and U18115 (N_18115,N_12234,N_12020);
or U18116 (N_18116,N_10032,N_12851);
and U18117 (N_18117,N_14901,N_12551);
or U18118 (N_18118,N_12810,N_14058);
xnor U18119 (N_18119,N_12767,N_10385);
or U18120 (N_18120,N_13364,N_13306);
and U18121 (N_18121,N_14872,N_11392);
nand U18122 (N_18122,N_12449,N_10095);
nor U18123 (N_18123,N_10003,N_10320);
nor U18124 (N_18124,N_12434,N_10934);
or U18125 (N_18125,N_14060,N_14552);
nand U18126 (N_18126,N_11929,N_11702);
and U18127 (N_18127,N_11313,N_12640);
or U18128 (N_18128,N_14502,N_11076);
nor U18129 (N_18129,N_12363,N_11373);
and U18130 (N_18130,N_12150,N_10437);
nor U18131 (N_18131,N_13447,N_14839);
nor U18132 (N_18132,N_11059,N_10435);
nand U18133 (N_18133,N_14737,N_10198);
and U18134 (N_18134,N_10330,N_11126);
or U18135 (N_18135,N_13168,N_11434);
or U18136 (N_18136,N_12754,N_11541);
nand U18137 (N_18137,N_13093,N_10338);
nand U18138 (N_18138,N_14224,N_10771);
and U18139 (N_18139,N_14020,N_13222);
and U18140 (N_18140,N_12802,N_10254);
nand U18141 (N_18141,N_10608,N_11773);
nor U18142 (N_18142,N_11441,N_12932);
or U18143 (N_18143,N_12300,N_14849);
nor U18144 (N_18144,N_10389,N_13872);
nor U18145 (N_18145,N_12649,N_14506);
and U18146 (N_18146,N_10609,N_10282);
nand U18147 (N_18147,N_13347,N_12391);
or U18148 (N_18148,N_11899,N_12694);
and U18149 (N_18149,N_11813,N_13938);
nor U18150 (N_18150,N_13815,N_10847);
or U18151 (N_18151,N_14493,N_11883);
nand U18152 (N_18152,N_11769,N_14132);
nand U18153 (N_18153,N_10323,N_12977);
nor U18154 (N_18154,N_11281,N_14373);
nor U18155 (N_18155,N_10809,N_12784);
nand U18156 (N_18156,N_10221,N_13615);
nand U18157 (N_18157,N_10476,N_14716);
nor U18158 (N_18158,N_11725,N_13927);
and U18159 (N_18159,N_10868,N_12468);
nand U18160 (N_18160,N_10903,N_12714);
nor U18161 (N_18161,N_12794,N_14944);
nor U18162 (N_18162,N_10713,N_14518);
nand U18163 (N_18163,N_11340,N_11963);
nor U18164 (N_18164,N_12439,N_12686);
nor U18165 (N_18165,N_11098,N_13393);
or U18166 (N_18166,N_13812,N_14954);
or U18167 (N_18167,N_13674,N_12959);
and U18168 (N_18168,N_10910,N_13969);
nand U18169 (N_18169,N_14117,N_14486);
nand U18170 (N_18170,N_12182,N_10802);
nor U18171 (N_18171,N_12773,N_12572);
nor U18172 (N_18172,N_12889,N_10855);
nor U18173 (N_18173,N_14058,N_11337);
nand U18174 (N_18174,N_11606,N_13481);
nand U18175 (N_18175,N_14818,N_14657);
and U18176 (N_18176,N_11993,N_12729);
or U18177 (N_18177,N_12338,N_13868);
and U18178 (N_18178,N_11095,N_12525);
nor U18179 (N_18179,N_11692,N_13654);
nor U18180 (N_18180,N_14416,N_10091);
and U18181 (N_18181,N_11446,N_14606);
and U18182 (N_18182,N_11558,N_11301);
nand U18183 (N_18183,N_12047,N_12220);
and U18184 (N_18184,N_13488,N_11032);
or U18185 (N_18185,N_11461,N_14369);
and U18186 (N_18186,N_14982,N_13713);
or U18187 (N_18187,N_11000,N_13463);
nor U18188 (N_18188,N_12193,N_14655);
nor U18189 (N_18189,N_14947,N_10688);
nor U18190 (N_18190,N_11230,N_10941);
nand U18191 (N_18191,N_10783,N_11063);
and U18192 (N_18192,N_11285,N_13289);
nand U18193 (N_18193,N_11059,N_13621);
and U18194 (N_18194,N_14429,N_14208);
and U18195 (N_18195,N_10725,N_11455);
or U18196 (N_18196,N_12787,N_14557);
nand U18197 (N_18197,N_13885,N_14566);
and U18198 (N_18198,N_11595,N_14580);
and U18199 (N_18199,N_11572,N_11732);
nor U18200 (N_18200,N_14308,N_14230);
or U18201 (N_18201,N_10241,N_10395);
and U18202 (N_18202,N_14116,N_11217);
nor U18203 (N_18203,N_14602,N_12060);
and U18204 (N_18204,N_12510,N_13390);
nand U18205 (N_18205,N_10728,N_13576);
or U18206 (N_18206,N_11373,N_11488);
nand U18207 (N_18207,N_11028,N_14103);
or U18208 (N_18208,N_12053,N_14605);
or U18209 (N_18209,N_13621,N_10307);
nor U18210 (N_18210,N_10059,N_12889);
and U18211 (N_18211,N_12783,N_11987);
or U18212 (N_18212,N_13463,N_10403);
and U18213 (N_18213,N_14827,N_14936);
nand U18214 (N_18214,N_13195,N_11263);
nor U18215 (N_18215,N_11999,N_10274);
or U18216 (N_18216,N_14708,N_12213);
nand U18217 (N_18217,N_14739,N_12502);
nand U18218 (N_18218,N_10474,N_14002);
nand U18219 (N_18219,N_12816,N_12988);
nand U18220 (N_18220,N_11301,N_12251);
nand U18221 (N_18221,N_12209,N_11288);
nor U18222 (N_18222,N_10359,N_14058);
nand U18223 (N_18223,N_13886,N_10779);
nor U18224 (N_18224,N_10708,N_10568);
or U18225 (N_18225,N_12369,N_13750);
or U18226 (N_18226,N_12633,N_14096);
or U18227 (N_18227,N_13773,N_10143);
and U18228 (N_18228,N_14931,N_14742);
and U18229 (N_18229,N_11730,N_10791);
nor U18230 (N_18230,N_11885,N_14923);
or U18231 (N_18231,N_10496,N_11105);
nor U18232 (N_18232,N_14578,N_11118);
xor U18233 (N_18233,N_11085,N_10482);
or U18234 (N_18234,N_11530,N_13005);
nand U18235 (N_18235,N_12115,N_14942);
and U18236 (N_18236,N_14091,N_14791);
xor U18237 (N_18237,N_12474,N_13222);
nand U18238 (N_18238,N_10965,N_14594);
or U18239 (N_18239,N_13105,N_11067);
nor U18240 (N_18240,N_13798,N_12168);
nand U18241 (N_18241,N_11951,N_13115);
or U18242 (N_18242,N_11572,N_14808);
nand U18243 (N_18243,N_10744,N_13502);
nor U18244 (N_18244,N_12237,N_12366);
nand U18245 (N_18245,N_10549,N_11934);
nor U18246 (N_18246,N_12382,N_14321);
and U18247 (N_18247,N_14486,N_14315);
nor U18248 (N_18248,N_10444,N_13121);
and U18249 (N_18249,N_12322,N_12732);
or U18250 (N_18250,N_14576,N_13153);
and U18251 (N_18251,N_12030,N_13351);
or U18252 (N_18252,N_12465,N_11993);
or U18253 (N_18253,N_14959,N_11527);
nor U18254 (N_18254,N_14630,N_13534);
xor U18255 (N_18255,N_13238,N_14279);
nor U18256 (N_18256,N_10295,N_14687);
and U18257 (N_18257,N_14220,N_12416);
or U18258 (N_18258,N_13201,N_12830);
or U18259 (N_18259,N_12190,N_10604);
and U18260 (N_18260,N_14864,N_13683);
nor U18261 (N_18261,N_10403,N_13414);
and U18262 (N_18262,N_14281,N_12429);
nor U18263 (N_18263,N_13408,N_11893);
and U18264 (N_18264,N_13081,N_11187);
nor U18265 (N_18265,N_11849,N_14824);
and U18266 (N_18266,N_12084,N_14038);
and U18267 (N_18267,N_13436,N_14758);
or U18268 (N_18268,N_11677,N_11809);
nand U18269 (N_18269,N_12137,N_14958);
or U18270 (N_18270,N_10334,N_12487);
nand U18271 (N_18271,N_14944,N_14970);
and U18272 (N_18272,N_14291,N_14724);
nand U18273 (N_18273,N_13273,N_11975);
and U18274 (N_18274,N_12849,N_11416);
or U18275 (N_18275,N_12602,N_11634);
or U18276 (N_18276,N_11823,N_12967);
nand U18277 (N_18277,N_14640,N_13671);
nor U18278 (N_18278,N_11061,N_14274);
and U18279 (N_18279,N_14506,N_11106);
nor U18280 (N_18280,N_10568,N_11565);
or U18281 (N_18281,N_12474,N_10954);
nor U18282 (N_18282,N_10885,N_13266);
nor U18283 (N_18283,N_11347,N_11642);
nor U18284 (N_18284,N_14373,N_14392);
or U18285 (N_18285,N_11082,N_12961);
and U18286 (N_18286,N_14846,N_14081);
nor U18287 (N_18287,N_14680,N_10358);
or U18288 (N_18288,N_13483,N_10196);
and U18289 (N_18289,N_14657,N_12939);
nor U18290 (N_18290,N_13286,N_12453);
nand U18291 (N_18291,N_11120,N_12660);
nand U18292 (N_18292,N_11237,N_11880);
nor U18293 (N_18293,N_11645,N_10794);
nand U18294 (N_18294,N_12702,N_11409);
nand U18295 (N_18295,N_12557,N_13676);
xnor U18296 (N_18296,N_13135,N_11072);
and U18297 (N_18297,N_11318,N_11231);
and U18298 (N_18298,N_13173,N_14552);
nand U18299 (N_18299,N_14833,N_12170);
xnor U18300 (N_18300,N_10127,N_14226);
and U18301 (N_18301,N_12682,N_13476);
and U18302 (N_18302,N_10268,N_14710);
nor U18303 (N_18303,N_10683,N_11193);
nand U18304 (N_18304,N_11445,N_12926);
nor U18305 (N_18305,N_12712,N_10937);
and U18306 (N_18306,N_12913,N_14064);
nor U18307 (N_18307,N_14219,N_13927);
and U18308 (N_18308,N_13771,N_11881);
nand U18309 (N_18309,N_13582,N_13455);
nand U18310 (N_18310,N_13748,N_11691);
nand U18311 (N_18311,N_11343,N_13010);
nand U18312 (N_18312,N_12341,N_11203);
nor U18313 (N_18313,N_12041,N_12353);
nand U18314 (N_18314,N_12526,N_10512);
nand U18315 (N_18315,N_10525,N_13764);
nand U18316 (N_18316,N_13855,N_11989);
or U18317 (N_18317,N_12266,N_12011);
xor U18318 (N_18318,N_13792,N_13734);
and U18319 (N_18319,N_11374,N_12790);
nor U18320 (N_18320,N_11652,N_14363);
nor U18321 (N_18321,N_13549,N_12386);
or U18322 (N_18322,N_12589,N_13133);
and U18323 (N_18323,N_14124,N_10763);
and U18324 (N_18324,N_12080,N_10855);
and U18325 (N_18325,N_11244,N_10833);
nor U18326 (N_18326,N_14582,N_11439);
nor U18327 (N_18327,N_12083,N_12226);
or U18328 (N_18328,N_12097,N_12700);
nand U18329 (N_18329,N_12735,N_11274);
and U18330 (N_18330,N_11861,N_11598);
nor U18331 (N_18331,N_13168,N_11374);
nand U18332 (N_18332,N_12860,N_13286);
nor U18333 (N_18333,N_10092,N_12739);
nand U18334 (N_18334,N_12141,N_13928);
nand U18335 (N_18335,N_12744,N_10991);
nor U18336 (N_18336,N_14700,N_14194);
or U18337 (N_18337,N_14533,N_11168);
or U18338 (N_18338,N_10892,N_12719);
nor U18339 (N_18339,N_13037,N_13333);
nor U18340 (N_18340,N_11632,N_11391);
and U18341 (N_18341,N_11917,N_14182);
nor U18342 (N_18342,N_10839,N_14339);
or U18343 (N_18343,N_12649,N_13712);
and U18344 (N_18344,N_11398,N_12834);
or U18345 (N_18345,N_13195,N_13921);
nand U18346 (N_18346,N_13002,N_13793);
or U18347 (N_18347,N_11739,N_12631);
and U18348 (N_18348,N_13337,N_13649);
and U18349 (N_18349,N_14534,N_11384);
or U18350 (N_18350,N_14687,N_11510);
nand U18351 (N_18351,N_12658,N_14634);
or U18352 (N_18352,N_14459,N_11024);
and U18353 (N_18353,N_12587,N_13650);
nand U18354 (N_18354,N_12120,N_14111);
or U18355 (N_18355,N_10148,N_14918);
nand U18356 (N_18356,N_10915,N_11882);
nand U18357 (N_18357,N_13458,N_14109);
and U18358 (N_18358,N_12394,N_10312);
nor U18359 (N_18359,N_13003,N_12076);
nand U18360 (N_18360,N_14270,N_10821);
or U18361 (N_18361,N_11965,N_10217);
and U18362 (N_18362,N_14884,N_12791);
nand U18363 (N_18363,N_14011,N_10294);
nor U18364 (N_18364,N_14521,N_11412);
or U18365 (N_18365,N_12930,N_13323);
nand U18366 (N_18366,N_14937,N_10230);
or U18367 (N_18367,N_10296,N_10739);
or U18368 (N_18368,N_10534,N_10676);
nand U18369 (N_18369,N_14760,N_13883);
nor U18370 (N_18370,N_11640,N_11571);
nor U18371 (N_18371,N_12488,N_11820);
and U18372 (N_18372,N_10270,N_10301);
nand U18373 (N_18373,N_11607,N_10336);
nand U18374 (N_18374,N_13739,N_10561);
nand U18375 (N_18375,N_13709,N_10341);
nand U18376 (N_18376,N_14460,N_13504);
and U18377 (N_18377,N_13603,N_12783);
and U18378 (N_18378,N_13617,N_10136);
or U18379 (N_18379,N_12532,N_14721);
nand U18380 (N_18380,N_11254,N_11800);
or U18381 (N_18381,N_11299,N_12178);
or U18382 (N_18382,N_10038,N_10293);
and U18383 (N_18383,N_11633,N_10464);
xnor U18384 (N_18384,N_11289,N_10276);
and U18385 (N_18385,N_14581,N_14130);
xnor U18386 (N_18386,N_12212,N_12975);
or U18387 (N_18387,N_11722,N_14423);
nor U18388 (N_18388,N_11030,N_12849);
nor U18389 (N_18389,N_14268,N_10393);
nor U18390 (N_18390,N_14160,N_10697);
nand U18391 (N_18391,N_11140,N_12956);
or U18392 (N_18392,N_10827,N_13046);
nand U18393 (N_18393,N_12261,N_14977);
nand U18394 (N_18394,N_14293,N_11518);
and U18395 (N_18395,N_12580,N_11314);
nor U18396 (N_18396,N_11693,N_12671);
and U18397 (N_18397,N_11413,N_14696);
nor U18398 (N_18398,N_13482,N_13244);
nand U18399 (N_18399,N_14914,N_10758);
or U18400 (N_18400,N_10497,N_14925);
nand U18401 (N_18401,N_13306,N_14385);
nor U18402 (N_18402,N_10107,N_11844);
or U18403 (N_18403,N_10122,N_14880);
nor U18404 (N_18404,N_14453,N_13663);
nor U18405 (N_18405,N_11269,N_10970);
and U18406 (N_18406,N_12094,N_13538);
and U18407 (N_18407,N_13780,N_14943);
or U18408 (N_18408,N_12144,N_10473);
and U18409 (N_18409,N_12231,N_11650);
xnor U18410 (N_18410,N_12528,N_12779);
nand U18411 (N_18411,N_13902,N_10812);
nor U18412 (N_18412,N_14668,N_10233);
nand U18413 (N_18413,N_10697,N_14985);
and U18414 (N_18414,N_11890,N_13838);
nand U18415 (N_18415,N_14277,N_14045);
nor U18416 (N_18416,N_11070,N_14727);
nor U18417 (N_18417,N_12049,N_14739);
nor U18418 (N_18418,N_13159,N_13225);
nand U18419 (N_18419,N_14758,N_11756);
nor U18420 (N_18420,N_14251,N_13206);
or U18421 (N_18421,N_14668,N_10727);
nor U18422 (N_18422,N_12230,N_14828);
and U18423 (N_18423,N_14040,N_14494);
nand U18424 (N_18424,N_10160,N_10553);
nor U18425 (N_18425,N_12895,N_12237);
nand U18426 (N_18426,N_14761,N_14109);
or U18427 (N_18427,N_13940,N_10732);
and U18428 (N_18428,N_12888,N_10309);
and U18429 (N_18429,N_14469,N_11595);
nand U18430 (N_18430,N_12766,N_10466);
and U18431 (N_18431,N_11095,N_10902);
nor U18432 (N_18432,N_10500,N_12355);
nor U18433 (N_18433,N_13272,N_11538);
nand U18434 (N_18434,N_12304,N_14220);
nor U18435 (N_18435,N_13945,N_13213);
or U18436 (N_18436,N_13854,N_13346);
or U18437 (N_18437,N_11094,N_11591);
and U18438 (N_18438,N_13553,N_13840);
and U18439 (N_18439,N_14822,N_10533);
and U18440 (N_18440,N_11261,N_11750);
nand U18441 (N_18441,N_14634,N_14626);
and U18442 (N_18442,N_11964,N_14315);
or U18443 (N_18443,N_12289,N_11035);
and U18444 (N_18444,N_13515,N_10297);
nand U18445 (N_18445,N_11368,N_14905);
and U18446 (N_18446,N_12879,N_13868);
nor U18447 (N_18447,N_13692,N_14833);
and U18448 (N_18448,N_14294,N_11668);
nor U18449 (N_18449,N_14862,N_10613);
nor U18450 (N_18450,N_14722,N_11348);
or U18451 (N_18451,N_11440,N_11839);
nor U18452 (N_18452,N_14218,N_11259);
nor U18453 (N_18453,N_10653,N_14322);
nor U18454 (N_18454,N_13050,N_11637);
or U18455 (N_18455,N_12158,N_14677);
nor U18456 (N_18456,N_10558,N_12084);
nand U18457 (N_18457,N_12643,N_14095);
or U18458 (N_18458,N_11336,N_13749);
nor U18459 (N_18459,N_14547,N_10999);
nand U18460 (N_18460,N_14664,N_12141);
and U18461 (N_18461,N_12948,N_11827);
nand U18462 (N_18462,N_13052,N_14257);
and U18463 (N_18463,N_10458,N_11985);
and U18464 (N_18464,N_14897,N_12250);
nand U18465 (N_18465,N_13911,N_11307);
or U18466 (N_18466,N_11918,N_10106);
and U18467 (N_18467,N_10798,N_14030);
or U18468 (N_18468,N_11133,N_10636);
and U18469 (N_18469,N_11254,N_12551);
nand U18470 (N_18470,N_12390,N_13622);
and U18471 (N_18471,N_13800,N_12038);
nand U18472 (N_18472,N_11690,N_11581);
nor U18473 (N_18473,N_14348,N_12276);
or U18474 (N_18474,N_12853,N_12599);
nand U18475 (N_18475,N_10592,N_10198);
or U18476 (N_18476,N_10314,N_10527);
nor U18477 (N_18477,N_14248,N_11855);
and U18478 (N_18478,N_10615,N_10891);
nor U18479 (N_18479,N_11783,N_13375);
and U18480 (N_18480,N_11104,N_10274);
or U18481 (N_18481,N_14567,N_14890);
or U18482 (N_18482,N_12873,N_13403);
or U18483 (N_18483,N_12981,N_12834);
or U18484 (N_18484,N_14323,N_12496);
and U18485 (N_18485,N_14697,N_13302);
nor U18486 (N_18486,N_12022,N_12965);
nor U18487 (N_18487,N_14018,N_13204);
or U18488 (N_18488,N_11013,N_14300);
and U18489 (N_18489,N_11423,N_10094);
and U18490 (N_18490,N_12521,N_11406);
or U18491 (N_18491,N_11074,N_13758);
nor U18492 (N_18492,N_10904,N_11381);
nand U18493 (N_18493,N_13268,N_13235);
or U18494 (N_18494,N_14564,N_14821);
nand U18495 (N_18495,N_14781,N_12160);
xnor U18496 (N_18496,N_14852,N_12370);
or U18497 (N_18497,N_11634,N_10644);
nand U18498 (N_18498,N_10655,N_12216);
nor U18499 (N_18499,N_12445,N_14021);
nor U18500 (N_18500,N_10948,N_13575);
or U18501 (N_18501,N_14943,N_10627);
nor U18502 (N_18502,N_11472,N_11847);
nor U18503 (N_18503,N_13689,N_14927);
or U18504 (N_18504,N_10984,N_14153);
xnor U18505 (N_18505,N_10958,N_11881);
nor U18506 (N_18506,N_12987,N_13531);
or U18507 (N_18507,N_13117,N_11260);
nor U18508 (N_18508,N_11584,N_14294);
nor U18509 (N_18509,N_12909,N_14080);
nor U18510 (N_18510,N_12610,N_13136);
nor U18511 (N_18511,N_14477,N_13084);
nor U18512 (N_18512,N_13405,N_12262);
and U18513 (N_18513,N_13251,N_11849);
or U18514 (N_18514,N_14710,N_10095);
and U18515 (N_18515,N_11508,N_12129);
and U18516 (N_18516,N_12064,N_12284);
and U18517 (N_18517,N_11550,N_11217);
nor U18518 (N_18518,N_14796,N_12055);
and U18519 (N_18519,N_14324,N_14391);
and U18520 (N_18520,N_13195,N_12969);
and U18521 (N_18521,N_11958,N_10897);
or U18522 (N_18522,N_10912,N_14822);
nand U18523 (N_18523,N_11297,N_11147);
xnor U18524 (N_18524,N_10723,N_10172);
nand U18525 (N_18525,N_13229,N_14360);
nor U18526 (N_18526,N_14692,N_11205);
xnor U18527 (N_18527,N_10456,N_12535);
nand U18528 (N_18528,N_12248,N_11300);
or U18529 (N_18529,N_12271,N_13550);
nand U18530 (N_18530,N_13949,N_11919);
nor U18531 (N_18531,N_14290,N_13793);
and U18532 (N_18532,N_14499,N_14267);
nand U18533 (N_18533,N_14899,N_13955);
and U18534 (N_18534,N_12430,N_14487);
or U18535 (N_18535,N_10527,N_12078);
or U18536 (N_18536,N_14163,N_11435);
nand U18537 (N_18537,N_13520,N_10619);
nor U18538 (N_18538,N_13874,N_12895);
nand U18539 (N_18539,N_13328,N_10799);
or U18540 (N_18540,N_14908,N_12233);
and U18541 (N_18541,N_10847,N_10467);
and U18542 (N_18542,N_12945,N_10895);
nand U18543 (N_18543,N_12732,N_13335);
and U18544 (N_18544,N_13577,N_12863);
and U18545 (N_18545,N_12176,N_12626);
and U18546 (N_18546,N_14325,N_10634);
nand U18547 (N_18547,N_12533,N_11135);
nand U18548 (N_18548,N_13733,N_10614);
nor U18549 (N_18549,N_11057,N_13954);
and U18550 (N_18550,N_14762,N_11228);
and U18551 (N_18551,N_11704,N_12823);
or U18552 (N_18552,N_11586,N_14432);
nand U18553 (N_18553,N_13783,N_14923);
and U18554 (N_18554,N_11248,N_12135);
nand U18555 (N_18555,N_11959,N_12066);
xor U18556 (N_18556,N_12606,N_12725);
nor U18557 (N_18557,N_13808,N_13582);
or U18558 (N_18558,N_10077,N_11394);
or U18559 (N_18559,N_14196,N_12972);
nor U18560 (N_18560,N_13399,N_11552);
or U18561 (N_18561,N_10548,N_11563);
nand U18562 (N_18562,N_12186,N_10673);
or U18563 (N_18563,N_12986,N_14030);
or U18564 (N_18564,N_12932,N_14482);
xnor U18565 (N_18565,N_12644,N_10312);
nand U18566 (N_18566,N_13049,N_12598);
and U18567 (N_18567,N_10776,N_13355);
nand U18568 (N_18568,N_12373,N_10741);
or U18569 (N_18569,N_13235,N_14770);
or U18570 (N_18570,N_14455,N_14351);
nor U18571 (N_18571,N_11903,N_10216);
or U18572 (N_18572,N_10831,N_10125);
nand U18573 (N_18573,N_14237,N_14129);
nor U18574 (N_18574,N_10808,N_14358);
xnor U18575 (N_18575,N_11285,N_14244);
and U18576 (N_18576,N_13212,N_14678);
and U18577 (N_18577,N_12021,N_10384);
or U18578 (N_18578,N_10584,N_14917);
and U18579 (N_18579,N_11217,N_11072);
or U18580 (N_18580,N_13406,N_10021);
and U18581 (N_18581,N_12997,N_12354);
nor U18582 (N_18582,N_10183,N_12664);
nor U18583 (N_18583,N_13767,N_13395);
or U18584 (N_18584,N_11037,N_11014);
and U18585 (N_18585,N_14917,N_13555);
or U18586 (N_18586,N_10211,N_10744);
and U18587 (N_18587,N_11676,N_12191);
nand U18588 (N_18588,N_11983,N_14124);
and U18589 (N_18589,N_13351,N_11457);
xor U18590 (N_18590,N_13292,N_13860);
or U18591 (N_18591,N_14914,N_14945);
nor U18592 (N_18592,N_10685,N_10265);
nor U18593 (N_18593,N_12038,N_11902);
nor U18594 (N_18594,N_11340,N_13115);
xor U18595 (N_18595,N_11749,N_10809);
nand U18596 (N_18596,N_13077,N_10316);
nor U18597 (N_18597,N_12909,N_14125);
or U18598 (N_18598,N_14155,N_11323);
nand U18599 (N_18599,N_11885,N_14348);
and U18600 (N_18600,N_10377,N_13434);
nand U18601 (N_18601,N_11668,N_12293);
nand U18602 (N_18602,N_12538,N_13243);
or U18603 (N_18603,N_10716,N_11783);
or U18604 (N_18604,N_13189,N_14543);
and U18605 (N_18605,N_12911,N_10510);
or U18606 (N_18606,N_10013,N_12974);
or U18607 (N_18607,N_10461,N_13031);
or U18608 (N_18608,N_13408,N_14844);
nor U18609 (N_18609,N_13933,N_12173);
nand U18610 (N_18610,N_13017,N_10383);
or U18611 (N_18611,N_11354,N_12246);
nand U18612 (N_18612,N_14540,N_12526);
nor U18613 (N_18613,N_13450,N_12757);
nand U18614 (N_18614,N_10989,N_10707);
or U18615 (N_18615,N_13213,N_13064);
nor U18616 (N_18616,N_12350,N_12837);
xnor U18617 (N_18617,N_10713,N_14045);
nor U18618 (N_18618,N_11315,N_14766);
nand U18619 (N_18619,N_10625,N_14656);
or U18620 (N_18620,N_10062,N_12432);
xnor U18621 (N_18621,N_14128,N_10554);
nand U18622 (N_18622,N_14756,N_10911);
xnor U18623 (N_18623,N_11680,N_12153);
nor U18624 (N_18624,N_10790,N_10351);
nor U18625 (N_18625,N_12333,N_13202);
nand U18626 (N_18626,N_13688,N_11707);
nor U18627 (N_18627,N_10273,N_11515);
or U18628 (N_18628,N_13812,N_14350);
and U18629 (N_18629,N_13670,N_11672);
or U18630 (N_18630,N_11195,N_14876);
or U18631 (N_18631,N_14766,N_11035);
or U18632 (N_18632,N_11237,N_10614);
and U18633 (N_18633,N_11462,N_13700);
and U18634 (N_18634,N_12978,N_10245);
nand U18635 (N_18635,N_10636,N_11495);
nor U18636 (N_18636,N_12129,N_14520);
or U18637 (N_18637,N_14802,N_11255);
nand U18638 (N_18638,N_13059,N_11864);
and U18639 (N_18639,N_12231,N_13993);
or U18640 (N_18640,N_14410,N_11965);
nor U18641 (N_18641,N_14304,N_11089);
nor U18642 (N_18642,N_10658,N_12113);
and U18643 (N_18643,N_12063,N_11292);
and U18644 (N_18644,N_11502,N_10775);
nand U18645 (N_18645,N_10450,N_11788);
nand U18646 (N_18646,N_11909,N_13225);
nor U18647 (N_18647,N_13785,N_12704);
or U18648 (N_18648,N_12624,N_12411);
and U18649 (N_18649,N_13787,N_10815);
nand U18650 (N_18650,N_14060,N_14124);
or U18651 (N_18651,N_13929,N_12877);
nor U18652 (N_18652,N_12327,N_13392);
nand U18653 (N_18653,N_11601,N_12539);
or U18654 (N_18654,N_10829,N_13423);
and U18655 (N_18655,N_13556,N_13449);
nor U18656 (N_18656,N_11679,N_10453);
and U18657 (N_18657,N_10775,N_13450);
and U18658 (N_18658,N_13890,N_14826);
and U18659 (N_18659,N_12353,N_14620);
nand U18660 (N_18660,N_12661,N_12510);
or U18661 (N_18661,N_11574,N_12182);
nor U18662 (N_18662,N_12860,N_12182);
nand U18663 (N_18663,N_10150,N_10463);
nor U18664 (N_18664,N_13586,N_14756);
nor U18665 (N_18665,N_10612,N_12407);
or U18666 (N_18666,N_14533,N_13959);
nor U18667 (N_18667,N_12574,N_10584);
and U18668 (N_18668,N_11057,N_11924);
and U18669 (N_18669,N_13970,N_11492);
xnor U18670 (N_18670,N_13813,N_14332);
or U18671 (N_18671,N_11856,N_11028);
and U18672 (N_18672,N_14652,N_10786);
or U18673 (N_18673,N_11813,N_10852);
and U18674 (N_18674,N_12028,N_10564);
or U18675 (N_18675,N_11659,N_12957);
nand U18676 (N_18676,N_11457,N_12527);
nor U18677 (N_18677,N_14385,N_13243);
or U18678 (N_18678,N_12909,N_12618);
nor U18679 (N_18679,N_11435,N_12209);
nand U18680 (N_18680,N_13424,N_12999);
or U18681 (N_18681,N_11305,N_14867);
or U18682 (N_18682,N_10556,N_14237);
nor U18683 (N_18683,N_14259,N_10867);
nor U18684 (N_18684,N_14108,N_10384);
nand U18685 (N_18685,N_12411,N_11111);
xnor U18686 (N_18686,N_12688,N_13977);
nor U18687 (N_18687,N_13433,N_12748);
nor U18688 (N_18688,N_12636,N_13230);
and U18689 (N_18689,N_14506,N_14254);
xor U18690 (N_18690,N_10020,N_11797);
or U18691 (N_18691,N_11535,N_10262);
or U18692 (N_18692,N_14371,N_11830);
or U18693 (N_18693,N_10278,N_11679);
and U18694 (N_18694,N_10593,N_11001);
or U18695 (N_18695,N_14778,N_14290);
nor U18696 (N_18696,N_13620,N_14628);
and U18697 (N_18697,N_12716,N_10184);
nor U18698 (N_18698,N_12090,N_14455);
and U18699 (N_18699,N_11480,N_10897);
or U18700 (N_18700,N_14937,N_14073);
nor U18701 (N_18701,N_14254,N_10193);
nor U18702 (N_18702,N_12592,N_14050);
nor U18703 (N_18703,N_12408,N_11694);
and U18704 (N_18704,N_10938,N_14639);
and U18705 (N_18705,N_11990,N_11873);
nor U18706 (N_18706,N_13248,N_11130);
nor U18707 (N_18707,N_14316,N_12085);
or U18708 (N_18708,N_12315,N_13919);
nand U18709 (N_18709,N_11952,N_14411);
and U18710 (N_18710,N_12059,N_10085);
xor U18711 (N_18711,N_14637,N_10847);
or U18712 (N_18712,N_14978,N_12260);
or U18713 (N_18713,N_13468,N_10237);
or U18714 (N_18714,N_11098,N_13092);
nor U18715 (N_18715,N_13956,N_10781);
nor U18716 (N_18716,N_14322,N_14213);
nand U18717 (N_18717,N_14774,N_11677);
and U18718 (N_18718,N_11225,N_13726);
nand U18719 (N_18719,N_12055,N_10054);
nor U18720 (N_18720,N_10011,N_12888);
nand U18721 (N_18721,N_10000,N_11841);
and U18722 (N_18722,N_14173,N_11158);
or U18723 (N_18723,N_14108,N_10512);
or U18724 (N_18724,N_10864,N_10115);
nand U18725 (N_18725,N_10063,N_10066);
nor U18726 (N_18726,N_11760,N_12622);
xor U18727 (N_18727,N_11829,N_14875);
and U18728 (N_18728,N_12804,N_10992);
nand U18729 (N_18729,N_13072,N_14516);
or U18730 (N_18730,N_14761,N_14727);
and U18731 (N_18731,N_14239,N_14679);
nor U18732 (N_18732,N_14582,N_12126);
nand U18733 (N_18733,N_14574,N_10291);
nand U18734 (N_18734,N_14526,N_12609);
nor U18735 (N_18735,N_12064,N_13649);
or U18736 (N_18736,N_10177,N_10988);
nand U18737 (N_18737,N_11799,N_10960);
nand U18738 (N_18738,N_12439,N_12667);
and U18739 (N_18739,N_10748,N_13045);
or U18740 (N_18740,N_12406,N_11584);
nand U18741 (N_18741,N_14416,N_13729);
or U18742 (N_18742,N_13963,N_14323);
nand U18743 (N_18743,N_14422,N_13864);
nor U18744 (N_18744,N_13769,N_11962);
or U18745 (N_18745,N_12450,N_14200);
or U18746 (N_18746,N_13078,N_12603);
nand U18747 (N_18747,N_10884,N_14694);
or U18748 (N_18748,N_12843,N_11961);
or U18749 (N_18749,N_10941,N_12210);
nand U18750 (N_18750,N_14622,N_12817);
and U18751 (N_18751,N_11267,N_11185);
nand U18752 (N_18752,N_12134,N_11731);
and U18753 (N_18753,N_11141,N_10797);
or U18754 (N_18754,N_11314,N_12599);
or U18755 (N_18755,N_13072,N_10983);
nand U18756 (N_18756,N_10501,N_10293);
nand U18757 (N_18757,N_12766,N_10314);
nand U18758 (N_18758,N_13296,N_14926);
or U18759 (N_18759,N_10935,N_13166);
nor U18760 (N_18760,N_11703,N_12086);
nor U18761 (N_18761,N_12413,N_13931);
and U18762 (N_18762,N_12133,N_12693);
nor U18763 (N_18763,N_14750,N_12551);
nand U18764 (N_18764,N_12595,N_10344);
or U18765 (N_18765,N_12122,N_12467);
nand U18766 (N_18766,N_13866,N_11322);
xnor U18767 (N_18767,N_11092,N_10236);
or U18768 (N_18768,N_13633,N_11729);
or U18769 (N_18769,N_14193,N_11233);
and U18770 (N_18770,N_13148,N_14645);
or U18771 (N_18771,N_13992,N_10218);
nor U18772 (N_18772,N_10776,N_10134);
nor U18773 (N_18773,N_11940,N_13003);
or U18774 (N_18774,N_13256,N_13106);
or U18775 (N_18775,N_10752,N_12745);
or U18776 (N_18776,N_14414,N_13498);
nor U18777 (N_18777,N_13684,N_14470);
and U18778 (N_18778,N_10725,N_11672);
or U18779 (N_18779,N_14742,N_13565);
or U18780 (N_18780,N_10315,N_10236);
and U18781 (N_18781,N_14881,N_14547);
and U18782 (N_18782,N_12427,N_12846);
or U18783 (N_18783,N_11879,N_10898);
nor U18784 (N_18784,N_10101,N_13561);
and U18785 (N_18785,N_13691,N_14123);
or U18786 (N_18786,N_12020,N_13957);
nor U18787 (N_18787,N_14835,N_14260);
or U18788 (N_18788,N_14487,N_14948);
and U18789 (N_18789,N_10778,N_12454);
and U18790 (N_18790,N_14573,N_11964);
nor U18791 (N_18791,N_14802,N_12920);
nand U18792 (N_18792,N_11531,N_14268);
nand U18793 (N_18793,N_14455,N_13610);
nand U18794 (N_18794,N_10713,N_11064);
nand U18795 (N_18795,N_10472,N_13845);
nor U18796 (N_18796,N_10978,N_14287);
or U18797 (N_18797,N_14100,N_12702);
or U18798 (N_18798,N_12650,N_10131);
or U18799 (N_18799,N_10143,N_10923);
nor U18800 (N_18800,N_11051,N_13263);
nand U18801 (N_18801,N_11112,N_14288);
and U18802 (N_18802,N_12815,N_11251);
nor U18803 (N_18803,N_13081,N_10608);
nor U18804 (N_18804,N_12866,N_14559);
nor U18805 (N_18805,N_13084,N_13736);
nor U18806 (N_18806,N_11651,N_13876);
nand U18807 (N_18807,N_13924,N_12784);
and U18808 (N_18808,N_11085,N_11965);
or U18809 (N_18809,N_12075,N_14594);
nor U18810 (N_18810,N_12475,N_14379);
or U18811 (N_18811,N_10406,N_13774);
and U18812 (N_18812,N_10429,N_13914);
and U18813 (N_18813,N_13309,N_12548);
and U18814 (N_18814,N_11663,N_14137);
nor U18815 (N_18815,N_13990,N_12369);
or U18816 (N_18816,N_12787,N_11379);
or U18817 (N_18817,N_10005,N_11691);
or U18818 (N_18818,N_14668,N_11854);
nand U18819 (N_18819,N_10402,N_14507);
nand U18820 (N_18820,N_12082,N_11833);
or U18821 (N_18821,N_11323,N_13570);
nor U18822 (N_18822,N_12582,N_11725);
nor U18823 (N_18823,N_13747,N_10451);
and U18824 (N_18824,N_13921,N_13775);
nor U18825 (N_18825,N_12919,N_10197);
nand U18826 (N_18826,N_12439,N_11125);
nand U18827 (N_18827,N_12187,N_13840);
or U18828 (N_18828,N_13224,N_12215);
and U18829 (N_18829,N_14576,N_11344);
and U18830 (N_18830,N_13811,N_12893);
nor U18831 (N_18831,N_11125,N_13444);
nand U18832 (N_18832,N_12059,N_10129);
nor U18833 (N_18833,N_13670,N_14991);
or U18834 (N_18834,N_12905,N_14811);
nand U18835 (N_18835,N_10840,N_10401);
and U18836 (N_18836,N_13070,N_14574);
xnor U18837 (N_18837,N_12484,N_11947);
and U18838 (N_18838,N_12182,N_13567);
nor U18839 (N_18839,N_12298,N_12802);
nand U18840 (N_18840,N_11388,N_13471);
or U18841 (N_18841,N_10900,N_12515);
nand U18842 (N_18842,N_10898,N_11454);
and U18843 (N_18843,N_12131,N_10399);
and U18844 (N_18844,N_10575,N_12447);
nor U18845 (N_18845,N_14281,N_11065);
or U18846 (N_18846,N_11747,N_14720);
nand U18847 (N_18847,N_11316,N_14143);
or U18848 (N_18848,N_10550,N_11665);
or U18849 (N_18849,N_10286,N_11955);
nand U18850 (N_18850,N_10092,N_12813);
nor U18851 (N_18851,N_13502,N_13760);
or U18852 (N_18852,N_10462,N_12784);
or U18853 (N_18853,N_10608,N_12823);
nor U18854 (N_18854,N_12172,N_13703);
nor U18855 (N_18855,N_11651,N_14746);
nor U18856 (N_18856,N_14640,N_12100);
nor U18857 (N_18857,N_13873,N_14127);
or U18858 (N_18858,N_13537,N_12120);
or U18859 (N_18859,N_12475,N_13289);
and U18860 (N_18860,N_14692,N_11493);
nand U18861 (N_18861,N_11703,N_10892);
nand U18862 (N_18862,N_12853,N_13256);
nand U18863 (N_18863,N_14380,N_11480);
nand U18864 (N_18864,N_14239,N_14710);
and U18865 (N_18865,N_12887,N_10649);
or U18866 (N_18866,N_10345,N_10741);
or U18867 (N_18867,N_14621,N_10684);
nor U18868 (N_18868,N_12514,N_12687);
nand U18869 (N_18869,N_13794,N_12250);
or U18870 (N_18870,N_12332,N_10718);
or U18871 (N_18871,N_11167,N_14688);
or U18872 (N_18872,N_14317,N_13361);
nand U18873 (N_18873,N_12155,N_11939);
xnor U18874 (N_18874,N_14641,N_14131);
nor U18875 (N_18875,N_11681,N_12285);
or U18876 (N_18876,N_11815,N_12634);
xnor U18877 (N_18877,N_14916,N_10682);
nand U18878 (N_18878,N_11874,N_13619);
and U18879 (N_18879,N_14665,N_13279);
nor U18880 (N_18880,N_10967,N_11478);
nor U18881 (N_18881,N_14021,N_13420);
nor U18882 (N_18882,N_13321,N_11330);
nand U18883 (N_18883,N_12338,N_11659);
or U18884 (N_18884,N_13940,N_14329);
nor U18885 (N_18885,N_12901,N_13359);
or U18886 (N_18886,N_14931,N_13603);
and U18887 (N_18887,N_11591,N_14392);
and U18888 (N_18888,N_10388,N_13849);
or U18889 (N_18889,N_12304,N_14320);
nor U18890 (N_18890,N_13837,N_11141);
nor U18891 (N_18891,N_12280,N_10254);
nor U18892 (N_18892,N_11033,N_12982);
or U18893 (N_18893,N_11436,N_10943);
nand U18894 (N_18894,N_14460,N_11696);
nand U18895 (N_18895,N_13340,N_13482);
nand U18896 (N_18896,N_13649,N_11469);
or U18897 (N_18897,N_11714,N_14565);
or U18898 (N_18898,N_10686,N_14265);
or U18899 (N_18899,N_11059,N_10566);
or U18900 (N_18900,N_13501,N_10730);
nand U18901 (N_18901,N_14838,N_11960);
or U18902 (N_18902,N_10692,N_14591);
or U18903 (N_18903,N_12659,N_12382);
and U18904 (N_18904,N_11019,N_10441);
or U18905 (N_18905,N_10087,N_14466);
and U18906 (N_18906,N_14160,N_13713);
and U18907 (N_18907,N_14737,N_13337);
or U18908 (N_18908,N_14671,N_13401);
nand U18909 (N_18909,N_11532,N_10399);
or U18910 (N_18910,N_10705,N_11621);
nor U18911 (N_18911,N_14058,N_11524);
nand U18912 (N_18912,N_10246,N_12619);
or U18913 (N_18913,N_10988,N_14649);
and U18914 (N_18914,N_10572,N_14990);
nor U18915 (N_18915,N_12074,N_14353);
nor U18916 (N_18916,N_12333,N_11235);
or U18917 (N_18917,N_11671,N_13482);
nand U18918 (N_18918,N_14283,N_13631);
nand U18919 (N_18919,N_12993,N_10413);
and U18920 (N_18920,N_10301,N_13189);
or U18921 (N_18921,N_12922,N_10827);
and U18922 (N_18922,N_11187,N_12523);
nand U18923 (N_18923,N_11580,N_11959);
or U18924 (N_18924,N_10155,N_10644);
nand U18925 (N_18925,N_12195,N_12567);
and U18926 (N_18926,N_12389,N_12931);
and U18927 (N_18927,N_11997,N_13260);
nor U18928 (N_18928,N_13071,N_13542);
or U18929 (N_18929,N_11913,N_12607);
and U18930 (N_18930,N_10290,N_11746);
or U18931 (N_18931,N_14441,N_11942);
or U18932 (N_18932,N_10467,N_13251);
nor U18933 (N_18933,N_12932,N_13578);
nor U18934 (N_18934,N_10621,N_11806);
nor U18935 (N_18935,N_10991,N_13545);
and U18936 (N_18936,N_12537,N_13699);
or U18937 (N_18937,N_12360,N_11486);
nor U18938 (N_18938,N_14767,N_14215);
nor U18939 (N_18939,N_14847,N_11617);
nor U18940 (N_18940,N_14177,N_14998);
nand U18941 (N_18941,N_12710,N_10069);
nor U18942 (N_18942,N_13100,N_12109);
nor U18943 (N_18943,N_14963,N_13091);
or U18944 (N_18944,N_14591,N_13302);
nand U18945 (N_18945,N_14788,N_12935);
xnor U18946 (N_18946,N_12906,N_14785);
nor U18947 (N_18947,N_13741,N_12431);
or U18948 (N_18948,N_10548,N_13919);
or U18949 (N_18949,N_10229,N_10587);
and U18950 (N_18950,N_13804,N_13454);
xnor U18951 (N_18951,N_12829,N_11509);
or U18952 (N_18952,N_12619,N_13167);
nand U18953 (N_18953,N_11807,N_10526);
or U18954 (N_18954,N_14131,N_11337);
nor U18955 (N_18955,N_10943,N_12939);
and U18956 (N_18956,N_13032,N_11289);
and U18957 (N_18957,N_12722,N_10968);
or U18958 (N_18958,N_14427,N_14695);
nor U18959 (N_18959,N_13364,N_13510);
nor U18960 (N_18960,N_11584,N_13156);
or U18961 (N_18961,N_12858,N_10148);
and U18962 (N_18962,N_10991,N_12957);
or U18963 (N_18963,N_12433,N_10475);
nand U18964 (N_18964,N_14645,N_11841);
or U18965 (N_18965,N_11234,N_14167);
or U18966 (N_18966,N_14476,N_13576);
and U18967 (N_18967,N_13731,N_13564);
nor U18968 (N_18968,N_14846,N_13797);
nand U18969 (N_18969,N_11686,N_10309);
and U18970 (N_18970,N_11880,N_14625);
nor U18971 (N_18971,N_12686,N_13634);
nor U18972 (N_18972,N_11232,N_11693);
nand U18973 (N_18973,N_13892,N_12332);
and U18974 (N_18974,N_11169,N_11143);
nor U18975 (N_18975,N_13794,N_12275);
nor U18976 (N_18976,N_10003,N_10405);
nand U18977 (N_18977,N_13510,N_12047);
nand U18978 (N_18978,N_12236,N_13266);
nor U18979 (N_18979,N_10350,N_14338);
nor U18980 (N_18980,N_12658,N_12757);
or U18981 (N_18981,N_12386,N_10264);
nor U18982 (N_18982,N_11798,N_14281);
nand U18983 (N_18983,N_14721,N_10903);
nand U18984 (N_18984,N_14516,N_12745);
nand U18985 (N_18985,N_10505,N_14625);
nor U18986 (N_18986,N_11405,N_13956);
and U18987 (N_18987,N_14527,N_13362);
nand U18988 (N_18988,N_13673,N_11745);
nand U18989 (N_18989,N_13237,N_11550);
and U18990 (N_18990,N_13916,N_13238);
and U18991 (N_18991,N_10788,N_14592);
nor U18992 (N_18992,N_10425,N_10821);
and U18993 (N_18993,N_11140,N_14516);
nor U18994 (N_18994,N_11687,N_10503);
or U18995 (N_18995,N_12046,N_10840);
nor U18996 (N_18996,N_10589,N_13584);
and U18997 (N_18997,N_11222,N_14837);
nor U18998 (N_18998,N_11242,N_14637);
and U18999 (N_18999,N_14458,N_13961);
or U19000 (N_19000,N_11191,N_14387);
nor U19001 (N_19001,N_10965,N_12949);
nor U19002 (N_19002,N_12347,N_12422);
and U19003 (N_19003,N_14636,N_13345);
nor U19004 (N_19004,N_14571,N_10457);
and U19005 (N_19005,N_10277,N_13460);
nor U19006 (N_19006,N_10310,N_14387);
nand U19007 (N_19007,N_10103,N_13016);
nand U19008 (N_19008,N_14588,N_14310);
nand U19009 (N_19009,N_12855,N_12277);
or U19010 (N_19010,N_12836,N_14855);
and U19011 (N_19011,N_14744,N_13059);
and U19012 (N_19012,N_14493,N_11888);
nor U19013 (N_19013,N_13542,N_12929);
nor U19014 (N_19014,N_10903,N_14104);
or U19015 (N_19015,N_13152,N_11265);
and U19016 (N_19016,N_11989,N_14739);
nor U19017 (N_19017,N_13647,N_11185);
nor U19018 (N_19018,N_14392,N_13224);
nor U19019 (N_19019,N_14366,N_14636);
nand U19020 (N_19020,N_12914,N_14404);
nor U19021 (N_19021,N_14456,N_13959);
and U19022 (N_19022,N_12483,N_14605);
or U19023 (N_19023,N_14310,N_12452);
nand U19024 (N_19024,N_14056,N_12537);
or U19025 (N_19025,N_11905,N_14749);
nor U19026 (N_19026,N_11131,N_13773);
nand U19027 (N_19027,N_12375,N_11444);
or U19028 (N_19028,N_12493,N_12647);
and U19029 (N_19029,N_14046,N_14579);
or U19030 (N_19030,N_12835,N_14972);
nor U19031 (N_19031,N_11587,N_12434);
nand U19032 (N_19032,N_11748,N_11848);
and U19033 (N_19033,N_14417,N_13641);
nand U19034 (N_19034,N_14747,N_12839);
nand U19035 (N_19035,N_13503,N_13727);
or U19036 (N_19036,N_13889,N_13017);
or U19037 (N_19037,N_13110,N_14749);
or U19038 (N_19038,N_11777,N_14989);
and U19039 (N_19039,N_12769,N_13863);
or U19040 (N_19040,N_10996,N_12834);
and U19041 (N_19041,N_10473,N_14138);
and U19042 (N_19042,N_12092,N_10078);
nand U19043 (N_19043,N_11090,N_11068);
or U19044 (N_19044,N_10388,N_12183);
or U19045 (N_19045,N_12236,N_11737);
nand U19046 (N_19046,N_14753,N_14658);
or U19047 (N_19047,N_11229,N_11656);
or U19048 (N_19048,N_11131,N_14262);
or U19049 (N_19049,N_10608,N_13883);
and U19050 (N_19050,N_12922,N_13005);
and U19051 (N_19051,N_14852,N_12205);
and U19052 (N_19052,N_10281,N_12595);
nor U19053 (N_19053,N_11894,N_14371);
nand U19054 (N_19054,N_14163,N_14330);
nor U19055 (N_19055,N_11823,N_12693);
nor U19056 (N_19056,N_11323,N_12577);
nor U19057 (N_19057,N_11283,N_11493);
nor U19058 (N_19058,N_12162,N_10709);
nor U19059 (N_19059,N_11984,N_14286);
or U19060 (N_19060,N_14398,N_11808);
xnor U19061 (N_19061,N_14865,N_12853);
nand U19062 (N_19062,N_13225,N_13824);
and U19063 (N_19063,N_11088,N_10539);
or U19064 (N_19064,N_13299,N_11944);
and U19065 (N_19065,N_10132,N_11233);
and U19066 (N_19066,N_12597,N_14821);
nor U19067 (N_19067,N_11605,N_11672);
nand U19068 (N_19068,N_12521,N_11166);
and U19069 (N_19069,N_12280,N_13734);
and U19070 (N_19070,N_11089,N_10558);
nor U19071 (N_19071,N_14842,N_13026);
and U19072 (N_19072,N_10930,N_10377);
and U19073 (N_19073,N_13398,N_11195);
xnor U19074 (N_19074,N_11363,N_12048);
or U19075 (N_19075,N_14940,N_14709);
and U19076 (N_19076,N_10218,N_10176);
nand U19077 (N_19077,N_12427,N_11275);
nor U19078 (N_19078,N_11894,N_11153);
nor U19079 (N_19079,N_11886,N_13119);
and U19080 (N_19080,N_10443,N_10463);
and U19081 (N_19081,N_12412,N_12070);
nor U19082 (N_19082,N_13968,N_10842);
nand U19083 (N_19083,N_10541,N_13587);
or U19084 (N_19084,N_11764,N_10184);
and U19085 (N_19085,N_11180,N_12599);
nand U19086 (N_19086,N_14358,N_13865);
nor U19087 (N_19087,N_10145,N_12934);
xor U19088 (N_19088,N_14631,N_13118);
or U19089 (N_19089,N_13216,N_10598);
or U19090 (N_19090,N_11714,N_11543);
or U19091 (N_19091,N_12488,N_13674);
nor U19092 (N_19092,N_13596,N_11133);
nor U19093 (N_19093,N_14681,N_14948);
nand U19094 (N_19094,N_12370,N_10460);
nor U19095 (N_19095,N_10167,N_14436);
or U19096 (N_19096,N_10319,N_14886);
nand U19097 (N_19097,N_13198,N_13569);
nor U19098 (N_19098,N_11571,N_12997);
nand U19099 (N_19099,N_13651,N_10967);
nor U19100 (N_19100,N_13013,N_14602);
xor U19101 (N_19101,N_10246,N_13921);
nand U19102 (N_19102,N_12965,N_13427);
nand U19103 (N_19103,N_12353,N_13248);
and U19104 (N_19104,N_14005,N_11876);
and U19105 (N_19105,N_12423,N_11054);
and U19106 (N_19106,N_11964,N_14166);
or U19107 (N_19107,N_12445,N_14074);
or U19108 (N_19108,N_11891,N_13969);
xnor U19109 (N_19109,N_13313,N_10236);
and U19110 (N_19110,N_12758,N_12857);
nor U19111 (N_19111,N_14116,N_12889);
and U19112 (N_19112,N_12235,N_13754);
nand U19113 (N_19113,N_10311,N_10246);
and U19114 (N_19114,N_10356,N_12881);
xor U19115 (N_19115,N_13624,N_11683);
nor U19116 (N_19116,N_10120,N_13651);
nor U19117 (N_19117,N_10568,N_10192);
or U19118 (N_19118,N_12399,N_10711);
nor U19119 (N_19119,N_11035,N_10774);
nor U19120 (N_19120,N_12410,N_12417);
nand U19121 (N_19121,N_13031,N_13287);
nor U19122 (N_19122,N_12825,N_10032);
nor U19123 (N_19123,N_13805,N_10161);
and U19124 (N_19124,N_11272,N_10178);
nand U19125 (N_19125,N_10210,N_11125);
or U19126 (N_19126,N_12016,N_10541);
nand U19127 (N_19127,N_13173,N_14049);
or U19128 (N_19128,N_13140,N_12242);
or U19129 (N_19129,N_10095,N_11203);
and U19130 (N_19130,N_10052,N_11451);
nand U19131 (N_19131,N_14735,N_13345);
nand U19132 (N_19132,N_10111,N_14023);
nor U19133 (N_19133,N_14878,N_12440);
nand U19134 (N_19134,N_10095,N_13966);
nand U19135 (N_19135,N_10582,N_12267);
and U19136 (N_19136,N_10220,N_11503);
xnor U19137 (N_19137,N_10624,N_11722);
and U19138 (N_19138,N_10257,N_13552);
and U19139 (N_19139,N_13984,N_10312);
and U19140 (N_19140,N_12158,N_13576);
nor U19141 (N_19141,N_12694,N_14859);
nor U19142 (N_19142,N_10363,N_13767);
or U19143 (N_19143,N_11900,N_14137);
or U19144 (N_19144,N_12647,N_10474);
or U19145 (N_19145,N_12387,N_14009);
nand U19146 (N_19146,N_14494,N_13977);
nor U19147 (N_19147,N_11095,N_14186);
and U19148 (N_19148,N_14111,N_13305);
and U19149 (N_19149,N_10634,N_14283);
and U19150 (N_19150,N_10359,N_11740);
or U19151 (N_19151,N_14417,N_10352);
and U19152 (N_19152,N_11417,N_13290);
or U19153 (N_19153,N_12374,N_12139);
nor U19154 (N_19154,N_14235,N_10961);
nor U19155 (N_19155,N_10529,N_14263);
nand U19156 (N_19156,N_14942,N_13020);
nand U19157 (N_19157,N_12935,N_14189);
nand U19158 (N_19158,N_12502,N_12570);
or U19159 (N_19159,N_14005,N_12971);
or U19160 (N_19160,N_11395,N_11709);
or U19161 (N_19161,N_12768,N_14511);
nor U19162 (N_19162,N_11365,N_12850);
and U19163 (N_19163,N_10082,N_11167);
and U19164 (N_19164,N_12388,N_13520);
nand U19165 (N_19165,N_12641,N_12256);
nor U19166 (N_19166,N_10618,N_14193);
nand U19167 (N_19167,N_12284,N_13269);
or U19168 (N_19168,N_14883,N_13397);
xor U19169 (N_19169,N_10135,N_11128);
and U19170 (N_19170,N_11415,N_14140);
and U19171 (N_19171,N_10699,N_13852);
and U19172 (N_19172,N_10015,N_10805);
and U19173 (N_19173,N_10739,N_10220);
nand U19174 (N_19174,N_13323,N_10752);
or U19175 (N_19175,N_12581,N_10561);
and U19176 (N_19176,N_14616,N_13294);
nor U19177 (N_19177,N_11904,N_13886);
or U19178 (N_19178,N_10152,N_14161);
or U19179 (N_19179,N_14047,N_14018);
nor U19180 (N_19180,N_12293,N_12779);
nor U19181 (N_19181,N_14885,N_12494);
and U19182 (N_19182,N_13618,N_10710);
nor U19183 (N_19183,N_13893,N_12249);
and U19184 (N_19184,N_12776,N_14937);
nand U19185 (N_19185,N_13404,N_10858);
nand U19186 (N_19186,N_14290,N_13880);
nand U19187 (N_19187,N_13015,N_11071);
nor U19188 (N_19188,N_12549,N_11793);
nand U19189 (N_19189,N_12887,N_13678);
or U19190 (N_19190,N_13966,N_11869);
xor U19191 (N_19191,N_14253,N_12474);
nand U19192 (N_19192,N_13413,N_13638);
nand U19193 (N_19193,N_11639,N_13380);
or U19194 (N_19194,N_14777,N_12830);
nand U19195 (N_19195,N_13425,N_10769);
nor U19196 (N_19196,N_11593,N_11697);
nand U19197 (N_19197,N_10736,N_11071);
and U19198 (N_19198,N_14619,N_12314);
nand U19199 (N_19199,N_14694,N_14565);
nor U19200 (N_19200,N_12486,N_14757);
and U19201 (N_19201,N_10154,N_14527);
nand U19202 (N_19202,N_11120,N_11997);
nor U19203 (N_19203,N_14013,N_12720);
or U19204 (N_19204,N_14983,N_11696);
nor U19205 (N_19205,N_12836,N_12034);
nor U19206 (N_19206,N_13748,N_10768);
or U19207 (N_19207,N_10315,N_14698);
xnor U19208 (N_19208,N_14774,N_12820);
nor U19209 (N_19209,N_12357,N_13530);
and U19210 (N_19210,N_11114,N_11696);
or U19211 (N_19211,N_11874,N_11855);
nand U19212 (N_19212,N_10186,N_14280);
nor U19213 (N_19213,N_10045,N_12910);
nand U19214 (N_19214,N_10518,N_11425);
nand U19215 (N_19215,N_14921,N_10614);
nor U19216 (N_19216,N_10657,N_10511);
nand U19217 (N_19217,N_10226,N_13779);
nor U19218 (N_19218,N_12151,N_14798);
xnor U19219 (N_19219,N_10721,N_13126);
nand U19220 (N_19220,N_11680,N_11950);
or U19221 (N_19221,N_10156,N_13901);
nand U19222 (N_19222,N_12463,N_10956);
nor U19223 (N_19223,N_14899,N_14279);
nand U19224 (N_19224,N_13184,N_12239);
nor U19225 (N_19225,N_10901,N_13568);
nor U19226 (N_19226,N_14707,N_13364);
and U19227 (N_19227,N_12253,N_10889);
nor U19228 (N_19228,N_10760,N_10652);
and U19229 (N_19229,N_10598,N_13820);
nand U19230 (N_19230,N_13101,N_11144);
nor U19231 (N_19231,N_12431,N_13293);
nor U19232 (N_19232,N_14119,N_11395);
and U19233 (N_19233,N_12453,N_12598);
xnor U19234 (N_19234,N_13529,N_12366);
nand U19235 (N_19235,N_10620,N_10682);
or U19236 (N_19236,N_11274,N_14768);
and U19237 (N_19237,N_10530,N_14745);
or U19238 (N_19238,N_12902,N_14671);
or U19239 (N_19239,N_14085,N_14649);
xor U19240 (N_19240,N_11950,N_11966);
and U19241 (N_19241,N_12677,N_14342);
nand U19242 (N_19242,N_13993,N_13371);
or U19243 (N_19243,N_11996,N_14935);
or U19244 (N_19244,N_14185,N_12199);
or U19245 (N_19245,N_12026,N_10887);
nand U19246 (N_19246,N_10778,N_13607);
and U19247 (N_19247,N_10617,N_10892);
or U19248 (N_19248,N_12922,N_13054);
or U19249 (N_19249,N_14604,N_10005);
nand U19250 (N_19250,N_14015,N_10188);
nor U19251 (N_19251,N_13927,N_12427);
and U19252 (N_19252,N_12526,N_11674);
nand U19253 (N_19253,N_11982,N_11868);
and U19254 (N_19254,N_13331,N_11654);
nor U19255 (N_19255,N_10389,N_12234);
nor U19256 (N_19256,N_14473,N_10185);
nor U19257 (N_19257,N_13616,N_10233);
and U19258 (N_19258,N_10207,N_13185);
and U19259 (N_19259,N_12438,N_12264);
or U19260 (N_19260,N_14112,N_10580);
nor U19261 (N_19261,N_14636,N_10970);
xnor U19262 (N_19262,N_13810,N_14456);
and U19263 (N_19263,N_12930,N_14783);
xor U19264 (N_19264,N_11888,N_12789);
nor U19265 (N_19265,N_10202,N_10227);
nor U19266 (N_19266,N_11939,N_11446);
and U19267 (N_19267,N_11300,N_13307);
nor U19268 (N_19268,N_10550,N_10203);
nor U19269 (N_19269,N_12244,N_12371);
or U19270 (N_19270,N_11639,N_14630);
and U19271 (N_19271,N_11876,N_12299);
nor U19272 (N_19272,N_12235,N_11281);
and U19273 (N_19273,N_12306,N_10178);
nand U19274 (N_19274,N_14761,N_14161);
nand U19275 (N_19275,N_14787,N_12427);
or U19276 (N_19276,N_12251,N_11023);
nand U19277 (N_19277,N_10472,N_10325);
or U19278 (N_19278,N_10969,N_13534);
xnor U19279 (N_19279,N_14970,N_11987);
and U19280 (N_19280,N_10280,N_10461);
or U19281 (N_19281,N_12385,N_10799);
nand U19282 (N_19282,N_14169,N_11627);
or U19283 (N_19283,N_14320,N_12098);
nand U19284 (N_19284,N_13305,N_14680);
nand U19285 (N_19285,N_14214,N_12035);
nand U19286 (N_19286,N_14839,N_11388);
or U19287 (N_19287,N_10015,N_12698);
and U19288 (N_19288,N_12225,N_14390);
nand U19289 (N_19289,N_13408,N_13314);
nor U19290 (N_19290,N_14562,N_14710);
nor U19291 (N_19291,N_12851,N_12941);
or U19292 (N_19292,N_14692,N_11939);
nand U19293 (N_19293,N_12546,N_12358);
xnor U19294 (N_19294,N_10849,N_11875);
or U19295 (N_19295,N_11557,N_12029);
nand U19296 (N_19296,N_13456,N_10661);
nand U19297 (N_19297,N_12483,N_10375);
nor U19298 (N_19298,N_14787,N_11003);
and U19299 (N_19299,N_10867,N_10713);
nand U19300 (N_19300,N_12529,N_10679);
and U19301 (N_19301,N_11237,N_11161);
or U19302 (N_19302,N_14561,N_10297);
and U19303 (N_19303,N_13283,N_13574);
nand U19304 (N_19304,N_10114,N_13412);
or U19305 (N_19305,N_11478,N_10923);
and U19306 (N_19306,N_14310,N_12202);
nor U19307 (N_19307,N_11503,N_11429);
and U19308 (N_19308,N_11718,N_11948);
nand U19309 (N_19309,N_14226,N_10915);
nor U19310 (N_19310,N_13428,N_14782);
or U19311 (N_19311,N_13752,N_12064);
nand U19312 (N_19312,N_10181,N_11426);
nor U19313 (N_19313,N_12178,N_14033);
nand U19314 (N_19314,N_10899,N_14900);
or U19315 (N_19315,N_10457,N_14561);
or U19316 (N_19316,N_14075,N_14127);
nand U19317 (N_19317,N_11934,N_10435);
nand U19318 (N_19318,N_12362,N_11618);
nor U19319 (N_19319,N_13789,N_14952);
nand U19320 (N_19320,N_11049,N_11471);
nor U19321 (N_19321,N_12313,N_12146);
or U19322 (N_19322,N_11214,N_11220);
nand U19323 (N_19323,N_14211,N_10003);
nand U19324 (N_19324,N_12726,N_11894);
xor U19325 (N_19325,N_12707,N_12062);
xor U19326 (N_19326,N_10964,N_11912);
nand U19327 (N_19327,N_13026,N_12335);
and U19328 (N_19328,N_13021,N_14368);
nand U19329 (N_19329,N_10904,N_12008);
and U19330 (N_19330,N_10634,N_13824);
nand U19331 (N_19331,N_11578,N_12071);
nor U19332 (N_19332,N_13952,N_11254);
xnor U19333 (N_19333,N_13599,N_11104);
nor U19334 (N_19334,N_10559,N_14701);
and U19335 (N_19335,N_14575,N_13512);
nand U19336 (N_19336,N_14752,N_12252);
and U19337 (N_19337,N_12911,N_13716);
nor U19338 (N_19338,N_14919,N_10317);
nor U19339 (N_19339,N_10031,N_12708);
or U19340 (N_19340,N_13597,N_14378);
nor U19341 (N_19341,N_12174,N_12446);
and U19342 (N_19342,N_12783,N_10165);
or U19343 (N_19343,N_14400,N_13844);
or U19344 (N_19344,N_11629,N_11184);
and U19345 (N_19345,N_11533,N_10152);
or U19346 (N_19346,N_11828,N_13741);
and U19347 (N_19347,N_14951,N_12955);
nor U19348 (N_19348,N_11394,N_14096);
nand U19349 (N_19349,N_13388,N_11039);
nor U19350 (N_19350,N_14462,N_14312);
nor U19351 (N_19351,N_12727,N_13133);
or U19352 (N_19352,N_14977,N_13975);
and U19353 (N_19353,N_14735,N_10047);
and U19354 (N_19354,N_11931,N_14176);
nand U19355 (N_19355,N_10308,N_14438);
xor U19356 (N_19356,N_11701,N_13070);
nor U19357 (N_19357,N_13887,N_10383);
or U19358 (N_19358,N_12920,N_12606);
nand U19359 (N_19359,N_10581,N_11291);
nand U19360 (N_19360,N_10614,N_14889);
and U19361 (N_19361,N_11623,N_13628);
and U19362 (N_19362,N_10281,N_12630);
and U19363 (N_19363,N_12946,N_14992);
or U19364 (N_19364,N_11136,N_13288);
nand U19365 (N_19365,N_13138,N_12836);
or U19366 (N_19366,N_12436,N_13765);
or U19367 (N_19367,N_14355,N_11326);
or U19368 (N_19368,N_14820,N_14784);
and U19369 (N_19369,N_13506,N_13577);
nor U19370 (N_19370,N_13253,N_12571);
nor U19371 (N_19371,N_10149,N_14718);
nor U19372 (N_19372,N_12862,N_13229);
nor U19373 (N_19373,N_11910,N_14982);
nand U19374 (N_19374,N_10423,N_11917);
xnor U19375 (N_19375,N_14268,N_14325);
or U19376 (N_19376,N_14643,N_14044);
nor U19377 (N_19377,N_10867,N_11090);
nand U19378 (N_19378,N_12181,N_10924);
or U19379 (N_19379,N_10842,N_12522);
nand U19380 (N_19380,N_14570,N_13282);
and U19381 (N_19381,N_10955,N_12438);
nand U19382 (N_19382,N_11294,N_10620);
nand U19383 (N_19383,N_13042,N_13780);
nor U19384 (N_19384,N_13375,N_11163);
nand U19385 (N_19385,N_12988,N_13314);
and U19386 (N_19386,N_14188,N_13875);
nor U19387 (N_19387,N_13864,N_13979);
nor U19388 (N_19388,N_12785,N_13349);
or U19389 (N_19389,N_10222,N_10308);
nor U19390 (N_19390,N_14021,N_10207);
nand U19391 (N_19391,N_12484,N_10198);
nor U19392 (N_19392,N_10048,N_12295);
nor U19393 (N_19393,N_13968,N_11023);
nor U19394 (N_19394,N_11694,N_14354);
and U19395 (N_19395,N_12038,N_10295);
or U19396 (N_19396,N_12803,N_13197);
xor U19397 (N_19397,N_13921,N_11771);
and U19398 (N_19398,N_14174,N_13221);
or U19399 (N_19399,N_14077,N_14941);
nor U19400 (N_19400,N_14718,N_14159);
and U19401 (N_19401,N_13635,N_10118);
nor U19402 (N_19402,N_12680,N_14527);
nor U19403 (N_19403,N_11648,N_14155);
and U19404 (N_19404,N_11458,N_12573);
or U19405 (N_19405,N_11370,N_12007);
or U19406 (N_19406,N_13746,N_14010);
and U19407 (N_19407,N_10722,N_13101);
or U19408 (N_19408,N_14454,N_11692);
nand U19409 (N_19409,N_14321,N_12666);
nand U19410 (N_19410,N_14973,N_12256);
or U19411 (N_19411,N_14487,N_10050);
and U19412 (N_19412,N_11710,N_11913);
nor U19413 (N_19413,N_10368,N_11682);
nor U19414 (N_19414,N_10432,N_12641);
nand U19415 (N_19415,N_13059,N_14607);
nand U19416 (N_19416,N_14400,N_12787);
nand U19417 (N_19417,N_11014,N_13314);
or U19418 (N_19418,N_11021,N_14301);
nand U19419 (N_19419,N_10756,N_14699);
and U19420 (N_19420,N_11124,N_12063);
and U19421 (N_19421,N_13214,N_10847);
nand U19422 (N_19422,N_14681,N_10326);
nand U19423 (N_19423,N_12160,N_12247);
nand U19424 (N_19424,N_11024,N_13638);
nand U19425 (N_19425,N_12808,N_12969);
xor U19426 (N_19426,N_13165,N_14940);
or U19427 (N_19427,N_12248,N_14736);
nand U19428 (N_19428,N_14659,N_14353);
nor U19429 (N_19429,N_11918,N_14558);
nor U19430 (N_19430,N_13140,N_13138);
nand U19431 (N_19431,N_12832,N_11180);
and U19432 (N_19432,N_14736,N_11968);
nor U19433 (N_19433,N_14785,N_14624);
nand U19434 (N_19434,N_13855,N_12965);
or U19435 (N_19435,N_11381,N_14300);
and U19436 (N_19436,N_10086,N_14707);
nor U19437 (N_19437,N_14905,N_12802);
or U19438 (N_19438,N_10804,N_14415);
nand U19439 (N_19439,N_11483,N_13681);
nor U19440 (N_19440,N_12545,N_11588);
nor U19441 (N_19441,N_13159,N_10617);
xnor U19442 (N_19442,N_13982,N_10236);
nand U19443 (N_19443,N_13130,N_10392);
and U19444 (N_19444,N_11808,N_14748);
or U19445 (N_19445,N_14097,N_14862);
or U19446 (N_19446,N_11364,N_14290);
nor U19447 (N_19447,N_10470,N_11509);
nor U19448 (N_19448,N_11883,N_10886);
nor U19449 (N_19449,N_12054,N_13062);
or U19450 (N_19450,N_13333,N_12853);
nand U19451 (N_19451,N_12562,N_13483);
nand U19452 (N_19452,N_11952,N_12814);
and U19453 (N_19453,N_14560,N_14532);
nor U19454 (N_19454,N_14874,N_13128);
and U19455 (N_19455,N_12236,N_10276);
nand U19456 (N_19456,N_10466,N_13267);
nor U19457 (N_19457,N_14066,N_11642);
nand U19458 (N_19458,N_12063,N_12669);
or U19459 (N_19459,N_14019,N_13702);
and U19460 (N_19460,N_10910,N_11684);
nor U19461 (N_19461,N_13488,N_14099);
nor U19462 (N_19462,N_11710,N_14852);
or U19463 (N_19463,N_12638,N_10448);
or U19464 (N_19464,N_13491,N_14089);
nand U19465 (N_19465,N_10909,N_10611);
and U19466 (N_19466,N_14283,N_14767);
xor U19467 (N_19467,N_13579,N_13866);
and U19468 (N_19468,N_13464,N_11411);
nand U19469 (N_19469,N_11624,N_14313);
nor U19470 (N_19470,N_11997,N_10267);
nor U19471 (N_19471,N_10954,N_10827);
nor U19472 (N_19472,N_11691,N_13593);
and U19473 (N_19473,N_11988,N_10507);
or U19474 (N_19474,N_11122,N_14545);
nor U19475 (N_19475,N_12962,N_14989);
and U19476 (N_19476,N_10341,N_14431);
nand U19477 (N_19477,N_13253,N_10419);
nand U19478 (N_19478,N_13222,N_12346);
or U19479 (N_19479,N_14975,N_13093);
nor U19480 (N_19480,N_10958,N_11014);
nor U19481 (N_19481,N_12183,N_13175);
and U19482 (N_19482,N_10569,N_12691);
nand U19483 (N_19483,N_12401,N_12526);
and U19484 (N_19484,N_14081,N_10506);
and U19485 (N_19485,N_10968,N_11485);
nor U19486 (N_19486,N_10817,N_13819);
nand U19487 (N_19487,N_13213,N_10472);
and U19488 (N_19488,N_11617,N_12684);
or U19489 (N_19489,N_11619,N_11404);
nand U19490 (N_19490,N_11319,N_14203);
or U19491 (N_19491,N_13155,N_13436);
and U19492 (N_19492,N_11001,N_13361);
or U19493 (N_19493,N_10036,N_10552);
nor U19494 (N_19494,N_10072,N_11448);
nand U19495 (N_19495,N_12444,N_12852);
or U19496 (N_19496,N_10063,N_11392);
and U19497 (N_19497,N_10270,N_12672);
nor U19498 (N_19498,N_14720,N_10552);
nor U19499 (N_19499,N_12427,N_14995);
nor U19500 (N_19500,N_10531,N_10898);
and U19501 (N_19501,N_10920,N_13881);
nor U19502 (N_19502,N_11334,N_10461);
nand U19503 (N_19503,N_13092,N_12541);
or U19504 (N_19504,N_14312,N_10656);
or U19505 (N_19505,N_10149,N_12930);
nor U19506 (N_19506,N_12234,N_11641);
and U19507 (N_19507,N_10815,N_11403);
xor U19508 (N_19508,N_13282,N_14441);
or U19509 (N_19509,N_14139,N_14301);
nand U19510 (N_19510,N_12320,N_14586);
nor U19511 (N_19511,N_12270,N_13364);
and U19512 (N_19512,N_11937,N_13715);
and U19513 (N_19513,N_11774,N_10412);
nor U19514 (N_19514,N_10782,N_11219);
xor U19515 (N_19515,N_12943,N_14464);
or U19516 (N_19516,N_11169,N_13186);
nand U19517 (N_19517,N_11951,N_13818);
or U19518 (N_19518,N_11380,N_11217);
or U19519 (N_19519,N_13847,N_14229);
or U19520 (N_19520,N_10262,N_14066);
or U19521 (N_19521,N_13902,N_14165);
nor U19522 (N_19522,N_12154,N_13158);
or U19523 (N_19523,N_10041,N_12483);
and U19524 (N_19524,N_14298,N_11725);
or U19525 (N_19525,N_11233,N_14292);
and U19526 (N_19526,N_12659,N_10468);
nor U19527 (N_19527,N_13026,N_12210);
nor U19528 (N_19528,N_11918,N_14779);
nand U19529 (N_19529,N_13141,N_11496);
or U19530 (N_19530,N_13866,N_13617);
nor U19531 (N_19531,N_13340,N_13356);
or U19532 (N_19532,N_12075,N_10072);
nand U19533 (N_19533,N_13773,N_10341);
nor U19534 (N_19534,N_12651,N_10575);
nor U19535 (N_19535,N_10848,N_12556);
and U19536 (N_19536,N_14134,N_12340);
or U19537 (N_19537,N_12609,N_11415);
or U19538 (N_19538,N_12184,N_14328);
and U19539 (N_19539,N_13169,N_10233);
nor U19540 (N_19540,N_14071,N_13694);
nor U19541 (N_19541,N_10211,N_11678);
nand U19542 (N_19542,N_10622,N_10981);
or U19543 (N_19543,N_12074,N_12167);
or U19544 (N_19544,N_13818,N_12624);
or U19545 (N_19545,N_11114,N_13638);
nand U19546 (N_19546,N_12250,N_13273);
nand U19547 (N_19547,N_11688,N_11179);
and U19548 (N_19548,N_10424,N_14833);
nand U19549 (N_19549,N_11801,N_10704);
nor U19550 (N_19550,N_14408,N_13810);
or U19551 (N_19551,N_12298,N_10976);
nor U19552 (N_19552,N_12104,N_11173);
and U19553 (N_19553,N_12190,N_13234);
nand U19554 (N_19554,N_13352,N_11403);
nand U19555 (N_19555,N_13678,N_10188);
nand U19556 (N_19556,N_11364,N_10198);
or U19557 (N_19557,N_11498,N_12882);
nor U19558 (N_19558,N_14026,N_13908);
nor U19559 (N_19559,N_10479,N_13382);
and U19560 (N_19560,N_10462,N_12652);
or U19561 (N_19561,N_13895,N_14541);
and U19562 (N_19562,N_12075,N_14852);
and U19563 (N_19563,N_11006,N_13149);
and U19564 (N_19564,N_12658,N_13288);
nor U19565 (N_19565,N_14410,N_14153);
and U19566 (N_19566,N_13194,N_12246);
and U19567 (N_19567,N_12579,N_14423);
nor U19568 (N_19568,N_13096,N_14963);
nor U19569 (N_19569,N_12036,N_12893);
or U19570 (N_19570,N_14525,N_11357);
nand U19571 (N_19571,N_13696,N_14081);
nor U19572 (N_19572,N_14155,N_13127);
nor U19573 (N_19573,N_10011,N_11698);
nor U19574 (N_19574,N_10230,N_13761);
or U19575 (N_19575,N_14883,N_14908);
or U19576 (N_19576,N_12293,N_13042);
nor U19577 (N_19577,N_13316,N_13507);
or U19578 (N_19578,N_10931,N_10879);
nor U19579 (N_19579,N_14550,N_11437);
nor U19580 (N_19580,N_10898,N_11911);
nor U19581 (N_19581,N_12973,N_14297);
or U19582 (N_19582,N_13860,N_12265);
or U19583 (N_19583,N_14213,N_13645);
and U19584 (N_19584,N_13119,N_11397);
nor U19585 (N_19585,N_13304,N_14224);
nor U19586 (N_19586,N_11056,N_13578);
nor U19587 (N_19587,N_12889,N_11115);
or U19588 (N_19588,N_14846,N_11166);
and U19589 (N_19589,N_13685,N_13962);
nand U19590 (N_19590,N_14429,N_14431);
nor U19591 (N_19591,N_14710,N_12301);
nand U19592 (N_19592,N_13023,N_14282);
or U19593 (N_19593,N_12529,N_10862);
nand U19594 (N_19594,N_11252,N_11247);
nor U19595 (N_19595,N_11483,N_11938);
and U19596 (N_19596,N_12136,N_12127);
and U19597 (N_19597,N_11183,N_11788);
nand U19598 (N_19598,N_10469,N_14943);
and U19599 (N_19599,N_13159,N_14338);
nor U19600 (N_19600,N_11434,N_12420);
and U19601 (N_19601,N_11077,N_12121);
or U19602 (N_19602,N_12129,N_10880);
nor U19603 (N_19603,N_12050,N_12260);
and U19604 (N_19604,N_11522,N_11610);
and U19605 (N_19605,N_10872,N_11804);
or U19606 (N_19606,N_14169,N_11836);
or U19607 (N_19607,N_12397,N_14459);
nand U19608 (N_19608,N_14638,N_12942);
nand U19609 (N_19609,N_11562,N_13568);
nor U19610 (N_19610,N_11569,N_14871);
or U19611 (N_19611,N_11157,N_10875);
and U19612 (N_19612,N_14667,N_10824);
nand U19613 (N_19613,N_10477,N_12386);
nand U19614 (N_19614,N_13502,N_13967);
nand U19615 (N_19615,N_11074,N_13295);
nor U19616 (N_19616,N_14458,N_10831);
nor U19617 (N_19617,N_12976,N_14306);
or U19618 (N_19618,N_13384,N_13753);
or U19619 (N_19619,N_11292,N_12258);
and U19620 (N_19620,N_13507,N_14577);
nand U19621 (N_19621,N_12363,N_10780);
nand U19622 (N_19622,N_14019,N_11311);
nand U19623 (N_19623,N_12436,N_14773);
or U19624 (N_19624,N_14015,N_13617);
nand U19625 (N_19625,N_13016,N_10197);
nor U19626 (N_19626,N_11893,N_11060);
or U19627 (N_19627,N_12114,N_14525);
nor U19628 (N_19628,N_12626,N_10693);
nand U19629 (N_19629,N_12323,N_11044);
nand U19630 (N_19630,N_14818,N_13216);
and U19631 (N_19631,N_11533,N_12839);
or U19632 (N_19632,N_10332,N_14235);
and U19633 (N_19633,N_14590,N_12365);
or U19634 (N_19634,N_13700,N_13765);
and U19635 (N_19635,N_11411,N_10822);
or U19636 (N_19636,N_13683,N_10651);
and U19637 (N_19637,N_12203,N_13161);
or U19638 (N_19638,N_10075,N_11438);
xor U19639 (N_19639,N_10727,N_12365);
nor U19640 (N_19640,N_13706,N_13783);
nor U19641 (N_19641,N_14498,N_14047);
or U19642 (N_19642,N_13783,N_12369);
or U19643 (N_19643,N_11731,N_12969);
or U19644 (N_19644,N_12833,N_10916);
or U19645 (N_19645,N_11207,N_13791);
nor U19646 (N_19646,N_14190,N_11251);
nor U19647 (N_19647,N_14104,N_10991);
and U19648 (N_19648,N_10783,N_10571);
or U19649 (N_19649,N_10402,N_12739);
nand U19650 (N_19650,N_10343,N_11323);
xor U19651 (N_19651,N_14500,N_14539);
or U19652 (N_19652,N_11998,N_12098);
and U19653 (N_19653,N_12344,N_13729);
or U19654 (N_19654,N_13168,N_13512);
nand U19655 (N_19655,N_10832,N_10119);
nor U19656 (N_19656,N_10183,N_12445);
or U19657 (N_19657,N_14362,N_11576);
nand U19658 (N_19658,N_13889,N_10986);
nor U19659 (N_19659,N_11974,N_13205);
and U19660 (N_19660,N_10741,N_11511);
nor U19661 (N_19661,N_12764,N_12546);
and U19662 (N_19662,N_13461,N_10212);
nand U19663 (N_19663,N_11787,N_10528);
or U19664 (N_19664,N_14085,N_10274);
nor U19665 (N_19665,N_12411,N_12688);
nand U19666 (N_19666,N_10573,N_11037);
nor U19667 (N_19667,N_12552,N_12647);
or U19668 (N_19668,N_13693,N_14817);
nand U19669 (N_19669,N_10518,N_14405);
or U19670 (N_19670,N_12611,N_14552);
nor U19671 (N_19671,N_10687,N_11967);
nand U19672 (N_19672,N_10951,N_14004);
and U19673 (N_19673,N_10209,N_10850);
and U19674 (N_19674,N_14120,N_12746);
nand U19675 (N_19675,N_13344,N_14889);
nor U19676 (N_19676,N_10032,N_12819);
nor U19677 (N_19677,N_13851,N_10383);
nand U19678 (N_19678,N_10718,N_10263);
nand U19679 (N_19679,N_14062,N_13879);
or U19680 (N_19680,N_11950,N_12712);
nand U19681 (N_19681,N_12625,N_11893);
nand U19682 (N_19682,N_11234,N_13820);
nor U19683 (N_19683,N_14471,N_11868);
and U19684 (N_19684,N_13776,N_10198);
or U19685 (N_19685,N_10669,N_14429);
nor U19686 (N_19686,N_14004,N_10884);
or U19687 (N_19687,N_14748,N_10184);
nand U19688 (N_19688,N_13170,N_14859);
nand U19689 (N_19689,N_10458,N_11412);
or U19690 (N_19690,N_11132,N_11701);
nand U19691 (N_19691,N_13898,N_12175);
or U19692 (N_19692,N_13373,N_10934);
nand U19693 (N_19693,N_14625,N_13360);
xnor U19694 (N_19694,N_13606,N_10553);
nand U19695 (N_19695,N_14789,N_11034);
and U19696 (N_19696,N_13904,N_10097);
nor U19697 (N_19697,N_13600,N_11549);
or U19698 (N_19698,N_11298,N_13029);
nor U19699 (N_19699,N_13198,N_14169);
and U19700 (N_19700,N_11545,N_14706);
or U19701 (N_19701,N_10454,N_10178);
and U19702 (N_19702,N_13599,N_13116);
and U19703 (N_19703,N_13896,N_12421);
or U19704 (N_19704,N_14021,N_11817);
nor U19705 (N_19705,N_13489,N_13487);
or U19706 (N_19706,N_14541,N_10278);
nor U19707 (N_19707,N_10196,N_13195);
nor U19708 (N_19708,N_10152,N_10442);
nor U19709 (N_19709,N_11764,N_11412);
and U19710 (N_19710,N_11206,N_12833);
xor U19711 (N_19711,N_11189,N_11914);
nand U19712 (N_19712,N_13249,N_12213);
and U19713 (N_19713,N_10641,N_10673);
and U19714 (N_19714,N_11801,N_12790);
nand U19715 (N_19715,N_10475,N_12897);
nor U19716 (N_19716,N_14085,N_13581);
or U19717 (N_19717,N_12649,N_13399);
nor U19718 (N_19718,N_10644,N_13160);
or U19719 (N_19719,N_11816,N_12355);
nand U19720 (N_19720,N_11756,N_11850);
and U19721 (N_19721,N_10916,N_14665);
and U19722 (N_19722,N_12270,N_14871);
nor U19723 (N_19723,N_10761,N_11056);
and U19724 (N_19724,N_12532,N_11148);
or U19725 (N_19725,N_11434,N_12212);
nor U19726 (N_19726,N_12246,N_10971);
or U19727 (N_19727,N_10412,N_10528);
nand U19728 (N_19728,N_14446,N_13233);
and U19729 (N_19729,N_10395,N_10656);
or U19730 (N_19730,N_12024,N_10391);
and U19731 (N_19731,N_12637,N_12227);
nor U19732 (N_19732,N_14767,N_13792);
and U19733 (N_19733,N_14491,N_12632);
or U19734 (N_19734,N_11603,N_11227);
and U19735 (N_19735,N_13919,N_10757);
and U19736 (N_19736,N_13046,N_14128);
nand U19737 (N_19737,N_13450,N_11356);
or U19738 (N_19738,N_14898,N_11574);
nand U19739 (N_19739,N_12164,N_12217);
or U19740 (N_19740,N_10915,N_14514);
or U19741 (N_19741,N_10082,N_11968);
or U19742 (N_19742,N_11906,N_13603);
nor U19743 (N_19743,N_10703,N_14697);
nor U19744 (N_19744,N_13446,N_14367);
and U19745 (N_19745,N_10697,N_13785);
nand U19746 (N_19746,N_14068,N_14297);
nand U19747 (N_19747,N_10183,N_12743);
and U19748 (N_19748,N_11431,N_12587);
and U19749 (N_19749,N_13710,N_14486);
nand U19750 (N_19750,N_10649,N_11722);
nor U19751 (N_19751,N_10367,N_14370);
and U19752 (N_19752,N_11409,N_14428);
and U19753 (N_19753,N_10744,N_11523);
nand U19754 (N_19754,N_14835,N_14251);
or U19755 (N_19755,N_11732,N_12291);
or U19756 (N_19756,N_14269,N_11426);
nor U19757 (N_19757,N_14254,N_12335);
or U19758 (N_19758,N_11956,N_13519);
nand U19759 (N_19759,N_10911,N_12982);
nand U19760 (N_19760,N_11379,N_13451);
nand U19761 (N_19761,N_13537,N_13279);
nor U19762 (N_19762,N_13201,N_13017);
or U19763 (N_19763,N_11532,N_10238);
nor U19764 (N_19764,N_11913,N_12993);
and U19765 (N_19765,N_13240,N_10418);
xor U19766 (N_19766,N_13218,N_14007);
nor U19767 (N_19767,N_12398,N_12914);
nand U19768 (N_19768,N_11304,N_10955);
and U19769 (N_19769,N_12200,N_13574);
nand U19770 (N_19770,N_13250,N_10128);
nor U19771 (N_19771,N_11037,N_13236);
or U19772 (N_19772,N_11835,N_14037);
nand U19773 (N_19773,N_12550,N_10202);
or U19774 (N_19774,N_12174,N_13512);
and U19775 (N_19775,N_14122,N_11679);
or U19776 (N_19776,N_14323,N_14232);
nor U19777 (N_19777,N_10124,N_10484);
nand U19778 (N_19778,N_12733,N_10286);
or U19779 (N_19779,N_10898,N_12816);
and U19780 (N_19780,N_11370,N_12763);
and U19781 (N_19781,N_12858,N_11055);
and U19782 (N_19782,N_11670,N_11224);
nand U19783 (N_19783,N_14255,N_12114);
or U19784 (N_19784,N_12368,N_11932);
nor U19785 (N_19785,N_14592,N_11141);
nand U19786 (N_19786,N_13067,N_14020);
nand U19787 (N_19787,N_13147,N_13519);
and U19788 (N_19788,N_11387,N_10479);
nor U19789 (N_19789,N_11125,N_13834);
nor U19790 (N_19790,N_11241,N_12717);
or U19791 (N_19791,N_12308,N_13327);
nor U19792 (N_19792,N_13159,N_14044);
nor U19793 (N_19793,N_11327,N_14713);
nand U19794 (N_19794,N_12233,N_12263);
or U19795 (N_19795,N_10359,N_12910);
or U19796 (N_19796,N_10230,N_10120);
nor U19797 (N_19797,N_14196,N_10604);
and U19798 (N_19798,N_14159,N_11938);
and U19799 (N_19799,N_14953,N_10228);
nand U19800 (N_19800,N_12642,N_11851);
nand U19801 (N_19801,N_10809,N_11928);
nand U19802 (N_19802,N_11016,N_11628);
nor U19803 (N_19803,N_12077,N_11533);
nor U19804 (N_19804,N_11088,N_13241);
nand U19805 (N_19805,N_12904,N_11932);
nor U19806 (N_19806,N_11914,N_10888);
nand U19807 (N_19807,N_10880,N_14823);
nand U19808 (N_19808,N_10337,N_11201);
and U19809 (N_19809,N_10463,N_12439);
and U19810 (N_19810,N_10295,N_10766);
nand U19811 (N_19811,N_10542,N_13679);
or U19812 (N_19812,N_12129,N_13443);
nand U19813 (N_19813,N_14464,N_11222);
nand U19814 (N_19814,N_10159,N_10803);
nand U19815 (N_19815,N_13057,N_10384);
or U19816 (N_19816,N_13835,N_12278);
nor U19817 (N_19817,N_10846,N_14116);
and U19818 (N_19818,N_14999,N_14420);
nand U19819 (N_19819,N_11496,N_12719);
or U19820 (N_19820,N_11539,N_10557);
or U19821 (N_19821,N_12107,N_13146);
nand U19822 (N_19822,N_11718,N_11473);
nor U19823 (N_19823,N_14496,N_11924);
and U19824 (N_19824,N_13148,N_13151);
xor U19825 (N_19825,N_10475,N_10114);
and U19826 (N_19826,N_12997,N_12031);
or U19827 (N_19827,N_13647,N_10477);
nor U19828 (N_19828,N_11860,N_14009);
nand U19829 (N_19829,N_14250,N_11130);
nor U19830 (N_19830,N_10114,N_11112);
nand U19831 (N_19831,N_10947,N_14858);
nand U19832 (N_19832,N_14498,N_12528);
or U19833 (N_19833,N_10020,N_10258);
nand U19834 (N_19834,N_11017,N_13700);
nand U19835 (N_19835,N_12021,N_14727);
nor U19836 (N_19836,N_14493,N_10904);
and U19837 (N_19837,N_14772,N_14357);
nand U19838 (N_19838,N_12480,N_12295);
nand U19839 (N_19839,N_12808,N_14511);
nor U19840 (N_19840,N_11846,N_14944);
nand U19841 (N_19841,N_14831,N_11971);
or U19842 (N_19842,N_10824,N_12938);
nor U19843 (N_19843,N_12751,N_11182);
nor U19844 (N_19844,N_10932,N_14163);
and U19845 (N_19845,N_13334,N_10406);
nor U19846 (N_19846,N_12124,N_10456);
nand U19847 (N_19847,N_13587,N_11075);
nor U19848 (N_19848,N_11534,N_10517);
or U19849 (N_19849,N_13729,N_11995);
and U19850 (N_19850,N_13641,N_12102);
or U19851 (N_19851,N_12296,N_12589);
nor U19852 (N_19852,N_13015,N_12717);
and U19853 (N_19853,N_11057,N_12239);
nand U19854 (N_19854,N_14478,N_13058);
nand U19855 (N_19855,N_11749,N_14695);
nand U19856 (N_19856,N_13127,N_12177);
or U19857 (N_19857,N_12559,N_11264);
nand U19858 (N_19858,N_13849,N_12464);
and U19859 (N_19859,N_11204,N_12512);
nand U19860 (N_19860,N_11227,N_12473);
and U19861 (N_19861,N_12124,N_14997);
nand U19862 (N_19862,N_12897,N_12058);
or U19863 (N_19863,N_14070,N_14418);
nand U19864 (N_19864,N_14523,N_11731);
nand U19865 (N_19865,N_11215,N_11384);
and U19866 (N_19866,N_13863,N_10679);
and U19867 (N_19867,N_10455,N_14856);
and U19868 (N_19868,N_13957,N_10735);
or U19869 (N_19869,N_12541,N_11265);
and U19870 (N_19870,N_14189,N_14731);
nand U19871 (N_19871,N_11819,N_12147);
nor U19872 (N_19872,N_11829,N_11855);
nor U19873 (N_19873,N_11995,N_13503);
nand U19874 (N_19874,N_14731,N_12332);
nor U19875 (N_19875,N_11935,N_10985);
nand U19876 (N_19876,N_13173,N_11113);
nor U19877 (N_19877,N_13714,N_13472);
nor U19878 (N_19878,N_13922,N_11673);
nand U19879 (N_19879,N_10670,N_10878);
nor U19880 (N_19880,N_10247,N_12416);
nor U19881 (N_19881,N_12697,N_12110);
and U19882 (N_19882,N_12414,N_13214);
nand U19883 (N_19883,N_13519,N_10177);
nor U19884 (N_19884,N_10963,N_14862);
nor U19885 (N_19885,N_10085,N_10500);
or U19886 (N_19886,N_11948,N_13426);
nor U19887 (N_19887,N_11432,N_11661);
nand U19888 (N_19888,N_12201,N_13071);
and U19889 (N_19889,N_13423,N_14563);
xor U19890 (N_19890,N_10025,N_14902);
nand U19891 (N_19891,N_12189,N_13241);
nor U19892 (N_19892,N_10145,N_10072);
nand U19893 (N_19893,N_11085,N_10022);
nor U19894 (N_19894,N_12493,N_12054);
xor U19895 (N_19895,N_14053,N_13112);
nand U19896 (N_19896,N_11195,N_11392);
nor U19897 (N_19897,N_13333,N_12667);
nand U19898 (N_19898,N_10446,N_12967);
and U19899 (N_19899,N_13067,N_13745);
and U19900 (N_19900,N_12594,N_13596);
nor U19901 (N_19901,N_12021,N_11091);
nor U19902 (N_19902,N_14500,N_11282);
nor U19903 (N_19903,N_13779,N_14273);
or U19904 (N_19904,N_13466,N_11596);
nand U19905 (N_19905,N_10141,N_10890);
or U19906 (N_19906,N_11280,N_11286);
and U19907 (N_19907,N_11951,N_11652);
nor U19908 (N_19908,N_13741,N_11736);
or U19909 (N_19909,N_12348,N_13459);
or U19910 (N_19910,N_12679,N_12665);
and U19911 (N_19911,N_11043,N_14770);
nand U19912 (N_19912,N_11311,N_12318);
nand U19913 (N_19913,N_10059,N_14395);
and U19914 (N_19914,N_11005,N_12456);
and U19915 (N_19915,N_10824,N_13417);
nor U19916 (N_19916,N_12869,N_13982);
nand U19917 (N_19917,N_10062,N_10328);
nor U19918 (N_19918,N_14321,N_14920);
nand U19919 (N_19919,N_13118,N_11989);
nor U19920 (N_19920,N_13084,N_14098);
nor U19921 (N_19921,N_12019,N_11232);
and U19922 (N_19922,N_12709,N_14826);
or U19923 (N_19923,N_10216,N_11502);
and U19924 (N_19924,N_14225,N_14251);
or U19925 (N_19925,N_11296,N_12891);
nor U19926 (N_19926,N_13454,N_10221);
nand U19927 (N_19927,N_10629,N_10005);
or U19928 (N_19928,N_11493,N_14776);
nand U19929 (N_19929,N_13550,N_10314);
and U19930 (N_19930,N_10642,N_12246);
nor U19931 (N_19931,N_14775,N_14159);
nor U19932 (N_19932,N_13438,N_10800);
or U19933 (N_19933,N_14290,N_11605);
or U19934 (N_19934,N_11054,N_11505);
or U19935 (N_19935,N_13571,N_11111);
or U19936 (N_19936,N_10374,N_14255);
and U19937 (N_19937,N_13910,N_14104);
or U19938 (N_19938,N_12036,N_10671);
nor U19939 (N_19939,N_11405,N_13476);
nor U19940 (N_19940,N_12890,N_11153);
nand U19941 (N_19941,N_14121,N_11687);
or U19942 (N_19942,N_12187,N_10951);
nor U19943 (N_19943,N_14938,N_14941);
and U19944 (N_19944,N_12859,N_13543);
and U19945 (N_19945,N_11063,N_11747);
nand U19946 (N_19946,N_13470,N_10876);
nor U19947 (N_19947,N_14661,N_12329);
nor U19948 (N_19948,N_14940,N_14641);
or U19949 (N_19949,N_10570,N_14831);
nand U19950 (N_19950,N_12433,N_13431);
nor U19951 (N_19951,N_13658,N_11389);
or U19952 (N_19952,N_13581,N_11264);
or U19953 (N_19953,N_10438,N_10896);
or U19954 (N_19954,N_11971,N_11423);
or U19955 (N_19955,N_12930,N_14985);
nor U19956 (N_19956,N_11374,N_12722);
nor U19957 (N_19957,N_12623,N_12779);
nor U19958 (N_19958,N_13518,N_10007);
nand U19959 (N_19959,N_14855,N_14810);
or U19960 (N_19960,N_10312,N_10405);
nand U19961 (N_19961,N_14251,N_11135);
nand U19962 (N_19962,N_12682,N_12365);
xnor U19963 (N_19963,N_12119,N_11253);
nor U19964 (N_19964,N_13127,N_14630);
and U19965 (N_19965,N_13329,N_12678);
nor U19966 (N_19966,N_12415,N_12008);
and U19967 (N_19967,N_13777,N_10636);
or U19968 (N_19968,N_13442,N_11351);
or U19969 (N_19969,N_14826,N_11230);
nand U19970 (N_19970,N_10087,N_11342);
and U19971 (N_19971,N_10763,N_12657);
or U19972 (N_19972,N_10626,N_12011);
or U19973 (N_19973,N_11941,N_12271);
nor U19974 (N_19974,N_10067,N_13495);
nand U19975 (N_19975,N_11904,N_12550);
and U19976 (N_19976,N_12735,N_10314);
nand U19977 (N_19977,N_11143,N_12577);
xnor U19978 (N_19978,N_13541,N_11321);
and U19979 (N_19979,N_14165,N_14062);
and U19980 (N_19980,N_10009,N_13022);
or U19981 (N_19981,N_13729,N_11761);
and U19982 (N_19982,N_14841,N_11064);
and U19983 (N_19983,N_12722,N_13300);
or U19984 (N_19984,N_13981,N_11534);
and U19985 (N_19985,N_10862,N_10511);
and U19986 (N_19986,N_13377,N_13919);
or U19987 (N_19987,N_11404,N_13799);
xnor U19988 (N_19988,N_13417,N_11374);
or U19989 (N_19989,N_12796,N_11948);
and U19990 (N_19990,N_11195,N_12059);
or U19991 (N_19991,N_14344,N_10579);
and U19992 (N_19992,N_10393,N_13117);
xor U19993 (N_19993,N_13866,N_10686);
nand U19994 (N_19994,N_11360,N_14329);
nand U19995 (N_19995,N_10084,N_10457);
or U19996 (N_19996,N_14410,N_11310);
nand U19997 (N_19997,N_14069,N_12027);
nor U19998 (N_19998,N_11412,N_11008);
xor U19999 (N_19999,N_11095,N_13918);
nand UO_0 (O_0,N_17979,N_17020);
nand UO_1 (O_1,N_17490,N_18712);
or UO_2 (O_2,N_15773,N_17242);
nor UO_3 (O_3,N_19424,N_15251);
or UO_4 (O_4,N_15245,N_17489);
nor UO_5 (O_5,N_18729,N_17905);
or UO_6 (O_6,N_15350,N_16400);
xnor UO_7 (O_7,N_19959,N_18796);
nor UO_8 (O_8,N_15386,N_17740);
nand UO_9 (O_9,N_17478,N_19930);
nand UO_10 (O_10,N_18091,N_17361);
nor UO_11 (O_11,N_17147,N_18614);
nand UO_12 (O_12,N_15624,N_17276);
nand UO_13 (O_13,N_19301,N_17501);
or UO_14 (O_14,N_15201,N_17323);
nor UO_15 (O_15,N_16052,N_19974);
xor UO_16 (O_16,N_18871,N_19780);
nand UO_17 (O_17,N_16957,N_15105);
and UO_18 (O_18,N_18173,N_18792);
or UO_19 (O_19,N_15462,N_18211);
nor UO_20 (O_20,N_19793,N_16197);
and UO_21 (O_21,N_17707,N_18361);
nand UO_22 (O_22,N_16723,N_16256);
and UO_23 (O_23,N_16598,N_17856);
nor UO_24 (O_24,N_19988,N_17952);
nand UO_25 (O_25,N_17082,N_17860);
xor UO_26 (O_26,N_18937,N_18772);
and UO_27 (O_27,N_19734,N_16394);
nor UO_28 (O_28,N_16322,N_17434);
or UO_29 (O_29,N_15067,N_15921);
nand UO_30 (O_30,N_17731,N_17822);
nor UO_31 (O_31,N_18856,N_17817);
and UO_32 (O_32,N_17439,N_19513);
and UO_33 (O_33,N_18543,N_18390);
nand UO_34 (O_34,N_19772,N_18953);
nor UO_35 (O_35,N_16129,N_19716);
or UO_36 (O_36,N_15411,N_16631);
or UO_37 (O_37,N_19078,N_17304);
nand UO_38 (O_38,N_18059,N_15015);
and UO_39 (O_39,N_15709,N_18236);
or UO_40 (O_40,N_17787,N_15284);
and UO_41 (O_41,N_17330,N_16128);
or UO_42 (O_42,N_17638,N_15515);
nor UO_43 (O_43,N_17256,N_16318);
xnor UO_44 (O_44,N_18031,N_16717);
and UO_45 (O_45,N_16618,N_16564);
nand UO_46 (O_46,N_19564,N_19099);
and UO_47 (O_47,N_19444,N_18261);
nand UO_48 (O_48,N_17072,N_18174);
or UO_49 (O_49,N_15333,N_17032);
and UO_50 (O_50,N_16011,N_17764);
nand UO_51 (O_51,N_17680,N_15871);
or UO_52 (O_52,N_15638,N_16445);
or UO_53 (O_53,N_17840,N_15435);
and UO_54 (O_54,N_19139,N_16758);
or UO_55 (O_55,N_15394,N_16730);
nor UO_56 (O_56,N_19536,N_16436);
and UO_57 (O_57,N_15780,N_18528);
or UO_58 (O_58,N_18355,N_18582);
nand UO_59 (O_59,N_18363,N_15484);
or UO_60 (O_60,N_16440,N_18298);
and UO_61 (O_61,N_15948,N_16025);
or UO_62 (O_62,N_17073,N_15879);
nand UO_63 (O_63,N_17423,N_17228);
nand UO_64 (O_64,N_15819,N_16625);
and UO_65 (O_65,N_16022,N_17530);
or UO_66 (O_66,N_19830,N_18897);
and UO_67 (O_67,N_16677,N_17108);
and UO_68 (O_68,N_16066,N_16845);
and UO_69 (O_69,N_18012,N_15905);
and UO_70 (O_70,N_19459,N_16594);
nor UO_71 (O_71,N_17296,N_16107);
or UO_72 (O_72,N_15226,N_17468);
or UO_73 (O_73,N_18379,N_17332);
nor UO_74 (O_74,N_17404,N_19533);
or UO_75 (O_75,N_15177,N_16049);
nand UO_76 (O_76,N_18376,N_19198);
and UO_77 (O_77,N_17949,N_16497);
nor UO_78 (O_78,N_18967,N_18210);
nor UO_79 (O_79,N_15283,N_18748);
nand UO_80 (O_80,N_19377,N_18891);
nand UO_81 (O_81,N_17966,N_19895);
nand UO_82 (O_82,N_15485,N_16061);
or UO_83 (O_83,N_15764,N_18693);
nand UO_84 (O_84,N_17903,N_19876);
or UO_85 (O_85,N_16888,N_18997);
xnor UO_86 (O_86,N_15397,N_16471);
nor UO_87 (O_87,N_16691,N_15393);
nand UO_88 (O_88,N_19381,N_15282);
nor UO_89 (O_89,N_16161,N_19719);
nand UO_90 (O_90,N_19640,N_18027);
and UO_91 (O_91,N_18787,N_16282);
nand UO_92 (O_92,N_17174,N_18654);
and UO_93 (O_93,N_18512,N_18542);
nand UO_94 (O_94,N_19018,N_15606);
nor UO_95 (O_95,N_15334,N_15714);
nand UO_96 (O_96,N_18500,N_16600);
or UO_97 (O_97,N_19315,N_15431);
or UO_98 (O_98,N_18392,N_15957);
and UO_99 (O_99,N_16513,N_16079);
nor UO_100 (O_100,N_19567,N_17533);
nand UO_101 (O_101,N_15254,N_19909);
xor UO_102 (O_102,N_17114,N_16818);
and UO_103 (O_103,N_15155,N_18521);
nor UO_104 (O_104,N_19217,N_17570);
nor UO_105 (O_105,N_16718,N_19280);
nor UO_106 (O_106,N_16287,N_19294);
nor UO_107 (O_107,N_16329,N_17368);
and UO_108 (O_108,N_16667,N_17844);
and UO_109 (O_109,N_15724,N_15924);
and UO_110 (O_110,N_16170,N_18869);
nand UO_111 (O_111,N_16449,N_17327);
and UO_112 (O_112,N_15037,N_19265);
or UO_113 (O_113,N_16964,N_17759);
and UO_114 (O_114,N_18313,N_19200);
nand UO_115 (O_115,N_16909,N_18889);
nor UO_116 (O_116,N_19641,N_17239);
and UO_117 (O_117,N_17871,N_19642);
and UO_118 (O_118,N_17843,N_18064);
nor UO_119 (O_119,N_15576,N_18080);
or UO_120 (O_120,N_15558,N_15331);
and UO_121 (O_121,N_18700,N_18062);
or UO_122 (O_122,N_19553,N_17988);
and UO_123 (O_123,N_15969,N_17061);
and UO_124 (O_124,N_17075,N_17666);
nor UO_125 (O_125,N_19562,N_16408);
nor UO_126 (O_126,N_18836,N_16807);
nor UO_127 (O_127,N_16599,N_18968);
nand UO_128 (O_128,N_16726,N_17269);
and UO_129 (O_129,N_19418,N_19173);
and UO_130 (O_130,N_19020,N_17411);
nor UO_131 (O_131,N_18074,N_15549);
nor UO_132 (O_132,N_15707,N_16505);
or UO_133 (O_133,N_19657,N_16099);
and UO_134 (O_134,N_18550,N_17661);
and UO_135 (O_135,N_18447,N_19838);
nor UO_136 (O_136,N_19388,N_17292);
nor UO_137 (O_137,N_16850,N_18398);
nor UO_138 (O_138,N_19523,N_16166);
nand UO_139 (O_139,N_19321,N_16611);
or UO_140 (O_140,N_15867,N_17804);
nor UO_141 (O_141,N_16949,N_16110);
and UO_142 (O_142,N_19621,N_18234);
nand UO_143 (O_143,N_17083,N_17647);
or UO_144 (O_144,N_19349,N_15071);
and UO_145 (O_145,N_18526,N_19060);
nor UO_146 (O_146,N_19005,N_17706);
nand UO_147 (O_147,N_19894,N_18982);
nand UO_148 (O_148,N_18405,N_15341);
or UO_149 (O_149,N_17322,N_16870);
and UO_150 (O_150,N_19798,N_15263);
nand UO_151 (O_151,N_16160,N_17435);
nand UO_152 (O_152,N_17145,N_15162);
or UO_153 (O_153,N_19287,N_19162);
nor UO_154 (O_154,N_17152,N_19061);
nand UO_155 (O_155,N_16262,N_18513);
or UO_156 (O_156,N_17649,N_19378);
nand UO_157 (O_157,N_18292,N_15951);
nor UO_158 (O_158,N_15255,N_15956);
or UO_159 (O_159,N_18706,N_16290);
nor UO_160 (O_160,N_16158,N_17633);
and UO_161 (O_161,N_18439,N_16180);
or UO_162 (O_162,N_17645,N_16386);
nor UO_163 (O_163,N_19805,N_19240);
nand UO_164 (O_164,N_16062,N_15719);
nor UO_165 (O_165,N_16184,N_18134);
nand UO_166 (O_166,N_16847,N_18715);
xor UO_167 (O_167,N_17862,N_18731);
and UO_168 (O_168,N_18456,N_17282);
nor UO_169 (O_169,N_19209,N_17915);
nand UO_170 (O_170,N_18849,N_19991);
nor UO_171 (O_171,N_15117,N_18746);
nor UO_172 (O_172,N_18077,N_17102);
and UO_173 (O_173,N_15895,N_17688);
and UO_174 (O_174,N_15191,N_16200);
or UO_175 (O_175,N_17247,N_18834);
and UO_176 (O_176,N_19690,N_17819);
nor UO_177 (O_177,N_17271,N_18221);
or UO_178 (O_178,N_17662,N_17350);
or UO_179 (O_179,N_19762,N_17413);
nand UO_180 (O_180,N_16995,N_19861);
nand UO_181 (O_181,N_18214,N_19134);
nor UO_182 (O_182,N_15733,N_18204);
or UO_183 (O_183,N_17041,N_15355);
or UO_184 (O_184,N_18309,N_16579);
nor UO_185 (O_185,N_18331,N_18400);
and UO_186 (O_186,N_17326,N_15232);
nand UO_187 (O_187,N_17297,N_19445);
or UO_188 (O_188,N_17829,N_19434);
or UO_189 (O_189,N_15963,N_16260);
nand UO_190 (O_190,N_18039,N_18703);
or UO_191 (O_191,N_15593,N_19620);
nor UO_192 (O_192,N_17336,N_18140);
or UO_193 (O_193,N_17216,N_17250);
xor UO_194 (O_194,N_16751,N_17425);
nand UO_195 (O_195,N_17803,N_18556);
or UO_196 (O_196,N_18795,N_17572);
nand UO_197 (O_197,N_18935,N_18287);
nand UO_198 (O_198,N_18319,N_15241);
and UO_199 (O_199,N_16443,N_17451);
and UO_200 (O_200,N_18955,N_15135);
nand UO_201 (O_201,N_17943,N_17655);
nand UO_202 (O_202,N_17436,N_19634);
and UO_203 (O_203,N_19897,N_15800);
nand UO_204 (O_204,N_17798,N_15463);
or UO_205 (O_205,N_17582,N_19518);
and UO_206 (O_206,N_18831,N_18719);
or UO_207 (O_207,N_17038,N_18219);
nand UO_208 (O_208,N_15659,N_15829);
or UO_209 (O_209,N_15290,N_19295);
or UO_210 (O_210,N_18994,N_15227);
nor UO_211 (O_211,N_19834,N_15058);
xnor UO_212 (O_212,N_16413,N_19215);
and UO_213 (O_213,N_18382,N_17566);
and UO_214 (O_214,N_17702,N_15204);
or UO_215 (O_215,N_16696,N_18264);
nor UO_216 (O_216,N_16966,N_19627);
or UO_217 (O_217,N_19852,N_19013);
nor UO_218 (O_218,N_18776,N_17396);
xor UO_219 (O_219,N_18675,N_17026);
nand UO_220 (O_220,N_19307,N_16946);
or UO_221 (O_221,N_17710,N_15766);
and UO_222 (O_222,N_15933,N_15493);
nand UO_223 (O_223,N_16164,N_15377);
xor UO_224 (O_224,N_18182,N_15955);
nor UO_225 (O_225,N_15340,N_18718);
xor UO_226 (O_226,N_17895,N_17818);
nand UO_227 (O_227,N_15189,N_18397);
nor UO_228 (O_228,N_17660,N_16346);
nor UO_229 (O_229,N_18651,N_17331);
or UO_230 (O_230,N_16988,N_15876);
nand UO_231 (O_231,N_19653,N_18307);
or UO_232 (O_232,N_17508,N_16634);
nand UO_233 (O_233,N_18815,N_17022);
or UO_234 (O_234,N_15185,N_18489);
nor UO_235 (O_235,N_15922,N_17932);
nand UO_236 (O_236,N_16962,N_15214);
and UO_237 (O_237,N_15433,N_15588);
and UO_238 (O_238,N_15115,N_17811);
nor UO_239 (O_239,N_15501,N_16183);
nor UO_240 (O_240,N_16476,N_16019);
nand UO_241 (O_241,N_19763,N_19969);
and UO_242 (O_242,N_16029,N_15392);
nand UO_243 (O_243,N_15578,N_19046);
or UO_244 (O_244,N_16253,N_19971);
or UO_245 (O_245,N_18471,N_18760);
nand UO_246 (O_246,N_17976,N_18862);
nand UO_247 (O_247,N_15869,N_19565);
nor UO_248 (O_248,N_18765,N_19591);
nor UO_249 (O_249,N_15008,N_15672);
nand UO_250 (O_250,N_16215,N_17616);
nor UO_251 (O_251,N_15423,N_16866);
nor UO_252 (O_252,N_19765,N_19302);
or UO_253 (O_253,N_15321,N_18939);
or UO_254 (O_254,N_18216,N_16193);
or UO_255 (O_255,N_19499,N_19733);
xnor UO_256 (O_256,N_19398,N_15775);
nor UO_257 (O_257,N_15090,N_18387);
or UO_258 (O_258,N_18433,N_16570);
nand UO_259 (O_259,N_19184,N_19407);
nand UO_260 (O_260,N_18227,N_19243);
nor UO_261 (O_261,N_17236,N_19975);
and UO_262 (O_262,N_15646,N_18738);
or UO_263 (O_263,N_16125,N_15381);
or UO_264 (O_264,N_18047,N_17595);
or UO_265 (O_265,N_15344,N_19192);
and UO_266 (O_266,N_19428,N_16101);
and UO_267 (O_267,N_16067,N_19421);
and UO_268 (O_268,N_15452,N_16776);
and UO_269 (O_269,N_19552,N_17450);
or UO_270 (O_270,N_19892,N_15998);
nor UO_271 (O_271,N_16994,N_19741);
nand UO_272 (O_272,N_19460,N_18951);
nor UO_273 (O_273,N_19055,N_17823);
or UO_274 (O_274,N_18095,N_16787);
and UO_275 (O_275,N_19555,N_16156);
and UO_276 (O_276,N_15249,N_18959);
or UO_277 (O_277,N_17786,N_16465);
nand UO_278 (O_278,N_18318,N_17054);
or UO_279 (O_279,N_18549,N_19609);
or UO_280 (O_280,N_18567,N_18372);
nor UO_281 (O_281,N_18021,N_19746);
or UO_282 (O_282,N_16093,N_19976);
nand UO_283 (O_283,N_18666,N_15562);
nand UO_284 (O_284,N_15403,N_16786);
and UO_285 (O_285,N_19457,N_18716);
nor UO_286 (O_286,N_18350,N_15474);
and UO_287 (O_287,N_19776,N_17963);
nor UO_288 (O_288,N_15026,N_18302);
nor UO_289 (O_289,N_16402,N_18791);
nor UO_290 (O_290,N_16323,N_15522);
and UO_291 (O_291,N_15720,N_19116);
nand UO_292 (O_292,N_17921,N_16433);
and UO_293 (O_293,N_18035,N_18168);
or UO_294 (O_294,N_17343,N_18936);
or UO_295 (O_295,N_19433,N_16147);
and UO_296 (O_296,N_17733,N_16586);
nand UO_297 (O_297,N_16675,N_15968);
and UO_298 (O_298,N_17371,N_17308);
and UO_299 (O_299,N_16334,N_16356);
nand UO_300 (O_300,N_17768,N_18535);
nor UO_301 (O_301,N_19264,N_19827);
and UO_302 (O_302,N_16021,N_17049);
and UO_303 (O_303,N_17567,N_15095);
nand UO_304 (O_304,N_16913,N_18083);
nor UO_305 (O_305,N_17264,N_15271);
nand UO_306 (O_306,N_19574,N_15286);
and UO_307 (O_307,N_15877,N_19255);
nor UO_308 (O_308,N_18341,N_17477);
nor UO_309 (O_309,N_18065,N_18463);
nand UO_310 (O_310,N_15936,N_18591);
nor UO_311 (O_311,N_15415,N_19468);
or UO_312 (O_312,N_17188,N_17092);
or UO_313 (O_313,N_17409,N_16367);
nand UO_314 (O_314,N_17491,N_16778);
nand UO_315 (O_315,N_17709,N_15838);
nor UO_316 (O_316,N_15616,N_16848);
and UO_317 (O_317,N_19203,N_15985);
and UO_318 (O_318,N_18629,N_16792);
or UO_319 (O_319,N_15508,N_18745);
nor UO_320 (O_320,N_17968,N_15175);
nor UO_321 (O_321,N_18152,N_16591);
or UO_322 (O_322,N_15088,N_17134);
and UO_323 (O_323,N_15890,N_19011);
and UO_324 (O_324,N_16742,N_19389);
nand UO_325 (O_325,N_18212,N_18749);
nor UO_326 (O_326,N_17469,N_16975);
nand UO_327 (O_327,N_18884,N_18407);
nor UO_328 (O_328,N_19496,N_18594);
nor UO_329 (O_329,N_17769,N_18491);
and UO_330 (O_330,N_15020,N_17744);
and UO_331 (O_331,N_16373,N_15518);
and UO_332 (O_332,N_15738,N_19906);
nand UO_333 (O_333,N_19232,N_17160);
and UO_334 (O_334,N_16908,N_15061);
and UO_335 (O_335,N_15866,N_15247);
or UO_336 (O_336,N_18838,N_19115);
and UO_337 (O_337,N_19836,N_16381);
nor UO_338 (O_338,N_15529,N_16243);
nor UO_339 (O_339,N_17187,N_17745);
and UO_340 (O_340,N_18317,N_17512);
and UO_341 (O_341,N_17266,N_16627);
or UO_342 (O_342,N_18695,N_16420);
or UO_343 (O_343,N_17640,N_15833);
and UO_344 (O_344,N_19954,N_18819);
and UO_345 (O_345,N_18984,N_18511);
nand UO_346 (O_346,N_15378,N_16605);
and UO_347 (O_347,N_18873,N_18123);
nand UO_348 (O_348,N_17931,N_19105);
or UO_349 (O_349,N_18435,N_17000);
nor UO_350 (O_350,N_17715,N_15285);
nand UO_351 (O_351,N_17283,N_18411);
or UO_352 (O_352,N_15427,N_19214);
nor UO_353 (O_353,N_17675,N_16468);
or UO_354 (O_354,N_15461,N_15305);
or UO_355 (O_355,N_16005,N_17626);
and UO_356 (O_356,N_16280,N_17265);
nor UO_357 (O_357,N_15821,N_19664);
and UO_358 (O_358,N_16017,N_16727);
or UO_359 (O_359,N_15600,N_17421);
nand UO_360 (O_360,N_15240,N_19787);
nand UO_361 (O_361,N_15499,N_18283);
nand UO_362 (O_362,N_15059,N_19384);
nand UO_363 (O_363,N_19871,N_18046);
nand UO_364 (O_364,N_17651,N_15010);
or UO_365 (O_365,N_15584,N_15478);
or UO_366 (O_366,N_15111,N_17213);
and UO_367 (O_367,N_15784,N_19800);
or UO_368 (O_368,N_16526,N_18342);
nor UO_369 (O_369,N_15170,N_15671);
xnor UO_370 (O_370,N_19500,N_16740);
nor UO_371 (O_371,N_15868,N_16151);
nor UO_372 (O_372,N_16583,N_18410);
nor UO_373 (O_373,N_19299,N_16623);
xnor UO_374 (O_374,N_18938,N_19411);
and UO_375 (O_375,N_17620,N_18139);
and UO_376 (O_376,N_15791,N_16135);
nor UO_377 (O_377,N_19990,N_15760);
nand UO_378 (O_378,N_17554,N_15676);
nand UO_379 (O_379,N_15443,N_17701);
or UO_380 (O_380,N_15222,N_15291);
nor UO_381 (O_381,N_16455,N_18965);
and UO_382 (O_382,N_15424,N_19029);
or UO_383 (O_383,N_15212,N_16555);
nand UO_384 (O_384,N_15744,N_17101);
and UO_385 (O_385,N_17021,N_19212);
nor UO_386 (O_386,N_18522,N_16084);
xor UO_387 (O_387,N_19363,N_18890);
nor UO_388 (O_388,N_18899,N_16142);
nand UO_389 (O_389,N_15633,N_19366);
nor UO_390 (O_390,N_18624,N_19718);
nand UO_391 (O_391,N_19174,N_17958);
and UO_392 (O_392,N_16519,N_18220);
and UO_393 (O_393,N_15181,N_17464);
nor UO_394 (O_394,N_19675,N_17796);
or UO_395 (O_395,N_19782,N_18101);
and UO_396 (O_396,N_19274,N_15533);
nor UO_397 (O_397,N_15995,N_19604);
nand UO_398 (O_398,N_15006,N_19545);
or UO_399 (O_399,N_15408,N_17547);
nor UO_400 (O_400,N_17964,N_16242);
nor UO_401 (O_401,N_15373,N_15831);
nand UO_402 (O_402,N_17791,N_18885);
and UO_403 (O_403,N_17034,N_17233);
nand UO_404 (O_404,N_16991,N_16003);
nand UO_405 (O_405,N_16722,N_16517);
nand UO_406 (O_406,N_17606,N_19491);
or UO_407 (O_407,N_17603,N_17474);
or UO_408 (O_408,N_15409,N_18677);
nor UO_409 (O_409,N_15345,N_16921);
and UO_410 (O_410,N_18284,N_19072);
and UO_411 (O_411,N_16672,N_17012);
or UO_412 (O_412,N_18115,N_15747);
nand UO_413 (O_413,N_17728,N_19695);
nand UO_414 (O_414,N_15056,N_18327);
nand UO_415 (O_415,N_16560,N_18306);
nand UO_416 (O_416,N_18243,N_18517);
nand UO_417 (O_417,N_17646,N_15063);
nor UO_418 (O_418,N_15685,N_19835);
nand UO_419 (O_419,N_15092,N_17154);
or UO_420 (O_420,N_19104,N_18085);
or UO_421 (O_421,N_16910,N_18539);
nor UO_422 (O_422,N_18037,N_17393);
nand UO_423 (O_423,N_15662,N_18497);
nor UO_424 (O_424,N_19027,N_18373);
and UO_425 (O_425,N_16499,N_16933);
nor UO_426 (O_426,N_19204,N_15993);
nand UO_427 (O_427,N_16635,N_18852);
or UO_428 (O_428,N_18430,N_19179);
or UO_429 (O_429,N_18256,N_17004);
nand UO_430 (O_430,N_19683,N_15050);
and UO_431 (O_431,N_16026,N_16543);
and UO_432 (O_432,N_19159,N_16601);
nand UO_433 (O_433,N_16869,N_18366);
and UO_434 (O_434,N_19968,N_15530);
nor UO_435 (O_435,N_18653,N_17043);
and UO_436 (O_436,N_18126,N_16856);
nor UO_437 (O_437,N_16640,N_16662);
nand UO_438 (O_438,N_18895,N_19638);
or UO_439 (O_439,N_15052,N_16620);
or UO_440 (O_440,N_16324,N_17929);
nand UO_441 (O_441,N_15076,N_17590);
or UO_442 (O_442,N_18725,N_19477);
nor UO_443 (O_443,N_15964,N_15012);
or UO_444 (O_444,N_19032,N_15627);
and UO_445 (O_445,N_16546,N_15704);
or UO_446 (O_446,N_19516,N_16438);
nand UO_447 (O_447,N_17426,N_15069);
and UO_448 (O_448,N_16755,N_19939);
xor UO_449 (O_449,N_15299,N_15252);
nor UO_450 (O_450,N_15464,N_19030);
or UO_451 (O_451,N_18036,N_19369);
nand UO_452 (O_452,N_18380,N_17010);
or UO_453 (O_453,N_17180,N_19917);
xor UO_454 (O_454,N_16883,N_18178);
nand UO_455 (O_455,N_15797,N_18782);
xor UO_456 (O_456,N_16550,N_15601);
nand UO_457 (O_457,N_15644,N_17738);
or UO_458 (O_458,N_16757,N_15690);
nor UO_459 (O_459,N_16508,N_15771);
and UO_460 (O_460,N_16312,N_16055);
xnor UO_461 (O_461,N_16340,N_18605);
and UO_462 (O_462,N_19858,N_16265);
nand UO_463 (O_463,N_18262,N_19651);
nand UO_464 (O_464,N_19033,N_16320);
xnor UO_465 (O_465,N_16141,N_18222);
nand UO_466 (O_466,N_16511,N_17475);
nand UO_467 (O_467,N_19228,N_19182);
nand UO_468 (O_468,N_17581,N_16784);
nand UO_469 (O_469,N_19401,N_16458);
nor UO_470 (O_470,N_16439,N_19448);
nand UO_471 (O_471,N_18509,N_17084);
or UO_472 (O_472,N_17055,N_15119);
nand UO_473 (O_473,N_17011,N_15035);
nor UO_474 (O_474,N_19826,N_15091);
or UO_475 (O_475,N_16596,N_17016);
or UO_476 (O_476,N_18930,N_15148);
or UO_477 (O_477,N_18124,N_15278);
nand UO_478 (O_478,N_19235,N_15713);
nand UO_479 (O_479,N_18466,N_19790);
or UO_480 (O_480,N_17085,N_16925);
nor UO_481 (O_481,N_15336,N_17109);
nand UO_482 (O_482,N_16626,N_15294);
or UO_483 (O_483,N_18799,N_16266);
or UO_484 (O_484,N_18980,N_19332);
and UO_485 (O_485,N_18590,N_17432);
or UO_486 (O_486,N_18141,N_19374);
nand UO_487 (O_487,N_16573,N_16024);
nand UO_488 (O_488,N_15314,N_16940);
nand UO_489 (O_489,N_18877,N_19272);
or UO_490 (O_490,N_19393,N_18086);
nor UO_491 (O_491,N_19558,N_18272);
nor UO_492 (O_492,N_19336,N_17850);
nor UO_493 (O_493,N_18747,N_19514);
nand UO_494 (O_494,N_17639,N_17219);
or UO_495 (O_495,N_18417,N_18763);
and UO_496 (O_496,N_15681,N_15539);
nand UO_497 (O_497,N_19994,N_15749);
nor UO_498 (O_498,N_15650,N_19122);
nand UO_499 (O_499,N_16085,N_19247);
nand UO_500 (O_500,N_17604,N_15500);
and UO_501 (O_501,N_18465,N_16681);
nand UO_502 (O_502,N_17462,N_15666);
or UO_503 (O_503,N_19660,N_19313);
or UO_504 (O_504,N_17782,N_17483);
and UO_505 (O_505,N_16059,N_17303);
nand UO_506 (O_506,N_15108,N_17365);
or UO_507 (O_507,N_16371,N_19537);
or UO_508 (O_508,N_16404,N_19813);
or UO_509 (O_509,N_17500,N_17267);
or UO_510 (O_510,N_15398,N_15310);
nor UO_511 (O_511,N_16911,N_17254);
and UO_512 (O_512,N_16965,N_19051);
nor UO_513 (O_513,N_16122,N_16349);
or UO_514 (O_514,N_18383,N_18681);
nor UO_515 (O_515,N_18562,N_16781);
xor UO_516 (O_516,N_15239,N_19796);
nand UO_517 (O_517,N_19035,N_19158);
nor UO_518 (O_518,N_18902,N_16480);
nor UO_519 (O_519,N_15425,N_15384);
and UO_520 (O_520,N_15698,N_15237);
nand UO_521 (O_521,N_16031,N_15628);
or UO_522 (O_522,N_19327,N_18584);
nor UO_523 (O_523,N_17433,N_16470);
and UO_524 (O_524,N_17677,N_17637);
nand UO_525 (O_525,N_17238,N_15759);
or UO_526 (O_526,N_15146,N_15978);
or UO_527 (O_527,N_17904,N_15575);
nor UO_528 (O_528,N_17611,N_16944);
nor UO_529 (O_529,N_19419,N_16587);
nor UO_530 (O_530,N_19960,N_19902);
nor UO_531 (O_531,N_18505,N_17153);
nand UO_532 (O_532,N_16407,N_16429);
nor UO_533 (O_533,N_19087,N_18067);
nor UO_534 (O_534,N_16703,N_17695);
and UO_535 (O_535,N_19546,N_16130);
or UO_536 (O_536,N_17515,N_16922);
nor UO_537 (O_537,N_19385,N_19819);
nor UO_538 (O_538,N_19316,N_18072);
or UO_539 (O_539,N_17445,N_15366);
or UO_540 (O_540,N_19368,N_19949);
nor UO_541 (O_541,N_19186,N_16143);
or UO_542 (O_542,N_18347,N_17193);
nand UO_543 (O_543,N_18474,N_19279);
nor UO_544 (O_544,N_18051,N_16315);
nor UO_545 (O_545,N_16531,N_15113);
nand UO_546 (O_546,N_15416,N_15445);
or UO_547 (O_547,N_18609,N_16399);
and UO_548 (O_548,N_18003,N_18002);
nor UO_549 (O_549,N_17800,N_15141);
xor UO_550 (O_550,N_16043,N_18579);
nand UO_551 (O_551,N_18736,N_17897);
and UO_552 (O_552,N_19245,N_15228);
or UO_553 (O_553,N_15728,N_17992);
or UO_554 (O_554,N_15894,N_15731);
and UO_555 (O_555,N_18741,N_16858);
nor UO_556 (O_556,N_16985,N_16298);
and UO_557 (O_557,N_18668,N_17284);
nor UO_558 (O_558,N_18825,N_15571);
xnor UO_559 (O_559,N_16203,N_15789);
and UO_560 (O_560,N_17067,N_19014);
nor UO_561 (O_561,N_17588,N_18162);
nor UO_562 (O_562,N_19870,N_17845);
nand UO_563 (O_563,N_16907,N_17730);
or UO_564 (O_564,N_17914,N_15893);
or UO_565 (O_565,N_17941,N_17293);
or UO_566 (O_566,N_17058,N_16409);
and UO_567 (O_567,N_19578,N_15811);
nand UO_568 (O_568,N_16923,N_18266);
and UO_569 (O_569,N_16876,N_16917);
nand UO_570 (O_570,N_19399,N_18110);
or UO_571 (O_571,N_17987,N_17749);
or UO_572 (O_572,N_17316,N_17984);
nand UO_573 (O_573,N_18113,N_16418);
and UO_574 (O_574,N_18111,N_17178);
nand UO_575 (O_575,N_18479,N_16768);
or UO_576 (O_576,N_17935,N_15420);
nor UO_577 (O_577,N_16355,N_19237);
nor UO_578 (O_578,N_19037,N_17560);
nor UO_579 (O_579,N_18109,N_16196);
nor UO_580 (O_580,N_15243,N_19599);
nor UO_581 (O_581,N_15973,N_16089);
xor UO_582 (O_582,N_17600,N_19082);
nor UO_583 (O_583,N_16393,N_19106);
or UO_584 (O_584,N_18345,N_17005);
nor UO_585 (O_585,N_19168,N_19259);
and UO_586 (O_586,N_15883,N_18336);
nor UO_587 (O_587,N_18329,N_17071);
or UO_588 (O_588,N_18920,N_17937);
nand UO_589 (O_589,N_16421,N_18612);
nand UO_590 (O_590,N_19488,N_17237);
nand UO_591 (O_591,N_19617,N_17877);
nor UO_592 (O_592,N_16832,N_15958);
or UO_593 (O_593,N_17928,N_19824);
nor UO_594 (O_594,N_17780,N_19251);
xnor UO_595 (O_595,N_19862,N_17068);
nor UO_596 (O_596,N_15174,N_19946);
and UO_597 (O_597,N_15917,N_16780);
nor UO_598 (O_598,N_15861,N_18241);
or UO_599 (O_599,N_19770,N_17790);
and UO_600 (O_600,N_15428,N_17214);
and UO_601 (O_601,N_19847,N_16118);
and UO_602 (O_602,N_19497,N_16139);
nand UO_603 (O_603,N_16624,N_16425);
and UO_604 (O_604,N_16976,N_15834);
nand UO_605 (O_605,N_19090,N_15954);
or UO_606 (O_606,N_18940,N_15209);
nand UO_607 (O_607,N_16844,N_16827);
and UO_608 (O_608,N_15472,N_18040);
nor UO_609 (O_609,N_18194,N_18784);
or UO_610 (O_610,N_15358,N_15696);
or UO_611 (O_611,N_15788,N_17942);
nand UO_612 (O_612,N_15765,N_16384);
and UO_613 (O_613,N_15083,N_17682);
nand UO_614 (O_614,N_19219,N_19036);
nand UO_615 (O_615,N_16636,N_18643);
nand UO_616 (O_616,N_19885,N_19364);
nand UO_617 (O_617,N_19757,N_15642);
or UO_618 (O_618,N_17203,N_17035);
or UO_619 (O_619,N_19597,N_15318);
nand UO_620 (O_620,N_17466,N_18710);
or UO_621 (O_621,N_18401,N_16506);
or UO_622 (O_622,N_15051,N_19205);
nor UO_623 (O_623,N_19193,N_16617);
nor UO_624 (O_624,N_18974,N_19242);
or UO_625 (O_625,N_15487,N_16091);
nor UO_626 (O_626,N_19880,N_15886);
and UO_627 (O_627,N_17132,N_18788);
and UO_628 (O_628,N_16841,N_18233);
and UO_629 (O_629,N_18503,N_16589);
nor UO_630 (O_630,N_18580,N_16545);
and UO_631 (O_631,N_15517,N_19804);
or UO_632 (O_632,N_17610,N_19652);
nor UO_633 (O_633,N_16057,N_19281);
and UO_634 (O_634,N_19676,N_19841);
nor UO_635 (O_635,N_16715,N_15967);
and UO_636 (O_636,N_16086,N_19955);
nand UO_637 (O_637,N_18759,N_19811);
and UO_638 (O_638,N_17954,N_15972);
nor UO_639 (O_639,N_19107,N_16572);
nor UO_640 (O_640,N_19588,N_19334);
nand UO_641 (O_641,N_17105,N_17096);
nand UO_642 (O_642,N_16169,N_16163);
nor UO_643 (O_643,N_18857,N_15123);
nand UO_644 (O_644,N_16152,N_16688);
or UO_645 (O_645,N_17857,N_18481);
nand UO_646 (O_646,N_18228,N_17318);
and UO_647 (O_647,N_16738,N_19887);
nor UO_648 (O_648,N_17431,N_19408);
and UO_649 (O_649,N_18742,N_15068);
and UO_650 (O_650,N_18082,N_19995);
nor UO_651 (O_651,N_17644,N_15631);
nor UO_652 (O_652,N_15114,N_15401);
and UO_653 (O_653,N_19402,N_17143);
nand UO_654 (O_654,N_17641,N_18724);
nand UO_655 (O_655,N_17389,N_15561);
or UO_656 (O_656,N_16770,N_17789);
nand UO_657 (O_657,N_18802,N_16803);
nor UO_658 (O_658,N_17215,N_15595);
and UO_659 (O_659,N_16548,N_18705);
nor UO_660 (O_660,N_17830,N_19413);
and UO_661 (O_661,N_17384,N_17699);
nand UO_662 (O_662,N_16915,N_16889);
and UO_663 (O_663,N_19803,N_16552);
or UO_664 (O_664,N_16732,N_19981);
nand UO_665 (O_665,N_15632,N_16405);
and UO_666 (O_666,N_15405,N_15983);
nand UO_667 (O_667,N_16588,N_17151);
nand UO_668 (O_668,N_18041,N_17452);
nand UO_669 (O_669,N_15581,N_15557);
or UO_670 (O_670,N_18364,N_17225);
nor UO_671 (O_671,N_19561,N_19121);
nor UO_672 (O_672,N_17329,N_15001);
nor UO_673 (O_673,N_17399,N_17459);
nand UO_674 (O_674,N_16370,N_19964);
nand UO_675 (O_675,N_18694,N_18158);
nand UO_676 (O_676,N_15154,N_15805);
nand UO_677 (O_677,N_15695,N_15904);
nor UO_678 (O_678,N_15842,N_17696);
nand UO_679 (O_679,N_19935,N_15412);
and UO_680 (O_680,N_19067,N_15622);
nor UO_681 (O_681,N_18138,N_18679);
nor UO_682 (O_682,N_15437,N_19973);
or UO_683 (O_683,N_19893,N_16068);
or UO_684 (O_684,N_15441,N_15322);
nand UO_685 (O_685,N_16698,N_19525);
or UO_686 (O_686,N_15176,N_15107);
nor UO_687 (O_687,N_15928,N_15959);
and UO_688 (O_688,N_19111,N_19387);
or UO_689 (O_689,N_15093,N_18828);
and UO_690 (O_690,N_16446,N_17832);
nor UO_691 (O_691,N_19155,N_19998);
or UO_692 (O_692,N_17140,N_19484);
xnor UO_693 (O_693,N_17165,N_19859);
nor UO_694 (O_694,N_18797,N_15637);
nand UO_695 (O_695,N_18734,N_18807);
or UO_696 (O_696,N_19019,N_18658);
or UO_697 (O_697,N_18673,N_16830);
and UO_698 (O_698,N_16452,N_15888);
or UO_699 (O_699,N_17150,N_16013);
nand UO_700 (O_700,N_15297,N_15475);
and UO_701 (O_701,N_15077,N_16167);
or UO_702 (O_702,N_16348,N_18837);
nand UO_703 (O_703,N_17230,N_17347);
or UO_704 (O_704,N_18551,N_16802);
or UO_705 (O_705,N_15289,N_17636);
nand UO_706 (O_706,N_15810,N_16679);
and UO_707 (O_707,N_17319,N_18449);
nand UO_708 (O_708,N_17360,N_17561);
and UO_709 (O_709,N_15145,N_18106);
and UO_710 (O_710,N_17476,N_18050);
nor UO_711 (O_711,N_19278,N_18687);
nand UO_712 (O_712,N_18983,N_19950);
or UO_713 (O_713,N_18723,N_16817);
or UO_714 (O_714,N_16686,N_15535);
nor UO_715 (O_715,N_19926,N_16796);
nor UO_716 (O_716,N_16423,N_18993);
nor UO_717 (O_717,N_17808,N_17886);
or UO_718 (O_718,N_16947,N_19766);
or UO_719 (O_719,N_18142,N_16250);
nand UO_720 (O_720,N_19330,N_16642);
or UO_721 (O_721,N_19570,N_16561);
nand UO_722 (O_722,N_16114,N_18811);
xnor UO_723 (O_723,N_16009,N_16008);
nand UO_724 (O_724,N_17418,N_17039);
or UO_725 (O_725,N_19794,N_17549);
and UO_726 (O_726,N_18130,N_16603);
or UO_727 (O_727,N_16704,N_19735);
or UO_728 (O_728,N_18335,N_19260);
nand UO_729 (O_729,N_19475,N_18625);
or UO_730 (O_730,N_15150,N_18377);
or UO_731 (O_731,N_18801,N_15567);
nor UO_732 (O_732,N_18552,N_19679);
nor UO_733 (O_733,N_19085,N_19463);
nor UO_734 (O_734,N_15447,N_16479);
nor UO_735 (O_735,N_15498,N_18870);
or UO_736 (O_736,N_17118,N_19605);
nor UO_737 (O_737,N_17841,N_16115);
nand UO_738 (O_738,N_18645,N_15617);
nor UO_739 (O_739,N_19869,N_17485);
nor UO_740 (O_740,N_16406,N_19635);
or UO_741 (O_741,N_19684,N_17587);
nor UO_742 (O_742,N_17869,N_16053);
nor UO_743 (O_743,N_18167,N_18515);
nor UO_744 (O_744,N_15808,N_19022);
or UO_745 (O_745,N_18961,N_16431);
or UO_746 (O_746,N_18617,N_18969);
or UO_747 (O_747,N_18330,N_18218);
nand UO_748 (O_748,N_15368,N_15167);
nor UO_749 (O_749,N_19972,N_15178);
and UO_750 (O_750,N_17957,N_16345);
and UO_751 (O_751,N_15513,N_18502);
nor UO_752 (O_752,N_17720,N_18388);
nor UO_753 (O_753,N_18754,N_16816);
or UO_754 (O_754,N_15246,N_16647);
nor UO_755 (O_755,N_19569,N_18548);
nand UO_756 (O_756,N_15363,N_18348);
nor UO_757 (O_757,N_17471,N_18013);
nand UO_758 (O_758,N_19490,N_16228);
nor UO_759 (O_759,N_19978,N_15062);
nand UO_760 (O_760,N_15741,N_17148);
or UO_761 (O_761,N_19650,N_18998);
nor UO_762 (O_762,N_17784,N_15796);
and UO_763 (O_763,N_15551,N_16221);
nand UO_764 (O_764,N_19547,N_19430);
nand UO_765 (O_765,N_16245,N_17351);
nor UO_766 (O_766,N_16368,N_15717);
nand UO_767 (O_767,N_17854,N_17366);
nor UO_768 (O_768,N_16457,N_18946);
nor UO_769 (O_769,N_19817,N_18324);
or UO_770 (O_770,N_19786,N_17372);
nor UO_771 (O_771,N_16220,N_17985);
nand UO_772 (O_772,N_16684,N_16774);
nand UO_773 (O_773,N_15526,N_18911);
nor UO_774 (O_774,N_15233,N_17511);
and UO_775 (O_775,N_15860,N_19028);
and UO_776 (O_776,N_19257,N_15203);
or UO_777 (O_777,N_18574,N_17615);
and UO_778 (O_778,N_16811,N_18295);
nor UO_779 (O_779,N_18577,N_16668);
or UO_780 (O_780,N_15367,N_17597);
or UO_781 (O_781,N_16006,N_18650);
and UO_782 (O_782,N_18835,N_18616);
or UO_783 (O_783,N_19322,N_16797);
or UO_784 (O_784,N_16953,N_16853);
and UO_785 (O_785,N_17195,N_16891);
or UO_786 (O_786,N_17300,N_15057);
nor UO_787 (O_787,N_17046,N_15049);
nand UO_788 (O_788,N_18744,N_19934);
or UO_789 (O_789,N_18581,N_18058);
nand UO_790 (O_790,N_15665,N_15453);
or UO_791 (O_791,N_18827,N_17053);
nand UO_792 (O_792,N_19231,N_18894);
or UO_793 (O_793,N_19338,N_17531);
or UO_794 (O_794,N_17458,N_16880);
or UO_795 (O_795,N_17933,N_19070);
nand UO_796 (O_796,N_18589,N_17299);
or UO_797 (O_797,N_17760,N_15312);
xnor UO_798 (O_798,N_18972,N_16772);
nand UO_799 (O_799,N_15136,N_18660);
nor UO_800 (O_800,N_18674,N_15975);
or UO_801 (O_801,N_17013,N_18855);
xor UO_802 (O_802,N_18758,N_18728);
nor UO_803 (O_803,N_16388,N_18164);
nand UO_804 (O_804,N_19822,N_16481);
nor UO_805 (O_805,N_17821,N_17212);
and UO_806 (O_806,N_17810,N_15837);
and UO_807 (O_807,N_17839,N_18144);
nor UO_808 (O_808,N_15828,N_15686);
xnor UO_809 (O_809,N_16277,N_18572);
nand UO_810 (O_810,N_19380,N_18785);
or UO_811 (O_811,N_17437,N_19449);
or UO_812 (O_812,N_15065,N_15158);
and UO_813 (O_813,N_19713,N_15740);
nand UO_814 (O_814,N_19271,N_15763);
or UO_815 (O_815,N_18464,N_18823);
nor UO_816 (O_816,N_18777,N_16828);
and UO_817 (O_817,N_19818,N_15122);
or UO_818 (O_818,N_19504,N_16338);
nand UO_819 (O_819,N_17183,N_18120);
or UO_820 (O_820,N_16790,N_17163);
or UO_821 (O_821,N_16609,N_18853);
nand UO_822 (O_822,N_15839,N_17755);
nor UO_823 (O_823,N_17605,N_19130);
nand UO_824 (O_824,N_18495,N_16899);
and UO_825 (O_825,N_17983,N_19343);
nand UO_826 (O_826,N_15899,N_18621);
and UO_827 (O_827,N_16191,N_19807);
or UO_828 (O_828,N_16906,N_17495);
or UO_829 (O_829,N_17113,N_18022);
nor UO_830 (O_830,N_17320,N_15352);
or UO_831 (O_831,N_15772,N_15147);
or UO_832 (O_832,N_15528,N_19443);
nor UO_833 (O_833,N_17685,N_16461);
and UO_834 (O_834,N_17408,N_18177);
or UO_835 (O_835,N_15103,N_18709);
and UO_836 (O_836,N_15537,N_16934);
or UO_837 (O_837,N_15307,N_16012);
nor UO_838 (O_838,N_15836,N_15126);
nand UO_839 (O_839,N_16205,N_16098);
nor UO_840 (O_840,N_19062,N_16317);
nor UO_841 (O_841,N_17521,N_16812);
or UO_842 (O_842,N_19789,N_18114);
or UO_843 (O_843,N_17936,N_18970);
nand UO_844 (O_844,N_18189,N_16222);
xor UO_845 (O_845,N_19396,N_19309);
and UO_846 (O_846,N_15813,N_16498);
and UO_847 (O_847,N_16254,N_16534);
and UO_848 (O_848,N_19758,N_16719);
nand UO_849 (O_849,N_15046,N_15906);
or UO_850 (O_850,N_18879,N_19135);
xor UO_851 (O_851,N_18667,N_16924);
nor UO_852 (O_852,N_17668,N_16747);
nand UO_853 (O_853,N_16469,N_17161);
nand UO_854 (O_854,N_15598,N_16155);
or UO_855 (O_855,N_19845,N_19097);
and UO_856 (O_856,N_16657,N_15809);
and UO_857 (O_857,N_17774,N_16762);
nor UO_858 (O_858,N_17534,N_15544);
xor UO_859 (O_859,N_17608,N_15516);
nor UO_860 (O_860,N_17024,N_16963);
nand UO_861 (O_861,N_16397,N_19607);
nor UO_862 (O_862,N_16240,N_19630);
and UO_863 (O_863,N_17920,N_16584);
nand UO_864 (O_864,N_16693,N_19276);
nand UO_865 (O_865,N_19613,N_16919);
or UO_866 (O_866,N_16283,N_19535);
nor UO_867 (O_867,N_16996,N_15977);
nor UO_868 (O_868,N_16311,N_15389);
or UO_869 (O_869,N_15276,N_19273);
and UO_870 (O_870,N_19532,N_19216);
nor UO_871 (O_871,N_18992,N_15540);
nand UO_872 (O_872,N_18730,N_18954);
xnor UO_873 (O_873,N_19201,N_17077);
or UO_874 (O_874,N_17901,N_18628);
and UO_875 (O_875,N_18420,N_18049);
and UO_876 (O_876,N_17257,N_16485);
or UO_877 (O_877,N_16496,N_18422);
and UO_878 (O_878,N_15726,N_16931);
nor UO_879 (O_879,N_17948,N_16375);
nor UO_880 (O_880,N_19524,N_18232);
xor UO_881 (O_881,N_15945,N_18312);
nor UO_882 (O_882,N_18184,N_15072);
nand UO_883 (O_883,N_19452,N_19124);
and UO_884 (O_884,N_18274,N_15362);
nor UO_885 (O_885,N_16671,N_18816);
nand UO_886 (O_886,N_18603,N_17625);
nor UO_887 (O_887,N_15524,N_19707);
or UO_888 (O_888,N_19120,N_18926);
and UO_889 (O_889,N_15468,N_17244);
nor UO_890 (O_890,N_18780,N_17492);
or UO_891 (O_891,N_16523,N_19125);
nand UO_892 (O_892,N_17623,N_16559);
xor UO_893 (O_893,N_16836,N_17947);
nor UO_894 (O_894,N_15317,N_18267);
and UO_895 (O_895,N_16632,N_19697);
or UO_896 (O_896,N_16553,N_16864);
nand UO_897 (O_897,N_18803,N_15000);
nor UO_898 (O_898,N_15440,N_18242);
nand UO_899 (O_899,N_15481,N_19031);
xor UO_900 (O_900,N_19092,N_16663);
or UO_901 (O_901,N_15319,N_17571);
nor UO_902 (O_902,N_15974,N_18247);
nor UO_903 (O_903,N_17349,N_18052);
or UO_904 (O_904,N_17031,N_18919);
or UO_905 (O_905,N_18136,N_16501);
and UO_906 (O_906,N_15075,N_19469);
nand UO_907 (O_907,N_15268,N_18310);
nand UO_908 (O_908,N_17170,N_15892);
and UO_909 (O_909,N_16678,N_18029);
nand UO_910 (O_910,N_16072,N_18135);
or UO_911 (O_911,N_15495,N_15762);
and UO_912 (O_912,N_19624,N_17540);
and UO_913 (O_913,N_16893,N_18244);
and UO_914 (O_914,N_15815,N_16120);
nor UO_915 (O_915,N_17123,N_15096);
nand UO_916 (O_916,N_15027,N_16544);
nor UO_917 (O_917,N_15774,N_16670);
and UO_918 (O_918,N_15846,N_19109);
and UO_919 (O_919,N_17858,N_17757);
nand UO_920 (O_920,N_19566,N_16258);
nor UO_921 (O_921,N_17441,N_16750);
nor UO_922 (O_922,N_15548,N_15986);
nand UO_923 (O_923,N_15300,N_16432);
nor UO_924 (O_924,N_15949,N_18648);
or UO_925 (O_925,N_17729,N_16038);
nand UO_926 (O_926,N_17222,N_19732);
and UO_927 (O_927,N_16267,N_16430);
or UO_928 (O_928,N_16687,N_18360);
or UO_929 (O_929,N_16813,N_16540);
nor UO_930 (O_930,N_16269,N_19575);
or UO_931 (O_931,N_16301,N_19953);
or UO_932 (O_932,N_18848,N_19866);
and UO_933 (O_933,N_16753,N_15654);
xnor UO_934 (O_934,N_16576,N_18104);
and UO_935 (O_935,N_15281,N_15611);
nor UO_936 (O_936,N_17898,N_15161);
nor UO_937 (O_937,N_15320,N_15469);
or UO_938 (O_938,N_18904,N_15238);
or UO_939 (O_939,N_15242,N_18541);
and UO_940 (O_940,N_19596,N_16357);
nand UO_941 (O_941,N_17375,N_16119);
nand UO_942 (O_942,N_18132,N_18636);
nand UO_943 (O_943,N_16536,N_16185);
and UO_944 (O_944,N_16252,N_18563);
nand UO_945 (O_945,N_19600,N_18547);
and UO_946 (O_946,N_16113,N_18297);
and UO_947 (O_947,N_16326,N_16754);
and UO_948 (O_948,N_16097,N_17252);
nand UO_949 (O_949,N_17025,N_18451);
nand UO_950 (O_950,N_17044,N_17691);
nand UO_951 (O_951,N_19728,N_18100);
nor UO_952 (O_952,N_16415,N_16477);
and UO_953 (O_953,N_16478,N_17993);
nor UO_954 (O_954,N_18595,N_19277);
nand UO_955 (O_955,N_15043,N_18057);
nor UO_956 (O_956,N_18402,N_19021);
nor UO_957 (O_957,N_15620,N_16018);
nor UO_958 (O_958,N_18598,N_18523);
or UO_959 (O_959,N_16302,N_16377);
nand UO_960 (O_960,N_17902,N_17982);
nor UO_961 (O_961,N_19864,N_19303);
nor UO_962 (O_962,N_19610,N_15293);
nand UO_963 (O_963,N_17658,N_19096);
and UO_964 (O_964,N_18119,N_19367);
or UO_965 (O_965,N_19053,N_18670);
nor UO_966 (O_966,N_15430,N_17874);
and UO_967 (O_967,N_18771,N_16782);
nor UO_968 (O_968,N_19840,N_19850);
nand UO_969 (O_969,N_19521,N_19471);
nor UO_970 (O_970,N_16999,N_18842);
nand UO_971 (O_971,N_16343,N_16264);
and UO_972 (O_972,N_18818,N_17556);
xnor UO_973 (O_973,N_19996,N_15976);
or UO_974 (O_974,N_19785,N_19354);
nand UO_975 (O_975,N_16798,N_15301);
or UO_976 (O_976,N_19357,N_15094);
nand UO_977 (O_977,N_15653,N_16938);
nor UO_978 (O_978,N_18001,N_15931);
or UO_979 (O_979,N_16374,N_18909);
and UO_980 (O_980,N_17557,N_17714);
and UO_981 (O_981,N_15932,N_19439);
nand UO_982 (O_982,N_17261,N_18180);
nor UO_983 (O_983,N_18956,N_17607);
nand UO_984 (O_984,N_15053,N_17835);
and UO_985 (O_985,N_19136,N_17062);
nor UO_986 (O_986,N_16482,N_19297);
nand UO_987 (O_987,N_18804,N_17428);
or UO_988 (O_988,N_17986,N_16956);
nand UO_989 (O_989,N_18534,N_18587);
nor UO_990 (O_990,N_19857,N_16063);
nand UO_991 (O_991,N_17761,N_19505);
or UO_992 (O_992,N_18320,N_18412);
nor UO_993 (O_993,N_15667,N_17613);
nand UO_994 (O_994,N_17872,N_17772);
or UO_995 (O_995,N_19306,N_17340);
or UO_996 (O_996,N_15887,N_15912);
nand UO_997 (O_997,N_16208,N_17325);
and UO_998 (O_998,N_18424,N_15521);
nand UO_999 (O_999,N_17367,N_19291);
nor UO_1000 (O_1000,N_17137,N_16614);
nor UO_1001 (O_1001,N_15031,N_18864);
nand UO_1002 (O_1002,N_19425,N_19681);
xor UO_1003 (O_1003,N_18664,N_16537);
nor UO_1004 (O_1004,N_18116,N_18009);
nor UO_1005 (O_1005,N_15234,N_19750);
or UO_1006 (O_1006,N_17497,N_17618);
xor UO_1007 (O_1007,N_19721,N_19517);
and UO_1008 (O_1008,N_17771,N_19922);
and UO_1009 (O_1009,N_17907,N_16633);
and UO_1010 (O_1010,N_15070,N_19152);
and UO_1011 (O_1011,N_16701,N_18947);
nand UO_1012 (O_1012,N_15602,N_19703);
and UO_1013 (O_1013,N_16278,N_17959);
nand UO_1014 (O_1014,N_15639,N_16948);
nor UO_1015 (O_1015,N_16045,N_19113);
or UO_1016 (O_1016,N_15547,N_15674);
or UO_1017 (O_1017,N_17596,N_15047);
or UO_1018 (O_1018,N_15721,N_17383);
xor UO_1019 (O_1019,N_17208,N_15250);
and UO_1020 (O_1020,N_19100,N_18773);
and UO_1021 (O_1021,N_18484,N_19706);
or UO_1022 (O_1022,N_15306,N_17103);
nand UO_1023 (O_1023,N_15505,N_17179);
and UO_1024 (O_1024,N_15718,N_15802);
and UO_1025 (O_1025,N_16749,N_16105);
nor UO_1026 (O_1026,N_16843,N_18185);
or UO_1027 (O_1027,N_19170,N_15661);
nor UO_1028 (O_1028,N_18131,N_18735);
nand UO_1029 (O_1029,N_19693,N_17217);
nand UO_1030 (O_1030,N_19557,N_16788);
xor UO_1031 (O_1031,N_18005,N_16145);
and UO_1032 (O_1032,N_16779,N_19944);
and UO_1033 (O_1033,N_19519,N_16967);
or UO_1034 (O_1034,N_19180,N_19006);
nor UO_1035 (O_1035,N_16785,N_19211);
nand UO_1036 (O_1036,N_16460,N_19310);
nand UO_1037 (O_1037,N_19806,N_19692);
and UO_1038 (O_1038,N_15248,N_16775);
or UO_1039 (O_1039,N_15900,N_16181);
and UO_1040 (O_1040,N_19878,N_17467);
and UO_1041 (O_1041,N_15213,N_15349);
nand UO_1042 (O_1042,N_17339,N_17580);
and UO_1043 (O_1043,N_15583,N_16767);
or UO_1044 (O_1044,N_17040,N_15577);
and UO_1045 (O_1045,N_15634,N_18631);
nor UO_1046 (O_1046,N_15748,N_19286);
nand UO_1047 (O_1047,N_17776,N_17111);
and UO_1048 (O_1048,N_15923,N_19967);
nand UO_1049 (O_1049,N_15303,N_17394);
nor UO_1050 (O_1050,N_18416,N_17667);
nand UO_1051 (O_1051,N_17306,N_19304);
nand UO_1052 (O_1052,N_18395,N_19755);
or UO_1053 (O_1053,N_16527,N_19091);
and UO_1054 (O_1054,N_15328,N_15937);
and UO_1055 (O_1055,N_18389,N_18450);
nor UO_1056 (O_1056,N_15467,N_16186);
nor UO_1057 (O_1057,N_15756,N_19009);
nand UO_1058 (O_1058,N_17578,N_17910);
nor UO_1059 (O_1059,N_17045,N_19710);
nor UO_1060 (O_1060,N_18840,N_19874);
or UO_1061 (O_1061,N_17562,N_15502);
nor UO_1062 (O_1062,N_16108,N_15872);
and UO_1063 (O_1063,N_19447,N_18000);
nand UO_1064 (O_1064,N_16892,N_17232);
and UO_1065 (O_1065,N_16739,N_17392);
nand UO_1066 (O_1066,N_19915,N_16664);
nand UO_1067 (O_1067,N_19194,N_15229);
or UO_1068 (O_1068,N_16823,N_19779);
or UO_1069 (O_1069,N_16855,N_18483);
or UO_1070 (O_1070,N_17552,N_19079);
or UO_1071 (O_1071,N_18755,N_19700);
xor UO_1072 (O_1072,N_15066,N_17659);
nand UO_1073 (O_1073,N_15757,N_15196);
nand UO_1074 (O_1074,N_17243,N_15660);
xor UO_1075 (O_1075,N_16319,N_19054);
nor UO_1076 (O_1076,N_19123,N_15417);
nor UO_1077 (O_1077,N_15550,N_16244);
or UO_1078 (O_1078,N_15663,N_16769);
or UO_1079 (O_1079,N_17259,N_18246);
and UO_1080 (O_1080,N_19756,N_15361);
nand UO_1081 (O_1081,N_17377,N_16488);
and UO_1082 (O_1082,N_17532,N_16492);
nand UO_1083 (O_1083,N_19714,N_15223);
nor UO_1084 (O_1084,N_16928,N_19199);
xnor UO_1085 (O_1085,N_19506,N_16234);
nor UO_1086 (O_1086,N_16539,N_16525);
nand UO_1087 (O_1087,N_19891,N_18806);
nand UO_1088 (O_1088,N_15338,N_15370);
nand UO_1089 (O_1089,N_19914,N_15697);
nor UO_1090 (O_1090,N_17104,N_15353);
nand UO_1091 (O_1091,N_18386,N_15116);
and UO_1092 (O_1092,N_18767,N_15280);
or UO_1093 (O_1093,N_16467,N_17589);
or UO_1094 (O_1094,N_16366,N_16690);
nand UO_1095 (O_1095,N_18406,N_16182);
and UO_1096 (O_1096,N_17412,N_15640);
or UO_1097 (O_1097,N_17781,N_16973);
nor UO_1098 (O_1098,N_19000,N_18976);
and UO_1099 (O_1099,N_17194,N_15391);
and UO_1100 (O_1100,N_17223,N_19730);
and UO_1101 (O_1101,N_16124,N_16520);
nor UO_1102 (O_1102,N_19848,N_16970);
nor UO_1103 (O_1103,N_17014,N_19511);
and UO_1104 (O_1104,N_15034,N_18254);
or UO_1105 (O_1105,N_17009,N_17385);
and UO_1106 (O_1106,N_17249,N_17363);
nor UO_1107 (O_1107,N_16424,N_15457);
nor UO_1108 (O_1108,N_15701,N_17310);
and UO_1109 (O_1109,N_19153,N_18314);
or UO_1110 (O_1110,N_19951,N_18898);
nand UO_1111 (O_1111,N_17894,N_16354);
and UO_1112 (O_1112,N_17403,N_17069);
nand UO_1113 (O_1113,N_19747,N_16733);
nor UO_1114 (O_1114,N_19961,N_19666);
nor UO_1115 (O_1115,N_17006,N_18508);
and UO_1116 (O_1116,N_19414,N_18932);
or UO_1117 (O_1117,N_19081,N_18030);
nand UO_1118 (O_1118,N_17378,N_19065);
nand UO_1119 (O_1119,N_16709,N_17609);
and UO_1120 (O_1120,N_19042,N_17619);
nor UO_1121 (O_1121,N_15491,N_16360);
or UO_1122 (O_1122,N_17875,N_17079);
or UO_1123 (O_1123,N_17281,N_16083);
nor UO_1124 (O_1124,N_16783,N_15850);
nor UO_1125 (O_1125,N_18475,N_18602);
or UO_1126 (O_1126,N_18321,N_16204);
or UO_1127 (O_1127,N_15820,N_15455);
and UO_1128 (O_1128,N_16724,N_19470);
or UO_1129 (O_1129,N_16303,N_18084);
nand UO_1130 (O_1130,N_15106,N_17258);
and UO_1131 (O_1131,N_17970,N_18568);
nor UO_1132 (O_1132,N_16877,N_19598);
and UO_1133 (O_1133,N_16879,N_16736);
and UO_1134 (O_1134,N_16218,N_15855);
nor UO_1135 (O_1135,N_16665,N_15711);
or UO_1136 (O_1136,N_19879,N_17735);
or UO_1137 (O_1137,N_19375,N_19712);
and UO_1138 (O_1138,N_18558,N_18841);
nand UO_1139 (O_1139,N_17100,N_16273);
or UO_1140 (O_1140,N_19285,N_17940);
nor UO_1141 (O_1141,N_19095,N_16187);
nor UO_1142 (O_1142,N_19383,N_15563);
and UO_1143 (O_1143,N_19590,N_18356);
or UO_1144 (O_1144,N_15220,N_18544);
and UO_1145 (O_1145,N_16551,N_15700);
and UO_1146 (O_1146,N_15326,N_17029);
and UO_1147 (O_1147,N_19768,N_16745);
nor UO_1148 (O_1148,N_15984,N_15560);
and UO_1149 (O_1149,N_17899,N_18334);
xnor UO_1150 (O_1150,N_18990,N_17263);
nor UO_1151 (O_1151,N_16351,N_17672);
and UO_1152 (O_1152,N_16316,N_15874);
or UO_1153 (O_1153,N_16064,N_16077);
or UO_1154 (O_1154,N_19839,N_15910);
or UO_1155 (O_1155,N_16814,N_16109);
xnor UO_1156 (O_1156,N_16510,N_17321);
or UO_1157 (O_1157,N_16820,N_16459);
nor UO_1158 (O_1158,N_19258,N_15994);
or UO_1159 (O_1159,N_17357,N_16096);
nand UO_1160 (O_1160,N_16047,N_19510);
and UO_1161 (O_1161,N_15777,N_15807);
or UO_1162 (O_1162,N_18183,N_19149);
or UO_1163 (O_1163,N_18434,N_17815);
xnor UO_1164 (O_1164,N_19126,N_17825);
and UO_1165 (O_1165,N_16930,N_17887);
nand UO_1166 (O_1166,N_16327,N_19250);
or UO_1167 (O_1167,N_15211,N_18737);
or UO_1168 (O_1168,N_15546,N_18875);
and UO_1169 (O_1169,N_16000,N_16515);
nand UO_1170 (O_1170,N_15060,N_18689);
xor UO_1171 (O_1171,N_19077,N_18618);
or UO_1172 (O_1172,N_18311,N_15699);
or UO_1173 (O_1173,N_17268,N_19429);
or UO_1174 (O_1174,N_15514,N_17479);
nor UO_1175 (O_1175,N_15990,N_19161);
or UO_1176 (O_1176,N_17652,N_16176);
and UO_1177 (O_1177,N_19584,N_18750);
nand UO_1178 (O_1178,N_17388,N_17726);
nand UO_1179 (O_1179,N_15396,N_17496);
or UO_1180 (O_1180,N_16387,N_18516);
and UO_1181 (O_1181,N_19221,N_18188);
and UO_1182 (O_1182,N_16815,N_19810);
and UO_1183 (O_1183,N_19889,N_17719);
nand UO_1184 (O_1184,N_19431,N_19187);
or UO_1185 (O_1185,N_16819,N_18604);
or UO_1186 (O_1186,N_17628,N_17516);
and UO_1187 (O_1187,N_17064,N_15404);
or UO_1188 (O_1188,N_16516,N_15216);
nand UO_1189 (O_1189,N_15376,N_18545);
or UO_1190 (O_1190,N_18941,N_17313);
nor UO_1191 (O_1191,N_16286,N_19543);
xnor UO_1192 (O_1192,N_19875,N_18720);
and UO_1193 (O_1193,N_16337,N_15843);
nor UO_1194 (O_1194,N_15579,N_18979);
and UO_1195 (O_1195,N_18462,N_17315);
nor UO_1196 (O_1196,N_15609,N_18915);
or UO_1197 (O_1197,N_15971,N_16680);
nor UO_1198 (O_1198,N_15988,N_19928);
and UO_1199 (O_1199,N_16752,N_16652);
nor UO_1200 (O_1200,N_15552,N_18861);
nor UO_1201 (O_1201,N_18190,N_15365);
nand UO_1202 (O_1202,N_18626,N_17346);
or UO_1203 (O_1203,N_19881,N_17227);
or UO_1204 (O_1204,N_19860,N_18496);
and UO_1205 (O_1205,N_15758,N_19825);
nor UO_1206 (O_1206,N_18977,N_16512);
nand UO_1207 (O_1207,N_16493,N_16676);
and UO_1208 (O_1208,N_19751,N_19956);
and UO_1209 (O_1209,N_19643,N_19673);
or UO_1210 (O_1210,N_18991,N_18357);
nor UO_1211 (O_1211,N_15799,N_15793);
nor UO_1212 (O_1212,N_17911,N_15635);
nand UO_1213 (O_1213,N_18273,N_17751);
nand UO_1214 (O_1214,N_19008,N_15827);
nand UO_1215 (O_1215,N_15804,N_18829);
and UO_1216 (O_1216,N_16980,N_16997);
nand UO_1217 (O_1217,N_19544,N_19358);
or UO_1218 (O_1218,N_17341,N_19705);
nand UO_1219 (O_1219,N_17893,N_19038);
and UO_1220 (O_1220,N_19464,N_17747);
and UO_1221 (O_1221,N_16941,N_19138);
nand UO_1222 (O_1222,N_15275,N_15287);
nor UO_1223 (O_1223,N_15002,N_15100);
nand UO_1224 (O_1224,N_19239,N_18351);
xor UO_1225 (O_1225,N_19466,N_17380);
nand UO_1226 (O_1226,N_16835,N_18105);
and UO_1227 (O_1227,N_18962,N_17778);
nand UO_1228 (O_1228,N_17448,N_19050);
nor UO_1229 (O_1229,N_18237,N_16619);
nor UO_1230 (O_1230,N_19921,N_19625);
or UO_1231 (O_1231,N_17087,N_19577);
nor UO_1232 (O_1232,N_17756,N_16070);
or UO_1233 (O_1233,N_18384,N_17967);
nand UO_1234 (O_1234,N_15573,N_19151);
nand UO_1235 (O_1235,N_18396,N_17737);
or UO_1236 (O_1236,N_15101,N_16137);
nand UO_1237 (O_1237,N_19663,N_15636);
and UO_1238 (O_1238,N_17427,N_19144);
nor UO_1239 (O_1239,N_19183,N_19611);
xnor UO_1240 (O_1240,N_17352,N_18202);
and UO_1241 (O_1241,N_16039,N_18832);
or UO_1242 (O_1242,N_16263,N_18786);
nor UO_1243 (O_1243,N_16937,N_18343);
and UO_1244 (O_1244,N_16448,N_19275);
and UO_1245 (O_1245,N_19615,N_15965);
nand UO_1246 (O_1246,N_15200,N_17057);
or UO_1247 (O_1247,N_17990,N_19941);
nand UO_1248 (O_1248,N_16352,N_15118);
and UO_1249 (O_1249,N_18315,N_17334);
or UO_1250 (O_1250,N_16378,N_17177);
xor UO_1251 (O_1251,N_18800,N_17816);
nor UO_1252 (O_1252,N_19458,N_16385);
nor UO_1253 (O_1253,N_19854,N_17328);
or UO_1254 (O_1254,N_17186,N_18646);
nor UO_1255 (O_1255,N_16628,N_16729);
nand UO_1256 (O_1256,N_16148,N_19128);
or UO_1257 (O_1257,N_16027,N_18743);
nor UO_1258 (O_1258,N_17220,N_15682);
nand UO_1259 (O_1259,N_15130,N_15716);
and UO_1260 (O_1260,N_16209,N_16342);
or UO_1261 (O_1261,N_16058,N_16621);
and UO_1262 (O_1262,N_19465,N_16335);
nand UO_1263 (O_1263,N_16138,N_18271);
or UO_1264 (O_1264,N_18217,N_18371);
nand UO_1265 (O_1265,N_15351,N_16653);
and UO_1266 (O_1266,N_16289,N_15471);
or UO_1267 (O_1267,N_17246,N_16650);
nor UO_1268 (O_1268,N_19534,N_19292);
and UO_1269 (O_1269,N_15689,N_18436);
xor UO_1270 (O_1270,N_16728,N_16574);
nand UO_1271 (O_1271,N_15183,N_16177);
or UO_1272 (O_1272,N_18291,N_18425);
nor UO_1273 (O_1273,N_18929,N_19253);
or UO_1274 (O_1274,N_15705,N_17989);
nor UO_1275 (O_1275,N_18060,N_17553);
and UO_1276 (O_1276,N_18987,N_15603);
nand UO_1277 (O_1277,N_18293,N_19069);
and UO_1278 (O_1278,N_17622,N_15693);
or UO_1279 (O_1279,N_17494,N_16585);
nand UO_1280 (O_1280,N_18672,N_16453);
nand UO_1281 (O_1281,N_18122,N_19602);
or UO_1282 (O_1282,N_16054,N_17689);
and UO_1283 (O_1283,N_18444,N_17820);
nand UO_1284 (O_1284,N_19816,N_15442);
nand UO_1285 (O_1285,N_16694,N_15342);
nor UO_1286 (O_1286,N_19058,N_18075);
and UO_1287 (O_1287,N_19164,N_19461);
nor UO_1288 (O_1288,N_19983,N_18399);
and UO_1289 (O_1289,N_19262,N_16361);
nand UO_1290 (O_1290,N_17923,N_19331);
nor UO_1291 (O_1291,N_18102,N_19137);
nand UO_1292 (O_1292,N_19832,N_17317);
nor UO_1293 (O_1293,N_18714,N_17969);
nand UO_1294 (O_1294,N_18691,N_16708);
nand UO_1295 (O_1295,N_19391,N_18437);
and UO_1296 (O_1296,N_16831,N_19372);
nand UO_1297 (O_1297,N_18443,N_18501);
nor UO_1298 (O_1298,N_15125,N_18707);
and UO_1299 (O_1299,N_17704,N_17836);
or UO_1300 (O_1300,N_17338,N_15844);
nor UO_1301 (O_1301,N_19853,N_19680);
nand UO_1302 (O_1302,N_19195,N_18157);
nand UO_1303 (O_1303,N_17191,N_16359);
nor UO_1304 (O_1304,N_17493,N_17664);
and UO_1305 (O_1305,N_17487,N_17690);
nand UO_1306 (O_1306,N_17575,N_17722);
nor UO_1307 (O_1307,N_19539,N_19682);
nand UO_1308 (O_1308,N_18079,N_19480);
and UO_1309 (O_1309,N_19335,N_15269);
or UO_1310 (O_1310,N_18868,N_18045);
and UO_1311 (O_1311,N_19319,N_15678);
nor UO_1312 (O_1312,N_18966,N_17663);
and UO_1313 (O_1313,N_16528,N_19507);
and UO_1314 (O_1314,N_15298,N_16629);
xor UO_1315 (O_1315,N_19141,N_16905);
and UO_1316 (O_1316,N_15357,N_16685);
nor UO_1317 (O_1317,N_19797,N_15630);
nor UO_1318 (O_1318,N_17023,N_18866);
nor UO_1319 (O_1319,N_19784,N_17594);
and UO_1320 (O_1320,N_19658,N_17614);
or UO_1321 (O_1321,N_18151,N_17253);
nand UO_1322 (O_1322,N_16646,N_19931);
nor UO_1323 (O_1323,N_18239,N_17900);
and UO_1324 (O_1324,N_18671,N_18453);
nand UO_1325 (O_1325,N_18613,N_15555);
xor UO_1326 (O_1326,N_19233,N_15110);
xor UO_1327 (O_1327,N_17362,N_16237);
or UO_1328 (O_1328,N_19325,N_19482);
nor UO_1329 (O_1329,N_19932,N_19769);
nor UO_1330 (O_1330,N_18032,N_18809);
nor UO_1331 (O_1331,N_16473,N_15897);
and UO_1332 (O_1332,N_19017,N_16575);
nand UO_1333 (O_1333,N_15776,N_15970);
nand UO_1334 (O_1334,N_15489,N_17172);
or UO_1335 (O_1335,N_15520,N_17224);
or UO_1336 (O_1336,N_18583,N_18934);
and UO_1337 (O_1337,N_19289,N_17260);
nor UO_1338 (O_1338,N_15823,N_15929);
or UO_1339 (O_1339,N_18978,N_18494);
nor UO_1340 (O_1340,N_15597,N_17712);
nand UO_1341 (O_1341,N_18918,N_16117);
or UO_1342 (O_1342,N_17444,N_16490);
or UO_1343 (O_1343,N_19759,N_15032);
and UO_1344 (O_1344,N_17273,N_19872);
or UO_1345 (O_1345,N_16087,N_19977);
and UO_1346 (O_1346,N_19945,N_17925);
nor UO_1347 (O_1347,N_18820,N_18066);
nand UO_1348 (O_1348,N_17406,N_18971);
nand UO_1349 (O_1349,N_15084,N_18669);
and UO_1350 (O_1350,N_18913,N_18339);
or UO_1351 (O_1351,N_19163,N_15947);
and UO_1352 (O_1352,N_18507,N_18299);
or UO_1353 (O_1353,N_19843,N_19495);
or UO_1354 (O_1354,N_18428,N_16236);
or UO_1355 (O_1355,N_16861,N_17307);
or UO_1356 (O_1356,N_16249,N_16577);
or UO_1357 (O_1357,N_19742,N_19563);
xnor UO_1358 (O_1358,N_17390,N_18565);
or UO_1359 (O_1359,N_17708,N_19777);
or UO_1360 (O_1360,N_18928,N_15184);
nor UO_1361 (O_1361,N_16689,N_18362);
and UO_1362 (O_1362,N_18510,N_18346);
or UO_1363 (O_1363,N_18943,N_18469);
nor UO_1364 (O_1364,N_15190,N_16808);
and UO_1365 (O_1365,N_17847,N_17922);
xor UO_1366 (O_1366,N_18063,N_15841);
or UO_1367 (O_1367,N_17142,N_19189);
nand UO_1368 (O_1368,N_18958,N_17364);
or UO_1369 (O_1369,N_19146,N_18019);
nor UO_1370 (O_1370,N_18423,N_18282);
nand UO_1371 (O_1371,N_16390,N_15348);
and UO_1372 (O_1372,N_17890,N_17302);
or UO_1373 (O_1373,N_17345,N_16175);
nand UO_1374 (O_1374,N_18251,N_19731);
and UO_1375 (O_1375,N_18844,N_17370);
and UO_1376 (O_1376,N_15140,N_18192);
nand UO_1377 (O_1377,N_19549,N_18559);
nand UO_1378 (O_1378,N_15215,N_17783);
nor UO_1379 (O_1379,N_15166,N_17951);
nor UO_1380 (O_1380,N_19594,N_16214);
nor UO_1381 (O_1381,N_15139,N_17033);
nand UO_1382 (O_1382,N_19373,N_16095);
or UO_1383 (O_1383,N_18764,N_15569);
nand UO_1384 (O_1384,N_15323,N_16225);
nor UO_1385 (O_1385,N_16363,N_15664);
and UO_1386 (O_1386,N_17158,N_15356);
nor UO_1387 (O_1387,N_17291,N_19362);
or UO_1388 (O_1388,N_15079,N_16945);
or UO_1389 (O_1389,N_17449,N_15466);
nor UO_1390 (O_1390,N_15055,N_15016);
or UO_1391 (O_1391,N_16030,N_17091);
or UO_1392 (O_1392,N_15806,N_19526);
and UO_1393 (O_1393,N_18656,N_19720);
nand UO_1394 (O_1394,N_18896,N_19145);
nor UO_1395 (O_1395,N_19837,N_17938);
nand UO_1396 (O_1396,N_17074,N_18632);
and UO_1397 (O_1397,N_17248,N_16961);
or UO_1398 (O_1398,N_15372,N_15710);
and UO_1399 (O_1399,N_16857,N_19993);
nand UO_1400 (O_1400,N_15265,N_16350);
xnor UO_1401 (O_1401,N_19300,N_18518);
nand UO_1402 (O_1402,N_18973,N_15735);
nand UO_1403 (O_1403,N_17348,N_16557);
and UO_1404 (O_1404,N_16834,N_17592);
and UO_1405 (O_1405,N_18661,N_17853);
nand UO_1406 (O_1406,N_16136,N_17960);
nand UO_1407 (O_1407,N_15669,N_17551);
or UO_1408 (O_1408,N_17585,N_19197);
or UO_1409 (O_1409,N_17913,N_16474);
nor UO_1410 (O_1410,N_15156,N_15375);
or UO_1411 (O_1411,N_15677,N_15848);
and UO_1412 (O_1412,N_15864,N_18308);
nor UO_1413 (O_1413,N_19340,N_19489);
and UO_1414 (O_1414,N_16132,N_15822);
and UO_1415 (O_1415,N_19963,N_17245);
or UO_1416 (O_1416,N_17742,N_19715);
or UO_1417 (O_1417,N_19933,N_17176);
nor UO_1418 (O_1418,N_18858,N_18025);
and UO_1419 (O_1419,N_19001,N_18181);
nand UO_1420 (O_1420,N_18881,N_17838);
or UO_1421 (O_1421,N_17076,N_16711);
nor UO_1422 (O_1422,N_17405,N_16896);
nand UO_1423 (O_1423,N_19435,N_16353);
nand UO_1424 (O_1424,N_17536,N_19098);
and UO_1425 (O_1425,N_18006,N_15712);
or UO_1426 (O_1426,N_19515,N_18839);
and UO_1427 (O_1427,N_16224,N_17030);
and UO_1428 (O_1428,N_15460,N_15590);
and UO_1429 (O_1429,N_16002,N_15295);
or UO_1430 (O_1430,N_15767,N_16737);
nor UO_1431 (O_1431,N_16971,N_15612);
and UO_1432 (O_1432,N_16881,N_15279);
or UO_1433 (O_1433,N_16226,N_17864);
or UO_1434 (O_1434,N_18223,N_17734);
nand UO_1435 (O_1435,N_19883,N_18300);
nor UO_1436 (O_1436,N_19942,N_18053);
nor UO_1437 (O_1437,N_19210,N_16521);
or UO_1438 (O_1438,N_19142,N_19236);
nor UO_1439 (O_1439,N_19403,N_16414);
nand UO_1440 (O_1440,N_17443,N_16450);
nor UO_1441 (O_1441,N_19531,N_16916);
nor UO_1442 (O_1442,N_16530,N_15702);
or UO_1443 (O_1443,N_19554,N_19831);
and UO_1444 (O_1444,N_18369,N_17270);
nor UO_1445 (O_1445,N_16074,N_19927);
or UO_1446 (O_1446,N_19958,N_17717);
and UO_1447 (O_1447,N_18770,N_17359);
nand UO_1448 (O_1448,N_15192,N_16504);
and UO_1449 (O_1449,N_17826,N_16804);
nor UO_1450 (O_1450,N_17586,N_17851);
nor UO_1451 (O_1451,N_16247,N_16867);
or UO_1452 (O_1452,N_19882,N_19985);
and UO_1453 (O_1453,N_18289,N_16116);
nand UO_1454 (O_1454,N_15480,N_19010);
or UO_1455 (O_1455,N_15625,N_15981);
nand UO_1456 (O_1456,N_18378,N_18702);
or UO_1457 (O_1457,N_15172,N_19520);
nand UO_1458 (O_1458,N_19672,N_18044);
nor UO_1459 (O_1459,N_15486,N_16959);
xnor UO_1460 (O_1460,N_16659,N_17683);
nor UO_1461 (O_1461,N_19094,N_18921);
or UO_1462 (O_1462,N_18004,N_19453);
and UO_1463 (O_1463,N_19618,N_17880);
nor UO_1464 (O_1464,N_19783,N_15459);
nor UO_1465 (O_1465,N_17202,N_17514);
or UO_1466 (O_1466,N_19270,N_18294);
and UO_1467 (O_1467,N_19626,N_15085);
xor UO_1468 (O_1468,N_19623,N_15210);
nor UO_1469 (O_1469,N_17945,N_15504);
nor UO_1470 (O_1470,N_15743,N_18487);
nor UO_1471 (O_1471,N_17093,N_15694);
or UO_1472 (O_1472,N_15080,N_16613);
nand UO_1473 (O_1473,N_16532,N_19737);
nor UO_1474 (O_1474,N_16347,N_19648);
and UO_1475 (O_1475,N_15891,N_17457);
or UO_1476 (O_1476,N_15751,N_18685);
nand UO_1477 (O_1477,N_16207,N_17097);
nor UO_1478 (O_1478,N_15128,N_19361);
nand UO_1479 (O_1479,N_17159,N_16422);
nand UO_1480 (O_1480,N_16714,N_19350);
and UO_1481 (O_1481,N_17980,N_16216);
nor UO_1482 (O_1482,N_17181,N_16648);
and UO_1483 (O_1483,N_15082,N_17520);
and UO_1484 (O_1484,N_17324,N_17133);
nand UO_1485 (O_1485,N_18206,N_19438);
nor UO_1486 (O_1486,N_19456,N_15675);
nand UO_1487 (O_1487,N_19436,N_16365);
nand UO_1488 (O_1488,N_19736,N_18892);
nand UO_1489 (O_1489,N_15138,N_16992);
or UO_1490 (O_1490,N_16339,N_15304);
nand UO_1491 (O_1491,N_18847,N_18248);
nor UO_1492 (O_1492,N_16305,N_19118);
and UO_1493 (O_1493,N_15400,N_19724);
xnor UO_1494 (O_1494,N_17996,N_17121);
nand UO_1495 (O_1495,N_19269,N_16954);
and UO_1496 (O_1496,N_16238,N_17848);
or UO_1497 (O_1497,N_19169,N_19263);
nand UO_1498 (O_1498,N_17078,N_19647);
and UO_1499 (O_1499,N_18413,N_18531);
and UO_1500 (O_1500,N_16071,N_17732);
or UO_1501 (O_1501,N_18514,N_16456);
and UO_1502 (O_1502,N_18775,N_19503);
and UO_1503 (O_1503,N_18607,N_15629);
and UO_1504 (O_1504,N_17117,N_16529);
and UO_1505 (O_1505,N_18205,N_18768);
nand UO_1506 (O_1506,N_17739,N_17289);
nand UO_1507 (O_1507,N_16695,N_18476);
and UO_1508 (O_1508,N_18623,N_15102);
nand UO_1509 (O_1509,N_18326,N_17358);
and UO_1510 (O_1510,N_17927,N_18352);
or UO_1511 (O_1511,N_16157,N_19318);
or UO_1512 (O_1512,N_19542,N_15332);
nor UO_1513 (O_1513,N_19140,N_15205);
xor UO_1514 (O_1514,N_15112,N_16604);
nor UO_1515 (O_1515,N_18170,N_19744);
and UO_1516 (O_1516,N_15028,N_16304);
or UO_1517 (O_1517,N_19711,N_19474);
nor UO_1518 (O_1518,N_15483,N_16463);
nor UO_1519 (O_1519,N_15873,N_15149);
nor UO_1520 (O_1520,N_15997,N_17961);
or UO_1521 (O_1521,N_19207,N_15770);
or UO_1522 (O_1522,N_17112,N_19218);
xor UO_1523 (O_1523,N_17505,N_18288);
or UO_1524 (O_1524,N_15159,N_17813);
xor UO_1525 (O_1525,N_17802,N_16261);
nor UO_1526 (O_1526,N_18649,N_16968);
nor UO_1527 (O_1527,N_16041,N_18586);
or UO_1528 (O_1528,N_18166,N_18662);
nor UO_1529 (O_1529,N_15680,N_16257);
and UO_1530 (O_1530,N_18097,N_15109);
and UO_1531 (O_1531,N_16514,N_18960);
or UO_1532 (O_1532,N_15692,N_17762);
nand UO_1533 (O_1533,N_18981,N_18761);
and UO_1534 (O_1534,N_16563,N_18880);
nor UO_1535 (O_1535,N_16189,N_15256);
nand UO_1536 (O_1536,N_18391,N_17241);
and UO_1537 (O_1537,N_17994,N_18038);
and UO_1538 (O_1538,N_19685,N_17503);
and UO_1539 (O_1539,N_18325,N_19317);
or UO_1540 (O_1540,N_17065,N_16310);
or UO_1541 (O_1541,N_17795,N_19406);
or UO_1542 (O_1542,N_16364,N_18859);
xor UO_1543 (O_1543,N_19586,N_16826);
nor UO_1544 (O_1544,N_16878,N_17417);
or UO_1545 (O_1545,N_18647,N_18620);
nand UO_1546 (O_1546,N_15264,N_17089);
and UO_1547 (O_1547,N_15121,N_18779);
and UO_1548 (O_1548,N_19346,N_16637);
nand UO_1549 (O_1549,N_19849,N_18249);
and UO_1550 (O_1550,N_19394,N_18358);
nor UO_1551 (O_1551,N_17440,N_17128);
and UO_1552 (O_1552,N_15380,N_18944);
nor UO_1553 (O_1553,N_16884,N_17855);
and UO_1554 (O_1554,N_19698,N_15914);
nor UO_1555 (O_1555,N_16172,N_16851);
nand UO_1556 (O_1556,N_19671,N_15683);
or UO_1557 (O_1557,N_19924,N_17697);
nor UO_1558 (O_1558,N_16764,N_18812);
or UO_1559 (O_1559,N_15364,N_18986);
nor UO_1560 (O_1560,N_18570,N_19478);
and UO_1561 (O_1561,N_19808,N_19999);
nor UO_1562 (O_1562,N_16712,N_15996);
nor UO_1563 (O_1563,N_17674,N_16379);
nand UO_1564 (O_1564,N_16969,N_16800);
and UO_1565 (O_1565,N_18129,N_18056);
nor UO_1566 (O_1566,N_19957,N_15909);
nand UO_1567 (O_1567,N_18540,N_16014);
and UO_1568 (O_1568,N_15619,N_19440);
and UO_1569 (O_1569,N_16325,N_18193);
nand UO_1570 (O_1570,N_15473,N_17454);
nor UO_1571 (O_1571,N_16756,N_15643);
or UO_1572 (O_1572,N_19213,N_17415);
and UO_1573 (O_1573,N_15511,N_17665);
nor UO_1574 (O_1574,N_16993,N_18908);
and UO_1575 (O_1575,N_16890,N_17545);
nand UO_1576 (O_1576,N_18995,N_17275);
nor UO_1577 (O_1577,N_17486,N_17231);
or UO_1578 (O_1578,N_19548,N_19360);
or UO_1579 (O_1579,N_17125,N_15044);
or UO_1580 (O_1580,N_19833,N_16464);
nand UO_1581 (O_1581,N_18560,N_18945);
nand UO_1582 (O_1582,N_15885,N_17766);
and UO_1583 (O_1583,N_18201,N_19738);
nand UO_1584 (O_1584,N_15649,N_19987);
nor UO_1585 (O_1585,N_16538,N_15769);
nor UO_1586 (O_1586,N_15880,N_19003);
xnor UO_1587 (O_1587,N_16874,N_19687);
or UO_1588 (O_1588,N_17538,N_17337);
or UO_1589 (O_1589,N_15755,N_17480);
nor UO_1590 (O_1590,N_17168,N_19472);
or UO_1591 (O_1591,N_16942,N_16198);
nand UO_1592 (O_1592,N_15684,N_19966);
and UO_1593 (O_1593,N_18014,N_15157);
or UO_1594 (O_1594,N_15168,N_16987);
nand UO_1595 (O_1595,N_16565,N_18270);
nor UO_1596 (O_1596,N_19108,N_19234);
nor UO_1597 (O_1597,N_15857,N_15450);
nand UO_1598 (O_1598,N_19589,N_19176);
nor UO_1599 (O_1599,N_16885,N_17721);
and UO_1600 (O_1600,N_15688,N_19057);
or UO_1601 (O_1601,N_16895,N_18460);
and UO_1602 (O_1602,N_17373,N_19007);
nand UO_1603 (O_1603,N_18533,N_17210);
nor UO_1604 (O_1604,N_17422,N_17419);
and UO_1605 (O_1605,N_15004,N_19093);
nor UO_1606 (O_1606,N_15889,N_17653);
or UO_1607 (O_1607,N_19185,N_18529);
nand UO_1608 (O_1608,N_18161,N_18268);
nor UO_1609 (O_1609,N_16562,N_16168);
nor UO_1610 (O_1610,N_16955,N_15798);
nor UO_1611 (O_1611,N_15503,N_16159);
and UO_1612 (O_1612,N_18445,N_18906);
or UO_1613 (O_1613,N_18323,N_15041);
xor UO_1614 (O_1614,N_19855,N_16943);
and UO_1615 (O_1615,N_17746,N_18952);
nand UO_1616 (O_1616,N_16771,N_19370);
nor UO_1617 (O_1617,N_18863,N_16765);
nand UO_1618 (O_1618,N_19012,N_19522);
and UO_1619 (O_1619,N_19686,N_16903);
nor UO_1620 (O_1620,N_18699,N_17599);
and UO_1621 (O_1621,N_18769,N_16076);
and UO_1622 (O_1622,N_18655,N_18338);
nor UO_1623 (O_1623,N_17995,N_18633);
and UO_1624 (O_1624,N_19157,N_15553);
nor UO_1625 (O_1625,N_17885,N_19481);
nor UO_1626 (O_1626,N_17559,N_15732);
nand UO_1627 (O_1627,N_17481,N_18564);
nand UO_1628 (O_1628,N_17379,N_16092);
and UO_1629 (O_1629,N_18280,N_15444);
nand UO_1630 (O_1630,N_16150,N_18452);
and UO_1631 (O_1631,N_17482,N_16535);
nor UO_1632 (O_1632,N_15007,N_15907);
nand UO_1633 (O_1633,N_15618,N_15626);
nand UO_1634 (O_1634,N_18337,N_19654);
and UO_1635 (O_1635,N_18488,N_17643);
and UO_1636 (O_1636,N_16036,N_16744);
and UO_1637 (O_1637,N_16524,N_18596);
or UO_1638 (O_1638,N_19823,N_15706);
or UO_1639 (O_1639,N_19308,N_18826);
or UO_1640 (O_1640,N_16271,N_15734);
and UO_1641 (O_1641,N_15814,N_16201);
nor UO_1642 (O_1642,N_18733,N_18442);
and UO_1643 (O_1643,N_16190,N_16410);
nor UO_1644 (O_1644,N_16806,N_15449);
and UO_1645 (O_1645,N_19422,N_16666);
or UO_1646 (O_1646,N_18798,N_15230);
and UO_1647 (O_1647,N_18942,N_19492);
and UO_1648 (O_1648,N_18301,N_15754);
nor UO_1649 (O_1649,N_17235,N_16571);
nor UO_1650 (O_1650,N_18601,N_18393);
nand UO_1651 (O_1651,N_18076,N_17189);
nor UO_1652 (O_1652,N_18789,N_16417);
or UO_1653 (O_1653,N_18092,N_17182);
and UO_1654 (O_1654,N_15354,N_17579);
nand UO_1655 (O_1655,N_18914,N_15013);
or UO_1656 (O_1656,N_19181,N_17723);
nand UO_1657 (O_1657,N_15235,N_16056);
and UO_1658 (O_1658,N_17420,N_19248);
or UO_1659 (O_1659,N_17262,N_19708);
and UO_1660 (O_1660,N_15652,N_16741);
or UO_1661 (O_1661,N_15507,N_16500);
or UO_1662 (O_1662,N_17354,N_16914);
nand UO_1663 (O_1663,N_17624,N_15244);
nand UO_1664 (O_1664,N_15418,N_19745);
or UO_1665 (O_1665,N_16759,N_16082);
and UO_1666 (O_1666,N_15011,N_15512);
xor UO_1667 (O_1667,N_16398,N_17965);
nand UO_1668 (O_1668,N_19467,N_19002);
nand UO_1669 (O_1669,N_19509,N_19244);
nand UO_1670 (O_1670,N_18427,N_18107);
nand UO_1671 (O_1671,N_19423,N_18208);
or UO_1672 (O_1672,N_17912,N_18468);
nor UO_1673 (O_1673,N_16622,N_15585);
and UO_1674 (O_1674,N_15952,N_16140);
nor UO_1675 (O_1675,N_18016,N_18933);
nand UO_1676 (O_1676,N_17544,N_17234);
and UO_1677 (O_1677,N_17681,N_18663);
nor UO_1678 (O_1678,N_18068,N_17455);
or UO_1679 (O_1679,N_17401,N_15036);
and UO_1680 (O_1680,N_17277,N_17059);
nand UO_1681 (O_1681,N_19089,N_18482);
or UO_1682 (O_1682,N_19877,N_15097);
nand UO_1683 (O_1683,N_17398,N_19938);
nor UO_1684 (O_1684,N_16766,N_17693);
nor UO_1685 (O_1685,N_18143,N_18642);
nor UO_1686 (O_1686,N_18900,N_18781);
nand UO_1687 (O_1687,N_16902,N_16721);
or UO_1688 (O_1688,N_18635,N_18571);
and UO_1689 (O_1689,N_17694,N_19177);
or UO_1690 (O_1690,N_17205,N_17801);
or UO_1691 (O_1691,N_15448,N_15745);
nor UO_1692 (O_1692,N_17977,N_16810);
nand UO_1693 (O_1693,N_17576,N_16050);
nand UO_1694 (O_1694,N_18473,N_19175);
and UO_1695 (O_1695,N_17525,N_19701);
or UO_1696 (O_1696,N_16979,N_19920);
nand UO_1697 (O_1697,N_17978,N_17648);
nor UO_1698 (O_1698,N_18619,N_19619);
nor UO_1699 (O_1699,N_16518,N_19629);
nor UO_1700 (O_1700,N_15817,N_17192);
nor UO_1701 (O_1701,N_19409,N_18615);
and UO_1702 (O_1702,N_17295,N_18790);
nand UO_1703 (O_1703,N_17548,N_16702);
or UO_1704 (O_1704,N_18340,N_18592);
nor UO_1705 (O_1705,N_17190,N_15231);
nand UO_1706 (O_1706,N_16020,N_18637);
xor UO_1707 (O_1707,N_16720,N_17251);
and UO_1708 (O_1708,N_17369,N_18250);
nor UO_1709 (O_1709,N_18010,N_17916);
and UO_1710 (O_1710,N_17048,N_18048);
nor UO_1711 (O_1711,N_15262,N_17498);
or UO_1712 (O_1712,N_17290,N_16651);
nor UO_1713 (O_1713,N_18985,N_16578);
or UO_1714 (O_1714,N_18432,N_15992);
and UO_1715 (O_1715,N_16123,N_15267);
nand UO_1716 (O_1716,N_16660,N_15198);
or UO_1717 (O_1717,N_16395,N_15207);
nand UO_1718 (O_1718,N_18071,N_18467);
or UO_1719 (O_1719,N_16217,N_18454);
xor UO_1720 (O_1720,N_15941,N_16307);
nor UO_1721 (O_1721,N_19230,N_15781);
nand UO_1722 (O_1722,N_18034,N_17200);
or UO_1723 (O_1723,N_19508,N_15878);
and UO_1724 (O_1724,N_19073,N_19865);
or UO_1725 (O_1725,N_15488,N_17876);
or UO_1726 (O_1726,N_15651,N_15982);
nor UO_1727 (O_1727,N_19743,N_15074);
or UO_1728 (O_1728,N_15131,N_19667);
or UO_1729 (O_1729,N_19015,N_16389);
nor UO_1730 (O_1730,N_19190,N_15939);
nand UO_1731 (O_1731,N_18441,N_16369);
or UO_1732 (O_1732,N_16549,N_15274);
nor UO_1733 (O_1733,N_19039,N_16016);
nor UO_1734 (O_1734,N_15308,N_19298);
nand UO_1735 (O_1735,N_15039,N_19801);
and UO_1736 (O_1736,N_17867,N_15343);
or UO_1737 (O_1737,N_15587,N_17670);
or UO_1738 (O_1738,N_18652,N_17868);
and UO_1739 (O_1739,N_16472,N_18774);
nor UO_1740 (O_1740,N_15033,N_15379);
or UO_1741 (O_1741,N_16154,N_16268);
nand UO_1742 (O_1742,N_17593,N_19923);
nor UO_1743 (O_1743,N_18999,N_17908);
nor UO_1744 (O_1744,N_16007,N_18538);
nor UO_1745 (O_1745,N_17926,N_18394);
nand UO_1746 (O_1746,N_15591,N_19628);
nor UO_1747 (O_1747,N_19498,N_15395);
nor UO_1748 (O_1748,N_19614,N_15930);
and UO_1749 (O_1749,N_15825,N_15432);
nand UO_1750 (O_1750,N_17621,N_15566);
and UO_1751 (O_1751,N_18499,N_18370);
nor UO_1752 (O_1752,N_15938,N_17122);
and UO_1753 (O_1753,N_15915,N_16595);
and UO_1754 (O_1754,N_15944,N_18225);
nand UO_1755 (O_1755,N_18569,N_15554);
and UO_1756 (O_1756,N_15852,N_17763);
nand UO_1757 (O_1757,N_16809,N_17882);
and UO_1758 (O_1758,N_18766,N_15311);
nand UO_1759 (O_1759,N_16886,N_16731);
nand UO_1760 (O_1760,N_19656,N_18519);
nand UO_1761 (O_1761,N_17703,N_15589);
nor UO_1762 (O_1762,N_18555,N_19699);
and UO_1763 (O_1763,N_17888,N_17617);
and UO_1764 (O_1764,N_15195,N_16649);
and UO_1765 (O_1765,N_16069,N_19344);
nor UO_1766 (O_1766,N_15439,N_18426);
or UO_1767 (O_1767,N_19863,N_17748);
nor UO_1768 (O_1768,N_15656,N_17523);
nor UO_1769 (O_1769,N_17955,N_15003);
nand UO_1770 (O_1770,N_15479,N_19048);
or UO_1771 (O_1771,N_16297,N_17827);
xnor UO_1772 (O_1772,N_15038,N_15556);
and UO_1773 (O_1773,N_18121,N_15613);
or UO_1774 (O_1774,N_19226,N_18925);
nor UO_1775 (O_1775,N_19802,N_16112);
or UO_1776 (O_1776,N_15610,N_17669);
nand UO_1777 (O_1777,N_17221,N_16868);
or UO_1778 (O_1778,N_16977,N_18093);
and UO_1779 (O_1779,N_17833,N_17461);
nand UO_1780 (O_1780,N_19903,N_16926);
nor UO_1781 (O_1781,N_15257,N_18606);
nor UO_1782 (O_1782,N_15752,N_17504);
nor UO_1783 (O_1783,N_17086,N_19645);
and UO_1784 (O_1784,N_19606,N_19929);
nand UO_1785 (O_1785,N_15143,N_16789);
nand UO_1786 (O_1786,N_15570,N_18359);
nor UO_1787 (O_1787,N_16210,N_16088);
nor UO_1788 (O_1788,N_16763,N_15881);
nor UO_1789 (O_1789,N_17971,N_16713);
or UO_1790 (O_1790,N_17312,N_18732);
nor UO_1791 (O_1791,N_19311,N_17240);
or UO_1792 (O_1792,N_18721,N_17953);
nand UO_1793 (O_1793,N_15592,N_19129);
or UO_1794 (O_1794,N_19293,N_16503);
nor UO_1795 (O_1795,N_17812,N_15882);
nand UO_1796 (O_1796,N_19086,N_16336);
nand UO_1797 (O_1797,N_19820,N_16743);
or UO_1798 (O_1798,N_16568,N_16328);
or UO_1799 (O_1799,N_17724,N_17080);
nand UO_1800 (O_1800,N_17612,N_15236);
and UO_1801 (O_1801,N_15803,N_16392);
nor UO_1802 (O_1802,N_16376,N_18957);
xor UO_1803 (O_1803,N_15648,N_15324);
nand UO_1804 (O_1804,N_18015,N_16645);
and UO_1805 (O_1805,N_19479,N_16793);
nand UO_1806 (O_1806,N_17499,N_15470);
or UO_1807 (O_1807,N_19760,N_17770);
nor UO_1808 (O_1808,N_18215,N_15374);
and UO_1809 (O_1809,N_19416,N_19473);
or UO_1810 (O_1810,N_19919,N_19962);
or UO_1811 (O_1811,N_17463,N_16608);
and UO_1812 (O_1812,N_15545,N_17414);
nand UO_1813 (O_1813,N_16491,N_17001);
and UO_1814 (O_1814,N_19337,N_18409);
nor UO_1815 (O_1815,N_18882,N_17700);
nor UO_1816 (O_1816,N_16974,N_17305);
nor UO_1817 (O_1817,N_18098,N_18255);
nand UO_1818 (O_1818,N_15388,N_17003);
nor UO_1819 (O_1819,N_16044,N_18599);
or UO_1820 (O_1820,N_18975,N_15792);
nor UO_1821 (O_1821,N_15725,N_15586);
or UO_1822 (O_1822,N_15302,N_19131);
and UO_1823 (O_1823,N_16582,N_19324);
or UO_1824 (O_1824,N_19404,N_19446);
or UO_1825 (O_1825,N_18690,N_16165);
and UO_1826 (O_1826,N_16230,N_15187);
nor UO_1827 (O_1827,N_18278,N_15451);
nand UO_1828 (O_1828,N_18810,N_18414);
nand UO_1829 (O_1829,N_19333,N_17906);
and UO_1830 (O_1830,N_15987,N_15926);
nor UO_1831 (O_1831,N_18860,N_15456);
and UO_1832 (O_1832,N_15186,N_16606);
or UO_1833 (O_1833,N_16697,N_15225);
nand UO_1834 (O_1834,N_15040,N_19476);
and UO_1835 (O_1835,N_19102,N_15847);
nand UO_1836 (O_1836,N_15795,N_17206);
or UO_1837 (O_1837,N_17527,N_15329);
or UO_1838 (O_1838,N_16331,N_16451);
nand UO_1839 (O_1839,N_17070,N_18657);
nand UO_1840 (O_1840,N_16416,N_17185);
nand UO_1841 (O_1841,N_19045,N_18883);
or UO_1842 (O_1842,N_17679,N_19080);
nor UO_1843 (O_1843,N_15313,N_16295);
or UO_1844 (O_1844,N_17705,N_15790);
and UO_1845 (O_1845,N_17162,N_18275);
or UO_1846 (O_1846,N_18794,N_17460);
and UO_1847 (O_1847,N_16040,N_16255);
nor UO_1848 (O_1848,N_17837,N_15527);
nor UO_1849 (O_1849,N_17314,N_18385);
nor UO_1850 (O_1850,N_18989,N_19451);
nor UO_1851 (O_1851,N_15582,N_19224);
nand UO_1852 (O_1852,N_18196,N_17298);
nor UO_1853 (O_1853,N_17438,N_15496);
and UO_1854 (O_1854,N_19583,N_18265);
nand UO_1855 (O_1855,N_19426,N_15402);
and UO_1856 (O_1856,N_19246,N_17502);
or UO_1857 (O_1857,N_17524,N_15296);
or UO_1858 (O_1858,N_17017,N_17765);
nor UO_1859 (O_1859,N_17591,N_15913);
nand UO_1860 (O_1860,N_17676,N_19791);
or UO_1861 (O_1861,N_16842,N_18722);
and UO_1862 (O_1862,N_19622,N_18948);
nor UO_1863 (O_1863,N_16706,N_17311);
and UO_1864 (O_1864,N_16638,N_19965);
nor UO_1865 (O_1865,N_16382,N_15490);
or UO_1866 (O_1866,N_15142,N_19208);
nor UO_1867 (O_1867,N_15098,N_17288);
nand UO_1868 (O_1868,N_19749,N_18830);
nor UO_1869 (O_1869,N_19040,N_18493);
nand UO_1870 (O_1870,N_15925,N_19912);
or UO_1871 (O_1871,N_19320,N_17881);
and UO_1872 (O_1872,N_15991,N_18461);
nand UO_1873 (O_1873,N_18213,N_17335);
or UO_1874 (O_1874,N_17814,N_19702);
or UO_1875 (O_1875,N_15927,N_19147);
or UO_1876 (O_1876,N_15482,N_17442);
nand UO_1877 (O_1877,N_19873,N_18226);
and UO_1878 (O_1878,N_15859,N_18257);
xor UO_1879 (O_1879,N_16219,N_18698);
and UO_1880 (O_1880,N_18713,N_19661);
nand UO_1881 (O_1881,N_17754,N_17374);
and UO_1882 (O_1882,N_15359,N_16065);
nand UO_1883 (O_1883,N_19171,N_18354);
and UO_1884 (O_1884,N_15224,N_19908);
and UO_1885 (O_1885,N_16153,N_15801);
nor UO_1886 (O_1886,N_18905,N_15087);
nor UO_1887 (O_1887,N_19678,N_18711);
nor UO_1888 (O_1888,N_16435,N_19103);
nand UO_1889 (O_1889,N_16372,N_17287);
and UO_1890 (O_1890,N_15266,N_19970);
nor UO_1891 (O_1891,N_19178,N_17716);
nand UO_1892 (O_1892,N_18089,N_17506);
and UO_1893 (O_1893,N_19284,N_18146);
nor UO_1894 (O_1894,N_19314,N_16849);
or UO_1895 (O_1895,N_18125,N_18020);
or UO_1896 (O_1896,N_19305,N_18263);
or UO_1897 (O_1897,N_15962,N_19867);
or UO_1898 (O_1898,N_17286,N_19752);
nor UO_1899 (O_1899,N_16292,N_17939);
nand UO_1900 (O_1900,N_19528,N_16428);
or UO_1901 (O_1901,N_19395,N_15180);
or UO_1902 (O_1902,N_18176,N_16746);
nor UO_1903 (O_1903,N_19165,N_15347);
or UO_1904 (O_1904,N_19068,N_18996);
or UO_1905 (O_1905,N_16111,N_16299);
nand UO_1906 (O_1906,N_17272,N_15851);
and UO_1907 (O_1907,N_18117,N_18349);
or UO_1908 (O_1908,N_19788,N_16986);
nand UO_1909 (O_1909,N_16950,N_15715);
or UO_1910 (O_1910,N_16862,N_17711);
or UO_1911 (O_1911,N_16281,N_15335);
xnor UO_1912 (O_1912,N_18403,N_17107);
and UO_1913 (O_1913,N_18203,N_19261);
nor UO_1914 (O_1914,N_19886,N_15369);
nand UO_1915 (O_1915,N_17333,N_19225);
and UO_1916 (O_1916,N_15708,N_17226);
and UO_1917 (O_1917,N_19143,N_19851);
or UO_1918 (O_1918,N_17095,N_16655);
nand UO_1919 (O_1919,N_15670,N_18187);
nand UO_1920 (O_1920,N_16046,N_15946);
nor UO_1921 (O_1921,N_16547,N_19556);
or UO_1922 (O_1922,N_17157,N_16981);
or UO_1923 (O_1923,N_19341,N_18575);
or UO_1924 (O_1924,N_16542,N_15382);
nor UO_1925 (O_1925,N_17891,N_16509);
nand UO_1926 (O_1926,N_18446,N_17919);
and UO_1927 (O_1927,N_19778,N_15019);
nor UO_1928 (O_1928,N_16309,N_19940);
and UO_1929 (O_1929,N_15942,N_19427);
nor UO_1930 (O_1930,N_19342,N_17635);
and UO_1931 (O_1931,N_16901,N_15608);
and UO_1932 (O_1932,N_18279,N_19842);
and UO_1933 (O_1933,N_15565,N_15193);
xor UO_1934 (O_1934,N_19603,N_18726);
or UO_1935 (O_1935,N_19282,N_16978);
or UO_1936 (O_1936,N_18485,N_16859);
nand UO_1937 (O_1937,N_17956,N_15564);
or UO_1938 (O_1938,N_16427,N_18333);
and UO_1939 (O_1939,N_18480,N_15615);
or UO_1940 (O_1940,N_17028,N_18155);
and UO_1941 (O_1941,N_17473,N_15259);
nand UO_1942 (O_1942,N_17018,N_17794);
nand UO_1943 (O_1943,N_15943,N_15742);
or UO_1944 (O_1944,N_18532,N_17824);
nor UO_1945 (O_1945,N_19052,N_15144);
and UO_1946 (O_1946,N_17453,N_16602);
or UO_1947 (O_1947,N_19047,N_16447);
or UO_1948 (O_1948,N_17509,N_16705);
nand UO_1949 (O_1949,N_15017,N_15337);
nor UO_1950 (O_1950,N_18238,N_16241);
nor UO_1951 (O_1951,N_15920,N_15870);
nor UO_1952 (O_1952,N_18353,N_17171);
or UO_1953 (O_1953,N_17793,N_17924);
or UO_1954 (O_1954,N_18778,N_19352);
nor UO_1955 (O_1955,N_16051,N_19150);
and UO_1956 (O_1956,N_19571,N_15727);
nor UO_1957 (O_1957,N_15604,N_19828);
or UO_1958 (O_1958,N_15458,N_16522);
xor UO_1959 (O_1959,N_15124,N_17229);
nor UO_1960 (O_1960,N_16558,N_17060);
or UO_1961 (O_1961,N_15919,N_15371);
nor UO_1962 (O_1962,N_19339,N_16028);
nand UO_1963 (O_1963,N_15830,N_19455);
nand UO_1964 (O_1964,N_16707,N_18851);
nor UO_1965 (O_1965,N_16674,N_18924);
or UO_1966 (O_1966,N_17519,N_18440);
and UO_1967 (O_1967,N_16229,N_15903);
and UO_1968 (O_1968,N_19916,N_16777);
and UO_1969 (O_1969,N_15188,N_19071);
nor UO_1970 (O_1970,N_17725,N_18209);
nor UO_1971 (O_1971,N_19376,N_18682);
nand UO_1972 (O_1972,N_19725,N_16821);
or UO_1973 (O_1973,N_19739,N_15330);
and UO_1974 (O_1974,N_16211,N_17002);
and UO_1975 (O_1975,N_18530,N_15253);
nand UO_1976 (O_1976,N_17047,N_18727);
nand UO_1977 (O_1977,N_18073,N_18640);
nand UO_1978 (O_1978,N_15794,N_19390);
and UO_1979 (O_1979,N_19312,N_16419);
nor UO_1980 (O_1980,N_19512,N_18043);
or UO_1981 (O_1981,N_19829,N_17946);
nand UO_1982 (O_1982,N_19132,N_17896);
and UO_1983 (O_1983,N_18676,N_17950);
nor UO_1984 (O_1984,N_15534,N_18684);
nor UO_1985 (O_1985,N_18404,N_18199);
nor UO_1986 (O_1986,N_16837,N_16643);
nor UO_1987 (O_1987,N_18112,N_16149);
nand UO_1988 (O_1988,N_17997,N_18783);
nand UO_1989 (O_1989,N_19527,N_15494);
nor UO_1990 (O_1990,N_16275,N_16033);
or UO_1991 (O_1991,N_19637,N_16960);
xnor UO_1992 (O_1992,N_18611,N_17727);
or UO_1993 (O_1993,N_16593,N_16484);
or UO_1994 (O_1994,N_19662,N_19400);
or UO_1995 (O_1995,N_19896,N_18090);
nor UO_1996 (O_1996,N_15729,N_16223);
nand UO_1997 (O_1997,N_15025,N_19084);
and UO_1998 (O_1998,N_17601,N_19726);
nand UO_1999 (O_1999,N_17204,N_16081);
nand UO_2000 (O_2000,N_15477,N_19365);
nand UO_2001 (O_2001,N_18096,N_17807);
or UO_2002 (O_2002,N_19016,N_16920);
nand UO_2003 (O_2003,N_18316,N_18845);
and UO_2004 (O_2004,N_19110,N_15089);
nor UO_2005 (O_2005,N_17974,N_16330);
or UO_2006 (O_2006,N_15390,N_15022);
nand UO_2007 (O_2007,N_15419,N_16144);
nor UO_2008 (O_2008,N_17353,N_15739);
or UO_2009 (O_2009,N_17430,N_18160);
or UO_2010 (O_2010,N_19114,N_17120);
nor UO_2011 (O_2011,N_18191,N_18159);
nor UO_2012 (O_2012,N_19815,N_17395);
and UO_2013 (O_2013,N_17831,N_16502);
and UO_2014 (O_2014,N_15853,N_15024);
and UO_2015 (O_2015,N_17686,N_19326);
or UO_2016 (O_2016,N_19356,N_18365);
nand UO_2017 (O_2017,N_15164,N_16918);
and UO_2018 (O_2018,N_19898,N_19064);
nand UO_2019 (O_2019,N_18492,N_19612);
and UO_2020 (O_2020,N_17488,N_19722);
or UO_2021 (O_2021,N_19948,N_15446);
nor UO_2022 (O_2022,N_16581,N_18150);
nand UO_2023 (O_2023,N_18285,N_16080);
or UO_2024 (O_2024,N_18753,N_15199);
nand UO_2025 (O_2025,N_15426,N_17584);
nand UO_2026 (O_2026,N_19486,N_19160);
and UO_2027 (O_2027,N_19256,N_17139);
or UO_2028 (O_2028,N_16401,N_17386);
nor UO_2029 (O_2029,N_17416,N_18644);
nand UO_2030 (O_2030,N_19025,N_19982);
and UO_2031 (O_2031,N_16075,N_17019);
and UO_2032 (O_2032,N_17037,N_18793);
or UO_2033 (O_2033,N_17852,N_18525);
nand UO_2034 (O_2034,N_15580,N_19133);
xnor UO_2035 (O_2035,N_19677,N_19729);
nor UO_2036 (O_2036,N_16541,N_15730);
or UO_2037 (O_2037,N_18069,N_18680);
and UO_2038 (O_2038,N_19034,N_18949);
or UO_2039 (O_2039,N_16034,N_17753);
and UO_2040 (O_2040,N_18197,N_19601);
nor UO_2041 (O_2041,N_19761,N_17526);
and UO_2042 (O_2042,N_16259,N_17173);
or UO_2043 (O_2043,N_16829,N_15163);
nand UO_2044 (O_2044,N_19041,N_19252);
nand UO_2045 (O_2045,N_17917,N_19056);
nand UO_2046 (O_2046,N_16824,N_16284);
or UO_2047 (O_2047,N_16761,N_18520);
and UO_2048 (O_2048,N_15173,N_19268);
and UO_2049 (O_2049,N_18498,N_17522);
nor UO_2050 (O_2050,N_17407,N_16306);
nand UO_2051 (O_2051,N_16042,N_17743);
and UO_2052 (O_2052,N_19483,N_17866);
nor UO_2053 (O_2053,N_16396,N_19792);
nand UO_2054 (O_2054,N_19632,N_19220);
nand UO_2055 (O_2055,N_16838,N_16313);
nand UO_2056 (O_2056,N_16162,N_16437);
nor UO_2057 (O_2057,N_17657,N_15966);
nor UO_2058 (O_2058,N_15277,N_19773);
or UO_2059 (O_2059,N_15151,N_18854);
nand UO_2060 (O_2060,N_15434,N_18276);
or UO_2061 (O_2061,N_19348,N_16195);
and UO_2062 (O_2062,N_17131,N_16682);
nor UO_2063 (O_2063,N_19154,N_17631);
or UO_2064 (O_2064,N_15787,N_16426);
or UO_2065 (O_2065,N_16854,N_19254);
nand UO_2066 (O_2066,N_17301,N_17381);
nand UO_2067 (O_2067,N_17402,N_18431);
nor UO_2068 (O_2068,N_15783,N_18094);
or UO_2069 (O_2069,N_16795,N_16462);
or UO_2070 (O_2070,N_18536,N_19223);
nand UO_2071 (O_2071,N_19386,N_15042);
and UO_2072 (O_2072,N_16929,N_17119);
nor UO_2073 (O_2073,N_16760,N_18186);
or UO_2074 (O_2074,N_18846,N_17564);
and UO_2075 (O_2075,N_18762,N_16206);
nand UO_2076 (O_2076,N_18537,N_19580);
or UO_2077 (O_2077,N_18156,N_18504);
nand UO_2078 (O_2078,N_16001,N_19890);
and UO_2079 (O_2079,N_16403,N_18231);
xnor UO_2080 (O_2080,N_18527,N_16010);
nor UO_2081 (O_2081,N_17036,N_16274);
or UO_2082 (O_2082,N_15691,N_15854);
or UO_2083 (O_2083,N_18042,N_17849);
or UO_2084 (O_2084,N_19355,N_15605);
nor UO_2085 (O_2085,N_17015,N_19382);
or UO_2086 (O_2086,N_16865,N_17127);
and UO_2087 (O_2087,N_15543,N_18910);
nand UO_2088 (O_2088,N_16233,N_17278);
and UO_2089 (O_2089,N_19665,N_16294);
or UO_2090 (O_2090,N_18701,N_15999);
nand UO_2091 (O_2091,N_15217,N_18367);
and UO_2092 (O_2092,N_18912,N_19821);
and UO_2093 (O_2093,N_16882,N_17775);
and UO_2094 (O_2094,N_16661,N_18017);
nor UO_2095 (O_2095,N_17999,N_15422);
nor UO_2096 (O_2096,N_16871,N_19986);
nor UO_2097 (O_2097,N_19694,N_18922);
or UO_2098 (O_2098,N_16188,N_18252);
or UO_2099 (O_2099,N_17201,N_18245);
nor UO_2100 (O_2100,N_15641,N_16799);
or UO_2101 (O_2101,N_15029,N_19290);
nand UO_2102 (O_2102,N_19083,N_18011);
nor UO_2103 (O_2103,N_18224,N_15206);
nand UO_2104 (O_2104,N_16489,N_18296);
or UO_2105 (O_2105,N_16494,N_18448);
nor UO_2106 (O_2106,N_16444,N_15054);
or UO_2107 (O_2107,N_19644,N_16411);
and UO_2108 (O_2108,N_18717,N_18137);
and UO_2109 (O_2109,N_16610,N_18258);
and UO_2110 (O_2110,N_16037,N_19781);
nor UO_2111 (O_2111,N_16380,N_18303);
or UO_2112 (O_2112,N_18688,N_19127);
or UO_2113 (O_2113,N_15413,N_16090);
or UO_2114 (O_2114,N_17513,N_15339);
nand UO_2115 (O_2115,N_17918,N_19023);
xnor UO_2116 (O_2116,N_18739,N_18696);
and UO_2117 (O_2117,N_15572,N_19191);
and UO_2118 (O_2118,N_16344,N_17510);
nor UO_2119 (O_2119,N_16442,N_15346);
or UO_2120 (O_2120,N_17627,N_16134);
or UO_2121 (O_2121,N_18964,N_17883);
nor UO_2122 (O_2122,N_19984,N_16173);
nor UO_2123 (O_2123,N_18903,N_16246);
and UO_2124 (O_2124,N_15383,N_17563);
and UO_2125 (O_2125,N_18950,N_18808);
and UO_2126 (O_2126,N_15687,N_18822);
or UO_2127 (O_2127,N_17870,N_19812);
or UO_2128 (O_2128,N_19579,N_15325);
and UO_2129 (O_2129,N_15816,N_16951);
nor UO_2130 (O_2130,N_18665,N_16833);
nor UO_2131 (O_2131,N_17196,N_17602);
nor UO_2132 (O_2132,N_16607,N_18081);
and UO_2133 (O_2133,N_15165,N_19989);
or UO_2134 (O_2134,N_15531,N_15623);
nor UO_2135 (O_2135,N_18171,N_17382);
nand UO_2136 (O_2136,N_16673,N_19856);
and UO_2137 (O_2137,N_17081,N_17767);
nand UO_2138 (O_2138,N_19441,N_16133);
nand UO_2139 (O_2139,N_18259,N_16927);
nand UO_2140 (O_2140,N_17809,N_16683);
nor UO_2141 (O_2141,N_15523,N_18087);
nand UO_2142 (O_2142,N_19717,N_18290);
nand UO_2143 (O_2143,N_15292,N_19487);
or UO_2144 (O_2144,N_19283,N_15525);
nor UO_2145 (O_2145,N_18198,N_15655);
and UO_2146 (O_2146,N_17758,N_18070);
or UO_2147 (O_2147,N_16293,N_19156);
and UO_2148 (O_2148,N_16773,N_17861);
or UO_2149 (O_2149,N_15429,N_18876);
nand UO_2150 (O_2150,N_19296,N_17528);
and UO_2151 (O_2151,N_17537,N_19024);
nor UO_2152 (O_2152,N_18281,N_19351);
nand UO_2153 (O_2153,N_15826,N_17741);
and UO_2154 (O_2154,N_15309,N_17546);
nor UO_2155 (O_2155,N_17650,N_16912);
or UO_2156 (O_2156,N_19063,N_19844);
nor UO_2157 (O_2157,N_19572,N_17094);
nand UO_2158 (O_2158,N_16873,N_17542);
or UO_2159 (O_2159,N_17387,N_15045);
nand UO_2160 (O_2160,N_18886,N_15407);
or UO_2161 (O_2161,N_18641,N_19172);
or UO_2162 (O_2162,N_15768,N_15179);
nor UO_2163 (O_2163,N_19329,N_17274);
nor UO_2164 (O_2164,N_18008,N_17671);
nand UO_2165 (O_2165,N_15497,N_19775);
or UO_2166 (O_2166,N_17846,N_17410);
and UO_2167 (O_2167,N_15902,N_17630);
or UO_2168 (O_2168,N_16580,N_17397);
or UO_2169 (O_2169,N_16078,N_19397);
nand UO_2170 (O_2170,N_19353,N_15169);
nand UO_2171 (O_2171,N_19420,N_16507);
nand UO_2172 (O_2172,N_18457,N_16174);
or UO_2173 (O_2173,N_18634,N_16300);
nor UO_2174 (O_2174,N_15410,N_19560);
nand UO_2175 (O_2175,N_17777,N_16441);
nand UO_2176 (O_2176,N_16023,N_17355);
nor UO_2177 (O_2177,N_19347,N_18917);
nor UO_2178 (O_2178,N_16990,N_15989);
and UO_2179 (O_2179,N_18118,N_18588);
and UO_2180 (O_2180,N_17391,N_15454);
nand UO_2181 (O_2181,N_19229,N_17166);
and UO_2182 (O_2182,N_15510,N_17156);
nand UO_2183 (O_2183,N_18878,N_19910);
and UO_2184 (O_2184,N_19649,N_17678);
and UO_2185 (O_2185,N_18328,N_15849);
xnor UO_2186 (O_2186,N_15916,N_19943);
or UO_2187 (O_2187,N_19088,N_16102);
nand UO_2188 (O_2188,N_19540,N_15219);
nor UO_2189 (O_2189,N_17052,N_19753);
or UO_2190 (O_2190,N_17884,N_17654);
or UO_2191 (O_2191,N_16178,N_16235);
or UO_2192 (O_2192,N_16285,N_16669);
or UO_2193 (O_2193,N_17063,N_17279);
nor UO_2194 (O_2194,N_19328,N_17736);
xnor UO_2195 (O_2195,N_15865,N_18169);
and UO_2196 (O_2196,N_18344,N_15568);
nand UO_2197 (O_2197,N_15785,N_17136);
nand UO_2198 (O_2198,N_18585,N_15657);
nor UO_2199 (O_2199,N_15018,N_18145);
nor UO_2200 (O_2200,N_16569,N_19573);
and UO_2201 (O_2201,N_17197,N_15658);
or UO_2202 (O_2202,N_15782,N_18546);
or UO_2203 (O_2203,N_15875,N_18813);
or UO_2204 (O_2204,N_18033,N_17859);
or UO_2205 (O_2205,N_18103,N_16894);
xor UO_2206 (O_2206,N_18927,N_17465);
nand UO_2207 (O_2207,N_15898,N_15596);
or UO_2208 (O_2208,N_16227,N_17805);
and UO_2209 (O_2209,N_16004,N_18007);
nand UO_2210 (O_2210,N_17863,N_17687);
nand UO_2211 (O_2211,N_15414,N_17164);
nor UO_2212 (O_2212,N_17110,N_17280);
xnor UO_2213 (O_2213,N_19723,N_17198);
nor UO_2214 (O_2214,N_17569,N_18148);
nor UO_2215 (O_2215,N_19674,N_15750);
nor UO_2216 (O_2216,N_16100,N_17779);
nand UO_2217 (O_2217,N_18028,N_16805);
nor UO_2218 (O_2218,N_18817,N_18078);
nand UO_2219 (O_2219,N_19493,N_17106);
or UO_2220 (O_2220,N_16852,N_17889);
nand UO_2221 (O_2221,N_15594,N_17342);
nor UO_2222 (O_2222,N_16644,N_16597);
nand UO_2223 (O_2223,N_16179,N_16658);
nand UO_2224 (O_2224,N_18415,N_18368);
nor UO_2225 (O_2225,N_19502,N_16202);
and UO_2226 (O_2226,N_15901,N_16248);
or UO_2227 (O_2227,N_15086,N_18638);
nor UO_2228 (O_2228,N_16748,N_19167);
nand UO_2229 (O_2229,N_16308,N_18740);
nand UO_2230 (O_2230,N_17007,N_16630);
xor UO_2231 (O_2231,N_18867,N_16983);
and UO_2232 (O_2232,N_19582,N_15532);
nor UO_2233 (O_2233,N_19913,N_19188);
xnor UO_2234 (O_2234,N_16839,N_18843);
and UO_2235 (O_2235,N_17027,N_18553);
nand UO_2236 (O_2236,N_18627,N_19727);
or UO_2237 (O_2237,N_18893,N_19049);
nand UO_2238 (O_2238,N_15171,N_18566);
nand UO_2239 (O_2239,N_17169,N_17834);
and UO_2240 (O_2240,N_17656,N_15137);
or UO_2241 (O_2241,N_17209,N_15979);
nand UO_2242 (O_2242,N_19937,N_18195);
nor UO_2243 (O_2243,N_15153,N_16863);
or UO_2244 (O_2244,N_19764,N_17842);
or UO_2245 (O_2245,N_17750,N_18486);
nand UO_2246 (O_2246,N_19359,N_17484);
or UO_2247 (O_2247,N_16192,N_18147);
nor UO_2248 (O_2248,N_18163,N_16641);
and UO_2249 (O_2249,N_17129,N_18478);
or UO_2250 (O_2250,N_19911,N_18127);
and UO_2251 (O_2251,N_18814,N_16296);
nand UO_2252 (O_2252,N_15911,N_19688);
nand UO_2253 (O_2253,N_16794,N_19112);
and UO_2254 (O_2254,N_18988,N_19249);
and UO_2255 (O_2255,N_19119,N_19925);
nand UO_2256 (O_2256,N_19437,N_17098);
xnor UO_2257 (O_2257,N_15761,N_17138);
nor UO_2258 (O_2258,N_19748,N_16612);
or UO_2259 (O_2259,N_18133,N_19795);
nand UO_2260 (O_2260,N_15261,N_16554);
and UO_2261 (O_2261,N_19551,N_19059);
nand UO_2262 (O_2262,N_17517,N_15465);
nand UO_2263 (O_2263,N_15935,N_18708);
nor UO_2264 (O_2264,N_18923,N_15273);
or UO_2265 (O_2265,N_16126,N_18757);
nand UO_2266 (O_2266,N_15078,N_15647);
nor UO_2267 (O_2267,N_19043,N_15980);
and UO_2268 (O_2268,N_18824,N_18470);
or UO_2269 (O_2269,N_17218,N_16533);
nand UO_2270 (O_2270,N_15064,N_18506);
nand UO_2271 (O_2271,N_19530,N_18175);
and UO_2272 (O_2272,N_19148,N_19323);
nor UO_2273 (O_2273,N_15536,N_19076);
nor UO_2274 (O_2274,N_18286,N_19415);
or UO_2275 (O_2275,N_15221,N_16232);
and UO_2276 (O_2276,N_18154,N_15812);
and UO_2277 (O_2277,N_18888,N_15258);
nor UO_2278 (O_2278,N_15778,N_18421);
and UO_2279 (O_2279,N_16846,N_18023);
nor UO_2280 (O_2280,N_16900,N_18931);
nand UO_2281 (O_2281,N_16487,N_15736);
and UO_2282 (O_2282,N_17356,N_15014);
nor UO_2283 (O_2283,N_15509,N_15542);
and UO_2284 (O_2284,N_17573,N_19905);
nand UO_2285 (O_2285,N_16279,N_18260);
nand UO_2286 (O_2286,N_16982,N_15021);
and UO_2287 (O_2287,N_16333,N_19670);
nor UO_2288 (O_2288,N_17909,N_17376);
and UO_2289 (O_2289,N_19288,N_18573);
or UO_2290 (O_2290,N_19074,N_18576);
nor UO_2291 (O_2291,N_17873,N_19581);
or UO_2292 (O_2292,N_17558,N_16692);
and UO_2293 (O_2293,N_18704,N_17568);
nor UO_2294 (O_2294,N_16321,N_19501);
and UO_2295 (O_2295,N_15673,N_18639);
and UO_2296 (O_2296,N_15009,N_18179);
nor UO_2297 (O_2297,N_19608,N_19655);
or UO_2298 (O_2298,N_15541,N_19771);
nor UO_2299 (O_2299,N_16567,N_18253);
nor UO_2300 (O_2300,N_15272,N_17167);
nor UO_2301 (O_2301,N_15934,N_19392);
and UO_2302 (O_2302,N_15960,N_19774);
nor UO_2303 (O_2303,N_17056,N_17642);
and UO_2304 (O_2304,N_19616,N_19814);
nand UO_2305 (O_2305,N_19997,N_17752);
and UO_2306 (O_2306,N_15835,N_18108);
or UO_2307 (O_2307,N_16288,N_18061);
nor UO_2308 (O_2308,N_15385,N_17535);
nand UO_2309 (O_2309,N_19936,N_18229);
or UO_2310 (O_2310,N_19101,N_19767);
and UO_2311 (O_2311,N_17155,N_18752);
nor UO_2312 (O_2312,N_17550,N_18322);
nand UO_2313 (O_2313,N_18683,N_18165);
nand UO_2314 (O_2314,N_17713,N_17583);
nand UO_2315 (O_2315,N_16556,N_19901);
and UO_2316 (O_2316,N_18455,N_16048);
and UO_2317 (O_2317,N_18610,N_16341);
nor UO_2318 (O_2318,N_16656,N_18304);
or UO_2319 (O_2319,N_15856,N_17797);
or UO_2320 (O_2320,N_15127,N_16939);
or UO_2321 (O_2321,N_15884,N_16860);
nand UO_2322 (O_2322,N_18375,N_18561);
or UO_2323 (O_2323,N_19568,N_15387);
and UO_2324 (O_2324,N_16654,N_16590);
nor UO_2325 (O_2325,N_18200,N_19633);
and UO_2326 (O_2326,N_15679,N_18207);
and UO_2327 (O_2327,N_19631,N_18472);
nand UO_2328 (O_2328,N_16822,N_19947);
nand UO_2329 (O_2329,N_16616,N_16212);
and UO_2330 (O_2330,N_19044,N_15208);
nand UO_2331 (O_2331,N_18381,N_15862);
or UO_2332 (O_2332,N_18678,N_19075);
nor UO_2333 (O_2333,N_18593,N_15607);
or UO_2334 (O_2334,N_17008,N_17211);
nor UO_2335 (O_2335,N_15845,N_15438);
nand UO_2336 (O_2336,N_17785,N_19238);
or UO_2337 (O_2337,N_19227,N_15182);
and UO_2338 (O_2338,N_17446,N_19004);
or UO_2339 (O_2339,N_19659,N_16486);
nand UO_2340 (O_2340,N_18622,N_15492);
xor UO_2341 (O_2341,N_15316,N_19868);
nand UO_2342 (O_2342,N_15197,N_19241);
and UO_2343 (O_2343,N_16710,N_17135);
and UO_2344 (O_2344,N_16495,N_16015);
or UO_2345 (O_2345,N_19979,N_16989);
nand UO_2346 (O_2346,N_18438,N_17124);
and UO_2347 (O_2347,N_19646,N_16104);
nand UO_2348 (O_2348,N_18630,N_18332);
or UO_2349 (O_2349,N_18459,N_17632);
and UO_2350 (O_2350,N_18756,N_15645);
nand UO_2351 (O_2351,N_17088,N_17972);
or UO_2352 (O_2352,N_19696,N_15574);
or UO_2353 (O_2353,N_18018,N_17773);
and UO_2354 (O_2354,N_17629,N_15005);
and UO_2355 (O_2355,N_16412,N_16454);
nand UO_2356 (O_2356,N_19636,N_17066);
nand UO_2357 (O_2357,N_19166,N_15858);
nor UO_2358 (O_2358,N_18429,N_19593);
nand UO_2359 (O_2359,N_15559,N_16194);
nand UO_2360 (O_2360,N_16332,N_15288);
nand UO_2361 (O_2361,N_17539,N_16615);
or UO_2362 (O_2362,N_16199,N_19538);
nand UO_2363 (O_2363,N_16362,N_19371);
nand UO_2364 (O_2364,N_15030,N_16131);
nor UO_2365 (O_2365,N_19576,N_17099);
nor UO_2366 (O_2366,N_15918,N_19494);
or UO_2367 (O_2367,N_17555,N_16483);
nand UO_2368 (O_2368,N_18916,N_18557);
nor UO_2369 (O_2369,N_19196,N_15270);
nor UO_2370 (O_2370,N_18277,N_17892);
or UO_2371 (O_2371,N_16952,N_18055);
nor UO_2372 (O_2372,N_15133,N_15746);
nor UO_2373 (O_2373,N_15202,N_18751);
nor UO_2374 (O_2374,N_19907,N_15099);
nand UO_2375 (O_2375,N_19754,N_15120);
or UO_2376 (O_2376,N_17684,N_15104);
and UO_2377 (O_2377,N_15614,N_15940);
and UO_2378 (O_2378,N_19899,N_17981);
nand UO_2379 (O_2379,N_19026,N_17565);
nand UO_2380 (O_2380,N_19266,N_16825);
or UO_2381 (O_2381,N_17574,N_19689);
nor UO_2382 (O_2382,N_18963,N_19432);
nand UO_2383 (O_2383,N_19992,N_18054);
and UO_2384 (O_2384,N_16566,N_17184);
and UO_2385 (O_2385,N_16592,N_15519);
xnor UO_2386 (O_2386,N_17879,N_18149);
nor UO_2387 (O_2387,N_16898,N_16239);
xnor UO_2388 (O_2388,N_18697,N_18887);
and UO_2389 (O_2389,N_18088,N_17507);
and UO_2390 (O_2390,N_16734,N_18374);
and UO_2391 (O_2391,N_18128,N_18477);
or UO_2392 (O_2392,N_17865,N_18269);
or UO_2393 (O_2393,N_19585,N_16735);
nand UO_2394 (O_2394,N_17126,N_16391);
xor UO_2395 (O_2395,N_19206,N_15668);
nor UO_2396 (O_2396,N_19740,N_15315);
and UO_2397 (O_2397,N_16121,N_17543);
nand UO_2398 (O_2398,N_15134,N_19541);
or UO_2399 (O_2399,N_15863,N_16434);
or UO_2400 (O_2400,N_15753,N_17692);
nor UO_2401 (O_2401,N_15723,N_19405);
or UO_2402 (O_2402,N_17991,N_17541);
and UO_2403 (O_2403,N_16872,N_18659);
nand UO_2404 (O_2404,N_19952,N_15129);
or UO_2405 (O_2405,N_17141,N_19846);
and UO_2406 (O_2406,N_19412,N_17792);
and UO_2407 (O_2407,N_17207,N_19918);
or UO_2408 (O_2408,N_19709,N_18907);
and UO_2409 (O_2409,N_17175,N_16272);
and UO_2410 (O_2410,N_16060,N_16639);
nand UO_2411 (O_2411,N_17470,N_16032);
and UO_2412 (O_2412,N_17998,N_17447);
and UO_2413 (O_2413,N_17529,N_17042);
and UO_2414 (O_2414,N_16716,N_17673);
nand UO_2415 (O_2415,N_17051,N_17934);
and UO_2416 (O_2416,N_17973,N_16791);
or UO_2417 (O_2417,N_17199,N_15840);
nand UO_2418 (O_2418,N_17472,N_16904);
and UO_2419 (O_2419,N_15023,N_15599);
or UO_2420 (O_2420,N_17090,N_19485);
nand UO_2421 (O_2421,N_17456,N_16998);
nor UO_2422 (O_2422,N_16314,N_16146);
nand UO_2423 (O_2423,N_16887,N_18821);
and UO_2424 (O_2424,N_18024,N_16106);
and UO_2425 (O_2425,N_17294,N_15421);
and UO_2426 (O_2426,N_19379,N_18578);
nand UO_2427 (O_2427,N_18490,N_19668);
nor UO_2428 (O_2428,N_18153,N_18419);
nor UO_2429 (O_2429,N_16270,N_17788);
or UO_2430 (O_2430,N_15073,N_18600);
and UO_2431 (O_2431,N_17975,N_18597);
or UO_2432 (O_2432,N_17116,N_15703);
xor UO_2433 (O_2433,N_18686,N_18172);
nor UO_2434 (O_2434,N_19592,N_18850);
nand UO_2435 (O_2435,N_19900,N_16073);
and UO_2436 (O_2436,N_16251,N_17285);
nand UO_2437 (O_2437,N_18554,N_19904);
or UO_2438 (O_2438,N_15786,N_18418);
nand UO_2439 (O_2439,N_16984,N_15538);
nand UO_2440 (O_2440,N_15908,N_16291);
or UO_2441 (O_2441,N_15824,N_19550);
nor UO_2442 (O_2442,N_17115,N_19454);
and UO_2443 (O_2443,N_16213,N_19559);
nor UO_2444 (O_2444,N_19267,N_15260);
and UO_2445 (O_2445,N_15961,N_15218);
nor UO_2446 (O_2446,N_15896,N_15152);
nor UO_2447 (O_2447,N_16875,N_17718);
nand UO_2448 (O_2448,N_16358,N_19417);
and UO_2449 (O_2449,N_15506,N_16958);
nor UO_2450 (O_2450,N_18865,N_15953);
and UO_2451 (O_2451,N_19529,N_18833);
nand UO_2452 (O_2452,N_19809,N_17050);
and UO_2453 (O_2453,N_15399,N_17518);
nand UO_2454 (O_2454,N_19117,N_15436);
nor UO_2455 (O_2455,N_18230,N_17828);
xor UO_2456 (O_2456,N_16094,N_16103);
nand UO_2457 (O_2457,N_17130,N_15360);
or UO_2458 (O_2458,N_16231,N_19704);
nor UO_2459 (O_2459,N_17146,N_15818);
nor UO_2460 (O_2460,N_17962,N_16932);
nand UO_2461 (O_2461,N_15832,N_19799);
and UO_2462 (O_2462,N_19222,N_18872);
or UO_2463 (O_2463,N_15327,N_18805);
or UO_2464 (O_2464,N_16466,N_17400);
and UO_2465 (O_2465,N_16475,N_18458);
nor UO_2466 (O_2466,N_15950,N_16383);
xor UO_2467 (O_2467,N_18408,N_15737);
nor UO_2468 (O_2468,N_16897,N_19450);
nand UO_2469 (O_2469,N_15194,N_17344);
and UO_2470 (O_2470,N_19691,N_15081);
or UO_2471 (O_2471,N_17149,N_16276);
and UO_2472 (O_2472,N_17598,N_17944);
nor UO_2473 (O_2473,N_19888,N_18692);
xnor UO_2474 (O_2474,N_19669,N_18305);
nor UO_2475 (O_2475,N_17577,N_16840);
and UO_2476 (O_2476,N_17429,N_19442);
nor UO_2477 (O_2477,N_19884,N_17634);
and UO_2478 (O_2478,N_17799,N_16801);
nand UO_2479 (O_2479,N_17806,N_16171);
nand UO_2480 (O_2480,N_17698,N_18026);
and UO_2481 (O_2481,N_16725,N_16935);
nand UO_2482 (O_2482,N_16127,N_19587);
nor UO_2483 (O_2483,N_18240,N_19595);
and UO_2484 (O_2484,N_15048,N_15132);
or UO_2485 (O_2485,N_19202,N_17144);
nand UO_2486 (O_2486,N_19980,N_15406);
nand UO_2487 (O_2487,N_15722,N_18874);
or UO_2488 (O_2488,N_16972,N_18524);
xnor UO_2489 (O_2489,N_15621,N_17878);
nor UO_2490 (O_2490,N_18901,N_19410);
and UO_2491 (O_2491,N_18099,N_19639);
nand UO_2492 (O_2492,N_17309,N_15476);
and UO_2493 (O_2493,N_16936,N_15779);
and UO_2494 (O_2494,N_18235,N_19345);
xnor UO_2495 (O_2495,N_17255,N_16699);
or UO_2496 (O_2496,N_19462,N_16035);
nor UO_2497 (O_2497,N_17424,N_16700);
or UO_2498 (O_2498,N_17930,N_18608);
or UO_2499 (O_2499,N_19066,N_15160);
endmodule