module basic_1500_15000_2000_15_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_178,In_233);
or U1 (N_1,In_848,In_492);
and U2 (N_2,In_725,In_459);
or U3 (N_3,In_743,In_778);
nor U4 (N_4,In_1348,In_977);
xnor U5 (N_5,In_1241,In_1382);
or U6 (N_6,In_1069,In_936);
and U7 (N_7,In_791,In_1456);
nand U8 (N_8,In_984,In_1391);
and U9 (N_9,In_240,In_904);
nand U10 (N_10,In_625,In_786);
nand U11 (N_11,In_793,In_1002);
nand U12 (N_12,In_466,In_79);
and U13 (N_13,In_1200,In_324);
or U14 (N_14,In_511,In_728);
nor U15 (N_15,In_276,In_767);
nor U16 (N_16,In_171,In_1025);
and U17 (N_17,In_1027,In_880);
and U18 (N_18,In_92,In_1203);
nand U19 (N_19,In_1379,In_199);
and U20 (N_20,In_1048,In_953);
and U21 (N_21,In_735,In_773);
or U22 (N_22,In_495,In_869);
or U23 (N_23,In_1091,In_678);
xnor U24 (N_24,In_437,In_690);
nand U25 (N_25,In_980,In_1285);
xor U26 (N_26,In_390,In_343);
xor U27 (N_27,In_284,In_1433);
xor U28 (N_28,In_841,In_1442);
nand U29 (N_29,In_1330,In_760);
xnor U30 (N_30,In_71,In_1491);
or U31 (N_31,In_361,In_1314);
nand U32 (N_32,In_95,In_1394);
xnor U33 (N_33,In_372,In_1232);
nor U34 (N_34,In_729,In_562);
and U35 (N_35,In_1411,In_1070);
nor U36 (N_36,In_1323,In_1169);
nor U37 (N_37,In_380,In_400);
or U38 (N_38,In_1135,In_1039);
or U39 (N_39,In_1041,In_603);
or U40 (N_40,In_70,In_109);
or U41 (N_41,In_15,In_216);
xnor U42 (N_42,In_815,In_471);
or U43 (N_43,In_98,In_682);
or U44 (N_44,In_1472,In_812);
or U45 (N_45,In_427,In_1176);
nand U46 (N_46,In_863,In_589);
nor U47 (N_47,In_247,In_269);
nor U48 (N_48,In_438,In_648);
or U49 (N_49,In_1020,In_1036);
xnor U50 (N_50,In_765,In_1454);
and U51 (N_51,In_691,In_948);
or U52 (N_52,In_127,In_218);
nand U53 (N_53,In_1123,In_1354);
or U54 (N_54,In_1292,In_148);
and U55 (N_55,In_619,In_1356);
or U56 (N_56,In_330,In_851);
nand U57 (N_57,In_584,In_111);
nand U58 (N_58,In_701,In_248);
nand U59 (N_59,In_813,In_1358);
xor U60 (N_60,In_420,In_886);
and U61 (N_61,In_1440,In_277);
nand U62 (N_62,In_933,In_1298);
nand U63 (N_63,In_794,In_1265);
or U64 (N_64,In_925,In_810);
nor U65 (N_65,In_181,In_1045);
nand U66 (N_66,In_480,In_961);
nor U67 (N_67,In_1450,In_297);
nand U68 (N_68,In_775,In_852);
or U69 (N_69,In_1403,In_833);
nand U70 (N_70,In_858,In_431);
xnor U71 (N_71,In_369,In_300);
and U72 (N_72,In_1238,In_103);
and U73 (N_73,In_2,In_644);
or U74 (N_74,In_456,In_789);
and U75 (N_75,In_1395,In_1386);
xor U76 (N_76,In_999,In_604);
nand U77 (N_77,In_751,In_164);
or U78 (N_78,In_874,In_558);
nor U79 (N_79,In_496,In_22);
nor U80 (N_80,In_721,In_637);
nand U81 (N_81,In_843,In_43);
nor U82 (N_82,In_1088,In_110);
and U83 (N_83,In_94,In_479);
nor U84 (N_84,In_387,In_1233);
or U85 (N_85,In_453,In_32);
nand U86 (N_86,In_531,In_707);
nor U87 (N_87,In_692,In_1335);
or U88 (N_88,In_757,In_261);
nor U89 (N_89,In_772,In_1311);
nand U90 (N_90,In_266,In_972);
and U91 (N_91,In_344,In_83);
and U92 (N_92,In_184,In_1026);
nor U93 (N_93,In_238,In_1243);
nand U94 (N_94,In_1283,In_1365);
xnor U95 (N_95,In_870,In_124);
nand U96 (N_96,In_1464,In_1195);
or U97 (N_97,In_1306,In_561);
xnor U98 (N_98,In_846,In_1353);
nand U99 (N_99,In_954,In_887);
xor U100 (N_100,In_1484,In_195);
or U101 (N_101,In_1370,In_879);
nand U102 (N_102,In_150,In_1420);
xor U103 (N_103,In_1287,In_1159);
nand U104 (N_104,In_667,In_436);
nor U105 (N_105,In_1217,In_900);
xor U106 (N_106,In_602,In_175);
and U107 (N_107,In_1104,In_123);
nand U108 (N_108,In_1368,In_366);
nor U109 (N_109,In_1384,In_1174);
and U110 (N_110,In_236,In_967);
nand U111 (N_111,In_287,In_264);
xnor U112 (N_112,In_401,In_742);
and U113 (N_113,In_1250,In_307);
xor U114 (N_114,In_1166,In_393);
or U115 (N_115,In_86,In_906);
and U116 (N_116,In_173,In_635);
and U117 (N_117,In_926,In_52);
nor U118 (N_118,In_1385,In_1448);
nor U119 (N_119,In_1219,In_1300);
and U120 (N_120,In_740,In_1101);
nor U121 (N_121,In_590,In_1278);
nor U122 (N_122,In_1255,In_413);
and U123 (N_123,In_458,In_213);
and U124 (N_124,In_769,In_566);
xnor U125 (N_125,In_1383,In_352);
nor U126 (N_126,In_280,In_271);
nand U127 (N_127,In_816,In_1156);
nand U128 (N_128,In_1415,In_1162);
nand U129 (N_129,In_314,In_824);
and U130 (N_130,In_1266,In_1142);
xnor U131 (N_131,In_1149,In_345);
and U132 (N_132,In_1270,In_1342);
or U133 (N_133,In_1252,In_623);
nand U134 (N_134,In_265,In_770);
nor U135 (N_135,In_342,In_859);
nor U136 (N_136,In_430,In_446);
or U137 (N_137,In_1230,In_1102);
nor U138 (N_138,In_48,In_696);
and U139 (N_139,In_541,In_463);
nand U140 (N_140,In_785,In_677);
nor U141 (N_141,In_597,In_397);
nand U142 (N_142,In_1380,In_726);
nand U143 (N_143,In_534,In_285);
nor U144 (N_144,In_1161,In_1204);
xnor U145 (N_145,In_717,In_1444);
or U146 (N_146,In_1181,In_334);
nor U147 (N_147,In_358,In_731);
nand U148 (N_148,In_513,In_1167);
nand U149 (N_149,In_99,In_371);
or U150 (N_150,In_179,In_1184);
nand U151 (N_151,In_473,In_1077);
or U152 (N_152,In_1202,In_647);
or U153 (N_153,In_31,In_655);
xor U154 (N_154,In_565,In_790);
and U155 (N_155,In_1488,In_620);
or U156 (N_156,In_1117,In_553);
nor U157 (N_157,In_1254,In_36);
nand U158 (N_158,In_613,In_1486);
nor U159 (N_159,In_362,In_423);
nand U160 (N_160,In_1482,In_806);
or U161 (N_161,In_1136,In_152);
and U162 (N_162,In_34,In_581);
and U163 (N_163,In_258,In_1453);
or U164 (N_164,In_820,In_1303);
xnor U165 (N_165,In_1115,In_381);
nand U166 (N_166,In_481,In_802);
and U167 (N_167,In_807,In_549);
nand U168 (N_168,In_777,In_836);
and U169 (N_169,In_1201,In_235);
nand U170 (N_170,In_272,In_1302);
nand U171 (N_171,In_808,In_39);
nor U172 (N_172,In_1079,In_1044);
nor U173 (N_173,In_1223,In_1248);
nand U174 (N_174,In_659,In_850);
nand U175 (N_175,In_20,In_364);
nand U176 (N_176,In_503,In_162);
nor U177 (N_177,In_1017,In_85);
or U178 (N_178,In_931,In_1053);
nand U179 (N_179,In_141,In_571);
xnor U180 (N_180,In_1022,In_1057);
or U181 (N_181,In_640,In_694);
or U182 (N_182,In_712,In_395);
nor U183 (N_183,In_305,In_291);
nor U184 (N_184,In_651,In_24);
nand U185 (N_185,In_222,In_895);
nor U186 (N_186,In_1094,In_1180);
xor U187 (N_187,In_1112,In_1496);
and U188 (N_188,In_744,In_1362);
nor U189 (N_189,In_1492,In_1421);
or U190 (N_190,In_142,In_1494);
xnor U191 (N_191,In_551,In_1452);
or U192 (N_192,In_1163,In_243);
or U193 (N_193,In_595,In_924);
nand U194 (N_194,In_392,In_897);
and U195 (N_195,In_74,In_660);
and U196 (N_196,In_55,In_733);
or U197 (N_197,In_512,In_185);
xnor U198 (N_198,In_875,In_662);
nor U199 (N_199,In_1092,In_599);
and U200 (N_200,In_125,In_434);
and U201 (N_201,In_295,In_348);
nand U202 (N_202,In_814,In_1175);
xnor U203 (N_203,In_1465,In_835);
xnor U204 (N_204,In_1046,In_1436);
nor U205 (N_205,In_629,In_1468);
and U206 (N_206,In_988,In_1324);
nor U207 (N_207,In_630,In_1304);
nor U208 (N_208,In_282,In_255);
or U209 (N_209,In_1445,In_1376);
xor U210 (N_210,In_335,In_405);
or U211 (N_211,In_828,In_302);
and U212 (N_212,In_776,In_166);
nand U213 (N_213,In_831,In_1032);
or U214 (N_214,In_1308,In_902);
nand U215 (N_215,In_256,In_1439);
nand U216 (N_216,In_464,In_1349);
and U217 (N_217,In_593,In_1253);
nand U218 (N_218,In_616,In_940);
nor U219 (N_219,In_766,In_1);
xnor U220 (N_220,In_1000,In_44);
nand U221 (N_221,In_1011,In_102);
or U222 (N_222,In_560,In_665);
nand U223 (N_223,In_1033,In_636);
or U224 (N_224,In_354,In_645);
or U225 (N_225,In_1222,In_1327);
xor U226 (N_226,In_29,In_546);
nor U227 (N_227,In_1108,In_847);
or U228 (N_228,In_1145,In_1013);
or U229 (N_229,In_1319,In_1393);
xnor U230 (N_230,In_1090,In_1364);
nor U231 (N_231,In_1082,In_505);
nor U232 (N_232,In_129,In_618);
nor U233 (N_233,In_469,In_674);
and U234 (N_234,In_861,In_1279);
nand U235 (N_235,In_842,In_37);
xnor U236 (N_236,In_117,In_928);
nand U237 (N_237,In_1332,In_1305);
or U238 (N_238,In_1430,In_965);
nor U239 (N_239,In_122,In_270);
and U240 (N_240,In_732,In_3);
or U241 (N_241,In_1224,In_33);
nand U242 (N_242,In_433,In_622);
nor U243 (N_243,In_356,In_1211);
xnor U244 (N_244,In_1274,In_13);
or U245 (N_245,In_871,In_1478);
nor U246 (N_246,In_12,In_1009);
nand U247 (N_247,In_476,In_782);
nand U248 (N_248,In_1346,In_1414);
or U249 (N_249,In_1471,In_781);
nand U250 (N_250,In_347,In_527);
or U251 (N_251,In_730,In_706);
nand U252 (N_252,In_498,In_245);
and U253 (N_253,In_1441,In_153);
and U254 (N_254,In_488,In_779);
or U255 (N_255,In_719,In_329);
or U256 (N_256,In_508,In_909);
nor U257 (N_257,In_196,In_693);
or U258 (N_258,In_950,In_143);
nor U259 (N_259,In_507,In_1231);
nand U260 (N_260,In_1047,In_722);
nand U261 (N_261,In_359,In_56);
and U262 (N_262,In_614,In_19);
nor U263 (N_263,In_891,In_1185);
nor U264 (N_264,In_1271,In_1343);
nand U265 (N_265,In_955,In_225);
nor U266 (N_266,In_144,In_1240);
or U267 (N_267,In_943,In_580);
nand U268 (N_268,In_45,In_17);
nor U269 (N_269,In_1320,In_1133);
or U270 (N_270,In_226,In_987);
nand U271 (N_271,In_1351,In_72);
nor U272 (N_272,In_537,In_296);
or U273 (N_273,In_1297,In_1316);
and U274 (N_274,In_714,In_191);
and U275 (N_275,In_1205,In_1338);
nand U276 (N_276,In_823,In_215);
nor U277 (N_277,In_100,In_42);
nand U278 (N_278,In_242,In_1155);
and U279 (N_279,In_1100,In_1144);
and U280 (N_280,In_1097,In_1409);
nand U281 (N_281,In_478,In_440);
or U282 (N_282,In_819,In_576);
nand U283 (N_283,In_327,In_1268);
or U284 (N_284,In_681,In_115);
or U285 (N_285,In_1473,In_1193);
nor U286 (N_286,In_1416,In_1059);
nor U287 (N_287,In_1321,In_567);
nand U288 (N_288,In_1431,In_254);
and U289 (N_289,In_176,In_1010);
or U290 (N_290,In_130,In_403);
or U291 (N_291,In_239,In_539);
nand U292 (N_292,In_1493,In_1328);
nand U293 (N_293,In_448,In_339);
nand U294 (N_294,In_518,In_994);
nand U295 (N_295,In_862,In_1212);
nand U296 (N_296,In_1260,In_809);
or U297 (N_297,In_151,In_997);
nand U298 (N_298,In_522,In_985);
nor U299 (N_299,In_155,In_992);
nor U300 (N_300,In_1138,In_1438);
or U301 (N_301,In_121,In_154);
nor U302 (N_302,In_587,In_1178);
or U303 (N_303,In_723,In_177);
and U304 (N_304,In_1085,In_490);
and U305 (N_305,In_556,In_1256);
nand U306 (N_306,In_550,In_385);
and U307 (N_307,In_652,In_1463);
or U308 (N_308,In_419,In_375);
and U309 (N_309,In_1375,In_586);
and U310 (N_310,In_796,In_856);
nor U311 (N_311,In_1281,In_941);
nand U312 (N_312,In_1006,In_220);
nand U313 (N_313,In_727,In_1004);
nor U314 (N_314,In_156,In_684);
nor U315 (N_315,In_552,In_351);
and U316 (N_316,In_801,In_461);
or U317 (N_317,In_749,In_1063);
and U318 (N_318,In_1434,In_396);
nor U319 (N_319,In_529,In_1018);
xnor U320 (N_320,In_410,In_452);
or U321 (N_321,In_570,In_10);
or U322 (N_322,In_963,In_612);
nor U323 (N_323,In_829,In_1127);
and U324 (N_324,In_1336,In_1483);
and U325 (N_325,In_698,In_736);
nand U326 (N_326,In_1043,In_1150);
or U327 (N_327,In_908,In_1152);
xor U328 (N_328,In_485,In_1151);
nand U329 (N_329,In_0,In_415);
nor U330 (N_330,In_800,In_292);
or U331 (N_331,In_1098,In_1289);
or U332 (N_332,In_1273,In_989);
or U333 (N_333,In_1113,In_864);
or U334 (N_334,In_439,In_9);
nor U335 (N_335,In_946,In_425);
nand U336 (N_336,In_533,In_517);
and U337 (N_337,In_670,In_4);
and U338 (N_338,In_1401,In_1008);
nand U339 (N_339,In_1242,In_116);
or U340 (N_340,In_1019,In_326);
nand U341 (N_341,In_873,In_536);
nor U342 (N_342,In_407,In_911);
or U343 (N_343,In_1470,In_982);
xor U344 (N_344,In_418,In_1106);
and U345 (N_345,In_697,In_249);
or U346 (N_346,In_288,In_394);
or U347 (N_347,In_145,In_956);
or U348 (N_348,In_1446,In_26);
nor U349 (N_349,In_46,In_598);
or U350 (N_350,In_878,In_1239);
or U351 (N_351,In_50,In_1272);
and U352 (N_352,In_1132,In_82);
nand U353 (N_353,In_204,In_376);
or U354 (N_354,In_606,In_1124);
nand U355 (N_355,In_1139,In_1055);
or U356 (N_356,In_1475,In_1194);
and U357 (N_357,In_1425,In_308);
nand U358 (N_358,In_1387,In_208);
or U359 (N_359,In_84,In_542);
nand U360 (N_360,In_1315,In_140);
and U361 (N_361,In_474,In_1359);
nand U362 (N_362,In_675,In_61);
xnor U363 (N_363,In_1012,In_1143);
nand U364 (N_364,In_1207,In_1076);
nor U365 (N_365,In_1390,In_379);
nand U366 (N_366,In_1128,In_161);
or U367 (N_367,In_658,In_221);
nand U368 (N_368,In_686,In_1107);
and U369 (N_369,In_237,In_408);
nand U370 (N_370,In_641,In_1220);
or U371 (N_371,In_914,In_460);
or U372 (N_372,In_457,In_1227);
or U373 (N_373,In_1427,In_332);
nor U374 (N_374,In_455,In_710);
and U375 (N_375,In_654,In_554);
and U376 (N_376,In_1126,In_1003);
nor U377 (N_377,In_594,In_1408);
nand U378 (N_378,In_197,In_1392);
and U379 (N_379,In_388,In_1075);
or U380 (N_380,In_234,In_1058);
nand U381 (N_381,In_839,In_788);
nor U382 (N_382,In_1301,In_336);
nand U383 (N_383,In_319,In_1487);
nor U384 (N_384,In_840,In_857);
or U385 (N_385,In_1423,In_47);
nand U386 (N_386,In_1485,In_1345);
nor U387 (N_387,In_268,In_1410);
nand U388 (N_388,In_210,In_798);
and U389 (N_389,In_1405,In_1312);
or U390 (N_390,In_1131,In_49);
nor U391 (N_391,In_206,In_320);
nand U392 (N_392,In_502,In_827);
and U393 (N_393,In_1280,In_532);
nor U394 (N_394,In_544,In_1049);
nand U395 (N_395,In_783,In_306);
xnor U396 (N_396,In_165,In_1397);
or U397 (N_397,In_1286,In_572);
or U398 (N_398,In_958,In_484);
nand U399 (N_399,In_991,In_849);
nor U400 (N_400,In_350,In_412);
or U401 (N_401,In_1209,In_1062);
nor U402 (N_402,In_718,In_1313);
and U403 (N_403,In_1457,In_715);
or U404 (N_404,In_298,In_611);
nor U405 (N_405,In_695,In_90);
and U406 (N_406,In_1284,In_169);
nand U407 (N_407,In_929,In_201);
or U408 (N_408,In_1072,In_108);
or U409 (N_409,In_617,In_979);
or U410 (N_410,In_974,In_938);
or U411 (N_411,In_526,In_106);
nand U412 (N_412,In_462,In_608);
and U413 (N_413,In_569,In_609);
or U414 (N_414,In_1089,In_889);
or U415 (N_415,In_1015,In_657);
or U416 (N_416,In_57,In_628);
and U417 (N_417,In_1038,In_600);
and U418 (N_418,In_1105,In_1388);
nand U419 (N_419,In_523,In_355);
nand U420 (N_420,In_942,In_1299);
and U421 (N_421,In_883,In_756);
nor U422 (N_422,In_1495,In_406);
and U423 (N_423,In_1035,In_912);
or U424 (N_424,In_750,In_1235);
nor U425 (N_425,In_1141,In_192);
and U426 (N_426,In_668,In_855);
or U427 (N_427,In_653,In_450);
nand U428 (N_428,In_1218,In_318);
or U429 (N_429,In_1074,In_905);
or U430 (N_430,In_1014,In_409);
nand U431 (N_431,In_250,In_817);
or U432 (N_432,In_278,In_69);
nand U433 (N_433,In_771,In_952);
or U434 (N_434,In_601,In_370);
and U435 (N_435,In_1129,In_1054);
nor U436 (N_436,In_1310,In_1190);
or U437 (N_437,In_795,In_205);
nor U438 (N_438,In_1398,In_441);
or U439 (N_439,In_892,In_559);
and U440 (N_440,In_834,In_762);
or U441 (N_441,In_40,In_983);
or U442 (N_442,In_411,In_525);
nor U443 (N_443,In_1083,In_624);
nand U444 (N_444,In_1052,In_232);
or U445 (N_445,In_182,In_1462);
and U446 (N_446,In_1093,In_6);
and U447 (N_447,In_1114,In_1296);
xnor U448 (N_448,In_377,In_759);
nand U449 (N_449,In_7,In_1418);
nand U450 (N_450,In_649,In_968);
xor U451 (N_451,In_244,In_428);
or U452 (N_452,In_1479,In_1366);
and U453 (N_453,In_451,In_337);
nand U454 (N_454,In_632,In_313);
and U455 (N_455,In_489,In_1412);
nor U456 (N_456,In_1435,In_995);
nand U457 (N_457,In_1341,In_564);
and U458 (N_458,In_1029,In_1179);
nor U459 (N_459,In_317,In_1307);
and U460 (N_460,In_228,In_530);
xor U461 (N_461,In_607,In_180);
or U462 (N_462,In_1067,In_1363);
nand U463 (N_463,In_753,In_1459);
or U464 (N_464,In_91,In_916);
and U465 (N_465,In_310,In_704);
and U466 (N_466,In_646,In_229);
nand U467 (N_467,In_399,In_1153);
and U468 (N_468,In_1005,In_1206);
and U469 (N_469,In_1171,In_214);
and U470 (N_470,In_207,In_818);
and U471 (N_471,In_1337,In_93);
and U472 (N_472,In_890,In_1078);
and U473 (N_473,In_68,In_1121);
nand U474 (N_474,In_444,In_573);
or U475 (N_475,In_1417,In_1118);
xor U476 (N_476,In_1317,In_309);
and U477 (N_477,In_1367,In_1196);
or U478 (N_478,In_132,In_1476);
and U479 (N_479,In_315,In_21);
nor U480 (N_480,In_519,In_365);
nor U481 (N_481,In_1361,In_1269);
and U482 (N_482,In_475,In_780);
nor U483 (N_483,In_231,In_1490);
and U484 (N_484,In_1389,In_510);
and U485 (N_485,In_993,In_884);
nand U486 (N_486,In_1165,In_976);
and U487 (N_487,In_200,In_1023);
nor U488 (N_488,In_1068,In_135);
or U489 (N_489,In_325,In_579);
and U490 (N_490,In_1229,In_1396);
nor U491 (N_491,In_80,In_520);
nand U492 (N_492,In_1371,In_1400);
or U493 (N_493,In_923,In_1237);
or U494 (N_494,In_51,In_913);
nor U495 (N_495,In_1455,In_1001);
nor U496 (N_496,In_230,In_1251);
or U497 (N_497,In_1419,In_755);
or U498 (N_498,In_190,In_761);
and U499 (N_499,In_1110,In_1111);
and U500 (N_500,In_1489,In_872);
and U501 (N_501,In_784,In_866);
nor U502 (N_502,In_787,In_515);
and U503 (N_503,In_937,In_557);
nand U504 (N_504,In_643,In_1191);
nand U505 (N_505,In_768,In_81);
xnor U506 (N_506,In_257,In_73);
and U507 (N_507,In_838,In_799);
and U508 (N_508,In_758,In_907);
and U509 (N_509,In_1099,In_1183);
or U510 (N_510,In_134,In_1333);
nor U511 (N_511,In_126,In_501);
nor U512 (N_512,In_107,In_391);
or U513 (N_513,In_592,In_1428);
and U514 (N_514,In_1173,In_754);
nand U515 (N_515,In_830,In_960);
or U516 (N_516,In_1172,In_605);
or U517 (N_517,In_118,In_1116);
or U518 (N_518,In_170,In_312);
or U519 (N_519,In_1061,In_241);
nor U520 (N_520,In_971,In_1016);
and U521 (N_521,In_521,In_1051);
nand U522 (N_522,In_1261,In_639);
nor U523 (N_523,In_650,In_899);
and U524 (N_524,In_1234,In_574);
nor U525 (N_525,In_188,In_1007);
nand U526 (N_526,In_998,In_1037);
nor U527 (N_527,In_89,In_194);
nand U528 (N_528,In_1066,In_360);
nand U529 (N_529,In_1399,In_138);
and U530 (N_530,In_1182,In_88);
or U531 (N_531,In_187,In_713);
nand U532 (N_532,In_30,In_1168);
nand U533 (N_533,In_1215,In_23);
or U534 (N_534,In_930,In_62);
nor U535 (N_535,In_59,In_54);
and U536 (N_536,In_1056,In_417);
xor U537 (N_537,In_1334,In_1498);
nor U538 (N_538,In_981,In_443);
nor U539 (N_539,In_699,In_1481);
nor U540 (N_540,In_724,In_867);
or U541 (N_541,In_1373,In_664);
nor U542 (N_542,In_934,In_1458);
xnor U543 (N_543,In_87,In_575);
or U544 (N_544,In_267,In_432);
nand U545 (N_545,In_1221,In_1322);
and U546 (N_546,In_1146,In_1164);
and U547 (N_547,In_555,In_16);
and U548 (N_548,In_738,In_1426);
and U549 (N_549,In_363,In_331);
nor U550 (N_550,In_881,In_734);
or U551 (N_551,In_104,In_414);
or U552 (N_552,In_346,In_514);
nor U553 (N_553,In_1461,In_445);
and U554 (N_554,In_633,In_825);
xor U555 (N_555,In_545,In_1350);
and U556 (N_556,In_1451,In_882);
or U557 (N_557,In_969,In_638);
and U558 (N_558,In_301,In_66);
nand U559 (N_559,In_128,In_1360);
and U560 (N_560,In_634,In_426);
xnor U561 (N_561,In_1357,In_877);
nand U562 (N_562,In_223,In_1267);
nand U563 (N_563,In_1187,In_1377);
or U564 (N_564,In_1344,In_1247);
nand U565 (N_565,In_671,In_826);
and U566 (N_566,In_563,In_1262);
or U567 (N_567,In_1443,In_1480);
or U568 (N_568,In_1404,In_1065);
xor U569 (N_569,In_367,In_688);
nand U570 (N_570,In_389,In_131);
and U571 (N_571,In_1294,In_1024);
and U572 (N_572,In_1244,In_1402);
nor U573 (N_573,In_745,In_922);
or U574 (N_574,In_535,In_304);
nor U575 (N_575,In_716,In_1080);
and U576 (N_576,In_1050,In_666);
xor U577 (N_577,In_1060,In_1154);
and U578 (N_578,In_853,In_959);
and U579 (N_579,In_449,In_1340);
or U580 (N_580,In_8,In_113);
xnor U581 (N_581,In_661,In_1326);
xor U582 (N_582,In_1103,In_917);
nand U583 (N_583,In_1210,In_333);
nand U584 (N_584,In_168,In_374);
and U585 (N_585,In_316,In_477);
or U586 (N_586,In_38,In_158);
or U587 (N_587,In_516,In_1449);
nand U588 (N_588,In_626,In_1125);
nor U589 (N_589,In_1245,In_506);
nor U590 (N_590,In_1147,In_894);
nor U591 (N_591,In_491,In_212);
or U592 (N_592,In_119,In_378);
and U593 (N_593,In_146,In_1120);
nor U594 (N_594,In_700,In_1130);
or U595 (N_595,In_281,In_1466);
nand U596 (N_596,In_1021,In_741);
and U597 (N_597,In_447,In_203);
or U598 (N_598,In_468,In_353);
xnor U599 (N_599,In_1214,In_1407);
and U600 (N_600,In_77,In_1263);
nand U601 (N_601,In_582,In_357);
or U602 (N_602,In_687,In_1122);
or U603 (N_603,In_837,In_328);
and U604 (N_604,In_865,In_709);
xor U605 (N_605,In_1339,In_1369);
nand U606 (N_606,In_1071,In_860);
or U607 (N_607,In_1216,In_1087);
nor U608 (N_608,In_1040,In_918);
and U609 (N_609,In_465,In_896);
xnor U610 (N_610,In_67,In_435);
and U611 (N_611,In_680,In_1309);
and U612 (N_612,In_975,In_472);
xor U613 (N_613,In_548,In_822);
or U614 (N_614,In_1095,In_547);
or U615 (N_615,In_1086,In_373);
or U616 (N_616,In_186,In_1264);
or U617 (N_617,In_1028,In_27);
nand U618 (N_618,In_673,In_504);
and U619 (N_619,In_227,In_947);
nand U620 (N_620,In_1460,In_167);
and U621 (N_621,In_75,In_583);
nand U622 (N_622,In_509,In_424);
and U623 (N_623,In_1225,In_159);
xnor U624 (N_624,In_1236,In_290);
and U625 (N_625,In_493,In_76);
nand U626 (N_626,In_803,In_252);
or U627 (N_627,In_18,In_1374);
nand U628 (N_628,In_921,In_898);
nand U629 (N_629,In_211,In_703);
nor U630 (N_630,In_136,In_683);
nor U631 (N_631,In_811,In_990);
nor U632 (N_632,In_1497,In_1197);
or U633 (N_633,In_1276,In_97);
nor U634 (N_634,In_1355,In_1474);
nor U635 (N_635,In_1325,In_966);
nand U636 (N_636,In_217,In_1198);
and U637 (N_637,In_627,In_1290);
nand U638 (N_638,In_944,In_578);
nand U639 (N_639,In_1199,In_1378);
or U640 (N_640,In_568,In_538);
nor U641 (N_641,In_274,In_1189);
nand U642 (N_642,In_845,In_663);
xor U643 (N_643,In_64,In_676);
nand U644 (N_644,In_286,In_747);
or U645 (N_645,In_65,In_540);
and U646 (N_646,In_1148,In_935);
and U647 (N_647,In_183,In_147);
nor U648 (N_648,In_1432,In_705);
nand U649 (N_649,In_1246,In_708);
nand U650 (N_650,In_1137,In_1257);
and U651 (N_651,In_299,In_486);
nor U652 (N_652,In_1208,In_137);
nor U653 (N_653,In_96,In_383);
and U654 (N_654,In_340,In_341);
xor U655 (N_655,In_1140,In_764);
and U656 (N_656,In_1499,In_1081);
nand U657 (N_657,In_35,In_202);
and U658 (N_658,In_1158,In_382);
nand U659 (N_659,In_467,In_1293);
nor U660 (N_660,In_172,In_832);
nor U661 (N_661,In_279,In_1259);
nand U662 (N_662,In_669,In_792);
xnor U663 (N_663,In_1258,In_888);
nand U664 (N_664,In_1192,In_679);
or U665 (N_665,In_1170,In_251);
or U666 (N_666,In_1073,In_262);
nor U667 (N_667,In_774,In_1186);
or U668 (N_668,In_454,In_112);
or U669 (N_669,In_901,In_1295);
nor U670 (N_670,In_1477,In_1291);
or U671 (N_671,In_876,In_283);
nor U672 (N_672,In_1437,In_752);
nor U673 (N_673,In_1157,In_157);
nor U674 (N_674,In_631,In_964);
nand U675 (N_675,In_949,In_483);
nand U676 (N_676,In_5,In_416);
or U677 (N_677,In_368,In_672);
or U678 (N_678,In_1413,In_1277);
nand U679 (N_679,In_421,In_101);
and U680 (N_680,In_402,In_263);
xnor U681 (N_681,In_748,In_114);
or U682 (N_682,In_945,In_14);
or U683 (N_683,In_259,In_163);
and U684 (N_684,In_885,In_932);
or U685 (N_685,In_805,In_384);
and U686 (N_686,In_821,In_844);
nand U687 (N_687,In_1318,In_893);
or U688 (N_688,In_209,In_1331);
and U689 (N_689,In_854,In_53);
or U690 (N_690,In_685,In_289);
nand U691 (N_691,In_1372,In_273);
and U692 (N_692,In_919,In_189);
nand U693 (N_693,In_429,In_1381);
nor U694 (N_694,In_1109,In_139);
xor U695 (N_695,In_1347,In_927);
or U696 (N_696,In_1228,In_978);
or U697 (N_697,In_1249,In_1329);
or U698 (N_698,In_910,In_1275);
xor U699 (N_699,In_1030,In_224);
xnor U700 (N_700,In_260,In_321);
nand U701 (N_701,In_610,In_58);
xnor U702 (N_702,In_615,In_303);
or U703 (N_703,In_1282,In_915);
or U704 (N_704,In_275,In_499);
nand U705 (N_705,In_160,In_487);
or U706 (N_706,In_1469,In_763);
nor U707 (N_707,In_621,In_689);
and U708 (N_708,In_133,In_1288);
xnor U709 (N_709,In_1406,In_1031);
nand U710 (N_710,In_25,In_193);
nand U711 (N_711,In_804,In_398);
or U712 (N_712,In_404,In_1177);
or U713 (N_713,In_1447,In_497);
nand U714 (N_714,In_585,In_422);
and U715 (N_715,In_349,In_939);
xor U716 (N_716,In_970,In_711);
nor U717 (N_717,In_219,In_1042);
xnor U718 (N_718,In_386,In_500);
or U719 (N_719,In_591,In_323);
nor U720 (N_720,In_1064,In_41);
nand U721 (N_721,In_868,In_524);
nor U722 (N_722,In_253,In_1160);
or U723 (N_723,In_442,In_1467);
or U724 (N_724,In_528,In_920);
xor U725 (N_725,In_338,In_482);
nand U726 (N_726,In_1119,In_494);
nand U727 (N_727,In_962,In_577);
nand U728 (N_728,In_78,In_105);
or U729 (N_729,In_1422,In_957);
xor U730 (N_730,In_1084,In_311);
xor U731 (N_731,In_588,In_1213);
and U732 (N_732,In_1226,In_322);
nand U733 (N_733,In_1188,In_951);
nand U734 (N_734,In_596,In_903);
nor U735 (N_735,In_1134,In_996);
or U736 (N_736,In_1034,In_543);
and U737 (N_737,In_120,In_198);
xor U738 (N_738,In_246,In_797);
nor U739 (N_739,In_470,In_294);
nor U740 (N_740,In_1424,In_60);
and U741 (N_741,In_1352,In_656);
or U742 (N_742,In_174,In_149);
and U743 (N_743,In_63,In_1429);
xor U744 (N_744,In_28,In_737);
and U745 (N_745,In_11,In_702);
and U746 (N_746,In_973,In_746);
xor U747 (N_747,In_986,In_739);
and U748 (N_748,In_720,In_642);
and U749 (N_749,In_1096,In_293);
nor U750 (N_750,In_969,In_494);
and U751 (N_751,In_1377,In_1004);
or U752 (N_752,In_2,In_1272);
xnor U753 (N_753,In_1476,In_31);
nand U754 (N_754,In_882,In_439);
and U755 (N_755,In_291,In_1465);
xnor U756 (N_756,In_360,In_153);
nor U757 (N_757,In_129,In_376);
nand U758 (N_758,In_599,In_986);
nor U759 (N_759,In_1076,In_1309);
nor U760 (N_760,In_820,In_1250);
nor U761 (N_761,In_1464,In_626);
or U762 (N_762,In_1334,In_120);
and U763 (N_763,In_591,In_835);
nand U764 (N_764,In_1278,In_43);
nor U765 (N_765,In_819,In_538);
nor U766 (N_766,In_1436,In_1125);
nor U767 (N_767,In_250,In_725);
or U768 (N_768,In_1096,In_653);
nand U769 (N_769,In_1078,In_776);
and U770 (N_770,In_643,In_868);
nor U771 (N_771,In_592,In_800);
nand U772 (N_772,In_863,In_480);
nor U773 (N_773,In_382,In_41);
or U774 (N_774,In_934,In_254);
xnor U775 (N_775,In_304,In_525);
xnor U776 (N_776,In_1137,In_739);
nor U777 (N_777,In_593,In_73);
and U778 (N_778,In_1473,In_1031);
and U779 (N_779,In_215,In_649);
or U780 (N_780,In_1472,In_923);
or U781 (N_781,In_683,In_779);
and U782 (N_782,In_1398,In_651);
or U783 (N_783,In_1114,In_1077);
nand U784 (N_784,In_1115,In_133);
xor U785 (N_785,In_848,In_776);
nor U786 (N_786,In_759,In_1271);
or U787 (N_787,In_559,In_1035);
nor U788 (N_788,In_269,In_51);
nand U789 (N_789,In_365,In_1146);
nand U790 (N_790,In_1175,In_1307);
or U791 (N_791,In_1137,In_1154);
nand U792 (N_792,In_563,In_1196);
nand U793 (N_793,In_1290,In_152);
and U794 (N_794,In_279,In_1118);
or U795 (N_795,In_413,In_673);
or U796 (N_796,In_575,In_287);
and U797 (N_797,In_303,In_1402);
or U798 (N_798,In_359,In_293);
nand U799 (N_799,In_1191,In_1101);
nor U800 (N_800,In_1458,In_1362);
xor U801 (N_801,In_629,In_669);
or U802 (N_802,In_46,In_335);
nor U803 (N_803,In_944,In_835);
or U804 (N_804,In_1100,In_56);
nand U805 (N_805,In_205,In_145);
nor U806 (N_806,In_1313,In_329);
nor U807 (N_807,In_371,In_472);
and U808 (N_808,In_252,In_1008);
nor U809 (N_809,In_998,In_396);
and U810 (N_810,In_1485,In_98);
nor U811 (N_811,In_1410,In_611);
and U812 (N_812,In_854,In_429);
xnor U813 (N_813,In_1344,In_1326);
nand U814 (N_814,In_1305,In_258);
or U815 (N_815,In_329,In_1300);
and U816 (N_816,In_1077,In_680);
and U817 (N_817,In_1273,In_687);
and U818 (N_818,In_442,In_1052);
nor U819 (N_819,In_435,In_1396);
nor U820 (N_820,In_1495,In_1204);
nor U821 (N_821,In_710,In_1400);
nor U822 (N_822,In_993,In_191);
nand U823 (N_823,In_4,In_229);
nor U824 (N_824,In_474,In_534);
xor U825 (N_825,In_618,In_88);
xor U826 (N_826,In_1382,In_1138);
nand U827 (N_827,In_1387,In_1097);
nor U828 (N_828,In_226,In_497);
and U829 (N_829,In_1067,In_280);
or U830 (N_830,In_617,In_308);
xnor U831 (N_831,In_728,In_245);
nor U832 (N_832,In_883,In_361);
nor U833 (N_833,In_1450,In_673);
and U834 (N_834,In_269,In_1183);
nor U835 (N_835,In_967,In_1057);
and U836 (N_836,In_1149,In_155);
nand U837 (N_837,In_916,In_89);
and U838 (N_838,In_1354,In_1222);
and U839 (N_839,In_640,In_1389);
nand U840 (N_840,In_899,In_122);
nor U841 (N_841,In_233,In_236);
nor U842 (N_842,In_1130,In_371);
nand U843 (N_843,In_585,In_1413);
or U844 (N_844,In_1320,In_620);
or U845 (N_845,In_116,In_360);
or U846 (N_846,In_1022,In_928);
and U847 (N_847,In_975,In_245);
nand U848 (N_848,In_300,In_1101);
nor U849 (N_849,In_9,In_954);
or U850 (N_850,In_159,In_1378);
or U851 (N_851,In_337,In_1417);
nand U852 (N_852,In_974,In_1220);
or U853 (N_853,In_1102,In_359);
nor U854 (N_854,In_959,In_1384);
nand U855 (N_855,In_555,In_1067);
nand U856 (N_856,In_1146,In_1296);
nand U857 (N_857,In_499,In_240);
nand U858 (N_858,In_1208,In_130);
or U859 (N_859,In_533,In_69);
and U860 (N_860,In_374,In_1029);
and U861 (N_861,In_668,In_769);
or U862 (N_862,In_667,In_1339);
nand U863 (N_863,In_261,In_78);
and U864 (N_864,In_738,In_1475);
and U865 (N_865,In_1014,In_1171);
nand U866 (N_866,In_1489,In_265);
and U867 (N_867,In_1084,In_244);
nand U868 (N_868,In_283,In_457);
nand U869 (N_869,In_899,In_862);
nand U870 (N_870,In_701,In_157);
and U871 (N_871,In_906,In_991);
or U872 (N_872,In_516,In_368);
and U873 (N_873,In_721,In_257);
nand U874 (N_874,In_350,In_813);
nand U875 (N_875,In_1071,In_621);
xor U876 (N_876,In_293,In_1185);
xor U877 (N_877,In_1185,In_154);
nor U878 (N_878,In_495,In_284);
nand U879 (N_879,In_1426,In_1363);
or U880 (N_880,In_1186,In_1227);
nand U881 (N_881,In_1461,In_90);
nand U882 (N_882,In_476,In_724);
and U883 (N_883,In_677,In_740);
and U884 (N_884,In_610,In_612);
nand U885 (N_885,In_1396,In_1105);
xnor U886 (N_886,In_356,In_805);
or U887 (N_887,In_289,In_438);
or U888 (N_888,In_402,In_485);
nand U889 (N_889,In_802,In_87);
nor U890 (N_890,In_1173,In_526);
nand U891 (N_891,In_908,In_963);
xor U892 (N_892,In_698,In_47);
xor U893 (N_893,In_370,In_578);
nand U894 (N_894,In_405,In_871);
nand U895 (N_895,In_1372,In_523);
or U896 (N_896,In_324,In_680);
nand U897 (N_897,In_679,In_1241);
or U898 (N_898,In_1164,In_21);
and U899 (N_899,In_839,In_658);
nand U900 (N_900,In_414,In_290);
nor U901 (N_901,In_1241,In_1238);
and U902 (N_902,In_943,In_240);
nor U903 (N_903,In_433,In_726);
nand U904 (N_904,In_665,In_450);
xor U905 (N_905,In_1303,In_1027);
or U906 (N_906,In_1041,In_1264);
and U907 (N_907,In_152,In_553);
or U908 (N_908,In_1293,In_223);
or U909 (N_909,In_1394,In_353);
nand U910 (N_910,In_1033,In_655);
and U911 (N_911,In_1202,In_823);
nand U912 (N_912,In_295,In_945);
and U913 (N_913,In_1148,In_858);
and U914 (N_914,In_408,In_355);
nand U915 (N_915,In_933,In_85);
nor U916 (N_916,In_473,In_390);
nand U917 (N_917,In_489,In_750);
or U918 (N_918,In_179,In_588);
and U919 (N_919,In_154,In_269);
nand U920 (N_920,In_1283,In_1247);
nand U921 (N_921,In_629,In_106);
or U922 (N_922,In_1293,In_961);
nor U923 (N_923,In_731,In_772);
or U924 (N_924,In_824,In_1324);
xor U925 (N_925,In_386,In_1219);
nand U926 (N_926,In_60,In_636);
or U927 (N_927,In_1092,In_685);
nand U928 (N_928,In_351,In_703);
nor U929 (N_929,In_1415,In_828);
and U930 (N_930,In_221,In_267);
nor U931 (N_931,In_312,In_121);
xnor U932 (N_932,In_579,In_1477);
or U933 (N_933,In_606,In_225);
nor U934 (N_934,In_621,In_561);
nand U935 (N_935,In_1101,In_941);
nor U936 (N_936,In_1118,In_953);
or U937 (N_937,In_151,In_240);
and U938 (N_938,In_1227,In_496);
xnor U939 (N_939,In_1069,In_149);
nor U940 (N_940,In_980,In_1488);
and U941 (N_941,In_1084,In_744);
nor U942 (N_942,In_1088,In_1147);
nor U943 (N_943,In_1418,In_574);
and U944 (N_944,In_1237,In_619);
nand U945 (N_945,In_476,In_382);
or U946 (N_946,In_19,In_11);
or U947 (N_947,In_844,In_82);
nand U948 (N_948,In_1137,In_648);
xor U949 (N_949,In_398,In_1458);
nor U950 (N_950,In_1454,In_963);
or U951 (N_951,In_514,In_1347);
xnor U952 (N_952,In_526,In_672);
and U953 (N_953,In_244,In_809);
or U954 (N_954,In_99,In_613);
or U955 (N_955,In_829,In_250);
nor U956 (N_956,In_447,In_399);
and U957 (N_957,In_916,In_743);
nor U958 (N_958,In_1252,In_628);
or U959 (N_959,In_920,In_402);
nand U960 (N_960,In_425,In_751);
nor U961 (N_961,In_366,In_559);
or U962 (N_962,In_1450,In_662);
and U963 (N_963,In_1086,In_211);
or U964 (N_964,In_755,In_408);
or U965 (N_965,In_1077,In_217);
xnor U966 (N_966,In_1174,In_1166);
nand U967 (N_967,In_29,In_726);
nand U968 (N_968,In_1353,In_159);
nand U969 (N_969,In_53,In_1354);
nor U970 (N_970,In_623,In_1120);
or U971 (N_971,In_324,In_1253);
and U972 (N_972,In_1378,In_945);
and U973 (N_973,In_357,In_406);
and U974 (N_974,In_1243,In_1273);
nand U975 (N_975,In_857,In_743);
or U976 (N_976,In_686,In_1081);
nand U977 (N_977,In_897,In_1478);
nand U978 (N_978,In_364,In_101);
nor U979 (N_979,In_937,In_309);
and U980 (N_980,In_221,In_953);
nand U981 (N_981,In_127,In_422);
or U982 (N_982,In_1409,In_250);
or U983 (N_983,In_83,In_755);
nand U984 (N_984,In_1155,In_519);
xnor U985 (N_985,In_889,In_805);
nand U986 (N_986,In_1304,In_311);
and U987 (N_987,In_904,In_378);
nand U988 (N_988,In_1174,In_131);
nor U989 (N_989,In_966,In_151);
or U990 (N_990,In_21,In_979);
nand U991 (N_991,In_136,In_1472);
or U992 (N_992,In_979,In_1047);
nand U993 (N_993,In_242,In_1023);
nor U994 (N_994,In_205,In_950);
and U995 (N_995,In_231,In_1344);
nor U996 (N_996,In_1009,In_939);
and U997 (N_997,In_1190,In_71);
and U998 (N_998,In_581,In_998);
nor U999 (N_999,In_828,In_986);
and U1000 (N_1000,N_425,N_726);
nand U1001 (N_1001,N_739,N_776);
and U1002 (N_1002,N_873,N_701);
nor U1003 (N_1003,N_638,N_67);
and U1004 (N_1004,N_202,N_811);
nor U1005 (N_1005,N_161,N_254);
or U1006 (N_1006,N_824,N_499);
nor U1007 (N_1007,N_595,N_549);
nor U1008 (N_1008,N_479,N_120);
nor U1009 (N_1009,N_505,N_7);
xor U1010 (N_1010,N_673,N_236);
and U1011 (N_1011,N_466,N_548);
nand U1012 (N_1012,N_614,N_582);
nand U1013 (N_1013,N_325,N_795);
or U1014 (N_1014,N_152,N_749);
xor U1015 (N_1015,N_37,N_40);
nand U1016 (N_1016,N_289,N_184);
and U1017 (N_1017,N_200,N_24);
xnor U1018 (N_1018,N_208,N_767);
or U1019 (N_1019,N_344,N_193);
xor U1020 (N_1020,N_970,N_819);
or U1021 (N_1021,N_231,N_287);
and U1022 (N_1022,N_887,N_69);
nand U1023 (N_1023,N_411,N_115);
nor U1024 (N_1024,N_833,N_451);
or U1025 (N_1025,N_654,N_89);
or U1026 (N_1026,N_503,N_492);
nor U1027 (N_1027,N_636,N_41);
nand U1028 (N_1028,N_381,N_319);
and U1029 (N_1029,N_153,N_628);
nand U1030 (N_1030,N_218,N_394);
and U1031 (N_1031,N_408,N_495);
or U1032 (N_1032,N_64,N_511);
and U1033 (N_1033,N_368,N_662);
or U1034 (N_1034,N_642,N_99);
or U1035 (N_1035,N_758,N_409);
nor U1036 (N_1036,N_332,N_295);
nand U1037 (N_1037,N_732,N_509);
and U1038 (N_1038,N_351,N_216);
or U1039 (N_1039,N_723,N_23);
nand U1040 (N_1040,N_306,N_592);
nor U1041 (N_1041,N_555,N_382);
and U1042 (N_1042,N_276,N_817);
or U1043 (N_1043,N_488,N_744);
nand U1044 (N_1044,N_514,N_303);
or U1045 (N_1045,N_27,N_757);
nor U1046 (N_1046,N_682,N_828);
nand U1047 (N_1047,N_455,N_362);
or U1048 (N_1048,N_49,N_170);
nor U1049 (N_1049,N_196,N_489);
or U1050 (N_1050,N_162,N_201);
or U1051 (N_1051,N_794,N_58);
nand U1052 (N_1052,N_279,N_943);
or U1053 (N_1053,N_535,N_852);
or U1054 (N_1054,N_357,N_546);
and U1055 (N_1055,N_888,N_78);
nand U1056 (N_1056,N_10,N_54);
or U1057 (N_1057,N_537,N_727);
and U1058 (N_1058,N_724,N_728);
or U1059 (N_1059,N_653,N_905);
or U1060 (N_1060,N_940,N_646);
nor U1061 (N_1061,N_483,N_796);
or U1062 (N_1062,N_334,N_480);
nand U1063 (N_1063,N_597,N_650);
nand U1064 (N_1064,N_624,N_211);
and U1065 (N_1065,N_150,N_688);
nand U1066 (N_1066,N_615,N_453);
and U1067 (N_1067,N_786,N_11);
or U1068 (N_1068,N_834,N_130);
or U1069 (N_1069,N_219,N_553);
or U1070 (N_1070,N_346,N_174);
and U1071 (N_1071,N_341,N_875);
and U1072 (N_1072,N_730,N_9);
or U1073 (N_1073,N_447,N_526);
nand U1074 (N_1074,N_281,N_707);
or U1075 (N_1075,N_275,N_979);
and U1076 (N_1076,N_826,N_228);
xnor U1077 (N_1077,N_671,N_814);
nor U1078 (N_1078,N_105,N_223);
or U1079 (N_1079,N_482,N_802);
and U1080 (N_1080,N_342,N_191);
nand U1081 (N_1081,N_810,N_770);
nand U1082 (N_1082,N_804,N_156);
nand U1083 (N_1083,N_554,N_73);
and U1084 (N_1084,N_608,N_854);
nand U1085 (N_1085,N_571,N_911);
and U1086 (N_1086,N_370,N_709);
nor U1087 (N_1087,N_348,N_221);
or U1088 (N_1088,N_622,N_415);
and U1089 (N_1089,N_820,N_884);
nor U1090 (N_1090,N_969,N_591);
or U1091 (N_1091,N_630,N_422);
or U1092 (N_1092,N_782,N_383);
and U1093 (N_1093,N_789,N_961);
and U1094 (N_1094,N_111,N_318);
nor U1095 (N_1095,N_542,N_423);
and U1096 (N_1096,N_373,N_987);
and U1097 (N_1097,N_367,N_832);
or U1098 (N_1098,N_915,N_551);
nor U1099 (N_1099,N_570,N_108);
or U1100 (N_1100,N_107,N_683);
nor U1101 (N_1101,N_641,N_541);
nand U1102 (N_1102,N_545,N_155);
or U1103 (N_1103,N_702,N_518);
and U1104 (N_1104,N_151,N_647);
and U1105 (N_1105,N_528,N_890);
xor U1106 (N_1106,N_398,N_585);
nand U1107 (N_1107,N_934,N_572);
nand U1108 (N_1108,N_859,N_574);
nand U1109 (N_1109,N_407,N_611);
and U1110 (N_1110,N_185,N_697);
or U1111 (N_1111,N_777,N_72);
xnor U1112 (N_1112,N_807,N_896);
and U1113 (N_1113,N_791,N_61);
nor U1114 (N_1114,N_224,N_259);
or U1115 (N_1115,N_243,N_720);
nor U1116 (N_1116,N_903,N_544);
and U1117 (N_1117,N_874,N_717);
nand U1118 (N_1118,N_16,N_285);
or U1119 (N_1119,N_298,N_81);
nand U1120 (N_1120,N_138,N_392);
or U1121 (N_1121,N_891,N_696);
nand U1122 (N_1122,N_129,N_240);
and U1123 (N_1123,N_456,N_869);
nand U1124 (N_1124,N_803,N_206);
or U1125 (N_1125,N_606,N_320);
nand U1126 (N_1126,N_780,N_312);
nor U1127 (N_1127,N_265,N_75);
nand U1128 (N_1128,N_908,N_633);
nand U1129 (N_1129,N_360,N_993);
nor U1130 (N_1130,N_388,N_841);
xnor U1131 (N_1131,N_241,N_779);
nor U1132 (N_1132,N_847,N_435);
or U1133 (N_1133,N_670,N_798);
nor U1134 (N_1134,N_17,N_771);
and U1135 (N_1135,N_266,N_271);
nor U1136 (N_1136,N_634,N_858);
nand U1137 (N_1137,N_234,N_924);
and U1138 (N_1138,N_831,N_716);
nand U1139 (N_1139,N_906,N_50);
xnor U1140 (N_1140,N_272,N_563);
and U1141 (N_1141,N_586,N_374);
nand U1142 (N_1142,N_736,N_559);
and U1143 (N_1143,N_645,N_496);
nor U1144 (N_1144,N_666,N_57);
xor U1145 (N_1145,N_255,N_998);
xnor U1146 (N_1146,N_406,N_567);
and U1147 (N_1147,N_439,N_989);
and U1148 (N_1148,N_159,N_643);
nor U1149 (N_1149,N_768,N_898);
nand U1150 (N_1150,N_278,N_909);
nand U1151 (N_1151,N_785,N_816);
or U1152 (N_1152,N_790,N_366);
or U1153 (N_1153,N_267,N_534);
nand U1154 (N_1154,N_166,N_431);
and U1155 (N_1155,N_395,N_253);
or U1156 (N_1156,N_878,N_599);
nor U1157 (N_1157,N_126,N_291);
and U1158 (N_1158,N_45,N_230);
nor U1159 (N_1159,N_763,N_371);
nand U1160 (N_1160,N_521,N_568);
nand U1161 (N_1161,N_941,N_632);
xor U1162 (N_1162,N_601,N_114);
nor U1163 (N_1163,N_335,N_870);
nor U1164 (N_1164,N_617,N_147);
xor U1165 (N_1165,N_593,N_311);
nand U1166 (N_1166,N_583,N_494);
nand U1167 (N_1167,N_775,N_353);
and U1168 (N_1168,N_519,N_48);
and U1169 (N_1169,N_498,N_283);
nor U1170 (N_1170,N_930,N_217);
xor U1171 (N_1171,N_327,N_565);
nand U1172 (N_1172,N_540,N_379);
and U1173 (N_1173,N_486,N_404);
xor U1174 (N_1174,N_957,N_292);
xnor U1175 (N_1175,N_516,N_558);
or U1176 (N_1176,N_310,N_117);
or U1177 (N_1177,N_835,N_385);
nand U1178 (N_1178,N_512,N_765);
nand U1179 (N_1179,N_109,N_317);
nor U1180 (N_1180,N_714,N_995);
and U1181 (N_1181,N_354,N_783);
nand U1182 (N_1182,N_358,N_607);
nor U1183 (N_1183,N_748,N_121);
nand U1184 (N_1184,N_467,N_475);
and U1185 (N_1185,N_119,N_70);
or U1186 (N_1186,N_444,N_245);
and U1187 (N_1187,N_644,N_856);
and U1188 (N_1188,N_880,N_925);
nor U1189 (N_1189,N_524,N_501);
or U1190 (N_1190,N_186,N_754);
nor U1191 (N_1191,N_257,N_38);
nand U1192 (N_1192,N_323,N_840);
xnor U1193 (N_1193,N_487,N_116);
or U1194 (N_1194,N_967,N_146);
nand U1195 (N_1195,N_515,N_756);
or U1196 (N_1196,N_60,N_88);
nand U1197 (N_1197,N_753,N_784);
nor U1198 (N_1198,N_82,N_263);
nor U1199 (N_1199,N_894,N_700);
or U1200 (N_1200,N_440,N_465);
and U1201 (N_1201,N_377,N_421);
nor U1202 (N_1202,N_523,N_350);
or U1203 (N_1203,N_235,N_889);
or U1204 (N_1204,N_806,N_418);
or U1205 (N_1205,N_866,N_13);
or U1206 (N_1206,N_659,N_953);
nand U1207 (N_1207,N_77,N_139);
nor U1208 (N_1208,N_284,N_403);
nor U1209 (N_1209,N_171,N_977);
or U1210 (N_1210,N_990,N_2);
or U1211 (N_1211,N_883,N_68);
or U1212 (N_1212,N_532,N_165);
nand U1213 (N_1213,N_842,N_996);
and U1214 (N_1214,N_25,N_157);
nor U1215 (N_1215,N_110,N_74);
or U1216 (N_1216,N_212,N_297);
nor U1217 (N_1217,N_315,N_436);
or U1218 (N_1218,N_937,N_920);
nand U1219 (N_1219,N_590,N_893);
and U1220 (N_1220,N_735,N_106);
and U1221 (N_1221,N_799,N_131);
nor U1222 (N_1222,N_530,N_427);
or U1223 (N_1223,N_584,N_476);
nand U1224 (N_1224,N_946,N_461);
and U1225 (N_1225,N_743,N_750);
nor U1226 (N_1226,N_364,N_222);
nand U1227 (N_1227,N_91,N_745);
nor U1228 (N_1228,N_945,N_839);
xnor U1229 (N_1229,N_14,N_651);
nor U1230 (N_1230,N_288,N_661);
xnor U1231 (N_1231,N_621,N_649);
and U1232 (N_1232,N_261,N_752);
nand U1233 (N_1233,N_179,N_113);
xnor U1234 (N_1234,N_26,N_849);
nand U1235 (N_1235,N_347,N_207);
nor U1236 (N_1236,N_602,N_746);
nand U1237 (N_1237,N_656,N_47);
nor U1238 (N_1238,N_917,N_102);
and U1239 (N_1239,N_268,N_97);
nor U1240 (N_1240,N_386,N_187);
and U1241 (N_1241,N_604,N_135);
xnor U1242 (N_1242,N_703,N_616);
nand U1243 (N_1243,N_982,N_500);
or U1244 (N_1244,N_349,N_900);
and U1245 (N_1245,N_414,N_902);
nor U1246 (N_1246,N_689,N_539);
nor U1247 (N_1247,N_705,N_913);
and U1248 (N_1248,N_363,N_892);
nand U1249 (N_1249,N_331,N_4);
or U1250 (N_1250,N_952,N_478);
or U1251 (N_1251,N_664,N_19);
or U1252 (N_1252,N_658,N_862);
nor U1253 (N_1253,N_299,N_619);
xor U1254 (N_1254,N_983,N_781);
xor U1255 (N_1255,N_964,N_922);
and U1256 (N_1256,N_426,N_79);
and U1257 (N_1257,N_98,N_313);
nor U1258 (N_1258,N_942,N_424);
and U1259 (N_1259,N_536,N_189);
xor U1260 (N_1260,N_182,N_53);
nand U1261 (N_1261,N_871,N_912);
or U1262 (N_1262,N_137,N_410);
nand U1263 (N_1263,N_837,N_239);
and U1264 (N_1264,N_626,N_927);
and U1265 (N_1265,N_721,N_256);
xor U1266 (N_1266,N_262,N_471);
or U1267 (N_1267,N_657,N_419);
or U1268 (N_1268,N_576,N_329);
nand U1269 (N_1269,N_868,N_742);
or U1270 (N_1270,N_976,N_985);
nor U1271 (N_1271,N_477,N_864);
nand U1272 (N_1272,N_899,N_968);
or U1273 (N_1273,N_845,N_710);
or U1274 (N_1274,N_933,N_956);
nor U1275 (N_1275,N_33,N_788);
and U1276 (N_1276,N_252,N_361);
and U1277 (N_1277,N_1,N_460);
or U1278 (N_1278,N_823,N_144);
nor U1279 (N_1279,N_958,N_397);
nor U1280 (N_1280,N_627,N_39);
nand U1281 (N_1281,N_822,N_20);
xor U1282 (N_1282,N_454,N_877);
and U1283 (N_1283,N_926,N_543);
or U1284 (N_1284,N_220,N_692);
nand U1285 (N_1285,N_35,N_981);
nand U1286 (N_1286,N_324,N_936);
or U1287 (N_1287,N_603,N_588);
and U1288 (N_1288,N_100,N_225);
nor U1289 (N_1289,N_145,N_294);
and U1290 (N_1290,N_508,N_430);
nor U1291 (N_1291,N_813,N_6);
nand U1292 (N_1292,N_391,N_938);
or U1293 (N_1293,N_300,N_733);
or U1294 (N_1294,N_774,N_95);
nor U1295 (N_1295,N_204,N_143);
and U1296 (N_1296,N_339,N_413);
or U1297 (N_1297,N_801,N_274);
and U1298 (N_1298,N_248,N_939);
or U1299 (N_1299,N_134,N_176);
nor U1300 (N_1300,N_984,N_90);
and U1301 (N_1301,N_154,N_715);
nand U1302 (N_1302,N_836,N_797);
and U1303 (N_1303,N_578,N_264);
or U1304 (N_1304,N_125,N_694);
and U1305 (N_1305,N_336,N_429);
or U1306 (N_1306,N_846,N_322);
nor U1307 (N_1307,N_538,N_610);
and U1308 (N_1308,N_389,N_459);
nor U1309 (N_1309,N_376,N_46);
and U1310 (N_1310,N_962,N_506);
and U1311 (N_1311,N_473,N_844);
nand U1312 (N_1312,N_860,N_463);
nor U1313 (N_1313,N_598,N_605);
nand U1314 (N_1314,N_734,N_485);
nor U1315 (N_1315,N_809,N_932);
and U1316 (N_1316,N_773,N_469);
nand U1317 (N_1317,N_199,N_928);
and U1318 (N_1318,N_772,N_44);
nand U1319 (N_1319,N_635,N_302);
nor U1320 (N_1320,N_921,N_674);
nand U1321 (N_1321,N_194,N_850);
or U1322 (N_1322,N_513,N_491);
nor U1323 (N_1323,N_258,N_973);
xnor U1324 (N_1324,N_691,N_183);
nor U1325 (N_1325,N_464,N_246);
nor U1326 (N_1326,N_612,N_988);
or U1327 (N_1327,N_321,N_195);
and U1328 (N_1328,N_55,N_148);
nand U1329 (N_1329,N_882,N_84);
or U1330 (N_1330,N_133,N_269);
or U1331 (N_1331,N_399,N_497);
nand U1332 (N_1332,N_448,N_762);
and U1333 (N_1333,N_520,N_560);
and U1334 (N_1334,N_879,N_764);
and U1335 (N_1335,N_450,N_992);
and U1336 (N_1336,N_980,N_978);
or U1337 (N_1337,N_793,N_569);
or U1338 (N_1338,N_872,N_711);
nand U1339 (N_1339,N_226,N_975);
and U1340 (N_1340,N_755,N_529);
nor U1341 (N_1341,N_690,N_101);
or U1342 (N_1342,N_227,N_618);
and U1343 (N_1343,N_865,N_305);
xor U1344 (N_1344,N_830,N_999);
nor U1345 (N_1345,N_947,N_32);
and U1346 (N_1346,N_173,N_966);
or U1347 (N_1347,N_525,N_140);
and U1348 (N_1348,N_326,N_85);
nand U1349 (N_1349,N_986,N_93);
nor U1350 (N_1350,N_393,N_180);
or U1351 (N_1351,N_695,N_307);
xor U1352 (N_1352,N_449,N_759);
or U1353 (N_1353,N_270,N_242);
nand U1354 (N_1354,N_722,N_507);
nor U1355 (N_1355,N_867,N_778);
or U1356 (N_1356,N_719,N_31);
nor U1357 (N_1357,N_198,N_34);
nor U1358 (N_1358,N_63,N_290);
or U1359 (N_1359,N_71,N_5);
and U1360 (N_1360,N_693,N_343);
xnor U1361 (N_1361,N_564,N_678);
or U1362 (N_1362,N_175,N_600);
nand U1363 (N_1363,N_330,N_623);
and U1364 (N_1364,N_594,N_587);
nand U1365 (N_1365,N_197,N_965);
or U1366 (N_1366,N_960,N_522);
and U1367 (N_1367,N_205,N_337);
or U1368 (N_1368,N_92,N_484);
or U1369 (N_1369,N_401,N_760);
and U1370 (N_1370,N_229,N_686);
xor U1371 (N_1371,N_527,N_396);
xnor U1372 (N_1372,N_766,N_997);
or U1373 (N_1373,N_445,N_687);
and U1374 (N_1374,N_713,N_954);
nand U1375 (N_1375,N_729,N_675);
xor U1376 (N_1376,N_123,N_169);
nor U1377 (N_1377,N_356,N_167);
nand U1378 (N_1378,N_918,N_280);
xor U1379 (N_1379,N_213,N_128);
nand U1380 (N_1380,N_127,N_629);
nand U1381 (N_1381,N_96,N_316);
or U1382 (N_1382,N_631,N_718);
nand U1383 (N_1383,N_493,N_384);
and U1384 (N_1384,N_561,N_359);
nor U1385 (N_1385,N_375,N_405);
xnor U1386 (N_1386,N_818,N_437);
nor U1387 (N_1387,N_712,N_94);
nand U1388 (N_1388,N_446,N_669);
xnor U1389 (N_1389,N_800,N_141);
and U1390 (N_1390,N_725,N_149);
and U1391 (N_1391,N_738,N_249);
or U1392 (N_1392,N_706,N_441);
or U1393 (N_1393,N_369,N_52);
and U1394 (N_1394,N_637,N_390);
nand U1395 (N_1395,N_308,N_103);
and U1396 (N_1396,N_639,N_28);
and U1397 (N_1397,N_432,N_438);
or U1398 (N_1398,N_0,N_955);
or U1399 (N_1399,N_827,N_950);
nand U1400 (N_1400,N_681,N_552);
nor U1401 (N_1401,N_462,N_620);
or U1402 (N_1402,N_660,N_829);
or U1403 (N_1403,N_136,N_843);
nand U1404 (N_1404,N_769,N_190);
xnor U1405 (N_1405,N_36,N_277);
and U1406 (N_1406,N_314,N_247);
nor U1407 (N_1407,N_273,N_677);
nand U1408 (N_1408,N_66,N_886);
or U1409 (N_1409,N_931,N_417);
nand U1410 (N_1410,N_881,N_8);
and U1411 (N_1411,N_472,N_244);
nand U1412 (N_1412,N_181,N_238);
or U1413 (N_1413,N_365,N_761);
and U1414 (N_1414,N_345,N_557);
or U1415 (N_1415,N_914,N_29);
nor U1416 (N_1416,N_87,N_805);
nand U1417 (N_1417,N_672,N_355);
nor U1418 (N_1418,N_580,N_625);
or U1419 (N_1419,N_338,N_470);
nor U1420 (N_1420,N_192,N_160);
or U1421 (N_1421,N_210,N_80);
and U1422 (N_1422,N_203,N_885);
xor U1423 (N_1423,N_504,N_340);
nor U1424 (N_1424,N_118,N_22);
or U1425 (N_1425,N_163,N_412);
or U1426 (N_1426,N_589,N_974);
and U1427 (N_1427,N_517,N_468);
nand U1428 (N_1428,N_502,N_851);
and U1429 (N_1429,N_86,N_352);
and U1430 (N_1430,N_876,N_51);
or U1431 (N_1431,N_853,N_944);
and U1432 (N_1432,N_609,N_333);
nand U1433 (N_1433,N_907,N_232);
and U1434 (N_1434,N_910,N_56);
nor U1435 (N_1435,N_474,N_923);
or U1436 (N_1436,N_815,N_533);
nor U1437 (N_1437,N_655,N_663);
nand U1438 (N_1438,N_665,N_648);
and U1439 (N_1439,N_698,N_104);
or U1440 (N_1440,N_65,N_296);
nor U1441 (N_1441,N_897,N_177);
or U1442 (N_1442,N_935,N_821);
or U1443 (N_1443,N_904,N_42);
nor U1444 (N_1444,N_458,N_948);
nor U1445 (N_1445,N_579,N_43);
and U1446 (N_1446,N_158,N_963);
and U1447 (N_1447,N_59,N_510);
nand U1448 (N_1448,N_699,N_452);
and U1449 (N_1449,N_848,N_12);
nor U1450 (N_1450,N_838,N_215);
or U1451 (N_1451,N_282,N_142);
xor U1452 (N_1452,N_420,N_684);
xnor U1453 (N_1453,N_188,N_15);
nand U1454 (N_1454,N_372,N_575);
or U1455 (N_1455,N_613,N_951);
nor U1456 (N_1456,N_83,N_3);
nand U1457 (N_1457,N_30,N_237);
or U1458 (N_1458,N_680,N_667);
and U1459 (N_1459,N_566,N_741);
nand U1460 (N_1460,N_443,N_562);
or U1461 (N_1461,N_676,N_233);
and U1462 (N_1462,N_18,N_679);
xor U1463 (N_1463,N_573,N_808);
or U1464 (N_1464,N_402,N_214);
and U1465 (N_1465,N_704,N_971);
nor U1466 (N_1466,N_972,N_164);
and U1467 (N_1467,N_434,N_577);
or U1468 (N_1468,N_301,N_251);
and U1469 (N_1469,N_916,N_708);
nor U1470 (N_1470,N_328,N_919);
and U1471 (N_1471,N_792,N_428);
nand U1472 (N_1472,N_178,N_861);
nand U1473 (N_1473,N_652,N_685);
and U1474 (N_1474,N_901,N_112);
and U1475 (N_1475,N_668,N_209);
or U1476 (N_1476,N_731,N_378);
nor U1477 (N_1477,N_387,N_751);
xor U1478 (N_1478,N_433,N_293);
nor U1479 (N_1479,N_857,N_124);
nor U1480 (N_1480,N_286,N_122);
or U1481 (N_1481,N_400,N_416);
and U1482 (N_1482,N_949,N_991);
nand U1483 (N_1483,N_442,N_812);
or U1484 (N_1484,N_929,N_490);
and U1485 (N_1485,N_260,N_747);
xnor U1486 (N_1486,N_596,N_994);
nand U1487 (N_1487,N_787,N_855);
or U1488 (N_1488,N_457,N_380);
or U1489 (N_1489,N_863,N_547);
or U1490 (N_1490,N_132,N_959);
or U1491 (N_1491,N_581,N_825);
and U1492 (N_1492,N_740,N_309);
or U1493 (N_1493,N_556,N_250);
and U1494 (N_1494,N_737,N_172);
xnor U1495 (N_1495,N_168,N_550);
nor U1496 (N_1496,N_531,N_76);
and U1497 (N_1497,N_481,N_62);
or U1498 (N_1498,N_304,N_640);
and U1499 (N_1499,N_21,N_895);
or U1500 (N_1500,N_236,N_577);
xor U1501 (N_1501,N_909,N_38);
nor U1502 (N_1502,N_666,N_901);
and U1503 (N_1503,N_38,N_624);
nor U1504 (N_1504,N_196,N_834);
nand U1505 (N_1505,N_839,N_793);
xnor U1506 (N_1506,N_705,N_364);
or U1507 (N_1507,N_140,N_845);
nor U1508 (N_1508,N_857,N_757);
nand U1509 (N_1509,N_980,N_560);
nor U1510 (N_1510,N_609,N_154);
xnor U1511 (N_1511,N_296,N_717);
nand U1512 (N_1512,N_661,N_310);
xnor U1513 (N_1513,N_807,N_441);
or U1514 (N_1514,N_32,N_397);
and U1515 (N_1515,N_142,N_441);
or U1516 (N_1516,N_334,N_501);
nor U1517 (N_1517,N_890,N_415);
nor U1518 (N_1518,N_353,N_132);
nor U1519 (N_1519,N_713,N_866);
or U1520 (N_1520,N_83,N_229);
xnor U1521 (N_1521,N_541,N_108);
or U1522 (N_1522,N_438,N_278);
xor U1523 (N_1523,N_310,N_528);
and U1524 (N_1524,N_228,N_707);
and U1525 (N_1525,N_171,N_63);
xnor U1526 (N_1526,N_961,N_632);
or U1527 (N_1527,N_204,N_653);
and U1528 (N_1528,N_940,N_643);
or U1529 (N_1529,N_877,N_114);
xor U1530 (N_1530,N_892,N_789);
and U1531 (N_1531,N_902,N_464);
nand U1532 (N_1532,N_971,N_312);
nand U1533 (N_1533,N_997,N_642);
or U1534 (N_1534,N_950,N_181);
nor U1535 (N_1535,N_528,N_986);
and U1536 (N_1536,N_224,N_111);
nor U1537 (N_1537,N_381,N_14);
or U1538 (N_1538,N_150,N_259);
and U1539 (N_1539,N_925,N_240);
or U1540 (N_1540,N_633,N_399);
nand U1541 (N_1541,N_852,N_864);
nor U1542 (N_1542,N_738,N_655);
or U1543 (N_1543,N_627,N_229);
and U1544 (N_1544,N_196,N_753);
and U1545 (N_1545,N_298,N_209);
xor U1546 (N_1546,N_201,N_336);
or U1547 (N_1547,N_955,N_993);
nand U1548 (N_1548,N_328,N_91);
and U1549 (N_1549,N_493,N_480);
nand U1550 (N_1550,N_21,N_307);
or U1551 (N_1551,N_111,N_259);
and U1552 (N_1552,N_745,N_323);
nor U1553 (N_1553,N_708,N_145);
nor U1554 (N_1554,N_146,N_548);
nor U1555 (N_1555,N_498,N_566);
and U1556 (N_1556,N_112,N_794);
or U1557 (N_1557,N_391,N_591);
nand U1558 (N_1558,N_609,N_309);
or U1559 (N_1559,N_490,N_733);
nand U1560 (N_1560,N_213,N_332);
or U1561 (N_1561,N_743,N_738);
and U1562 (N_1562,N_99,N_333);
and U1563 (N_1563,N_869,N_115);
and U1564 (N_1564,N_622,N_854);
nand U1565 (N_1565,N_120,N_920);
xnor U1566 (N_1566,N_934,N_730);
xor U1567 (N_1567,N_750,N_924);
xor U1568 (N_1568,N_352,N_77);
nand U1569 (N_1569,N_416,N_729);
or U1570 (N_1570,N_383,N_271);
nor U1571 (N_1571,N_784,N_641);
xor U1572 (N_1572,N_288,N_922);
nor U1573 (N_1573,N_152,N_379);
nor U1574 (N_1574,N_609,N_290);
nand U1575 (N_1575,N_735,N_118);
or U1576 (N_1576,N_570,N_598);
xnor U1577 (N_1577,N_163,N_211);
nand U1578 (N_1578,N_517,N_265);
nand U1579 (N_1579,N_549,N_191);
xnor U1580 (N_1580,N_409,N_297);
and U1581 (N_1581,N_153,N_279);
or U1582 (N_1582,N_521,N_360);
nand U1583 (N_1583,N_855,N_375);
nand U1584 (N_1584,N_596,N_444);
and U1585 (N_1585,N_309,N_244);
nand U1586 (N_1586,N_893,N_945);
or U1587 (N_1587,N_641,N_988);
nor U1588 (N_1588,N_357,N_750);
or U1589 (N_1589,N_490,N_87);
and U1590 (N_1590,N_187,N_650);
nand U1591 (N_1591,N_346,N_571);
nor U1592 (N_1592,N_764,N_125);
nor U1593 (N_1593,N_809,N_30);
nor U1594 (N_1594,N_20,N_403);
xnor U1595 (N_1595,N_114,N_609);
and U1596 (N_1596,N_753,N_63);
xnor U1597 (N_1597,N_377,N_834);
and U1598 (N_1598,N_765,N_99);
xor U1599 (N_1599,N_300,N_590);
or U1600 (N_1600,N_869,N_684);
and U1601 (N_1601,N_22,N_177);
or U1602 (N_1602,N_427,N_390);
nand U1603 (N_1603,N_466,N_726);
xor U1604 (N_1604,N_572,N_435);
nor U1605 (N_1605,N_818,N_198);
and U1606 (N_1606,N_606,N_955);
or U1607 (N_1607,N_317,N_23);
nand U1608 (N_1608,N_273,N_194);
xnor U1609 (N_1609,N_952,N_552);
or U1610 (N_1610,N_831,N_420);
nand U1611 (N_1611,N_111,N_696);
nor U1612 (N_1612,N_865,N_934);
or U1613 (N_1613,N_505,N_986);
or U1614 (N_1614,N_818,N_668);
nor U1615 (N_1615,N_786,N_79);
and U1616 (N_1616,N_85,N_477);
or U1617 (N_1617,N_298,N_177);
or U1618 (N_1618,N_653,N_389);
nand U1619 (N_1619,N_989,N_81);
or U1620 (N_1620,N_618,N_252);
nand U1621 (N_1621,N_899,N_456);
or U1622 (N_1622,N_254,N_655);
nor U1623 (N_1623,N_193,N_503);
nor U1624 (N_1624,N_495,N_537);
and U1625 (N_1625,N_539,N_765);
or U1626 (N_1626,N_513,N_151);
or U1627 (N_1627,N_198,N_346);
nand U1628 (N_1628,N_801,N_726);
and U1629 (N_1629,N_608,N_89);
nand U1630 (N_1630,N_231,N_58);
nor U1631 (N_1631,N_881,N_72);
nand U1632 (N_1632,N_235,N_676);
or U1633 (N_1633,N_512,N_756);
nand U1634 (N_1634,N_272,N_328);
or U1635 (N_1635,N_717,N_46);
or U1636 (N_1636,N_200,N_768);
and U1637 (N_1637,N_895,N_891);
xor U1638 (N_1638,N_638,N_20);
nand U1639 (N_1639,N_43,N_756);
and U1640 (N_1640,N_715,N_383);
nand U1641 (N_1641,N_543,N_765);
nor U1642 (N_1642,N_180,N_889);
and U1643 (N_1643,N_446,N_397);
and U1644 (N_1644,N_309,N_867);
nand U1645 (N_1645,N_773,N_614);
or U1646 (N_1646,N_67,N_899);
or U1647 (N_1647,N_920,N_318);
and U1648 (N_1648,N_560,N_757);
and U1649 (N_1649,N_514,N_302);
xnor U1650 (N_1650,N_10,N_127);
and U1651 (N_1651,N_853,N_922);
and U1652 (N_1652,N_32,N_799);
nor U1653 (N_1653,N_386,N_259);
and U1654 (N_1654,N_937,N_902);
and U1655 (N_1655,N_140,N_996);
xor U1656 (N_1656,N_600,N_666);
or U1657 (N_1657,N_109,N_186);
or U1658 (N_1658,N_917,N_626);
nand U1659 (N_1659,N_340,N_619);
or U1660 (N_1660,N_250,N_99);
nor U1661 (N_1661,N_64,N_577);
and U1662 (N_1662,N_497,N_881);
and U1663 (N_1663,N_194,N_744);
and U1664 (N_1664,N_574,N_403);
or U1665 (N_1665,N_300,N_354);
and U1666 (N_1666,N_749,N_521);
or U1667 (N_1667,N_618,N_714);
and U1668 (N_1668,N_801,N_14);
nand U1669 (N_1669,N_14,N_944);
nand U1670 (N_1670,N_472,N_660);
nor U1671 (N_1671,N_462,N_148);
or U1672 (N_1672,N_871,N_48);
xor U1673 (N_1673,N_314,N_875);
and U1674 (N_1674,N_371,N_228);
nand U1675 (N_1675,N_292,N_233);
nor U1676 (N_1676,N_995,N_39);
nand U1677 (N_1677,N_714,N_654);
nor U1678 (N_1678,N_375,N_275);
nand U1679 (N_1679,N_140,N_349);
and U1680 (N_1680,N_860,N_584);
and U1681 (N_1681,N_463,N_715);
nand U1682 (N_1682,N_501,N_678);
or U1683 (N_1683,N_332,N_277);
and U1684 (N_1684,N_463,N_586);
nor U1685 (N_1685,N_230,N_507);
nor U1686 (N_1686,N_880,N_273);
xnor U1687 (N_1687,N_440,N_913);
nand U1688 (N_1688,N_105,N_75);
nor U1689 (N_1689,N_579,N_344);
and U1690 (N_1690,N_375,N_7);
and U1691 (N_1691,N_800,N_782);
and U1692 (N_1692,N_654,N_341);
and U1693 (N_1693,N_79,N_146);
nor U1694 (N_1694,N_562,N_281);
xor U1695 (N_1695,N_95,N_517);
or U1696 (N_1696,N_165,N_476);
or U1697 (N_1697,N_983,N_387);
or U1698 (N_1698,N_975,N_697);
nand U1699 (N_1699,N_70,N_820);
and U1700 (N_1700,N_268,N_853);
nor U1701 (N_1701,N_975,N_924);
and U1702 (N_1702,N_857,N_300);
nor U1703 (N_1703,N_912,N_836);
or U1704 (N_1704,N_840,N_624);
and U1705 (N_1705,N_66,N_802);
or U1706 (N_1706,N_945,N_54);
and U1707 (N_1707,N_469,N_984);
xnor U1708 (N_1708,N_596,N_435);
and U1709 (N_1709,N_984,N_975);
xnor U1710 (N_1710,N_7,N_496);
nand U1711 (N_1711,N_853,N_859);
nor U1712 (N_1712,N_494,N_114);
nand U1713 (N_1713,N_914,N_486);
and U1714 (N_1714,N_461,N_469);
nor U1715 (N_1715,N_685,N_516);
nor U1716 (N_1716,N_890,N_475);
or U1717 (N_1717,N_846,N_695);
nand U1718 (N_1718,N_77,N_308);
or U1719 (N_1719,N_359,N_942);
and U1720 (N_1720,N_907,N_420);
and U1721 (N_1721,N_535,N_822);
and U1722 (N_1722,N_439,N_91);
xnor U1723 (N_1723,N_243,N_93);
xor U1724 (N_1724,N_792,N_789);
nand U1725 (N_1725,N_357,N_854);
nor U1726 (N_1726,N_888,N_544);
and U1727 (N_1727,N_993,N_216);
nand U1728 (N_1728,N_693,N_594);
or U1729 (N_1729,N_774,N_293);
nor U1730 (N_1730,N_190,N_412);
and U1731 (N_1731,N_572,N_778);
or U1732 (N_1732,N_321,N_3);
and U1733 (N_1733,N_647,N_187);
nor U1734 (N_1734,N_104,N_94);
or U1735 (N_1735,N_548,N_708);
nor U1736 (N_1736,N_17,N_623);
and U1737 (N_1737,N_378,N_579);
or U1738 (N_1738,N_555,N_271);
nand U1739 (N_1739,N_101,N_575);
and U1740 (N_1740,N_727,N_14);
or U1741 (N_1741,N_114,N_911);
nor U1742 (N_1742,N_131,N_268);
nor U1743 (N_1743,N_88,N_741);
nand U1744 (N_1744,N_713,N_22);
or U1745 (N_1745,N_270,N_403);
xor U1746 (N_1746,N_459,N_375);
nor U1747 (N_1747,N_257,N_768);
xnor U1748 (N_1748,N_113,N_57);
nand U1749 (N_1749,N_113,N_370);
nor U1750 (N_1750,N_491,N_480);
and U1751 (N_1751,N_857,N_530);
nand U1752 (N_1752,N_353,N_631);
nand U1753 (N_1753,N_554,N_121);
nand U1754 (N_1754,N_189,N_232);
nand U1755 (N_1755,N_49,N_190);
nor U1756 (N_1756,N_678,N_471);
or U1757 (N_1757,N_241,N_672);
nand U1758 (N_1758,N_752,N_872);
and U1759 (N_1759,N_849,N_684);
nor U1760 (N_1760,N_82,N_336);
nor U1761 (N_1761,N_748,N_435);
and U1762 (N_1762,N_538,N_971);
and U1763 (N_1763,N_683,N_651);
and U1764 (N_1764,N_967,N_274);
or U1765 (N_1765,N_648,N_961);
nor U1766 (N_1766,N_993,N_861);
nor U1767 (N_1767,N_354,N_976);
and U1768 (N_1768,N_508,N_488);
and U1769 (N_1769,N_366,N_906);
nor U1770 (N_1770,N_538,N_139);
and U1771 (N_1771,N_938,N_820);
nor U1772 (N_1772,N_336,N_815);
and U1773 (N_1773,N_669,N_808);
or U1774 (N_1774,N_395,N_988);
or U1775 (N_1775,N_721,N_735);
or U1776 (N_1776,N_957,N_585);
and U1777 (N_1777,N_236,N_924);
nor U1778 (N_1778,N_845,N_262);
nand U1779 (N_1779,N_820,N_449);
or U1780 (N_1780,N_556,N_322);
xor U1781 (N_1781,N_236,N_483);
nor U1782 (N_1782,N_817,N_822);
or U1783 (N_1783,N_159,N_371);
nor U1784 (N_1784,N_192,N_436);
and U1785 (N_1785,N_188,N_606);
or U1786 (N_1786,N_792,N_500);
nand U1787 (N_1787,N_438,N_186);
nand U1788 (N_1788,N_506,N_160);
nand U1789 (N_1789,N_474,N_375);
nand U1790 (N_1790,N_725,N_330);
or U1791 (N_1791,N_382,N_510);
or U1792 (N_1792,N_603,N_288);
and U1793 (N_1793,N_963,N_560);
nor U1794 (N_1794,N_179,N_524);
or U1795 (N_1795,N_623,N_160);
or U1796 (N_1796,N_971,N_795);
or U1797 (N_1797,N_351,N_25);
xnor U1798 (N_1798,N_749,N_323);
or U1799 (N_1799,N_294,N_107);
nand U1800 (N_1800,N_229,N_559);
nor U1801 (N_1801,N_371,N_311);
and U1802 (N_1802,N_354,N_208);
and U1803 (N_1803,N_377,N_796);
and U1804 (N_1804,N_575,N_481);
nor U1805 (N_1805,N_737,N_221);
nor U1806 (N_1806,N_457,N_383);
nor U1807 (N_1807,N_736,N_607);
nand U1808 (N_1808,N_154,N_490);
xnor U1809 (N_1809,N_815,N_796);
nor U1810 (N_1810,N_627,N_813);
or U1811 (N_1811,N_192,N_948);
nand U1812 (N_1812,N_320,N_943);
and U1813 (N_1813,N_540,N_545);
nor U1814 (N_1814,N_296,N_292);
or U1815 (N_1815,N_492,N_608);
or U1816 (N_1816,N_601,N_647);
nor U1817 (N_1817,N_218,N_352);
nand U1818 (N_1818,N_166,N_283);
nor U1819 (N_1819,N_545,N_0);
and U1820 (N_1820,N_895,N_316);
nand U1821 (N_1821,N_287,N_595);
and U1822 (N_1822,N_691,N_840);
nand U1823 (N_1823,N_616,N_964);
nor U1824 (N_1824,N_373,N_897);
xor U1825 (N_1825,N_84,N_421);
or U1826 (N_1826,N_929,N_993);
xor U1827 (N_1827,N_298,N_369);
and U1828 (N_1828,N_92,N_865);
or U1829 (N_1829,N_155,N_516);
nand U1830 (N_1830,N_122,N_756);
nand U1831 (N_1831,N_539,N_221);
nor U1832 (N_1832,N_540,N_781);
or U1833 (N_1833,N_438,N_701);
and U1834 (N_1834,N_933,N_762);
and U1835 (N_1835,N_879,N_669);
nand U1836 (N_1836,N_541,N_100);
nor U1837 (N_1837,N_939,N_902);
nand U1838 (N_1838,N_224,N_616);
or U1839 (N_1839,N_609,N_578);
nor U1840 (N_1840,N_797,N_463);
nand U1841 (N_1841,N_730,N_977);
nor U1842 (N_1842,N_354,N_158);
nand U1843 (N_1843,N_886,N_380);
and U1844 (N_1844,N_717,N_969);
nor U1845 (N_1845,N_681,N_414);
xnor U1846 (N_1846,N_963,N_609);
nor U1847 (N_1847,N_766,N_424);
xnor U1848 (N_1848,N_949,N_319);
or U1849 (N_1849,N_674,N_900);
nand U1850 (N_1850,N_364,N_990);
nor U1851 (N_1851,N_176,N_934);
or U1852 (N_1852,N_583,N_43);
nand U1853 (N_1853,N_393,N_782);
or U1854 (N_1854,N_306,N_36);
or U1855 (N_1855,N_235,N_32);
or U1856 (N_1856,N_386,N_257);
nor U1857 (N_1857,N_681,N_675);
nor U1858 (N_1858,N_95,N_730);
nor U1859 (N_1859,N_436,N_832);
and U1860 (N_1860,N_886,N_622);
xor U1861 (N_1861,N_628,N_482);
nand U1862 (N_1862,N_641,N_502);
and U1863 (N_1863,N_815,N_17);
and U1864 (N_1864,N_697,N_314);
and U1865 (N_1865,N_348,N_822);
nand U1866 (N_1866,N_173,N_285);
or U1867 (N_1867,N_257,N_736);
nor U1868 (N_1868,N_696,N_367);
xor U1869 (N_1869,N_238,N_641);
or U1870 (N_1870,N_331,N_718);
xor U1871 (N_1871,N_712,N_239);
nand U1872 (N_1872,N_585,N_731);
nor U1873 (N_1873,N_227,N_478);
xor U1874 (N_1874,N_311,N_952);
xnor U1875 (N_1875,N_371,N_53);
nand U1876 (N_1876,N_912,N_90);
nor U1877 (N_1877,N_643,N_169);
and U1878 (N_1878,N_846,N_943);
nor U1879 (N_1879,N_944,N_23);
or U1880 (N_1880,N_62,N_386);
xnor U1881 (N_1881,N_345,N_496);
xnor U1882 (N_1882,N_499,N_334);
and U1883 (N_1883,N_752,N_454);
and U1884 (N_1884,N_642,N_269);
or U1885 (N_1885,N_782,N_168);
xnor U1886 (N_1886,N_720,N_340);
nand U1887 (N_1887,N_385,N_252);
nand U1888 (N_1888,N_88,N_489);
and U1889 (N_1889,N_851,N_35);
and U1890 (N_1890,N_862,N_473);
nor U1891 (N_1891,N_463,N_71);
nor U1892 (N_1892,N_935,N_398);
nand U1893 (N_1893,N_330,N_55);
and U1894 (N_1894,N_407,N_185);
or U1895 (N_1895,N_723,N_71);
and U1896 (N_1896,N_170,N_124);
or U1897 (N_1897,N_213,N_713);
nor U1898 (N_1898,N_129,N_678);
nor U1899 (N_1899,N_299,N_96);
nand U1900 (N_1900,N_702,N_255);
or U1901 (N_1901,N_691,N_313);
nor U1902 (N_1902,N_931,N_59);
xnor U1903 (N_1903,N_129,N_5);
or U1904 (N_1904,N_384,N_799);
xor U1905 (N_1905,N_57,N_886);
and U1906 (N_1906,N_493,N_241);
or U1907 (N_1907,N_424,N_230);
xnor U1908 (N_1908,N_449,N_163);
or U1909 (N_1909,N_62,N_182);
nand U1910 (N_1910,N_709,N_347);
or U1911 (N_1911,N_554,N_511);
or U1912 (N_1912,N_172,N_32);
nor U1913 (N_1913,N_669,N_117);
or U1914 (N_1914,N_678,N_491);
or U1915 (N_1915,N_254,N_544);
and U1916 (N_1916,N_932,N_900);
nor U1917 (N_1917,N_953,N_483);
or U1918 (N_1918,N_297,N_641);
xor U1919 (N_1919,N_590,N_705);
nor U1920 (N_1920,N_596,N_903);
nor U1921 (N_1921,N_965,N_482);
nor U1922 (N_1922,N_744,N_965);
or U1923 (N_1923,N_952,N_565);
nand U1924 (N_1924,N_437,N_339);
nor U1925 (N_1925,N_469,N_856);
or U1926 (N_1926,N_650,N_829);
or U1927 (N_1927,N_68,N_548);
and U1928 (N_1928,N_89,N_329);
or U1929 (N_1929,N_880,N_630);
and U1930 (N_1930,N_822,N_457);
nand U1931 (N_1931,N_6,N_127);
xnor U1932 (N_1932,N_323,N_195);
or U1933 (N_1933,N_654,N_20);
nor U1934 (N_1934,N_653,N_679);
or U1935 (N_1935,N_191,N_7);
nor U1936 (N_1936,N_572,N_832);
xor U1937 (N_1937,N_251,N_918);
and U1938 (N_1938,N_660,N_938);
and U1939 (N_1939,N_577,N_748);
or U1940 (N_1940,N_606,N_858);
xnor U1941 (N_1941,N_581,N_809);
or U1942 (N_1942,N_25,N_452);
nand U1943 (N_1943,N_745,N_210);
nor U1944 (N_1944,N_175,N_388);
nand U1945 (N_1945,N_234,N_694);
nand U1946 (N_1946,N_865,N_390);
nand U1947 (N_1947,N_586,N_106);
nor U1948 (N_1948,N_679,N_758);
xnor U1949 (N_1949,N_33,N_514);
and U1950 (N_1950,N_340,N_985);
xor U1951 (N_1951,N_998,N_28);
nor U1952 (N_1952,N_221,N_545);
nand U1953 (N_1953,N_146,N_748);
nor U1954 (N_1954,N_652,N_603);
nand U1955 (N_1955,N_475,N_817);
and U1956 (N_1956,N_366,N_894);
xnor U1957 (N_1957,N_453,N_882);
nor U1958 (N_1958,N_413,N_289);
and U1959 (N_1959,N_655,N_245);
nand U1960 (N_1960,N_441,N_828);
xnor U1961 (N_1961,N_475,N_166);
or U1962 (N_1962,N_17,N_994);
nor U1963 (N_1963,N_674,N_953);
nor U1964 (N_1964,N_439,N_919);
and U1965 (N_1965,N_700,N_818);
or U1966 (N_1966,N_89,N_698);
nand U1967 (N_1967,N_637,N_365);
nor U1968 (N_1968,N_389,N_471);
nand U1969 (N_1969,N_159,N_866);
xnor U1970 (N_1970,N_143,N_658);
xnor U1971 (N_1971,N_449,N_519);
nor U1972 (N_1972,N_50,N_596);
xor U1973 (N_1973,N_665,N_582);
or U1974 (N_1974,N_650,N_610);
and U1975 (N_1975,N_565,N_88);
and U1976 (N_1976,N_162,N_806);
nor U1977 (N_1977,N_315,N_27);
nor U1978 (N_1978,N_690,N_42);
nor U1979 (N_1979,N_154,N_634);
xnor U1980 (N_1980,N_382,N_193);
or U1981 (N_1981,N_665,N_354);
xnor U1982 (N_1982,N_104,N_604);
nor U1983 (N_1983,N_127,N_956);
xor U1984 (N_1984,N_7,N_437);
nand U1985 (N_1985,N_620,N_548);
nand U1986 (N_1986,N_124,N_286);
or U1987 (N_1987,N_469,N_279);
nor U1988 (N_1988,N_210,N_343);
nor U1989 (N_1989,N_625,N_968);
nor U1990 (N_1990,N_835,N_347);
nand U1991 (N_1991,N_488,N_57);
nor U1992 (N_1992,N_155,N_590);
and U1993 (N_1993,N_393,N_528);
nor U1994 (N_1994,N_631,N_581);
and U1995 (N_1995,N_755,N_565);
or U1996 (N_1996,N_672,N_928);
or U1997 (N_1997,N_237,N_221);
nand U1998 (N_1998,N_684,N_772);
nor U1999 (N_1999,N_899,N_951);
nor U2000 (N_2000,N_1331,N_1288);
and U2001 (N_2001,N_1004,N_1676);
nor U2002 (N_2002,N_1069,N_1140);
nor U2003 (N_2003,N_1397,N_1709);
or U2004 (N_2004,N_1792,N_1366);
or U2005 (N_2005,N_1728,N_1243);
nand U2006 (N_2006,N_1665,N_1409);
or U2007 (N_2007,N_1099,N_1384);
xor U2008 (N_2008,N_1463,N_1458);
and U2009 (N_2009,N_1509,N_1442);
xor U2010 (N_2010,N_1577,N_1159);
nor U2011 (N_2011,N_1008,N_1380);
and U2012 (N_2012,N_1926,N_1937);
nand U2013 (N_2013,N_1848,N_1347);
or U2014 (N_2014,N_1921,N_1217);
or U2015 (N_2015,N_1328,N_1223);
or U2016 (N_2016,N_1268,N_1492);
nand U2017 (N_2017,N_1662,N_1777);
nor U2018 (N_2018,N_1459,N_1659);
nand U2019 (N_2019,N_1947,N_1863);
and U2020 (N_2020,N_1918,N_1977);
nor U2021 (N_2021,N_1816,N_1600);
or U2022 (N_2022,N_1575,N_1833);
nor U2023 (N_2023,N_1529,N_1982);
or U2024 (N_2024,N_1359,N_1907);
and U2025 (N_2025,N_1252,N_1202);
xnor U2026 (N_2026,N_1299,N_1681);
or U2027 (N_2027,N_1456,N_1788);
or U2028 (N_2028,N_1352,N_1037);
nor U2029 (N_2029,N_1919,N_1087);
or U2030 (N_2030,N_1849,N_1995);
or U2031 (N_2031,N_1689,N_1856);
nor U2032 (N_2032,N_1307,N_1452);
nand U2033 (N_2033,N_1860,N_1864);
or U2034 (N_2034,N_1758,N_1542);
or U2035 (N_2035,N_1284,N_1932);
or U2036 (N_2036,N_1572,N_1478);
and U2037 (N_2037,N_1412,N_1127);
nor U2038 (N_2038,N_1764,N_1346);
and U2039 (N_2039,N_1097,N_1319);
nor U2040 (N_2040,N_1260,N_1820);
nand U2041 (N_2041,N_1813,N_1762);
nand U2042 (N_2042,N_1535,N_1016);
or U2043 (N_2043,N_1592,N_1169);
nor U2044 (N_2044,N_1528,N_1510);
or U2045 (N_2045,N_1167,N_1385);
xnor U2046 (N_2046,N_1315,N_1886);
and U2047 (N_2047,N_1095,N_1779);
nor U2048 (N_2048,N_1695,N_1828);
nand U2049 (N_2049,N_1609,N_1013);
and U2050 (N_2050,N_1742,N_1663);
or U2051 (N_2051,N_1046,N_1445);
xor U2052 (N_2052,N_1636,N_1292);
nor U2053 (N_2053,N_1059,N_1207);
nand U2054 (N_2054,N_1946,N_1226);
and U2055 (N_2055,N_1321,N_1556);
nand U2056 (N_2056,N_1558,N_1085);
nand U2057 (N_2057,N_1578,N_1249);
nand U2058 (N_2058,N_1938,N_1765);
nor U2059 (N_2059,N_1736,N_1330);
nand U2060 (N_2060,N_1618,N_1550);
or U2061 (N_2061,N_1158,N_1376);
nand U2062 (N_2062,N_1287,N_1690);
and U2063 (N_2063,N_1621,N_1061);
and U2064 (N_2064,N_1964,N_1810);
nor U2065 (N_2065,N_1274,N_1721);
and U2066 (N_2066,N_1162,N_1317);
and U2067 (N_2067,N_1596,N_1824);
nand U2068 (N_2068,N_1519,N_1116);
and U2069 (N_2069,N_1474,N_1587);
nand U2070 (N_2070,N_1924,N_1190);
and U2071 (N_2071,N_1969,N_1030);
xnor U2072 (N_2072,N_1897,N_1832);
xnor U2073 (N_2073,N_1922,N_1804);
nand U2074 (N_2074,N_1763,N_1067);
nand U2075 (N_2075,N_1144,N_1204);
nor U2076 (N_2076,N_1774,N_1790);
nor U2077 (N_2077,N_1554,N_1232);
nand U2078 (N_2078,N_1381,N_1271);
and U2079 (N_2079,N_1383,N_1872);
nor U2080 (N_2080,N_1679,N_1137);
and U2081 (N_2081,N_1340,N_1212);
or U2082 (N_2082,N_1266,N_1312);
and U2083 (N_2083,N_1814,N_1120);
nand U2084 (N_2084,N_1858,N_1084);
nand U2085 (N_2085,N_1267,N_1595);
xor U2086 (N_2086,N_1342,N_1576);
and U2087 (N_2087,N_1058,N_1318);
and U2088 (N_2088,N_1219,N_1983);
xor U2089 (N_2089,N_1700,N_1781);
or U2090 (N_2090,N_1976,N_1564);
nor U2091 (N_2091,N_1605,N_1791);
nand U2092 (N_2092,N_1211,N_1094);
xnor U2093 (N_2093,N_1082,N_1996);
or U2094 (N_2094,N_1074,N_1654);
or U2095 (N_2095,N_1105,N_1138);
or U2096 (N_2096,N_1582,N_1155);
or U2097 (N_2097,N_1165,N_1063);
nand U2098 (N_2098,N_1987,N_1834);
nor U2099 (N_2099,N_1205,N_1688);
nand U2100 (N_2100,N_1959,N_1917);
and U2101 (N_2101,N_1153,N_1460);
and U2102 (N_2102,N_1320,N_1745);
xnor U2103 (N_2103,N_1770,N_1766);
nand U2104 (N_2104,N_1939,N_1694);
nor U2105 (N_2105,N_1594,N_1571);
xnor U2106 (N_2106,N_1607,N_1150);
nor U2107 (N_2107,N_1610,N_1102);
nor U2108 (N_2108,N_1379,N_1769);
nand U2109 (N_2109,N_1422,N_1933);
nand U2110 (N_2110,N_1705,N_1324);
or U2111 (N_2111,N_1850,N_1086);
and U2112 (N_2112,N_1998,N_1454);
xnor U2113 (N_2113,N_1163,N_1544);
and U2114 (N_2114,N_1551,N_1634);
nand U2115 (N_2115,N_1425,N_1493);
or U2116 (N_2116,N_1489,N_1348);
or U2117 (N_2117,N_1555,N_1613);
nor U2118 (N_2118,N_1809,N_1434);
or U2119 (N_2119,N_1691,N_1432);
nand U2120 (N_2120,N_1275,N_1685);
nor U2121 (N_2121,N_1078,N_1899);
nor U2122 (N_2122,N_1988,N_1991);
nor U2123 (N_2123,N_1088,N_1044);
or U2124 (N_2124,N_1981,N_1377);
xor U2125 (N_2125,N_1026,N_1704);
or U2126 (N_2126,N_1638,N_1986);
or U2127 (N_2127,N_1538,N_1608);
nor U2128 (N_2128,N_1483,N_1438);
or U2129 (N_2129,N_1282,N_1540);
nand U2130 (N_2130,N_1869,N_1221);
or U2131 (N_2131,N_1053,N_1786);
and U2132 (N_2132,N_1787,N_1815);
nor U2133 (N_2133,N_1301,N_1802);
xnor U2134 (N_2134,N_1229,N_1714);
nor U2135 (N_2135,N_1602,N_1258);
or U2136 (N_2136,N_1270,N_1149);
nor U2137 (N_2137,N_1943,N_1754);
xnor U2138 (N_2138,N_1753,N_1356);
and U2139 (N_2139,N_1593,N_1011);
nand U2140 (N_2140,N_1142,N_1389);
and U2141 (N_2141,N_1336,N_1390);
xor U2142 (N_2142,N_1928,N_1300);
nor U2143 (N_2143,N_1416,N_1072);
nand U2144 (N_2144,N_1083,N_1701);
nand U2145 (N_2145,N_1123,N_1503);
and U2146 (N_2146,N_1130,N_1748);
or U2147 (N_2147,N_1308,N_1374);
or U2148 (N_2148,N_1811,N_1896);
and U2149 (N_2149,N_1890,N_1606);
and U2150 (N_2150,N_1857,N_1294);
nor U2151 (N_2151,N_1451,N_1885);
and U2152 (N_2152,N_1744,N_1513);
nand U2153 (N_2153,N_1974,N_1712);
nand U2154 (N_2154,N_1189,N_1901);
or U2155 (N_2155,N_1498,N_1341);
nor U2156 (N_2156,N_1990,N_1773);
nor U2157 (N_2157,N_1399,N_1029);
xnor U2158 (N_2158,N_1673,N_1338);
nand U2159 (N_2159,N_1414,N_1043);
nor U2160 (N_2160,N_1584,N_1491);
and U2161 (N_2161,N_1629,N_1883);
and U2162 (N_2162,N_1831,N_1994);
or U2163 (N_2163,N_1724,N_1524);
nand U2164 (N_2164,N_1539,N_1224);
or U2165 (N_2165,N_1984,N_1291);
nor U2166 (N_2166,N_1512,N_1898);
nor U2167 (N_2167,N_1351,N_1104);
nand U2168 (N_2168,N_1716,N_1041);
and U2169 (N_2169,N_1435,N_1670);
or U2170 (N_2170,N_1180,N_1141);
nand U2171 (N_2171,N_1014,N_1655);
and U2172 (N_2172,N_1119,N_1822);
xnor U2173 (N_2173,N_1598,N_1424);
nand U2174 (N_2174,N_1240,N_1192);
xor U2175 (N_2175,N_1749,N_1601);
nand U2176 (N_2176,N_1126,N_1365);
nor U2177 (N_2177,N_1426,N_1682);
and U2178 (N_2178,N_1361,N_1923);
or U2179 (N_2179,N_1680,N_1747);
and U2180 (N_2180,N_1428,N_1148);
xor U2181 (N_2181,N_1891,N_1045);
and U2182 (N_2182,N_1664,N_1406);
and U2183 (N_2183,N_1278,N_1100);
and U2184 (N_2184,N_1040,N_1635);
nand U2185 (N_2185,N_1620,N_1625);
nand U2186 (N_2186,N_1382,N_1047);
nand U2187 (N_2187,N_1281,N_1561);
and U2188 (N_2188,N_1837,N_1722);
nor U2189 (N_2189,N_1051,N_1835);
and U2190 (N_2190,N_1942,N_1725);
or U2191 (N_2191,N_1372,N_1841);
nor U2192 (N_2192,N_1929,N_1633);
nor U2193 (N_2193,N_1265,N_1952);
and U2194 (N_2194,N_1882,N_1332);
nand U2195 (N_2195,N_1209,N_1256);
or U2196 (N_2196,N_1298,N_1657);
nor U2197 (N_2197,N_1954,N_1089);
and U2198 (N_2198,N_1639,N_1971);
and U2199 (N_2199,N_1836,N_1980);
and U2200 (N_2200,N_1549,N_1027);
nor U2201 (N_2201,N_1056,N_1198);
and U2202 (N_2202,N_1168,N_1808);
nand U2203 (N_2203,N_1829,N_1526);
nand U2204 (N_2204,N_1533,N_1234);
or U2205 (N_2205,N_1050,N_1182);
or U2206 (N_2206,N_1711,N_1874);
nor U2207 (N_2207,N_1036,N_1652);
or U2208 (N_2208,N_1909,N_1855);
nor U2209 (N_2209,N_1368,N_1669);
nor U2210 (N_2210,N_1840,N_1798);
or U2211 (N_2211,N_1586,N_1285);
nand U2212 (N_2212,N_1293,N_1847);
or U2213 (N_2213,N_1737,N_1877);
or U2214 (N_2214,N_1499,N_1830);
nor U2215 (N_2215,N_1279,N_1230);
and U2216 (N_2216,N_1257,N_1778);
and U2217 (N_2217,N_1464,N_1490);
or U2218 (N_2218,N_1968,N_1131);
and U2219 (N_2219,N_1443,N_1839);
nor U2220 (N_2220,N_1075,N_1589);
or U2221 (N_2221,N_1989,N_1201);
nor U2222 (N_2222,N_1235,N_1552);
nand U2223 (N_2223,N_1070,N_1719);
nand U2224 (N_2224,N_1247,N_1878);
nor U2225 (N_2225,N_1220,N_1865);
nor U2226 (N_2226,N_1852,N_1283);
nand U2227 (N_2227,N_1910,N_1517);
or U2228 (N_2228,N_1170,N_1420);
nand U2229 (N_2229,N_1966,N_1920);
or U2230 (N_2230,N_1628,N_1945);
and U2231 (N_2231,N_1449,N_1296);
nand U2232 (N_2232,N_1448,N_1112);
and U2233 (N_2233,N_1683,N_1427);
or U2234 (N_2234,N_1617,N_1767);
and U2235 (N_2235,N_1181,N_1873);
and U2236 (N_2236,N_1161,N_1881);
nand U2237 (N_2237,N_1091,N_1914);
nor U2238 (N_2238,N_1644,N_1054);
and U2239 (N_2239,N_1641,N_1780);
and U2240 (N_2240,N_1818,N_1530);
and U2241 (N_2241,N_1861,N_1151);
nand U2242 (N_2242,N_1471,N_1073);
and U2243 (N_2243,N_1122,N_1080);
and U2244 (N_2244,N_1823,N_1941);
nand U2245 (N_2245,N_1115,N_1031);
nand U2246 (N_2246,N_1065,N_1132);
nand U2247 (N_2247,N_1674,N_1286);
nor U2248 (N_2248,N_1647,N_1194);
nand U2249 (N_2249,N_1160,N_1183);
and U2250 (N_2250,N_1485,N_1912);
nor U2251 (N_2251,N_1525,N_1066);
nand U2252 (N_2252,N_1500,N_1532);
nand U2253 (N_2253,N_1482,N_1433);
or U2254 (N_2254,N_1911,N_1410);
and U2255 (N_2255,N_1166,N_1955);
nand U2256 (N_2256,N_1559,N_1187);
nand U2257 (N_2257,N_1807,N_1106);
or U2258 (N_2258,N_1060,N_1430);
and U2259 (N_2259,N_1775,N_1128);
and U2260 (N_2260,N_1472,N_1009);
or U2261 (N_2261,N_1186,N_1147);
nor U2262 (N_2262,N_1591,N_1951);
nand U2263 (N_2263,N_1337,N_1827);
nor U2264 (N_2264,N_1603,N_1854);
nor U2265 (N_2265,N_1845,N_1007);
nor U2266 (N_2266,N_1251,N_1751);
or U2267 (N_2267,N_1903,N_1311);
nand U2268 (N_2268,N_1686,N_1470);
or U2269 (N_2269,N_1562,N_1304);
or U2270 (N_2270,N_1507,N_1739);
and U2271 (N_2271,N_1653,N_1269);
nor U2272 (N_2272,N_1501,N_1473);
nand U2273 (N_2273,N_1323,N_1805);
or U2274 (N_2274,N_1488,N_1868);
xnor U2275 (N_2275,N_1494,N_1081);
xnor U2276 (N_2276,N_1684,N_1667);
or U2277 (N_2277,N_1396,N_1876);
xnor U2278 (N_2278,N_1255,N_1042);
xnor U2279 (N_2279,N_1543,N_1071);
nand U2280 (N_2280,N_1803,N_1113);
and U2281 (N_2281,N_1092,N_1157);
nand U2282 (N_2282,N_1978,N_1817);
or U2283 (N_2283,N_1570,N_1110);
nand U2284 (N_2284,N_1429,N_1010);
nand U2285 (N_2285,N_1152,N_1146);
nor U2286 (N_2286,N_1580,N_1391);
xor U2287 (N_2287,N_1394,N_1948);
nand U2288 (N_2288,N_1892,N_1843);
and U2289 (N_2289,N_1431,N_1581);
nor U2290 (N_2290,N_1545,N_1757);
nand U2291 (N_2291,N_1447,N_1992);
and U2292 (N_2292,N_1273,N_1314);
and U2293 (N_2293,N_1560,N_1768);
nor U2294 (N_2294,N_1076,N_1611);
nand U2295 (N_2295,N_1590,N_1355);
or U2296 (N_2296,N_1098,N_1760);
or U2297 (N_2297,N_1569,N_1838);
nand U2298 (N_2298,N_1970,N_1349);
xnor U2299 (N_2299,N_1867,N_1801);
nand U2300 (N_2300,N_1949,N_1495);
and U2301 (N_2301,N_1585,N_1184);
and U2302 (N_2302,N_1048,N_1261);
nor U2303 (N_2303,N_1916,N_1965);
or U2304 (N_2304,N_1859,N_1797);
or U2305 (N_2305,N_1436,N_1795);
and U2306 (N_2306,N_1668,N_1537);
and U2307 (N_2307,N_1164,N_1661);
nor U2308 (N_2308,N_1677,N_1627);
nor U2309 (N_2309,N_1440,N_1437);
and U2310 (N_2310,N_1846,N_1962);
nor U2311 (N_2311,N_1276,N_1637);
or U2312 (N_2312,N_1772,N_1729);
nand U2313 (N_2313,N_1514,N_1109);
nor U2314 (N_2314,N_1913,N_1640);
nand U2315 (N_2315,N_1518,N_1821);
nand U2316 (N_2316,N_1334,N_1310);
nor U2317 (N_2317,N_1371,N_1782);
or U2318 (N_2318,N_1021,N_1333);
nor U2319 (N_2319,N_1107,N_1386);
xor U2320 (N_2320,N_1401,N_1210);
and U2321 (N_2321,N_1237,N_1958);
and U2322 (N_2322,N_1723,N_1233);
nor U2323 (N_2323,N_1935,N_1708);
nor U2324 (N_2324,N_1395,N_1566);
nor U2325 (N_2325,N_1111,N_1173);
nor U2326 (N_2326,N_1521,N_1776);
or U2327 (N_2327,N_1019,N_1696);
or U2328 (N_2328,N_1002,N_1573);
and U2329 (N_2329,N_1335,N_1236);
nor U2330 (N_2330,N_1364,N_1614);
nand U2331 (N_2331,N_1402,N_1504);
and U2332 (N_2332,N_1523,N_1651);
nor U2333 (N_2333,N_1322,N_1692);
or U2334 (N_2334,N_1761,N_1936);
nor U2335 (N_2335,N_1370,N_1049);
and U2336 (N_2336,N_1703,N_1666);
or U2337 (N_2337,N_1387,N_1441);
nor U2338 (N_2338,N_1248,N_1185);
nand U2339 (N_2339,N_1175,N_1497);
and U2340 (N_2340,N_1527,N_1302);
and U2341 (N_2341,N_1400,N_1746);
or U2342 (N_2342,N_1902,N_1579);
or U2343 (N_2343,N_1238,N_1623);
nand U2344 (N_2344,N_1015,N_1702);
nor U2345 (N_2345,N_1289,N_1693);
nand U2346 (N_2346,N_1612,N_1024);
nor U2347 (N_2347,N_1630,N_1888);
or U2348 (N_2348,N_1875,N_1417);
nor U2349 (N_2349,N_1531,N_1656);
nand U2350 (N_2350,N_1461,N_1297);
nand U2351 (N_2351,N_1905,N_1496);
nor U2352 (N_2352,N_1956,N_1957);
or U2353 (N_2353,N_1218,N_1930);
and U2354 (N_2354,N_1177,N_1353);
nand U2355 (N_2355,N_1678,N_1502);
xor U2356 (N_2356,N_1622,N_1893);
nor U2357 (N_2357,N_1812,N_1343);
and U2358 (N_2358,N_1135,N_1154);
nor U2359 (N_2359,N_1960,N_1731);
nor U2360 (N_2360,N_1367,N_1407);
and U2361 (N_2361,N_1032,N_1193);
nand U2362 (N_2362,N_1973,N_1643);
nand U2363 (N_2363,N_1200,N_1423);
and U2364 (N_2364,N_1262,N_1462);
and U2365 (N_2365,N_1931,N_1467);
nand U2366 (N_2366,N_1479,N_1028);
and U2367 (N_2367,N_1900,N_1726);
and U2368 (N_2368,N_1730,N_1378);
nand U2369 (N_2369,N_1870,N_1415);
and U2370 (N_2370,N_1191,N_1624);
nand U2371 (N_2371,N_1362,N_1179);
nand U2372 (N_2372,N_1124,N_1213);
or U2373 (N_2373,N_1477,N_1125);
nor U2374 (N_2374,N_1534,N_1536);
nand U2375 (N_2375,N_1649,N_1894);
nor U2376 (N_2376,N_1411,N_1079);
and U2377 (N_2377,N_1565,N_1906);
nand U2378 (N_2378,N_1963,N_1844);
nand U2379 (N_2379,N_1825,N_1216);
nor U2380 (N_2380,N_1068,N_1631);
nor U2381 (N_2381,N_1129,N_1508);
or U2382 (N_2382,N_1171,N_1143);
and U2383 (N_2383,N_1806,N_1419);
and U2384 (N_2384,N_1979,N_1866);
and U2385 (N_2385,N_1784,N_1468);
or U2386 (N_2386,N_1604,N_1174);
xnor U2387 (N_2387,N_1196,N_1214);
or U2388 (N_2388,N_1064,N_1972);
and U2389 (N_2389,N_1208,N_1567);
nand U2390 (N_2390,N_1290,N_1642);
xor U2391 (N_2391,N_1457,N_1453);
nand U2392 (N_2392,N_1718,N_1759);
and U2393 (N_2393,N_1715,N_1093);
xor U2394 (N_2394,N_1363,N_1658);
or U2395 (N_2395,N_1789,N_1734);
and U2396 (N_2396,N_1139,N_1038);
nor U2397 (N_2397,N_1574,N_1675);
or U2398 (N_2398,N_1506,N_1853);
and U2399 (N_2399,N_1800,N_1915);
or U2400 (N_2400,N_1259,N_1993);
and U2401 (N_2401,N_1699,N_1246);
xnor U2402 (N_2402,N_1887,N_1062);
nand U2403 (N_2403,N_1090,N_1020);
nand U2404 (N_2404,N_1339,N_1583);
nand U2405 (N_2405,N_1710,N_1199);
and U2406 (N_2406,N_1985,N_1012);
nand U2407 (N_2407,N_1392,N_1819);
nor U2408 (N_2408,N_1557,N_1360);
and U2409 (N_2409,N_1871,N_1487);
and U2410 (N_2410,N_1309,N_1316);
nand U2411 (N_2411,N_1313,N_1404);
and U2412 (N_2412,N_1466,N_1619);
or U2413 (N_2413,N_1953,N_1785);
nand U2414 (N_2414,N_1927,N_1961);
or U2415 (N_2415,N_1727,N_1421);
nor U2416 (N_2416,N_1717,N_1553);
and U2417 (N_2417,N_1178,N_1000);
nand U2418 (N_2418,N_1103,N_1967);
and U2419 (N_2419,N_1206,N_1597);
xnor U2420 (N_2420,N_1568,N_1136);
or U2421 (N_2421,N_1475,N_1741);
or U2422 (N_2422,N_1001,N_1999);
xnor U2423 (N_2423,N_1344,N_1783);
or U2424 (N_2424,N_1484,N_1195);
xor U2425 (N_2425,N_1541,N_1121);
and U2426 (N_2426,N_1904,N_1950);
and U2427 (N_2427,N_1215,N_1203);
nor U2428 (N_2428,N_1017,N_1733);
or U2429 (N_2429,N_1720,N_1862);
or U2430 (N_2430,N_1231,N_1118);
xnor U2431 (N_2431,N_1743,N_1280);
or U2432 (N_2432,N_1481,N_1035);
nor U2433 (N_2433,N_1697,N_1239);
nor U2434 (N_2434,N_1975,N_1277);
nand U2435 (N_2435,N_1616,N_1176);
nand U2436 (N_2436,N_1398,N_1706);
nor U2437 (N_2437,N_1908,N_1563);
nand U2438 (N_2438,N_1546,N_1188);
and U2439 (N_2439,N_1826,N_1241);
or U2440 (N_2440,N_1707,N_1306);
nand U2441 (N_2441,N_1439,N_1303);
and U2442 (N_2442,N_1511,N_1735);
nor U2443 (N_2443,N_1851,N_1626);
or U2444 (N_2444,N_1096,N_1895);
or U2445 (N_2445,N_1884,N_1632);
nor U2446 (N_2446,N_1879,N_1057);
nand U2447 (N_2447,N_1465,N_1752);
nand U2448 (N_2448,N_1944,N_1295);
nor U2449 (N_2449,N_1418,N_1687);
or U2450 (N_2450,N_1345,N_1101);
and U2451 (N_2451,N_1516,N_1548);
xnor U2452 (N_2452,N_1393,N_1227);
or U2453 (N_2453,N_1671,N_1444);
or U2454 (N_2454,N_1272,N_1172);
nand U2455 (N_2455,N_1034,N_1476);
nor U2456 (N_2456,N_1455,N_1756);
xor U2457 (N_2457,N_1794,N_1842);
xnor U2458 (N_2458,N_1520,N_1515);
nor U2459 (N_2459,N_1052,N_1242);
and U2460 (N_2460,N_1645,N_1750);
nor U2461 (N_2461,N_1264,N_1329);
or U2462 (N_2462,N_1698,N_1650);
nand U2463 (N_2463,N_1388,N_1055);
nand U2464 (N_2464,N_1672,N_1023);
nand U2465 (N_2465,N_1522,N_1713);
and U2466 (N_2466,N_1225,N_1997);
nor U2467 (N_2467,N_1022,N_1039);
xor U2468 (N_2468,N_1796,N_1646);
xnor U2469 (N_2469,N_1732,N_1505);
or U2470 (N_2470,N_1660,N_1486);
or U2471 (N_2471,N_1588,N_1108);
xor U2472 (N_2472,N_1134,N_1354);
and U2473 (N_2473,N_1003,N_1771);
nand U2474 (N_2474,N_1880,N_1648);
and U2475 (N_2475,N_1077,N_1547);
nor U2476 (N_2476,N_1133,N_1755);
or U2477 (N_2477,N_1033,N_1925);
or U2478 (N_2478,N_1117,N_1403);
and U2479 (N_2479,N_1253,N_1738);
nand U2480 (N_2480,N_1250,N_1254);
nand U2481 (N_2481,N_1889,N_1025);
and U2482 (N_2482,N_1375,N_1327);
nand U2483 (N_2483,N_1934,N_1305);
and U2484 (N_2484,N_1006,N_1799);
and U2485 (N_2485,N_1326,N_1469);
nand U2486 (N_2486,N_1450,N_1263);
xor U2487 (N_2487,N_1350,N_1480);
or U2488 (N_2488,N_1145,N_1156);
nand U2489 (N_2489,N_1197,N_1615);
and U2490 (N_2490,N_1740,N_1405);
and U2491 (N_2491,N_1369,N_1373);
and U2492 (N_2492,N_1357,N_1793);
nand U2493 (N_2493,N_1325,N_1408);
nor U2494 (N_2494,N_1222,N_1005);
xor U2495 (N_2495,N_1940,N_1245);
nor U2496 (N_2496,N_1358,N_1244);
and U2497 (N_2497,N_1446,N_1599);
nor U2498 (N_2498,N_1228,N_1018);
or U2499 (N_2499,N_1413,N_1114);
nand U2500 (N_2500,N_1992,N_1504);
and U2501 (N_2501,N_1079,N_1703);
nor U2502 (N_2502,N_1941,N_1912);
nor U2503 (N_2503,N_1305,N_1494);
and U2504 (N_2504,N_1198,N_1197);
nand U2505 (N_2505,N_1692,N_1430);
nor U2506 (N_2506,N_1045,N_1994);
nand U2507 (N_2507,N_1350,N_1354);
nand U2508 (N_2508,N_1014,N_1560);
or U2509 (N_2509,N_1927,N_1192);
and U2510 (N_2510,N_1051,N_1674);
or U2511 (N_2511,N_1795,N_1642);
and U2512 (N_2512,N_1353,N_1449);
or U2513 (N_2513,N_1789,N_1134);
xor U2514 (N_2514,N_1562,N_1865);
nor U2515 (N_2515,N_1964,N_1819);
or U2516 (N_2516,N_1877,N_1308);
or U2517 (N_2517,N_1954,N_1538);
xnor U2518 (N_2518,N_1622,N_1440);
xnor U2519 (N_2519,N_1502,N_1901);
nand U2520 (N_2520,N_1736,N_1556);
xor U2521 (N_2521,N_1084,N_1412);
and U2522 (N_2522,N_1448,N_1473);
and U2523 (N_2523,N_1297,N_1626);
or U2524 (N_2524,N_1229,N_1653);
nor U2525 (N_2525,N_1127,N_1051);
and U2526 (N_2526,N_1047,N_1022);
or U2527 (N_2527,N_1274,N_1244);
and U2528 (N_2528,N_1635,N_1688);
or U2529 (N_2529,N_1141,N_1647);
nor U2530 (N_2530,N_1283,N_1289);
and U2531 (N_2531,N_1438,N_1619);
or U2532 (N_2532,N_1682,N_1120);
nor U2533 (N_2533,N_1059,N_1045);
and U2534 (N_2534,N_1269,N_1043);
or U2535 (N_2535,N_1294,N_1874);
or U2536 (N_2536,N_1867,N_1814);
nand U2537 (N_2537,N_1902,N_1502);
and U2538 (N_2538,N_1508,N_1551);
nand U2539 (N_2539,N_1454,N_1330);
nand U2540 (N_2540,N_1816,N_1498);
nand U2541 (N_2541,N_1490,N_1129);
or U2542 (N_2542,N_1388,N_1294);
and U2543 (N_2543,N_1135,N_1293);
and U2544 (N_2544,N_1701,N_1879);
xnor U2545 (N_2545,N_1450,N_1119);
or U2546 (N_2546,N_1959,N_1431);
nor U2547 (N_2547,N_1704,N_1440);
and U2548 (N_2548,N_1726,N_1636);
and U2549 (N_2549,N_1374,N_1392);
or U2550 (N_2550,N_1394,N_1715);
nand U2551 (N_2551,N_1029,N_1219);
nand U2552 (N_2552,N_1589,N_1110);
xnor U2553 (N_2553,N_1973,N_1971);
nor U2554 (N_2554,N_1111,N_1049);
xnor U2555 (N_2555,N_1428,N_1967);
and U2556 (N_2556,N_1055,N_1737);
or U2557 (N_2557,N_1483,N_1761);
nor U2558 (N_2558,N_1745,N_1915);
nor U2559 (N_2559,N_1647,N_1087);
xnor U2560 (N_2560,N_1497,N_1461);
nand U2561 (N_2561,N_1696,N_1340);
nand U2562 (N_2562,N_1059,N_1859);
nand U2563 (N_2563,N_1819,N_1722);
or U2564 (N_2564,N_1352,N_1819);
and U2565 (N_2565,N_1127,N_1433);
and U2566 (N_2566,N_1702,N_1327);
or U2567 (N_2567,N_1768,N_1697);
nand U2568 (N_2568,N_1954,N_1384);
and U2569 (N_2569,N_1030,N_1207);
nand U2570 (N_2570,N_1675,N_1882);
and U2571 (N_2571,N_1983,N_1240);
or U2572 (N_2572,N_1316,N_1763);
nand U2573 (N_2573,N_1859,N_1836);
nor U2574 (N_2574,N_1688,N_1724);
nand U2575 (N_2575,N_1719,N_1649);
nand U2576 (N_2576,N_1130,N_1549);
or U2577 (N_2577,N_1123,N_1397);
nor U2578 (N_2578,N_1498,N_1881);
nor U2579 (N_2579,N_1016,N_1145);
nand U2580 (N_2580,N_1833,N_1098);
and U2581 (N_2581,N_1881,N_1680);
nor U2582 (N_2582,N_1316,N_1829);
nand U2583 (N_2583,N_1309,N_1823);
nor U2584 (N_2584,N_1511,N_1829);
and U2585 (N_2585,N_1631,N_1441);
nand U2586 (N_2586,N_1543,N_1941);
nand U2587 (N_2587,N_1850,N_1835);
and U2588 (N_2588,N_1468,N_1596);
nor U2589 (N_2589,N_1606,N_1066);
or U2590 (N_2590,N_1555,N_1015);
nand U2591 (N_2591,N_1506,N_1054);
nand U2592 (N_2592,N_1580,N_1636);
nand U2593 (N_2593,N_1911,N_1247);
xor U2594 (N_2594,N_1014,N_1527);
or U2595 (N_2595,N_1670,N_1681);
and U2596 (N_2596,N_1394,N_1974);
and U2597 (N_2597,N_1333,N_1773);
and U2598 (N_2598,N_1358,N_1004);
xor U2599 (N_2599,N_1130,N_1311);
and U2600 (N_2600,N_1933,N_1996);
nor U2601 (N_2601,N_1320,N_1267);
or U2602 (N_2602,N_1752,N_1548);
nor U2603 (N_2603,N_1343,N_1685);
xnor U2604 (N_2604,N_1948,N_1479);
nand U2605 (N_2605,N_1978,N_1332);
nand U2606 (N_2606,N_1543,N_1948);
and U2607 (N_2607,N_1308,N_1230);
xor U2608 (N_2608,N_1976,N_1377);
nand U2609 (N_2609,N_1236,N_1655);
xor U2610 (N_2610,N_1480,N_1081);
and U2611 (N_2611,N_1915,N_1809);
nand U2612 (N_2612,N_1356,N_1846);
or U2613 (N_2613,N_1940,N_1126);
or U2614 (N_2614,N_1582,N_1656);
xnor U2615 (N_2615,N_1191,N_1252);
and U2616 (N_2616,N_1955,N_1518);
nand U2617 (N_2617,N_1217,N_1059);
and U2618 (N_2618,N_1094,N_1478);
nor U2619 (N_2619,N_1575,N_1336);
or U2620 (N_2620,N_1449,N_1696);
xor U2621 (N_2621,N_1330,N_1421);
nand U2622 (N_2622,N_1310,N_1134);
nor U2623 (N_2623,N_1480,N_1623);
nand U2624 (N_2624,N_1968,N_1698);
nor U2625 (N_2625,N_1590,N_1225);
nor U2626 (N_2626,N_1474,N_1202);
and U2627 (N_2627,N_1403,N_1605);
nand U2628 (N_2628,N_1171,N_1830);
nand U2629 (N_2629,N_1863,N_1123);
nor U2630 (N_2630,N_1117,N_1916);
and U2631 (N_2631,N_1579,N_1089);
and U2632 (N_2632,N_1778,N_1091);
or U2633 (N_2633,N_1827,N_1450);
and U2634 (N_2634,N_1114,N_1536);
and U2635 (N_2635,N_1873,N_1623);
nand U2636 (N_2636,N_1458,N_1569);
and U2637 (N_2637,N_1404,N_1720);
and U2638 (N_2638,N_1206,N_1820);
and U2639 (N_2639,N_1588,N_1901);
and U2640 (N_2640,N_1809,N_1485);
nor U2641 (N_2641,N_1122,N_1107);
xnor U2642 (N_2642,N_1298,N_1121);
and U2643 (N_2643,N_1689,N_1099);
or U2644 (N_2644,N_1460,N_1158);
xor U2645 (N_2645,N_1389,N_1769);
or U2646 (N_2646,N_1509,N_1304);
nor U2647 (N_2647,N_1875,N_1470);
nor U2648 (N_2648,N_1405,N_1901);
or U2649 (N_2649,N_1738,N_1316);
nor U2650 (N_2650,N_1960,N_1494);
nand U2651 (N_2651,N_1747,N_1587);
nand U2652 (N_2652,N_1892,N_1418);
nand U2653 (N_2653,N_1442,N_1817);
or U2654 (N_2654,N_1818,N_1431);
and U2655 (N_2655,N_1234,N_1144);
xor U2656 (N_2656,N_1393,N_1488);
or U2657 (N_2657,N_1752,N_1275);
nand U2658 (N_2658,N_1812,N_1635);
and U2659 (N_2659,N_1860,N_1704);
nand U2660 (N_2660,N_1718,N_1819);
and U2661 (N_2661,N_1951,N_1169);
or U2662 (N_2662,N_1727,N_1013);
or U2663 (N_2663,N_1297,N_1024);
and U2664 (N_2664,N_1203,N_1207);
xnor U2665 (N_2665,N_1279,N_1210);
nand U2666 (N_2666,N_1300,N_1988);
nand U2667 (N_2667,N_1723,N_1833);
nand U2668 (N_2668,N_1689,N_1973);
xor U2669 (N_2669,N_1869,N_1551);
and U2670 (N_2670,N_1486,N_1760);
xor U2671 (N_2671,N_1955,N_1974);
xor U2672 (N_2672,N_1795,N_1421);
nor U2673 (N_2673,N_1113,N_1770);
nand U2674 (N_2674,N_1787,N_1990);
nor U2675 (N_2675,N_1043,N_1737);
nand U2676 (N_2676,N_1354,N_1414);
xor U2677 (N_2677,N_1184,N_1152);
or U2678 (N_2678,N_1174,N_1593);
xor U2679 (N_2679,N_1287,N_1976);
and U2680 (N_2680,N_1754,N_1653);
xor U2681 (N_2681,N_1702,N_1594);
or U2682 (N_2682,N_1792,N_1282);
nor U2683 (N_2683,N_1667,N_1047);
xor U2684 (N_2684,N_1039,N_1104);
or U2685 (N_2685,N_1220,N_1177);
and U2686 (N_2686,N_1892,N_1917);
or U2687 (N_2687,N_1651,N_1302);
nor U2688 (N_2688,N_1855,N_1717);
or U2689 (N_2689,N_1727,N_1172);
or U2690 (N_2690,N_1139,N_1180);
or U2691 (N_2691,N_1921,N_1047);
xnor U2692 (N_2692,N_1100,N_1191);
nand U2693 (N_2693,N_1832,N_1912);
nor U2694 (N_2694,N_1743,N_1573);
nand U2695 (N_2695,N_1547,N_1240);
xnor U2696 (N_2696,N_1793,N_1582);
nand U2697 (N_2697,N_1388,N_1886);
or U2698 (N_2698,N_1307,N_1899);
nor U2699 (N_2699,N_1591,N_1007);
nand U2700 (N_2700,N_1157,N_1693);
and U2701 (N_2701,N_1535,N_1035);
nand U2702 (N_2702,N_1769,N_1175);
xnor U2703 (N_2703,N_1998,N_1109);
or U2704 (N_2704,N_1125,N_1518);
and U2705 (N_2705,N_1668,N_1042);
or U2706 (N_2706,N_1380,N_1604);
or U2707 (N_2707,N_1833,N_1257);
nand U2708 (N_2708,N_1711,N_1474);
nor U2709 (N_2709,N_1469,N_1358);
and U2710 (N_2710,N_1129,N_1955);
nor U2711 (N_2711,N_1687,N_1328);
and U2712 (N_2712,N_1228,N_1480);
nand U2713 (N_2713,N_1128,N_1295);
or U2714 (N_2714,N_1514,N_1587);
or U2715 (N_2715,N_1294,N_1948);
xnor U2716 (N_2716,N_1267,N_1714);
nand U2717 (N_2717,N_1953,N_1258);
and U2718 (N_2718,N_1826,N_1923);
nand U2719 (N_2719,N_1262,N_1898);
nor U2720 (N_2720,N_1968,N_1467);
nand U2721 (N_2721,N_1546,N_1622);
xnor U2722 (N_2722,N_1935,N_1219);
or U2723 (N_2723,N_1716,N_1198);
and U2724 (N_2724,N_1763,N_1788);
or U2725 (N_2725,N_1961,N_1893);
and U2726 (N_2726,N_1031,N_1524);
nor U2727 (N_2727,N_1986,N_1740);
nor U2728 (N_2728,N_1984,N_1258);
xnor U2729 (N_2729,N_1213,N_1918);
xnor U2730 (N_2730,N_1991,N_1812);
or U2731 (N_2731,N_1203,N_1823);
nor U2732 (N_2732,N_1765,N_1319);
nand U2733 (N_2733,N_1925,N_1721);
and U2734 (N_2734,N_1830,N_1083);
nor U2735 (N_2735,N_1209,N_1520);
or U2736 (N_2736,N_1489,N_1877);
nor U2737 (N_2737,N_1228,N_1687);
nor U2738 (N_2738,N_1017,N_1799);
and U2739 (N_2739,N_1070,N_1987);
or U2740 (N_2740,N_1689,N_1802);
and U2741 (N_2741,N_1382,N_1977);
or U2742 (N_2742,N_1617,N_1301);
and U2743 (N_2743,N_1499,N_1384);
or U2744 (N_2744,N_1591,N_1417);
and U2745 (N_2745,N_1883,N_1779);
and U2746 (N_2746,N_1123,N_1953);
and U2747 (N_2747,N_1770,N_1085);
nand U2748 (N_2748,N_1169,N_1298);
nor U2749 (N_2749,N_1460,N_1685);
and U2750 (N_2750,N_1871,N_1674);
xnor U2751 (N_2751,N_1835,N_1556);
and U2752 (N_2752,N_1303,N_1945);
xnor U2753 (N_2753,N_1866,N_1694);
xnor U2754 (N_2754,N_1469,N_1237);
xnor U2755 (N_2755,N_1456,N_1622);
or U2756 (N_2756,N_1845,N_1107);
and U2757 (N_2757,N_1747,N_1278);
nor U2758 (N_2758,N_1557,N_1159);
nor U2759 (N_2759,N_1968,N_1198);
nor U2760 (N_2760,N_1335,N_1778);
nand U2761 (N_2761,N_1149,N_1876);
or U2762 (N_2762,N_1727,N_1309);
and U2763 (N_2763,N_1405,N_1452);
xor U2764 (N_2764,N_1082,N_1234);
or U2765 (N_2765,N_1504,N_1804);
or U2766 (N_2766,N_1307,N_1247);
and U2767 (N_2767,N_1655,N_1747);
and U2768 (N_2768,N_1468,N_1884);
or U2769 (N_2769,N_1418,N_1360);
or U2770 (N_2770,N_1383,N_1966);
nor U2771 (N_2771,N_1981,N_1004);
or U2772 (N_2772,N_1884,N_1125);
and U2773 (N_2773,N_1003,N_1116);
or U2774 (N_2774,N_1700,N_1312);
or U2775 (N_2775,N_1281,N_1504);
xnor U2776 (N_2776,N_1218,N_1051);
or U2777 (N_2777,N_1772,N_1410);
xor U2778 (N_2778,N_1244,N_1618);
xnor U2779 (N_2779,N_1880,N_1840);
nor U2780 (N_2780,N_1101,N_1890);
nor U2781 (N_2781,N_1992,N_1198);
and U2782 (N_2782,N_1727,N_1058);
nand U2783 (N_2783,N_1802,N_1982);
or U2784 (N_2784,N_1729,N_1408);
and U2785 (N_2785,N_1308,N_1300);
nand U2786 (N_2786,N_1029,N_1804);
nand U2787 (N_2787,N_1571,N_1645);
nand U2788 (N_2788,N_1343,N_1309);
xor U2789 (N_2789,N_1678,N_1836);
and U2790 (N_2790,N_1028,N_1932);
nor U2791 (N_2791,N_1577,N_1091);
and U2792 (N_2792,N_1757,N_1432);
nor U2793 (N_2793,N_1223,N_1915);
nand U2794 (N_2794,N_1392,N_1772);
or U2795 (N_2795,N_1824,N_1324);
nor U2796 (N_2796,N_1689,N_1662);
xor U2797 (N_2797,N_1180,N_1586);
nor U2798 (N_2798,N_1159,N_1283);
nand U2799 (N_2799,N_1027,N_1799);
nand U2800 (N_2800,N_1208,N_1981);
and U2801 (N_2801,N_1933,N_1636);
and U2802 (N_2802,N_1286,N_1425);
and U2803 (N_2803,N_1830,N_1909);
nor U2804 (N_2804,N_1343,N_1224);
nand U2805 (N_2805,N_1247,N_1871);
or U2806 (N_2806,N_1383,N_1280);
and U2807 (N_2807,N_1277,N_1410);
nor U2808 (N_2808,N_1429,N_1877);
xnor U2809 (N_2809,N_1615,N_1018);
nor U2810 (N_2810,N_1745,N_1820);
and U2811 (N_2811,N_1917,N_1333);
nor U2812 (N_2812,N_1973,N_1163);
nor U2813 (N_2813,N_1187,N_1828);
or U2814 (N_2814,N_1375,N_1215);
nor U2815 (N_2815,N_1086,N_1867);
nor U2816 (N_2816,N_1937,N_1327);
nor U2817 (N_2817,N_1102,N_1881);
nor U2818 (N_2818,N_1345,N_1446);
nand U2819 (N_2819,N_1289,N_1661);
nor U2820 (N_2820,N_1437,N_1954);
nor U2821 (N_2821,N_1475,N_1975);
nand U2822 (N_2822,N_1005,N_1387);
nor U2823 (N_2823,N_1164,N_1488);
or U2824 (N_2824,N_1184,N_1875);
or U2825 (N_2825,N_1427,N_1467);
or U2826 (N_2826,N_1243,N_1146);
or U2827 (N_2827,N_1004,N_1229);
nand U2828 (N_2828,N_1127,N_1269);
xor U2829 (N_2829,N_1206,N_1533);
nor U2830 (N_2830,N_1684,N_1880);
nand U2831 (N_2831,N_1736,N_1778);
nor U2832 (N_2832,N_1819,N_1326);
nand U2833 (N_2833,N_1069,N_1804);
nand U2834 (N_2834,N_1923,N_1758);
or U2835 (N_2835,N_1107,N_1488);
xor U2836 (N_2836,N_1506,N_1882);
and U2837 (N_2837,N_1179,N_1341);
nor U2838 (N_2838,N_1499,N_1625);
or U2839 (N_2839,N_1996,N_1836);
and U2840 (N_2840,N_1401,N_1605);
nor U2841 (N_2841,N_1412,N_1985);
and U2842 (N_2842,N_1721,N_1377);
xnor U2843 (N_2843,N_1807,N_1741);
xor U2844 (N_2844,N_1940,N_1725);
nor U2845 (N_2845,N_1596,N_1862);
nor U2846 (N_2846,N_1127,N_1235);
and U2847 (N_2847,N_1427,N_1566);
xnor U2848 (N_2848,N_1804,N_1683);
or U2849 (N_2849,N_1252,N_1023);
nor U2850 (N_2850,N_1635,N_1315);
or U2851 (N_2851,N_1907,N_1835);
nor U2852 (N_2852,N_1838,N_1885);
nor U2853 (N_2853,N_1987,N_1380);
nor U2854 (N_2854,N_1982,N_1731);
and U2855 (N_2855,N_1201,N_1589);
or U2856 (N_2856,N_1765,N_1183);
or U2857 (N_2857,N_1587,N_1233);
nor U2858 (N_2858,N_1263,N_1535);
nor U2859 (N_2859,N_1010,N_1106);
xnor U2860 (N_2860,N_1493,N_1400);
or U2861 (N_2861,N_1248,N_1698);
and U2862 (N_2862,N_1943,N_1898);
nand U2863 (N_2863,N_1129,N_1948);
nor U2864 (N_2864,N_1301,N_1156);
and U2865 (N_2865,N_1884,N_1324);
and U2866 (N_2866,N_1798,N_1964);
nand U2867 (N_2867,N_1045,N_1560);
and U2868 (N_2868,N_1414,N_1285);
or U2869 (N_2869,N_1305,N_1860);
or U2870 (N_2870,N_1845,N_1331);
nand U2871 (N_2871,N_1643,N_1706);
xor U2872 (N_2872,N_1768,N_1426);
nor U2873 (N_2873,N_1338,N_1480);
nor U2874 (N_2874,N_1976,N_1697);
nor U2875 (N_2875,N_1886,N_1366);
or U2876 (N_2876,N_1875,N_1955);
nor U2877 (N_2877,N_1010,N_1586);
nand U2878 (N_2878,N_1538,N_1273);
nor U2879 (N_2879,N_1735,N_1512);
nor U2880 (N_2880,N_1031,N_1460);
nor U2881 (N_2881,N_1541,N_1183);
nor U2882 (N_2882,N_1340,N_1937);
nor U2883 (N_2883,N_1409,N_1092);
nand U2884 (N_2884,N_1377,N_1227);
nand U2885 (N_2885,N_1731,N_1794);
and U2886 (N_2886,N_1332,N_1192);
or U2887 (N_2887,N_1203,N_1116);
xor U2888 (N_2888,N_1383,N_1614);
or U2889 (N_2889,N_1925,N_1692);
nor U2890 (N_2890,N_1702,N_1395);
or U2891 (N_2891,N_1591,N_1185);
nor U2892 (N_2892,N_1891,N_1008);
and U2893 (N_2893,N_1150,N_1589);
nand U2894 (N_2894,N_1260,N_1681);
nor U2895 (N_2895,N_1099,N_1589);
nor U2896 (N_2896,N_1780,N_1387);
xor U2897 (N_2897,N_1659,N_1262);
or U2898 (N_2898,N_1047,N_1511);
nand U2899 (N_2899,N_1449,N_1902);
or U2900 (N_2900,N_1606,N_1054);
xor U2901 (N_2901,N_1959,N_1844);
nor U2902 (N_2902,N_1272,N_1375);
and U2903 (N_2903,N_1720,N_1398);
xor U2904 (N_2904,N_1519,N_1097);
nor U2905 (N_2905,N_1479,N_1561);
xor U2906 (N_2906,N_1304,N_1967);
and U2907 (N_2907,N_1634,N_1672);
nor U2908 (N_2908,N_1311,N_1426);
nor U2909 (N_2909,N_1387,N_1680);
nor U2910 (N_2910,N_1615,N_1104);
nor U2911 (N_2911,N_1391,N_1395);
nand U2912 (N_2912,N_1505,N_1487);
nor U2913 (N_2913,N_1924,N_1456);
nand U2914 (N_2914,N_1387,N_1335);
or U2915 (N_2915,N_1444,N_1615);
and U2916 (N_2916,N_1365,N_1604);
and U2917 (N_2917,N_1221,N_1641);
nand U2918 (N_2918,N_1141,N_1019);
and U2919 (N_2919,N_1020,N_1501);
nand U2920 (N_2920,N_1120,N_1330);
nor U2921 (N_2921,N_1262,N_1446);
nor U2922 (N_2922,N_1518,N_1130);
or U2923 (N_2923,N_1064,N_1136);
or U2924 (N_2924,N_1848,N_1395);
or U2925 (N_2925,N_1168,N_1801);
and U2926 (N_2926,N_1529,N_1790);
xor U2927 (N_2927,N_1463,N_1370);
xor U2928 (N_2928,N_1472,N_1511);
and U2929 (N_2929,N_1274,N_1311);
nand U2930 (N_2930,N_1315,N_1205);
nand U2931 (N_2931,N_1484,N_1712);
or U2932 (N_2932,N_1849,N_1648);
or U2933 (N_2933,N_1391,N_1742);
nor U2934 (N_2934,N_1292,N_1478);
and U2935 (N_2935,N_1438,N_1360);
and U2936 (N_2936,N_1033,N_1945);
or U2937 (N_2937,N_1151,N_1636);
and U2938 (N_2938,N_1607,N_1455);
or U2939 (N_2939,N_1476,N_1047);
or U2940 (N_2940,N_1943,N_1604);
nor U2941 (N_2941,N_1894,N_1202);
and U2942 (N_2942,N_1666,N_1354);
or U2943 (N_2943,N_1014,N_1782);
or U2944 (N_2944,N_1289,N_1664);
and U2945 (N_2945,N_1533,N_1421);
nor U2946 (N_2946,N_1032,N_1197);
nand U2947 (N_2947,N_1561,N_1741);
nand U2948 (N_2948,N_1189,N_1707);
nor U2949 (N_2949,N_1321,N_1980);
nand U2950 (N_2950,N_1589,N_1376);
nor U2951 (N_2951,N_1586,N_1351);
nor U2952 (N_2952,N_1486,N_1416);
nand U2953 (N_2953,N_1653,N_1520);
nor U2954 (N_2954,N_1020,N_1781);
or U2955 (N_2955,N_1071,N_1962);
and U2956 (N_2956,N_1508,N_1172);
nand U2957 (N_2957,N_1930,N_1862);
and U2958 (N_2958,N_1315,N_1035);
nand U2959 (N_2959,N_1314,N_1655);
nor U2960 (N_2960,N_1589,N_1658);
or U2961 (N_2961,N_1162,N_1119);
or U2962 (N_2962,N_1099,N_1868);
or U2963 (N_2963,N_1317,N_1153);
nor U2964 (N_2964,N_1810,N_1872);
or U2965 (N_2965,N_1943,N_1581);
and U2966 (N_2966,N_1388,N_1713);
or U2967 (N_2967,N_1829,N_1307);
and U2968 (N_2968,N_1217,N_1391);
nor U2969 (N_2969,N_1065,N_1739);
nor U2970 (N_2970,N_1584,N_1660);
xor U2971 (N_2971,N_1506,N_1249);
nand U2972 (N_2972,N_1944,N_1832);
nand U2973 (N_2973,N_1738,N_1511);
or U2974 (N_2974,N_1071,N_1311);
and U2975 (N_2975,N_1462,N_1689);
nor U2976 (N_2976,N_1849,N_1836);
nand U2977 (N_2977,N_1308,N_1912);
or U2978 (N_2978,N_1340,N_1654);
nor U2979 (N_2979,N_1918,N_1569);
and U2980 (N_2980,N_1791,N_1747);
or U2981 (N_2981,N_1128,N_1068);
or U2982 (N_2982,N_1285,N_1016);
and U2983 (N_2983,N_1344,N_1420);
or U2984 (N_2984,N_1274,N_1853);
nor U2985 (N_2985,N_1523,N_1932);
or U2986 (N_2986,N_1747,N_1757);
or U2987 (N_2987,N_1057,N_1378);
and U2988 (N_2988,N_1071,N_1288);
and U2989 (N_2989,N_1915,N_1097);
xnor U2990 (N_2990,N_1019,N_1745);
nand U2991 (N_2991,N_1695,N_1425);
nor U2992 (N_2992,N_1504,N_1022);
or U2993 (N_2993,N_1512,N_1364);
nand U2994 (N_2994,N_1668,N_1018);
and U2995 (N_2995,N_1233,N_1819);
and U2996 (N_2996,N_1515,N_1271);
nand U2997 (N_2997,N_1064,N_1324);
nand U2998 (N_2998,N_1038,N_1788);
or U2999 (N_2999,N_1758,N_1771);
nor U3000 (N_3000,N_2630,N_2015);
and U3001 (N_3001,N_2969,N_2991);
nor U3002 (N_3002,N_2654,N_2536);
and U3003 (N_3003,N_2049,N_2677);
nand U3004 (N_3004,N_2873,N_2135);
nor U3005 (N_3005,N_2762,N_2201);
xnor U3006 (N_3006,N_2980,N_2611);
or U3007 (N_3007,N_2352,N_2697);
or U3008 (N_3008,N_2792,N_2406);
nand U3009 (N_3009,N_2585,N_2649);
nor U3010 (N_3010,N_2220,N_2417);
or U3011 (N_3011,N_2271,N_2750);
nand U3012 (N_3012,N_2653,N_2850);
and U3013 (N_3013,N_2771,N_2217);
nand U3014 (N_3014,N_2313,N_2885);
nand U3015 (N_3015,N_2027,N_2727);
nor U3016 (N_3016,N_2460,N_2328);
xnor U3017 (N_3017,N_2495,N_2317);
or U3018 (N_3018,N_2411,N_2517);
nor U3019 (N_3019,N_2290,N_2811);
xnor U3020 (N_3020,N_2337,N_2810);
and U3021 (N_3021,N_2799,N_2302);
or U3022 (N_3022,N_2544,N_2367);
nand U3023 (N_3023,N_2702,N_2205);
nor U3024 (N_3024,N_2211,N_2509);
and U3025 (N_3025,N_2715,N_2721);
nand U3026 (N_3026,N_2741,N_2722);
xnor U3027 (N_3027,N_2320,N_2599);
nand U3028 (N_3028,N_2005,N_2783);
or U3029 (N_3029,N_2159,N_2160);
or U3030 (N_3030,N_2202,N_2403);
and U3031 (N_3031,N_2474,N_2747);
and U3032 (N_3032,N_2760,N_2842);
nand U3033 (N_3033,N_2034,N_2666);
or U3034 (N_3034,N_2289,N_2609);
or U3035 (N_3035,N_2634,N_2689);
nor U3036 (N_3036,N_2108,N_2746);
or U3037 (N_3037,N_2351,N_2790);
and U3038 (N_3038,N_2710,N_2934);
nor U3039 (N_3039,N_2864,N_2006);
nand U3040 (N_3040,N_2208,N_2481);
and U3041 (N_3041,N_2923,N_2553);
nand U3042 (N_3042,N_2911,N_2943);
or U3043 (N_3043,N_2789,N_2977);
nand U3044 (N_3044,N_2636,N_2733);
nand U3045 (N_3045,N_2392,N_2322);
nand U3046 (N_3046,N_2619,N_2974);
nand U3047 (N_3047,N_2142,N_2079);
nand U3048 (N_3048,N_2145,N_2755);
and U3049 (N_3049,N_2307,N_2359);
or U3050 (N_3050,N_2652,N_2239);
and U3051 (N_3051,N_2028,N_2759);
xnor U3052 (N_3052,N_2554,N_2833);
or U3053 (N_3053,N_2578,N_2321);
and U3054 (N_3054,N_2989,N_2304);
nor U3055 (N_3055,N_2797,N_2502);
and U3056 (N_3056,N_2254,N_2470);
nand U3057 (N_3057,N_2880,N_2272);
or U3058 (N_3058,N_2489,N_2287);
nand U3059 (N_3059,N_2156,N_2749);
nand U3060 (N_3060,N_2099,N_2516);
or U3061 (N_3061,N_2175,N_2176);
or U3062 (N_3062,N_2354,N_2572);
xnor U3063 (N_3063,N_2106,N_2729);
nand U3064 (N_3064,N_2580,N_2889);
or U3065 (N_3065,N_2523,N_2920);
nand U3066 (N_3066,N_2828,N_2679);
or U3067 (N_3067,N_2555,N_2737);
and U3068 (N_3068,N_2266,N_2625);
nand U3069 (N_3069,N_2624,N_2957);
nand U3070 (N_3070,N_2541,N_2298);
xnor U3071 (N_3071,N_2694,N_2812);
or U3072 (N_3072,N_2404,N_2471);
xor U3073 (N_3073,N_2238,N_2023);
or U3074 (N_3074,N_2641,N_2731);
and U3075 (N_3075,N_2848,N_2025);
and U3076 (N_3076,N_2081,N_2745);
nor U3077 (N_3077,N_2425,N_2912);
or U3078 (N_3078,N_2146,N_2192);
nor U3079 (N_3079,N_2919,N_2103);
or U3080 (N_3080,N_2659,N_2177);
or U3081 (N_3081,N_2959,N_2498);
nand U3082 (N_3082,N_2942,N_2396);
nor U3083 (N_3083,N_2904,N_2844);
nand U3084 (N_3084,N_2595,N_2821);
nor U3085 (N_3085,N_2091,N_2700);
nand U3086 (N_3086,N_2087,N_2093);
nor U3087 (N_3087,N_2968,N_2798);
and U3088 (N_3088,N_2843,N_2781);
and U3089 (N_3089,N_2469,N_2874);
xor U3090 (N_3090,N_2228,N_2273);
nand U3091 (N_3091,N_2092,N_2558);
and U3092 (N_3092,N_2251,N_2350);
or U3093 (N_3093,N_2846,N_2308);
or U3094 (N_3094,N_2382,N_2455);
or U3095 (N_3095,N_2493,N_2144);
xnor U3096 (N_3096,N_2983,N_2375);
nand U3097 (N_3097,N_2956,N_2349);
nand U3098 (N_3098,N_2535,N_2708);
nand U3099 (N_3099,N_2219,N_2736);
and U3100 (N_3100,N_2610,N_2086);
nand U3101 (N_3101,N_2608,N_2181);
nor U3102 (N_3102,N_2235,N_2180);
nand U3103 (N_3103,N_2297,N_2899);
and U3104 (N_3104,N_2960,N_2420);
nand U3105 (N_3105,N_2607,N_2267);
nand U3106 (N_3106,N_2987,N_2114);
and U3107 (N_3107,N_2263,N_2627);
or U3108 (N_3108,N_2426,N_2947);
nand U3109 (N_3109,N_2701,N_2463);
nand U3110 (N_3110,N_2130,N_2838);
or U3111 (N_3111,N_2587,N_2095);
nand U3112 (N_3112,N_2647,N_2327);
nor U3113 (N_3113,N_2152,N_2340);
nand U3114 (N_3114,N_2073,N_2293);
nor U3115 (N_3115,N_2391,N_2237);
nor U3116 (N_3116,N_2836,N_2451);
nor U3117 (N_3117,N_2061,N_2914);
and U3118 (N_3118,N_2837,N_2094);
and U3119 (N_3119,N_2900,N_2633);
nand U3120 (N_3120,N_2526,N_2077);
or U3121 (N_3121,N_2941,N_2164);
nand U3122 (N_3122,N_2954,N_2256);
xor U3123 (N_3123,N_2024,N_2245);
or U3124 (N_3124,N_2815,N_2813);
or U3125 (N_3125,N_2043,N_2961);
or U3126 (N_3126,N_2300,N_2591);
nand U3127 (N_3127,N_2070,N_2170);
nand U3128 (N_3128,N_2774,N_2550);
and U3129 (N_3129,N_2962,N_2851);
nor U3130 (N_3130,N_2058,N_2318);
nand U3131 (N_3131,N_2906,N_2910);
nor U3132 (N_3132,N_2832,N_2125);
nand U3133 (N_3133,N_2068,N_2496);
xor U3134 (N_3134,N_2089,N_2944);
xnor U3135 (N_3135,N_2384,N_2705);
and U3136 (N_3136,N_2998,N_2744);
or U3137 (N_3137,N_2690,N_2497);
nand U3138 (N_3138,N_2743,N_2414);
nand U3139 (N_3139,N_2286,N_2724);
nor U3140 (N_3140,N_2664,N_2617);
and U3141 (N_3141,N_2213,N_2029);
or U3142 (N_3142,N_2676,N_2150);
or U3143 (N_3143,N_2547,N_2379);
nor U3144 (N_3144,N_2818,N_2780);
nor U3145 (N_3145,N_2827,N_2695);
or U3146 (N_3146,N_2820,N_2712);
xnor U3147 (N_3147,N_2675,N_2107);
or U3148 (N_3148,N_2126,N_2937);
or U3149 (N_3149,N_2405,N_2728);
xor U3150 (N_3150,N_2198,N_2357);
or U3151 (N_3151,N_2226,N_2370);
and U3152 (N_3152,N_2949,N_2215);
and U3153 (N_3153,N_2133,N_2990);
and U3154 (N_3154,N_2168,N_2197);
and U3155 (N_3155,N_2557,N_2791);
or U3156 (N_3156,N_2522,N_2723);
and U3157 (N_3157,N_2975,N_2112);
nor U3158 (N_3158,N_2036,N_2967);
and U3159 (N_3159,N_2199,N_2871);
and U3160 (N_3160,N_2867,N_2395);
nor U3161 (N_3161,N_2698,N_2886);
or U3162 (N_3162,N_2770,N_2007);
and U3163 (N_3163,N_2753,N_2807);
nand U3164 (N_3164,N_2763,N_2174);
nor U3165 (N_3165,N_2720,N_2629);
nand U3166 (N_3166,N_2993,N_2589);
and U3167 (N_3167,N_2803,N_2637);
and U3168 (N_3168,N_2806,N_2277);
or U3169 (N_3169,N_2567,N_2090);
nor U3170 (N_3170,N_2343,N_2852);
and U3171 (N_3171,N_2538,N_2921);
nand U3172 (N_3172,N_2346,N_2682);
nand U3173 (N_3173,N_2031,N_2527);
nand U3174 (N_3174,N_2067,N_2441);
nor U3175 (N_3175,N_2928,N_2978);
nand U3176 (N_3176,N_2853,N_2628);
nor U3177 (N_3177,N_2862,N_2787);
xnor U3178 (N_3178,N_2696,N_2645);
nor U3179 (N_3179,N_2229,N_2157);
or U3180 (N_3180,N_2953,N_2345);
or U3181 (N_3181,N_2971,N_2190);
or U3182 (N_3182,N_2568,N_2913);
nor U3183 (N_3183,N_2571,N_2042);
or U3184 (N_3184,N_2856,N_2519);
and U3185 (N_3185,N_2458,N_2877);
or U3186 (N_3186,N_2464,N_2639);
and U3187 (N_3187,N_2866,N_2952);
nand U3188 (N_3188,N_2258,N_2825);
nand U3189 (N_3189,N_2830,N_2504);
nor U3190 (N_3190,N_2686,N_2888);
nor U3191 (N_3191,N_2713,N_2431);
or U3192 (N_3192,N_2592,N_2562);
or U3193 (N_3193,N_2531,N_2415);
nor U3194 (N_3194,N_2981,N_2530);
xnor U3195 (N_3195,N_2369,N_2779);
nor U3196 (N_3196,N_2480,N_2879);
nor U3197 (N_3197,N_2863,N_2410);
and U3198 (N_3198,N_2102,N_2261);
nor U3199 (N_3199,N_2390,N_2932);
nand U3200 (N_3200,N_2930,N_2616);
nor U3201 (N_3201,N_2687,N_2761);
nor U3202 (N_3202,N_2010,N_2224);
or U3203 (N_3203,N_2421,N_2584);
or U3204 (N_3204,N_2784,N_2450);
xnor U3205 (N_3205,N_2507,N_2332);
or U3206 (N_3206,N_2494,N_2878);
and U3207 (N_3207,N_2111,N_2559);
or U3208 (N_3208,N_2373,N_2683);
or U3209 (N_3209,N_2603,N_2206);
nor U3210 (N_3210,N_2400,N_2075);
nor U3211 (N_3211,N_2845,N_2247);
and U3212 (N_3212,N_2193,N_2839);
or U3213 (N_3213,N_2336,N_2642);
nor U3214 (N_3214,N_2734,N_2809);
nand U3215 (N_3215,N_2309,N_2231);
or U3216 (N_3216,N_2333,N_2422);
nor U3217 (N_3217,N_2210,N_2204);
xor U3218 (N_3218,N_2292,N_2071);
or U3219 (N_3219,N_2284,N_2021);
nor U3220 (N_3220,N_2935,N_2882);
and U3221 (N_3221,N_2262,N_2281);
nand U3222 (N_3222,N_2374,N_2822);
or U3223 (N_3223,N_2182,N_2691);
nand U3224 (N_3224,N_2950,N_2312);
xnor U3225 (N_3225,N_2468,N_2487);
nand U3226 (N_3226,N_2823,N_2618);
and U3227 (N_3227,N_2044,N_2966);
or U3228 (N_3228,N_2604,N_2363);
nor U3229 (N_3229,N_2566,N_2100);
nand U3230 (N_3230,N_2051,N_2593);
nand U3231 (N_3231,N_2548,N_2194);
xor U3232 (N_3232,N_2581,N_2896);
nand U3233 (N_3233,N_2802,N_2511);
nand U3234 (N_3234,N_2065,N_2173);
nand U3235 (N_3235,N_2518,N_2052);
or U3236 (N_3236,N_2521,N_2499);
xnor U3237 (N_3237,N_2917,N_2965);
nor U3238 (N_3238,N_2478,N_2129);
or U3239 (N_3239,N_2143,N_2785);
nor U3240 (N_3240,N_2163,N_2264);
nor U3241 (N_3241,N_2681,N_2155);
nand U3242 (N_3242,N_2161,N_2964);
xor U3243 (N_3243,N_2362,N_2057);
nor U3244 (N_3244,N_2438,N_2655);
or U3245 (N_3245,N_2925,N_2085);
nor U3246 (N_3246,N_2001,N_2280);
and U3247 (N_3247,N_2819,N_2795);
nand U3248 (N_3248,N_2053,N_2355);
and U3249 (N_3249,N_2137,N_2241);
xnor U3250 (N_3250,N_2936,N_2808);
or U3251 (N_3251,N_2758,N_2520);
and U3252 (N_3252,N_2735,N_2804);
xor U3253 (N_3253,N_2560,N_2598);
nor U3254 (N_3254,N_2897,N_2492);
nor U3255 (N_3255,N_2751,N_2658);
xor U3256 (N_3256,N_2184,N_2166);
xnor U3257 (N_3257,N_2412,N_2994);
or U3258 (N_3258,N_2847,N_2565);
nor U3259 (N_3259,N_2465,N_2668);
nor U3260 (N_3260,N_2019,N_2446);
nand U3261 (N_3261,N_2119,N_2684);
nand U3262 (N_3262,N_2646,N_2982);
or U3263 (N_3263,N_2169,N_2260);
or U3264 (N_3264,N_2831,N_2663);
nor U3265 (N_3265,N_2013,N_2621);
or U3266 (N_3266,N_2269,N_2236);
or U3267 (N_3267,N_2457,N_2657);
and U3268 (N_3268,N_2062,N_2009);
and U3269 (N_3269,N_2301,N_2244);
or U3270 (N_3270,N_2117,N_2265);
or U3271 (N_3271,N_2250,N_2927);
xor U3272 (N_3272,N_2933,N_2669);
xnor U3273 (N_3273,N_2105,N_2101);
xnor U3274 (N_3274,N_2861,N_2054);
or U3275 (N_3275,N_2326,N_2121);
nand U3276 (N_3276,N_2992,N_2167);
xor U3277 (N_3277,N_2767,N_2951);
nand U3278 (N_3278,N_2829,N_2738);
xnor U3279 (N_3279,N_2014,N_2040);
xor U3280 (N_3280,N_2945,N_2324);
xor U3281 (N_3281,N_2685,N_2366);
nor U3282 (N_3282,N_2012,N_2556);
nand U3283 (N_3283,N_2786,N_2626);
or U3284 (N_3284,N_2486,N_2752);
nand U3285 (N_3285,N_2134,N_2742);
or U3286 (N_3286,N_2872,N_2552);
and U3287 (N_3287,N_2389,N_2574);
nor U3288 (N_3288,N_2672,N_2793);
or U3289 (N_3289,N_2656,N_2314);
nor U3290 (N_3290,N_2946,N_2881);
xor U3291 (N_3291,N_2338,N_2388);
nand U3292 (N_3292,N_2467,N_2894);
or U3293 (N_3293,N_2564,N_2123);
nor U3294 (N_3294,N_2462,N_2335);
nor U3295 (N_3295,N_2569,N_2171);
xnor U3296 (N_3296,N_2582,N_2719);
nand U3297 (N_3297,N_2632,N_2183);
or U3298 (N_3298,N_2597,N_2017);
nand U3299 (N_3299,N_2323,N_2063);
nand U3300 (N_3300,N_2360,N_2141);
nor U3301 (N_3301,N_2124,N_2283);
nor U3302 (N_3302,N_2948,N_2865);
nor U3303 (N_3303,N_2573,N_2586);
and U3304 (N_3304,N_2704,N_2246);
xnor U3305 (N_3305,N_2452,N_2903);
nor U3306 (N_3306,N_2242,N_2613);
and U3307 (N_3307,N_2387,N_2003);
and U3308 (N_3308,N_2394,N_2310);
nor U3309 (N_3309,N_2240,N_2282);
nand U3310 (N_3310,N_2503,N_2748);
and U3311 (N_3311,N_2315,N_2187);
nor U3312 (N_3312,N_2596,N_2651);
and U3313 (N_3313,N_2334,N_2033);
xor U3314 (N_3314,N_2110,N_2778);
xor U3315 (N_3315,N_2243,N_2038);
or U3316 (N_3316,N_2475,N_2643);
or U3317 (N_3317,N_2383,N_2311);
nand U3318 (N_3318,N_2186,N_2409);
nand U3319 (N_3319,N_2064,N_2158);
and U3320 (N_3320,N_2329,N_2435);
or U3321 (N_3321,N_2365,N_2147);
nor U3322 (N_3322,N_2154,N_2078);
nor U3323 (N_3323,N_2008,N_2139);
and U3324 (N_3324,N_2252,N_2386);
nor U3325 (N_3325,N_2249,N_2660);
xor U3326 (N_3326,N_2041,N_2726);
nand U3327 (N_3327,N_2270,N_2303);
nand U3328 (N_3328,N_2225,N_2459);
or U3329 (N_3329,N_2901,N_2506);
nand U3330 (N_3330,N_2344,N_2407);
nor U3331 (N_3331,N_2995,N_2047);
or U3332 (N_3332,N_2418,N_2234);
nor U3333 (N_3333,N_2428,N_2500);
and U3334 (N_3334,N_2233,N_2445);
nand U3335 (N_3335,N_2491,N_2620);
nand U3336 (N_3336,N_2178,N_2288);
or U3337 (N_3337,N_2551,N_2255);
nand U3338 (N_3338,N_2188,N_2988);
nor U3339 (N_3339,N_2542,N_2257);
and U3340 (N_3340,N_2074,N_2893);
nand U3341 (N_3341,N_2413,N_2443);
or U3342 (N_3342,N_2179,N_2353);
nand U3343 (N_3343,N_2640,N_2050);
or U3344 (N_3344,N_2032,N_2537);
and U3345 (N_3345,N_2018,N_2035);
nor U3346 (N_3346,N_2875,N_2929);
nor U3347 (N_3347,N_2601,N_2766);
nand U3348 (N_3348,N_2514,N_2706);
and U3349 (N_3349,N_2138,N_2148);
or U3350 (N_3350,N_2069,N_2466);
nand U3351 (N_3351,N_2841,N_2275);
nand U3352 (N_3352,N_2898,N_2230);
xor U3353 (N_3353,N_2826,N_2577);
or U3354 (N_3354,N_2136,N_2423);
nor U3355 (N_3355,N_2772,N_2510);
or U3356 (N_3356,N_2268,N_2473);
nand U3357 (N_3357,N_2088,N_2484);
or U3358 (N_3358,N_2732,N_2754);
nand U3359 (N_3359,N_2020,N_2399);
and U3360 (N_3360,N_2483,N_2397);
and U3361 (N_3361,N_2606,N_2059);
nor U3362 (N_3362,N_2223,N_2140);
nor U3363 (N_3363,N_2776,N_2768);
or U3364 (N_3364,N_2623,N_2570);
nor U3365 (N_3365,N_2765,N_2097);
and U3366 (N_3366,N_2539,N_2891);
nor U3367 (N_3367,N_2840,N_2756);
and U3368 (N_3368,N_2638,N_2549);
and U3369 (N_3369,N_2940,N_2393);
xnor U3370 (N_3370,N_2533,N_2859);
and U3371 (N_3371,N_2296,N_2172);
xnor U3372 (N_3372,N_2543,N_2773);
nand U3373 (N_3373,N_2931,N_2440);
and U3374 (N_3374,N_2860,N_2892);
or U3375 (N_3375,N_2000,N_2870);
and U3376 (N_3376,N_2600,N_2294);
nand U3377 (N_3377,N_2805,N_2472);
nor U3378 (N_3378,N_2817,N_2680);
xor U3379 (N_3379,N_2515,N_2434);
and U3380 (N_3380,N_2490,N_2248);
or U3381 (N_3381,N_2788,N_2524);
nand U3382 (N_3382,N_2424,N_2376);
and U3383 (N_3383,N_2045,N_2084);
nor U3384 (N_3384,N_2325,N_2330);
or U3385 (N_3385,N_2816,N_2650);
nand U3386 (N_3386,N_2939,N_2381);
or U3387 (N_3387,N_2890,N_2699);
nand U3388 (N_3388,N_2730,N_2476);
nand U3389 (N_3389,N_2276,N_2725);
xor U3390 (N_3390,N_2908,N_2358);
nand U3391 (N_3391,N_2253,N_2916);
nor U3392 (N_3392,N_2835,N_2703);
nand U3393 (N_3393,N_2529,N_2740);
nor U3394 (N_3394,N_2212,N_2361);
or U3395 (N_3395,N_2576,N_2707);
or U3396 (N_3396,N_2115,N_2887);
nand U3397 (N_3397,N_2671,N_2060);
xor U3398 (N_3398,N_2191,N_2113);
nor U3399 (N_3399,N_2056,N_2082);
nand U3400 (N_3400,N_2165,N_2454);
nand U3401 (N_3401,N_2717,N_2644);
nand U3402 (N_3402,N_2918,N_2274);
xor U3403 (N_3403,N_2777,N_2341);
nand U3404 (N_3404,N_2149,N_2532);
and U3405 (N_3405,N_2963,N_2782);
nor U3406 (N_3406,N_2973,N_2814);
or U3407 (N_3407,N_2026,N_2858);
xor U3408 (N_3408,N_2528,N_2594);
nor U3409 (N_3409,N_2437,N_2590);
nor U3410 (N_3410,N_2377,N_2222);
nor U3411 (N_3411,N_2039,N_2104);
or U3412 (N_3412,N_2512,N_2076);
nand U3413 (N_3413,N_2128,N_2485);
nor U3414 (N_3414,N_2227,N_2153);
and U3415 (N_3415,N_2444,N_2976);
nor U3416 (N_3416,N_2316,N_2120);
or U3417 (N_3417,N_2022,N_2209);
and U3418 (N_3418,N_2970,N_2456);
and U3419 (N_3419,N_2540,N_2449);
or U3420 (N_3420,N_2200,N_2667);
or U3421 (N_3421,N_2716,N_2151);
nor U3422 (N_3422,N_2356,N_2259);
and U3423 (N_3423,N_2757,N_2408);
nand U3424 (N_3424,N_2291,N_2347);
and U3425 (N_3425,N_2857,N_2801);
or U3426 (N_3426,N_2203,N_2924);
or U3427 (N_3427,N_2402,N_2378);
nor U3428 (N_3428,N_2999,N_2185);
xnor U3429 (N_3429,N_2380,N_2055);
nor U3430 (N_3430,N_2678,N_2909);
and U3431 (N_3431,N_2218,N_2868);
and U3432 (N_3432,N_2648,N_2331);
nor U3433 (N_3433,N_2011,N_2907);
nand U3434 (N_3434,N_2615,N_2299);
and U3435 (N_3435,N_2665,N_2688);
nor U3436 (N_3436,N_2895,N_2714);
or U3437 (N_3437,N_2364,N_2372);
xor U3438 (N_3438,N_2563,N_2692);
or U3439 (N_3439,N_2534,N_2419);
nor U3440 (N_3440,N_2368,N_2986);
nor U3441 (N_3441,N_2479,N_2769);
or U3442 (N_3442,N_2118,N_2232);
or U3443 (N_3443,N_2579,N_2216);
nor U3444 (N_3444,N_2046,N_2072);
or U3445 (N_3445,N_2207,N_2453);
nand U3446 (N_3446,N_2066,N_2305);
or U3447 (N_3447,N_2588,N_2834);
nand U3448 (N_3448,N_2972,N_2116);
or U3449 (N_3449,N_2824,N_2214);
or U3450 (N_3450,N_2984,N_2739);
and U3451 (N_3451,N_2477,N_2278);
nor U3452 (N_3452,N_2670,N_2693);
or U3453 (N_3453,N_2096,N_2561);
nor U3454 (N_3454,N_2439,N_2635);
or U3455 (N_3455,N_2436,N_2622);
or U3456 (N_3456,N_2342,N_2575);
nand U3457 (N_3457,N_2433,N_2221);
or U3458 (N_3458,N_2796,N_2285);
nand U3459 (N_3459,N_2955,N_2416);
and U3460 (N_3460,N_2132,N_2884);
xor U3461 (N_3461,N_2505,N_2427);
xnor U3462 (N_3462,N_2849,N_2162);
nor U3463 (N_3463,N_2306,N_2016);
nand U3464 (N_3464,N_2545,N_2508);
nor U3465 (N_3465,N_2996,N_2429);
or U3466 (N_3466,N_2631,N_2546);
or U3467 (N_3467,N_2002,N_2905);
or U3468 (N_3468,N_2876,N_2958);
nor U3469 (N_3469,N_2869,N_2430);
and U3470 (N_3470,N_2048,N_2662);
or U3471 (N_3471,N_2605,N_2122);
nor U3472 (N_3472,N_2189,N_2501);
or U3473 (N_3473,N_2711,N_2709);
and U3474 (N_3474,N_2602,N_2902);
and U3475 (N_3475,N_2398,N_2488);
and U3476 (N_3476,N_2915,N_2080);
nor U3477 (N_3477,N_2371,N_2348);
and U3478 (N_3478,N_2513,N_2922);
and U3479 (N_3479,N_2674,N_2083);
and U3480 (N_3480,N_2401,N_2525);
or U3481 (N_3481,N_2030,N_2764);
nor U3482 (N_3482,N_2800,N_2883);
nand U3483 (N_3483,N_2037,N_2997);
nand U3484 (N_3484,N_2279,N_2775);
or U3485 (N_3485,N_2583,N_2098);
nor U3486 (N_3486,N_2612,N_2004);
or U3487 (N_3487,N_2339,N_2985);
nor U3488 (N_3488,N_2447,N_2979);
nand U3489 (N_3489,N_2854,N_2482);
xnor U3490 (N_3490,N_2319,N_2614);
nand U3491 (N_3491,N_2718,N_2127);
or U3492 (N_3492,N_2385,N_2938);
or U3493 (N_3493,N_2196,N_2442);
nand U3494 (N_3494,N_2661,N_2295);
nand U3495 (N_3495,N_2432,N_2448);
nor U3496 (N_3496,N_2855,N_2673);
and U3497 (N_3497,N_2461,N_2926);
nand U3498 (N_3498,N_2794,N_2195);
and U3499 (N_3499,N_2131,N_2109);
or U3500 (N_3500,N_2618,N_2887);
or U3501 (N_3501,N_2843,N_2366);
and U3502 (N_3502,N_2900,N_2419);
or U3503 (N_3503,N_2239,N_2501);
nand U3504 (N_3504,N_2578,N_2043);
and U3505 (N_3505,N_2182,N_2601);
nand U3506 (N_3506,N_2738,N_2048);
nor U3507 (N_3507,N_2787,N_2598);
and U3508 (N_3508,N_2676,N_2762);
or U3509 (N_3509,N_2699,N_2286);
and U3510 (N_3510,N_2815,N_2791);
or U3511 (N_3511,N_2497,N_2976);
and U3512 (N_3512,N_2732,N_2513);
xnor U3513 (N_3513,N_2852,N_2523);
and U3514 (N_3514,N_2140,N_2576);
or U3515 (N_3515,N_2639,N_2475);
xor U3516 (N_3516,N_2987,N_2950);
nor U3517 (N_3517,N_2266,N_2404);
nand U3518 (N_3518,N_2817,N_2974);
or U3519 (N_3519,N_2772,N_2167);
nor U3520 (N_3520,N_2597,N_2614);
and U3521 (N_3521,N_2478,N_2796);
nor U3522 (N_3522,N_2291,N_2356);
nand U3523 (N_3523,N_2740,N_2973);
nor U3524 (N_3524,N_2143,N_2706);
and U3525 (N_3525,N_2627,N_2751);
xnor U3526 (N_3526,N_2695,N_2743);
nand U3527 (N_3527,N_2798,N_2146);
nor U3528 (N_3528,N_2155,N_2209);
nor U3529 (N_3529,N_2278,N_2276);
or U3530 (N_3530,N_2151,N_2857);
and U3531 (N_3531,N_2323,N_2904);
nor U3532 (N_3532,N_2004,N_2293);
or U3533 (N_3533,N_2741,N_2291);
or U3534 (N_3534,N_2703,N_2341);
nor U3535 (N_3535,N_2390,N_2952);
nor U3536 (N_3536,N_2883,N_2607);
xnor U3537 (N_3537,N_2918,N_2022);
nor U3538 (N_3538,N_2299,N_2429);
xor U3539 (N_3539,N_2035,N_2047);
nor U3540 (N_3540,N_2700,N_2919);
nor U3541 (N_3541,N_2274,N_2386);
nor U3542 (N_3542,N_2322,N_2566);
xor U3543 (N_3543,N_2895,N_2728);
and U3544 (N_3544,N_2528,N_2989);
nand U3545 (N_3545,N_2684,N_2188);
xor U3546 (N_3546,N_2645,N_2022);
and U3547 (N_3547,N_2340,N_2533);
nor U3548 (N_3548,N_2921,N_2901);
and U3549 (N_3549,N_2637,N_2167);
nand U3550 (N_3550,N_2402,N_2093);
or U3551 (N_3551,N_2541,N_2782);
or U3552 (N_3552,N_2901,N_2676);
xnor U3553 (N_3553,N_2664,N_2060);
nand U3554 (N_3554,N_2006,N_2755);
and U3555 (N_3555,N_2564,N_2277);
nand U3556 (N_3556,N_2925,N_2814);
nor U3557 (N_3557,N_2359,N_2099);
or U3558 (N_3558,N_2370,N_2879);
nor U3559 (N_3559,N_2776,N_2040);
and U3560 (N_3560,N_2119,N_2046);
and U3561 (N_3561,N_2929,N_2883);
and U3562 (N_3562,N_2616,N_2596);
nand U3563 (N_3563,N_2846,N_2122);
nand U3564 (N_3564,N_2653,N_2769);
xor U3565 (N_3565,N_2489,N_2039);
and U3566 (N_3566,N_2331,N_2884);
or U3567 (N_3567,N_2061,N_2247);
nand U3568 (N_3568,N_2285,N_2848);
nand U3569 (N_3569,N_2197,N_2821);
or U3570 (N_3570,N_2047,N_2058);
and U3571 (N_3571,N_2404,N_2394);
nor U3572 (N_3572,N_2947,N_2132);
xnor U3573 (N_3573,N_2844,N_2120);
nand U3574 (N_3574,N_2002,N_2454);
nor U3575 (N_3575,N_2545,N_2774);
or U3576 (N_3576,N_2877,N_2430);
or U3577 (N_3577,N_2053,N_2475);
nand U3578 (N_3578,N_2216,N_2679);
and U3579 (N_3579,N_2136,N_2291);
and U3580 (N_3580,N_2417,N_2468);
and U3581 (N_3581,N_2512,N_2342);
nand U3582 (N_3582,N_2587,N_2028);
nor U3583 (N_3583,N_2248,N_2683);
or U3584 (N_3584,N_2757,N_2350);
nor U3585 (N_3585,N_2952,N_2063);
nand U3586 (N_3586,N_2578,N_2861);
nand U3587 (N_3587,N_2381,N_2605);
or U3588 (N_3588,N_2366,N_2742);
nand U3589 (N_3589,N_2909,N_2143);
or U3590 (N_3590,N_2524,N_2432);
nand U3591 (N_3591,N_2520,N_2977);
nand U3592 (N_3592,N_2928,N_2476);
nand U3593 (N_3593,N_2680,N_2132);
nand U3594 (N_3594,N_2341,N_2837);
nand U3595 (N_3595,N_2411,N_2522);
nor U3596 (N_3596,N_2548,N_2532);
nor U3597 (N_3597,N_2387,N_2335);
or U3598 (N_3598,N_2927,N_2459);
and U3599 (N_3599,N_2805,N_2323);
xnor U3600 (N_3600,N_2505,N_2327);
nor U3601 (N_3601,N_2429,N_2560);
or U3602 (N_3602,N_2575,N_2173);
nor U3603 (N_3603,N_2601,N_2126);
nand U3604 (N_3604,N_2168,N_2245);
and U3605 (N_3605,N_2266,N_2869);
or U3606 (N_3606,N_2429,N_2546);
or U3607 (N_3607,N_2734,N_2004);
and U3608 (N_3608,N_2396,N_2905);
nand U3609 (N_3609,N_2091,N_2228);
or U3610 (N_3610,N_2926,N_2247);
xnor U3611 (N_3611,N_2512,N_2945);
or U3612 (N_3612,N_2127,N_2619);
nor U3613 (N_3613,N_2674,N_2841);
nor U3614 (N_3614,N_2900,N_2690);
nand U3615 (N_3615,N_2560,N_2065);
nand U3616 (N_3616,N_2815,N_2010);
nand U3617 (N_3617,N_2044,N_2768);
nand U3618 (N_3618,N_2709,N_2254);
nor U3619 (N_3619,N_2096,N_2896);
and U3620 (N_3620,N_2798,N_2541);
nand U3621 (N_3621,N_2125,N_2984);
nand U3622 (N_3622,N_2187,N_2345);
nand U3623 (N_3623,N_2465,N_2233);
or U3624 (N_3624,N_2642,N_2198);
nor U3625 (N_3625,N_2840,N_2394);
and U3626 (N_3626,N_2670,N_2216);
nor U3627 (N_3627,N_2427,N_2300);
or U3628 (N_3628,N_2674,N_2517);
xnor U3629 (N_3629,N_2889,N_2384);
nor U3630 (N_3630,N_2499,N_2130);
and U3631 (N_3631,N_2921,N_2690);
xnor U3632 (N_3632,N_2843,N_2423);
or U3633 (N_3633,N_2048,N_2111);
or U3634 (N_3634,N_2265,N_2647);
xor U3635 (N_3635,N_2701,N_2934);
nor U3636 (N_3636,N_2688,N_2539);
nor U3637 (N_3637,N_2845,N_2554);
nor U3638 (N_3638,N_2639,N_2747);
and U3639 (N_3639,N_2351,N_2914);
or U3640 (N_3640,N_2876,N_2436);
and U3641 (N_3641,N_2497,N_2712);
nand U3642 (N_3642,N_2466,N_2050);
nor U3643 (N_3643,N_2583,N_2715);
or U3644 (N_3644,N_2433,N_2599);
nand U3645 (N_3645,N_2511,N_2589);
or U3646 (N_3646,N_2840,N_2672);
nand U3647 (N_3647,N_2656,N_2870);
xor U3648 (N_3648,N_2729,N_2644);
xor U3649 (N_3649,N_2499,N_2908);
xnor U3650 (N_3650,N_2612,N_2969);
and U3651 (N_3651,N_2243,N_2065);
nand U3652 (N_3652,N_2816,N_2854);
nor U3653 (N_3653,N_2699,N_2651);
and U3654 (N_3654,N_2769,N_2241);
or U3655 (N_3655,N_2458,N_2242);
or U3656 (N_3656,N_2587,N_2388);
and U3657 (N_3657,N_2385,N_2536);
nand U3658 (N_3658,N_2233,N_2418);
or U3659 (N_3659,N_2492,N_2138);
nor U3660 (N_3660,N_2300,N_2365);
or U3661 (N_3661,N_2807,N_2276);
or U3662 (N_3662,N_2505,N_2780);
and U3663 (N_3663,N_2811,N_2385);
nor U3664 (N_3664,N_2250,N_2157);
nor U3665 (N_3665,N_2673,N_2297);
or U3666 (N_3666,N_2375,N_2496);
nand U3667 (N_3667,N_2396,N_2534);
nor U3668 (N_3668,N_2728,N_2830);
nor U3669 (N_3669,N_2135,N_2563);
and U3670 (N_3670,N_2658,N_2777);
nand U3671 (N_3671,N_2969,N_2150);
and U3672 (N_3672,N_2676,N_2291);
xor U3673 (N_3673,N_2155,N_2436);
nor U3674 (N_3674,N_2968,N_2851);
nor U3675 (N_3675,N_2184,N_2657);
nor U3676 (N_3676,N_2401,N_2889);
or U3677 (N_3677,N_2358,N_2285);
xor U3678 (N_3678,N_2063,N_2917);
and U3679 (N_3679,N_2605,N_2884);
and U3680 (N_3680,N_2216,N_2863);
nand U3681 (N_3681,N_2527,N_2937);
and U3682 (N_3682,N_2103,N_2644);
and U3683 (N_3683,N_2931,N_2183);
and U3684 (N_3684,N_2989,N_2539);
nand U3685 (N_3685,N_2382,N_2095);
and U3686 (N_3686,N_2110,N_2002);
or U3687 (N_3687,N_2836,N_2874);
xor U3688 (N_3688,N_2486,N_2286);
nor U3689 (N_3689,N_2545,N_2977);
nor U3690 (N_3690,N_2941,N_2877);
and U3691 (N_3691,N_2380,N_2210);
or U3692 (N_3692,N_2164,N_2340);
nor U3693 (N_3693,N_2641,N_2389);
nand U3694 (N_3694,N_2422,N_2164);
and U3695 (N_3695,N_2989,N_2140);
xnor U3696 (N_3696,N_2543,N_2443);
and U3697 (N_3697,N_2102,N_2643);
nand U3698 (N_3698,N_2842,N_2892);
nor U3699 (N_3699,N_2863,N_2148);
or U3700 (N_3700,N_2018,N_2176);
and U3701 (N_3701,N_2069,N_2884);
and U3702 (N_3702,N_2300,N_2309);
nand U3703 (N_3703,N_2302,N_2130);
nor U3704 (N_3704,N_2153,N_2475);
or U3705 (N_3705,N_2737,N_2394);
nand U3706 (N_3706,N_2468,N_2239);
or U3707 (N_3707,N_2992,N_2106);
nand U3708 (N_3708,N_2509,N_2671);
nor U3709 (N_3709,N_2291,N_2620);
xor U3710 (N_3710,N_2088,N_2653);
nand U3711 (N_3711,N_2045,N_2337);
or U3712 (N_3712,N_2180,N_2509);
nor U3713 (N_3713,N_2625,N_2507);
or U3714 (N_3714,N_2978,N_2989);
nor U3715 (N_3715,N_2296,N_2229);
nor U3716 (N_3716,N_2410,N_2247);
nand U3717 (N_3717,N_2138,N_2926);
nor U3718 (N_3718,N_2151,N_2794);
nand U3719 (N_3719,N_2220,N_2252);
and U3720 (N_3720,N_2996,N_2304);
or U3721 (N_3721,N_2137,N_2634);
or U3722 (N_3722,N_2370,N_2109);
nand U3723 (N_3723,N_2892,N_2064);
and U3724 (N_3724,N_2129,N_2704);
or U3725 (N_3725,N_2673,N_2841);
or U3726 (N_3726,N_2627,N_2613);
or U3727 (N_3727,N_2643,N_2687);
xnor U3728 (N_3728,N_2354,N_2787);
nand U3729 (N_3729,N_2519,N_2683);
nor U3730 (N_3730,N_2436,N_2195);
nor U3731 (N_3731,N_2856,N_2103);
nand U3732 (N_3732,N_2510,N_2910);
nand U3733 (N_3733,N_2416,N_2669);
nor U3734 (N_3734,N_2080,N_2064);
and U3735 (N_3735,N_2463,N_2180);
and U3736 (N_3736,N_2008,N_2502);
and U3737 (N_3737,N_2967,N_2276);
and U3738 (N_3738,N_2061,N_2592);
nand U3739 (N_3739,N_2906,N_2702);
or U3740 (N_3740,N_2974,N_2249);
nand U3741 (N_3741,N_2402,N_2169);
xor U3742 (N_3742,N_2313,N_2241);
nand U3743 (N_3743,N_2322,N_2923);
xor U3744 (N_3744,N_2634,N_2644);
nor U3745 (N_3745,N_2560,N_2710);
nand U3746 (N_3746,N_2603,N_2884);
nand U3747 (N_3747,N_2458,N_2212);
nor U3748 (N_3748,N_2261,N_2873);
or U3749 (N_3749,N_2981,N_2258);
or U3750 (N_3750,N_2048,N_2694);
nor U3751 (N_3751,N_2210,N_2232);
xnor U3752 (N_3752,N_2428,N_2726);
and U3753 (N_3753,N_2713,N_2200);
or U3754 (N_3754,N_2122,N_2280);
or U3755 (N_3755,N_2016,N_2243);
nand U3756 (N_3756,N_2579,N_2974);
nor U3757 (N_3757,N_2450,N_2280);
or U3758 (N_3758,N_2687,N_2711);
or U3759 (N_3759,N_2198,N_2841);
nand U3760 (N_3760,N_2348,N_2205);
xnor U3761 (N_3761,N_2570,N_2706);
nor U3762 (N_3762,N_2400,N_2104);
nor U3763 (N_3763,N_2200,N_2618);
nand U3764 (N_3764,N_2640,N_2117);
and U3765 (N_3765,N_2324,N_2389);
nor U3766 (N_3766,N_2289,N_2702);
nor U3767 (N_3767,N_2609,N_2752);
and U3768 (N_3768,N_2065,N_2095);
nor U3769 (N_3769,N_2044,N_2590);
nand U3770 (N_3770,N_2786,N_2047);
nand U3771 (N_3771,N_2469,N_2068);
and U3772 (N_3772,N_2678,N_2390);
nand U3773 (N_3773,N_2520,N_2237);
or U3774 (N_3774,N_2598,N_2037);
and U3775 (N_3775,N_2882,N_2513);
and U3776 (N_3776,N_2588,N_2211);
nor U3777 (N_3777,N_2653,N_2931);
and U3778 (N_3778,N_2214,N_2627);
nor U3779 (N_3779,N_2757,N_2489);
or U3780 (N_3780,N_2742,N_2394);
nor U3781 (N_3781,N_2361,N_2028);
and U3782 (N_3782,N_2043,N_2339);
and U3783 (N_3783,N_2416,N_2879);
nor U3784 (N_3784,N_2548,N_2500);
nor U3785 (N_3785,N_2455,N_2243);
nand U3786 (N_3786,N_2912,N_2457);
nand U3787 (N_3787,N_2894,N_2837);
nand U3788 (N_3788,N_2953,N_2817);
xnor U3789 (N_3789,N_2235,N_2520);
or U3790 (N_3790,N_2997,N_2090);
and U3791 (N_3791,N_2980,N_2932);
or U3792 (N_3792,N_2711,N_2752);
nor U3793 (N_3793,N_2229,N_2310);
and U3794 (N_3794,N_2094,N_2531);
or U3795 (N_3795,N_2317,N_2958);
or U3796 (N_3796,N_2521,N_2043);
nor U3797 (N_3797,N_2908,N_2317);
or U3798 (N_3798,N_2423,N_2698);
nand U3799 (N_3799,N_2692,N_2341);
nor U3800 (N_3800,N_2726,N_2807);
nand U3801 (N_3801,N_2054,N_2243);
nor U3802 (N_3802,N_2814,N_2638);
nor U3803 (N_3803,N_2431,N_2383);
nand U3804 (N_3804,N_2334,N_2658);
xor U3805 (N_3805,N_2612,N_2484);
and U3806 (N_3806,N_2291,N_2248);
xor U3807 (N_3807,N_2403,N_2378);
or U3808 (N_3808,N_2040,N_2076);
nor U3809 (N_3809,N_2588,N_2547);
nand U3810 (N_3810,N_2961,N_2160);
nor U3811 (N_3811,N_2799,N_2724);
nand U3812 (N_3812,N_2960,N_2572);
nand U3813 (N_3813,N_2744,N_2020);
nand U3814 (N_3814,N_2561,N_2785);
and U3815 (N_3815,N_2255,N_2133);
nand U3816 (N_3816,N_2537,N_2730);
nand U3817 (N_3817,N_2134,N_2611);
and U3818 (N_3818,N_2150,N_2693);
nor U3819 (N_3819,N_2149,N_2067);
or U3820 (N_3820,N_2059,N_2143);
and U3821 (N_3821,N_2354,N_2888);
nand U3822 (N_3822,N_2878,N_2055);
or U3823 (N_3823,N_2923,N_2386);
xor U3824 (N_3824,N_2023,N_2631);
nand U3825 (N_3825,N_2307,N_2516);
nand U3826 (N_3826,N_2776,N_2330);
nor U3827 (N_3827,N_2472,N_2914);
or U3828 (N_3828,N_2645,N_2828);
and U3829 (N_3829,N_2963,N_2528);
or U3830 (N_3830,N_2207,N_2410);
nor U3831 (N_3831,N_2014,N_2658);
nor U3832 (N_3832,N_2729,N_2444);
and U3833 (N_3833,N_2318,N_2978);
xor U3834 (N_3834,N_2566,N_2573);
nor U3835 (N_3835,N_2375,N_2668);
nor U3836 (N_3836,N_2493,N_2366);
and U3837 (N_3837,N_2669,N_2903);
or U3838 (N_3838,N_2261,N_2752);
nor U3839 (N_3839,N_2200,N_2890);
nor U3840 (N_3840,N_2322,N_2301);
nor U3841 (N_3841,N_2380,N_2635);
nand U3842 (N_3842,N_2945,N_2062);
and U3843 (N_3843,N_2324,N_2549);
nand U3844 (N_3844,N_2959,N_2752);
or U3845 (N_3845,N_2525,N_2364);
nand U3846 (N_3846,N_2370,N_2729);
or U3847 (N_3847,N_2914,N_2159);
nand U3848 (N_3848,N_2238,N_2021);
nor U3849 (N_3849,N_2139,N_2448);
nand U3850 (N_3850,N_2920,N_2632);
nor U3851 (N_3851,N_2928,N_2426);
or U3852 (N_3852,N_2567,N_2630);
xnor U3853 (N_3853,N_2611,N_2386);
nor U3854 (N_3854,N_2033,N_2999);
nand U3855 (N_3855,N_2559,N_2170);
or U3856 (N_3856,N_2450,N_2779);
or U3857 (N_3857,N_2851,N_2687);
and U3858 (N_3858,N_2755,N_2973);
nor U3859 (N_3859,N_2471,N_2856);
nand U3860 (N_3860,N_2366,N_2904);
nand U3861 (N_3861,N_2118,N_2686);
nor U3862 (N_3862,N_2240,N_2693);
nand U3863 (N_3863,N_2274,N_2512);
or U3864 (N_3864,N_2662,N_2813);
nor U3865 (N_3865,N_2700,N_2645);
or U3866 (N_3866,N_2473,N_2054);
or U3867 (N_3867,N_2992,N_2285);
nor U3868 (N_3868,N_2036,N_2958);
nand U3869 (N_3869,N_2911,N_2922);
or U3870 (N_3870,N_2537,N_2612);
nand U3871 (N_3871,N_2580,N_2656);
nor U3872 (N_3872,N_2234,N_2681);
and U3873 (N_3873,N_2794,N_2000);
or U3874 (N_3874,N_2759,N_2689);
nor U3875 (N_3875,N_2475,N_2318);
or U3876 (N_3876,N_2927,N_2159);
or U3877 (N_3877,N_2602,N_2093);
and U3878 (N_3878,N_2157,N_2891);
or U3879 (N_3879,N_2957,N_2837);
nor U3880 (N_3880,N_2869,N_2196);
nor U3881 (N_3881,N_2749,N_2601);
nor U3882 (N_3882,N_2775,N_2469);
nand U3883 (N_3883,N_2902,N_2146);
or U3884 (N_3884,N_2259,N_2396);
nor U3885 (N_3885,N_2274,N_2890);
and U3886 (N_3886,N_2334,N_2694);
nand U3887 (N_3887,N_2888,N_2106);
xnor U3888 (N_3888,N_2097,N_2574);
nor U3889 (N_3889,N_2787,N_2942);
and U3890 (N_3890,N_2726,N_2125);
nor U3891 (N_3891,N_2826,N_2694);
or U3892 (N_3892,N_2340,N_2299);
and U3893 (N_3893,N_2602,N_2984);
nor U3894 (N_3894,N_2106,N_2836);
nor U3895 (N_3895,N_2770,N_2293);
nand U3896 (N_3896,N_2900,N_2587);
and U3897 (N_3897,N_2920,N_2617);
nor U3898 (N_3898,N_2460,N_2583);
nor U3899 (N_3899,N_2847,N_2993);
and U3900 (N_3900,N_2911,N_2857);
and U3901 (N_3901,N_2047,N_2782);
nand U3902 (N_3902,N_2539,N_2100);
or U3903 (N_3903,N_2616,N_2960);
xnor U3904 (N_3904,N_2771,N_2657);
and U3905 (N_3905,N_2015,N_2980);
and U3906 (N_3906,N_2074,N_2850);
or U3907 (N_3907,N_2036,N_2368);
nor U3908 (N_3908,N_2774,N_2230);
and U3909 (N_3909,N_2926,N_2338);
or U3910 (N_3910,N_2881,N_2170);
or U3911 (N_3911,N_2734,N_2660);
or U3912 (N_3912,N_2514,N_2677);
nand U3913 (N_3913,N_2243,N_2638);
nand U3914 (N_3914,N_2130,N_2006);
and U3915 (N_3915,N_2751,N_2164);
and U3916 (N_3916,N_2263,N_2515);
and U3917 (N_3917,N_2682,N_2110);
nor U3918 (N_3918,N_2011,N_2988);
and U3919 (N_3919,N_2899,N_2195);
and U3920 (N_3920,N_2018,N_2451);
or U3921 (N_3921,N_2094,N_2982);
and U3922 (N_3922,N_2015,N_2073);
or U3923 (N_3923,N_2822,N_2997);
or U3924 (N_3924,N_2112,N_2373);
xnor U3925 (N_3925,N_2510,N_2316);
nor U3926 (N_3926,N_2079,N_2160);
and U3927 (N_3927,N_2053,N_2971);
xor U3928 (N_3928,N_2536,N_2670);
xnor U3929 (N_3929,N_2472,N_2602);
nand U3930 (N_3930,N_2583,N_2386);
xor U3931 (N_3931,N_2336,N_2833);
xor U3932 (N_3932,N_2912,N_2000);
or U3933 (N_3933,N_2629,N_2490);
nor U3934 (N_3934,N_2315,N_2399);
nand U3935 (N_3935,N_2650,N_2501);
nor U3936 (N_3936,N_2034,N_2887);
nand U3937 (N_3937,N_2426,N_2339);
nor U3938 (N_3938,N_2092,N_2267);
or U3939 (N_3939,N_2521,N_2526);
nand U3940 (N_3940,N_2871,N_2490);
nor U3941 (N_3941,N_2795,N_2606);
and U3942 (N_3942,N_2202,N_2692);
and U3943 (N_3943,N_2148,N_2427);
nor U3944 (N_3944,N_2126,N_2142);
nor U3945 (N_3945,N_2297,N_2371);
and U3946 (N_3946,N_2840,N_2639);
nand U3947 (N_3947,N_2772,N_2451);
or U3948 (N_3948,N_2139,N_2577);
nor U3949 (N_3949,N_2070,N_2504);
and U3950 (N_3950,N_2103,N_2818);
nand U3951 (N_3951,N_2339,N_2056);
nand U3952 (N_3952,N_2951,N_2789);
and U3953 (N_3953,N_2417,N_2655);
or U3954 (N_3954,N_2063,N_2124);
or U3955 (N_3955,N_2162,N_2291);
nand U3956 (N_3956,N_2874,N_2258);
nor U3957 (N_3957,N_2454,N_2025);
nand U3958 (N_3958,N_2425,N_2335);
nand U3959 (N_3959,N_2795,N_2856);
nand U3960 (N_3960,N_2101,N_2152);
or U3961 (N_3961,N_2585,N_2131);
or U3962 (N_3962,N_2503,N_2795);
or U3963 (N_3963,N_2971,N_2526);
or U3964 (N_3964,N_2868,N_2040);
nand U3965 (N_3965,N_2635,N_2012);
nor U3966 (N_3966,N_2705,N_2927);
nand U3967 (N_3967,N_2001,N_2235);
or U3968 (N_3968,N_2832,N_2298);
nand U3969 (N_3969,N_2857,N_2575);
xor U3970 (N_3970,N_2011,N_2072);
and U3971 (N_3971,N_2968,N_2625);
nand U3972 (N_3972,N_2182,N_2325);
nand U3973 (N_3973,N_2264,N_2518);
or U3974 (N_3974,N_2927,N_2622);
or U3975 (N_3975,N_2237,N_2280);
nand U3976 (N_3976,N_2027,N_2771);
xnor U3977 (N_3977,N_2875,N_2576);
or U3978 (N_3978,N_2374,N_2919);
and U3979 (N_3979,N_2231,N_2414);
and U3980 (N_3980,N_2077,N_2887);
nor U3981 (N_3981,N_2081,N_2039);
or U3982 (N_3982,N_2210,N_2023);
nand U3983 (N_3983,N_2985,N_2117);
and U3984 (N_3984,N_2569,N_2755);
nor U3985 (N_3985,N_2202,N_2043);
nor U3986 (N_3986,N_2686,N_2925);
nand U3987 (N_3987,N_2730,N_2972);
or U3988 (N_3988,N_2869,N_2263);
nand U3989 (N_3989,N_2846,N_2458);
nor U3990 (N_3990,N_2891,N_2474);
or U3991 (N_3991,N_2763,N_2057);
nor U3992 (N_3992,N_2957,N_2413);
nand U3993 (N_3993,N_2630,N_2218);
or U3994 (N_3994,N_2286,N_2779);
nor U3995 (N_3995,N_2375,N_2155);
or U3996 (N_3996,N_2195,N_2097);
xor U3997 (N_3997,N_2384,N_2774);
and U3998 (N_3998,N_2970,N_2342);
nor U3999 (N_3999,N_2498,N_2699);
and U4000 (N_4000,N_3721,N_3652);
xnor U4001 (N_4001,N_3846,N_3364);
nor U4002 (N_4002,N_3768,N_3182);
nand U4003 (N_4003,N_3709,N_3510);
or U4004 (N_4004,N_3617,N_3308);
or U4005 (N_4005,N_3203,N_3581);
or U4006 (N_4006,N_3130,N_3782);
nand U4007 (N_4007,N_3775,N_3329);
xnor U4008 (N_4008,N_3878,N_3834);
nor U4009 (N_4009,N_3994,N_3697);
nand U4010 (N_4010,N_3419,N_3309);
or U4011 (N_4011,N_3330,N_3351);
and U4012 (N_4012,N_3444,N_3409);
xor U4013 (N_4013,N_3575,N_3648);
xnor U4014 (N_4014,N_3109,N_3734);
or U4015 (N_4015,N_3475,N_3976);
nand U4016 (N_4016,N_3081,N_3959);
nor U4017 (N_4017,N_3772,N_3625);
nor U4018 (N_4018,N_3894,N_3265);
or U4019 (N_4019,N_3525,N_3277);
nor U4020 (N_4020,N_3234,N_3074);
nand U4021 (N_4021,N_3505,N_3570);
nor U4022 (N_4022,N_3369,N_3898);
nor U4023 (N_4023,N_3428,N_3835);
nand U4024 (N_4024,N_3354,N_3950);
or U4025 (N_4025,N_3091,N_3261);
xor U4026 (N_4026,N_3357,N_3170);
xor U4027 (N_4027,N_3229,N_3268);
and U4028 (N_4028,N_3181,N_3259);
nand U4029 (N_4029,N_3951,N_3741);
and U4030 (N_4030,N_3923,N_3387);
or U4031 (N_4031,N_3822,N_3438);
nand U4032 (N_4032,N_3703,N_3078);
or U4033 (N_4033,N_3820,N_3436);
nand U4034 (N_4034,N_3698,N_3283);
nand U4035 (N_4035,N_3889,N_3397);
nor U4036 (N_4036,N_3190,N_3803);
xor U4037 (N_4037,N_3016,N_3664);
or U4038 (N_4038,N_3430,N_3879);
and U4039 (N_4039,N_3727,N_3897);
or U4040 (N_4040,N_3928,N_3589);
nand U4041 (N_4041,N_3314,N_3723);
nand U4042 (N_4042,N_3830,N_3195);
nand U4043 (N_4043,N_3827,N_3967);
and U4044 (N_4044,N_3949,N_3205);
nor U4045 (N_4045,N_3416,N_3569);
nor U4046 (N_4046,N_3210,N_3502);
xnor U4047 (N_4047,N_3316,N_3383);
nand U4048 (N_4048,N_3607,N_3033);
and U4049 (N_4049,N_3871,N_3902);
nand U4050 (N_4050,N_3401,N_3676);
nor U4051 (N_4051,N_3113,N_3596);
nand U4052 (N_4052,N_3493,N_3453);
or U4053 (N_4053,N_3690,N_3577);
xnor U4054 (N_4054,N_3026,N_3576);
or U4055 (N_4055,N_3736,N_3619);
nand U4056 (N_4056,N_3228,N_3326);
and U4057 (N_4057,N_3471,N_3992);
or U4058 (N_4058,N_3915,N_3545);
or U4059 (N_4059,N_3748,N_3791);
or U4060 (N_4060,N_3754,N_3489);
or U4061 (N_4061,N_3536,N_3404);
nor U4062 (N_4062,N_3340,N_3437);
nor U4063 (N_4063,N_3646,N_3256);
and U4064 (N_4064,N_3456,N_3472);
nand U4065 (N_4065,N_3838,N_3629);
nand U4066 (N_4066,N_3937,N_3385);
and U4067 (N_4067,N_3013,N_3358);
or U4068 (N_4068,N_3974,N_3679);
xor U4069 (N_4069,N_3159,N_3299);
or U4070 (N_4070,N_3044,N_3626);
or U4071 (N_4071,N_3905,N_3029);
nor U4072 (N_4072,N_3080,N_3880);
and U4073 (N_4073,N_3944,N_3881);
nand U4074 (N_4074,N_3584,N_3360);
or U4075 (N_4075,N_3022,N_3262);
nand U4076 (N_4076,N_3675,N_3968);
or U4077 (N_4077,N_3090,N_3564);
nor U4078 (N_4078,N_3924,N_3290);
nor U4079 (N_4079,N_3238,N_3568);
nand U4080 (N_4080,N_3609,N_3621);
and U4081 (N_4081,N_3442,N_3796);
or U4082 (N_4082,N_3451,N_3530);
xor U4083 (N_4083,N_3491,N_3917);
or U4084 (N_4084,N_3647,N_3067);
nand U4085 (N_4085,N_3759,N_3247);
or U4086 (N_4086,N_3227,N_3126);
or U4087 (N_4087,N_3398,N_3958);
nor U4088 (N_4088,N_3426,N_3856);
and U4089 (N_4089,N_3455,N_3997);
nand U4090 (N_4090,N_3724,N_3231);
and U4091 (N_4091,N_3543,N_3563);
and U4092 (N_4092,N_3004,N_3555);
nand U4093 (N_4093,N_3207,N_3312);
nor U4094 (N_4094,N_3606,N_3274);
or U4095 (N_4095,N_3188,N_3868);
or U4096 (N_4096,N_3655,N_3494);
xor U4097 (N_4097,N_3267,N_3302);
or U4098 (N_4098,N_3192,N_3722);
and U4099 (N_4099,N_3281,N_3852);
and U4100 (N_4100,N_3125,N_3466);
and U4101 (N_4101,N_3597,N_3053);
or U4102 (N_4102,N_3191,N_3853);
nor U4103 (N_4103,N_3896,N_3972);
or U4104 (N_4104,N_3624,N_3659);
and U4105 (N_4105,N_3965,N_3264);
or U4106 (N_4106,N_3583,N_3099);
nor U4107 (N_4107,N_3272,N_3840);
nor U4108 (N_4108,N_3200,N_3497);
nand U4109 (N_4109,N_3052,N_3324);
or U4110 (N_4110,N_3356,N_3618);
nor U4111 (N_4111,N_3337,N_3071);
nor U4112 (N_4112,N_3289,N_3933);
or U4113 (N_4113,N_3925,N_3729);
or U4114 (N_4114,N_3640,N_3954);
nand U4115 (N_4115,N_3588,N_3580);
nor U4116 (N_4116,N_3402,N_3169);
or U4117 (N_4117,N_3632,N_3194);
or U4118 (N_4118,N_3458,N_3644);
or U4119 (N_4119,N_3197,N_3522);
and U4120 (N_4120,N_3161,N_3446);
nand U4121 (N_4121,N_3166,N_3391);
nor U4122 (N_4122,N_3237,N_3848);
and U4123 (N_4123,N_3677,N_3408);
nand U4124 (N_4124,N_3981,N_3135);
xnor U4125 (N_4125,N_3955,N_3149);
and U4126 (N_4126,N_3943,N_3151);
or U4127 (N_4127,N_3962,N_3064);
nand U4128 (N_4128,N_3084,N_3177);
nand U4129 (N_4129,N_3488,N_3296);
nand U4130 (N_4130,N_3480,N_3671);
nor U4131 (N_4131,N_3643,N_3167);
nand U4132 (N_4132,N_3684,N_3347);
or U4133 (N_4133,N_3328,N_3051);
nor U4134 (N_4134,N_3199,N_3323);
and U4135 (N_4135,N_3011,N_3552);
nor U4136 (N_4136,N_3622,N_3215);
nand U4137 (N_4137,N_3054,N_3836);
or U4138 (N_4138,N_3112,N_3929);
xor U4139 (N_4139,N_3062,N_3651);
nand U4140 (N_4140,N_3061,N_3799);
and U4141 (N_4141,N_3445,N_3027);
or U4142 (N_4142,N_3452,N_3219);
nor U4143 (N_4143,N_3457,N_3809);
or U4144 (N_4144,N_3932,N_3114);
or U4145 (N_4145,N_3183,N_3484);
nor U4146 (N_4146,N_3826,N_3399);
and U4147 (N_4147,N_3098,N_3270);
or U4148 (N_4148,N_3911,N_3174);
and U4149 (N_4149,N_3672,N_3198);
nand U4150 (N_4150,N_3311,N_3842);
and U4151 (N_4151,N_3030,N_3593);
or U4152 (N_4152,N_3212,N_3374);
and U4153 (N_4153,N_3845,N_3964);
nor U4154 (N_4154,N_3087,N_3823);
or U4155 (N_4155,N_3196,N_3854);
or U4156 (N_4156,N_3865,N_3146);
or U4157 (N_4157,N_3808,N_3828);
nor U4158 (N_4158,N_3470,N_3947);
or U4159 (N_4159,N_3434,N_3884);
xor U4160 (N_4160,N_3571,N_3656);
or U4161 (N_4161,N_3468,N_3635);
and U4162 (N_4162,N_3255,N_3757);
nor U4163 (N_4163,N_3591,N_3257);
nand U4164 (N_4164,N_3825,N_3774);
and U4165 (N_4165,N_3097,N_3165);
nor U4166 (N_4166,N_3031,N_3418);
nand U4167 (N_4167,N_3319,N_3710);
or U4168 (N_4168,N_3770,N_3800);
nand U4169 (N_4169,N_3859,N_3076);
nand U4170 (N_4170,N_3614,N_3831);
and U4171 (N_4171,N_3134,N_3100);
nand U4172 (N_4172,N_3393,N_3178);
nor U4173 (N_4173,N_3047,N_3473);
or U4174 (N_4174,N_3599,N_3005);
or U4175 (N_4175,N_3046,N_3738);
or U4176 (N_4176,N_3982,N_3737);
and U4177 (N_4177,N_3242,N_3221);
nand U4178 (N_4178,N_3740,N_3132);
nor U4179 (N_4179,N_3841,N_3668);
and U4180 (N_4180,N_3873,N_3887);
or U4181 (N_4181,N_3368,N_3818);
and U4182 (N_4182,N_3211,N_3006);
nand U4183 (N_4183,N_3235,N_3907);
nand U4184 (N_4184,N_3636,N_3193);
or U4185 (N_4185,N_3735,N_3674);
or U4186 (N_4186,N_3041,N_3998);
and U4187 (N_4187,N_3241,N_3540);
xor U4188 (N_4188,N_3714,N_3175);
xor U4189 (N_4189,N_3535,N_3156);
or U4190 (N_4190,N_3786,N_3295);
xnor U4191 (N_4191,N_3598,N_3077);
or U4192 (N_4192,N_3477,N_3527);
nand U4193 (N_4193,N_3948,N_3850);
nor U4194 (N_4194,N_3678,N_3699);
nand U4195 (N_4195,N_3223,N_3036);
nor U4196 (N_4196,N_3882,N_3055);
and U4197 (N_4197,N_3355,N_3345);
and U4198 (N_4198,N_3433,N_3544);
nor U4199 (N_4199,N_3155,N_3321);
nor U4200 (N_4200,N_3874,N_3127);
nor U4201 (N_4201,N_3789,N_3910);
nor U4202 (N_4202,N_3728,N_3681);
nor U4203 (N_4203,N_3578,N_3110);
xnor U4204 (N_4204,N_3481,N_3423);
nor U4205 (N_4205,N_3604,N_3978);
or U4206 (N_4206,N_3877,N_3032);
and U4207 (N_4207,N_3960,N_3285);
or U4208 (N_4208,N_3523,N_3339);
nand U4209 (N_4209,N_3260,N_3464);
and U4210 (N_4210,N_3245,N_3462);
nor U4211 (N_4211,N_3922,N_3798);
nor U4212 (N_4212,N_3993,N_3349);
nor U4213 (N_4213,N_3565,N_3008);
nor U4214 (N_4214,N_3692,N_3746);
and U4215 (N_4215,N_3269,N_3532);
nand U4216 (N_4216,N_3318,N_3507);
nand U4217 (N_4217,N_3720,N_3482);
nand U4218 (N_4218,N_3843,N_3551);
nand U4219 (N_4219,N_3454,N_3893);
and U4220 (N_4220,N_3131,N_3117);
nand U4221 (N_4221,N_3549,N_3913);
or U4222 (N_4222,N_3103,N_3204);
nand U4223 (N_4223,N_3939,N_3392);
nand U4224 (N_4224,N_3762,N_3766);
or U4225 (N_4225,N_3785,N_3400);
nor U4226 (N_4226,N_3375,N_3793);
xor U4227 (N_4227,N_3483,N_3612);
xor U4228 (N_4228,N_3298,N_3331);
nand U4229 (N_4229,N_3363,N_3524);
nand U4230 (N_4230,N_3163,N_3926);
nor U4231 (N_4231,N_3790,N_3142);
and U4232 (N_4232,N_3988,N_3560);
or U4233 (N_4233,N_3779,N_3615);
nand U4234 (N_4234,N_3633,N_3903);
or U4235 (N_4235,N_3427,N_3060);
nor U4236 (N_4236,N_3352,N_3582);
or U4237 (N_4237,N_3645,N_3554);
and U4238 (N_4238,N_3760,N_3660);
and U4239 (N_4239,N_3119,N_3348);
or U4240 (N_4240,N_3758,N_3857);
and U4241 (N_4241,N_3461,N_3743);
or U4242 (N_4242,N_3370,N_3001);
and U4243 (N_4243,N_3096,N_3176);
and U4244 (N_4244,N_3144,N_3070);
nand U4245 (N_4245,N_3058,N_3214);
or U4246 (N_4246,N_3528,N_3666);
nor U4247 (N_4247,N_3336,N_3403);
or U4248 (N_4248,N_3977,N_3875);
nand U4249 (N_4249,N_3908,N_3010);
xnor U4250 (N_4250,N_3499,N_3726);
nand U4251 (N_4251,N_3334,N_3143);
and U4252 (N_4252,N_3969,N_3009);
or U4253 (N_4253,N_3232,N_3325);
nor U4254 (N_4254,N_3899,N_3610);
or U4255 (N_4255,N_3919,N_3240);
nor U4256 (N_4256,N_3141,N_3556);
or U4257 (N_4257,N_3832,N_3755);
nand U4258 (N_4258,N_3258,N_3781);
nand U4259 (N_4259,N_3628,N_3095);
or U4260 (N_4260,N_3287,N_3670);
or U4261 (N_4261,N_3002,N_3322);
nand U4262 (N_4262,N_3007,N_3148);
xnor U4263 (N_4263,N_3202,N_3999);
nor U4264 (N_4264,N_3776,N_3485);
or U4265 (N_4265,N_3082,N_3373);
and U4266 (N_4266,N_3890,N_3686);
nand U4267 (N_4267,N_3459,N_3567);
and U4268 (N_4268,N_3927,N_3089);
nor U4269 (N_4269,N_3388,N_3572);
or U4270 (N_4270,N_3137,N_3023);
nand U4271 (N_4271,N_3696,N_3805);
and U4272 (N_4272,N_3980,N_3294);
and U4273 (N_4273,N_3815,N_3271);
or U4274 (N_4274,N_3814,N_3689);
nand U4275 (N_4275,N_3043,N_3465);
nor U4276 (N_4276,N_3763,N_3449);
and U4277 (N_4277,N_3605,N_3938);
and U4278 (N_4278,N_3384,N_3602);
xor U4279 (N_4279,N_3719,N_3557);
or U4280 (N_4280,N_3895,N_3380);
nor U4281 (N_4281,N_3467,N_3961);
xnor U4282 (N_4282,N_3120,N_3479);
nand U4283 (N_4283,N_3411,N_3486);
nand U4284 (N_4284,N_3780,N_3513);
nand U4285 (N_4285,N_3263,N_3286);
or U4286 (N_4286,N_3390,N_3844);
xnor U4287 (N_4287,N_3541,N_3833);
and U4288 (N_4288,N_3685,N_3802);
and U4289 (N_4289,N_3313,N_3806);
xnor U4290 (N_4290,N_3495,N_3105);
nand U4291 (N_4291,N_3707,N_3613);
nand U4292 (N_4292,N_3702,N_3788);
and U4293 (N_4293,N_3417,N_3885);
nor U4294 (N_4294,N_3088,N_3984);
or U4295 (N_4295,N_3303,N_3343);
nor U4296 (N_4296,N_3429,N_3000);
and U4297 (N_4297,N_3350,N_3413);
or U4298 (N_4298,N_3749,N_3600);
and U4299 (N_4299,N_3173,N_3377);
and U4300 (N_4300,N_3537,N_3509);
nor U4301 (N_4301,N_3435,N_3102);
or U4302 (N_4302,N_3079,N_3310);
nand U4303 (N_4303,N_3506,N_3139);
nor U4304 (N_4304,N_3744,N_3847);
and U4305 (N_4305,N_3548,N_3209);
or U4306 (N_4306,N_3003,N_3512);
nor U4307 (N_4307,N_3412,N_3957);
xnor U4308 (N_4308,N_3725,N_3851);
nor U4309 (N_4309,N_3152,N_3342);
and U4310 (N_4310,N_3837,N_3293);
and U4311 (N_4311,N_3371,N_3275);
xnor U4312 (N_4312,N_3276,N_3185);
and U4313 (N_4313,N_3138,N_3171);
xnor U4314 (N_4314,N_3093,N_3520);
nand U4315 (N_4315,N_3867,N_3121);
nand U4316 (N_4316,N_3996,N_3764);
nand U4317 (N_4317,N_3979,N_3226);
and U4318 (N_4318,N_3086,N_3028);
or U4319 (N_4319,N_3439,N_3233);
and U4320 (N_4320,N_3284,N_3189);
nor U4321 (N_4321,N_3057,N_3492);
and U4322 (N_4322,N_3590,N_3945);
or U4323 (N_4323,N_3346,N_3059);
nor U4324 (N_4324,N_3715,N_3048);
and U4325 (N_4325,N_3266,N_3886);
nor U4326 (N_4326,N_3519,N_3431);
and U4327 (N_4327,N_3115,N_3936);
nand U4328 (N_4328,N_3410,N_3920);
and U4329 (N_4329,N_3122,N_3731);
nand U4330 (N_4330,N_3012,N_3601);
nor U4331 (N_4331,N_3792,N_3683);
or U4332 (N_4332,N_3921,N_3991);
or U4333 (N_4333,N_3595,N_3653);
nand U4334 (N_4334,N_3250,N_3244);
nor U4335 (N_4335,N_3278,N_3111);
or U4336 (N_4336,N_3381,N_3251);
nand U4337 (N_4337,N_3585,N_3767);
xnor U4338 (N_4338,N_3118,N_3441);
and U4339 (N_4339,N_3990,N_3443);
and U4340 (N_4340,N_3634,N_3206);
nor U4341 (N_4341,N_3222,N_3918);
nand U4342 (N_4342,N_3795,N_3700);
nor U4343 (N_4343,N_3157,N_3708);
nand U4344 (N_4344,N_3382,N_3711);
nor U4345 (N_4345,N_3072,N_3168);
xor U4346 (N_4346,N_3420,N_3546);
nor U4347 (N_4347,N_3425,N_3498);
nand U4348 (N_4348,N_3288,N_3300);
xnor U4349 (N_4349,N_3306,N_3301);
nand U4350 (N_4350,N_3642,N_3305);
nand U4351 (N_4351,N_3273,N_3147);
and U4352 (N_4352,N_3804,N_3559);
nor U4353 (N_4353,N_3526,N_3989);
and U4354 (N_4354,N_3035,N_3034);
and U4355 (N_4355,N_3359,N_3050);
xor U4356 (N_4356,N_3562,N_3500);
nand U4357 (N_4357,N_3049,N_3778);
and U4358 (N_4358,N_3140,N_3765);
and U4359 (N_4359,N_3248,N_3504);
or U4360 (N_4360,N_3861,N_3773);
nor U4361 (N_4361,N_3586,N_3104);
and U4362 (N_4362,N_3732,N_3508);
and U4363 (N_4363,N_3254,N_3249);
or U4364 (N_4364,N_3930,N_3970);
nor U4365 (N_4365,N_3531,N_3956);
nand U4366 (N_4366,N_3213,N_3108);
nor U4367 (N_4367,N_3876,N_3106);
and U4368 (N_4368,N_3045,N_3320);
and U4369 (N_4369,N_3892,N_3065);
or U4370 (N_4370,N_3153,N_3372);
and U4371 (N_4371,N_3516,N_3931);
nor U4372 (N_4372,N_3953,N_3395);
nand U4373 (N_4373,N_3801,N_3389);
nand U4374 (N_4374,N_3718,N_3592);
nor U4375 (N_4375,N_3783,N_3904);
or U4376 (N_4376,N_3916,N_3218);
and U4377 (N_4377,N_3558,N_3367);
and U4378 (N_4378,N_3179,N_3745);
nor U4379 (N_4379,N_3864,N_3361);
and U4380 (N_4380,N_3150,N_3986);
or U4381 (N_4381,N_3158,N_3187);
and U4382 (N_4382,N_3641,N_3985);
nor U4383 (N_4383,N_3973,N_3474);
or U4384 (N_4384,N_3542,N_3378);
xnor U4385 (N_4385,N_3463,N_3573);
nor U4386 (N_4386,N_3888,N_3066);
nand U4387 (N_4387,N_3849,N_3243);
and U4388 (N_4388,N_3085,N_3338);
nand U4389 (N_4389,N_3771,N_3665);
nand U4390 (N_4390,N_3490,N_3693);
and U4391 (N_4391,N_3687,N_3657);
or U4392 (N_4392,N_3813,N_3704);
nor U4393 (N_4393,N_3129,N_3694);
or U4394 (N_4394,N_3335,N_3971);
nand U4395 (N_4395,N_3797,N_3824);
nor U4396 (N_4396,N_3811,N_3252);
nor U4397 (N_4397,N_3631,N_3891);
and U4398 (N_4398,N_3701,N_3807);
or U4399 (N_4399,N_3341,N_3638);
nand U4400 (N_4400,N_3422,N_3063);
nand U4401 (N_4401,N_3579,N_3332);
nor U4402 (N_4402,N_3405,N_3663);
xnor U4403 (N_4403,N_3821,N_3184);
nand U4404 (N_4404,N_3975,N_3935);
nand U4405 (N_4405,N_3021,N_3934);
and U4406 (N_4406,N_3630,N_3611);
and U4407 (N_4407,N_3817,N_3872);
nor U4408 (N_4408,N_3662,N_3107);
nand U4409 (N_4409,N_3810,N_3447);
or U4410 (N_4410,N_3503,N_3756);
nor U4411 (N_4411,N_3750,N_3414);
nand U4412 (N_4412,N_3862,N_3730);
or U4413 (N_4413,N_3366,N_3476);
and U4414 (N_4414,N_3230,N_3136);
nor U4415 (N_4415,N_3858,N_3075);
or U4416 (N_4416,N_3353,N_3855);
and U4417 (N_4417,N_3224,N_3501);
and U4418 (N_4418,N_3816,N_3469);
and U4419 (N_4419,N_3712,N_3386);
or U4420 (N_4420,N_3496,N_3421);
nor U4421 (N_4421,N_3717,N_3037);
xnor U4422 (N_4422,N_3553,N_3160);
and U4423 (N_4423,N_3292,N_3952);
nand U4424 (N_4424,N_3083,N_3761);
nand U4425 (N_4425,N_3667,N_3018);
nand U4426 (N_4426,N_3123,N_3963);
nand U4427 (N_4427,N_3432,N_3379);
nor U4428 (N_4428,N_3024,N_3521);
nand U4429 (N_4429,N_3518,N_3253);
xor U4430 (N_4430,N_3201,N_3747);
nor U4431 (N_4431,N_3594,N_3966);
xor U4432 (N_4432,N_3020,N_3220);
nand U4433 (N_4433,N_3517,N_3424);
nand U4434 (N_4434,N_3068,N_3787);
and U4435 (N_4435,N_3124,N_3673);
nand U4436 (N_4436,N_3533,N_3561);
nand U4437 (N_4437,N_3450,N_3019);
or U4438 (N_4438,N_3987,N_3829);
and U4439 (N_4439,N_3056,N_3069);
nor U4440 (N_4440,N_3128,N_3547);
nand U4441 (N_4441,N_3900,N_3706);
or U4442 (N_4442,N_3344,N_3236);
nand U4443 (N_4443,N_3940,N_3025);
nor U4444 (N_4444,N_3839,N_3376);
or U4445 (N_4445,N_3180,N_3282);
or U4446 (N_4446,N_3162,N_3883);
or U4447 (N_4447,N_3777,N_3909);
or U4448 (N_4448,N_3092,N_3487);
and U4449 (N_4449,N_3705,N_3733);
nand U4450 (N_4450,N_3440,N_3304);
and U4451 (N_4451,N_3616,N_3682);
or U4452 (N_4452,N_3534,N_3637);
or U4453 (N_4453,N_3751,N_3073);
or U4454 (N_4454,N_3574,N_3307);
and U4455 (N_4455,N_3394,N_3794);
nand U4456 (N_4456,N_3942,N_3291);
or U4457 (N_4457,N_3654,N_3154);
xor U4458 (N_4458,N_3186,N_3538);
nand U4459 (N_4459,N_3941,N_3739);
nor U4460 (N_4460,N_3297,N_3620);
and U4461 (N_4461,N_3627,N_3566);
or U4462 (N_4462,N_3742,N_3639);
nand U4463 (N_4463,N_3280,N_3669);
or U4464 (N_4464,N_3116,N_3650);
or U4465 (N_4465,N_3396,N_3014);
nor U4466 (N_4466,N_3623,N_3995);
or U4467 (N_4467,N_3914,N_3460);
nor U4468 (N_4468,N_3406,N_3946);
nor U4469 (N_4469,N_3015,N_3603);
nor U4470 (N_4470,N_3038,N_3860);
nand U4471 (N_4471,N_3333,N_3514);
nand U4472 (N_4472,N_3550,N_3101);
nand U4473 (N_4473,N_3094,N_3217);
nor U4474 (N_4474,N_3752,N_3819);
nor U4475 (N_4475,N_3172,N_3688);
nor U4476 (N_4476,N_3515,N_3415);
and U4477 (N_4477,N_3784,N_3362);
and U4478 (N_4478,N_3216,N_3769);
or U4479 (N_4479,N_3225,N_3407);
or U4480 (N_4480,N_3912,N_3661);
or U4481 (N_4481,N_3906,N_3866);
nor U4482 (N_4482,N_3145,N_3327);
nand U4483 (N_4483,N_3208,N_3587);
and U4484 (N_4484,N_3164,N_3901);
nor U4485 (N_4485,N_3695,N_3680);
or U4486 (N_4486,N_3608,N_3658);
nor U4487 (N_4487,N_3983,N_3529);
and U4488 (N_4488,N_3365,N_3315);
nor U4489 (N_4489,N_3511,N_3713);
nor U4490 (N_4490,N_3448,N_3869);
nor U4491 (N_4491,N_3649,N_3478);
or U4492 (N_4492,N_3246,N_3239);
nor U4493 (N_4493,N_3017,N_3279);
nor U4494 (N_4494,N_3863,N_3753);
and U4495 (N_4495,N_3133,N_3042);
nor U4496 (N_4496,N_3040,N_3317);
and U4497 (N_4497,N_3039,N_3716);
nor U4498 (N_4498,N_3870,N_3691);
or U4499 (N_4499,N_3812,N_3539);
or U4500 (N_4500,N_3552,N_3550);
or U4501 (N_4501,N_3869,N_3692);
nor U4502 (N_4502,N_3387,N_3271);
and U4503 (N_4503,N_3693,N_3782);
nor U4504 (N_4504,N_3720,N_3032);
and U4505 (N_4505,N_3388,N_3104);
and U4506 (N_4506,N_3085,N_3611);
nand U4507 (N_4507,N_3065,N_3299);
or U4508 (N_4508,N_3651,N_3733);
or U4509 (N_4509,N_3271,N_3978);
and U4510 (N_4510,N_3917,N_3576);
nand U4511 (N_4511,N_3301,N_3110);
nor U4512 (N_4512,N_3242,N_3902);
xor U4513 (N_4513,N_3289,N_3613);
xnor U4514 (N_4514,N_3252,N_3500);
or U4515 (N_4515,N_3813,N_3565);
nand U4516 (N_4516,N_3890,N_3156);
and U4517 (N_4517,N_3516,N_3987);
or U4518 (N_4518,N_3439,N_3624);
nor U4519 (N_4519,N_3658,N_3642);
and U4520 (N_4520,N_3910,N_3786);
and U4521 (N_4521,N_3144,N_3185);
nand U4522 (N_4522,N_3578,N_3118);
nand U4523 (N_4523,N_3475,N_3294);
nand U4524 (N_4524,N_3483,N_3087);
and U4525 (N_4525,N_3898,N_3984);
or U4526 (N_4526,N_3100,N_3620);
nor U4527 (N_4527,N_3404,N_3590);
xnor U4528 (N_4528,N_3270,N_3682);
or U4529 (N_4529,N_3685,N_3927);
or U4530 (N_4530,N_3119,N_3471);
nor U4531 (N_4531,N_3073,N_3716);
nand U4532 (N_4532,N_3673,N_3485);
nor U4533 (N_4533,N_3310,N_3505);
nor U4534 (N_4534,N_3018,N_3709);
nand U4535 (N_4535,N_3700,N_3133);
and U4536 (N_4536,N_3946,N_3693);
nor U4537 (N_4537,N_3840,N_3058);
and U4538 (N_4538,N_3669,N_3413);
nand U4539 (N_4539,N_3467,N_3421);
nor U4540 (N_4540,N_3796,N_3076);
nor U4541 (N_4541,N_3296,N_3400);
nor U4542 (N_4542,N_3187,N_3229);
and U4543 (N_4543,N_3218,N_3067);
nor U4544 (N_4544,N_3477,N_3597);
nand U4545 (N_4545,N_3236,N_3738);
or U4546 (N_4546,N_3366,N_3406);
and U4547 (N_4547,N_3495,N_3451);
or U4548 (N_4548,N_3697,N_3611);
and U4549 (N_4549,N_3201,N_3777);
nand U4550 (N_4550,N_3395,N_3643);
nor U4551 (N_4551,N_3577,N_3246);
or U4552 (N_4552,N_3998,N_3686);
and U4553 (N_4553,N_3540,N_3909);
nor U4554 (N_4554,N_3712,N_3877);
and U4555 (N_4555,N_3187,N_3914);
nor U4556 (N_4556,N_3719,N_3680);
and U4557 (N_4557,N_3919,N_3780);
nor U4558 (N_4558,N_3174,N_3478);
or U4559 (N_4559,N_3372,N_3414);
and U4560 (N_4560,N_3026,N_3960);
or U4561 (N_4561,N_3261,N_3669);
or U4562 (N_4562,N_3395,N_3308);
nand U4563 (N_4563,N_3729,N_3446);
or U4564 (N_4564,N_3796,N_3727);
nor U4565 (N_4565,N_3166,N_3922);
and U4566 (N_4566,N_3169,N_3552);
nor U4567 (N_4567,N_3034,N_3324);
nor U4568 (N_4568,N_3493,N_3347);
nor U4569 (N_4569,N_3002,N_3595);
and U4570 (N_4570,N_3691,N_3593);
and U4571 (N_4571,N_3439,N_3342);
xnor U4572 (N_4572,N_3557,N_3776);
xor U4573 (N_4573,N_3218,N_3154);
nor U4574 (N_4574,N_3448,N_3552);
nand U4575 (N_4575,N_3609,N_3089);
nor U4576 (N_4576,N_3596,N_3388);
and U4577 (N_4577,N_3459,N_3727);
xnor U4578 (N_4578,N_3457,N_3040);
or U4579 (N_4579,N_3806,N_3740);
and U4580 (N_4580,N_3060,N_3517);
and U4581 (N_4581,N_3522,N_3217);
nor U4582 (N_4582,N_3920,N_3737);
nand U4583 (N_4583,N_3698,N_3969);
nand U4584 (N_4584,N_3542,N_3596);
and U4585 (N_4585,N_3990,N_3117);
nor U4586 (N_4586,N_3806,N_3146);
nor U4587 (N_4587,N_3975,N_3149);
and U4588 (N_4588,N_3202,N_3939);
and U4589 (N_4589,N_3421,N_3826);
and U4590 (N_4590,N_3950,N_3139);
nand U4591 (N_4591,N_3400,N_3147);
and U4592 (N_4592,N_3625,N_3856);
or U4593 (N_4593,N_3449,N_3358);
and U4594 (N_4594,N_3054,N_3486);
or U4595 (N_4595,N_3950,N_3213);
nor U4596 (N_4596,N_3158,N_3105);
and U4597 (N_4597,N_3711,N_3936);
and U4598 (N_4598,N_3102,N_3084);
or U4599 (N_4599,N_3294,N_3257);
nor U4600 (N_4600,N_3241,N_3136);
and U4601 (N_4601,N_3895,N_3056);
nand U4602 (N_4602,N_3058,N_3308);
nor U4603 (N_4603,N_3641,N_3663);
nand U4604 (N_4604,N_3110,N_3488);
or U4605 (N_4605,N_3209,N_3056);
nor U4606 (N_4606,N_3061,N_3090);
nand U4607 (N_4607,N_3472,N_3019);
or U4608 (N_4608,N_3332,N_3839);
or U4609 (N_4609,N_3637,N_3071);
nand U4610 (N_4610,N_3144,N_3624);
nand U4611 (N_4611,N_3139,N_3345);
nor U4612 (N_4612,N_3735,N_3064);
and U4613 (N_4613,N_3524,N_3130);
nand U4614 (N_4614,N_3773,N_3781);
nand U4615 (N_4615,N_3968,N_3599);
nand U4616 (N_4616,N_3994,N_3280);
and U4617 (N_4617,N_3403,N_3463);
nor U4618 (N_4618,N_3448,N_3473);
or U4619 (N_4619,N_3392,N_3467);
nand U4620 (N_4620,N_3364,N_3852);
and U4621 (N_4621,N_3899,N_3513);
nor U4622 (N_4622,N_3819,N_3076);
or U4623 (N_4623,N_3029,N_3714);
or U4624 (N_4624,N_3705,N_3513);
or U4625 (N_4625,N_3331,N_3212);
and U4626 (N_4626,N_3535,N_3077);
nand U4627 (N_4627,N_3879,N_3771);
or U4628 (N_4628,N_3111,N_3958);
nand U4629 (N_4629,N_3409,N_3928);
and U4630 (N_4630,N_3973,N_3220);
or U4631 (N_4631,N_3829,N_3652);
xnor U4632 (N_4632,N_3541,N_3714);
and U4633 (N_4633,N_3794,N_3196);
nor U4634 (N_4634,N_3641,N_3794);
nor U4635 (N_4635,N_3982,N_3641);
xnor U4636 (N_4636,N_3415,N_3221);
and U4637 (N_4637,N_3439,N_3737);
nand U4638 (N_4638,N_3556,N_3970);
nand U4639 (N_4639,N_3654,N_3367);
and U4640 (N_4640,N_3691,N_3386);
or U4641 (N_4641,N_3426,N_3063);
nand U4642 (N_4642,N_3401,N_3855);
or U4643 (N_4643,N_3320,N_3807);
nand U4644 (N_4644,N_3227,N_3105);
or U4645 (N_4645,N_3518,N_3091);
nor U4646 (N_4646,N_3758,N_3362);
or U4647 (N_4647,N_3187,N_3493);
or U4648 (N_4648,N_3659,N_3781);
or U4649 (N_4649,N_3117,N_3301);
nor U4650 (N_4650,N_3407,N_3640);
nand U4651 (N_4651,N_3131,N_3823);
nor U4652 (N_4652,N_3325,N_3908);
nor U4653 (N_4653,N_3909,N_3422);
xnor U4654 (N_4654,N_3614,N_3348);
and U4655 (N_4655,N_3241,N_3445);
or U4656 (N_4656,N_3109,N_3725);
or U4657 (N_4657,N_3364,N_3549);
nor U4658 (N_4658,N_3800,N_3809);
nor U4659 (N_4659,N_3411,N_3315);
nor U4660 (N_4660,N_3060,N_3014);
and U4661 (N_4661,N_3859,N_3083);
and U4662 (N_4662,N_3625,N_3854);
nand U4663 (N_4663,N_3297,N_3862);
nor U4664 (N_4664,N_3731,N_3840);
nor U4665 (N_4665,N_3193,N_3652);
and U4666 (N_4666,N_3573,N_3939);
and U4667 (N_4667,N_3359,N_3961);
and U4668 (N_4668,N_3648,N_3409);
or U4669 (N_4669,N_3275,N_3613);
nand U4670 (N_4670,N_3707,N_3103);
nor U4671 (N_4671,N_3887,N_3403);
nand U4672 (N_4672,N_3391,N_3898);
nand U4673 (N_4673,N_3431,N_3953);
or U4674 (N_4674,N_3082,N_3207);
xor U4675 (N_4675,N_3050,N_3918);
or U4676 (N_4676,N_3142,N_3369);
and U4677 (N_4677,N_3197,N_3956);
nor U4678 (N_4678,N_3856,N_3265);
nand U4679 (N_4679,N_3224,N_3899);
and U4680 (N_4680,N_3611,N_3200);
nand U4681 (N_4681,N_3761,N_3635);
or U4682 (N_4682,N_3841,N_3580);
nand U4683 (N_4683,N_3167,N_3477);
nor U4684 (N_4684,N_3747,N_3089);
or U4685 (N_4685,N_3090,N_3583);
nand U4686 (N_4686,N_3368,N_3006);
or U4687 (N_4687,N_3975,N_3703);
or U4688 (N_4688,N_3240,N_3389);
and U4689 (N_4689,N_3744,N_3227);
and U4690 (N_4690,N_3991,N_3414);
nor U4691 (N_4691,N_3413,N_3440);
or U4692 (N_4692,N_3387,N_3418);
nor U4693 (N_4693,N_3899,N_3897);
or U4694 (N_4694,N_3360,N_3820);
nand U4695 (N_4695,N_3411,N_3439);
or U4696 (N_4696,N_3301,N_3826);
xor U4697 (N_4697,N_3088,N_3278);
nand U4698 (N_4698,N_3778,N_3712);
nor U4699 (N_4699,N_3549,N_3977);
nor U4700 (N_4700,N_3478,N_3818);
nor U4701 (N_4701,N_3333,N_3881);
nor U4702 (N_4702,N_3099,N_3247);
or U4703 (N_4703,N_3731,N_3075);
and U4704 (N_4704,N_3634,N_3083);
nand U4705 (N_4705,N_3776,N_3872);
xor U4706 (N_4706,N_3725,N_3025);
or U4707 (N_4707,N_3534,N_3574);
nor U4708 (N_4708,N_3576,N_3117);
or U4709 (N_4709,N_3108,N_3837);
or U4710 (N_4710,N_3213,N_3093);
nand U4711 (N_4711,N_3026,N_3676);
nand U4712 (N_4712,N_3833,N_3816);
and U4713 (N_4713,N_3217,N_3916);
xor U4714 (N_4714,N_3628,N_3291);
or U4715 (N_4715,N_3666,N_3697);
nor U4716 (N_4716,N_3121,N_3492);
nor U4717 (N_4717,N_3306,N_3369);
nor U4718 (N_4718,N_3460,N_3173);
nor U4719 (N_4719,N_3941,N_3300);
nand U4720 (N_4720,N_3265,N_3909);
nor U4721 (N_4721,N_3443,N_3505);
xnor U4722 (N_4722,N_3481,N_3633);
and U4723 (N_4723,N_3699,N_3152);
xnor U4724 (N_4724,N_3377,N_3533);
or U4725 (N_4725,N_3239,N_3009);
nand U4726 (N_4726,N_3754,N_3926);
nor U4727 (N_4727,N_3389,N_3743);
and U4728 (N_4728,N_3871,N_3593);
nand U4729 (N_4729,N_3437,N_3989);
nand U4730 (N_4730,N_3803,N_3906);
or U4731 (N_4731,N_3800,N_3719);
nand U4732 (N_4732,N_3044,N_3775);
nand U4733 (N_4733,N_3988,N_3921);
nand U4734 (N_4734,N_3803,N_3668);
and U4735 (N_4735,N_3406,N_3556);
nor U4736 (N_4736,N_3584,N_3125);
and U4737 (N_4737,N_3725,N_3243);
nand U4738 (N_4738,N_3741,N_3458);
and U4739 (N_4739,N_3426,N_3011);
nor U4740 (N_4740,N_3157,N_3799);
and U4741 (N_4741,N_3119,N_3892);
nor U4742 (N_4742,N_3427,N_3288);
nor U4743 (N_4743,N_3500,N_3490);
or U4744 (N_4744,N_3350,N_3242);
nand U4745 (N_4745,N_3989,N_3420);
and U4746 (N_4746,N_3232,N_3249);
and U4747 (N_4747,N_3866,N_3918);
xor U4748 (N_4748,N_3256,N_3995);
and U4749 (N_4749,N_3339,N_3958);
and U4750 (N_4750,N_3590,N_3569);
nor U4751 (N_4751,N_3021,N_3040);
nor U4752 (N_4752,N_3151,N_3846);
xor U4753 (N_4753,N_3599,N_3853);
nand U4754 (N_4754,N_3536,N_3853);
and U4755 (N_4755,N_3034,N_3819);
nand U4756 (N_4756,N_3891,N_3388);
or U4757 (N_4757,N_3939,N_3556);
and U4758 (N_4758,N_3825,N_3213);
nand U4759 (N_4759,N_3381,N_3153);
and U4760 (N_4760,N_3400,N_3619);
nor U4761 (N_4761,N_3329,N_3205);
nor U4762 (N_4762,N_3357,N_3991);
nand U4763 (N_4763,N_3274,N_3271);
nand U4764 (N_4764,N_3569,N_3646);
nor U4765 (N_4765,N_3241,N_3791);
nand U4766 (N_4766,N_3296,N_3475);
or U4767 (N_4767,N_3642,N_3120);
nand U4768 (N_4768,N_3243,N_3103);
nor U4769 (N_4769,N_3385,N_3316);
xor U4770 (N_4770,N_3951,N_3116);
and U4771 (N_4771,N_3256,N_3749);
nor U4772 (N_4772,N_3483,N_3842);
nor U4773 (N_4773,N_3522,N_3450);
nor U4774 (N_4774,N_3722,N_3956);
xnor U4775 (N_4775,N_3767,N_3748);
xnor U4776 (N_4776,N_3670,N_3488);
or U4777 (N_4777,N_3185,N_3389);
or U4778 (N_4778,N_3911,N_3695);
and U4779 (N_4779,N_3567,N_3748);
nor U4780 (N_4780,N_3306,N_3577);
nand U4781 (N_4781,N_3381,N_3757);
or U4782 (N_4782,N_3440,N_3723);
nand U4783 (N_4783,N_3707,N_3175);
and U4784 (N_4784,N_3530,N_3491);
nand U4785 (N_4785,N_3111,N_3493);
nand U4786 (N_4786,N_3132,N_3471);
xnor U4787 (N_4787,N_3947,N_3993);
and U4788 (N_4788,N_3305,N_3395);
and U4789 (N_4789,N_3188,N_3297);
or U4790 (N_4790,N_3566,N_3973);
or U4791 (N_4791,N_3083,N_3691);
nor U4792 (N_4792,N_3530,N_3105);
or U4793 (N_4793,N_3411,N_3715);
nand U4794 (N_4794,N_3909,N_3009);
and U4795 (N_4795,N_3608,N_3304);
or U4796 (N_4796,N_3267,N_3816);
or U4797 (N_4797,N_3859,N_3149);
nor U4798 (N_4798,N_3648,N_3346);
nor U4799 (N_4799,N_3733,N_3473);
nor U4800 (N_4800,N_3244,N_3368);
xor U4801 (N_4801,N_3737,N_3482);
and U4802 (N_4802,N_3647,N_3283);
nor U4803 (N_4803,N_3743,N_3408);
nor U4804 (N_4804,N_3516,N_3582);
nor U4805 (N_4805,N_3022,N_3101);
nand U4806 (N_4806,N_3852,N_3845);
nor U4807 (N_4807,N_3608,N_3165);
nand U4808 (N_4808,N_3484,N_3988);
xor U4809 (N_4809,N_3332,N_3428);
and U4810 (N_4810,N_3011,N_3448);
nand U4811 (N_4811,N_3707,N_3898);
nor U4812 (N_4812,N_3505,N_3806);
xor U4813 (N_4813,N_3994,N_3139);
and U4814 (N_4814,N_3014,N_3370);
nand U4815 (N_4815,N_3701,N_3653);
nor U4816 (N_4816,N_3806,N_3656);
and U4817 (N_4817,N_3008,N_3182);
nor U4818 (N_4818,N_3795,N_3901);
or U4819 (N_4819,N_3450,N_3233);
nand U4820 (N_4820,N_3152,N_3542);
and U4821 (N_4821,N_3882,N_3630);
and U4822 (N_4822,N_3959,N_3366);
or U4823 (N_4823,N_3926,N_3579);
and U4824 (N_4824,N_3814,N_3373);
and U4825 (N_4825,N_3088,N_3683);
nand U4826 (N_4826,N_3966,N_3044);
or U4827 (N_4827,N_3692,N_3676);
or U4828 (N_4828,N_3745,N_3800);
nand U4829 (N_4829,N_3555,N_3250);
nor U4830 (N_4830,N_3703,N_3466);
nor U4831 (N_4831,N_3929,N_3751);
xnor U4832 (N_4832,N_3068,N_3044);
nand U4833 (N_4833,N_3257,N_3848);
nand U4834 (N_4834,N_3246,N_3690);
nand U4835 (N_4835,N_3202,N_3394);
or U4836 (N_4836,N_3064,N_3073);
and U4837 (N_4837,N_3738,N_3803);
and U4838 (N_4838,N_3571,N_3200);
nor U4839 (N_4839,N_3779,N_3645);
or U4840 (N_4840,N_3973,N_3843);
or U4841 (N_4841,N_3183,N_3567);
nand U4842 (N_4842,N_3753,N_3026);
or U4843 (N_4843,N_3190,N_3473);
or U4844 (N_4844,N_3401,N_3980);
xor U4845 (N_4845,N_3571,N_3103);
nand U4846 (N_4846,N_3443,N_3904);
nor U4847 (N_4847,N_3736,N_3578);
nand U4848 (N_4848,N_3051,N_3463);
and U4849 (N_4849,N_3994,N_3022);
nor U4850 (N_4850,N_3246,N_3066);
xor U4851 (N_4851,N_3139,N_3036);
nor U4852 (N_4852,N_3503,N_3525);
or U4853 (N_4853,N_3983,N_3032);
or U4854 (N_4854,N_3303,N_3270);
xor U4855 (N_4855,N_3886,N_3098);
xnor U4856 (N_4856,N_3958,N_3163);
nor U4857 (N_4857,N_3676,N_3441);
nor U4858 (N_4858,N_3609,N_3883);
xor U4859 (N_4859,N_3850,N_3076);
xor U4860 (N_4860,N_3139,N_3136);
or U4861 (N_4861,N_3127,N_3483);
nand U4862 (N_4862,N_3157,N_3401);
nand U4863 (N_4863,N_3793,N_3237);
or U4864 (N_4864,N_3810,N_3943);
nand U4865 (N_4865,N_3465,N_3254);
or U4866 (N_4866,N_3153,N_3802);
xnor U4867 (N_4867,N_3867,N_3327);
and U4868 (N_4868,N_3473,N_3895);
nand U4869 (N_4869,N_3026,N_3352);
or U4870 (N_4870,N_3667,N_3184);
and U4871 (N_4871,N_3818,N_3675);
or U4872 (N_4872,N_3133,N_3851);
and U4873 (N_4873,N_3809,N_3006);
xnor U4874 (N_4874,N_3434,N_3433);
xnor U4875 (N_4875,N_3980,N_3777);
and U4876 (N_4876,N_3936,N_3873);
and U4877 (N_4877,N_3854,N_3866);
or U4878 (N_4878,N_3252,N_3869);
nor U4879 (N_4879,N_3153,N_3271);
and U4880 (N_4880,N_3213,N_3568);
and U4881 (N_4881,N_3679,N_3580);
and U4882 (N_4882,N_3975,N_3253);
nand U4883 (N_4883,N_3778,N_3518);
nor U4884 (N_4884,N_3037,N_3298);
or U4885 (N_4885,N_3234,N_3389);
nor U4886 (N_4886,N_3778,N_3628);
and U4887 (N_4887,N_3296,N_3793);
or U4888 (N_4888,N_3556,N_3202);
xnor U4889 (N_4889,N_3136,N_3332);
nand U4890 (N_4890,N_3401,N_3885);
nand U4891 (N_4891,N_3297,N_3755);
or U4892 (N_4892,N_3381,N_3431);
nor U4893 (N_4893,N_3205,N_3917);
nand U4894 (N_4894,N_3785,N_3329);
and U4895 (N_4895,N_3866,N_3585);
nor U4896 (N_4896,N_3049,N_3123);
nor U4897 (N_4897,N_3979,N_3192);
or U4898 (N_4898,N_3703,N_3261);
or U4899 (N_4899,N_3744,N_3397);
nor U4900 (N_4900,N_3512,N_3724);
nand U4901 (N_4901,N_3354,N_3811);
nand U4902 (N_4902,N_3557,N_3715);
nor U4903 (N_4903,N_3800,N_3374);
nor U4904 (N_4904,N_3076,N_3965);
nor U4905 (N_4905,N_3719,N_3214);
xor U4906 (N_4906,N_3266,N_3388);
and U4907 (N_4907,N_3642,N_3783);
or U4908 (N_4908,N_3249,N_3542);
nand U4909 (N_4909,N_3651,N_3832);
or U4910 (N_4910,N_3351,N_3782);
nor U4911 (N_4911,N_3065,N_3696);
nand U4912 (N_4912,N_3589,N_3675);
nor U4913 (N_4913,N_3398,N_3021);
nor U4914 (N_4914,N_3814,N_3538);
or U4915 (N_4915,N_3496,N_3381);
xnor U4916 (N_4916,N_3184,N_3576);
xor U4917 (N_4917,N_3781,N_3018);
nand U4918 (N_4918,N_3433,N_3376);
and U4919 (N_4919,N_3454,N_3265);
nand U4920 (N_4920,N_3276,N_3946);
nor U4921 (N_4921,N_3989,N_3967);
xor U4922 (N_4922,N_3063,N_3638);
nor U4923 (N_4923,N_3905,N_3141);
or U4924 (N_4924,N_3809,N_3526);
or U4925 (N_4925,N_3740,N_3920);
xnor U4926 (N_4926,N_3975,N_3171);
xnor U4927 (N_4927,N_3182,N_3702);
and U4928 (N_4928,N_3626,N_3414);
nand U4929 (N_4929,N_3806,N_3729);
or U4930 (N_4930,N_3736,N_3858);
nor U4931 (N_4931,N_3038,N_3333);
or U4932 (N_4932,N_3969,N_3905);
nor U4933 (N_4933,N_3276,N_3022);
nand U4934 (N_4934,N_3216,N_3997);
nor U4935 (N_4935,N_3587,N_3282);
and U4936 (N_4936,N_3058,N_3426);
nor U4937 (N_4937,N_3357,N_3870);
and U4938 (N_4938,N_3321,N_3301);
and U4939 (N_4939,N_3081,N_3565);
nor U4940 (N_4940,N_3660,N_3181);
nor U4941 (N_4941,N_3420,N_3515);
nand U4942 (N_4942,N_3082,N_3938);
and U4943 (N_4943,N_3736,N_3526);
nor U4944 (N_4944,N_3297,N_3498);
or U4945 (N_4945,N_3950,N_3120);
nand U4946 (N_4946,N_3345,N_3839);
nor U4947 (N_4947,N_3708,N_3377);
and U4948 (N_4948,N_3886,N_3079);
or U4949 (N_4949,N_3385,N_3988);
nor U4950 (N_4950,N_3045,N_3924);
or U4951 (N_4951,N_3419,N_3386);
and U4952 (N_4952,N_3355,N_3919);
nand U4953 (N_4953,N_3962,N_3830);
and U4954 (N_4954,N_3016,N_3922);
xnor U4955 (N_4955,N_3388,N_3771);
nor U4956 (N_4956,N_3843,N_3906);
nand U4957 (N_4957,N_3458,N_3253);
nand U4958 (N_4958,N_3462,N_3120);
nand U4959 (N_4959,N_3862,N_3405);
nor U4960 (N_4960,N_3154,N_3447);
nand U4961 (N_4961,N_3649,N_3704);
or U4962 (N_4962,N_3776,N_3636);
nor U4963 (N_4963,N_3019,N_3770);
and U4964 (N_4964,N_3317,N_3362);
nand U4965 (N_4965,N_3011,N_3056);
and U4966 (N_4966,N_3633,N_3727);
xnor U4967 (N_4967,N_3628,N_3228);
nor U4968 (N_4968,N_3397,N_3161);
or U4969 (N_4969,N_3210,N_3479);
and U4970 (N_4970,N_3364,N_3824);
nand U4971 (N_4971,N_3555,N_3328);
xnor U4972 (N_4972,N_3466,N_3917);
and U4973 (N_4973,N_3978,N_3997);
nand U4974 (N_4974,N_3477,N_3751);
or U4975 (N_4975,N_3912,N_3987);
and U4976 (N_4976,N_3277,N_3892);
and U4977 (N_4977,N_3771,N_3004);
and U4978 (N_4978,N_3557,N_3968);
or U4979 (N_4979,N_3127,N_3315);
nor U4980 (N_4980,N_3024,N_3078);
xor U4981 (N_4981,N_3063,N_3162);
nand U4982 (N_4982,N_3738,N_3734);
nor U4983 (N_4983,N_3794,N_3652);
nand U4984 (N_4984,N_3580,N_3199);
xnor U4985 (N_4985,N_3157,N_3874);
and U4986 (N_4986,N_3485,N_3413);
or U4987 (N_4987,N_3474,N_3927);
and U4988 (N_4988,N_3009,N_3588);
or U4989 (N_4989,N_3810,N_3260);
nand U4990 (N_4990,N_3262,N_3302);
xnor U4991 (N_4991,N_3959,N_3129);
and U4992 (N_4992,N_3244,N_3712);
nand U4993 (N_4993,N_3066,N_3813);
or U4994 (N_4994,N_3369,N_3347);
nand U4995 (N_4995,N_3733,N_3203);
or U4996 (N_4996,N_3300,N_3155);
nand U4997 (N_4997,N_3324,N_3863);
and U4998 (N_4998,N_3635,N_3120);
and U4999 (N_4999,N_3128,N_3388);
or U5000 (N_5000,N_4339,N_4857);
xor U5001 (N_5001,N_4297,N_4400);
nor U5002 (N_5002,N_4625,N_4072);
nand U5003 (N_5003,N_4269,N_4337);
and U5004 (N_5004,N_4418,N_4587);
or U5005 (N_5005,N_4827,N_4138);
nand U5006 (N_5006,N_4494,N_4540);
nor U5007 (N_5007,N_4941,N_4755);
nand U5008 (N_5008,N_4955,N_4136);
and U5009 (N_5009,N_4772,N_4325);
nor U5010 (N_5010,N_4626,N_4383);
and U5011 (N_5011,N_4988,N_4863);
nand U5012 (N_5012,N_4791,N_4491);
and U5013 (N_5013,N_4807,N_4855);
and U5014 (N_5014,N_4679,N_4966);
and U5015 (N_5015,N_4630,N_4634);
or U5016 (N_5016,N_4476,N_4263);
nor U5017 (N_5017,N_4194,N_4907);
nand U5018 (N_5018,N_4454,N_4799);
nand U5019 (N_5019,N_4188,N_4474);
nor U5020 (N_5020,N_4356,N_4722);
nor U5021 (N_5021,N_4856,N_4990);
nor U5022 (N_5022,N_4522,N_4889);
nor U5023 (N_5023,N_4153,N_4227);
nor U5024 (N_5024,N_4007,N_4960);
nor U5025 (N_5025,N_4437,N_4352);
xor U5026 (N_5026,N_4436,N_4228);
nor U5027 (N_5027,N_4224,N_4719);
nor U5028 (N_5028,N_4659,N_4554);
nor U5029 (N_5029,N_4117,N_4578);
and U5030 (N_5030,N_4528,N_4979);
nor U5031 (N_5031,N_4078,N_4651);
and U5032 (N_5032,N_4694,N_4756);
xnor U5033 (N_5033,N_4585,N_4823);
and U5034 (N_5034,N_4940,N_4777);
or U5035 (N_5035,N_4477,N_4861);
nor U5036 (N_5036,N_4558,N_4850);
or U5037 (N_5037,N_4134,N_4318);
xnor U5038 (N_5038,N_4408,N_4283);
nor U5039 (N_5039,N_4206,N_4902);
nor U5040 (N_5040,N_4100,N_4164);
and U5041 (N_5041,N_4716,N_4853);
and U5042 (N_5042,N_4743,N_4961);
nand U5043 (N_5043,N_4820,N_4598);
and U5044 (N_5044,N_4232,N_4407);
and U5045 (N_5045,N_4537,N_4236);
or U5046 (N_5046,N_4552,N_4358);
nand U5047 (N_5047,N_4316,N_4958);
or U5048 (N_5048,N_4333,N_4879);
nor U5049 (N_5049,N_4700,N_4049);
and U5050 (N_5050,N_4524,N_4357);
xor U5051 (N_5051,N_4299,N_4306);
or U5052 (N_5052,N_4565,N_4945);
or U5053 (N_5053,N_4124,N_4122);
and U5054 (N_5054,N_4146,N_4214);
nor U5055 (N_5055,N_4709,N_4096);
nor U5056 (N_5056,N_4387,N_4233);
nor U5057 (N_5057,N_4635,N_4847);
nor U5058 (N_5058,N_4697,N_4390);
nand U5059 (N_5059,N_4413,N_4562);
nor U5060 (N_5060,N_4180,N_4652);
and U5061 (N_5061,N_4597,N_4244);
nor U5062 (N_5062,N_4076,N_4074);
or U5063 (N_5063,N_4954,N_4790);
and U5064 (N_5064,N_4584,N_4415);
nor U5065 (N_5065,N_4456,N_4040);
nand U5066 (N_5066,N_4484,N_4069);
or U5067 (N_5067,N_4929,N_4726);
or U5068 (N_5068,N_4167,N_4329);
and U5069 (N_5069,N_4278,N_4953);
nor U5070 (N_5070,N_4090,N_4720);
nand U5071 (N_5071,N_4057,N_4257);
nand U5072 (N_5072,N_4241,N_4615);
nor U5073 (N_5073,N_4810,N_4775);
nor U5074 (N_5074,N_4774,N_4691);
and U5075 (N_5075,N_4821,N_4669);
xor U5076 (N_5076,N_4922,N_4721);
nor U5077 (N_5077,N_4305,N_4406);
nor U5078 (N_5078,N_4489,N_4588);
or U5079 (N_5079,N_4412,N_4896);
and U5080 (N_5080,N_4898,N_4166);
and U5081 (N_5081,N_4171,N_4788);
nand U5082 (N_5082,N_4841,N_4758);
and U5083 (N_5083,N_4193,N_4053);
nor U5084 (N_5084,N_4943,N_4910);
nand U5085 (N_5085,N_4208,N_4302);
nand U5086 (N_5086,N_4473,N_4198);
xnor U5087 (N_5087,N_4009,N_4906);
nor U5088 (N_5088,N_4899,N_4946);
nand U5089 (N_5089,N_4673,N_4569);
nor U5090 (N_5090,N_4353,N_4020);
nor U5091 (N_5091,N_4919,N_4277);
and U5092 (N_5092,N_4493,N_4523);
or U5093 (N_5093,N_4817,N_4285);
nor U5094 (N_5094,N_4080,N_4660);
or U5095 (N_5095,N_4846,N_4315);
nor U5096 (N_5096,N_4905,N_4570);
nand U5097 (N_5097,N_4925,N_4939);
and U5098 (N_5098,N_4087,N_4986);
or U5099 (N_5099,N_4314,N_4472);
and U5100 (N_5100,N_4388,N_4092);
or U5101 (N_5101,N_4551,N_4867);
nor U5102 (N_5102,N_4935,N_4710);
or U5103 (N_5103,N_4842,N_4414);
and U5104 (N_5104,N_4301,N_4114);
nand U5105 (N_5105,N_4382,N_4028);
nand U5106 (N_5106,N_4079,N_4157);
nand U5107 (N_5107,N_4931,N_4816);
nor U5108 (N_5108,N_4463,N_4970);
nor U5109 (N_5109,N_4852,N_4094);
and U5110 (N_5110,N_4796,N_4223);
nor U5111 (N_5111,N_4497,N_4077);
nor U5112 (N_5112,N_4336,N_4311);
or U5113 (N_5113,N_4753,N_4005);
nand U5114 (N_5114,N_4848,N_4065);
and U5115 (N_5115,N_4894,N_4482);
nand U5116 (N_5116,N_4828,N_4765);
and U5117 (N_5117,N_4086,N_4971);
nor U5118 (N_5118,N_4964,N_4617);
nor U5119 (N_5119,N_4851,N_4411);
nand U5120 (N_5120,N_4624,N_4176);
nand U5121 (N_5121,N_4204,N_4581);
or U5122 (N_5122,N_4441,N_4460);
and U5123 (N_5123,N_4284,N_4023);
and U5124 (N_5124,N_4000,N_4831);
nor U5125 (N_5125,N_4212,N_4667);
nand U5126 (N_5126,N_4490,N_4151);
nand U5127 (N_5127,N_4419,N_4701);
nor U5128 (N_5128,N_4409,N_4286);
nor U5129 (N_5129,N_4127,N_4025);
nand U5130 (N_5130,N_4976,N_4534);
or U5131 (N_5131,N_4862,N_4328);
and U5132 (N_5132,N_4260,N_4590);
nand U5133 (N_5133,N_4422,N_4677);
and U5134 (N_5134,N_4112,N_4818);
nand U5135 (N_5135,N_4641,N_4977);
nand U5136 (N_5136,N_4152,N_4429);
or U5137 (N_5137,N_4637,N_4368);
nor U5138 (N_5138,N_4448,N_4380);
or U5139 (N_5139,N_4201,N_4261);
or U5140 (N_5140,N_4398,N_4968);
nand U5141 (N_5141,N_4169,N_4690);
nand U5142 (N_5142,N_4962,N_4944);
and U5143 (N_5143,N_4243,N_4844);
xor U5144 (N_5144,N_4759,N_4052);
nand U5145 (N_5145,N_4825,N_4500);
or U5146 (N_5146,N_4869,N_4391);
nand U5147 (N_5147,N_4705,N_4304);
nand U5148 (N_5148,N_4684,N_4310);
nand U5149 (N_5149,N_4526,N_4004);
and U5150 (N_5150,N_4001,N_4525);
and U5151 (N_5151,N_4070,N_4779);
or U5152 (N_5152,N_4854,N_4133);
nor U5153 (N_5153,N_4707,N_4567);
nand U5154 (N_5154,N_4068,N_4423);
xnor U5155 (N_5155,N_4268,N_4140);
nor U5156 (N_5156,N_4274,N_4773);
and U5157 (N_5157,N_4681,N_4645);
xor U5158 (N_5158,N_4596,N_4903);
or U5159 (N_5159,N_4512,N_4126);
and U5160 (N_5160,N_4048,N_4991);
nor U5161 (N_5161,N_4104,N_4678);
nor U5162 (N_5162,N_4348,N_4202);
xor U5163 (N_5163,N_4544,N_4378);
and U5164 (N_5164,N_4583,N_4331);
and U5165 (N_5165,N_4047,N_4303);
nor U5166 (N_5166,N_4217,N_4006);
nor U5167 (N_5167,N_4804,N_4431);
nor U5168 (N_5168,N_4452,N_4289);
or U5169 (N_5169,N_4930,N_4873);
and U5170 (N_5170,N_4926,N_4599);
nand U5171 (N_5171,N_4981,N_4162);
nand U5172 (N_5172,N_4345,N_4764);
nand U5173 (N_5173,N_4824,N_4298);
and U5174 (N_5174,N_4095,N_4366);
or U5175 (N_5175,N_4075,N_4513);
xnor U5176 (N_5176,N_4658,N_4475);
and U5177 (N_5177,N_4837,N_4531);
and U5178 (N_5178,N_4341,N_4480);
nand U5179 (N_5179,N_4781,N_4119);
and U5180 (N_5180,N_4222,N_4974);
or U5181 (N_5181,N_4254,N_4184);
nor U5182 (N_5182,N_4952,N_4003);
nor U5183 (N_5183,N_4296,N_4642);
xnor U5184 (N_5184,N_4511,N_4170);
nor U5185 (N_5185,N_4547,N_4687);
or U5186 (N_5186,N_4835,N_4754);
and U5187 (N_5187,N_4739,N_4782);
nor U5188 (N_5188,N_4665,N_4682);
xor U5189 (N_5189,N_4727,N_4410);
or U5190 (N_5190,N_4251,N_4886);
and U5191 (N_5191,N_4030,N_4793);
nor U5192 (N_5192,N_4438,N_4015);
nand U5193 (N_5193,N_4211,N_4083);
or U5194 (N_5194,N_4874,N_4120);
nor U5195 (N_5195,N_4255,N_4912);
and U5196 (N_5196,N_4091,N_4364);
and U5197 (N_5197,N_4614,N_4458);
and U5198 (N_5198,N_4225,N_4989);
nor U5199 (N_5199,N_4736,N_4320);
or U5200 (N_5200,N_4757,N_4291);
and U5201 (N_5201,N_4605,N_4913);
or U5202 (N_5202,N_4787,N_4093);
xnor U5203 (N_5203,N_4447,N_4864);
nand U5204 (N_5204,N_4059,N_4027);
or U5205 (N_5205,N_4063,N_4768);
and U5206 (N_5206,N_4231,N_4692);
or U5207 (N_5207,N_4518,N_4041);
and U5208 (N_5208,N_4037,N_4771);
nand U5209 (N_5209,N_4393,N_4182);
nor U5210 (N_5210,N_4440,N_4502);
nor U5211 (N_5211,N_4538,N_4733);
or U5212 (N_5212,N_4603,N_4610);
xnor U5213 (N_5213,N_4156,N_4375);
nand U5214 (N_5214,N_4056,N_4664);
nand U5215 (N_5215,N_4612,N_4340);
and U5216 (N_5216,N_4872,N_4420);
nor U5217 (N_5217,N_4483,N_4143);
nor U5218 (N_5218,N_4891,N_4563);
xor U5219 (N_5219,N_4885,N_4108);
nor U5220 (N_5220,N_4282,N_4287);
and U5221 (N_5221,N_4948,N_4714);
nand U5222 (N_5222,N_4611,N_4703);
or U5223 (N_5223,N_4717,N_4139);
and U5224 (N_5224,N_4253,N_4392);
or U5225 (N_5225,N_4309,N_4742);
or U5226 (N_5226,N_4495,N_4085);
nand U5227 (N_5227,N_4330,N_4618);
and U5228 (N_5228,N_4267,N_4859);
nand U5229 (N_5229,N_4479,N_4099);
and U5230 (N_5230,N_4631,N_4121);
and U5231 (N_5231,N_4026,N_4809);
nand U5232 (N_5232,N_4516,N_4917);
or U5233 (N_5233,N_4887,N_4882);
nand U5234 (N_5234,N_4784,N_4973);
and U5235 (N_5235,N_4209,N_4623);
xor U5236 (N_5236,N_4181,N_4459);
and U5237 (N_5237,N_4744,N_4633);
nand U5238 (N_5238,N_4783,N_4347);
xnor U5239 (N_5239,N_4520,N_4235);
or U5240 (N_5240,N_4312,N_4464);
and U5241 (N_5241,N_4672,N_4795);
nor U5242 (N_5242,N_4355,N_4485);
and U5243 (N_5243,N_4179,N_4385);
nand U5244 (N_5244,N_4349,N_4279);
and U5245 (N_5245,N_4332,N_4792);
or U5246 (N_5246,N_4376,N_4504);
nand U5247 (N_5247,N_4741,N_4865);
xor U5248 (N_5248,N_4498,N_4510);
or U5249 (N_5249,N_4671,N_4486);
nor U5250 (N_5250,N_4019,N_4055);
and U5251 (N_5251,N_4826,N_4369);
xor U5252 (N_5252,N_4499,N_4323);
or U5253 (N_5253,N_4688,N_4668);
xor U5254 (N_5254,N_4858,N_4555);
nand U5255 (N_5255,N_4933,N_4435);
and U5256 (N_5256,N_4881,N_4514);
nor U5257 (N_5257,N_4165,N_4060);
nor U5258 (N_5258,N_4579,N_4556);
nand U5259 (N_5259,N_4295,N_4785);
nand U5260 (N_5260,N_4770,N_4521);
xnor U5261 (N_5261,N_4740,N_4592);
or U5262 (N_5262,N_4084,N_4014);
nand U5263 (N_5263,N_4798,N_4909);
nand U5264 (N_5264,N_4866,N_4923);
nand U5265 (N_5265,N_4342,N_4920);
nand U5266 (N_5266,N_4533,N_4515);
nor U5267 (N_5267,N_4158,N_4806);
nor U5268 (N_5268,N_4417,N_4519);
nand U5269 (N_5269,N_4994,N_4892);
and U5270 (N_5270,N_4262,N_4646);
or U5271 (N_5271,N_4980,N_4911);
nor U5272 (N_5272,N_4566,N_4381);
xor U5273 (N_5273,N_4426,N_4527);
or U5274 (N_5274,N_4478,N_4921);
and U5275 (N_5275,N_4876,N_4187);
or U5276 (N_5276,N_4405,N_4686);
and U5277 (N_5277,N_4481,N_4589);
and U5278 (N_5278,N_4750,N_4838);
and U5279 (N_5279,N_4992,N_4042);
or U5280 (N_5280,N_4871,N_4256);
or U5281 (N_5281,N_4934,N_4622);
and U5282 (N_5282,N_4800,N_4549);
nand U5283 (N_5283,N_4238,N_4443);
or U5284 (N_5284,N_4789,N_4932);
or U5285 (N_5285,N_4372,N_4959);
and U5286 (N_5286,N_4367,N_4942);
nor U5287 (N_5287,N_4361,N_4662);
xor U5288 (N_5288,N_4629,N_4338);
or U5289 (N_5289,N_4430,N_4593);
or U5290 (N_5290,N_4160,N_4730);
or U5291 (N_5291,N_4239,N_4109);
nor U5292 (N_5292,N_4103,N_4322);
nor U5293 (N_5293,N_4829,N_4878);
nand U5294 (N_5294,N_4021,N_4794);
and U5295 (N_5295,N_4895,N_4220);
and U5296 (N_5296,N_4805,N_4706);
nand U5297 (N_5297,N_4273,N_4313);
and U5298 (N_5298,N_4998,N_4729);
and U5299 (N_5299,N_4321,N_4748);
nor U5300 (N_5300,N_4543,N_4702);
nor U5301 (N_5301,N_4967,N_4008);
or U5302 (N_5302,N_4031,N_4288);
and U5303 (N_5303,N_4914,N_4234);
xor U5304 (N_5304,N_4843,N_4997);
and U5305 (N_5305,N_4833,N_4421);
nand U5306 (N_5306,N_4762,N_4029);
xnor U5307 (N_5307,N_4602,N_4428);
xnor U5308 (N_5308,N_4307,N_4246);
or U5309 (N_5309,N_4836,N_4033);
and U5310 (N_5310,N_4893,N_4432);
and U5311 (N_5311,N_4613,N_4427);
nor U5312 (N_5312,N_4880,N_4814);
xor U5313 (N_5313,N_4760,N_4761);
nand U5314 (N_5314,N_4649,N_4638);
nand U5315 (N_5315,N_4319,N_4130);
nand U5316 (N_5316,N_4449,N_4123);
nand U5317 (N_5317,N_4207,N_4402);
nor U5318 (N_5318,N_4245,N_4216);
nand U5319 (N_5319,N_4975,N_4767);
nor U5320 (N_5320,N_4695,N_4446);
nand U5321 (N_5321,N_4632,N_4689);
nor U5322 (N_5322,N_4168,N_4110);
or U5323 (N_5323,N_4469,N_4987);
and U5324 (N_5324,N_4735,N_4424);
nor U5325 (N_5325,N_4191,N_4149);
nand U5326 (N_5326,N_4606,N_4901);
and U5327 (N_5327,N_4657,N_4517);
and U5328 (N_5328,N_4397,N_4496);
nand U5329 (N_5329,N_4751,N_4106);
and U5330 (N_5330,N_4680,N_4264);
nor U5331 (N_5331,N_4354,N_4465);
nand U5332 (N_5332,N_4404,N_4746);
and U5333 (N_5333,N_4248,N_4265);
nand U5334 (N_5334,N_4653,N_4035);
and U5335 (N_5335,N_4993,N_4704);
nand U5336 (N_5336,N_4039,N_4591);
nand U5337 (N_5337,N_4118,N_4275);
xor U5338 (N_5338,N_4786,N_4113);
nand U5339 (N_5339,N_4178,N_4281);
or U5340 (N_5340,N_4766,N_4373);
xnor U5341 (N_5341,N_4073,N_4032);
or U5342 (N_5342,N_4928,N_4403);
xor U5343 (N_5343,N_4548,N_4737);
nor U5344 (N_5344,N_4002,N_4131);
and U5345 (N_5345,N_4557,N_4956);
xnor U5346 (N_5346,N_4346,N_4969);
xnor U5347 (N_5347,N_4362,N_4965);
or U5348 (N_5348,N_4142,N_4230);
nand U5349 (N_5349,N_4190,N_4067);
and U5350 (N_5350,N_4957,N_4155);
nand U5351 (N_5351,N_4868,N_4636);
or U5352 (N_5352,N_4144,N_4334);
nand U5353 (N_5353,N_4038,N_4609);
or U5354 (N_5354,N_4937,N_4066);
or U5355 (N_5355,N_4145,N_4963);
nor U5356 (N_5356,N_4947,N_4883);
or U5357 (N_5357,N_4399,N_4434);
and U5358 (N_5358,N_4640,N_4501);
or U5359 (N_5359,N_4226,N_4999);
nor U5360 (N_5360,N_4620,N_4259);
or U5361 (N_5361,N_4467,N_4471);
and U5362 (N_5362,N_4175,N_4416);
or U5363 (N_5363,N_4763,N_4012);
and U5364 (N_5364,N_4173,N_4218);
or U5365 (N_5365,N_4016,N_4860);
nand U5366 (N_5366,N_4125,N_4568);
nor U5367 (N_5367,N_4487,N_4249);
and U5368 (N_5368,N_4877,N_4738);
and U5369 (N_5369,N_4200,N_4985);
nor U5370 (N_5370,N_4654,N_4082);
or U5371 (N_5371,N_4050,N_4508);
nand U5372 (N_5372,N_4335,N_4834);
or U5373 (N_5373,N_4455,N_4189);
xnor U5374 (N_5374,N_4685,N_4071);
nor U5375 (N_5375,N_4666,N_4683);
and U5376 (N_5376,N_4749,N_4229);
nand U5377 (N_5377,N_4832,N_4177);
and U5378 (N_5378,N_4575,N_4148);
nand U5379 (N_5379,N_4845,N_4324);
or U5380 (N_5380,N_4453,N_4221);
and U5381 (N_5381,N_4608,N_4822);
or U5382 (N_5382,N_4270,N_4728);
nand U5383 (N_5383,N_4237,N_4102);
nor U5384 (N_5384,N_4343,N_4101);
or U5385 (N_5385,N_4509,N_4560);
xnor U5386 (N_5386,N_4205,N_4159);
nand U5387 (N_5387,N_4559,N_4370);
and U5388 (N_5388,N_4022,N_4545);
and U5389 (N_5389,N_4745,N_4813);
xor U5390 (N_5390,N_4293,N_4344);
nand U5391 (N_5391,N_4747,N_4197);
nand U5392 (N_5392,N_4644,N_4199);
nor U5393 (N_5393,N_4811,N_4192);
or U5394 (N_5394,N_4377,N_4051);
nor U5395 (N_5395,N_4462,N_4918);
nand U5396 (N_5396,N_4445,N_4776);
nand U5397 (N_5397,N_4210,N_4492);
and U5398 (N_5398,N_4619,N_4280);
nand U5399 (N_5399,N_4196,N_4013);
and U5400 (N_5400,N_4442,N_4389);
nand U5401 (N_5401,N_4650,N_4154);
nand U5402 (N_5402,N_4088,N_4550);
or U5403 (N_5403,N_4815,N_4470);
and U5404 (N_5404,N_4732,N_4916);
or U5405 (N_5405,N_4535,N_4185);
nor U5406 (N_5406,N_4542,N_4529);
and U5407 (N_5407,N_4163,N_4573);
nor U5408 (N_5408,N_4107,N_4507);
or U5409 (N_5409,N_4582,N_4081);
or U5410 (N_5410,N_4656,N_4819);
nand U5411 (N_5411,N_4564,N_4384);
and U5412 (N_5412,N_4017,N_4539);
and U5413 (N_5413,N_4951,N_4116);
nor U5414 (N_5414,N_4129,N_4780);
or U5415 (N_5415,N_4699,N_4884);
and U5416 (N_5416,N_4276,N_4219);
nor U5417 (N_5417,N_4983,N_4718);
nand U5418 (N_5418,N_4674,N_4054);
xnor U5419 (N_5419,N_4300,N_4505);
and U5420 (N_5420,N_4978,N_4247);
or U5421 (N_5421,N_4503,N_4250);
nand U5422 (N_5422,N_4174,N_4639);
or U5423 (N_5423,N_4996,N_4949);
or U5424 (N_5424,N_4812,N_4802);
nand U5425 (N_5425,N_4044,N_4574);
nand U5426 (N_5426,N_4290,N_4924);
and U5427 (N_5427,N_4723,N_4128);
and U5428 (N_5428,N_4594,N_4797);
nand U5429 (N_5429,N_4995,N_4663);
nand U5430 (N_5430,N_4708,N_4141);
and U5431 (N_5431,N_4731,N_4984);
and U5432 (N_5432,N_4450,N_4936);
xor U5433 (N_5433,N_4425,N_4371);
nor U5434 (N_5434,N_4062,N_4266);
nor U5435 (N_5435,N_4532,N_4972);
nand U5436 (N_5436,N_4135,N_4461);
or U5437 (N_5437,N_4840,N_4897);
or U5438 (N_5438,N_4386,N_4530);
nand U5439 (N_5439,N_4888,N_4577);
or U5440 (N_5440,N_4360,N_4488);
and U5441 (N_5441,N_4046,N_4801);
and U5442 (N_5442,N_4670,N_4132);
nand U5443 (N_5443,N_4830,N_4725);
and U5444 (N_5444,N_4308,N_4724);
nand U5445 (N_5445,N_4713,N_4401);
nand U5446 (N_5446,N_4875,N_4379);
nor U5447 (N_5447,N_4213,N_4466);
and U5448 (N_5448,N_4536,N_4698);
or U5449 (N_5449,N_4571,N_4778);
or U5450 (N_5450,N_4576,N_4849);
nor U5451 (N_5451,N_4572,N_4938);
and U5452 (N_5452,N_4676,N_4147);
or U5453 (N_5453,N_4506,N_4111);
nor U5454 (N_5454,N_4024,N_4607);
and U5455 (N_5455,N_4186,N_4272);
nor U5456 (N_5456,N_4870,N_4058);
or U5457 (N_5457,N_4769,N_4271);
nand U5458 (N_5458,N_4627,N_4444);
nand U5459 (N_5459,N_4715,N_4655);
or U5460 (N_5460,N_4105,N_4580);
and U5461 (N_5461,N_4097,N_4900);
or U5462 (N_5462,N_4904,N_4365);
xor U5463 (N_5463,N_4252,N_4395);
nor U5464 (N_5464,N_4661,N_4711);
and U5465 (N_5465,N_4541,N_4115);
or U5466 (N_5466,N_4010,N_4693);
xnor U5467 (N_5467,N_4439,N_4927);
or U5468 (N_5468,N_4433,N_4161);
xor U5469 (N_5469,N_4172,N_4240);
and U5470 (N_5470,N_4045,N_4752);
nor U5471 (N_5471,N_4808,N_4908);
nand U5472 (N_5472,N_4195,N_4890);
nor U5473 (N_5473,N_4394,N_4327);
xnor U5474 (N_5474,N_4150,N_4839);
and U5475 (N_5475,N_4561,N_4011);
or U5476 (N_5476,N_4018,N_4215);
and U5477 (N_5477,N_4696,N_4317);
or U5478 (N_5478,N_4803,N_4468);
and U5479 (N_5479,N_4616,N_4915);
and U5480 (N_5480,N_4183,N_4712);
or U5481 (N_5481,N_4034,N_4137);
nand U5482 (N_5482,N_4098,N_4457);
or U5483 (N_5483,N_4374,N_4451);
and U5484 (N_5484,N_4601,N_4258);
and U5485 (N_5485,N_4242,N_4950);
nand U5486 (N_5486,N_4294,N_4628);
and U5487 (N_5487,N_4586,N_4621);
nor U5488 (N_5488,N_4064,N_4675);
nand U5489 (N_5489,N_4350,N_4036);
nand U5490 (N_5490,N_4203,N_4363);
and U5491 (N_5491,N_4396,N_4292);
nand U5492 (N_5492,N_4604,N_4351);
or U5493 (N_5493,N_4359,N_4595);
and U5494 (N_5494,N_4546,N_4089);
nand U5495 (N_5495,N_4982,N_4061);
and U5496 (N_5496,N_4647,N_4043);
nand U5497 (N_5497,N_4734,N_4553);
nor U5498 (N_5498,N_4643,N_4600);
nand U5499 (N_5499,N_4326,N_4648);
or U5500 (N_5500,N_4985,N_4814);
and U5501 (N_5501,N_4856,N_4179);
or U5502 (N_5502,N_4767,N_4141);
and U5503 (N_5503,N_4193,N_4851);
nand U5504 (N_5504,N_4242,N_4560);
and U5505 (N_5505,N_4132,N_4830);
or U5506 (N_5506,N_4193,N_4556);
and U5507 (N_5507,N_4598,N_4215);
nand U5508 (N_5508,N_4356,N_4072);
and U5509 (N_5509,N_4146,N_4273);
nor U5510 (N_5510,N_4465,N_4440);
or U5511 (N_5511,N_4507,N_4042);
or U5512 (N_5512,N_4490,N_4890);
or U5513 (N_5513,N_4908,N_4181);
nand U5514 (N_5514,N_4162,N_4365);
nor U5515 (N_5515,N_4139,N_4752);
nand U5516 (N_5516,N_4432,N_4569);
nor U5517 (N_5517,N_4477,N_4781);
and U5518 (N_5518,N_4999,N_4583);
nor U5519 (N_5519,N_4444,N_4834);
nor U5520 (N_5520,N_4333,N_4520);
nor U5521 (N_5521,N_4523,N_4191);
nand U5522 (N_5522,N_4416,N_4796);
nor U5523 (N_5523,N_4375,N_4916);
nor U5524 (N_5524,N_4855,N_4490);
nand U5525 (N_5525,N_4489,N_4647);
nand U5526 (N_5526,N_4798,N_4985);
nand U5527 (N_5527,N_4662,N_4450);
and U5528 (N_5528,N_4284,N_4055);
and U5529 (N_5529,N_4621,N_4771);
xnor U5530 (N_5530,N_4585,N_4534);
and U5531 (N_5531,N_4987,N_4853);
and U5532 (N_5532,N_4965,N_4141);
nand U5533 (N_5533,N_4729,N_4285);
or U5534 (N_5534,N_4457,N_4920);
xor U5535 (N_5535,N_4681,N_4313);
nor U5536 (N_5536,N_4555,N_4130);
nand U5537 (N_5537,N_4931,N_4796);
xnor U5538 (N_5538,N_4601,N_4434);
and U5539 (N_5539,N_4235,N_4420);
nand U5540 (N_5540,N_4092,N_4747);
and U5541 (N_5541,N_4302,N_4675);
nor U5542 (N_5542,N_4969,N_4955);
xnor U5543 (N_5543,N_4573,N_4147);
and U5544 (N_5544,N_4440,N_4710);
nand U5545 (N_5545,N_4428,N_4159);
xnor U5546 (N_5546,N_4175,N_4669);
xnor U5547 (N_5547,N_4763,N_4278);
nor U5548 (N_5548,N_4671,N_4963);
nand U5549 (N_5549,N_4659,N_4930);
or U5550 (N_5550,N_4167,N_4999);
or U5551 (N_5551,N_4918,N_4105);
nor U5552 (N_5552,N_4333,N_4956);
nor U5553 (N_5553,N_4864,N_4172);
and U5554 (N_5554,N_4590,N_4366);
xnor U5555 (N_5555,N_4564,N_4699);
or U5556 (N_5556,N_4007,N_4801);
nor U5557 (N_5557,N_4995,N_4326);
or U5558 (N_5558,N_4479,N_4938);
or U5559 (N_5559,N_4204,N_4525);
nor U5560 (N_5560,N_4992,N_4341);
nand U5561 (N_5561,N_4707,N_4590);
and U5562 (N_5562,N_4982,N_4938);
nand U5563 (N_5563,N_4576,N_4464);
xnor U5564 (N_5564,N_4000,N_4901);
nor U5565 (N_5565,N_4399,N_4693);
nand U5566 (N_5566,N_4442,N_4125);
or U5567 (N_5567,N_4244,N_4848);
nand U5568 (N_5568,N_4042,N_4935);
nor U5569 (N_5569,N_4987,N_4025);
and U5570 (N_5570,N_4824,N_4908);
nand U5571 (N_5571,N_4484,N_4677);
or U5572 (N_5572,N_4205,N_4384);
nor U5573 (N_5573,N_4159,N_4172);
nor U5574 (N_5574,N_4952,N_4076);
and U5575 (N_5575,N_4061,N_4619);
nor U5576 (N_5576,N_4082,N_4304);
nand U5577 (N_5577,N_4675,N_4734);
nand U5578 (N_5578,N_4911,N_4353);
or U5579 (N_5579,N_4670,N_4193);
nor U5580 (N_5580,N_4017,N_4012);
nand U5581 (N_5581,N_4881,N_4116);
nand U5582 (N_5582,N_4845,N_4917);
nor U5583 (N_5583,N_4434,N_4411);
nand U5584 (N_5584,N_4949,N_4907);
nand U5585 (N_5585,N_4985,N_4470);
or U5586 (N_5586,N_4198,N_4974);
nor U5587 (N_5587,N_4186,N_4735);
nand U5588 (N_5588,N_4706,N_4963);
and U5589 (N_5589,N_4284,N_4477);
or U5590 (N_5590,N_4406,N_4781);
and U5591 (N_5591,N_4425,N_4995);
or U5592 (N_5592,N_4274,N_4040);
nand U5593 (N_5593,N_4740,N_4656);
or U5594 (N_5594,N_4335,N_4495);
nand U5595 (N_5595,N_4756,N_4220);
nand U5596 (N_5596,N_4835,N_4253);
xor U5597 (N_5597,N_4807,N_4617);
nand U5598 (N_5598,N_4714,N_4861);
nand U5599 (N_5599,N_4934,N_4260);
nand U5600 (N_5600,N_4095,N_4241);
nand U5601 (N_5601,N_4847,N_4494);
and U5602 (N_5602,N_4361,N_4629);
nor U5603 (N_5603,N_4916,N_4298);
and U5604 (N_5604,N_4632,N_4886);
nor U5605 (N_5605,N_4641,N_4256);
nand U5606 (N_5606,N_4890,N_4975);
nand U5607 (N_5607,N_4935,N_4013);
nor U5608 (N_5608,N_4456,N_4099);
nand U5609 (N_5609,N_4180,N_4565);
xor U5610 (N_5610,N_4182,N_4923);
nor U5611 (N_5611,N_4690,N_4428);
and U5612 (N_5612,N_4011,N_4356);
and U5613 (N_5613,N_4929,N_4692);
xnor U5614 (N_5614,N_4784,N_4871);
or U5615 (N_5615,N_4887,N_4661);
or U5616 (N_5616,N_4380,N_4771);
nand U5617 (N_5617,N_4967,N_4267);
xor U5618 (N_5618,N_4717,N_4896);
and U5619 (N_5619,N_4320,N_4375);
or U5620 (N_5620,N_4990,N_4346);
or U5621 (N_5621,N_4821,N_4952);
nor U5622 (N_5622,N_4652,N_4193);
and U5623 (N_5623,N_4486,N_4316);
xor U5624 (N_5624,N_4791,N_4735);
nor U5625 (N_5625,N_4733,N_4525);
and U5626 (N_5626,N_4083,N_4525);
and U5627 (N_5627,N_4601,N_4829);
xnor U5628 (N_5628,N_4821,N_4517);
nand U5629 (N_5629,N_4677,N_4883);
or U5630 (N_5630,N_4023,N_4547);
nand U5631 (N_5631,N_4185,N_4708);
nand U5632 (N_5632,N_4760,N_4058);
and U5633 (N_5633,N_4528,N_4471);
or U5634 (N_5634,N_4892,N_4215);
nand U5635 (N_5635,N_4701,N_4604);
nor U5636 (N_5636,N_4914,N_4218);
nand U5637 (N_5637,N_4856,N_4458);
nand U5638 (N_5638,N_4092,N_4487);
nand U5639 (N_5639,N_4045,N_4434);
nor U5640 (N_5640,N_4889,N_4861);
xor U5641 (N_5641,N_4624,N_4559);
xnor U5642 (N_5642,N_4976,N_4233);
and U5643 (N_5643,N_4794,N_4836);
nor U5644 (N_5644,N_4790,N_4607);
nor U5645 (N_5645,N_4587,N_4344);
or U5646 (N_5646,N_4851,N_4582);
or U5647 (N_5647,N_4543,N_4839);
nor U5648 (N_5648,N_4596,N_4197);
nor U5649 (N_5649,N_4205,N_4386);
nand U5650 (N_5650,N_4069,N_4343);
nor U5651 (N_5651,N_4332,N_4589);
and U5652 (N_5652,N_4148,N_4660);
or U5653 (N_5653,N_4095,N_4443);
and U5654 (N_5654,N_4675,N_4741);
and U5655 (N_5655,N_4237,N_4180);
nor U5656 (N_5656,N_4220,N_4878);
nor U5657 (N_5657,N_4182,N_4838);
or U5658 (N_5658,N_4610,N_4437);
and U5659 (N_5659,N_4016,N_4357);
nand U5660 (N_5660,N_4191,N_4309);
and U5661 (N_5661,N_4497,N_4942);
nand U5662 (N_5662,N_4972,N_4868);
nor U5663 (N_5663,N_4438,N_4511);
nor U5664 (N_5664,N_4986,N_4604);
or U5665 (N_5665,N_4638,N_4598);
nor U5666 (N_5666,N_4646,N_4363);
nand U5667 (N_5667,N_4857,N_4268);
or U5668 (N_5668,N_4239,N_4566);
nor U5669 (N_5669,N_4901,N_4265);
nor U5670 (N_5670,N_4542,N_4690);
nand U5671 (N_5671,N_4692,N_4116);
xnor U5672 (N_5672,N_4294,N_4614);
nand U5673 (N_5673,N_4758,N_4685);
nor U5674 (N_5674,N_4023,N_4563);
nand U5675 (N_5675,N_4659,N_4828);
nor U5676 (N_5676,N_4904,N_4932);
or U5677 (N_5677,N_4468,N_4348);
nand U5678 (N_5678,N_4702,N_4931);
nand U5679 (N_5679,N_4277,N_4034);
xnor U5680 (N_5680,N_4277,N_4017);
and U5681 (N_5681,N_4795,N_4936);
nand U5682 (N_5682,N_4338,N_4413);
nor U5683 (N_5683,N_4799,N_4741);
nor U5684 (N_5684,N_4570,N_4088);
xnor U5685 (N_5685,N_4226,N_4898);
nand U5686 (N_5686,N_4717,N_4226);
nand U5687 (N_5687,N_4924,N_4730);
and U5688 (N_5688,N_4083,N_4112);
and U5689 (N_5689,N_4628,N_4946);
or U5690 (N_5690,N_4916,N_4841);
and U5691 (N_5691,N_4387,N_4439);
nor U5692 (N_5692,N_4230,N_4137);
or U5693 (N_5693,N_4791,N_4371);
nor U5694 (N_5694,N_4651,N_4069);
or U5695 (N_5695,N_4399,N_4129);
xnor U5696 (N_5696,N_4865,N_4545);
nand U5697 (N_5697,N_4529,N_4903);
nand U5698 (N_5698,N_4954,N_4547);
and U5699 (N_5699,N_4104,N_4063);
nor U5700 (N_5700,N_4001,N_4074);
xor U5701 (N_5701,N_4313,N_4645);
nand U5702 (N_5702,N_4251,N_4097);
and U5703 (N_5703,N_4765,N_4110);
nor U5704 (N_5704,N_4088,N_4122);
or U5705 (N_5705,N_4360,N_4705);
nand U5706 (N_5706,N_4505,N_4035);
or U5707 (N_5707,N_4743,N_4062);
nor U5708 (N_5708,N_4304,N_4137);
or U5709 (N_5709,N_4717,N_4245);
nand U5710 (N_5710,N_4799,N_4946);
nor U5711 (N_5711,N_4670,N_4770);
and U5712 (N_5712,N_4414,N_4637);
and U5713 (N_5713,N_4326,N_4158);
or U5714 (N_5714,N_4847,N_4588);
or U5715 (N_5715,N_4346,N_4366);
and U5716 (N_5716,N_4470,N_4519);
nor U5717 (N_5717,N_4413,N_4942);
and U5718 (N_5718,N_4084,N_4604);
nand U5719 (N_5719,N_4887,N_4693);
or U5720 (N_5720,N_4554,N_4668);
or U5721 (N_5721,N_4464,N_4110);
nor U5722 (N_5722,N_4732,N_4255);
and U5723 (N_5723,N_4723,N_4029);
nor U5724 (N_5724,N_4685,N_4923);
or U5725 (N_5725,N_4148,N_4237);
or U5726 (N_5726,N_4102,N_4782);
or U5727 (N_5727,N_4920,N_4953);
nand U5728 (N_5728,N_4302,N_4968);
and U5729 (N_5729,N_4066,N_4586);
nand U5730 (N_5730,N_4123,N_4800);
nor U5731 (N_5731,N_4094,N_4273);
xnor U5732 (N_5732,N_4927,N_4820);
and U5733 (N_5733,N_4264,N_4606);
xor U5734 (N_5734,N_4915,N_4289);
and U5735 (N_5735,N_4561,N_4626);
nor U5736 (N_5736,N_4703,N_4751);
nand U5737 (N_5737,N_4338,N_4711);
or U5738 (N_5738,N_4292,N_4052);
nor U5739 (N_5739,N_4425,N_4080);
and U5740 (N_5740,N_4980,N_4845);
nor U5741 (N_5741,N_4655,N_4876);
nand U5742 (N_5742,N_4127,N_4040);
and U5743 (N_5743,N_4340,N_4866);
nand U5744 (N_5744,N_4486,N_4845);
nand U5745 (N_5745,N_4002,N_4643);
and U5746 (N_5746,N_4395,N_4064);
and U5747 (N_5747,N_4876,N_4058);
nand U5748 (N_5748,N_4435,N_4585);
and U5749 (N_5749,N_4688,N_4167);
xor U5750 (N_5750,N_4125,N_4937);
or U5751 (N_5751,N_4522,N_4661);
nand U5752 (N_5752,N_4990,N_4302);
or U5753 (N_5753,N_4960,N_4037);
or U5754 (N_5754,N_4524,N_4261);
or U5755 (N_5755,N_4955,N_4927);
nor U5756 (N_5756,N_4818,N_4139);
and U5757 (N_5757,N_4847,N_4084);
and U5758 (N_5758,N_4632,N_4757);
and U5759 (N_5759,N_4445,N_4540);
nor U5760 (N_5760,N_4882,N_4040);
nand U5761 (N_5761,N_4388,N_4246);
and U5762 (N_5762,N_4300,N_4844);
or U5763 (N_5763,N_4580,N_4195);
and U5764 (N_5764,N_4101,N_4188);
nor U5765 (N_5765,N_4492,N_4801);
and U5766 (N_5766,N_4638,N_4730);
or U5767 (N_5767,N_4276,N_4827);
or U5768 (N_5768,N_4487,N_4785);
or U5769 (N_5769,N_4072,N_4043);
nor U5770 (N_5770,N_4643,N_4539);
nor U5771 (N_5771,N_4358,N_4203);
nor U5772 (N_5772,N_4434,N_4275);
or U5773 (N_5773,N_4894,N_4066);
nor U5774 (N_5774,N_4046,N_4522);
nor U5775 (N_5775,N_4081,N_4167);
nand U5776 (N_5776,N_4527,N_4824);
nor U5777 (N_5777,N_4277,N_4529);
nor U5778 (N_5778,N_4547,N_4097);
or U5779 (N_5779,N_4093,N_4143);
or U5780 (N_5780,N_4824,N_4185);
and U5781 (N_5781,N_4040,N_4159);
or U5782 (N_5782,N_4971,N_4908);
xnor U5783 (N_5783,N_4659,N_4657);
nor U5784 (N_5784,N_4380,N_4077);
nand U5785 (N_5785,N_4933,N_4418);
or U5786 (N_5786,N_4927,N_4469);
and U5787 (N_5787,N_4045,N_4288);
nor U5788 (N_5788,N_4367,N_4578);
nor U5789 (N_5789,N_4691,N_4934);
xor U5790 (N_5790,N_4563,N_4516);
xor U5791 (N_5791,N_4297,N_4038);
or U5792 (N_5792,N_4960,N_4183);
nor U5793 (N_5793,N_4503,N_4842);
nor U5794 (N_5794,N_4640,N_4139);
and U5795 (N_5795,N_4460,N_4911);
or U5796 (N_5796,N_4151,N_4788);
xnor U5797 (N_5797,N_4926,N_4731);
nor U5798 (N_5798,N_4030,N_4768);
or U5799 (N_5799,N_4688,N_4822);
nor U5800 (N_5800,N_4702,N_4687);
and U5801 (N_5801,N_4538,N_4832);
nand U5802 (N_5802,N_4664,N_4934);
nand U5803 (N_5803,N_4578,N_4602);
and U5804 (N_5804,N_4343,N_4129);
and U5805 (N_5805,N_4142,N_4012);
nor U5806 (N_5806,N_4420,N_4302);
nor U5807 (N_5807,N_4609,N_4928);
nor U5808 (N_5808,N_4385,N_4017);
nand U5809 (N_5809,N_4703,N_4286);
nand U5810 (N_5810,N_4587,N_4493);
xor U5811 (N_5811,N_4004,N_4051);
xor U5812 (N_5812,N_4020,N_4325);
or U5813 (N_5813,N_4331,N_4036);
or U5814 (N_5814,N_4924,N_4307);
and U5815 (N_5815,N_4078,N_4247);
xor U5816 (N_5816,N_4509,N_4079);
xor U5817 (N_5817,N_4408,N_4237);
or U5818 (N_5818,N_4253,N_4057);
nor U5819 (N_5819,N_4621,N_4265);
and U5820 (N_5820,N_4274,N_4488);
nand U5821 (N_5821,N_4348,N_4108);
and U5822 (N_5822,N_4273,N_4036);
nor U5823 (N_5823,N_4404,N_4563);
and U5824 (N_5824,N_4839,N_4702);
xnor U5825 (N_5825,N_4905,N_4782);
and U5826 (N_5826,N_4878,N_4025);
or U5827 (N_5827,N_4095,N_4431);
nor U5828 (N_5828,N_4948,N_4411);
or U5829 (N_5829,N_4545,N_4081);
and U5830 (N_5830,N_4063,N_4043);
and U5831 (N_5831,N_4088,N_4620);
and U5832 (N_5832,N_4630,N_4962);
or U5833 (N_5833,N_4801,N_4185);
nor U5834 (N_5834,N_4045,N_4569);
nand U5835 (N_5835,N_4677,N_4037);
xnor U5836 (N_5836,N_4204,N_4580);
nor U5837 (N_5837,N_4585,N_4495);
nand U5838 (N_5838,N_4577,N_4922);
nand U5839 (N_5839,N_4594,N_4518);
xnor U5840 (N_5840,N_4852,N_4737);
and U5841 (N_5841,N_4317,N_4254);
or U5842 (N_5842,N_4306,N_4813);
nand U5843 (N_5843,N_4737,N_4147);
nor U5844 (N_5844,N_4287,N_4681);
xor U5845 (N_5845,N_4489,N_4417);
or U5846 (N_5846,N_4620,N_4813);
or U5847 (N_5847,N_4497,N_4717);
or U5848 (N_5848,N_4389,N_4159);
or U5849 (N_5849,N_4044,N_4463);
and U5850 (N_5850,N_4833,N_4471);
and U5851 (N_5851,N_4803,N_4059);
nor U5852 (N_5852,N_4367,N_4377);
nand U5853 (N_5853,N_4116,N_4163);
nor U5854 (N_5854,N_4587,N_4928);
xnor U5855 (N_5855,N_4255,N_4208);
and U5856 (N_5856,N_4301,N_4054);
nor U5857 (N_5857,N_4310,N_4885);
nand U5858 (N_5858,N_4169,N_4424);
nand U5859 (N_5859,N_4124,N_4600);
nand U5860 (N_5860,N_4495,N_4362);
and U5861 (N_5861,N_4840,N_4530);
xor U5862 (N_5862,N_4170,N_4766);
nor U5863 (N_5863,N_4710,N_4947);
nor U5864 (N_5864,N_4352,N_4697);
or U5865 (N_5865,N_4036,N_4166);
nand U5866 (N_5866,N_4047,N_4281);
nor U5867 (N_5867,N_4867,N_4168);
nor U5868 (N_5868,N_4199,N_4316);
nand U5869 (N_5869,N_4289,N_4584);
xor U5870 (N_5870,N_4933,N_4991);
nand U5871 (N_5871,N_4885,N_4946);
or U5872 (N_5872,N_4757,N_4104);
xor U5873 (N_5873,N_4160,N_4573);
nand U5874 (N_5874,N_4981,N_4637);
or U5875 (N_5875,N_4649,N_4705);
or U5876 (N_5876,N_4157,N_4000);
and U5877 (N_5877,N_4168,N_4950);
and U5878 (N_5878,N_4238,N_4552);
nor U5879 (N_5879,N_4262,N_4496);
or U5880 (N_5880,N_4505,N_4956);
or U5881 (N_5881,N_4720,N_4439);
and U5882 (N_5882,N_4159,N_4780);
nor U5883 (N_5883,N_4183,N_4144);
nand U5884 (N_5884,N_4920,N_4008);
nand U5885 (N_5885,N_4229,N_4758);
or U5886 (N_5886,N_4758,N_4081);
nand U5887 (N_5887,N_4315,N_4190);
nand U5888 (N_5888,N_4441,N_4532);
nand U5889 (N_5889,N_4751,N_4528);
and U5890 (N_5890,N_4329,N_4872);
and U5891 (N_5891,N_4027,N_4847);
nor U5892 (N_5892,N_4906,N_4448);
or U5893 (N_5893,N_4234,N_4249);
nor U5894 (N_5894,N_4805,N_4298);
or U5895 (N_5895,N_4510,N_4759);
nand U5896 (N_5896,N_4263,N_4495);
nand U5897 (N_5897,N_4990,N_4431);
xnor U5898 (N_5898,N_4214,N_4338);
nand U5899 (N_5899,N_4419,N_4132);
and U5900 (N_5900,N_4334,N_4993);
nand U5901 (N_5901,N_4486,N_4864);
and U5902 (N_5902,N_4354,N_4864);
nor U5903 (N_5903,N_4138,N_4321);
or U5904 (N_5904,N_4611,N_4470);
or U5905 (N_5905,N_4112,N_4831);
nor U5906 (N_5906,N_4686,N_4441);
nor U5907 (N_5907,N_4309,N_4728);
nor U5908 (N_5908,N_4346,N_4227);
nand U5909 (N_5909,N_4919,N_4887);
nor U5910 (N_5910,N_4120,N_4438);
nor U5911 (N_5911,N_4762,N_4730);
and U5912 (N_5912,N_4435,N_4556);
or U5913 (N_5913,N_4405,N_4616);
nand U5914 (N_5914,N_4654,N_4197);
or U5915 (N_5915,N_4501,N_4152);
xor U5916 (N_5916,N_4186,N_4655);
nand U5917 (N_5917,N_4024,N_4248);
or U5918 (N_5918,N_4906,N_4834);
and U5919 (N_5919,N_4422,N_4453);
nand U5920 (N_5920,N_4921,N_4109);
or U5921 (N_5921,N_4937,N_4205);
and U5922 (N_5922,N_4573,N_4887);
nor U5923 (N_5923,N_4493,N_4558);
nor U5924 (N_5924,N_4057,N_4598);
nand U5925 (N_5925,N_4729,N_4133);
and U5926 (N_5926,N_4756,N_4874);
xnor U5927 (N_5927,N_4120,N_4047);
xor U5928 (N_5928,N_4955,N_4620);
and U5929 (N_5929,N_4259,N_4328);
or U5930 (N_5930,N_4818,N_4622);
nand U5931 (N_5931,N_4767,N_4523);
or U5932 (N_5932,N_4064,N_4868);
xnor U5933 (N_5933,N_4329,N_4916);
nor U5934 (N_5934,N_4257,N_4084);
or U5935 (N_5935,N_4955,N_4559);
and U5936 (N_5936,N_4451,N_4735);
nor U5937 (N_5937,N_4178,N_4256);
and U5938 (N_5938,N_4304,N_4780);
nand U5939 (N_5939,N_4416,N_4666);
or U5940 (N_5940,N_4555,N_4606);
or U5941 (N_5941,N_4282,N_4049);
and U5942 (N_5942,N_4175,N_4637);
nand U5943 (N_5943,N_4370,N_4873);
xnor U5944 (N_5944,N_4933,N_4402);
and U5945 (N_5945,N_4408,N_4469);
or U5946 (N_5946,N_4184,N_4099);
or U5947 (N_5947,N_4149,N_4288);
or U5948 (N_5948,N_4826,N_4714);
nor U5949 (N_5949,N_4185,N_4749);
nor U5950 (N_5950,N_4029,N_4947);
nand U5951 (N_5951,N_4173,N_4937);
and U5952 (N_5952,N_4069,N_4054);
nand U5953 (N_5953,N_4970,N_4804);
and U5954 (N_5954,N_4898,N_4358);
nor U5955 (N_5955,N_4797,N_4864);
nand U5956 (N_5956,N_4815,N_4996);
and U5957 (N_5957,N_4173,N_4264);
and U5958 (N_5958,N_4098,N_4899);
xnor U5959 (N_5959,N_4520,N_4921);
nor U5960 (N_5960,N_4908,N_4441);
or U5961 (N_5961,N_4228,N_4916);
nand U5962 (N_5962,N_4829,N_4005);
nor U5963 (N_5963,N_4199,N_4703);
nor U5964 (N_5964,N_4254,N_4348);
or U5965 (N_5965,N_4894,N_4314);
or U5966 (N_5966,N_4302,N_4280);
or U5967 (N_5967,N_4623,N_4317);
and U5968 (N_5968,N_4528,N_4504);
nand U5969 (N_5969,N_4146,N_4448);
xor U5970 (N_5970,N_4856,N_4520);
nor U5971 (N_5971,N_4756,N_4701);
nand U5972 (N_5972,N_4207,N_4567);
and U5973 (N_5973,N_4573,N_4686);
or U5974 (N_5974,N_4211,N_4516);
and U5975 (N_5975,N_4086,N_4605);
nand U5976 (N_5976,N_4734,N_4680);
or U5977 (N_5977,N_4315,N_4538);
or U5978 (N_5978,N_4440,N_4324);
nor U5979 (N_5979,N_4568,N_4025);
nand U5980 (N_5980,N_4543,N_4477);
or U5981 (N_5981,N_4098,N_4236);
nor U5982 (N_5982,N_4165,N_4421);
or U5983 (N_5983,N_4923,N_4497);
and U5984 (N_5984,N_4250,N_4147);
nor U5985 (N_5985,N_4154,N_4892);
or U5986 (N_5986,N_4092,N_4185);
or U5987 (N_5987,N_4559,N_4382);
and U5988 (N_5988,N_4409,N_4442);
nor U5989 (N_5989,N_4630,N_4545);
or U5990 (N_5990,N_4519,N_4093);
and U5991 (N_5991,N_4792,N_4276);
or U5992 (N_5992,N_4655,N_4799);
or U5993 (N_5993,N_4494,N_4757);
nand U5994 (N_5994,N_4306,N_4342);
or U5995 (N_5995,N_4102,N_4752);
nor U5996 (N_5996,N_4602,N_4779);
and U5997 (N_5997,N_4847,N_4162);
nor U5998 (N_5998,N_4677,N_4371);
nor U5999 (N_5999,N_4049,N_4403);
or U6000 (N_6000,N_5276,N_5088);
and U6001 (N_6001,N_5178,N_5454);
nand U6002 (N_6002,N_5445,N_5770);
nor U6003 (N_6003,N_5412,N_5760);
nand U6004 (N_6004,N_5366,N_5346);
nand U6005 (N_6005,N_5420,N_5994);
and U6006 (N_6006,N_5391,N_5958);
and U6007 (N_6007,N_5358,N_5004);
nand U6008 (N_6008,N_5446,N_5064);
or U6009 (N_6009,N_5757,N_5462);
and U6010 (N_6010,N_5525,N_5006);
or U6011 (N_6011,N_5061,N_5865);
nor U6012 (N_6012,N_5126,N_5599);
nor U6013 (N_6013,N_5794,N_5014);
and U6014 (N_6014,N_5233,N_5259);
or U6015 (N_6015,N_5904,N_5452);
and U6016 (N_6016,N_5868,N_5364);
nor U6017 (N_6017,N_5010,N_5931);
xnor U6018 (N_6018,N_5636,N_5155);
and U6019 (N_6019,N_5830,N_5813);
xor U6020 (N_6020,N_5734,N_5221);
nor U6021 (N_6021,N_5528,N_5068);
and U6022 (N_6022,N_5102,N_5226);
nor U6023 (N_6023,N_5993,N_5926);
nor U6024 (N_6024,N_5437,N_5078);
xnor U6025 (N_6025,N_5207,N_5218);
and U6026 (N_6026,N_5209,N_5272);
or U6027 (N_6027,N_5918,N_5369);
nor U6028 (N_6028,N_5986,N_5568);
nor U6029 (N_6029,N_5562,N_5302);
nor U6030 (N_6030,N_5729,N_5516);
nor U6031 (N_6031,N_5312,N_5775);
and U6032 (N_6032,N_5878,N_5638);
or U6033 (N_6033,N_5845,N_5159);
and U6034 (N_6034,N_5786,N_5717);
nand U6035 (N_6035,N_5566,N_5778);
nor U6036 (N_6036,N_5246,N_5242);
or U6037 (N_6037,N_5811,N_5493);
nor U6038 (N_6038,N_5457,N_5721);
or U6039 (N_6039,N_5058,N_5506);
and U6040 (N_6040,N_5213,N_5381);
and U6041 (N_6041,N_5645,N_5376);
or U6042 (N_6042,N_5664,N_5567);
xnor U6043 (N_6043,N_5923,N_5572);
or U6044 (N_6044,N_5417,N_5719);
nand U6045 (N_6045,N_5237,N_5486);
and U6046 (N_6046,N_5753,N_5593);
or U6047 (N_6047,N_5428,N_5507);
and U6048 (N_6048,N_5948,N_5955);
nand U6049 (N_6049,N_5468,N_5589);
or U6050 (N_6050,N_5470,N_5192);
or U6051 (N_6051,N_5502,N_5125);
and U6052 (N_6052,N_5592,N_5025);
or U6053 (N_6053,N_5530,N_5034);
and U6054 (N_6054,N_5885,N_5066);
nand U6055 (N_6055,N_5017,N_5890);
or U6056 (N_6056,N_5810,N_5691);
nand U6057 (N_6057,N_5104,N_5804);
or U6058 (N_6058,N_5925,N_5084);
and U6059 (N_6059,N_5657,N_5617);
nor U6060 (N_6060,N_5888,N_5090);
nor U6061 (N_6061,N_5724,N_5011);
nor U6062 (N_6062,N_5912,N_5311);
and U6063 (N_6063,N_5114,N_5487);
or U6064 (N_6064,N_5602,N_5712);
and U6065 (N_6065,N_5124,N_5135);
nand U6066 (N_6066,N_5190,N_5863);
nor U6067 (N_6067,N_5012,N_5464);
or U6068 (N_6068,N_5591,N_5901);
or U6069 (N_6069,N_5151,N_5648);
or U6070 (N_6070,N_5386,N_5429);
nor U6071 (N_6071,N_5939,N_5536);
nor U6072 (N_6072,N_5387,N_5363);
and U6073 (N_6073,N_5289,N_5979);
or U6074 (N_6074,N_5920,N_5158);
xor U6075 (N_6075,N_5057,N_5937);
xor U6076 (N_6076,N_5582,N_5651);
nor U6077 (N_6077,N_5320,N_5248);
nand U6078 (N_6078,N_5324,N_5145);
or U6079 (N_6079,N_5326,N_5230);
nand U6080 (N_6080,N_5534,N_5328);
or U6081 (N_6081,N_5876,N_5570);
nand U6082 (N_6082,N_5623,N_5492);
and U6083 (N_6083,N_5755,N_5726);
nor U6084 (N_6084,N_5673,N_5267);
and U6085 (N_6085,N_5989,N_5401);
nand U6086 (N_6086,N_5569,N_5303);
nor U6087 (N_6087,N_5508,N_5288);
xor U6088 (N_6088,N_5577,N_5730);
and U6089 (N_6089,N_5718,N_5667);
xnor U6090 (N_6090,N_5972,N_5640);
and U6091 (N_6091,N_5783,N_5161);
or U6092 (N_6092,N_5800,N_5587);
nor U6093 (N_6093,N_5849,N_5060);
nand U6094 (N_6094,N_5173,N_5344);
nand U6095 (N_6095,N_5130,N_5910);
xnor U6096 (N_6096,N_5764,N_5030);
nand U6097 (N_6097,N_5037,N_5893);
xnor U6098 (N_6098,N_5273,N_5999);
xor U6099 (N_6099,N_5574,N_5015);
xnor U6100 (N_6100,N_5922,N_5049);
nand U6101 (N_6101,N_5152,N_5002);
and U6102 (N_6102,N_5678,N_5216);
or U6103 (N_6103,N_5414,N_5463);
and U6104 (N_6104,N_5631,N_5991);
nor U6105 (N_6105,N_5785,N_5440);
nand U6106 (N_6106,N_5857,N_5708);
nand U6107 (N_6107,N_5504,N_5194);
xnor U6108 (N_6108,N_5399,N_5789);
nand U6109 (N_6109,N_5204,N_5756);
and U6110 (N_6110,N_5711,N_5828);
nor U6111 (N_6111,N_5716,N_5984);
nand U6112 (N_6112,N_5680,N_5983);
and U6113 (N_6113,N_5634,N_5632);
or U6114 (N_6114,N_5908,N_5879);
or U6115 (N_6115,N_5982,N_5129);
and U6116 (N_6116,N_5685,N_5681);
xnor U6117 (N_6117,N_5515,N_5971);
xnor U6118 (N_6118,N_5117,N_5059);
and U6119 (N_6119,N_5367,N_5086);
or U6120 (N_6120,N_5927,N_5001);
nand U6121 (N_6121,N_5843,N_5545);
nand U6122 (N_6122,N_5877,N_5539);
and U6123 (N_6123,N_5278,N_5028);
nor U6124 (N_6124,N_5250,N_5781);
nand U6125 (N_6125,N_5924,N_5873);
nand U6126 (N_6126,N_5389,N_5024);
and U6127 (N_6127,N_5674,N_5662);
and U6128 (N_6128,N_5338,N_5720);
and U6129 (N_6129,N_5820,N_5222);
or U6130 (N_6130,N_5047,N_5089);
and U6131 (N_6131,N_5180,N_5336);
nor U6132 (N_6132,N_5296,N_5062);
nor U6133 (N_6133,N_5601,N_5985);
and U6134 (N_6134,N_5436,N_5294);
xnor U6135 (N_6135,N_5600,N_5043);
or U6136 (N_6136,N_5342,N_5175);
and U6137 (N_6137,N_5777,N_5941);
nand U6138 (N_6138,N_5481,N_5735);
xor U6139 (N_6139,N_5263,N_5141);
and U6140 (N_6140,N_5837,N_5398);
nand U6141 (N_6141,N_5966,N_5395);
and U6142 (N_6142,N_5167,N_5531);
xnor U6143 (N_6143,N_5279,N_5021);
xnor U6144 (N_6144,N_5578,N_5065);
xor U6145 (N_6145,N_5921,N_5622);
nand U6146 (N_6146,N_5836,N_5038);
xnor U6147 (N_6147,N_5191,N_5643);
or U6148 (N_6148,N_5693,N_5829);
and U6149 (N_6149,N_5476,N_5677);
and U6150 (N_6150,N_5103,N_5430);
or U6151 (N_6151,N_5671,N_5360);
nand U6152 (N_6152,N_5241,N_5073);
nor U6153 (N_6153,N_5611,N_5082);
and U6154 (N_6154,N_5236,N_5461);
or U6155 (N_6155,N_5140,N_5650);
nand U6156 (N_6156,N_5198,N_5579);
xor U6157 (N_6157,N_5251,N_5137);
and U6158 (N_6158,N_5413,N_5256);
or U6159 (N_6159,N_5313,N_5113);
nand U6160 (N_6160,N_5070,N_5348);
nor U6161 (N_6161,N_5654,N_5659);
and U6162 (N_6162,N_5598,N_5826);
xnor U6163 (N_6163,N_5505,N_5975);
or U6164 (N_6164,N_5341,N_5844);
xor U6165 (N_6165,N_5548,N_5040);
nand U6166 (N_6166,N_5776,N_5701);
nor U6167 (N_6167,N_5423,N_5479);
and U6168 (N_6168,N_5620,N_5425);
or U6169 (N_6169,N_5854,N_5707);
or U6170 (N_6170,N_5238,N_5254);
nand U6171 (N_6171,N_5408,N_5887);
or U6172 (N_6172,N_5377,N_5963);
xor U6173 (N_6173,N_5833,N_5694);
nor U6174 (N_6174,N_5968,N_5848);
nand U6175 (N_6175,N_5977,N_5980);
xnor U6176 (N_6176,N_5016,N_5343);
nand U6177 (N_6177,N_5831,N_5818);
or U6178 (N_6178,N_5146,N_5488);
nor U6179 (N_6179,N_5390,N_5660);
and U6180 (N_6180,N_5003,N_5882);
or U6181 (N_6181,N_5590,N_5200);
nand U6182 (N_6182,N_5339,N_5450);
nand U6183 (N_6183,N_5766,N_5957);
nor U6184 (N_6184,N_5841,N_5079);
nand U6185 (N_6185,N_5610,N_5409);
or U6186 (N_6186,N_5281,N_5944);
and U6187 (N_6187,N_5415,N_5959);
nand U6188 (N_6188,N_5867,N_5471);
nand U6189 (N_6189,N_5754,N_5935);
nor U6190 (N_6190,N_5150,N_5261);
or U6191 (N_6191,N_5709,N_5499);
nand U6192 (N_6192,N_5297,N_5337);
and U6193 (N_6193,N_5350,N_5112);
nor U6194 (N_6194,N_5370,N_5223);
nor U6195 (N_6195,N_5949,N_5048);
xor U6196 (N_6196,N_5235,N_5981);
or U6197 (N_6197,N_5228,N_5309);
and U6198 (N_6198,N_5635,N_5700);
and U6199 (N_6199,N_5584,N_5005);
nor U6200 (N_6200,N_5875,N_5298);
or U6201 (N_6201,N_5380,N_5052);
and U6202 (N_6202,N_5892,N_5886);
xnor U6203 (N_6203,N_5306,N_5606);
xnor U6204 (N_6204,N_5356,N_5434);
or U6205 (N_6205,N_5771,N_5675);
and U6206 (N_6206,N_5688,N_5029);
and U6207 (N_6207,N_5243,N_5856);
and U6208 (N_6208,N_5624,N_5746);
nor U6209 (N_6209,N_5109,N_5551);
xor U6210 (N_6210,N_5115,N_5484);
or U6211 (N_6211,N_5575,N_5197);
or U6212 (N_6212,N_5092,N_5116);
and U6213 (N_6213,N_5858,N_5665);
or U6214 (N_6214,N_5774,N_5422);
or U6215 (N_6215,N_5123,N_5407);
and U6216 (N_6216,N_5214,N_5588);
nor U6217 (N_6217,N_5862,N_5449);
nor U6218 (N_6218,N_5613,N_5133);
xnor U6219 (N_6219,N_5809,N_5768);
nor U6220 (N_6220,N_5308,N_5797);
nand U6221 (N_6221,N_5332,N_5704);
and U6222 (N_6222,N_5725,N_5368);
nor U6223 (N_6223,N_5603,N_5523);
or U6224 (N_6224,N_5521,N_5345);
nor U6225 (N_6225,N_5518,N_5458);
nor U6226 (N_6226,N_5105,N_5748);
nand U6227 (N_6227,N_5046,N_5318);
or U6228 (N_6228,N_5555,N_5814);
nand U6229 (N_6229,N_5072,N_5633);
or U6230 (N_6230,N_5134,N_5576);
xnor U6231 (N_6231,N_5396,N_5702);
or U6232 (N_6232,N_5444,N_5581);
and U6233 (N_6233,N_5615,N_5639);
nand U6234 (N_6234,N_5619,N_5542);
and U6235 (N_6235,N_5362,N_5162);
and U6236 (N_6236,N_5751,N_5965);
nand U6237 (N_6237,N_5535,N_5988);
nor U6238 (N_6238,N_5397,N_5628);
nor U6239 (N_6239,N_5782,N_5400);
and U6240 (N_6240,N_5189,N_5911);
nor U6241 (N_6241,N_5375,N_5268);
or U6242 (N_6242,N_5871,N_5987);
nand U6243 (N_6243,N_5179,N_5032);
and U6244 (N_6244,N_5008,N_5497);
xnor U6245 (N_6245,N_5322,N_5524);
and U6246 (N_6246,N_5050,N_5282);
nand U6247 (N_6247,N_5443,N_5177);
and U6248 (N_6248,N_5442,N_5496);
and U6249 (N_6249,N_5127,N_5169);
nand U6250 (N_6250,N_5349,N_5299);
and U6251 (N_6251,N_5790,N_5883);
nand U6252 (N_6252,N_5874,N_5802);
nand U6253 (N_6253,N_5745,N_5821);
or U6254 (N_6254,N_5494,N_5347);
or U6255 (N_6255,N_5131,N_5930);
and U6256 (N_6256,N_5365,N_5946);
and U6257 (N_6257,N_5621,N_5947);
nor U6258 (N_6258,N_5096,N_5201);
or U6259 (N_6259,N_5128,N_5148);
nor U6260 (N_6260,N_5439,N_5459);
nand U6261 (N_6261,N_5609,N_5938);
or U6262 (N_6262,N_5077,N_5477);
or U6263 (N_6263,N_5315,N_5792);
nor U6264 (N_6264,N_5331,N_5284);
nor U6265 (N_6265,N_5041,N_5835);
nand U6266 (N_6266,N_5646,N_5889);
nor U6267 (N_6267,N_5329,N_5174);
nand U6268 (N_6268,N_5679,N_5739);
and U6269 (N_6269,N_5998,N_5954);
or U6270 (N_6270,N_5325,N_5630);
nor U6271 (N_6271,N_5182,N_5618);
or U6272 (N_6272,N_5163,N_5512);
nand U6273 (N_6273,N_5549,N_5193);
nand U6274 (N_6274,N_5027,N_5184);
or U6275 (N_6275,N_5157,N_5265);
nor U6276 (N_6276,N_5663,N_5894);
or U6277 (N_6277,N_5044,N_5456);
xnor U6278 (N_6278,N_5208,N_5895);
nand U6279 (N_6279,N_5661,N_5293);
nand U6280 (N_6280,N_5101,N_5727);
nand U6281 (N_6281,N_5817,N_5107);
or U6282 (N_6282,N_5394,N_5608);
nand U6283 (N_6283,N_5563,N_5733);
nor U6284 (N_6284,N_5206,N_5406);
xor U6285 (N_6285,N_5290,N_5538);
and U6286 (N_6286,N_5300,N_5168);
or U6287 (N_6287,N_5652,N_5378);
nor U6288 (N_6288,N_5546,N_5763);
xor U6289 (N_6289,N_5035,N_5352);
nor U6290 (N_6290,N_5232,N_5249);
or U6291 (N_6291,N_5383,N_5564);
nor U6292 (N_6292,N_5418,N_5909);
or U6293 (N_6293,N_5698,N_5353);
nor U6294 (N_6294,N_5153,N_5808);
nor U6295 (N_6295,N_5132,N_5950);
xnor U6296 (N_6296,N_5503,N_5188);
or U6297 (N_6297,N_5310,N_5424);
nor U6298 (N_6298,N_5996,N_5929);
xor U6299 (N_6299,N_5847,N_5314);
xnor U6300 (N_6300,N_5093,N_5710);
nand U6301 (N_6301,N_5327,N_5713);
nor U6302 (N_6302,N_5286,N_5485);
nor U6303 (N_6303,N_5779,N_5795);
nand U6304 (N_6304,N_5697,N_5585);
nor U6305 (N_6305,N_5834,N_5953);
and U6306 (N_6306,N_5703,N_5832);
and U6307 (N_6307,N_5211,N_5421);
nand U6308 (N_6308,N_5732,N_5758);
nor U6309 (N_6309,N_5683,N_5340);
xor U6310 (N_6310,N_5670,N_5898);
nand U6311 (N_6311,N_5840,N_5740);
xnor U6312 (N_6312,N_5627,N_5851);
or U6313 (N_6313,N_5405,N_5304);
nand U6314 (N_6314,N_5081,N_5166);
nand U6315 (N_6315,N_5260,N_5100);
or U6316 (N_6316,N_5956,N_5203);
xnor U6317 (N_6317,N_5097,N_5372);
nand U6318 (N_6318,N_5769,N_5687);
and U6319 (N_6319,N_5234,N_5543);
or U6320 (N_6320,N_5335,N_5447);
and U6321 (N_6321,N_5007,N_5385);
nor U6322 (N_6322,N_5076,N_5045);
xor U6323 (N_6323,N_5672,N_5165);
nand U6324 (N_6324,N_5765,N_5692);
nand U6325 (N_6325,N_5815,N_5743);
xnor U6326 (N_6326,N_5772,N_5520);
nor U6327 (N_6327,N_5571,N_5215);
xor U6328 (N_6328,N_5558,N_5705);
and U6329 (N_6329,N_5527,N_5491);
nor U6330 (N_6330,N_5000,N_5074);
or U6331 (N_6331,N_5316,N_5108);
nand U6332 (N_6332,N_5605,N_5501);
nor U6333 (N_6333,N_5067,N_5351);
nor U6334 (N_6334,N_5056,N_5791);
nor U6335 (N_6335,N_5480,N_5554);
nor U6336 (N_6336,N_5411,N_5855);
nand U6337 (N_6337,N_5747,N_5714);
or U6338 (N_6338,N_5750,N_5827);
and U6339 (N_6339,N_5960,N_5839);
or U6340 (N_6340,N_5269,N_5160);
and U6341 (N_6341,N_5026,N_5547);
nor U6342 (N_6342,N_5036,N_5870);
or U6343 (N_6343,N_5181,N_5690);
and U6344 (N_6344,N_5934,N_5942);
nor U6345 (N_6345,N_5402,N_5916);
and U6346 (N_6346,N_5932,N_5974);
nand U6347 (N_6347,N_5388,N_5951);
and U6348 (N_6348,N_5280,N_5244);
or U6349 (N_6349,N_5881,N_5872);
nand U6350 (N_6350,N_5597,N_5292);
and U6351 (N_6351,N_5333,N_5098);
nand U6352 (N_6352,N_5842,N_5187);
xor U6353 (N_6353,N_5513,N_5807);
nand U6354 (N_6354,N_5330,N_5933);
nor U6355 (N_6355,N_5906,N_5202);
nand U6356 (N_6356,N_5099,N_5051);
or U6357 (N_6357,N_5964,N_5039);
or U6358 (N_6358,N_5361,N_5095);
or U6359 (N_6359,N_5453,N_5668);
and U6360 (N_6360,N_5451,N_5642);
or U6361 (N_6361,N_5416,N_5533);
nor U6362 (N_6362,N_5122,N_5357);
and U6363 (N_6363,N_5738,N_5438);
nand U6364 (N_6364,N_5156,N_5225);
nor U6365 (N_6365,N_5149,N_5196);
and U6366 (N_6366,N_5291,N_5441);
or U6367 (N_6367,N_5860,N_5616);
or U6368 (N_6368,N_5580,N_5255);
nor U6369 (N_6369,N_5915,N_5728);
or U6370 (N_6370,N_5419,N_5928);
nor U6371 (N_6371,N_5607,N_5559);
xor U6372 (N_6372,N_5379,N_5120);
nor U6373 (N_6373,N_5147,N_5253);
nand U6374 (N_6374,N_5803,N_5796);
nand U6375 (N_6375,N_5371,N_5426);
and U6376 (N_6376,N_5392,N_5219);
and U6377 (N_6377,N_5220,N_5943);
and U6378 (N_6378,N_5354,N_5655);
and U6379 (N_6379,N_5676,N_5583);
and U6380 (N_6380,N_5245,N_5699);
nand U6381 (N_6381,N_5071,N_5784);
nor U6382 (N_6382,N_5695,N_5798);
and U6383 (N_6383,N_5277,N_5239);
nor U6384 (N_6384,N_5247,N_5864);
nor U6385 (N_6385,N_5307,N_5271);
nor U6386 (N_6386,N_5185,N_5541);
nor U6387 (N_6387,N_5094,N_5227);
or U6388 (N_6388,N_5121,N_5500);
or U6389 (N_6389,N_5788,N_5472);
or U6390 (N_6390,N_5522,N_5106);
nor U6391 (N_6391,N_5478,N_5475);
nand U6392 (N_6392,N_5962,N_5722);
nand U6393 (N_6393,N_5069,N_5940);
nand U6394 (N_6394,N_5715,N_5767);
or U6395 (N_6395,N_5460,N_5517);
nand U6396 (N_6396,N_5080,N_5427);
or U6397 (N_6397,N_5305,N_5301);
or U6398 (N_6398,N_5264,N_5509);
nand U6399 (N_6399,N_5838,N_5969);
and U6400 (N_6400,N_5596,N_5033);
and U6401 (N_6401,N_5917,N_5262);
and U6402 (N_6402,N_5176,N_5142);
xnor U6403 (N_6403,N_5164,N_5819);
xor U6404 (N_6404,N_5706,N_5139);
nand U6405 (N_6405,N_5075,N_5224);
nand U6406 (N_6406,N_5022,N_5474);
xnor U6407 (N_6407,N_5612,N_5055);
and U6408 (N_6408,N_5321,N_5270);
or U6409 (N_6409,N_5853,N_5111);
and U6410 (N_6410,N_5519,N_5274);
and U6411 (N_6411,N_5323,N_5295);
or U6412 (N_6412,N_5283,N_5550);
nand U6413 (N_6413,N_5850,N_5063);
or U6414 (N_6414,N_5658,N_5656);
nor U6415 (N_6415,N_5054,N_5317);
or U6416 (N_6416,N_5552,N_5087);
or U6417 (N_6417,N_5467,N_5759);
or U6418 (N_6418,N_5689,N_5556);
or U6419 (N_6419,N_5085,N_5171);
xor U6420 (N_6420,N_5240,N_5952);
nand U6421 (N_6421,N_5641,N_5604);
or U6422 (N_6422,N_5919,N_5170);
nand U6423 (N_6423,N_5905,N_5540);
xnor U6424 (N_6424,N_5644,N_5696);
or U6425 (N_6425,N_5978,N_5629);
or U6426 (N_6426,N_5009,N_5976);
or U6427 (N_6427,N_5205,N_5560);
or U6428 (N_6428,N_5172,N_5465);
and U6429 (N_6429,N_5537,N_5666);
or U6430 (N_6430,N_5359,N_5565);
nor U6431 (N_6431,N_5744,N_5433);
nor U6432 (N_6432,N_5532,N_5053);
and U6433 (N_6433,N_5019,N_5586);
and U6434 (N_6434,N_5773,N_5403);
nor U6435 (N_6435,N_5490,N_5903);
and U6436 (N_6436,N_5762,N_5897);
nor U6437 (N_6437,N_5899,N_5186);
nor U6438 (N_6438,N_5824,N_5900);
nor U6439 (N_6439,N_5780,N_5801);
or U6440 (N_6440,N_5431,N_5143);
nand U6441 (N_6441,N_5787,N_5266);
nor U6442 (N_6442,N_5514,N_5020);
nor U6443 (N_6443,N_5119,N_5374);
nor U6444 (N_6444,N_5995,N_5432);
nand U6445 (N_6445,N_5285,N_5510);
and U6446 (N_6446,N_5884,N_5553);
nor U6447 (N_6447,N_5287,N_5217);
or U6448 (N_6448,N_5455,N_5384);
nand U6449 (N_6449,N_5031,N_5210);
nor U6450 (N_6450,N_5752,N_5682);
and U6451 (N_6451,N_5866,N_5625);
nor U6452 (N_6452,N_5823,N_5183);
or U6453 (N_6453,N_5669,N_5647);
nand U6454 (N_6454,N_5936,N_5653);
xor U6455 (N_6455,N_5907,N_5257);
nand U6456 (N_6456,N_5880,N_5258);
and U6457 (N_6457,N_5561,N_5448);
nor U6458 (N_6458,N_5466,N_5118);
and U6459 (N_6459,N_5355,N_5869);
nor U6460 (N_6460,N_5806,N_5483);
xor U6461 (N_6461,N_5961,N_5846);
or U6462 (N_6462,N_5825,N_5489);
or U6463 (N_6463,N_5761,N_5473);
nor U6464 (N_6464,N_5812,N_5741);
nand U6465 (N_6465,N_5231,N_5731);
nand U6466 (N_6466,N_5637,N_5737);
nand U6467 (N_6467,N_5091,N_5018);
and U6468 (N_6468,N_5042,N_5435);
or U6469 (N_6469,N_5154,N_5229);
xnor U6470 (N_6470,N_5852,N_5023);
nand U6471 (N_6471,N_5393,N_5382);
and U6472 (N_6472,N_5110,N_5945);
nor U6473 (N_6473,N_5373,N_5723);
nor U6474 (N_6474,N_5212,N_5199);
nor U6475 (N_6475,N_5973,N_5799);
and U6476 (N_6476,N_5902,N_5970);
xor U6477 (N_6477,N_5822,N_5404);
or U6478 (N_6478,N_5742,N_5793);
and U6479 (N_6479,N_5482,N_5896);
nor U6480 (N_6480,N_5967,N_5511);
and U6481 (N_6481,N_5083,N_5686);
or U6482 (N_6482,N_5749,N_5861);
xor U6483 (N_6483,N_5410,N_5891);
or U6484 (N_6484,N_5626,N_5992);
nor U6485 (N_6485,N_5544,N_5805);
or U6486 (N_6486,N_5469,N_5138);
or U6487 (N_6487,N_5816,N_5319);
and U6488 (N_6488,N_5913,N_5594);
and U6489 (N_6489,N_5252,N_5859);
nand U6490 (N_6490,N_5914,N_5334);
xnor U6491 (N_6491,N_5649,N_5495);
nand U6492 (N_6492,N_5990,N_5573);
nor U6493 (N_6493,N_5013,N_5684);
or U6494 (N_6494,N_5498,N_5195);
or U6495 (N_6495,N_5595,N_5275);
nor U6496 (N_6496,N_5529,N_5557);
nor U6497 (N_6497,N_5614,N_5144);
xor U6498 (N_6498,N_5997,N_5736);
nand U6499 (N_6499,N_5526,N_5136);
xor U6500 (N_6500,N_5266,N_5576);
nand U6501 (N_6501,N_5085,N_5322);
nand U6502 (N_6502,N_5501,N_5751);
nor U6503 (N_6503,N_5397,N_5711);
and U6504 (N_6504,N_5925,N_5634);
xnor U6505 (N_6505,N_5992,N_5760);
nand U6506 (N_6506,N_5629,N_5396);
or U6507 (N_6507,N_5122,N_5987);
or U6508 (N_6508,N_5866,N_5972);
nand U6509 (N_6509,N_5902,N_5448);
and U6510 (N_6510,N_5543,N_5257);
nor U6511 (N_6511,N_5578,N_5801);
or U6512 (N_6512,N_5088,N_5582);
and U6513 (N_6513,N_5953,N_5220);
and U6514 (N_6514,N_5675,N_5861);
or U6515 (N_6515,N_5245,N_5060);
and U6516 (N_6516,N_5446,N_5989);
nand U6517 (N_6517,N_5011,N_5179);
nand U6518 (N_6518,N_5376,N_5738);
or U6519 (N_6519,N_5885,N_5193);
nor U6520 (N_6520,N_5172,N_5375);
nor U6521 (N_6521,N_5282,N_5531);
and U6522 (N_6522,N_5482,N_5425);
nand U6523 (N_6523,N_5802,N_5121);
xor U6524 (N_6524,N_5358,N_5676);
nor U6525 (N_6525,N_5288,N_5820);
nor U6526 (N_6526,N_5501,N_5806);
xor U6527 (N_6527,N_5593,N_5129);
and U6528 (N_6528,N_5294,N_5463);
xor U6529 (N_6529,N_5265,N_5111);
or U6530 (N_6530,N_5411,N_5988);
or U6531 (N_6531,N_5736,N_5926);
nand U6532 (N_6532,N_5794,N_5191);
or U6533 (N_6533,N_5745,N_5709);
or U6534 (N_6534,N_5208,N_5576);
nor U6535 (N_6535,N_5591,N_5886);
or U6536 (N_6536,N_5171,N_5020);
and U6537 (N_6537,N_5670,N_5145);
or U6538 (N_6538,N_5620,N_5612);
or U6539 (N_6539,N_5576,N_5158);
or U6540 (N_6540,N_5629,N_5451);
nand U6541 (N_6541,N_5557,N_5225);
or U6542 (N_6542,N_5873,N_5779);
nor U6543 (N_6543,N_5048,N_5074);
nor U6544 (N_6544,N_5486,N_5983);
and U6545 (N_6545,N_5749,N_5817);
nand U6546 (N_6546,N_5373,N_5974);
and U6547 (N_6547,N_5090,N_5428);
and U6548 (N_6548,N_5659,N_5717);
or U6549 (N_6549,N_5530,N_5552);
and U6550 (N_6550,N_5245,N_5362);
nor U6551 (N_6551,N_5135,N_5648);
nor U6552 (N_6552,N_5073,N_5825);
nand U6553 (N_6553,N_5171,N_5603);
nor U6554 (N_6554,N_5919,N_5727);
xor U6555 (N_6555,N_5678,N_5945);
or U6556 (N_6556,N_5368,N_5886);
or U6557 (N_6557,N_5626,N_5963);
and U6558 (N_6558,N_5757,N_5179);
nand U6559 (N_6559,N_5256,N_5509);
xnor U6560 (N_6560,N_5867,N_5098);
nor U6561 (N_6561,N_5313,N_5849);
xor U6562 (N_6562,N_5930,N_5031);
or U6563 (N_6563,N_5646,N_5553);
or U6564 (N_6564,N_5616,N_5634);
and U6565 (N_6565,N_5994,N_5045);
nor U6566 (N_6566,N_5938,N_5298);
nor U6567 (N_6567,N_5508,N_5749);
or U6568 (N_6568,N_5865,N_5584);
or U6569 (N_6569,N_5977,N_5463);
nand U6570 (N_6570,N_5120,N_5378);
nor U6571 (N_6571,N_5819,N_5808);
or U6572 (N_6572,N_5003,N_5732);
nor U6573 (N_6573,N_5918,N_5247);
or U6574 (N_6574,N_5081,N_5541);
or U6575 (N_6575,N_5432,N_5211);
and U6576 (N_6576,N_5520,N_5940);
xor U6577 (N_6577,N_5334,N_5961);
nand U6578 (N_6578,N_5328,N_5711);
or U6579 (N_6579,N_5828,N_5521);
or U6580 (N_6580,N_5118,N_5157);
xor U6581 (N_6581,N_5924,N_5961);
or U6582 (N_6582,N_5363,N_5425);
nand U6583 (N_6583,N_5017,N_5699);
or U6584 (N_6584,N_5596,N_5471);
or U6585 (N_6585,N_5230,N_5404);
or U6586 (N_6586,N_5226,N_5773);
or U6587 (N_6587,N_5687,N_5507);
xor U6588 (N_6588,N_5918,N_5618);
nor U6589 (N_6589,N_5758,N_5135);
nand U6590 (N_6590,N_5149,N_5653);
or U6591 (N_6591,N_5373,N_5497);
nor U6592 (N_6592,N_5290,N_5960);
or U6593 (N_6593,N_5835,N_5305);
and U6594 (N_6594,N_5154,N_5477);
nor U6595 (N_6595,N_5430,N_5064);
or U6596 (N_6596,N_5894,N_5702);
nand U6597 (N_6597,N_5751,N_5230);
xnor U6598 (N_6598,N_5483,N_5220);
nor U6599 (N_6599,N_5940,N_5614);
nand U6600 (N_6600,N_5291,N_5681);
or U6601 (N_6601,N_5900,N_5283);
or U6602 (N_6602,N_5220,N_5792);
and U6603 (N_6603,N_5316,N_5174);
and U6604 (N_6604,N_5488,N_5825);
and U6605 (N_6605,N_5516,N_5168);
nand U6606 (N_6606,N_5513,N_5583);
nand U6607 (N_6607,N_5792,N_5802);
nand U6608 (N_6608,N_5178,N_5998);
nor U6609 (N_6609,N_5431,N_5707);
and U6610 (N_6610,N_5076,N_5131);
and U6611 (N_6611,N_5969,N_5783);
nor U6612 (N_6612,N_5418,N_5491);
or U6613 (N_6613,N_5208,N_5247);
and U6614 (N_6614,N_5570,N_5452);
nand U6615 (N_6615,N_5634,N_5397);
and U6616 (N_6616,N_5866,N_5923);
nor U6617 (N_6617,N_5587,N_5348);
nand U6618 (N_6618,N_5206,N_5536);
xnor U6619 (N_6619,N_5815,N_5168);
xnor U6620 (N_6620,N_5683,N_5853);
nor U6621 (N_6621,N_5611,N_5932);
and U6622 (N_6622,N_5526,N_5811);
nor U6623 (N_6623,N_5066,N_5098);
or U6624 (N_6624,N_5491,N_5828);
or U6625 (N_6625,N_5138,N_5359);
nand U6626 (N_6626,N_5768,N_5510);
nor U6627 (N_6627,N_5561,N_5829);
or U6628 (N_6628,N_5981,N_5158);
xnor U6629 (N_6629,N_5643,N_5239);
nor U6630 (N_6630,N_5259,N_5830);
nand U6631 (N_6631,N_5532,N_5141);
nor U6632 (N_6632,N_5560,N_5323);
nor U6633 (N_6633,N_5187,N_5208);
or U6634 (N_6634,N_5689,N_5200);
and U6635 (N_6635,N_5864,N_5166);
xor U6636 (N_6636,N_5241,N_5781);
or U6637 (N_6637,N_5016,N_5082);
nor U6638 (N_6638,N_5694,N_5266);
and U6639 (N_6639,N_5285,N_5882);
nand U6640 (N_6640,N_5741,N_5182);
nor U6641 (N_6641,N_5039,N_5562);
or U6642 (N_6642,N_5307,N_5316);
xor U6643 (N_6643,N_5935,N_5679);
xor U6644 (N_6644,N_5257,N_5314);
nor U6645 (N_6645,N_5319,N_5050);
nor U6646 (N_6646,N_5393,N_5159);
or U6647 (N_6647,N_5803,N_5337);
or U6648 (N_6648,N_5679,N_5830);
xor U6649 (N_6649,N_5631,N_5206);
and U6650 (N_6650,N_5549,N_5619);
or U6651 (N_6651,N_5588,N_5128);
xnor U6652 (N_6652,N_5770,N_5399);
or U6653 (N_6653,N_5186,N_5707);
xor U6654 (N_6654,N_5712,N_5861);
nand U6655 (N_6655,N_5379,N_5937);
nor U6656 (N_6656,N_5513,N_5531);
nor U6657 (N_6657,N_5076,N_5975);
nor U6658 (N_6658,N_5229,N_5557);
and U6659 (N_6659,N_5158,N_5630);
or U6660 (N_6660,N_5520,N_5051);
or U6661 (N_6661,N_5354,N_5425);
xor U6662 (N_6662,N_5939,N_5395);
and U6663 (N_6663,N_5515,N_5692);
nand U6664 (N_6664,N_5463,N_5475);
nand U6665 (N_6665,N_5995,N_5759);
and U6666 (N_6666,N_5783,N_5884);
xor U6667 (N_6667,N_5472,N_5343);
nand U6668 (N_6668,N_5654,N_5774);
or U6669 (N_6669,N_5580,N_5003);
and U6670 (N_6670,N_5287,N_5724);
or U6671 (N_6671,N_5968,N_5574);
or U6672 (N_6672,N_5474,N_5043);
nor U6673 (N_6673,N_5330,N_5792);
nand U6674 (N_6674,N_5695,N_5467);
and U6675 (N_6675,N_5561,N_5639);
nand U6676 (N_6676,N_5567,N_5519);
nand U6677 (N_6677,N_5586,N_5329);
nor U6678 (N_6678,N_5492,N_5450);
xor U6679 (N_6679,N_5622,N_5414);
and U6680 (N_6680,N_5441,N_5526);
and U6681 (N_6681,N_5842,N_5263);
nor U6682 (N_6682,N_5783,N_5766);
and U6683 (N_6683,N_5448,N_5678);
nand U6684 (N_6684,N_5855,N_5774);
or U6685 (N_6685,N_5633,N_5943);
and U6686 (N_6686,N_5499,N_5355);
or U6687 (N_6687,N_5144,N_5668);
nor U6688 (N_6688,N_5878,N_5838);
and U6689 (N_6689,N_5737,N_5361);
or U6690 (N_6690,N_5413,N_5636);
nor U6691 (N_6691,N_5843,N_5798);
xnor U6692 (N_6692,N_5258,N_5977);
nor U6693 (N_6693,N_5613,N_5511);
and U6694 (N_6694,N_5074,N_5054);
or U6695 (N_6695,N_5354,N_5789);
and U6696 (N_6696,N_5399,N_5269);
and U6697 (N_6697,N_5643,N_5977);
and U6698 (N_6698,N_5924,N_5091);
or U6699 (N_6699,N_5534,N_5613);
or U6700 (N_6700,N_5835,N_5912);
nor U6701 (N_6701,N_5509,N_5888);
nand U6702 (N_6702,N_5627,N_5841);
or U6703 (N_6703,N_5090,N_5434);
xor U6704 (N_6704,N_5452,N_5237);
nor U6705 (N_6705,N_5969,N_5222);
or U6706 (N_6706,N_5117,N_5124);
nor U6707 (N_6707,N_5561,N_5802);
or U6708 (N_6708,N_5705,N_5810);
nor U6709 (N_6709,N_5667,N_5897);
and U6710 (N_6710,N_5118,N_5786);
and U6711 (N_6711,N_5009,N_5722);
and U6712 (N_6712,N_5251,N_5036);
and U6713 (N_6713,N_5768,N_5498);
nand U6714 (N_6714,N_5235,N_5395);
nor U6715 (N_6715,N_5106,N_5428);
nor U6716 (N_6716,N_5386,N_5006);
and U6717 (N_6717,N_5628,N_5134);
and U6718 (N_6718,N_5355,N_5164);
and U6719 (N_6719,N_5997,N_5928);
nor U6720 (N_6720,N_5263,N_5018);
and U6721 (N_6721,N_5206,N_5555);
nand U6722 (N_6722,N_5043,N_5495);
nor U6723 (N_6723,N_5341,N_5504);
nand U6724 (N_6724,N_5391,N_5493);
or U6725 (N_6725,N_5506,N_5442);
and U6726 (N_6726,N_5387,N_5560);
nand U6727 (N_6727,N_5600,N_5160);
or U6728 (N_6728,N_5937,N_5595);
and U6729 (N_6729,N_5038,N_5375);
and U6730 (N_6730,N_5505,N_5592);
and U6731 (N_6731,N_5447,N_5535);
and U6732 (N_6732,N_5920,N_5518);
nor U6733 (N_6733,N_5050,N_5000);
nor U6734 (N_6734,N_5444,N_5400);
or U6735 (N_6735,N_5438,N_5726);
nor U6736 (N_6736,N_5841,N_5331);
nand U6737 (N_6737,N_5559,N_5954);
or U6738 (N_6738,N_5098,N_5579);
nor U6739 (N_6739,N_5639,N_5619);
nor U6740 (N_6740,N_5215,N_5556);
nand U6741 (N_6741,N_5197,N_5920);
or U6742 (N_6742,N_5750,N_5833);
nand U6743 (N_6743,N_5117,N_5030);
nand U6744 (N_6744,N_5020,N_5523);
nor U6745 (N_6745,N_5571,N_5695);
nor U6746 (N_6746,N_5284,N_5147);
nand U6747 (N_6747,N_5851,N_5430);
or U6748 (N_6748,N_5731,N_5086);
or U6749 (N_6749,N_5177,N_5336);
nand U6750 (N_6750,N_5262,N_5076);
nand U6751 (N_6751,N_5634,N_5300);
nand U6752 (N_6752,N_5163,N_5675);
nor U6753 (N_6753,N_5499,N_5871);
xor U6754 (N_6754,N_5198,N_5682);
nor U6755 (N_6755,N_5774,N_5019);
nor U6756 (N_6756,N_5216,N_5245);
and U6757 (N_6757,N_5634,N_5931);
or U6758 (N_6758,N_5955,N_5364);
nor U6759 (N_6759,N_5576,N_5938);
or U6760 (N_6760,N_5985,N_5803);
nor U6761 (N_6761,N_5338,N_5669);
nor U6762 (N_6762,N_5960,N_5647);
and U6763 (N_6763,N_5299,N_5075);
nand U6764 (N_6764,N_5165,N_5310);
nand U6765 (N_6765,N_5452,N_5678);
nor U6766 (N_6766,N_5144,N_5280);
or U6767 (N_6767,N_5732,N_5387);
xor U6768 (N_6768,N_5909,N_5760);
and U6769 (N_6769,N_5070,N_5424);
xor U6770 (N_6770,N_5286,N_5723);
and U6771 (N_6771,N_5061,N_5550);
and U6772 (N_6772,N_5674,N_5597);
or U6773 (N_6773,N_5497,N_5508);
and U6774 (N_6774,N_5666,N_5774);
nand U6775 (N_6775,N_5612,N_5305);
or U6776 (N_6776,N_5837,N_5040);
and U6777 (N_6777,N_5111,N_5961);
xor U6778 (N_6778,N_5795,N_5566);
nor U6779 (N_6779,N_5976,N_5604);
and U6780 (N_6780,N_5459,N_5249);
nand U6781 (N_6781,N_5363,N_5530);
xor U6782 (N_6782,N_5081,N_5885);
nand U6783 (N_6783,N_5842,N_5893);
or U6784 (N_6784,N_5597,N_5061);
or U6785 (N_6785,N_5001,N_5802);
and U6786 (N_6786,N_5712,N_5241);
xnor U6787 (N_6787,N_5694,N_5350);
and U6788 (N_6788,N_5101,N_5367);
nor U6789 (N_6789,N_5495,N_5499);
nand U6790 (N_6790,N_5137,N_5120);
nor U6791 (N_6791,N_5361,N_5824);
or U6792 (N_6792,N_5375,N_5276);
or U6793 (N_6793,N_5212,N_5155);
nor U6794 (N_6794,N_5614,N_5419);
and U6795 (N_6795,N_5971,N_5402);
nand U6796 (N_6796,N_5413,N_5045);
nor U6797 (N_6797,N_5527,N_5004);
nor U6798 (N_6798,N_5417,N_5774);
and U6799 (N_6799,N_5626,N_5162);
nor U6800 (N_6800,N_5738,N_5720);
xnor U6801 (N_6801,N_5399,N_5210);
or U6802 (N_6802,N_5358,N_5454);
and U6803 (N_6803,N_5748,N_5330);
nand U6804 (N_6804,N_5052,N_5078);
nand U6805 (N_6805,N_5339,N_5011);
xor U6806 (N_6806,N_5251,N_5618);
nand U6807 (N_6807,N_5015,N_5020);
xnor U6808 (N_6808,N_5881,N_5685);
or U6809 (N_6809,N_5763,N_5092);
nand U6810 (N_6810,N_5325,N_5110);
nand U6811 (N_6811,N_5861,N_5611);
nand U6812 (N_6812,N_5311,N_5017);
nor U6813 (N_6813,N_5268,N_5675);
nand U6814 (N_6814,N_5094,N_5012);
and U6815 (N_6815,N_5609,N_5266);
and U6816 (N_6816,N_5341,N_5508);
nor U6817 (N_6817,N_5529,N_5266);
and U6818 (N_6818,N_5982,N_5746);
and U6819 (N_6819,N_5486,N_5172);
xor U6820 (N_6820,N_5140,N_5341);
and U6821 (N_6821,N_5109,N_5016);
nand U6822 (N_6822,N_5766,N_5499);
xor U6823 (N_6823,N_5697,N_5063);
nand U6824 (N_6824,N_5723,N_5411);
nand U6825 (N_6825,N_5755,N_5673);
and U6826 (N_6826,N_5709,N_5125);
nand U6827 (N_6827,N_5771,N_5108);
nand U6828 (N_6828,N_5428,N_5982);
or U6829 (N_6829,N_5634,N_5980);
or U6830 (N_6830,N_5453,N_5661);
nand U6831 (N_6831,N_5805,N_5636);
nor U6832 (N_6832,N_5237,N_5705);
and U6833 (N_6833,N_5531,N_5688);
nor U6834 (N_6834,N_5985,N_5302);
and U6835 (N_6835,N_5644,N_5629);
nor U6836 (N_6836,N_5405,N_5496);
xnor U6837 (N_6837,N_5305,N_5672);
nor U6838 (N_6838,N_5977,N_5509);
nand U6839 (N_6839,N_5911,N_5457);
nor U6840 (N_6840,N_5472,N_5803);
nor U6841 (N_6841,N_5168,N_5893);
xor U6842 (N_6842,N_5599,N_5882);
or U6843 (N_6843,N_5496,N_5517);
or U6844 (N_6844,N_5730,N_5748);
nor U6845 (N_6845,N_5558,N_5735);
xor U6846 (N_6846,N_5667,N_5639);
nor U6847 (N_6847,N_5801,N_5696);
and U6848 (N_6848,N_5597,N_5255);
and U6849 (N_6849,N_5533,N_5409);
and U6850 (N_6850,N_5007,N_5699);
or U6851 (N_6851,N_5324,N_5736);
nor U6852 (N_6852,N_5545,N_5805);
or U6853 (N_6853,N_5461,N_5828);
and U6854 (N_6854,N_5021,N_5155);
nor U6855 (N_6855,N_5048,N_5985);
nor U6856 (N_6856,N_5717,N_5218);
xnor U6857 (N_6857,N_5155,N_5452);
nor U6858 (N_6858,N_5766,N_5261);
and U6859 (N_6859,N_5486,N_5655);
nand U6860 (N_6860,N_5227,N_5064);
nand U6861 (N_6861,N_5576,N_5118);
nor U6862 (N_6862,N_5489,N_5711);
nor U6863 (N_6863,N_5995,N_5441);
xor U6864 (N_6864,N_5326,N_5865);
or U6865 (N_6865,N_5839,N_5742);
nor U6866 (N_6866,N_5255,N_5475);
nand U6867 (N_6867,N_5174,N_5338);
nand U6868 (N_6868,N_5445,N_5968);
nor U6869 (N_6869,N_5338,N_5880);
or U6870 (N_6870,N_5883,N_5169);
or U6871 (N_6871,N_5941,N_5937);
nor U6872 (N_6872,N_5796,N_5012);
nand U6873 (N_6873,N_5300,N_5235);
or U6874 (N_6874,N_5165,N_5276);
nand U6875 (N_6875,N_5842,N_5520);
nand U6876 (N_6876,N_5294,N_5895);
nand U6877 (N_6877,N_5839,N_5145);
nand U6878 (N_6878,N_5659,N_5863);
or U6879 (N_6879,N_5785,N_5246);
and U6880 (N_6880,N_5179,N_5677);
nand U6881 (N_6881,N_5736,N_5605);
nor U6882 (N_6882,N_5826,N_5533);
nand U6883 (N_6883,N_5165,N_5980);
and U6884 (N_6884,N_5719,N_5810);
xnor U6885 (N_6885,N_5865,N_5301);
or U6886 (N_6886,N_5712,N_5274);
and U6887 (N_6887,N_5886,N_5561);
nor U6888 (N_6888,N_5981,N_5133);
nor U6889 (N_6889,N_5197,N_5864);
xor U6890 (N_6890,N_5127,N_5644);
and U6891 (N_6891,N_5024,N_5451);
or U6892 (N_6892,N_5024,N_5624);
and U6893 (N_6893,N_5749,N_5497);
nor U6894 (N_6894,N_5613,N_5650);
and U6895 (N_6895,N_5173,N_5188);
nand U6896 (N_6896,N_5060,N_5718);
and U6897 (N_6897,N_5212,N_5422);
nor U6898 (N_6898,N_5820,N_5695);
xnor U6899 (N_6899,N_5483,N_5617);
and U6900 (N_6900,N_5260,N_5890);
nor U6901 (N_6901,N_5638,N_5939);
nand U6902 (N_6902,N_5804,N_5391);
or U6903 (N_6903,N_5830,N_5169);
nand U6904 (N_6904,N_5174,N_5668);
or U6905 (N_6905,N_5317,N_5816);
nor U6906 (N_6906,N_5699,N_5260);
and U6907 (N_6907,N_5607,N_5030);
nand U6908 (N_6908,N_5627,N_5235);
nor U6909 (N_6909,N_5271,N_5803);
nand U6910 (N_6910,N_5519,N_5004);
and U6911 (N_6911,N_5514,N_5671);
xnor U6912 (N_6912,N_5028,N_5895);
or U6913 (N_6913,N_5420,N_5076);
nor U6914 (N_6914,N_5011,N_5255);
xor U6915 (N_6915,N_5088,N_5884);
nand U6916 (N_6916,N_5380,N_5841);
or U6917 (N_6917,N_5896,N_5407);
and U6918 (N_6918,N_5330,N_5743);
or U6919 (N_6919,N_5760,N_5020);
xnor U6920 (N_6920,N_5333,N_5719);
or U6921 (N_6921,N_5551,N_5807);
xor U6922 (N_6922,N_5927,N_5701);
nand U6923 (N_6923,N_5463,N_5583);
and U6924 (N_6924,N_5304,N_5022);
nor U6925 (N_6925,N_5671,N_5120);
nor U6926 (N_6926,N_5839,N_5134);
and U6927 (N_6927,N_5324,N_5978);
nor U6928 (N_6928,N_5453,N_5640);
nand U6929 (N_6929,N_5484,N_5297);
or U6930 (N_6930,N_5960,N_5566);
nor U6931 (N_6931,N_5573,N_5780);
nand U6932 (N_6932,N_5721,N_5208);
or U6933 (N_6933,N_5502,N_5227);
nor U6934 (N_6934,N_5314,N_5058);
or U6935 (N_6935,N_5054,N_5198);
or U6936 (N_6936,N_5701,N_5913);
or U6937 (N_6937,N_5769,N_5737);
or U6938 (N_6938,N_5170,N_5669);
xnor U6939 (N_6939,N_5197,N_5909);
and U6940 (N_6940,N_5580,N_5801);
nand U6941 (N_6941,N_5109,N_5203);
and U6942 (N_6942,N_5879,N_5407);
or U6943 (N_6943,N_5143,N_5422);
nand U6944 (N_6944,N_5180,N_5039);
nor U6945 (N_6945,N_5658,N_5697);
xnor U6946 (N_6946,N_5273,N_5061);
or U6947 (N_6947,N_5239,N_5407);
or U6948 (N_6948,N_5853,N_5818);
or U6949 (N_6949,N_5092,N_5961);
nor U6950 (N_6950,N_5144,N_5837);
and U6951 (N_6951,N_5041,N_5130);
xor U6952 (N_6952,N_5076,N_5331);
or U6953 (N_6953,N_5972,N_5794);
and U6954 (N_6954,N_5616,N_5790);
nand U6955 (N_6955,N_5548,N_5546);
nor U6956 (N_6956,N_5689,N_5800);
nand U6957 (N_6957,N_5733,N_5578);
nand U6958 (N_6958,N_5793,N_5614);
nor U6959 (N_6959,N_5969,N_5874);
and U6960 (N_6960,N_5097,N_5433);
nor U6961 (N_6961,N_5170,N_5612);
nor U6962 (N_6962,N_5821,N_5825);
nor U6963 (N_6963,N_5780,N_5962);
and U6964 (N_6964,N_5116,N_5411);
xor U6965 (N_6965,N_5650,N_5299);
and U6966 (N_6966,N_5747,N_5330);
xnor U6967 (N_6967,N_5046,N_5111);
or U6968 (N_6968,N_5950,N_5249);
nor U6969 (N_6969,N_5631,N_5258);
or U6970 (N_6970,N_5230,N_5915);
nand U6971 (N_6971,N_5659,N_5449);
and U6972 (N_6972,N_5308,N_5161);
or U6973 (N_6973,N_5556,N_5547);
and U6974 (N_6974,N_5848,N_5629);
nor U6975 (N_6975,N_5771,N_5943);
nand U6976 (N_6976,N_5717,N_5320);
and U6977 (N_6977,N_5645,N_5798);
nand U6978 (N_6978,N_5827,N_5969);
nor U6979 (N_6979,N_5907,N_5215);
xor U6980 (N_6980,N_5703,N_5441);
and U6981 (N_6981,N_5808,N_5977);
nor U6982 (N_6982,N_5318,N_5055);
xnor U6983 (N_6983,N_5029,N_5101);
and U6984 (N_6984,N_5998,N_5767);
or U6985 (N_6985,N_5171,N_5543);
nor U6986 (N_6986,N_5067,N_5600);
and U6987 (N_6987,N_5573,N_5049);
or U6988 (N_6988,N_5400,N_5069);
and U6989 (N_6989,N_5702,N_5023);
nor U6990 (N_6990,N_5723,N_5394);
nor U6991 (N_6991,N_5671,N_5854);
nor U6992 (N_6992,N_5914,N_5145);
and U6993 (N_6993,N_5884,N_5312);
or U6994 (N_6994,N_5695,N_5668);
and U6995 (N_6995,N_5442,N_5678);
nand U6996 (N_6996,N_5990,N_5562);
and U6997 (N_6997,N_5920,N_5042);
or U6998 (N_6998,N_5254,N_5811);
nor U6999 (N_6999,N_5983,N_5352);
nand U7000 (N_7000,N_6002,N_6986);
nand U7001 (N_7001,N_6227,N_6468);
nand U7002 (N_7002,N_6004,N_6566);
and U7003 (N_7003,N_6073,N_6912);
and U7004 (N_7004,N_6295,N_6683);
nand U7005 (N_7005,N_6250,N_6780);
nand U7006 (N_7006,N_6712,N_6045);
or U7007 (N_7007,N_6821,N_6260);
nand U7008 (N_7008,N_6306,N_6657);
and U7009 (N_7009,N_6554,N_6363);
nand U7010 (N_7010,N_6883,N_6461);
and U7011 (N_7011,N_6977,N_6587);
or U7012 (N_7012,N_6740,N_6823);
and U7013 (N_7013,N_6679,N_6943);
and U7014 (N_7014,N_6800,N_6789);
nand U7015 (N_7015,N_6117,N_6089);
and U7016 (N_7016,N_6463,N_6076);
or U7017 (N_7017,N_6484,N_6244);
and U7018 (N_7018,N_6005,N_6131);
nand U7019 (N_7019,N_6026,N_6187);
or U7020 (N_7020,N_6033,N_6339);
nand U7021 (N_7021,N_6776,N_6636);
nor U7022 (N_7022,N_6514,N_6826);
and U7023 (N_7023,N_6634,N_6469);
and U7024 (N_7024,N_6121,N_6689);
or U7025 (N_7025,N_6772,N_6997);
nor U7026 (N_7026,N_6752,N_6685);
nor U7027 (N_7027,N_6188,N_6980);
and U7028 (N_7028,N_6533,N_6923);
nor U7029 (N_7029,N_6944,N_6460);
nand U7030 (N_7030,N_6793,N_6629);
nor U7031 (N_7031,N_6788,N_6124);
xnor U7032 (N_7032,N_6704,N_6105);
xnor U7033 (N_7033,N_6720,N_6455);
xnor U7034 (N_7034,N_6050,N_6531);
and U7035 (N_7035,N_6995,N_6608);
nand U7036 (N_7036,N_6955,N_6583);
or U7037 (N_7037,N_6924,N_6770);
nand U7038 (N_7038,N_6413,N_6078);
or U7039 (N_7039,N_6388,N_6079);
and U7040 (N_7040,N_6946,N_6391);
and U7041 (N_7041,N_6537,N_6114);
or U7042 (N_7042,N_6046,N_6054);
nand U7043 (N_7043,N_6799,N_6062);
or U7044 (N_7044,N_6411,N_6327);
nor U7045 (N_7045,N_6971,N_6233);
nand U7046 (N_7046,N_6577,N_6156);
and U7047 (N_7047,N_6113,N_6624);
and U7048 (N_7048,N_6321,N_6653);
and U7049 (N_7049,N_6906,N_6612);
nor U7050 (N_7050,N_6769,N_6410);
nor U7051 (N_7051,N_6402,N_6508);
nand U7052 (N_7052,N_6319,N_6948);
or U7053 (N_7053,N_6690,N_6771);
xnor U7054 (N_7054,N_6070,N_6518);
nand U7055 (N_7055,N_6022,N_6103);
and U7056 (N_7056,N_6525,N_6497);
and U7057 (N_7057,N_6438,N_6506);
or U7058 (N_7058,N_6746,N_6169);
nand U7059 (N_7059,N_6096,N_6840);
or U7060 (N_7060,N_6648,N_6052);
and U7061 (N_7061,N_6546,N_6208);
and U7062 (N_7062,N_6697,N_6080);
and U7063 (N_7063,N_6847,N_6978);
or U7064 (N_7064,N_6757,N_6621);
and U7065 (N_7065,N_6386,N_6768);
nand U7066 (N_7066,N_6904,N_6729);
xor U7067 (N_7067,N_6684,N_6494);
or U7068 (N_7068,N_6705,N_6063);
and U7069 (N_7069,N_6818,N_6953);
xnor U7070 (N_7070,N_6365,N_6905);
or U7071 (N_7071,N_6110,N_6966);
and U7072 (N_7072,N_6011,N_6029);
or U7073 (N_7073,N_6722,N_6398);
xnor U7074 (N_7074,N_6500,N_6901);
or U7075 (N_7075,N_6220,N_6673);
xnor U7076 (N_7076,N_6628,N_6226);
xnor U7077 (N_7077,N_6568,N_6021);
nor U7078 (N_7078,N_6259,N_6238);
or U7079 (N_7079,N_6532,N_6559);
and U7080 (N_7080,N_6876,N_6359);
and U7081 (N_7081,N_6805,N_6444);
nor U7082 (N_7082,N_6256,N_6507);
nand U7083 (N_7083,N_6421,N_6197);
xor U7084 (N_7084,N_6926,N_6087);
nor U7085 (N_7085,N_6018,N_6782);
nor U7086 (N_7086,N_6938,N_6499);
nor U7087 (N_7087,N_6618,N_6833);
or U7088 (N_7088,N_6291,N_6877);
nor U7089 (N_7089,N_6606,N_6318);
nand U7090 (N_7090,N_6465,N_6387);
nand U7091 (N_7091,N_6517,N_6732);
nand U7092 (N_7092,N_6867,N_6257);
xor U7093 (N_7093,N_6146,N_6846);
nand U7094 (N_7094,N_6964,N_6343);
nand U7095 (N_7095,N_6707,N_6837);
xnor U7096 (N_7096,N_6708,N_6841);
and U7097 (N_7097,N_6936,N_6625);
nand U7098 (N_7098,N_6854,N_6686);
and U7099 (N_7099,N_6862,N_6892);
and U7100 (N_7100,N_6434,N_6389);
or U7101 (N_7101,N_6540,N_6158);
nand U7102 (N_7102,N_6842,N_6125);
and U7103 (N_7103,N_6392,N_6013);
xor U7104 (N_7104,N_6863,N_6151);
nand U7105 (N_7105,N_6878,N_6472);
xnor U7106 (N_7106,N_6298,N_6055);
and U7107 (N_7107,N_6613,N_6212);
nor U7108 (N_7108,N_6420,N_6916);
nor U7109 (N_7109,N_6322,N_6888);
or U7110 (N_7110,N_6326,N_6868);
nor U7111 (N_7111,N_6795,N_6317);
and U7112 (N_7112,N_6962,N_6639);
or U7113 (N_7113,N_6462,N_6817);
xnor U7114 (N_7114,N_6165,N_6860);
nand U7115 (N_7115,N_6541,N_6246);
and U7116 (N_7116,N_6214,N_6489);
and U7117 (N_7117,N_6490,N_6677);
nor U7118 (N_7118,N_6034,N_6399);
or U7119 (N_7119,N_6999,N_6443);
nor U7120 (N_7120,N_6237,N_6902);
or U7121 (N_7121,N_6945,N_6714);
or U7122 (N_7122,N_6739,N_6611);
nand U7123 (N_7123,N_6019,N_6652);
or U7124 (N_7124,N_6996,N_6148);
xnor U7125 (N_7125,N_6838,N_6601);
and U7126 (N_7126,N_6660,N_6929);
or U7127 (N_7127,N_6400,N_6377);
or U7128 (N_7128,N_6027,N_6135);
and U7129 (N_7129,N_6572,N_6798);
and U7130 (N_7130,N_6825,N_6213);
nor U7131 (N_7131,N_6643,N_6111);
nor U7132 (N_7132,N_6934,N_6965);
and U7133 (N_7133,N_6102,N_6483);
or U7134 (N_7134,N_6473,N_6510);
nor U7135 (N_7135,N_6272,N_6366);
and U7136 (N_7136,N_6567,N_6255);
and U7137 (N_7137,N_6098,N_6985);
nor U7138 (N_7138,N_6235,N_6196);
nor U7139 (N_7139,N_6157,N_6496);
nor U7140 (N_7140,N_6448,N_6030);
xor U7141 (N_7141,N_6819,N_6409);
nand U7142 (N_7142,N_6267,N_6287);
nand U7143 (N_7143,N_6703,N_6325);
and U7144 (N_7144,N_6289,N_6207);
nor U7145 (N_7145,N_6597,N_6861);
and U7146 (N_7146,N_6889,N_6312);
xnor U7147 (N_7147,N_6136,N_6718);
xor U7148 (N_7148,N_6812,N_6815);
nor U7149 (N_7149,N_6414,N_6006);
nor U7150 (N_7150,N_6616,N_6987);
or U7151 (N_7151,N_6794,N_6032);
nand U7152 (N_7152,N_6898,N_6632);
xnor U7153 (N_7153,N_6385,N_6894);
nand U7154 (N_7154,N_6334,N_6551);
and U7155 (N_7155,N_6759,N_6743);
nand U7156 (N_7156,N_6493,N_6236);
and U7157 (N_7157,N_6333,N_6038);
and U7158 (N_7158,N_6349,N_6442);
and U7159 (N_7159,N_6205,N_6337);
or U7160 (N_7160,N_6160,N_6266);
and U7161 (N_7161,N_6879,N_6139);
and U7162 (N_7162,N_6641,N_6808);
and U7163 (N_7163,N_6224,N_6573);
nand U7164 (N_7164,N_6311,N_6681);
and U7165 (N_7165,N_6661,N_6766);
nor U7166 (N_7166,N_6180,N_6633);
or U7167 (N_7167,N_6228,N_6249);
nor U7168 (N_7168,N_6345,N_6164);
or U7169 (N_7169,N_6492,N_6090);
or U7170 (N_7170,N_6579,N_6851);
or U7171 (N_7171,N_6774,N_6240);
and U7172 (N_7172,N_6723,N_6201);
nand U7173 (N_7173,N_6412,N_6893);
and U7174 (N_7174,N_6061,N_6353);
or U7175 (N_7175,N_6425,N_6453);
xor U7176 (N_7176,N_6756,N_6562);
nor U7177 (N_7177,N_6362,N_6575);
xnor U7178 (N_7178,N_6215,N_6764);
nand U7179 (N_7179,N_6149,N_6582);
nand U7180 (N_7180,N_6174,N_6171);
or U7181 (N_7181,N_6968,N_6041);
xnor U7182 (N_7182,N_6376,N_6503);
nor U7183 (N_7183,N_6431,N_6881);
or U7184 (N_7184,N_6430,N_6428);
and U7185 (N_7185,N_6302,N_6932);
or U7186 (N_7186,N_6976,N_6384);
nor U7187 (N_7187,N_6803,N_6390);
xnor U7188 (N_7188,N_6992,N_6544);
nand U7189 (N_7189,N_6591,N_6827);
and U7190 (N_7190,N_6107,N_6809);
nor U7191 (N_7191,N_6560,N_6719);
or U7192 (N_7192,N_6380,N_6667);
nand U7193 (N_7193,N_6942,N_6843);
nor U7194 (N_7194,N_6086,N_6513);
and U7195 (N_7195,N_6476,N_6580);
nor U7196 (N_7196,N_6713,N_6885);
and U7197 (N_7197,N_6527,N_6264);
xor U7198 (N_7198,N_6536,N_6432);
or U7199 (N_7199,N_6839,N_6535);
nor U7200 (N_7200,N_6137,N_6159);
or U7201 (N_7201,N_6736,N_6828);
nor U7202 (N_7202,N_6734,N_6277);
and U7203 (N_7203,N_6604,N_6074);
nand U7204 (N_7204,N_6176,N_6346);
and U7205 (N_7205,N_6694,N_6020);
nand U7206 (N_7206,N_6101,N_6261);
or U7207 (N_7207,N_6880,N_6669);
nand U7208 (N_7208,N_6891,N_6687);
and U7209 (N_7209,N_6057,N_6557);
nand U7210 (N_7210,N_6071,N_6920);
nor U7211 (N_7211,N_6143,N_6501);
and U7212 (N_7212,N_6569,N_6477);
xnor U7213 (N_7213,N_6806,N_6297);
and U7214 (N_7214,N_6441,N_6724);
nand U7215 (N_7215,N_6108,N_6913);
or U7216 (N_7216,N_6692,N_6265);
nand U7217 (N_7217,N_6014,N_6069);
nand U7218 (N_7218,N_6754,N_6104);
or U7219 (N_7219,N_6984,N_6012);
and U7220 (N_7220,N_6239,N_6225);
nor U7221 (N_7221,N_6585,N_6547);
nand U7222 (N_7222,N_6459,N_6662);
xor U7223 (N_7223,N_6664,N_6951);
nor U7224 (N_7224,N_6748,N_6128);
or U7225 (N_7225,N_6179,N_6900);
and U7226 (N_7226,N_6315,N_6347);
nand U7227 (N_7227,N_6275,N_6609);
or U7228 (N_7228,N_6897,N_6751);
nor U7229 (N_7229,N_6451,N_6232);
nand U7230 (N_7230,N_6674,N_6276);
and U7231 (N_7231,N_6593,N_6701);
nor U7232 (N_7232,N_6456,N_6822);
nand U7233 (N_7233,N_6738,N_6796);
or U7234 (N_7234,N_6859,N_6085);
nand U7235 (N_7235,N_6134,N_6711);
nand U7236 (N_7236,N_6749,N_6811);
nand U7237 (N_7237,N_6543,N_6163);
nor U7238 (N_7238,N_6274,N_6873);
nor U7239 (N_7239,N_6850,N_6969);
nor U7240 (N_7240,N_6449,N_6142);
and U7241 (N_7241,N_6024,N_6072);
nor U7242 (N_7242,N_6991,N_6007);
nand U7243 (N_7243,N_6241,N_6330);
nand U7244 (N_7244,N_6270,N_6427);
and U7245 (N_7245,N_6369,N_6963);
and U7246 (N_7246,N_6979,N_6150);
or U7247 (N_7247,N_6068,N_6252);
or U7248 (N_7248,N_6067,N_6300);
or U7249 (N_7249,N_6899,N_6132);
and U7250 (N_7250,N_6292,N_6283);
or U7251 (N_7251,N_6765,N_6166);
nand U7252 (N_7252,N_6930,N_6426);
or U7253 (N_7253,N_6871,N_6209);
and U7254 (N_7254,N_6548,N_6742);
nor U7255 (N_7255,N_6301,N_6576);
nand U7256 (N_7256,N_6478,N_6271);
nor U7257 (N_7257,N_6109,N_6790);
nand U7258 (N_7258,N_6269,N_6578);
or U7259 (N_7259,N_6288,N_6229);
nor U7260 (N_7260,N_6230,N_6895);
or U7261 (N_7261,N_6185,N_6282);
and U7262 (N_7262,N_6154,N_6316);
nand U7263 (N_7263,N_6623,N_6273);
nand U7264 (N_7264,N_6675,N_6730);
nand U7265 (N_7265,N_6872,N_6829);
xnor U7266 (N_7266,N_6475,N_6059);
nand U7267 (N_7267,N_6589,N_6360);
or U7268 (N_7268,N_6130,N_6933);
or U7269 (N_7269,N_6355,N_6263);
nor U7270 (N_7270,N_6524,N_6037);
and U7271 (N_7271,N_6908,N_6485);
nand U7272 (N_7272,N_6716,N_6922);
or U7273 (N_7273,N_6975,N_6915);
or U7274 (N_7274,N_6981,N_6401);
or U7275 (N_7275,N_6561,N_6191);
or U7276 (N_7276,N_6314,N_6910);
nor U7277 (N_7277,N_6053,N_6175);
or U7278 (N_7278,N_6064,N_6440);
and U7279 (N_7279,N_6830,N_6670);
and U7280 (N_7280,N_6354,N_6305);
nand U7281 (N_7281,N_6120,N_6042);
and U7282 (N_7282,N_6153,N_6170);
nor U7283 (N_7283,N_6422,N_6009);
and U7284 (N_7284,N_6727,N_6381);
or U7285 (N_7285,N_6173,N_6044);
and U7286 (N_7286,N_6656,N_6279);
nand U7287 (N_7287,N_6558,N_6530);
nor U7288 (N_7288,N_6351,N_6066);
nor U7289 (N_7289,N_6281,N_6186);
nor U7290 (N_7290,N_6299,N_6970);
or U7291 (N_7291,N_6504,N_6509);
xnor U7292 (N_7292,N_6393,N_6332);
xnor U7293 (N_7293,N_6590,N_6058);
or U7294 (N_7294,N_6309,N_6065);
nand U7295 (N_7295,N_6133,N_6855);
or U7296 (N_7296,N_6184,N_6082);
nor U7297 (N_7297,N_6408,N_6331);
nor U7298 (N_7298,N_6947,N_6152);
or U7299 (N_7299,N_6048,N_6199);
or U7300 (N_7300,N_6814,N_6047);
and U7301 (N_7301,N_6668,N_6595);
xor U7302 (N_7302,N_6731,N_6429);
or U7303 (N_7303,N_6710,N_6310);
nor U7304 (N_7304,N_6845,N_6520);
or U7305 (N_7305,N_6552,N_6417);
nor U7306 (N_7306,N_6647,N_6638);
and U7307 (N_7307,N_6890,N_6630);
and U7308 (N_7308,N_6418,N_6918);
nand U7309 (N_7309,N_6592,N_6745);
nor U7310 (N_7310,N_6141,N_6869);
or U7311 (N_7311,N_6198,N_6631);
or U7312 (N_7312,N_6907,N_6804);
nor U7313 (N_7313,N_6744,N_6379);
nand U7314 (N_7314,N_6234,N_6696);
nand U7315 (N_7315,N_6051,N_6294);
or U7316 (N_7316,N_6994,N_6698);
or U7317 (N_7317,N_6571,N_6396);
or U7318 (N_7318,N_6471,N_6663);
and U7319 (N_7319,N_6760,N_6581);
or U7320 (N_7320,N_6340,N_6017);
or U7321 (N_7321,N_6452,N_6556);
nor U7322 (N_7322,N_6161,N_6937);
nor U7323 (N_7323,N_6659,N_6177);
and U7324 (N_7324,N_6989,N_6832);
and U7325 (N_7325,N_6974,N_6761);
nor U7326 (N_7326,N_6563,N_6382);
nor U7327 (N_7327,N_6285,N_6848);
nand U7328 (N_7328,N_6786,N_6491);
nor U7329 (N_7329,N_6404,N_6534);
nor U7330 (N_7330,N_6627,N_6614);
and U7331 (N_7331,N_6555,N_6375);
or U7332 (N_7332,N_6338,N_6982);
nor U7333 (N_7333,N_6168,N_6522);
and U7334 (N_7334,N_6728,N_6983);
nand U7335 (N_7335,N_6099,N_6549);
nand U7336 (N_7336,N_6655,N_6364);
nand U7337 (N_7337,N_6824,N_6084);
or U7338 (N_7338,N_6092,N_6802);
nor U7339 (N_7339,N_6081,N_6747);
nor U7340 (N_7340,N_6335,N_6395);
xnor U7341 (N_7341,N_6293,N_6341);
nor U7342 (N_7342,N_6635,N_6792);
nand U7343 (N_7343,N_6043,N_6268);
nor U7344 (N_7344,N_6665,N_6466);
xor U7345 (N_7345,N_6129,N_6258);
and U7346 (N_7346,N_6884,N_6834);
nor U7347 (N_7347,N_6858,N_6077);
nand U7348 (N_7348,N_6486,N_6959);
nand U7349 (N_7349,N_6735,N_6758);
or U7350 (N_7350,N_6028,N_6370);
nor U7351 (N_7351,N_6015,N_6584);
nor U7352 (N_7352,N_6040,N_6374);
nand U7353 (N_7353,N_6642,N_6116);
nor U7354 (N_7354,N_6495,N_6775);
xor U7355 (N_7355,N_6419,N_6973);
or U7356 (N_7356,N_6357,N_6035);
xor U7357 (N_7357,N_6095,N_6622);
or U7358 (N_7358,N_6511,N_6539);
and U7359 (N_7359,N_6195,N_6680);
nor U7360 (N_7360,N_6248,N_6403);
nor U7361 (N_7361,N_6397,N_6515);
xor U7362 (N_7362,N_6935,N_6231);
or U7363 (N_7363,N_6816,N_6242);
or U7364 (N_7364,N_6882,N_6307);
and U7365 (N_7365,N_6886,N_6596);
nor U7366 (N_7366,N_6831,N_6836);
or U7367 (N_7367,N_6481,N_6529);
and U7368 (N_7368,N_6695,N_6324);
xnor U7369 (N_7369,N_6445,N_6849);
nand U7370 (N_7370,N_6039,N_6056);
nand U7371 (N_7371,N_6436,N_6182);
xnor U7372 (N_7372,N_6512,N_6783);
nor U7373 (N_7373,N_6243,N_6820);
and U7374 (N_7374,N_6619,N_6925);
xnor U7375 (N_7375,N_6693,N_6521);
nand U7376 (N_7376,N_6487,N_6866);
and U7377 (N_7377,N_6725,N_6280);
xnor U7378 (N_7378,N_6464,N_6870);
xnor U7379 (N_7379,N_6553,N_6542);
or U7380 (N_7380,N_6378,N_6864);
or U7381 (N_7381,N_6650,N_6123);
nor U7382 (N_7382,N_6147,N_6167);
nand U7383 (N_7383,N_6717,N_6447);
and U7384 (N_7384,N_6406,N_6100);
and U7385 (N_7385,N_6450,N_6474);
nand U7386 (N_7386,N_6348,N_6637);
nand U7387 (N_7387,N_6733,N_6344);
xnor U7388 (N_7388,N_6140,N_6887);
or U7389 (N_7389,N_6003,N_6190);
and U7390 (N_7390,N_6211,N_6875);
nand U7391 (N_7391,N_6144,N_6988);
xnor U7392 (N_7392,N_6939,N_6526);
or U7393 (N_7393,N_6763,N_6219);
and U7394 (N_7394,N_6896,N_6458);
nor U7395 (N_7395,N_6779,N_6954);
or U7396 (N_7396,N_6480,N_6336);
or U7397 (N_7397,N_6204,N_6919);
and U7398 (N_7398,N_6023,N_6538);
and U7399 (N_7399,N_6588,N_6262);
nor U7400 (N_7400,N_6853,N_6284);
or U7401 (N_7401,N_6488,N_6741);
xor U7402 (N_7402,N_6290,N_6328);
or U7403 (N_7403,N_6658,N_6036);
and U7404 (N_7404,N_6119,N_6367);
nor U7405 (N_7405,N_6115,N_6203);
nand U7406 (N_7406,N_6106,N_6405);
nor U7407 (N_7407,N_6183,N_6691);
nand U7408 (N_7408,N_6620,N_6990);
and U7409 (N_7409,N_6941,N_6903);
or U7410 (N_7410,N_6813,N_6138);
and U7411 (N_7411,N_6200,N_6254);
and U7412 (N_7412,N_6784,N_6193);
nor U7413 (N_7413,N_6646,N_6672);
nand U7414 (N_7414,N_6251,N_6599);
and U7415 (N_7415,N_6528,N_6961);
nor U7416 (N_7416,N_6126,N_6470);
xor U7417 (N_7417,N_6865,N_6371);
xor U7418 (N_7418,N_6956,N_6940);
and U7419 (N_7419,N_6570,N_6709);
or U7420 (N_7420,N_6702,N_6304);
or U7421 (N_7421,N_6433,N_6008);
nand U7422 (N_7422,N_6781,N_6206);
nor U7423 (N_7423,N_6181,N_6091);
nor U7424 (N_7424,N_6286,N_6454);
nor U7425 (N_7425,N_6617,N_6957);
nor U7426 (N_7426,N_6753,N_6810);
nor U7427 (N_7427,N_6112,N_6640);
and U7428 (N_7428,N_6651,N_6372);
nand U7429 (N_7429,N_6564,N_6688);
or U7430 (N_7430,N_6807,N_6031);
nor U7431 (N_7431,N_6607,N_6202);
nand U7432 (N_7432,N_6223,N_6253);
nand U7433 (N_7433,N_6615,N_6931);
or U7434 (N_7434,N_6407,N_6917);
and U7435 (N_7435,N_6600,N_6162);
and U7436 (N_7436,N_6358,N_6247);
and U7437 (N_7437,N_6516,N_6602);
xor U7438 (N_7438,N_6928,N_6210);
xor U7439 (N_7439,N_6671,N_6001);
or U7440 (N_7440,N_6178,N_6498);
and U7441 (N_7441,N_6356,N_6610);
nor U7442 (N_7442,N_6218,N_6172);
or U7443 (N_7443,N_6644,N_6323);
nor U7444 (N_7444,N_6145,N_6649);
nor U7445 (N_7445,N_6715,N_6565);
or U7446 (N_7446,N_6993,N_6394);
nor U7447 (N_7447,N_6801,N_6949);
xor U7448 (N_7448,N_6368,N_6967);
xor U7449 (N_7449,N_6313,N_6424);
and U7450 (N_7450,N_6479,N_6952);
nor U7451 (N_7451,N_6678,N_6329);
nor U7452 (N_7452,N_6155,N_6654);
xor U7453 (N_7453,N_6773,N_6245);
nor U7454 (N_7454,N_6519,N_6605);
or U7455 (N_7455,N_6852,N_6467);
or U7456 (N_7456,N_6350,N_6457);
or U7457 (N_7457,N_6755,N_6972);
or U7458 (N_7458,N_6192,N_6598);
nor U7459 (N_7459,N_6217,N_6097);
and U7460 (N_7460,N_6010,N_6909);
nand U7461 (N_7461,N_6093,N_6950);
nor U7462 (N_7462,N_6221,N_6000);
and U7463 (N_7463,N_6423,N_6296);
nand U7464 (N_7464,N_6088,N_6750);
and U7465 (N_7465,N_6446,N_6415);
or U7466 (N_7466,N_6785,N_6914);
and U7467 (N_7467,N_6856,N_6706);
nand U7468 (N_7468,N_6676,N_6721);
nand U7469 (N_7469,N_6958,N_6921);
or U7470 (N_7470,N_6194,N_6016);
or U7471 (N_7471,N_6586,N_6911);
nor U7472 (N_7472,N_6700,N_6797);
or U7473 (N_7473,N_6320,N_6626);
or U7474 (N_7474,N_6352,N_6222);
and U7475 (N_7475,N_6726,N_6189);
or U7476 (N_7476,N_6844,N_6603);
nor U7477 (N_7477,N_6278,N_6523);
xor U7478 (N_7478,N_6594,N_6127);
nor U7479 (N_7479,N_6857,N_6998);
nand U7480 (N_7480,N_6791,N_6482);
xnor U7481 (N_7481,N_6666,N_6361);
and U7482 (N_7482,N_6787,N_6435);
and U7483 (N_7483,N_6416,N_6383);
nor U7484 (N_7484,N_6960,N_6049);
nor U7485 (N_7485,N_6122,N_6762);
nand U7486 (N_7486,N_6342,N_6737);
nand U7487 (N_7487,N_6060,N_6094);
and U7488 (N_7488,N_6373,N_6682);
and U7489 (N_7489,N_6303,N_6545);
or U7490 (N_7490,N_6118,N_6927);
or U7491 (N_7491,N_6075,N_6778);
and U7492 (N_7492,N_6874,N_6645);
and U7493 (N_7493,N_6550,N_6574);
or U7494 (N_7494,N_6835,N_6437);
or U7495 (N_7495,N_6083,N_6767);
nor U7496 (N_7496,N_6216,N_6025);
or U7497 (N_7497,N_6699,N_6439);
xor U7498 (N_7498,N_6308,N_6777);
nand U7499 (N_7499,N_6502,N_6505);
nor U7500 (N_7500,N_6162,N_6479);
nor U7501 (N_7501,N_6535,N_6217);
or U7502 (N_7502,N_6600,N_6443);
or U7503 (N_7503,N_6087,N_6800);
xor U7504 (N_7504,N_6253,N_6042);
or U7505 (N_7505,N_6316,N_6451);
xnor U7506 (N_7506,N_6586,N_6081);
nand U7507 (N_7507,N_6164,N_6707);
nor U7508 (N_7508,N_6659,N_6085);
and U7509 (N_7509,N_6469,N_6053);
xnor U7510 (N_7510,N_6784,N_6445);
xnor U7511 (N_7511,N_6213,N_6883);
nor U7512 (N_7512,N_6900,N_6473);
or U7513 (N_7513,N_6488,N_6378);
and U7514 (N_7514,N_6193,N_6840);
nor U7515 (N_7515,N_6915,N_6683);
nor U7516 (N_7516,N_6595,N_6601);
nand U7517 (N_7517,N_6627,N_6554);
or U7518 (N_7518,N_6818,N_6426);
nand U7519 (N_7519,N_6497,N_6446);
xor U7520 (N_7520,N_6820,N_6135);
nor U7521 (N_7521,N_6345,N_6095);
or U7522 (N_7522,N_6727,N_6710);
or U7523 (N_7523,N_6686,N_6788);
nor U7524 (N_7524,N_6491,N_6650);
and U7525 (N_7525,N_6706,N_6419);
nor U7526 (N_7526,N_6841,N_6095);
nor U7527 (N_7527,N_6293,N_6842);
nor U7528 (N_7528,N_6219,N_6985);
nand U7529 (N_7529,N_6625,N_6335);
xnor U7530 (N_7530,N_6908,N_6785);
xor U7531 (N_7531,N_6714,N_6955);
nand U7532 (N_7532,N_6616,N_6771);
xor U7533 (N_7533,N_6651,N_6772);
xor U7534 (N_7534,N_6325,N_6066);
nand U7535 (N_7535,N_6774,N_6087);
xnor U7536 (N_7536,N_6175,N_6925);
and U7537 (N_7537,N_6663,N_6776);
nor U7538 (N_7538,N_6412,N_6560);
xor U7539 (N_7539,N_6173,N_6842);
nor U7540 (N_7540,N_6952,N_6789);
nor U7541 (N_7541,N_6104,N_6303);
nand U7542 (N_7542,N_6890,N_6909);
nor U7543 (N_7543,N_6413,N_6841);
nor U7544 (N_7544,N_6250,N_6790);
nor U7545 (N_7545,N_6650,N_6224);
nand U7546 (N_7546,N_6047,N_6599);
or U7547 (N_7547,N_6140,N_6191);
xnor U7548 (N_7548,N_6571,N_6642);
or U7549 (N_7549,N_6795,N_6617);
nor U7550 (N_7550,N_6546,N_6757);
xor U7551 (N_7551,N_6627,N_6171);
nor U7552 (N_7552,N_6011,N_6129);
nor U7553 (N_7553,N_6572,N_6067);
nor U7554 (N_7554,N_6877,N_6968);
and U7555 (N_7555,N_6250,N_6861);
nand U7556 (N_7556,N_6519,N_6357);
nor U7557 (N_7557,N_6268,N_6070);
or U7558 (N_7558,N_6365,N_6200);
or U7559 (N_7559,N_6150,N_6482);
and U7560 (N_7560,N_6832,N_6649);
and U7561 (N_7561,N_6489,N_6968);
or U7562 (N_7562,N_6043,N_6641);
or U7563 (N_7563,N_6443,N_6662);
nand U7564 (N_7564,N_6599,N_6831);
nand U7565 (N_7565,N_6565,N_6429);
and U7566 (N_7566,N_6655,N_6765);
xor U7567 (N_7567,N_6488,N_6450);
and U7568 (N_7568,N_6744,N_6098);
and U7569 (N_7569,N_6648,N_6081);
nand U7570 (N_7570,N_6166,N_6036);
nor U7571 (N_7571,N_6087,N_6756);
nand U7572 (N_7572,N_6151,N_6762);
or U7573 (N_7573,N_6066,N_6782);
nand U7574 (N_7574,N_6219,N_6651);
or U7575 (N_7575,N_6473,N_6782);
nand U7576 (N_7576,N_6417,N_6080);
nor U7577 (N_7577,N_6711,N_6066);
and U7578 (N_7578,N_6907,N_6833);
and U7579 (N_7579,N_6822,N_6967);
xnor U7580 (N_7580,N_6420,N_6557);
or U7581 (N_7581,N_6115,N_6237);
nor U7582 (N_7582,N_6925,N_6759);
and U7583 (N_7583,N_6486,N_6690);
nand U7584 (N_7584,N_6616,N_6776);
nand U7585 (N_7585,N_6503,N_6318);
nor U7586 (N_7586,N_6015,N_6257);
nand U7587 (N_7587,N_6612,N_6883);
nor U7588 (N_7588,N_6472,N_6368);
nor U7589 (N_7589,N_6280,N_6634);
and U7590 (N_7590,N_6048,N_6569);
or U7591 (N_7591,N_6037,N_6302);
nand U7592 (N_7592,N_6943,N_6710);
nor U7593 (N_7593,N_6546,N_6281);
nor U7594 (N_7594,N_6094,N_6724);
or U7595 (N_7595,N_6020,N_6463);
xor U7596 (N_7596,N_6467,N_6323);
nor U7597 (N_7597,N_6618,N_6604);
or U7598 (N_7598,N_6053,N_6246);
nand U7599 (N_7599,N_6032,N_6306);
nand U7600 (N_7600,N_6281,N_6992);
or U7601 (N_7601,N_6860,N_6932);
nor U7602 (N_7602,N_6434,N_6347);
nand U7603 (N_7603,N_6822,N_6267);
nor U7604 (N_7604,N_6703,N_6719);
or U7605 (N_7605,N_6167,N_6470);
and U7606 (N_7606,N_6419,N_6365);
nor U7607 (N_7607,N_6891,N_6079);
and U7608 (N_7608,N_6430,N_6719);
xor U7609 (N_7609,N_6064,N_6103);
and U7610 (N_7610,N_6455,N_6705);
and U7611 (N_7611,N_6702,N_6779);
or U7612 (N_7612,N_6256,N_6458);
nor U7613 (N_7613,N_6366,N_6821);
nand U7614 (N_7614,N_6896,N_6779);
nor U7615 (N_7615,N_6918,N_6712);
xnor U7616 (N_7616,N_6238,N_6798);
xor U7617 (N_7617,N_6253,N_6476);
nand U7618 (N_7618,N_6514,N_6534);
nor U7619 (N_7619,N_6616,N_6633);
or U7620 (N_7620,N_6549,N_6393);
nand U7621 (N_7621,N_6550,N_6001);
nor U7622 (N_7622,N_6433,N_6237);
or U7623 (N_7623,N_6448,N_6110);
or U7624 (N_7624,N_6392,N_6237);
and U7625 (N_7625,N_6688,N_6286);
or U7626 (N_7626,N_6319,N_6028);
nor U7627 (N_7627,N_6102,N_6266);
xnor U7628 (N_7628,N_6315,N_6927);
nor U7629 (N_7629,N_6773,N_6718);
nor U7630 (N_7630,N_6988,N_6567);
nand U7631 (N_7631,N_6712,N_6990);
or U7632 (N_7632,N_6920,N_6367);
and U7633 (N_7633,N_6945,N_6066);
and U7634 (N_7634,N_6821,N_6920);
and U7635 (N_7635,N_6276,N_6426);
or U7636 (N_7636,N_6035,N_6723);
or U7637 (N_7637,N_6428,N_6622);
or U7638 (N_7638,N_6696,N_6263);
nand U7639 (N_7639,N_6271,N_6252);
nor U7640 (N_7640,N_6906,N_6519);
xor U7641 (N_7641,N_6394,N_6501);
and U7642 (N_7642,N_6461,N_6388);
or U7643 (N_7643,N_6652,N_6262);
nand U7644 (N_7644,N_6202,N_6731);
nor U7645 (N_7645,N_6763,N_6996);
and U7646 (N_7646,N_6767,N_6930);
or U7647 (N_7647,N_6707,N_6674);
nand U7648 (N_7648,N_6545,N_6846);
nand U7649 (N_7649,N_6219,N_6589);
and U7650 (N_7650,N_6393,N_6898);
and U7651 (N_7651,N_6391,N_6491);
or U7652 (N_7652,N_6447,N_6786);
nand U7653 (N_7653,N_6795,N_6345);
and U7654 (N_7654,N_6889,N_6350);
or U7655 (N_7655,N_6773,N_6206);
or U7656 (N_7656,N_6517,N_6238);
and U7657 (N_7657,N_6304,N_6834);
and U7658 (N_7658,N_6356,N_6935);
and U7659 (N_7659,N_6382,N_6624);
xnor U7660 (N_7660,N_6698,N_6846);
nor U7661 (N_7661,N_6529,N_6894);
and U7662 (N_7662,N_6990,N_6013);
nand U7663 (N_7663,N_6272,N_6917);
and U7664 (N_7664,N_6115,N_6210);
nor U7665 (N_7665,N_6798,N_6532);
nor U7666 (N_7666,N_6010,N_6597);
and U7667 (N_7667,N_6359,N_6602);
xnor U7668 (N_7668,N_6269,N_6751);
nor U7669 (N_7669,N_6620,N_6227);
or U7670 (N_7670,N_6966,N_6438);
and U7671 (N_7671,N_6986,N_6884);
and U7672 (N_7672,N_6777,N_6247);
and U7673 (N_7673,N_6283,N_6611);
or U7674 (N_7674,N_6140,N_6675);
or U7675 (N_7675,N_6437,N_6865);
and U7676 (N_7676,N_6845,N_6779);
nor U7677 (N_7677,N_6615,N_6282);
nand U7678 (N_7678,N_6775,N_6646);
or U7679 (N_7679,N_6669,N_6247);
and U7680 (N_7680,N_6532,N_6245);
xor U7681 (N_7681,N_6795,N_6440);
or U7682 (N_7682,N_6771,N_6284);
xnor U7683 (N_7683,N_6242,N_6267);
and U7684 (N_7684,N_6319,N_6015);
nand U7685 (N_7685,N_6814,N_6952);
xnor U7686 (N_7686,N_6856,N_6388);
nand U7687 (N_7687,N_6736,N_6792);
and U7688 (N_7688,N_6029,N_6916);
nor U7689 (N_7689,N_6814,N_6760);
and U7690 (N_7690,N_6095,N_6793);
or U7691 (N_7691,N_6485,N_6061);
and U7692 (N_7692,N_6070,N_6869);
and U7693 (N_7693,N_6937,N_6093);
nand U7694 (N_7694,N_6799,N_6157);
or U7695 (N_7695,N_6882,N_6759);
or U7696 (N_7696,N_6727,N_6654);
nor U7697 (N_7697,N_6886,N_6628);
and U7698 (N_7698,N_6721,N_6548);
or U7699 (N_7699,N_6695,N_6245);
and U7700 (N_7700,N_6217,N_6211);
nand U7701 (N_7701,N_6579,N_6901);
or U7702 (N_7702,N_6203,N_6745);
nor U7703 (N_7703,N_6952,N_6659);
nand U7704 (N_7704,N_6212,N_6854);
or U7705 (N_7705,N_6733,N_6167);
or U7706 (N_7706,N_6329,N_6288);
nand U7707 (N_7707,N_6554,N_6364);
and U7708 (N_7708,N_6035,N_6530);
and U7709 (N_7709,N_6490,N_6137);
and U7710 (N_7710,N_6689,N_6832);
or U7711 (N_7711,N_6756,N_6344);
nand U7712 (N_7712,N_6452,N_6936);
xnor U7713 (N_7713,N_6772,N_6163);
and U7714 (N_7714,N_6375,N_6753);
nand U7715 (N_7715,N_6083,N_6616);
nor U7716 (N_7716,N_6604,N_6899);
nor U7717 (N_7717,N_6785,N_6031);
nand U7718 (N_7718,N_6109,N_6325);
nand U7719 (N_7719,N_6193,N_6343);
and U7720 (N_7720,N_6877,N_6774);
nor U7721 (N_7721,N_6431,N_6008);
nor U7722 (N_7722,N_6432,N_6242);
nand U7723 (N_7723,N_6107,N_6659);
nand U7724 (N_7724,N_6612,N_6674);
and U7725 (N_7725,N_6942,N_6431);
nor U7726 (N_7726,N_6114,N_6784);
or U7727 (N_7727,N_6636,N_6145);
and U7728 (N_7728,N_6385,N_6845);
and U7729 (N_7729,N_6966,N_6004);
nor U7730 (N_7730,N_6499,N_6253);
or U7731 (N_7731,N_6922,N_6525);
nor U7732 (N_7732,N_6721,N_6501);
nand U7733 (N_7733,N_6862,N_6006);
and U7734 (N_7734,N_6972,N_6297);
and U7735 (N_7735,N_6712,N_6742);
nor U7736 (N_7736,N_6755,N_6447);
nor U7737 (N_7737,N_6828,N_6387);
and U7738 (N_7738,N_6094,N_6896);
nand U7739 (N_7739,N_6168,N_6775);
and U7740 (N_7740,N_6865,N_6231);
nand U7741 (N_7741,N_6398,N_6303);
nand U7742 (N_7742,N_6499,N_6665);
nor U7743 (N_7743,N_6251,N_6762);
and U7744 (N_7744,N_6939,N_6625);
nor U7745 (N_7745,N_6746,N_6259);
and U7746 (N_7746,N_6104,N_6649);
and U7747 (N_7747,N_6044,N_6670);
nand U7748 (N_7748,N_6283,N_6549);
and U7749 (N_7749,N_6826,N_6759);
nor U7750 (N_7750,N_6706,N_6365);
xnor U7751 (N_7751,N_6085,N_6701);
and U7752 (N_7752,N_6812,N_6559);
nand U7753 (N_7753,N_6406,N_6662);
and U7754 (N_7754,N_6850,N_6359);
and U7755 (N_7755,N_6536,N_6902);
nor U7756 (N_7756,N_6957,N_6401);
nor U7757 (N_7757,N_6861,N_6091);
xor U7758 (N_7758,N_6166,N_6567);
and U7759 (N_7759,N_6221,N_6370);
nand U7760 (N_7760,N_6671,N_6875);
nor U7761 (N_7761,N_6443,N_6842);
and U7762 (N_7762,N_6930,N_6677);
or U7763 (N_7763,N_6461,N_6746);
xnor U7764 (N_7764,N_6325,N_6940);
or U7765 (N_7765,N_6947,N_6630);
nand U7766 (N_7766,N_6104,N_6765);
nor U7767 (N_7767,N_6079,N_6872);
and U7768 (N_7768,N_6873,N_6503);
nor U7769 (N_7769,N_6560,N_6400);
and U7770 (N_7770,N_6569,N_6391);
nand U7771 (N_7771,N_6529,N_6203);
and U7772 (N_7772,N_6792,N_6722);
and U7773 (N_7773,N_6790,N_6814);
or U7774 (N_7774,N_6146,N_6781);
xor U7775 (N_7775,N_6263,N_6768);
and U7776 (N_7776,N_6983,N_6677);
nand U7777 (N_7777,N_6617,N_6231);
nand U7778 (N_7778,N_6429,N_6102);
and U7779 (N_7779,N_6515,N_6070);
nand U7780 (N_7780,N_6001,N_6534);
nand U7781 (N_7781,N_6112,N_6284);
nand U7782 (N_7782,N_6333,N_6300);
nand U7783 (N_7783,N_6040,N_6632);
nand U7784 (N_7784,N_6026,N_6295);
xor U7785 (N_7785,N_6768,N_6255);
nand U7786 (N_7786,N_6613,N_6122);
or U7787 (N_7787,N_6607,N_6229);
nand U7788 (N_7788,N_6393,N_6743);
and U7789 (N_7789,N_6227,N_6014);
or U7790 (N_7790,N_6207,N_6913);
nor U7791 (N_7791,N_6170,N_6767);
and U7792 (N_7792,N_6317,N_6936);
nand U7793 (N_7793,N_6933,N_6677);
or U7794 (N_7794,N_6517,N_6229);
nor U7795 (N_7795,N_6995,N_6454);
nand U7796 (N_7796,N_6590,N_6869);
nand U7797 (N_7797,N_6315,N_6306);
and U7798 (N_7798,N_6797,N_6285);
nor U7799 (N_7799,N_6645,N_6513);
nor U7800 (N_7800,N_6528,N_6550);
nand U7801 (N_7801,N_6692,N_6819);
and U7802 (N_7802,N_6742,N_6656);
nand U7803 (N_7803,N_6075,N_6604);
nand U7804 (N_7804,N_6107,N_6417);
nor U7805 (N_7805,N_6442,N_6380);
or U7806 (N_7806,N_6442,N_6302);
nor U7807 (N_7807,N_6983,N_6117);
and U7808 (N_7808,N_6650,N_6455);
nand U7809 (N_7809,N_6649,N_6274);
xnor U7810 (N_7810,N_6746,N_6798);
nor U7811 (N_7811,N_6561,N_6984);
nand U7812 (N_7812,N_6523,N_6802);
xnor U7813 (N_7813,N_6111,N_6688);
and U7814 (N_7814,N_6073,N_6193);
xnor U7815 (N_7815,N_6137,N_6578);
and U7816 (N_7816,N_6901,N_6072);
or U7817 (N_7817,N_6855,N_6900);
nor U7818 (N_7818,N_6502,N_6345);
xnor U7819 (N_7819,N_6447,N_6802);
or U7820 (N_7820,N_6401,N_6496);
nor U7821 (N_7821,N_6807,N_6939);
or U7822 (N_7822,N_6260,N_6244);
or U7823 (N_7823,N_6477,N_6147);
or U7824 (N_7824,N_6524,N_6802);
xor U7825 (N_7825,N_6241,N_6747);
or U7826 (N_7826,N_6889,N_6875);
nor U7827 (N_7827,N_6210,N_6124);
and U7828 (N_7828,N_6182,N_6372);
nor U7829 (N_7829,N_6827,N_6416);
nand U7830 (N_7830,N_6288,N_6274);
and U7831 (N_7831,N_6244,N_6409);
nand U7832 (N_7832,N_6155,N_6061);
nand U7833 (N_7833,N_6974,N_6433);
nand U7834 (N_7834,N_6189,N_6019);
nor U7835 (N_7835,N_6683,N_6853);
nand U7836 (N_7836,N_6305,N_6382);
or U7837 (N_7837,N_6870,N_6088);
nor U7838 (N_7838,N_6387,N_6644);
or U7839 (N_7839,N_6791,N_6511);
nand U7840 (N_7840,N_6306,N_6365);
nor U7841 (N_7841,N_6741,N_6760);
and U7842 (N_7842,N_6220,N_6955);
nand U7843 (N_7843,N_6678,N_6003);
nand U7844 (N_7844,N_6232,N_6742);
nor U7845 (N_7845,N_6100,N_6250);
xnor U7846 (N_7846,N_6984,N_6416);
nand U7847 (N_7847,N_6142,N_6350);
nand U7848 (N_7848,N_6088,N_6589);
nor U7849 (N_7849,N_6399,N_6349);
or U7850 (N_7850,N_6627,N_6038);
and U7851 (N_7851,N_6480,N_6667);
or U7852 (N_7852,N_6717,N_6308);
or U7853 (N_7853,N_6484,N_6019);
nor U7854 (N_7854,N_6597,N_6854);
nand U7855 (N_7855,N_6851,N_6288);
and U7856 (N_7856,N_6599,N_6689);
nor U7857 (N_7857,N_6842,N_6697);
and U7858 (N_7858,N_6095,N_6665);
and U7859 (N_7859,N_6933,N_6305);
nor U7860 (N_7860,N_6735,N_6917);
or U7861 (N_7861,N_6176,N_6295);
nor U7862 (N_7862,N_6892,N_6137);
and U7863 (N_7863,N_6838,N_6468);
nand U7864 (N_7864,N_6991,N_6159);
xor U7865 (N_7865,N_6313,N_6340);
nand U7866 (N_7866,N_6226,N_6930);
nor U7867 (N_7867,N_6916,N_6041);
or U7868 (N_7868,N_6212,N_6042);
and U7869 (N_7869,N_6566,N_6743);
and U7870 (N_7870,N_6455,N_6316);
nand U7871 (N_7871,N_6494,N_6523);
and U7872 (N_7872,N_6684,N_6496);
nand U7873 (N_7873,N_6076,N_6583);
nor U7874 (N_7874,N_6972,N_6593);
or U7875 (N_7875,N_6472,N_6048);
or U7876 (N_7876,N_6961,N_6839);
nand U7877 (N_7877,N_6302,N_6795);
and U7878 (N_7878,N_6501,N_6726);
xor U7879 (N_7879,N_6802,N_6016);
nand U7880 (N_7880,N_6028,N_6170);
and U7881 (N_7881,N_6858,N_6886);
nand U7882 (N_7882,N_6067,N_6907);
or U7883 (N_7883,N_6935,N_6175);
or U7884 (N_7884,N_6100,N_6959);
xor U7885 (N_7885,N_6876,N_6277);
or U7886 (N_7886,N_6863,N_6538);
or U7887 (N_7887,N_6745,N_6271);
nor U7888 (N_7888,N_6050,N_6196);
nand U7889 (N_7889,N_6339,N_6202);
xnor U7890 (N_7890,N_6613,N_6509);
and U7891 (N_7891,N_6240,N_6944);
nor U7892 (N_7892,N_6052,N_6691);
and U7893 (N_7893,N_6257,N_6272);
and U7894 (N_7894,N_6410,N_6969);
or U7895 (N_7895,N_6986,N_6760);
nor U7896 (N_7896,N_6034,N_6256);
nand U7897 (N_7897,N_6040,N_6674);
or U7898 (N_7898,N_6267,N_6596);
or U7899 (N_7899,N_6706,N_6404);
nand U7900 (N_7900,N_6229,N_6886);
nand U7901 (N_7901,N_6973,N_6313);
or U7902 (N_7902,N_6881,N_6566);
nor U7903 (N_7903,N_6014,N_6891);
and U7904 (N_7904,N_6437,N_6042);
or U7905 (N_7905,N_6770,N_6841);
xnor U7906 (N_7906,N_6235,N_6985);
and U7907 (N_7907,N_6711,N_6137);
nor U7908 (N_7908,N_6458,N_6556);
nor U7909 (N_7909,N_6821,N_6567);
nand U7910 (N_7910,N_6516,N_6125);
xor U7911 (N_7911,N_6226,N_6271);
and U7912 (N_7912,N_6653,N_6566);
or U7913 (N_7913,N_6658,N_6014);
and U7914 (N_7914,N_6371,N_6116);
and U7915 (N_7915,N_6512,N_6756);
or U7916 (N_7916,N_6254,N_6073);
xnor U7917 (N_7917,N_6387,N_6936);
or U7918 (N_7918,N_6994,N_6227);
nor U7919 (N_7919,N_6272,N_6853);
or U7920 (N_7920,N_6654,N_6215);
nor U7921 (N_7921,N_6746,N_6384);
xor U7922 (N_7922,N_6689,N_6676);
nand U7923 (N_7923,N_6655,N_6142);
xnor U7924 (N_7924,N_6681,N_6047);
nor U7925 (N_7925,N_6311,N_6432);
nor U7926 (N_7926,N_6413,N_6382);
nand U7927 (N_7927,N_6418,N_6199);
or U7928 (N_7928,N_6781,N_6049);
xnor U7929 (N_7929,N_6201,N_6222);
nand U7930 (N_7930,N_6580,N_6015);
and U7931 (N_7931,N_6878,N_6346);
nand U7932 (N_7932,N_6451,N_6478);
nor U7933 (N_7933,N_6518,N_6846);
or U7934 (N_7934,N_6785,N_6998);
or U7935 (N_7935,N_6035,N_6551);
and U7936 (N_7936,N_6929,N_6442);
nand U7937 (N_7937,N_6939,N_6667);
or U7938 (N_7938,N_6325,N_6744);
nor U7939 (N_7939,N_6434,N_6988);
or U7940 (N_7940,N_6503,N_6123);
xor U7941 (N_7941,N_6967,N_6069);
nor U7942 (N_7942,N_6260,N_6444);
nor U7943 (N_7943,N_6137,N_6538);
xor U7944 (N_7944,N_6922,N_6647);
nor U7945 (N_7945,N_6105,N_6534);
and U7946 (N_7946,N_6321,N_6813);
and U7947 (N_7947,N_6521,N_6644);
nor U7948 (N_7948,N_6323,N_6795);
nor U7949 (N_7949,N_6888,N_6146);
nor U7950 (N_7950,N_6912,N_6933);
or U7951 (N_7951,N_6932,N_6106);
and U7952 (N_7952,N_6203,N_6581);
nand U7953 (N_7953,N_6955,N_6582);
and U7954 (N_7954,N_6114,N_6622);
and U7955 (N_7955,N_6810,N_6819);
nand U7956 (N_7956,N_6398,N_6571);
or U7957 (N_7957,N_6172,N_6646);
or U7958 (N_7958,N_6783,N_6918);
nor U7959 (N_7959,N_6172,N_6047);
nor U7960 (N_7960,N_6122,N_6209);
or U7961 (N_7961,N_6281,N_6888);
and U7962 (N_7962,N_6533,N_6196);
or U7963 (N_7963,N_6573,N_6478);
nor U7964 (N_7964,N_6952,N_6415);
nor U7965 (N_7965,N_6472,N_6144);
nand U7966 (N_7966,N_6674,N_6884);
nor U7967 (N_7967,N_6266,N_6246);
and U7968 (N_7968,N_6524,N_6600);
nand U7969 (N_7969,N_6518,N_6997);
nor U7970 (N_7970,N_6873,N_6695);
nor U7971 (N_7971,N_6896,N_6001);
and U7972 (N_7972,N_6659,N_6336);
nand U7973 (N_7973,N_6113,N_6357);
nor U7974 (N_7974,N_6041,N_6273);
and U7975 (N_7975,N_6503,N_6800);
nand U7976 (N_7976,N_6440,N_6270);
and U7977 (N_7977,N_6781,N_6642);
nand U7978 (N_7978,N_6504,N_6758);
and U7979 (N_7979,N_6068,N_6981);
nor U7980 (N_7980,N_6357,N_6200);
nor U7981 (N_7981,N_6169,N_6864);
xor U7982 (N_7982,N_6778,N_6606);
xor U7983 (N_7983,N_6808,N_6653);
and U7984 (N_7984,N_6052,N_6360);
nand U7985 (N_7985,N_6826,N_6882);
or U7986 (N_7986,N_6054,N_6876);
xor U7987 (N_7987,N_6987,N_6272);
or U7988 (N_7988,N_6405,N_6648);
nand U7989 (N_7989,N_6499,N_6486);
nand U7990 (N_7990,N_6223,N_6340);
and U7991 (N_7991,N_6102,N_6691);
and U7992 (N_7992,N_6427,N_6229);
nand U7993 (N_7993,N_6817,N_6930);
nand U7994 (N_7994,N_6154,N_6699);
xnor U7995 (N_7995,N_6802,N_6833);
nand U7996 (N_7996,N_6087,N_6982);
or U7997 (N_7997,N_6373,N_6253);
or U7998 (N_7998,N_6304,N_6681);
and U7999 (N_7999,N_6277,N_6667);
or U8000 (N_8000,N_7693,N_7969);
xnor U8001 (N_8001,N_7422,N_7747);
or U8002 (N_8002,N_7062,N_7712);
or U8003 (N_8003,N_7626,N_7997);
and U8004 (N_8004,N_7159,N_7613);
or U8005 (N_8005,N_7427,N_7357);
and U8006 (N_8006,N_7849,N_7746);
nor U8007 (N_8007,N_7800,N_7855);
nand U8008 (N_8008,N_7103,N_7483);
xor U8009 (N_8009,N_7112,N_7371);
nor U8010 (N_8010,N_7329,N_7199);
and U8011 (N_8011,N_7177,N_7525);
nand U8012 (N_8012,N_7869,N_7610);
nor U8013 (N_8013,N_7774,N_7081);
or U8014 (N_8014,N_7918,N_7479);
nor U8015 (N_8015,N_7531,N_7523);
nor U8016 (N_8016,N_7415,N_7729);
or U8017 (N_8017,N_7173,N_7735);
and U8018 (N_8018,N_7826,N_7416);
nor U8019 (N_8019,N_7827,N_7818);
and U8020 (N_8020,N_7726,N_7156);
and U8021 (N_8021,N_7792,N_7309);
xor U8022 (N_8022,N_7940,N_7488);
or U8023 (N_8023,N_7899,N_7717);
and U8024 (N_8024,N_7303,N_7473);
or U8025 (N_8025,N_7300,N_7544);
or U8026 (N_8026,N_7618,N_7344);
nor U8027 (N_8027,N_7314,N_7218);
xor U8028 (N_8028,N_7652,N_7897);
or U8029 (N_8029,N_7679,N_7226);
xnor U8030 (N_8030,N_7202,N_7882);
or U8031 (N_8031,N_7625,N_7343);
or U8032 (N_8032,N_7521,N_7588);
nor U8033 (N_8033,N_7541,N_7326);
nand U8034 (N_8034,N_7246,N_7280);
or U8035 (N_8035,N_7787,N_7537);
or U8036 (N_8036,N_7168,N_7130);
and U8037 (N_8037,N_7465,N_7619);
xnor U8038 (N_8038,N_7392,N_7509);
xor U8039 (N_8039,N_7606,N_7706);
or U8040 (N_8040,N_7578,N_7466);
or U8041 (N_8041,N_7359,N_7165);
xnor U8042 (N_8042,N_7086,N_7938);
nand U8043 (N_8043,N_7463,N_7437);
xnor U8044 (N_8044,N_7272,N_7066);
and U8045 (N_8045,N_7064,N_7189);
nand U8046 (N_8046,N_7347,N_7510);
or U8047 (N_8047,N_7454,N_7838);
xnor U8048 (N_8048,N_7829,N_7047);
nor U8049 (N_8049,N_7658,N_7305);
nor U8050 (N_8050,N_7991,N_7602);
nand U8051 (N_8051,N_7954,N_7023);
xnor U8052 (N_8052,N_7121,N_7724);
nand U8053 (N_8053,N_7327,N_7843);
and U8054 (N_8054,N_7686,N_7768);
or U8055 (N_8055,N_7024,N_7571);
nor U8056 (N_8056,N_7699,N_7029);
and U8057 (N_8057,N_7126,N_7580);
or U8058 (N_8058,N_7681,N_7119);
nor U8059 (N_8059,N_7232,N_7971);
and U8060 (N_8060,N_7780,N_7074);
nor U8061 (N_8061,N_7115,N_7338);
nand U8062 (N_8062,N_7900,N_7836);
xor U8063 (N_8063,N_7958,N_7663);
or U8064 (N_8064,N_7756,N_7822);
or U8065 (N_8065,N_7102,N_7834);
and U8066 (N_8066,N_7552,N_7017);
nor U8067 (N_8067,N_7754,N_7150);
nor U8068 (N_8068,N_7925,N_7803);
nor U8069 (N_8069,N_7727,N_7721);
nand U8070 (N_8070,N_7627,N_7773);
nand U8071 (N_8071,N_7378,N_7253);
or U8072 (N_8072,N_7381,N_7442);
nand U8073 (N_8073,N_7451,N_7315);
and U8074 (N_8074,N_7373,N_7157);
nor U8075 (N_8075,N_7453,N_7669);
or U8076 (N_8076,N_7399,N_7917);
or U8077 (N_8077,N_7198,N_7500);
nor U8078 (N_8078,N_7242,N_7876);
xnor U8079 (N_8079,N_7716,N_7894);
or U8080 (N_8080,N_7678,N_7527);
and U8081 (N_8081,N_7075,N_7247);
xor U8082 (N_8082,N_7092,N_7052);
xor U8083 (N_8083,N_7631,N_7937);
and U8084 (N_8084,N_7009,N_7425);
nand U8085 (N_8085,N_7128,N_7947);
nand U8086 (N_8086,N_7923,N_7944);
and U8087 (N_8087,N_7421,N_7603);
nor U8088 (N_8088,N_7733,N_7697);
and U8089 (N_8089,N_7409,N_7594);
xor U8090 (N_8090,N_7151,N_7161);
nand U8091 (N_8091,N_7375,N_7034);
or U8092 (N_8092,N_7858,N_7880);
and U8093 (N_8093,N_7291,N_7585);
nor U8094 (N_8094,N_7290,N_7931);
and U8095 (N_8095,N_7149,N_7820);
nor U8096 (N_8096,N_7258,N_7597);
nand U8097 (N_8097,N_7576,N_7720);
and U8098 (N_8098,N_7845,N_7654);
nor U8099 (N_8099,N_7030,N_7930);
nor U8100 (N_8100,N_7551,N_7348);
nor U8101 (N_8101,N_7601,N_7432);
nor U8102 (N_8102,N_7942,N_7659);
or U8103 (N_8103,N_7703,N_7864);
or U8104 (N_8104,N_7692,N_7705);
xor U8105 (N_8105,N_7445,N_7815);
and U8106 (N_8106,N_7817,N_7142);
and U8107 (N_8107,N_7194,N_7532);
nor U8108 (N_8108,N_7584,N_7837);
or U8109 (N_8109,N_7553,N_7210);
and U8110 (N_8110,N_7682,N_7653);
or U8111 (N_8111,N_7105,N_7251);
nor U8112 (N_8112,N_7609,N_7021);
or U8113 (N_8113,N_7046,N_7033);
nand U8114 (N_8114,N_7438,N_7436);
and U8115 (N_8115,N_7111,N_7857);
nand U8116 (N_8116,N_7561,N_7163);
and U8117 (N_8117,N_7129,N_7734);
or U8118 (N_8118,N_7006,N_7043);
nand U8119 (N_8119,N_7943,N_7885);
nor U8120 (N_8120,N_7002,N_7387);
and U8121 (N_8121,N_7700,N_7426);
or U8122 (N_8122,N_7223,N_7556);
xor U8123 (N_8123,N_7853,N_7494);
xnor U8124 (N_8124,N_7162,N_7896);
and U8125 (N_8125,N_7572,N_7536);
or U8126 (N_8126,N_7784,N_7760);
nand U8127 (N_8127,N_7228,N_7646);
xor U8128 (N_8128,N_7713,N_7830);
nand U8129 (N_8129,N_7833,N_7673);
nand U8130 (N_8130,N_7311,N_7898);
nor U8131 (N_8131,N_7263,N_7516);
nand U8132 (N_8132,N_7863,N_7252);
nand U8133 (N_8133,N_7546,N_7337);
or U8134 (N_8134,N_7179,N_7522);
nor U8135 (N_8135,N_7123,N_7502);
xor U8136 (N_8136,N_7797,N_7887);
and U8137 (N_8137,N_7981,N_7063);
and U8138 (N_8138,N_7292,N_7261);
and U8139 (N_8139,N_7020,N_7100);
nand U8140 (N_8140,N_7146,N_7262);
nand U8141 (N_8141,N_7404,N_7236);
nor U8142 (N_8142,N_7901,N_7846);
or U8143 (N_8143,N_7860,N_7091);
nand U8144 (N_8144,N_7751,N_7630);
or U8145 (N_8145,N_7213,N_7406);
or U8146 (N_8146,N_7053,N_7848);
xor U8147 (N_8147,N_7497,N_7979);
nand U8148 (N_8148,N_7785,N_7281);
and U8149 (N_8149,N_7358,N_7983);
or U8150 (N_8150,N_7147,N_7615);
and U8151 (N_8151,N_7195,N_7957);
and U8152 (N_8152,N_7928,N_7317);
and U8153 (N_8153,N_7568,N_7581);
or U8154 (N_8154,N_7059,N_7737);
xnor U8155 (N_8155,N_7336,N_7484);
nand U8156 (N_8156,N_7127,N_7569);
nand U8157 (N_8157,N_7040,N_7487);
nand U8158 (N_8158,N_7794,N_7999);
nand U8159 (N_8159,N_7968,N_7011);
xnor U8160 (N_8160,N_7139,N_7191);
or U8161 (N_8161,N_7694,N_7482);
and U8162 (N_8162,N_7424,N_7701);
xnor U8163 (N_8163,N_7916,N_7616);
nor U8164 (N_8164,N_7519,N_7816);
xor U8165 (N_8165,N_7459,N_7428);
nor U8166 (N_8166,N_7992,N_7757);
nand U8167 (N_8167,N_7206,N_7116);
or U8168 (N_8168,N_7443,N_7271);
nor U8169 (N_8169,N_7605,N_7665);
xor U8170 (N_8170,N_7219,N_7138);
and U8171 (N_8171,N_7675,N_7172);
or U8172 (N_8172,N_7240,N_7941);
nor U8173 (N_8173,N_7069,N_7078);
or U8174 (N_8174,N_7985,N_7810);
and U8175 (N_8175,N_7499,N_7225);
nor U8176 (N_8176,N_7645,N_7909);
and U8177 (N_8177,N_7554,N_7579);
and U8178 (N_8178,N_7691,N_7823);
nand U8179 (N_8179,N_7623,N_7963);
or U8180 (N_8180,N_7495,N_7976);
nor U8181 (N_8181,N_7286,N_7256);
and U8182 (N_8182,N_7014,N_7470);
nor U8183 (N_8183,N_7840,N_7352);
and U8184 (N_8184,N_7770,N_7158);
and U8185 (N_8185,N_7506,N_7423);
or U8186 (N_8186,N_7259,N_7513);
and U8187 (N_8187,N_7684,N_7084);
and U8188 (N_8188,N_7489,N_7458);
or U8189 (N_8189,N_7222,N_7617);
and U8190 (N_8190,N_7769,N_7695);
nor U8191 (N_8191,N_7176,N_7341);
and U8192 (N_8192,N_7964,N_7611);
nor U8193 (N_8193,N_7217,N_7389);
nor U8194 (N_8194,N_7961,N_7676);
nor U8195 (N_8195,N_7388,N_7257);
xnor U8196 (N_8196,N_7154,N_7362);
xor U8197 (N_8197,N_7595,N_7268);
nor U8198 (N_8198,N_7591,N_7071);
and U8199 (N_8199,N_7562,N_7211);
nand U8200 (N_8200,N_7793,N_7190);
xor U8201 (N_8201,N_7744,N_7790);
and U8202 (N_8202,N_7634,N_7779);
nand U8203 (N_8203,N_7614,N_7874);
nand U8204 (N_8204,N_7323,N_7235);
or U8205 (N_8205,N_7927,N_7902);
and U8206 (N_8206,N_7471,N_7660);
nand U8207 (N_8207,N_7316,N_7908);
nand U8208 (N_8208,N_7950,N_7032);
nor U8209 (N_8209,N_7227,N_7411);
xnor U8210 (N_8210,N_7913,N_7996);
nor U8211 (N_8211,N_7639,N_7915);
nor U8212 (N_8212,N_7312,N_7106);
and U8213 (N_8213,N_7277,N_7385);
nor U8214 (N_8214,N_7383,N_7035);
nor U8215 (N_8215,N_7590,N_7514);
nor U8216 (N_8216,N_7905,N_7450);
nand U8217 (N_8217,N_7197,N_7807);
and U8218 (N_8218,N_7956,N_7393);
or U8219 (N_8219,N_7145,N_7564);
nand U8220 (N_8220,N_7073,N_7866);
and U8221 (N_8221,N_7640,N_7775);
or U8222 (N_8222,N_7233,N_7125);
nor U8223 (N_8223,N_7267,N_7295);
nor U8224 (N_8224,N_7655,N_7798);
or U8225 (N_8225,N_7629,N_7299);
or U8226 (N_8226,N_7248,N_7216);
nor U8227 (N_8227,N_7320,N_7704);
or U8228 (N_8228,N_7641,N_7975);
and U8229 (N_8229,N_7175,N_7349);
nor U8230 (N_8230,N_7587,N_7080);
xor U8231 (N_8231,N_7056,N_7910);
or U8232 (N_8232,N_7637,N_7856);
nand U8233 (N_8233,N_7596,N_7766);
nor U8234 (N_8234,N_7265,N_7282);
nor U8235 (N_8235,N_7410,N_7632);
or U8236 (N_8236,N_7457,N_7408);
nor U8237 (N_8237,N_7668,N_7517);
and U8238 (N_8238,N_7397,N_7209);
and U8239 (N_8239,N_7906,N_7384);
and U8240 (N_8240,N_7872,N_7953);
or U8241 (N_8241,N_7831,N_7934);
nand U8242 (N_8242,N_7104,N_7351);
or U8243 (N_8243,N_7284,N_7708);
nand U8244 (N_8244,N_7504,N_7948);
nor U8245 (N_8245,N_7844,N_7369);
nor U8246 (N_8246,N_7143,N_7994);
or U8247 (N_8247,N_7288,N_7333);
and U8248 (N_8248,N_7360,N_7307);
and U8249 (N_8249,N_7865,N_7109);
and U8250 (N_8250,N_7714,N_7243);
and U8251 (N_8251,N_7003,N_7481);
or U8252 (N_8252,N_7061,N_7604);
nand U8253 (N_8253,N_7013,N_7196);
nor U8254 (N_8254,N_7220,N_7988);
and U8255 (N_8255,N_7503,N_7097);
nor U8256 (N_8256,N_7090,N_7842);
nand U8257 (N_8257,N_7296,N_7624);
or U8258 (N_8258,N_7980,N_7753);
nor U8259 (N_8259,N_7065,N_7814);
nor U8260 (N_8260,N_7742,N_7302);
nor U8261 (N_8261,N_7440,N_7083);
and U8262 (N_8262,N_7635,N_7401);
and U8263 (N_8263,N_7386,N_7044);
nand U8264 (N_8264,N_7741,N_7390);
or U8265 (N_8265,N_7926,N_7835);
nand U8266 (N_8266,N_7722,N_7117);
and U8267 (N_8267,N_7093,N_7832);
and U8268 (N_8268,N_7374,N_7702);
nand U8269 (N_8269,N_7873,N_7802);
nor U8270 (N_8270,N_7241,N_7435);
nor U8271 (N_8271,N_7085,N_7936);
nand U8272 (N_8272,N_7019,N_7847);
nand U8273 (N_8273,N_7322,N_7868);
or U8274 (N_8274,N_7368,N_7205);
and U8275 (N_8275,N_7862,N_7650);
nand U8276 (N_8276,N_7186,N_7528);
nor U8277 (N_8277,N_7412,N_7743);
nor U8278 (N_8278,N_7577,N_7952);
nand U8279 (N_8279,N_7042,N_7221);
xnor U8280 (N_8280,N_7345,N_7526);
nor U8281 (N_8281,N_7643,N_7407);
and U8282 (N_8282,N_7871,N_7318);
and U8283 (N_8283,N_7549,N_7728);
nand U8284 (N_8284,N_7372,N_7558);
nand U8285 (N_8285,N_7657,N_7054);
nand U8286 (N_8286,N_7474,N_7285);
or U8287 (N_8287,N_7400,N_7113);
or U8288 (N_8288,N_7745,N_7204);
xor U8289 (N_8289,N_7932,N_7077);
xor U8290 (N_8290,N_7464,N_7039);
or U8291 (N_8291,N_7539,N_7215);
nor U8292 (N_8292,N_7621,N_7171);
and U8293 (N_8293,N_7783,N_7808);
or U8294 (N_8294,N_7582,N_7680);
and U8295 (N_8295,N_7739,N_7007);
and U8296 (N_8296,N_7608,N_7430);
nor U8297 (N_8297,N_7662,N_7970);
nor U8298 (N_8298,N_7380,N_7183);
nor U8299 (N_8299,N_7912,N_7356);
and U8300 (N_8300,N_7824,N_7004);
xnor U8301 (N_8301,N_7907,N_7110);
or U8302 (N_8302,N_7405,N_7781);
nor U8303 (N_8303,N_7325,N_7575);
or U8304 (N_8304,N_7642,N_7306);
and U8305 (N_8305,N_7342,N_7886);
nand U8306 (N_8306,N_7759,N_7067);
nor U8307 (N_8307,N_7330,N_7439);
or U8308 (N_8308,N_7732,N_7192);
xor U8309 (N_8309,N_7238,N_7529);
nor U8310 (N_8310,N_7960,N_7565);
nor U8311 (N_8311,N_7607,N_7879);
or U8312 (N_8312,N_7018,N_7990);
nand U8313 (N_8313,N_7155,N_7518);
nand U8314 (N_8314,N_7244,N_7396);
and U8315 (N_8315,N_7841,N_7530);
or U8316 (N_8316,N_7612,N_7599);
or U8317 (N_8317,N_7730,N_7283);
nor U8318 (N_8318,N_7683,N_7167);
and U8319 (N_8319,N_7049,N_7332);
nand U8320 (N_8320,N_7972,N_7468);
xnor U8321 (N_8321,N_7715,N_7082);
nor U8322 (N_8322,N_7949,N_7542);
and U8323 (N_8323,N_7382,N_7016);
and U8324 (N_8324,N_7098,N_7805);
nor U8325 (N_8325,N_7891,N_7279);
nor U8326 (N_8326,N_7812,N_7939);
and U8327 (N_8327,N_7696,N_7446);
nand U8328 (N_8328,N_7012,N_7709);
nand U8329 (N_8329,N_7764,N_7789);
and U8330 (N_8330,N_7184,N_7328);
and U8331 (N_8331,N_7496,N_7791);
nor U8332 (N_8332,N_7429,N_7738);
or U8333 (N_8333,N_7174,N_7152);
nor U8334 (N_8334,N_7144,N_7188);
nand U8335 (N_8335,N_7447,N_7586);
nand U8336 (N_8336,N_7593,N_7978);
and U8337 (N_8337,N_7274,N_7293);
nand U8338 (N_8338,N_7828,N_7566);
or U8339 (N_8339,N_7710,N_7687);
nor U8340 (N_8340,N_7962,N_7633);
nand U8341 (N_8341,N_7986,N_7533);
or U8342 (N_8342,N_7418,N_7353);
or U8343 (N_8343,N_7058,N_7308);
and U8344 (N_8344,N_7460,N_7664);
nand U8345 (N_8345,N_7324,N_7298);
nand U8346 (N_8346,N_7545,N_7433);
and U8347 (N_8347,N_7480,N_7573);
xor U8348 (N_8348,N_7079,N_7124);
or U8349 (N_8349,N_7355,N_7788);
or U8350 (N_8350,N_7001,N_7469);
nor U8351 (N_8351,N_7543,N_7214);
nand U8352 (N_8352,N_7203,N_7984);
and U8353 (N_8353,N_7088,N_7230);
nor U8354 (N_8354,N_7060,N_7431);
nor U8355 (N_8355,N_7461,N_7786);
and U8356 (N_8356,N_7859,N_7289);
nand U8357 (N_8357,N_7776,N_7249);
xnor U8358 (N_8358,N_7131,N_7935);
and U8359 (N_8359,N_7041,N_7557);
nand U8360 (N_8360,N_7895,N_7141);
nand U8361 (N_8361,N_7666,N_7711);
nor U8362 (N_8362,N_7638,N_7795);
nand U8363 (N_8363,N_7099,N_7364);
and U8364 (N_8364,N_7995,N_7998);
and U8365 (N_8365,N_7672,N_7264);
nor U8366 (N_8366,N_7051,N_7136);
and U8367 (N_8367,N_7391,N_7763);
xor U8368 (N_8368,N_7881,N_7031);
and U8369 (N_8369,N_7574,N_7698);
nand U8370 (N_8370,N_7132,N_7477);
xor U8371 (N_8371,N_7765,N_7892);
nand U8372 (N_8372,N_7321,N_7493);
nor U8373 (N_8373,N_7234,N_7015);
and U8374 (N_8374,N_7255,N_7010);
nor U8375 (N_8375,N_7160,N_7982);
nor U8376 (N_8376,N_7107,N_7933);
or U8377 (N_8377,N_7740,N_7507);
or U8378 (N_8378,N_7164,N_7661);
nand U8379 (N_8379,N_7850,N_7890);
nand U8380 (N_8380,N_7670,N_7379);
or U8381 (N_8381,N_7883,N_7920);
nand U8382 (N_8382,N_7273,N_7335);
and U8383 (N_8383,N_7101,N_7598);
xnor U8384 (N_8384,N_7821,N_7122);
nand U8385 (N_8385,N_7402,N_7945);
or U8386 (N_8386,N_7087,N_7114);
nor U8387 (N_8387,N_7589,N_7297);
and U8388 (N_8388,N_7153,N_7647);
or U8389 (N_8389,N_7045,N_7778);
nor U8390 (N_8390,N_7354,N_7365);
nand U8391 (N_8391,N_7889,N_7475);
nor U8392 (N_8392,N_7313,N_7534);
and U8393 (N_8393,N_7548,N_7540);
nand U8394 (N_8394,N_7875,N_7538);
and U8395 (N_8395,N_7276,N_7520);
xor U8396 (N_8396,N_7550,N_7563);
or U8397 (N_8397,N_7515,N_7148);
or U8398 (N_8398,N_7187,N_7094);
or U8399 (N_8399,N_7208,N_7854);
or U8400 (N_8400,N_7361,N_7755);
or U8401 (N_8401,N_7570,N_7260);
xor U8402 (N_8402,N_7772,N_7310);
xnor U8403 (N_8403,N_7182,N_7254);
nor U8404 (N_8404,N_7644,N_7767);
nor U8405 (N_8405,N_7367,N_7560);
nand U8406 (N_8406,N_7478,N_7796);
nand U8407 (N_8407,N_7096,N_7485);
nand U8408 (N_8408,N_7758,N_7270);
and U8409 (N_8409,N_7370,N_7275);
or U8410 (N_8410,N_7505,N_7559);
nor U8411 (N_8411,N_7736,N_7076);
and U8412 (N_8412,N_7028,N_7250);
or U8413 (N_8413,N_7108,N_7376);
or U8414 (N_8414,N_7201,N_7877);
and U8415 (N_8415,N_7048,N_7535);
nor U8416 (N_8416,N_7839,N_7799);
nand U8417 (N_8417,N_7861,N_7748);
or U8418 (N_8418,N_7237,N_7946);
nor U8419 (N_8419,N_7068,N_7649);
and U8420 (N_8420,N_7777,N_7987);
or U8421 (N_8421,N_7319,N_7037);
nand U8422 (N_8422,N_7231,N_7870);
nor U8423 (N_8423,N_7977,N_7973);
or U8424 (N_8424,N_7118,N_7022);
nor U8425 (N_8425,N_7133,N_7725);
and U8426 (N_8426,N_7414,N_7903);
nor U8427 (N_8427,N_7914,N_7620);
nor U8428 (N_8428,N_7967,N_7904);
and U8429 (N_8429,N_7000,N_7547);
xnor U8430 (N_8430,N_7304,N_7269);
or U8431 (N_8431,N_7825,N_7867);
nor U8432 (N_8432,N_7512,N_7038);
or U8433 (N_8433,N_7181,N_7811);
nor U8434 (N_8434,N_7363,N_7462);
nand U8435 (N_8435,N_7398,N_7301);
or U8436 (N_8436,N_7524,N_7413);
nor U8437 (N_8437,N_7685,N_7771);
nor U8438 (N_8438,N_7366,N_7555);
nor U8439 (N_8439,N_7472,N_7731);
and U8440 (N_8440,N_7026,N_7921);
nand U8441 (N_8441,N_7137,N_7070);
nor U8442 (N_8442,N_7501,N_7974);
nand U8443 (N_8443,N_7648,N_7339);
nor U8444 (N_8444,N_7350,N_7919);
xor U8445 (N_8445,N_7813,N_7911);
or U8446 (N_8446,N_7656,N_7508);
or U8447 (N_8447,N_7434,N_7511);
and U8448 (N_8448,N_7718,N_7095);
nand U8449 (N_8449,N_7456,N_7628);
or U8450 (N_8450,N_7036,N_7417);
nor U8451 (N_8451,N_7072,N_7878);
and U8452 (N_8452,N_7888,N_7207);
or U8453 (N_8453,N_7027,N_7965);
and U8454 (N_8454,N_7170,N_7135);
and U8455 (N_8455,N_7804,N_7120);
xor U8456 (N_8456,N_7651,N_7334);
nor U8457 (N_8457,N_7394,N_7498);
or U8458 (N_8458,N_7592,N_7467);
or U8459 (N_8459,N_7448,N_7490);
nor U8460 (N_8460,N_7600,N_7331);
or U8461 (N_8461,N_7005,N_7441);
and U8462 (N_8462,N_7340,N_7622);
nand U8463 (N_8463,N_7134,N_7025);
nand U8464 (N_8464,N_7723,N_7050);
or U8465 (N_8465,N_7346,N_7245);
nor U8466 (N_8466,N_7924,N_7966);
nand U8467 (N_8467,N_7239,N_7761);
nand U8468 (N_8468,N_7455,N_7667);
nor U8469 (N_8469,N_7707,N_7951);
xnor U8470 (N_8470,N_7185,N_7801);
nor U8471 (N_8471,N_7166,N_7419);
nand U8472 (N_8472,N_7169,N_7224);
xnor U8473 (N_8473,N_7089,N_7806);
nor U8474 (N_8474,N_7444,N_7278);
xnor U8475 (N_8475,N_7486,N_7929);
or U8476 (N_8476,N_7055,N_7492);
or U8477 (N_8477,N_7377,N_7452);
nor U8478 (N_8478,N_7762,N_7567);
and U8479 (N_8479,N_7750,N_7395);
and U8480 (N_8480,N_7449,N_7403);
and U8481 (N_8481,N_7851,N_7229);
nor U8482 (N_8482,N_7719,N_7212);
nor U8483 (N_8483,N_7689,N_7852);
and U8484 (N_8484,N_7294,N_7287);
nor U8485 (N_8485,N_7476,N_7688);
or U8486 (N_8486,N_7420,N_7674);
and U8487 (N_8487,N_7193,N_7819);
or U8488 (N_8488,N_7671,N_7752);
nor U8489 (N_8489,N_7266,N_7677);
nor U8490 (N_8490,N_7491,N_7782);
or U8491 (N_8491,N_7955,N_7140);
nand U8492 (N_8492,N_7922,N_7749);
nor U8493 (N_8493,N_7884,N_7583);
and U8494 (N_8494,N_7008,N_7809);
or U8495 (N_8495,N_7993,N_7057);
or U8496 (N_8496,N_7893,N_7180);
nand U8497 (N_8497,N_7690,N_7989);
or U8498 (N_8498,N_7178,N_7636);
and U8499 (N_8499,N_7200,N_7959);
nand U8500 (N_8500,N_7030,N_7046);
or U8501 (N_8501,N_7263,N_7231);
nor U8502 (N_8502,N_7586,N_7161);
nand U8503 (N_8503,N_7087,N_7276);
and U8504 (N_8504,N_7770,N_7305);
nor U8505 (N_8505,N_7070,N_7396);
nand U8506 (N_8506,N_7771,N_7906);
and U8507 (N_8507,N_7963,N_7761);
and U8508 (N_8508,N_7092,N_7687);
xnor U8509 (N_8509,N_7323,N_7826);
nand U8510 (N_8510,N_7577,N_7759);
nor U8511 (N_8511,N_7567,N_7036);
or U8512 (N_8512,N_7965,N_7604);
nor U8513 (N_8513,N_7395,N_7132);
nand U8514 (N_8514,N_7763,N_7558);
or U8515 (N_8515,N_7480,N_7212);
xnor U8516 (N_8516,N_7741,N_7413);
nand U8517 (N_8517,N_7369,N_7198);
xnor U8518 (N_8518,N_7780,N_7806);
nand U8519 (N_8519,N_7929,N_7095);
nand U8520 (N_8520,N_7076,N_7016);
xor U8521 (N_8521,N_7744,N_7511);
and U8522 (N_8522,N_7435,N_7150);
xnor U8523 (N_8523,N_7918,N_7811);
and U8524 (N_8524,N_7051,N_7141);
and U8525 (N_8525,N_7603,N_7685);
and U8526 (N_8526,N_7483,N_7946);
nand U8527 (N_8527,N_7966,N_7692);
nand U8528 (N_8528,N_7723,N_7063);
or U8529 (N_8529,N_7933,N_7568);
xor U8530 (N_8530,N_7262,N_7789);
nand U8531 (N_8531,N_7131,N_7456);
nor U8532 (N_8532,N_7333,N_7739);
nor U8533 (N_8533,N_7134,N_7377);
and U8534 (N_8534,N_7349,N_7334);
nand U8535 (N_8535,N_7124,N_7051);
and U8536 (N_8536,N_7793,N_7753);
or U8537 (N_8537,N_7375,N_7724);
xnor U8538 (N_8538,N_7238,N_7452);
nand U8539 (N_8539,N_7433,N_7399);
or U8540 (N_8540,N_7153,N_7114);
and U8541 (N_8541,N_7588,N_7635);
xnor U8542 (N_8542,N_7743,N_7980);
nand U8543 (N_8543,N_7505,N_7002);
and U8544 (N_8544,N_7613,N_7867);
and U8545 (N_8545,N_7881,N_7060);
xor U8546 (N_8546,N_7149,N_7674);
nor U8547 (N_8547,N_7967,N_7675);
or U8548 (N_8548,N_7920,N_7018);
or U8549 (N_8549,N_7836,N_7644);
and U8550 (N_8550,N_7591,N_7330);
xor U8551 (N_8551,N_7945,N_7272);
xor U8552 (N_8552,N_7395,N_7827);
or U8553 (N_8553,N_7784,N_7169);
or U8554 (N_8554,N_7816,N_7254);
nor U8555 (N_8555,N_7771,N_7057);
or U8556 (N_8556,N_7473,N_7731);
and U8557 (N_8557,N_7138,N_7848);
nand U8558 (N_8558,N_7875,N_7861);
and U8559 (N_8559,N_7431,N_7828);
and U8560 (N_8560,N_7325,N_7333);
xor U8561 (N_8561,N_7710,N_7830);
nor U8562 (N_8562,N_7286,N_7213);
and U8563 (N_8563,N_7886,N_7491);
xor U8564 (N_8564,N_7600,N_7493);
nand U8565 (N_8565,N_7607,N_7767);
and U8566 (N_8566,N_7587,N_7205);
nand U8567 (N_8567,N_7305,N_7344);
and U8568 (N_8568,N_7414,N_7134);
nor U8569 (N_8569,N_7370,N_7790);
and U8570 (N_8570,N_7339,N_7333);
nand U8571 (N_8571,N_7378,N_7213);
nor U8572 (N_8572,N_7032,N_7019);
nor U8573 (N_8573,N_7266,N_7037);
nand U8574 (N_8574,N_7495,N_7075);
or U8575 (N_8575,N_7224,N_7891);
nor U8576 (N_8576,N_7847,N_7394);
nand U8577 (N_8577,N_7330,N_7473);
nor U8578 (N_8578,N_7063,N_7381);
nor U8579 (N_8579,N_7037,N_7922);
and U8580 (N_8580,N_7371,N_7898);
and U8581 (N_8581,N_7590,N_7877);
and U8582 (N_8582,N_7793,N_7159);
nand U8583 (N_8583,N_7083,N_7565);
or U8584 (N_8584,N_7151,N_7436);
nor U8585 (N_8585,N_7069,N_7172);
nor U8586 (N_8586,N_7057,N_7662);
nand U8587 (N_8587,N_7803,N_7008);
nand U8588 (N_8588,N_7943,N_7231);
nor U8589 (N_8589,N_7384,N_7005);
or U8590 (N_8590,N_7575,N_7217);
or U8591 (N_8591,N_7042,N_7273);
and U8592 (N_8592,N_7582,N_7876);
or U8593 (N_8593,N_7526,N_7236);
nand U8594 (N_8594,N_7157,N_7918);
and U8595 (N_8595,N_7944,N_7776);
or U8596 (N_8596,N_7180,N_7455);
xnor U8597 (N_8597,N_7141,N_7496);
nand U8598 (N_8598,N_7147,N_7358);
and U8599 (N_8599,N_7408,N_7503);
or U8600 (N_8600,N_7894,N_7088);
and U8601 (N_8601,N_7507,N_7250);
or U8602 (N_8602,N_7726,N_7428);
nor U8603 (N_8603,N_7263,N_7942);
or U8604 (N_8604,N_7809,N_7650);
nand U8605 (N_8605,N_7192,N_7666);
or U8606 (N_8606,N_7177,N_7243);
or U8607 (N_8607,N_7878,N_7799);
and U8608 (N_8608,N_7418,N_7329);
or U8609 (N_8609,N_7773,N_7110);
or U8610 (N_8610,N_7098,N_7353);
or U8611 (N_8611,N_7491,N_7906);
or U8612 (N_8612,N_7396,N_7482);
xnor U8613 (N_8613,N_7515,N_7271);
and U8614 (N_8614,N_7583,N_7456);
and U8615 (N_8615,N_7490,N_7648);
and U8616 (N_8616,N_7864,N_7692);
or U8617 (N_8617,N_7513,N_7478);
or U8618 (N_8618,N_7535,N_7520);
nand U8619 (N_8619,N_7674,N_7985);
or U8620 (N_8620,N_7525,N_7705);
and U8621 (N_8621,N_7618,N_7737);
or U8622 (N_8622,N_7982,N_7129);
nand U8623 (N_8623,N_7553,N_7634);
xor U8624 (N_8624,N_7720,N_7349);
nand U8625 (N_8625,N_7864,N_7429);
and U8626 (N_8626,N_7511,N_7921);
nand U8627 (N_8627,N_7894,N_7690);
nor U8628 (N_8628,N_7863,N_7623);
nand U8629 (N_8629,N_7315,N_7824);
nor U8630 (N_8630,N_7993,N_7853);
nor U8631 (N_8631,N_7839,N_7383);
nor U8632 (N_8632,N_7139,N_7070);
and U8633 (N_8633,N_7046,N_7482);
xnor U8634 (N_8634,N_7117,N_7186);
xor U8635 (N_8635,N_7932,N_7292);
nand U8636 (N_8636,N_7665,N_7647);
and U8637 (N_8637,N_7890,N_7895);
nor U8638 (N_8638,N_7364,N_7229);
and U8639 (N_8639,N_7807,N_7598);
xor U8640 (N_8640,N_7612,N_7613);
nor U8641 (N_8641,N_7260,N_7721);
xnor U8642 (N_8642,N_7262,N_7462);
nand U8643 (N_8643,N_7742,N_7254);
nor U8644 (N_8644,N_7939,N_7833);
and U8645 (N_8645,N_7177,N_7183);
or U8646 (N_8646,N_7371,N_7515);
xor U8647 (N_8647,N_7531,N_7241);
and U8648 (N_8648,N_7992,N_7795);
nand U8649 (N_8649,N_7818,N_7639);
and U8650 (N_8650,N_7277,N_7435);
and U8651 (N_8651,N_7513,N_7254);
xor U8652 (N_8652,N_7411,N_7728);
and U8653 (N_8653,N_7549,N_7278);
nor U8654 (N_8654,N_7816,N_7520);
or U8655 (N_8655,N_7676,N_7620);
or U8656 (N_8656,N_7934,N_7886);
xnor U8657 (N_8657,N_7967,N_7126);
nor U8658 (N_8658,N_7118,N_7263);
or U8659 (N_8659,N_7742,N_7810);
or U8660 (N_8660,N_7569,N_7250);
and U8661 (N_8661,N_7101,N_7352);
xnor U8662 (N_8662,N_7093,N_7875);
nor U8663 (N_8663,N_7244,N_7907);
nor U8664 (N_8664,N_7161,N_7497);
xnor U8665 (N_8665,N_7919,N_7687);
nor U8666 (N_8666,N_7542,N_7947);
or U8667 (N_8667,N_7721,N_7456);
nor U8668 (N_8668,N_7975,N_7231);
nand U8669 (N_8669,N_7742,N_7154);
xnor U8670 (N_8670,N_7879,N_7296);
and U8671 (N_8671,N_7151,N_7931);
nor U8672 (N_8672,N_7600,N_7845);
or U8673 (N_8673,N_7315,N_7519);
nand U8674 (N_8674,N_7850,N_7292);
or U8675 (N_8675,N_7595,N_7682);
or U8676 (N_8676,N_7150,N_7384);
nand U8677 (N_8677,N_7554,N_7862);
and U8678 (N_8678,N_7351,N_7044);
or U8679 (N_8679,N_7308,N_7064);
nor U8680 (N_8680,N_7097,N_7749);
and U8681 (N_8681,N_7791,N_7884);
or U8682 (N_8682,N_7556,N_7510);
or U8683 (N_8683,N_7394,N_7435);
and U8684 (N_8684,N_7174,N_7873);
or U8685 (N_8685,N_7491,N_7989);
xor U8686 (N_8686,N_7455,N_7335);
and U8687 (N_8687,N_7810,N_7321);
and U8688 (N_8688,N_7086,N_7117);
and U8689 (N_8689,N_7080,N_7336);
nand U8690 (N_8690,N_7279,N_7630);
nand U8691 (N_8691,N_7159,N_7576);
and U8692 (N_8692,N_7262,N_7169);
nor U8693 (N_8693,N_7493,N_7470);
and U8694 (N_8694,N_7421,N_7157);
or U8695 (N_8695,N_7515,N_7147);
nor U8696 (N_8696,N_7971,N_7881);
and U8697 (N_8697,N_7221,N_7538);
xnor U8698 (N_8698,N_7970,N_7474);
nand U8699 (N_8699,N_7147,N_7324);
nand U8700 (N_8700,N_7682,N_7900);
and U8701 (N_8701,N_7310,N_7375);
or U8702 (N_8702,N_7622,N_7034);
or U8703 (N_8703,N_7030,N_7000);
nor U8704 (N_8704,N_7102,N_7609);
nand U8705 (N_8705,N_7555,N_7054);
or U8706 (N_8706,N_7495,N_7185);
nand U8707 (N_8707,N_7184,N_7609);
and U8708 (N_8708,N_7877,N_7625);
or U8709 (N_8709,N_7806,N_7321);
nor U8710 (N_8710,N_7086,N_7941);
or U8711 (N_8711,N_7978,N_7165);
nor U8712 (N_8712,N_7252,N_7636);
xor U8713 (N_8713,N_7270,N_7237);
and U8714 (N_8714,N_7757,N_7181);
and U8715 (N_8715,N_7722,N_7806);
and U8716 (N_8716,N_7951,N_7491);
or U8717 (N_8717,N_7120,N_7428);
nand U8718 (N_8718,N_7980,N_7340);
and U8719 (N_8719,N_7760,N_7079);
xnor U8720 (N_8720,N_7384,N_7577);
nand U8721 (N_8721,N_7002,N_7175);
nor U8722 (N_8722,N_7938,N_7701);
and U8723 (N_8723,N_7729,N_7901);
and U8724 (N_8724,N_7262,N_7977);
nor U8725 (N_8725,N_7780,N_7170);
nor U8726 (N_8726,N_7621,N_7521);
and U8727 (N_8727,N_7745,N_7734);
or U8728 (N_8728,N_7454,N_7611);
and U8729 (N_8729,N_7843,N_7667);
nor U8730 (N_8730,N_7375,N_7125);
or U8731 (N_8731,N_7118,N_7112);
and U8732 (N_8732,N_7650,N_7757);
nand U8733 (N_8733,N_7985,N_7068);
and U8734 (N_8734,N_7201,N_7886);
or U8735 (N_8735,N_7362,N_7205);
and U8736 (N_8736,N_7456,N_7551);
nor U8737 (N_8737,N_7543,N_7884);
nand U8738 (N_8738,N_7010,N_7008);
and U8739 (N_8739,N_7288,N_7965);
nand U8740 (N_8740,N_7304,N_7830);
or U8741 (N_8741,N_7490,N_7605);
or U8742 (N_8742,N_7596,N_7297);
or U8743 (N_8743,N_7337,N_7142);
or U8744 (N_8744,N_7506,N_7015);
and U8745 (N_8745,N_7843,N_7645);
nor U8746 (N_8746,N_7604,N_7875);
and U8747 (N_8747,N_7798,N_7761);
nor U8748 (N_8748,N_7548,N_7444);
or U8749 (N_8749,N_7083,N_7278);
nand U8750 (N_8750,N_7930,N_7758);
nor U8751 (N_8751,N_7047,N_7801);
nor U8752 (N_8752,N_7061,N_7454);
nor U8753 (N_8753,N_7576,N_7730);
nor U8754 (N_8754,N_7001,N_7445);
and U8755 (N_8755,N_7880,N_7948);
nor U8756 (N_8756,N_7298,N_7174);
nor U8757 (N_8757,N_7237,N_7373);
nor U8758 (N_8758,N_7383,N_7901);
and U8759 (N_8759,N_7662,N_7135);
and U8760 (N_8760,N_7278,N_7862);
nand U8761 (N_8761,N_7401,N_7486);
xor U8762 (N_8762,N_7017,N_7257);
nand U8763 (N_8763,N_7965,N_7885);
nor U8764 (N_8764,N_7829,N_7192);
and U8765 (N_8765,N_7524,N_7781);
nor U8766 (N_8766,N_7681,N_7235);
nand U8767 (N_8767,N_7415,N_7522);
or U8768 (N_8768,N_7861,N_7094);
nor U8769 (N_8769,N_7958,N_7038);
xor U8770 (N_8770,N_7067,N_7678);
and U8771 (N_8771,N_7611,N_7691);
nand U8772 (N_8772,N_7844,N_7588);
xor U8773 (N_8773,N_7230,N_7020);
nand U8774 (N_8774,N_7620,N_7362);
or U8775 (N_8775,N_7812,N_7971);
and U8776 (N_8776,N_7123,N_7071);
or U8777 (N_8777,N_7169,N_7686);
nor U8778 (N_8778,N_7494,N_7912);
and U8779 (N_8779,N_7581,N_7605);
xnor U8780 (N_8780,N_7603,N_7800);
or U8781 (N_8781,N_7787,N_7232);
xor U8782 (N_8782,N_7885,N_7267);
xnor U8783 (N_8783,N_7480,N_7390);
nand U8784 (N_8784,N_7945,N_7646);
or U8785 (N_8785,N_7961,N_7564);
and U8786 (N_8786,N_7559,N_7024);
nor U8787 (N_8787,N_7332,N_7650);
or U8788 (N_8788,N_7162,N_7877);
and U8789 (N_8789,N_7416,N_7362);
nor U8790 (N_8790,N_7421,N_7539);
or U8791 (N_8791,N_7615,N_7120);
nand U8792 (N_8792,N_7111,N_7834);
nor U8793 (N_8793,N_7438,N_7840);
nand U8794 (N_8794,N_7049,N_7251);
nand U8795 (N_8795,N_7343,N_7694);
nor U8796 (N_8796,N_7593,N_7726);
xor U8797 (N_8797,N_7971,N_7226);
nor U8798 (N_8798,N_7143,N_7650);
nor U8799 (N_8799,N_7140,N_7192);
and U8800 (N_8800,N_7999,N_7934);
nor U8801 (N_8801,N_7823,N_7177);
or U8802 (N_8802,N_7065,N_7638);
xor U8803 (N_8803,N_7300,N_7910);
nand U8804 (N_8804,N_7263,N_7222);
or U8805 (N_8805,N_7017,N_7449);
nand U8806 (N_8806,N_7986,N_7721);
nor U8807 (N_8807,N_7868,N_7001);
and U8808 (N_8808,N_7939,N_7963);
or U8809 (N_8809,N_7119,N_7095);
nand U8810 (N_8810,N_7279,N_7073);
nor U8811 (N_8811,N_7650,N_7697);
or U8812 (N_8812,N_7434,N_7688);
nand U8813 (N_8813,N_7305,N_7141);
or U8814 (N_8814,N_7071,N_7002);
and U8815 (N_8815,N_7932,N_7780);
or U8816 (N_8816,N_7293,N_7413);
nor U8817 (N_8817,N_7972,N_7437);
and U8818 (N_8818,N_7477,N_7047);
or U8819 (N_8819,N_7309,N_7790);
nor U8820 (N_8820,N_7264,N_7304);
and U8821 (N_8821,N_7724,N_7639);
and U8822 (N_8822,N_7373,N_7374);
nor U8823 (N_8823,N_7081,N_7384);
nor U8824 (N_8824,N_7154,N_7306);
nand U8825 (N_8825,N_7778,N_7583);
and U8826 (N_8826,N_7970,N_7042);
nor U8827 (N_8827,N_7649,N_7258);
nor U8828 (N_8828,N_7143,N_7592);
and U8829 (N_8829,N_7003,N_7371);
or U8830 (N_8830,N_7526,N_7759);
xnor U8831 (N_8831,N_7624,N_7237);
nor U8832 (N_8832,N_7875,N_7576);
xor U8833 (N_8833,N_7878,N_7044);
or U8834 (N_8834,N_7062,N_7479);
nor U8835 (N_8835,N_7155,N_7993);
nand U8836 (N_8836,N_7672,N_7885);
and U8837 (N_8837,N_7125,N_7292);
or U8838 (N_8838,N_7007,N_7542);
or U8839 (N_8839,N_7327,N_7035);
nor U8840 (N_8840,N_7681,N_7558);
or U8841 (N_8841,N_7522,N_7050);
or U8842 (N_8842,N_7887,N_7923);
nor U8843 (N_8843,N_7678,N_7353);
or U8844 (N_8844,N_7494,N_7806);
nand U8845 (N_8845,N_7865,N_7462);
nand U8846 (N_8846,N_7514,N_7390);
xnor U8847 (N_8847,N_7677,N_7931);
and U8848 (N_8848,N_7973,N_7794);
nor U8849 (N_8849,N_7813,N_7228);
or U8850 (N_8850,N_7926,N_7792);
or U8851 (N_8851,N_7412,N_7380);
and U8852 (N_8852,N_7819,N_7878);
xnor U8853 (N_8853,N_7684,N_7851);
nor U8854 (N_8854,N_7336,N_7083);
xnor U8855 (N_8855,N_7351,N_7246);
and U8856 (N_8856,N_7796,N_7078);
nand U8857 (N_8857,N_7873,N_7870);
nor U8858 (N_8858,N_7773,N_7729);
nor U8859 (N_8859,N_7200,N_7309);
or U8860 (N_8860,N_7781,N_7707);
or U8861 (N_8861,N_7982,N_7016);
nor U8862 (N_8862,N_7549,N_7663);
nand U8863 (N_8863,N_7155,N_7367);
and U8864 (N_8864,N_7043,N_7641);
and U8865 (N_8865,N_7036,N_7652);
or U8866 (N_8866,N_7133,N_7562);
nor U8867 (N_8867,N_7095,N_7387);
xor U8868 (N_8868,N_7680,N_7333);
and U8869 (N_8869,N_7368,N_7016);
nor U8870 (N_8870,N_7798,N_7754);
or U8871 (N_8871,N_7240,N_7379);
nor U8872 (N_8872,N_7700,N_7872);
nand U8873 (N_8873,N_7973,N_7265);
nand U8874 (N_8874,N_7069,N_7307);
and U8875 (N_8875,N_7195,N_7411);
and U8876 (N_8876,N_7405,N_7091);
or U8877 (N_8877,N_7618,N_7885);
and U8878 (N_8878,N_7954,N_7036);
nand U8879 (N_8879,N_7016,N_7839);
nor U8880 (N_8880,N_7452,N_7487);
nor U8881 (N_8881,N_7934,N_7561);
nand U8882 (N_8882,N_7037,N_7212);
xor U8883 (N_8883,N_7901,N_7559);
or U8884 (N_8884,N_7562,N_7649);
or U8885 (N_8885,N_7042,N_7572);
nor U8886 (N_8886,N_7765,N_7450);
xnor U8887 (N_8887,N_7436,N_7784);
nor U8888 (N_8888,N_7057,N_7972);
and U8889 (N_8889,N_7181,N_7408);
or U8890 (N_8890,N_7636,N_7113);
nand U8891 (N_8891,N_7929,N_7725);
nor U8892 (N_8892,N_7715,N_7827);
xnor U8893 (N_8893,N_7626,N_7227);
or U8894 (N_8894,N_7339,N_7049);
or U8895 (N_8895,N_7446,N_7979);
nand U8896 (N_8896,N_7220,N_7148);
and U8897 (N_8897,N_7825,N_7989);
nand U8898 (N_8898,N_7680,N_7628);
and U8899 (N_8899,N_7579,N_7892);
nand U8900 (N_8900,N_7332,N_7149);
or U8901 (N_8901,N_7747,N_7127);
xor U8902 (N_8902,N_7808,N_7774);
and U8903 (N_8903,N_7839,N_7171);
xnor U8904 (N_8904,N_7571,N_7606);
nor U8905 (N_8905,N_7213,N_7344);
xor U8906 (N_8906,N_7309,N_7809);
or U8907 (N_8907,N_7905,N_7108);
nand U8908 (N_8908,N_7234,N_7568);
nor U8909 (N_8909,N_7507,N_7246);
xor U8910 (N_8910,N_7566,N_7261);
and U8911 (N_8911,N_7219,N_7545);
xor U8912 (N_8912,N_7395,N_7774);
and U8913 (N_8913,N_7895,N_7788);
and U8914 (N_8914,N_7678,N_7042);
and U8915 (N_8915,N_7848,N_7866);
nand U8916 (N_8916,N_7446,N_7175);
or U8917 (N_8917,N_7354,N_7211);
nand U8918 (N_8918,N_7671,N_7263);
and U8919 (N_8919,N_7785,N_7557);
nand U8920 (N_8920,N_7370,N_7114);
or U8921 (N_8921,N_7510,N_7528);
nand U8922 (N_8922,N_7814,N_7734);
nand U8923 (N_8923,N_7844,N_7052);
and U8924 (N_8924,N_7644,N_7285);
nand U8925 (N_8925,N_7327,N_7272);
nand U8926 (N_8926,N_7385,N_7522);
or U8927 (N_8927,N_7541,N_7727);
nand U8928 (N_8928,N_7157,N_7016);
and U8929 (N_8929,N_7114,N_7290);
nor U8930 (N_8930,N_7703,N_7531);
or U8931 (N_8931,N_7099,N_7577);
nand U8932 (N_8932,N_7378,N_7692);
xnor U8933 (N_8933,N_7355,N_7542);
nand U8934 (N_8934,N_7623,N_7535);
xnor U8935 (N_8935,N_7678,N_7787);
nor U8936 (N_8936,N_7025,N_7125);
or U8937 (N_8937,N_7567,N_7022);
nand U8938 (N_8938,N_7728,N_7462);
nor U8939 (N_8939,N_7712,N_7131);
nor U8940 (N_8940,N_7033,N_7438);
nor U8941 (N_8941,N_7911,N_7928);
and U8942 (N_8942,N_7708,N_7776);
xor U8943 (N_8943,N_7923,N_7273);
nand U8944 (N_8944,N_7004,N_7795);
nand U8945 (N_8945,N_7415,N_7034);
and U8946 (N_8946,N_7780,N_7759);
nor U8947 (N_8947,N_7261,N_7750);
nand U8948 (N_8948,N_7710,N_7277);
nand U8949 (N_8949,N_7868,N_7428);
nor U8950 (N_8950,N_7666,N_7845);
and U8951 (N_8951,N_7394,N_7408);
and U8952 (N_8952,N_7806,N_7049);
or U8953 (N_8953,N_7492,N_7020);
nand U8954 (N_8954,N_7089,N_7858);
xnor U8955 (N_8955,N_7257,N_7547);
xnor U8956 (N_8956,N_7040,N_7046);
and U8957 (N_8957,N_7014,N_7529);
and U8958 (N_8958,N_7469,N_7568);
nand U8959 (N_8959,N_7603,N_7057);
nor U8960 (N_8960,N_7373,N_7123);
xnor U8961 (N_8961,N_7215,N_7652);
nor U8962 (N_8962,N_7406,N_7597);
and U8963 (N_8963,N_7355,N_7789);
xor U8964 (N_8964,N_7050,N_7656);
nand U8965 (N_8965,N_7658,N_7120);
xnor U8966 (N_8966,N_7605,N_7991);
xor U8967 (N_8967,N_7978,N_7329);
or U8968 (N_8968,N_7149,N_7763);
or U8969 (N_8969,N_7014,N_7361);
nand U8970 (N_8970,N_7201,N_7612);
and U8971 (N_8971,N_7361,N_7848);
nor U8972 (N_8972,N_7192,N_7725);
and U8973 (N_8973,N_7768,N_7594);
xnor U8974 (N_8974,N_7434,N_7205);
nor U8975 (N_8975,N_7055,N_7108);
nand U8976 (N_8976,N_7178,N_7979);
and U8977 (N_8977,N_7856,N_7651);
nand U8978 (N_8978,N_7986,N_7888);
nand U8979 (N_8979,N_7002,N_7866);
nor U8980 (N_8980,N_7767,N_7545);
or U8981 (N_8981,N_7882,N_7982);
or U8982 (N_8982,N_7342,N_7461);
nor U8983 (N_8983,N_7319,N_7593);
or U8984 (N_8984,N_7015,N_7448);
nor U8985 (N_8985,N_7834,N_7390);
nor U8986 (N_8986,N_7609,N_7784);
nand U8987 (N_8987,N_7571,N_7796);
nand U8988 (N_8988,N_7438,N_7554);
and U8989 (N_8989,N_7602,N_7064);
or U8990 (N_8990,N_7838,N_7519);
nor U8991 (N_8991,N_7290,N_7928);
and U8992 (N_8992,N_7789,N_7350);
xor U8993 (N_8993,N_7753,N_7772);
xnor U8994 (N_8994,N_7542,N_7387);
nand U8995 (N_8995,N_7555,N_7092);
xor U8996 (N_8996,N_7529,N_7719);
nor U8997 (N_8997,N_7173,N_7499);
nand U8998 (N_8998,N_7580,N_7697);
and U8999 (N_8999,N_7956,N_7477);
or U9000 (N_9000,N_8456,N_8241);
nor U9001 (N_9001,N_8266,N_8222);
and U9002 (N_9002,N_8818,N_8661);
nor U9003 (N_9003,N_8270,N_8153);
nor U9004 (N_9004,N_8023,N_8985);
or U9005 (N_9005,N_8007,N_8318);
and U9006 (N_9006,N_8202,N_8416);
nor U9007 (N_9007,N_8472,N_8931);
and U9008 (N_9008,N_8957,N_8120);
nand U9009 (N_9009,N_8684,N_8148);
nand U9010 (N_9010,N_8110,N_8555);
and U9011 (N_9011,N_8531,N_8519);
and U9012 (N_9012,N_8838,N_8198);
and U9013 (N_9013,N_8921,N_8160);
or U9014 (N_9014,N_8207,N_8847);
and U9015 (N_9015,N_8724,N_8221);
nand U9016 (N_9016,N_8060,N_8471);
and U9017 (N_9017,N_8587,N_8974);
nand U9018 (N_9018,N_8473,N_8329);
nand U9019 (N_9019,N_8161,N_8457);
or U9020 (N_9020,N_8451,N_8956);
or U9021 (N_9021,N_8116,N_8622);
and U9022 (N_9022,N_8552,N_8828);
nand U9023 (N_9023,N_8439,N_8501);
and U9024 (N_9024,N_8182,N_8085);
and U9025 (N_9025,N_8577,N_8333);
nand U9026 (N_9026,N_8192,N_8480);
and U9027 (N_9027,N_8417,N_8132);
and U9028 (N_9028,N_8083,N_8466);
nand U9029 (N_9029,N_8789,N_8246);
xor U9030 (N_9030,N_8903,N_8156);
nor U9031 (N_9031,N_8721,N_8759);
nand U9032 (N_9032,N_8984,N_8168);
xor U9033 (N_9033,N_8337,N_8402);
nor U9034 (N_9034,N_8176,N_8961);
xor U9035 (N_9035,N_8093,N_8028);
nor U9036 (N_9036,N_8239,N_8939);
nor U9037 (N_9037,N_8302,N_8374);
or U9038 (N_9038,N_8748,N_8338);
and U9039 (N_9039,N_8716,N_8010);
nand U9040 (N_9040,N_8389,N_8428);
and U9041 (N_9041,N_8145,N_8042);
and U9042 (N_9042,N_8217,N_8522);
or U9043 (N_9043,N_8282,N_8248);
or U9044 (N_9044,N_8876,N_8867);
or U9045 (N_9045,N_8654,N_8163);
nand U9046 (N_9046,N_8914,N_8667);
and U9047 (N_9047,N_8226,N_8504);
xnor U9048 (N_9048,N_8840,N_8879);
nand U9049 (N_9049,N_8484,N_8181);
nor U9050 (N_9050,N_8170,N_8560);
and U9051 (N_9051,N_8663,N_8362);
and U9052 (N_9052,N_8200,N_8923);
xor U9053 (N_9053,N_8762,N_8741);
nand U9054 (N_9054,N_8218,N_8870);
xor U9055 (N_9055,N_8404,N_8185);
and U9056 (N_9056,N_8334,N_8765);
nand U9057 (N_9057,N_8286,N_8004);
nand U9058 (N_9058,N_8698,N_8506);
xnor U9059 (N_9059,N_8056,N_8420);
nor U9060 (N_9060,N_8029,N_8799);
nand U9061 (N_9061,N_8082,N_8142);
nand U9062 (N_9062,N_8498,N_8041);
nor U9063 (N_9063,N_8073,N_8014);
nand U9064 (N_9064,N_8938,N_8067);
or U9065 (N_9065,N_8631,N_8433);
and U9066 (N_9066,N_8108,N_8670);
and U9067 (N_9067,N_8856,N_8650);
and U9068 (N_9068,N_8089,N_8959);
nor U9069 (N_9069,N_8419,N_8933);
and U9070 (N_9070,N_8469,N_8682);
xnor U9071 (N_9071,N_8016,N_8360);
or U9072 (N_9072,N_8758,N_8250);
or U9073 (N_9073,N_8874,N_8666);
nor U9074 (N_9074,N_8717,N_8753);
or U9075 (N_9075,N_8539,N_8008);
or U9076 (N_9076,N_8940,N_8962);
and U9077 (N_9077,N_8924,N_8851);
xnor U9078 (N_9078,N_8837,N_8925);
nand U9079 (N_9079,N_8367,N_8269);
nor U9080 (N_9080,N_8779,N_8688);
nor U9081 (N_9081,N_8964,N_8482);
nand U9082 (N_9082,N_8517,N_8460);
or U9083 (N_9083,N_8604,N_8893);
nand U9084 (N_9084,N_8236,N_8836);
nand U9085 (N_9085,N_8092,N_8548);
or U9086 (N_9086,N_8628,N_8109);
nor U9087 (N_9087,N_8071,N_8995);
xor U9088 (N_9088,N_8958,N_8397);
xor U9089 (N_9089,N_8188,N_8065);
xor U9090 (N_9090,N_8880,N_8340);
nor U9091 (N_9091,N_8760,N_8474);
nor U9092 (N_9092,N_8502,N_8275);
nand U9093 (N_9093,N_8697,N_8079);
nor U9094 (N_9094,N_8393,N_8194);
xnor U9095 (N_9095,N_8590,N_8094);
nor U9096 (N_9096,N_8297,N_8518);
or U9097 (N_9097,N_8934,N_8048);
or U9098 (N_9098,N_8227,N_8570);
nand U9099 (N_9099,N_8904,N_8727);
and U9100 (N_9100,N_8898,N_8510);
nand U9101 (N_9101,N_8848,N_8154);
nor U9102 (N_9102,N_8115,N_8049);
and U9103 (N_9103,N_8003,N_8038);
nor U9104 (N_9104,N_8113,N_8339);
and U9105 (N_9105,N_8695,N_8277);
nand U9106 (N_9106,N_8965,N_8101);
nand U9107 (N_9107,N_8576,N_8033);
nand U9108 (N_9108,N_8950,N_8778);
xor U9109 (N_9109,N_8315,N_8750);
or U9110 (N_9110,N_8172,N_8827);
nor U9111 (N_9111,N_8189,N_8289);
xnor U9112 (N_9112,N_8969,N_8937);
nor U9113 (N_9113,N_8017,N_8791);
nor U9114 (N_9114,N_8512,N_8019);
or U9115 (N_9115,N_8771,N_8763);
nor U9116 (N_9116,N_8128,N_8565);
and U9117 (N_9117,N_8342,N_8784);
nor U9118 (N_9118,N_8767,N_8283);
and U9119 (N_9119,N_8866,N_8888);
xnor U9120 (N_9120,N_8465,N_8119);
and U9121 (N_9121,N_8230,N_8986);
xor U9122 (N_9122,N_8887,N_8310);
or U9123 (N_9123,N_8262,N_8728);
nand U9124 (N_9124,N_8359,N_8546);
nor U9125 (N_9125,N_8736,N_8523);
and U9126 (N_9126,N_8686,N_8414);
nor U9127 (N_9127,N_8975,N_8813);
nand U9128 (N_9128,N_8766,N_8634);
nor U9129 (N_9129,N_8782,N_8216);
or U9130 (N_9130,N_8449,N_8685);
nor U9131 (N_9131,N_8798,N_8701);
nor U9132 (N_9132,N_8910,N_8745);
nor U9133 (N_9133,N_8392,N_8316);
nand U9134 (N_9134,N_8309,N_8494);
or U9135 (N_9135,N_8882,N_8461);
nand U9136 (N_9136,N_8993,N_8279);
and U9137 (N_9137,N_8044,N_8353);
nand U9138 (N_9138,N_8488,N_8639);
nor U9139 (N_9139,N_8117,N_8186);
and U9140 (N_9140,N_8233,N_8369);
or U9141 (N_9141,N_8797,N_8356);
and U9142 (N_9142,N_8345,N_8107);
or U9143 (N_9143,N_8897,N_8139);
nand U9144 (N_9144,N_8579,N_8648);
or U9145 (N_9145,N_8875,N_8668);
nand U9146 (N_9146,N_8179,N_8994);
nor U9147 (N_9147,N_8258,N_8293);
or U9148 (N_9148,N_8377,N_8599);
nor U9149 (N_9149,N_8436,N_8061);
nor U9150 (N_9150,N_8647,N_8573);
nor U9151 (N_9151,N_8596,N_8803);
nand U9152 (N_9152,N_8845,N_8299);
nor U9153 (N_9153,N_8209,N_8410);
nand U9154 (N_9154,N_8497,N_8388);
and U9155 (N_9155,N_8746,N_8043);
or U9156 (N_9156,N_8706,N_8646);
and U9157 (N_9157,N_8303,N_8676);
xnor U9158 (N_9158,N_8140,N_8951);
or U9159 (N_9159,N_8991,N_8920);
nor U9160 (N_9160,N_8588,N_8863);
xnor U9161 (N_9161,N_8589,N_8507);
nand U9162 (N_9162,N_8199,N_8922);
or U9163 (N_9163,N_8908,N_8544);
or U9164 (N_9164,N_8205,N_8575);
xor U9165 (N_9165,N_8725,N_8260);
xnor U9166 (N_9166,N_8878,N_8540);
nand U9167 (N_9167,N_8702,N_8580);
and U9168 (N_9168,N_8642,N_8752);
nor U9169 (N_9169,N_8086,N_8679);
nand U9170 (N_9170,N_8820,N_8455);
nand U9171 (N_9171,N_8850,N_8475);
nand U9172 (N_9172,N_8602,N_8247);
xor U9173 (N_9173,N_8889,N_8059);
nor U9174 (N_9174,N_8772,N_8280);
and U9175 (N_9175,N_8672,N_8208);
and U9176 (N_9176,N_8582,N_8683);
nor U9177 (N_9177,N_8581,N_8643);
xor U9178 (N_9178,N_8967,N_8124);
or U9179 (N_9179,N_8627,N_8183);
nor U9180 (N_9180,N_8326,N_8332);
nor U9181 (N_9181,N_8268,N_8164);
and U9182 (N_9182,N_8385,N_8087);
or U9183 (N_9183,N_8430,N_8865);
nand U9184 (N_9184,N_8399,N_8853);
nor U9185 (N_9185,N_8788,N_8902);
xor U9186 (N_9186,N_8568,N_8615);
or U9187 (N_9187,N_8499,N_8786);
nor U9188 (N_9188,N_8320,N_8660);
or U9189 (N_9189,N_8372,N_8992);
and U9190 (N_9190,N_8256,N_8877);
nand U9191 (N_9191,N_8632,N_8585);
nor U9192 (N_9192,N_8295,N_8006);
and U9193 (N_9193,N_8562,N_8013);
nor U9194 (N_9194,N_8158,N_8122);
nor U9195 (N_9195,N_8452,N_8141);
nand U9196 (N_9196,N_8406,N_8737);
nand U9197 (N_9197,N_8550,N_8689);
or U9198 (N_9198,N_8960,N_8123);
and U9199 (N_9199,N_8816,N_8125);
xnor U9200 (N_9200,N_8046,N_8220);
and U9201 (N_9201,N_8438,N_8595);
nand U9202 (N_9202,N_8052,N_8988);
or U9203 (N_9203,N_8096,N_8613);
or U9204 (N_9204,N_8755,N_8396);
nand U9205 (N_9205,N_8244,N_8138);
xor U9206 (N_9206,N_8435,N_8674);
nand U9207 (N_9207,N_8535,N_8321);
nand U9208 (N_9208,N_8864,N_8722);
nand U9209 (N_9209,N_8257,N_8794);
nand U9210 (N_9210,N_8411,N_8121);
nand U9211 (N_9211,N_8401,N_8169);
or U9212 (N_9212,N_8729,N_8476);
xnor U9213 (N_9213,N_8942,N_8407);
or U9214 (N_9214,N_8743,N_8335);
nand U9215 (N_9215,N_8653,N_8486);
nor U9216 (N_9216,N_8932,N_8658);
or U9217 (N_9217,N_8155,N_8478);
nand U9218 (N_9218,N_8190,N_8586);
and U9219 (N_9219,N_8989,N_8883);
nand U9220 (N_9220,N_8445,N_8718);
nand U9221 (N_9221,N_8711,N_8584);
or U9222 (N_9222,N_8001,N_8618);
nor U9223 (N_9223,N_8796,N_8814);
nor U9224 (N_9224,N_8928,N_8561);
nand U9225 (N_9225,N_8600,N_8536);
nand U9226 (N_9226,N_8290,N_8780);
nor U9227 (N_9227,N_8030,N_8285);
or U9228 (N_9228,N_8609,N_8998);
nand U9229 (N_9229,N_8913,N_8841);
nand U9230 (N_9230,N_8355,N_8051);
nand U9231 (N_9231,N_8231,N_8212);
or U9232 (N_9232,N_8640,N_8930);
nor U9233 (N_9233,N_8025,N_8503);
nand U9234 (N_9234,N_8180,N_8637);
or U9235 (N_9235,N_8129,N_8949);
and U9236 (N_9236,N_8662,N_8294);
nand U9237 (N_9237,N_8306,N_8551);
xor U9238 (N_9238,N_8623,N_8206);
nand U9239 (N_9239,N_8413,N_8458);
nor U9240 (N_9240,N_8687,N_8483);
nand U9241 (N_9241,N_8621,N_8846);
nand U9242 (N_9242,N_8700,N_8542);
nand U9243 (N_9243,N_8532,N_8253);
or U9244 (N_9244,N_8733,N_8177);
nand U9245 (N_9245,N_8699,N_8464);
nand U9246 (N_9246,N_8204,N_8804);
or U9247 (N_9247,N_8418,N_8441);
nand U9248 (N_9248,N_8907,N_8592);
and U9249 (N_9249,N_8768,N_8792);
nand U9250 (N_9250,N_8130,N_8605);
and U9251 (N_9251,N_8971,N_8809);
or U9252 (N_9252,N_8431,N_8022);
and U9253 (N_9253,N_8157,N_8376);
nor U9254 (N_9254,N_8754,N_8395);
nor U9255 (N_9255,N_8261,N_8284);
nand U9256 (N_9256,N_8553,N_8739);
or U9257 (N_9257,N_8424,N_8228);
and U9258 (N_9258,N_8031,N_8968);
or U9259 (N_9259,N_8629,N_8298);
xor U9260 (N_9260,N_8505,N_8616);
or U9261 (N_9261,N_8134,N_8611);
or U9262 (N_9262,N_8747,N_8823);
or U9263 (N_9263,N_8649,N_8514);
or U9264 (N_9264,N_8980,N_8574);
nand U9265 (N_9265,N_8375,N_8098);
nand U9266 (N_9266,N_8520,N_8673);
nor U9267 (N_9267,N_8015,N_8425);
nor U9268 (N_9268,N_8533,N_8868);
and U9269 (N_9269,N_8147,N_8541);
and U9270 (N_9270,N_8636,N_8343);
or U9271 (N_9271,N_8076,N_8184);
xnor U9272 (N_9272,N_8825,N_8774);
nand U9273 (N_9273,N_8608,N_8528);
nor U9274 (N_9274,N_8513,N_8901);
and U9275 (N_9275,N_8324,N_8749);
xnor U9276 (N_9276,N_8254,N_8097);
and U9277 (N_9277,N_8252,N_8511);
and U9278 (N_9278,N_8669,N_8919);
or U9279 (N_9279,N_8111,N_8665);
and U9280 (N_9280,N_8652,N_8869);
nor U9281 (N_9281,N_8074,N_8987);
or U9282 (N_9282,N_8873,N_8091);
and U9283 (N_9283,N_8734,N_8485);
nor U9284 (N_9284,N_8776,N_8273);
nor U9285 (N_9285,N_8970,N_8444);
or U9286 (N_9286,N_8890,N_8516);
xor U9287 (N_9287,N_8296,N_8826);
nor U9288 (N_9288,N_8619,N_8287);
nand U9289 (N_9289,N_8265,N_8659);
nand U9290 (N_9290,N_8103,N_8459);
or U9291 (N_9291,N_8214,N_8744);
xor U9292 (N_9292,N_8149,N_8319);
nand U9293 (N_9293,N_8211,N_8235);
and U9294 (N_9294,N_8999,N_8807);
or U9295 (N_9295,N_8322,N_8291);
and U9296 (N_9296,N_8821,N_8187);
or U9297 (N_9297,N_8106,N_8645);
nand U9298 (N_9298,N_8055,N_8681);
or U9299 (N_9299,N_8824,N_8620);
xnor U9300 (N_9300,N_8812,N_8549);
nor U9301 (N_9301,N_8862,N_8426);
nand U9302 (N_9302,N_8713,N_8527);
nand U9303 (N_9303,N_8166,N_8943);
nand U9304 (N_9304,N_8446,N_8379);
xnor U9305 (N_9305,N_8331,N_8104);
nor U9306 (N_9306,N_8657,N_8948);
and U9307 (N_9307,N_8423,N_8210);
nand U9308 (N_9308,N_8735,N_8447);
or U9309 (N_9309,N_8229,N_8412);
nor U9310 (N_9310,N_8378,N_8020);
or U9311 (N_9311,N_8150,N_8448);
nor U9312 (N_9312,N_8770,N_8521);
and U9313 (N_9313,N_8656,N_8223);
and U9314 (N_9314,N_8740,N_8597);
and U9315 (N_9315,N_8126,N_8834);
nand U9316 (N_9316,N_8308,N_8363);
or U9317 (N_9317,N_8144,N_8136);
or U9318 (N_9318,N_8035,N_8278);
nor U9319 (N_9319,N_8057,N_8045);
xnor U9320 (N_9320,N_8387,N_8034);
and U9321 (N_9321,N_8714,N_8349);
or U9322 (N_9322,N_8066,N_8365);
xor U9323 (N_9323,N_8978,N_8313);
nand U9324 (N_9324,N_8040,N_8380);
and U9325 (N_9325,N_8373,N_8274);
nand U9326 (N_9326,N_8479,N_8572);
nor U9327 (N_9327,N_8556,N_8311);
nand U9328 (N_9328,N_8099,N_8614);
nand U9329 (N_9329,N_8197,N_8583);
or U9330 (N_9330,N_8612,N_8899);
and U9331 (N_9331,N_8243,N_8972);
and U9332 (N_9332,N_8368,N_8219);
nand U9333 (N_9333,N_8351,N_8203);
and U9334 (N_9334,N_8830,N_8167);
nor U9335 (N_9335,N_8708,N_8276);
nor U9336 (N_9336,N_8490,N_8347);
or U9337 (N_9337,N_8358,N_8118);
nand U9338 (N_9338,N_8977,N_8131);
nor U9339 (N_9339,N_8403,N_8976);
xor U9340 (N_9340,N_8346,N_8525);
nand U9341 (N_9341,N_8617,N_8053);
nand U9342 (N_9342,N_8644,N_8357);
xor U9343 (N_9343,N_8601,N_8801);
nor U9344 (N_9344,N_8947,N_8861);
nand U9345 (N_9345,N_8281,N_8300);
nor U9346 (N_9346,N_8245,N_8677);
nor U9347 (N_9347,N_8945,N_8839);
nor U9348 (N_9348,N_8983,N_8526);
nand U9349 (N_9349,N_8707,N_8751);
and U9350 (N_9350,N_8894,N_8064);
and U9351 (N_9351,N_8193,N_8072);
xnor U9352 (N_9352,N_8468,N_8831);
xnor U9353 (N_9353,N_8723,N_8543);
nand U9354 (N_9354,N_8641,N_8292);
nor U9355 (N_9355,N_8781,N_8886);
and U9356 (N_9356,N_8162,N_8386);
nand U9357 (N_9357,N_8063,N_8655);
nor U9358 (N_9358,N_8234,N_8058);
nor U9359 (N_9359,N_8070,N_8390);
nand U9360 (N_9360,N_8691,N_8050);
nand U9361 (N_9361,N_8165,N_8026);
and U9362 (N_9362,N_8196,N_8593);
nor U9363 (N_9363,N_8911,N_8090);
nand U9364 (N_9364,N_8328,N_8912);
or U9365 (N_9365,N_8371,N_8624);
nor U9366 (N_9366,N_8844,N_8981);
and U9367 (N_9367,N_8429,N_8381);
and U9368 (N_9368,N_8761,N_8421);
nand U9369 (N_9369,N_8069,N_8731);
and U9370 (N_9370,N_8537,N_8178);
or U9371 (N_9371,N_8493,N_8470);
or U9372 (N_9372,N_8800,N_8238);
or U9373 (N_9373,N_8327,N_8712);
nor U9374 (N_9374,N_8871,N_8341);
or U9375 (N_9375,N_8591,N_8915);
and U9376 (N_9376,N_8929,N_8242);
and U9377 (N_9377,N_8935,N_8500);
or U9378 (N_9378,N_8489,N_8720);
and U9379 (N_9379,N_8849,N_8810);
and U9380 (N_9380,N_8884,N_8626);
or U9381 (N_9381,N_8635,N_8726);
nor U9382 (N_9382,N_8775,N_8255);
or U9383 (N_9383,N_8078,N_8080);
and U9384 (N_9384,N_8213,N_8545);
and U9385 (N_9385,N_8440,N_8633);
nor U9386 (N_9386,N_8941,N_8927);
and U9387 (N_9387,N_8529,N_8307);
nand U9388 (N_9388,N_8742,N_8664);
nand U9389 (N_9389,N_8515,N_8829);
nand U9390 (N_9390,N_8557,N_8408);
xor U9391 (N_9391,N_8606,N_8009);
nor U9392 (N_9392,N_8370,N_8240);
and U9393 (N_9393,N_8764,N_8530);
nor U9394 (N_9394,N_8492,N_8769);
nand U9395 (N_9395,N_8793,N_8415);
nand U9396 (N_9396,N_8963,N_8084);
or U9397 (N_9397,N_8088,N_8361);
nand U9398 (N_9398,N_8996,N_8625);
and U9399 (N_9399,N_8690,N_8437);
or U9400 (N_9400,N_8566,N_8855);
nand U9401 (N_9401,N_8481,N_8578);
xnor U9402 (N_9402,N_8487,N_8534);
nor U9403 (N_9403,N_8264,N_8610);
nand U9404 (N_9404,N_8990,N_8000);
nor U9405 (N_9405,N_8671,N_8719);
xor U9406 (N_9406,N_8391,N_8558);
and U9407 (N_9407,N_8382,N_8005);
and U9408 (N_9408,N_8594,N_8100);
xnor U9409 (N_9409,N_8559,N_8495);
nand U9410 (N_9410,N_8738,N_8892);
and U9411 (N_9411,N_8095,N_8305);
and U9412 (N_9412,N_8806,N_8811);
nor U9413 (N_9413,N_8018,N_8271);
nor U9414 (N_9414,N_8491,N_8508);
nand U9415 (N_9415,N_8710,N_8857);
nand U9416 (N_9416,N_8409,N_8224);
nand U9417 (N_9417,N_8304,N_8068);
or U9418 (N_9418,N_8895,N_8979);
and U9419 (N_9419,N_8678,N_8705);
and U9420 (N_9420,N_8703,N_8146);
nor U9421 (N_9421,N_8819,N_8603);
nor U9422 (N_9422,N_8953,N_8936);
or U9423 (N_9423,N_8330,N_8062);
xnor U9424 (N_9424,N_8692,N_8900);
nand U9425 (N_9425,N_8790,N_8102);
or U9426 (N_9426,N_8288,N_8012);
nor U9427 (N_9427,N_8715,N_8075);
and U9428 (N_9428,N_8171,N_8916);
nor U9429 (N_9429,N_8127,N_8997);
nor U9430 (N_9430,N_8027,N_8795);
and U9431 (N_9431,N_8442,N_8047);
or U9432 (N_9432,N_8785,N_8251);
and U9433 (N_9433,N_8191,N_8860);
and U9434 (N_9434,N_8133,N_8854);
nand U9435 (N_9435,N_8694,N_8024);
or U9436 (N_9436,N_8201,N_8822);
xnor U9437 (N_9437,N_8450,N_8114);
nand U9438 (N_9438,N_8434,N_8852);
nand U9439 (N_9439,N_8859,N_8817);
and U9440 (N_9440,N_8272,N_8159);
nor U9441 (N_9441,N_8077,N_8301);
and U9442 (N_9442,N_8354,N_8263);
or U9443 (N_9443,N_8783,N_8384);
nor U9444 (N_9444,N_8554,N_8454);
nor U9445 (N_9445,N_8215,N_8477);
or U9446 (N_9446,N_8757,N_8344);
and U9447 (N_9447,N_8105,N_8598);
xor U9448 (N_9448,N_8756,N_8680);
and U9449 (N_9449,N_8805,N_8952);
nand U9450 (N_9450,N_8366,N_8039);
and U9451 (N_9451,N_8872,N_8467);
or U9452 (N_9452,N_8569,N_8842);
nand U9453 (N_9453,N_8267,N_8881);
nor U9454 (N_9454,N_8021,N_8773);
nor U9455 (N_9455,N_8259,N_8730);
nor U9456 (N_9456,N_8112,N_8607);
and U9457 (N_9457,N_8944,N_8808);
nand U9458 (N_9458,N_8400,N_8462);
nand U9459 (N_9459,N_8336,N_8917);
or U9460 (N_9460,N_8509,N_8463);
nor U9461 (N_9461,N_8966,N_8249);
or U9462 (N_9462,N_8563,N_8896);
and U9463 (N_9463,N_8524,N_8954);
nand U9464 (N_9464,N_8152,N_8906);
nor U9465 (N_9465,N_8054,N_8777);
nand U9466 (N_9466,N_8323,N_8815);
xor U9467 (N_9467,N_8630,N_8651);
or U9468 (N_9468,N_8443,N_8709);
nor U9469 (N_9469,N_8732,N_8453);
nand U9470 (N_9470,N_8002,N_8352);
or U9471 (N_9471,N_8232,N_8946);
and U9472 (N_9472,N_8858,N_8955);
nor U9473 (N_9473,N_8833,N_8137);
xnor U9474 (N_9474,N_8364,N_8918);
nand U9475 (N_9475,N_8432,N_8312);
or U9476 (N_9476,N_8394,N_8036);
and U9477 (N_9477,N_8174,N_8905);
nor U9478 (N_9478,N_8926,N_8225);
or U9479 (N_9479,N_8143,N_8696);
or U9480 (N_9480,N_8398,N_8151);
or U9481 (N_9481,N_8547,N_8422);
or U9482 (N_9482,N_8787,N_8675);
and U9483 (N_9483,N_8314,N_8496);
or U9484 (N_9484,N_8982,N_8317);
or U9485 (N_9485,N_8832,N_8885);
xor U9486 (N_9486,N_8383,N_8011);
and U9487 (N_9487,N_8032,N_8909);
nor U9488 (N_9488,N_8973,N_8081);
nand U9489 (N_9489,N_8348,N_8135);
and U9490 (N_9490,N_8173,N_8405);
or U9491 (N_9491,N_8564,N_8571);
or U9492 (N_9492,N_8891,N_8638);
and U9493 (N_9493,N_8427,N_8195);
and U9494 (N_9494,N_8567,N_8704);
and U9495 (N_9495,N_8538,N_8325);
nand U9496 (N_9496,N_8037,N_8802);
and U9497 (N_9497,N_8237,N_8175);
nand U9498 (N_9498,N_8350,N_8835);
or U9499 (N_9499,N_8693,N_8843);
nor U9500 (N_9500,N_8648,N_8511);
and U9501 (N_9501,N_8881,N_8989);
or U9502 (N_9502,N_8137,N_8012);
and U9503 (N_9503,N_8189,N_8863);
and U9504 (N_9504,N_8354,N_8835);
nand U9505 (N_9505,N_8905,N_8432);
or U9506 (N_9506,N_8908,N_8904);
and U9507 (N_9507,N_8660,N_8825);
and U9508 (N_9508,N_8540,N_8590);
nand U9509 (N_9509,N_8755,N_8495);
xor U9510 (N_9510,N_8166,N_8092);
nor U9511 (N_9511,N_8878,N_8697);
or U9512 (N_9512,N_8175,N_8289);
and U9513 (N_9513,N_8563,N_8137);
or U9514 (N_9514,N_8475,N_8571);
or U9515 (N_9515,N_8283,N_8709);
nor U9516 (N_9516,N_8624,N_8092);
nor U9517 (N_9517,N_8637,N_8380);
and U9518 (N_9518,N_8385,N_8277);
xor U9519 (N_9519,N_8014,N_8791);
or U9520 (N_9520,N_8158,N_8827);
and U9521 (N_9521,N_8074,N_8207);
nor U9522 (N_9522,N_8294,N_8793);
or U9523 (N_9523,N_8985,N_8872);
nand U9524 (N_9524,N_8962,N_8367);
nand U9525 (N_9525,N_8467,N_8903);
xor U9526 (N_9526,N_8478,N_8649);
nand U9527 (N_9527,N_8254,N_8441);
nor U9528 (N_9528,N_8595,N_8017);
nor U9529 (N_9529,N_8524,N_8899);
xnor U9530 (N_9530,N_8694,N_8781);
or U9531 (N_9531,N_8385,N_8144);
nand U9532 (N_9532,N_8101,N_8295);
nor U9533 (N_9533,N_8309,N_8774);
nand U9534 (N_9534,N_8244,N_8730);
nand U9535 (N_9535,N_8813,N_8849);
nor U9536 (N_9536,N_8667,N_8021);
nand U9537 (N_9537,N_8399,N_8468);
nand U9538 (N_9538,N_8480,N_8394);
nand U9539 (N_9539,N_8999,N_8100);
or U9540 (N_9540,N_8731,N_8498);
and U9541 (N_9541,N_8197,N_8976);
nand U9542 (N_9542,N_8599,N_8129);
or U9543 (N_9543,N_8334,N_8784);
nand U9544 (N_9544,N_8571,N_8349);
and U9545 (N_9545,N_8662,N_8532);
nand U9546 (N_9546,N_8607,N_8161);
or U9547 (N_9547,N_8562,N_8540);
and U9548 (N_9548,N_8528,N_8036);
nor U9549 (N_9549,N_8101,N_8978);
nand U9550 (N_9550,N_8538,N_8687);
and U9551 (N_9551,N_8699,N_8587);
and U9552 (N_9552,N_8355,N_8029);
nand U9553 (N_9553,N_8080,N_8858);
and U9554 (N_9554,N_8383,N_8734);
nand U9555 (N_9555,N_8705,N_8113);
nor U9556 (N_9556,N_8463,N_8564);
and U9557 (N_9557,N_8713,N_8235);
or U9558 (N_9558,N_8696,N_8473);
and U9559 (N_9559,N_8002,N_8877);
and U9560 (N_9560,N_8880,N_8821);
nand U9561 (N_9561,N_8750,N_8543);
nand U9562 (N_9562,N_8763,N_8624);
nor U9563 (N_9563,N_8010,N_8784);
nand U9564 (N_9564,N_8314,N_8272);
and U9565 (N_9565,N_8879,N_8550);
or U9566 (N_9566,N_8216,N_8747);
and U9567 (N_9567,N_8343,N_8205);
and U9568 (N_9568,N_8739,N_8789);
nand U9569 (N_9569,N_8756,N_8976);
nor U9570 (N_9570,N_8169,N_8479);
and U9571 (N_9571,N_8305,N_8350);
nor U9572 (N_9572,N_8114,N_8364);
nor U9573 (N_9573,N_8994,N_8082);
nor U9574 (N_9574,N_8931,N_8541);
and U9575 (N_9575,N_8564,N_8259);
nor U9576 (N_9576,N_8351,N_8070);
nor U9577 (N_9577,N_8469,N_8185);
or U9578 (N_9578,N_8501,N_8488);
nand U9579 (N_9579,N_8500,N_8411);
nand U9580 (N_9580,N_8412,N_8587);
nand U9581 (N_9581,N_8441,N_8857);
or U9582 (N_9582,N_8097,N_8444);
xnor U9583 (N_9583,N_8804,N_8781);
or U9584 (N_9584,N_8665,N_8870);
and U9585 (N_9585,N_8145,N_8305);
nor U9586 (N_9586,N_8980,N_8547);
xnor U9587 (N_9587,N_8109,N_8141);
nor U9588 (N_9588,N_8018,N_8454);
and U9589 (N_9589,N_8940,N_8550);
nand U9590 (N_9590,N_8966,N_8595);
and U9591 (N_9591,N_8059,N_8250);
xor U9592 (N_9592,N_8784,N_8386);
xnor U9593 (N_9593,N_8953,N_8915);
nor U9594 (N_9594,N_8339,N_8038);
nand U9595 (N_9595,N_8403,N_8887);
nand U9596 (N_9596,N_8538,N_8461);
nand U9597 (N_9597,N_8115,N_8319);
and U9598 (N_9598,N_8516,N_8186);
and U9599 (N_9599,N_8857,N_8999);
nor U9600 (N_9600,N_8667,N_8217);
nor U9601 (N_9601,N_8124,N_8376);
and U9602 (N_9602,N_8289,N_8883);
or U9603 (N_9603,N_8699,N_8691);
and U9604 (N_9604,N_8148,N_8812);
and U9605 (N_9605,N_8344,N_8202);
nor U9606 (N_9606,N_8448,N_8059);
and U9607 (N_9607,N_8800,N_8506);
nor U9608 (N_9608,N_8081,N_8980);
nor U9609 (N_9609,N_8715,N_8900);
or U9610 (N_9610,N_8831,N_8701);
nor U9611 (N_9611,N_8169,N_8322);
nand U9612 (N_9612,N_8527,N_8751);
nand U9613 (N_9613,N_8411,N_8785);
and U9614 (N_9614,N_8991,N_8178);
nor U9615 (N_9615,N_8070,N_8382);
xnor U9616 (N_9616,N_8341,N_8023);
and U9617 (N_9617,N_8579,N_8416);
nor U9618 (N_9618,N_8807,N_8432);
or U9619 (N_9619,N_8701,N_8316);
nand U9620 (N_9620,N_8354,N_8809);
and U9621 (N_9621,N_8052,N_8853);
nand U9622 (N_9622,N_8249,N_8525);
nor U9623 (N_9623,N_8326,N_8872);
nand U9624 (N_9624,N_8446,N_8332);
nor U9625 (N_9625,N_8131,N_8253);
nor U9626 (N_9626,N_8309,N_8156);
nand U9627 (N_9627,N_8939,N_8394);
xor U9628 (N_9628,N_8968,N_8873);
or U9629 (N_9629,N_8949,N_8476);
or U9630 (N_9630,N_8463,N_8702);
nor U9631 (N_9631,N_8415,N_8095);
and U9632 (N_9632,N_8271,N_8683);
and U9633 (N_9633,N_8549,N_8916);
nor U9634 (N_9634,N_8461,N_8584);
nand U9635 (N_9635,N_8972,N_8900);
and U9636 (N_9636,N_8018,N_8680);
and U9637 (N_9637,N_8048,N_8665);
or U9638 (N_9638,N_8133,N_8163);
or U9639 (N_9639,N_8063,N_8684);
and U9640 (N_9640,N_8215,N_8239);
nand U9641 (N_9641,N_8219,N_8090);
xor U9642 (N_9642,N_8415,N_8952);
and U9643 (N_9643,N_8705,N_8304);
or U9644 (N_9644,N_8660,N_8311);
or U9645 (N_9645,N_8915,N_8037);
nand U9646 (N_9646,N_8021,N_8307);
nand U9647 (N_9647,N_8889,N_8435);
nand U9648 (N_9648,N_8489,N_8240);
or U9649 (N_9649,N_8048,N_8515);
xnor U9650 (N_9650,N_8699,N_8237);
nor U9651 (N_9651,N_8891,N_8428);
nand U9652 (N_9652,N_8672,N_8852);
and U9653 (N_9653,N_8854,N_8192);
nor U9654 (N_9654,N_8141,N_8687);
or U9655 (N_9655,N_8047,N_8587);
nor U9656 (N_9656,N_8689,N_8029);
nor U9657 (N_9657,N_8658,N_8184);
nor U9658 (N_9658,N_8439,N_8378);
or U9659 (N_9659,N_8620,N_8583);
nor U9660 (N_9660,N_8937,N_8634);
nand U9661 (N_9661,N_8992,N_8565);
or U9662 (N_9662,N_8958,N_8086);
and U9663 (N_9663,N_8070,N_8544);
and U9664 (N_9664,N_8961,N_8734);
xnor U9665 (N_9665,N_8165,N_8819);
and U9666 (N_9666,N_8831,N_8398);
and U9667 (N_9667,N_8029,N_8513);
xnor U9668 (N_9668,N_8153,N_8129);
nor U9669 (N_9669,N_8608,N_8737);
nand U9670 (N_9670,N_8495,N_8680);
nand U9671 (N_9671,N_8099,N_8907);
nand U9672 (N_9672,N_8483,N_8748);
or U9673 (N_9673,N_8051,N_8126);
xor U9674 (N_9674,N_8991,N_8097);
and U9675 (N_9675,N_8759,N_8645);
nand U9676 (N_9676,N_8906,N_8163);
nor U9677 (N_9677,N_8392,N_8257);
and U9678 (N_9678,N_8856,N_8560);
and U9679 (N_9679,N_8104,N_8284);
and U9680 (N_9680,N_8221,N_8619);
nor U9681 (N_9681,N_8533,N_8728);
nand U9682 (N_9682,N_8351,N_8731);
or U9683 (N_9683,N_8526,N_8629);
nor U9684 (N_9684,N_8345,N_8556);
and U9685 (N_9685,N_8883,N_8642);
nor U9686 (N_9686,N_8189,N_8243);
nor U9687 (N_9687,N_8292,N_8564);
or U9688 (N_9688,N_8623,N_8187);
and U9689 (N_9689,N_8198,N_8591);
or U9690 (N_9690,N_8413,N_8563);
and U9691 (N_9691,N_8679,N_8702);
nor U9692 (N_9692,N_8299,N_8420);
and U9693 (N_9693,N_8234,N_8970);
nand U9694 (N_9694,N_8861,N_8506);
and U9695 (N_9695,N_8951,N_8190);
nand U9696 (N_9696,N_8335,N_8636);
nor U9697 (N_9697,N_8954,N_8758);
xor U9698 (N_9698,N_8221,N_8578);
or U9699 (N_9699,N_8492,N_8842);
or U9700 (N_9700,N_8101,N_8213);
or U9701 (N_9701,N_8465,N_8828);
nand U9702 (N_9702,N_8722,N_8760);
nand U9703 (N_9703,N_8017,N_8102);
nor U9704 (N_9704,N_8491,N_8385);
nor U9705 (N_9705,N_8928,N_8208);
xor U9706 (N_9706,N_8881,N_8394);
or U9707 (N_9707,N_8125,N_8595);
nand U9708 (N_9708,N_8618,N_8411);
or U9709 (N_9709,N_8013,N_8134);
nor U9710 (N_9710,N_8657,N_8128);
and U9711 (N_9711,N_8311,N_8449);
xor U9712 (N_9712,N_8632,N_8802);
nand U9713 (N_9713,N_8043,N_8090);
nand U9714 (N_9714,N_8725,N_8865);
nor U9715 (N_9715,N_8510,N_8579);
nand U9716 (N_9716,N_8363,N_8122);
nor U9717 (N_9717,N_8812,N_8911);
or U9718 (N_9718,N_8680,N_8291);
or U9719 (N_9719,N_8104,N_8600);
nand U9720 (N_9720,N_8332,N_8139);
nor U9721 (N_9721,N_8066,N_8172);
nand U9722 (N_9722,N_8494,N_8207);
nor U9723 (N_9723,N_8970,N_8827);
and U9724 (N_9724,N_8943,N_8875);
nand U9725 (N_9725,N_8761,N_8770);
or U9726 (N_9726,N_8482,N_8527);
nor U9727 (N_9727,N_8356,N_8258);
or U9728 (N_9728,N_8630,N_8890);
or U9729 (N_9729,N_8599,N_8402);
xnor U9730 (N_9730,N_8916,N_8091);
or U9731 (N_9731,N_8017,N_8925);
nand U9732 (N_9732,N_8614,N_8356);
or U9733 (N_9733,N_8784,N_8392);
nor U9734 (N_9734,N_8568,N_8985);
nand U9735 (N_9735,N_8695,N_8645);
or U9736 (N_9736,N_8298,N_8637);
or U9737 (N_9737,N_8574,N_8765);
xor U9738 (N_9738,N_8366,N_8601);
and U9739 (N_9739,N_8655,N_8283);
nand U9740 (N_9740,N_8502,N_8218);
nor U9741 (N_9741,N_8268,N_8197);
nor U9742 (N_9742,N_8719,N_8272);
nand U9743 (N_9743,N_8908,N_8676);
and U9744 (N_9744,N_8106,N_8284);
nand U9745 (N_9745,N_8644,N_8525);
and U9746 (N_9746,N_8561,N_8994);
or U9747 (N_9747,N_8940,N_8580);
xor U9748 (N_9748,N_8691,N_8654);
nand U9749 (N_9749,N_8152,N_8100);
or U9750 (N_9750,N_8878,N_8236);
xnor U9751 (N_9751,N_8611,N_8425);
nor U9752 (N_9752,N_8971,N_8392);
nand U9753 (N_9753,N_8532,N_8609);
xor U9754 (N_9754,N_8608,N_8809);
and U9755 (N_9755,N_8246,N_8396);
nor U9756 (N_9756,N_8882,N_8494);
nand U9757 (N_9757,N_8546,N_8381);
nor U9758 (N_9758,N_8558,N_8831);
xor U9759 (N_9759,N_8752,N_8277);
and U9760 (N_9760,N_8371,N_8351);
nand U9761 (N_9761,N_8677,N_8688);
nand U9762 (N_9762,N_8389,N_8357);
and U9763 (N_9763,N_8833,N_8679);
and U9764 (N_9764,N_8154,N_8714);
nor U9765 (N_9765,N_8938,N_8009);
nand U9766 (N_9766,N_8956,N_8290);
nand U9767 (N_9767,N_8755,N_8332);
nand U9768 (N_9768,N_8392,N_8124);
and U9769 (N_9769,N_8993,N_8049);
nand U9770 (N_9770,N_8370,N_8427);
nand U9771 (N_9771,N_8966,N_8524);
nand U9772 (N_9772,N_8018,N_8320);
and U9773 (N_9773,N_8167,N_8481);
xor U9774 (N_9774,N_8806,N_8867);
xnor U9775 (N_9775,N_8412,N_8915);
and U9776 (N_9776,N_8182,N_8240);
nand U9777 (N_9777,N_8660,N_8904);
and U9778 (N_9778,N_8823,N_8878);
nand U9779 (N_9779,N_8534,N_8547);
and U9780 (N_9780,N_8242,N_8786);
or U9781 (N_9781,N_8732,N_8949);
and U9782 (N_9782,N_8014,N_8521);
nand U9783 (N_9783,N_8578,N_8430);
or U9784 (N_9784,N_8938,N_8896);
nor U9785 (N_9785,N_8158,N_8176);
and U9786 (N_9786,N_8548,N_8387);
and U9787 (N_9787,N_8664,N_8708);
or U9788 (N_9788,N_8880,N_8206);
nand U9789 (N_9789,N_8806,N_8229);
or U9790 (N_9790,N_8487,N_8975);
nor U9791 (N_9791,N_8935,N_8735);
nand U9792 (N_9792,N_8346,N_8131);
nor U9793 (N_9793,N_8344,N_8103);
or U9794 (N_9794,N_8490,N_8298);
or U9795 (N_9795,N_8340,N_8806);
nand U9796 (N_9796,N_8669,N_8049);
or U9797 (N_9797,N_8789,N_8481);
nor U9798 (N_9798,N_8716,N_8126);
nand U9799 (N_9799,N_8243,N_8943);
xnor U9800 (N_9800,N_8253,N_8367);
nor U9801 (N_9801,N_8943,N_8803);
or U9802 (N_9802,N_8891,N_8701);
xor U9803 (N_9803,N_8290,N_8687);
or U9804 (N_9804,N_8025,N_8214);
or U9805 (N_9805,N_8833,N_8143);
xnor U9806 (N_9806,N_8148,N_8360);
and U9807 (N_9807,N_8900,N_8145);
and U9808 (N_9808,N_8831,N_8885);
or U9809 (N_9809,N_8886,N_8677);
nand U9810 (N_9810,N_8744,N_8481);
or U9811 (N_9811,N_8168,N_8076);
nand U9812 (N_9812,N_8995,N_8288);
nor U9813 (N_9813,N_8779,N_8152);
nor U9814 (N_9814,N_8491,N_8667);
and U9815 (N_9815,N_8515,N_8985);
or U9816 (N_9816,N_8516,N_8451);
or U9817 (N_9817,N_8206,N_8621);
and U9818 (N_9818,N_8471,N_8035);
or U9819 (N_9819,N_8870,N_8118);
or U9820 (N_9820,N_8310,N_8533);
and U9821 (N_9821,N_8664,N_8633);
nand U9822 (N_9822,N_8540,N_8970);
nor U9823 (N_9823,N_8746,N_8772);
nand U9824 (N_9824,N_8644,N_8307);
nand U9825 (N_9825,N_8758,N_8228);
or U9826 (N_9826,N_8285,N_8510);
nor U9827 (N_9827,N_8874,N_8636);
or U9828 (N_9828,N_8681,N_8040);
or U9829 (N_9829,N_8764,N_8396);
or U9830 (N_9830,N_8935,N_8523);
nand U9831 (N_9831,N_8080,N_8631);
or U9832 (N_9832,N_8662,N_8753);
nand U9833 (N_9833,N_8858,N_8193);
nor U9834 (N_9834,N_8755,N_8467);
nor U9835 (N_9835,N_8447,N_8339);
or U9836 (N_9836,N_8822,N_8943);
and U9837 (N_9837,N_8309,N_8238);
and U9838 (N_9838,N_8239,N_8722);
or U9839 (N_9839,N_8182,N_8261);
nor U9840 (N_9840,N_8863,N_8193);
xnor U9841 (N_9841,N_8705,N_8492);
and U9842 (N_9842,N_8714,N_8394);
nor U9843 (N_9843,N_8297,N_8755);
nand U9844 (N_9844,N_8368,N_8444);
nand U9845 (N_9845,N_8336,N_8868);
nor U9846 (N_9846,N_8604,N_8832);
nor U9847 (N_9847,N_8007,N_8204);
nand U9848 (N_9848,N_8417,N_8925);
nor U9849 (N_9849,N_8292,N_8783);
nand U9850 (N_9850,N_8011,N_8197);
and U9851 (N_9851,N_8378,N_8513);
nor U9852 (N_9852,N_8683,N_8728);
nand U9853 (N_9853,N_8310,N_8395);
and U9854 (N_9854,N_8521,N_8303);
xor U9855 (N_9855,N_8601,N_8668);
nand U9856 (N_9856,N_8041,N_8774);
nand U9857 (N_9857,N_8223,N_8130);
and U9858 (N_9858,N_8429,N_8140);
and U9859 (N_9859,N_8767,N_8305);
or U9860 (N_9860,N_8626,N_8086);
nor U9861 (N_9861,N_8254,N_8800);
nand U9862 (N_9862,N_8733,N_8631);
nor U9863 (N_9863,N_8064,N_8586);
nand U9864 (N_9864,N_8439,N_8655);
nor U9865 (N_9865,N_8940,N_8825);
nor U9866 (N_9866,N_8714,N_8133);
nand U9867 (N_9867,N_8344,N_8893);
nand U9868 (N_9868,N_8538,N_8915);
xor U9869 (N_9869,N_8937,N_8344);
nor U9870 (N_9870,N_8286,N_8308);
nand U9871 (N_9871,N_8970,N_8603);
nor U9872 (N_9872,N_8562,N_8857);
nand U9873 (N_9873,N_8576,N_8529);
nand U9874 (N_9874,N_8607,N_8351);
and U9875 (N_9875,N_8408,N_8240);
and U9876 (N_9876,N_8712,N_8991);
nand U9877 (N_9877,N_8801,N_8657);
and U9878 (N_9878,N_8157,N_8280);
and U9879 (N_9879,N_8599,N_8493);
and U9880 (N_9880,N_8375,N_8667);
and U9881 (N_9881,N_8215,N_8149);
or U9882 (N_9882,N_8247,N_8125);
or U9883 (N_9883,N_8863,N_8042);
or U9884 (N_9884,N_8345,N_8775);
xor U9885 (N_9885,N_8089,N_8719);
and U9886 (N_9886,N_8339,N_8350);
or U9887 (N_9887,N_8338,N_8278);
or U9888 (N_9888,N_8289,N_8231);
or U9889 (N_9889,N_8631,N_8144);
nand U9890 (N_9890,N_8077,N_8315);
or U9891 (N_9891,N_8048,N_8119);
and U9892 (N_9892,N_8168,N_8731);
or U9893 (N_9893,N_8378,N_8943);
nor U9894 (N_9894,N_8943,N_8630);
nor U9895 (N_9895,N_8225,N_8867);
and U9896 (N_9896,N_8303,N_8730);
nand U9897 (N_9897,N_8320,N_8063);
nand U9898 (N_9898,N_8011,N_8562);
or U9899 (N_9899,N_8039,N_8658);
nor U9900 (N_9900,N_8841,N_8828);
nor U9901 (N_9901,N_8383,N_8560);
nand U9902 (N_9902,N_8039,N_8483);
and U9903 (N_9903,N_8567,N_8763);
and U9904 (N_9904,N_8828,N_8360);
nand U9905 (N_9905,N_8211,N_8213);
or U9906 (N_9906,N_8593,N_8193);
nor U9907 (N_9907,N_8946,N_8123);
nor U9908 (N_9908,N_8736,N_8924);
nor U9909 (N_9909,N_8460,N_8135);
nand U9910 (N_9910,N_8702,N_8271);
nor U9911 (N_9911,N_8532,N_8255);
xor U9912 (N_9912,N_8441,N_8595);
nor U9913 (N_9913,N_8252,N_8990);
xor U9914 (N_9914,N_8547,N_8884);
nor U9915 (N_9915,N_8496,N_8980);
or U9916 (N_9916,N_8265,N_8111);
xnor U9917 (N_9917,N_8977,N_8589);
nor U9918 (N_9918,N_8853,N_8835);
xnor U9919 (N_9919,N_8481,N_8127);
nor U9920 (N_9920,N_8506,N_8765);
and U9921 (N_9921,N_8401,N_8192);
nor U9922 (N_9922,N_8641,N_8502);
nand U9923 (N_9923,N_8594,N_8816);
nand U9924 (N_9924,N_8636,N_8642);
nor U9925 (N_9925,N_8690,N_8858);
xnor U9926 (N_9926,N_8355,N_8554);
and U9927 (N_9927,N_8704,N_8062);
nand U9928 (N_9928,N_8783,N_8110);
nor U9929 (N_9929,N_8409,N_8370);
and U9930 (N_9930,N_8558,N_8501);
or U9931 (N_9931,N_8536,N_8285);
xor U9932 (N_9932,N_8829,N_8291);
nor U9933 (N_9933,N_8025,N_8768);
or U9934 (N_9934,N_8397,N_8926);
nor U9935 (N_9935,N_8729,N_8473);
or U9936 (N_9936,N_8530,N_8232);
or U9937 (N_9937,N_8796,N_8650);
nand U9938 (N_9938,N_8723,N_8002);
or U9939 (N_9939,N_8223,N_8371);
xor U9940 (N_9940,N_8523,N_8259);
and U9941 (N_9941,N_8825,N_8832);
or U9942 (N_9942,N_8870,N_8038);
nor U9943 (N_9943,N_8263,N_8131);
nand U9944 (N_9944,N_8596,N_8248);
xnor U9945 (N_9945,N_8587,N_8056);
and U9946 (N_9946,N_8519,N_8094);
or U9947 (N_9947,N_8153,N_8973);
nand U9948 (N_9948,N_8303,N_8335);
and U9949 (N_9949,N_8145,N_8858);
and U9950 (N_9950,N_8312,N_8723);
nand U9951 (N_9951,N_8721,N_8095);
or U9952 (N_9952,N_8263,N_8245);
and U9953 (N_9953,N_8102,N_8160);
or U9954 (N_9954,N_8252,N_8936);
nor U9955 (N_9955,N_8219,N_8751);
and U9956 (N_9956,N_8663,N_8523);
or U9957 (N_9957,N_8249,N_8654);
and U9958 (N_9958,N_8853,N_8765);
and U9959 (N_9959,N_8393,N_8774);
nor U9960 (N_9960,N_8438,N_8095);
and U9961 (N_9961,N_8403,N_8073);
nand U9962 (N_9962,N_8696,N_8303);
or U9963 (N_9963,N_8222,N_8662);
nand U9964 (N_9964,N_8500,N_8577);
xor U9965 (N_9965,N_8429,N_8157);
nand U9966 (N_9966,N_8630,N_8316);
and U9967 (N_9967,N_8884,N_8186);
and U9968 (N_9968,N_8602,N_8164);
nand U9969 (N_9969,N_8216,N_8245);
nor U9970 (N_9970,N_8918,N_8271);
nor U9971 (N_9971,N_8649,N_8523);
xnor U9972 (N_9972,N_8254,N_8572);
and U9973 (N_9973,N_8551,N_8443);
nand U9974 (N_9974,N_8175,N_8802);
or U9975 (N_9975,N_8367,N_8792);
and U9976 (N_9976,N_8390,N_8054);
and U9977 (N_9977,N_8704,N_8642);
nor U9978 (N_9978,N_8245,N_8342);
or U9979 (N_9979,N_8689,N_8221);
and U9980 (N_9980,N_8446,N_8427);
and U9981 (N_9981,N_8307,N_8811);
or U9982 (N_9982,N_8593,N_8891);
and U9983 (N_9983,N_8257,N_8474);
and U9984 (N_9984,N_8062,N_8655);
or U9985 (N_9985,N_8671,N_8303);
xnor U9986 (N_9986,N_8321,N_8744);
xor U9987 (N_9987,N_8458,N_8610);
and U9988 (N_9988,N_8571,N_8297);
nand U9989 (N_9989,N_8138,N_8029);
and U9990 (N_9990,N_8381,N_8600);
and U9991 (N_9991,N_8361,N_8405);
nand U9992 (N_9992,N_8284,N_8443);
xnor U9993 (N_9993,N_8482,N_8499);
nand U9994 (N_9994,N_8749,N_8933);
nor U9995 (N_9995,N_8835,N_8870);
nor U9996 (N_9996,N_8189,N_8520);
nand U9997 (N_9997,N_8214,N_8885);
or U9998 (N_9998,N_8471,N_8798);
and U9999 (N_9999,N_8473,N_8866);
nor U10000 (N_10000,N_9091,N_9622);
nand U10001 (N_10001,N_9853,N_9394);
nand U10002 (N_10002,N_9023,N_9199);
and U10003 (N_10003,N_9710,N_9180);
and U10004 (N_10004,N_9335,N_9107);
xnor U10005 (N_10005,N_9385,N_9550);
nand U10006 (N_10006,N_9342,N_9676);
xor U10007 (N_10007,N_9787,N_9174);
xnor U10008 (N_10008,N_9034,N_9879);
or U10009 (N_10009,N_9408,N_9451);
or U10010 (N_10010,N_9522,N_9055);
xor U10011 (N_10011,N_9286,N_9650);
and U10012 (N_10012,N_9299,N_9063);
xor U10013 (N_10013,N_9968,N_9581);
nor U10014 (N_10014,N_9726,N_9017);
or U10015 (N_10015,N_9035,N_9521);
nor U10016 (N_10016,N_9626,N_9586);
nand U10017 (N_10017,N_9992,N_9907);
and U10018 (N_10018,N_9250,N_9821);
or U10019 (N_10019,N_9936,N_9670);
or U10020 (N_10020,N_9865,N_9925);
nor U10021 (N_10021,N_9002,N_9763);
and U10022 (N_10022,N_9155,N_9212);
and U10023 (N_10023,N_9858,N_9437);
and U10024 (N_10024,N_9652,N_9556);
nand U10025 (N_10025,N_9530,N_9987);
nand U10026 (N_10026,N_9053,N_9756);
nand U10027 (N_10027,N_9897,N_9507);
nand U10028 (N_10028,N_9672,N_9344);
and U10029 (N_10029,N_9528,N_9237);
or U10030 (N_10030,N_9085,N_9825);
or U10031 (N_10031,N_9628,N_9599);
or U10032 (N_10032,N_9057,N_9312);
and U10033 (N_10033,N_9568,N_9957);
nor U10034 (N_10034,N_9014,N_9928);
and U10035 (N_10035,N_9187,N_9078);
and U10036 (N_10036,N_9460,N_9724);
and U10037 (N_10037,N_9478,N_9240);
or U10038 (N_10038,N_9243,N_9043);
nor U10039 (N_10039,N_9164,N_9177);
xor U10040 (N_10040,N_9816,N_9012);
and U10041 (N_10041,N_9480,N_9494);
nor U10042 (N_10042,N_9734,N_9130);
or U10043 (N_10043,N_9304,N_9148);
nand U10044 (N_10044,N_9838,N_9236);
or U10045 (N_10045,N_9254,N_9784);
and U10046 (N_10046,N_9452,N_9347);
nor U10047 (N_10047,N_9366,N_9737);
nor U10048 (N_10048,N_9955,N_9808);
nand U10049 (N_10049,N_9436,N_9569);
nand U10050 (N_10050,N_9706,N_9317);
or U10051 (N_10051,N_9336,N_9118);
nand U10052 (N_10052,N_9602,N_9917);
or U10053 (N_10053,N_9306,N_9506);
xor U10054 (N_10054,N_9900,N_9213);
and U10055 (N_10055,N_9662,N_9776);
nor U10056 (N_10056,N_9643,N_9051);
nand U10057 (N_10057,N_9360,N_9358);
or U10058 (N_10058,N_9890,N_9584);
and U10059 (N_10059,N_9944,N_9223);
nor U10060 (N_10060,N_9577,N_9631);
nor U10061 (N_10061,N_9975,N_9022);
nand U10062 (N_10062,N_9515,N_9860);
and U10063 (N_10063,N_9627,N_9463);
and U10064 (N_10064,N_9050,N_9178);
nor U10065 (N_10065,N_9100,N_9849);
nand U10066 (N_10066,N_9161,N_9994);
nand U10067 (N_10067,N_9242,N_9084);
and U10068 (N_10068,N_9030,N_9741);
nor U10069 (N_10069,N_9616,N_9321);
xor U10070 (N_10070,N_9378,N_9477);
xnor U10071 (N_10071,N_9603,N_9889);
and U10072 (N_10072,N_9758,N_9565);
xor U10073 (N_10073,N_9800,N_9723);
nand U10074 (N_10074,N_9722,N_9296);
nor U10075 (N_10075,N_9046,N_9818);
and U10076 (N_10076,N_9327,N_9893);
or U10077 (N_10077,N_9246,N_9634);
nor U10078 (N_10078,N_9420,N_9707);
nand U10079 (N_10079,N_9112,N_9618);
nor U10080 (N_10080,N_9266,N_9235);
nand U10081 (N_10081,N_9686,N_9807);
xor U10082 (N_10082,N_9961,N_9381);
or U10083 (N_10083,N_9127,N_9339);
nand U10084 (N_10084,N_9859,N_9457);
nor U10085 (N_10085,N_9110,N_9659);
nand U10086 (N_10086,N_9337,N_9224);
or U10087 (N_10087,N_9458,N_9731);
or U10088 (N_10088,N_9400,N_9273);
nand U10089 (N_10089,N_9422,N_9728);
nor U10090 (N_10090,N_9760,N_9911);
nor U10091 (N_10091,N_9594,N_9702);
xnor U10092 (N_10092,N_9139,N_9695);
and U10093 (N_10093,N_9667,N_9820);
or U10094 (N_10094,N_9145,N_9574);
nor U10095 (N_10095,N_9154,N_9000);
nor U10096 (N_10096,N_9472,N_9509);
and U10097 (N_10097,N_9720,N_9721);
and U10098 (N_10098,N_9923,N_9216);
nor U10099 (N_10099,N_9241,N_9952);
and U10100 (N_10100,N_9210,N_9276);
nor U10101 (N_10101,N_9045,N_9497);
or U10102 (N_10102,N_9697,N_9411);
and U10103 (N_10103,N_9260,N_9470);
or U10104 (N_10104,N_9138,N_9409);
xor U10105 (N_10105,N_9817,N_9914);
or U10106 (N_10106,N_9263,N_9134);
xnor U10107 (N_10107,N_9910,N_9732);
and U10108 (N_10108,N_9481,N_9555);
nand U10109 (N_10109,N_9028,N_9788);
and U10110 (N_10110,N_9326,N_9190);
or U10111 (N_10111,N_9692,N_9905);
nand U10112 (N_10112,N_9572,N_9249);
nand U10113 (N_10113,N_9694,N_9126);
and U10114 (N_10114,N_9730,N_9070);
nor U10115 (N_10115,N_9934,N_9488);
xor U10116 (N_10116,N_9208,N_9532);
nor U10117 (N_10117,N_9442,N_9729);
and U10118 (N_10118,N_9933,N_9736);
nand U10119 (N_10119,N_9739,N_9529);
and U10120 (N_10120,N_9974,N_9665);
nor U10121 (N_10121,N_9104,N_9330);
nand U10122 (N_10122,N_9517,N_9746);
nor U10123 (N_10123,N_9864,N_9289);
nor U10124 (N_10124,N_9450,N_9749);
nor U10125 (N_10125,N_9779,N_9931);
and U10126 (N_10126,N_9072,N_9356);
nor U10127 (N_10127,N_9412,N_9873);
nand U10128 (N_10128,N_9500,N_9150);
nand U10129 (N_10129,N_9402,N_9283);
xnor U10130 (N_10130,N_9432,N_9188);
nor U10131 (N_10131,N_9123,N_9691);
nor U10132 (N_10132,N_9384,N_9842);
nand U10133 (N_10133,N_9693,N_9365);
nor U10134 (N_10134,N_9062,N_9465);
nand U10135 (N_10135,N_9308,N_9950);
or U10136 (N_10136,N_9809,N_9999);
xnor U10137 (N_10137,N_9827,N_9226);
nor U10138 (N_10138,N_9526,N_9418);
and U10139 (N_10139,N_9593,N_9281);
and U10140 (N_10140,N_9553,N_9095);
and U10141 (N_10141,N_9832,N_9490);
or U10142 (N_10142,N_9646,N_9630);
or U10143 (N_10143,N_9074,N_9993);
or U10144 (N_10144,N_9752,N_9922);
and U10145 (N_10145,N_9124,N_9272);
or U10146 (N_10146,N_9839,N_9567);
nand U10147 (N_10147,N_9918,N_9990);
and U10148 (N_10148,N_9880,N_9921);
nand U10149 (N_10149,N_9775,N_9305);
or U10150 (N_10150,N_9082,N_9464);
or U10151 (N_10151,N_9343,N_9605);
or U10152 (N_10152,N_9533,N_9852);
or U10153 (N_10153,N_9875,N_9021);
nor U10154 (N_10154,N_9209,N_9225);
and U10155 (N_10155,N_9044,N_9878);
nor U10156 (N_10156,N_9795,N_9920);
xnor U10157 (N_10157,N_9782,N_9781);
nor U10158 (N_10158,N_9989,N_9279);
and U10159 (N_10159,N_9658,N_9774);
nor U10160 (N_10160,N_9166,N_9538);
or U10161 (N_10161,N_9217,N_9716);
nand U10162 (N_10162,N_9588,N_9566);
nor U10163 (N_10163,N_9290,N_9153);
nand U10164 (N_10164,N_9882,N_9881);
and U10165 (N_10165,N_9282,N_9613);
or U10166 (N_10166,N_9583,N_9980);
and U10167 (N_10167,N_9099,N_9743);
xor U10168 (N_10168,N_9128,N_9049);
nor U10169 (N_10169,N_9193,N_9162);
or U10170 (N_10170,N_9601,N_9709);
nor U10171 (N_10171,N_9619,N_9060);
nand U10172 (N_10172,N_9399,N_9799);
nand U10173 (N_10173,N_9669,N_9271);
and U10174 (N_10174,N_9229,N_9232);
or U10175 (N_10175,N_9704,N_9340);
nor U10176 (N_10176,N_9058,N_9194);
and U10177 (N_10177,N_9899,N_9684);
and U10178 (N_10178,N_9714,N_9847);
nand U10179 (N_10179,N_9578,N_9683);
or U10180 (N_10180,N_9003,N_9536);
nor U10181 (N_10181,N_9544,N_9186);
or U10182 (N_10182,N_9106,N_9037);
nand U10183 (N_10183,N_9906,N_9964);
nand U10184 (N_10184,N_9183,N_9495);
nand U10185 (N_10185,N_9636,N_9487);
nand U10186 (N_10186,N_9894,N_9625);
nor U10187 (N_10187,N_9372,N_9778);
nor U10188 (N_10188,N_9103,N_9170);
nand U10189 (N_10189,N_9198,N_9374);
nor U10190 (N_10190,N_9132,N_9587);
and U10191 (N_10191,N_9648,N_9168);
and U10192 (N_10192,N_9629,N_9649);
and U10193 (N_10193,N_9377,N_9551);
nor U10194 (N_10194,N_9125,N_9725);
nor U10195 (N_10195,N_9484,N_9514);
nor U10196 (N_10196,N_9328,N_9757);
and U10197 (N_10197,N_9831,N_9380);
and U10198 (N_10198,N_9024,N_9483);
and U10199 (N_10199,N_9080,N_9668);
xnor U10200 (N_10200,N_9397,N_9332);
nor U10201 (N_10201,N_9610,N_9753);
or U10202 (N_10202,N_9935,N_9401);
nor U10203 (N_10203,N_9047,N_9769);
xor U10204 (N_10204,N_9635,N_9215);
and U10205 (N_10205,N_9780,N_9115);
and U10206 (N_10206,N_9803,N_9580);
nor U10207 (N_10207,N_9883,N_9938);
nor U10208 (N_10208,N_9851,N_9267);
and U10209 (N_10209,N_9812,N_9025);
nor U10210 (N_10210,N_9268,N_9404);
nor U10211 (N_10211,N_9690,N_9227);
nand U10212 (N_10212,N_9558,N_9953);
xnor U10213 (N_10213,N_9762,N_9940);
nand U10214 (N_10214,N_9369,N_9773);
nor U10215 (N_10215,N_9158,N_9836);
nand U10216 (N_10216,N_9543,N_9203);
nor U10217 (N_10217,N_9449,N_9220);
and U10218 (N_10218,N_9681,N_9020);
nand U10219 (N_10219,N_9719,N_9396);
nand U10220 (N_10220,N_9948,N_9424);
nor U10221 (N_10221,N_9313,N_9230);
nand U10222 (N_10222,N_9231,N_9485);
or U10223 (N_10223,N_9856,N_9962);
nor U10224 (N_10224,N_9927,N_9073);
nor U10225 (N_10225,N_9007,N_9302);
and U10226 (N_10226,N_9981,N_9008);
nand U10227 (N_10227,N_9564,N_9175);
nor U10228 (N_10228,N_9791,N_9872);
or U10229 (N_10229,N_9006,N_9624);
nor U10230 (N_10230,N_9863,N_9407);
or U10231 (N_10231,N_9835,N_9523);
nand U10232 (N_10232,N_9205,N_9744);
nand U10233 (N_10233,N_9525,N_9552);
and U10234 (N_10234,N_9039,N_9674);
nand U10235 (N_10235,N_9245,N_9887);
and U10236 (N_10236,N_9687,N_9386);
xnor U10237 (N_10237,N_9383,N_9963);
nand U10238 (N_10238,N_9311,N_9785);
nor U10239 (N_10239,N_9376,N_9712);
and U10240 (N_10240,N_9958,N_9218);
and U10241 (N_10241,N_9951,N_9261);
nand U10242 (N_10242,N_9547,N_9733);
or U10243 (N_10243,N_9828,N_9391);
nand U10244 (N_10244,N_9755,N_9801);
or U10245 (N_10245,N_9367,N_9301);
nor U10246 (N_10246,N_9438,N_9997);
or U10247 (N_10247,N_9896,N_9867);
xor U10248 (N_10248,N_9575,N_9096);
nand U10249 (N_10249,N_9351,N_9454);
and U10250 (N_10250,N_9295,N_9696);
and U10251 (N_10251,N_9748,N_9429);
or U10252 (N_10252,N_9447,N_9040);
xnor U10253 (N_10253,N_9141,N_9278);
or U10254 (N_10254,N_9519,N_9761);
nor U10255 (N_10255,N_9173,N_9456);
and U10256 (N_10256,N_9647,N_9713);
and U10257 (N_10257,N_9909,N_9508);
nor U10258 (N_10258,N_9172,N_9094);
nand U10259 (N_10259,N_9109,N_9064);
nor U10260 (N_10260,N_9257,N_9065);
nor U10261 (N_10261,N_9623,N_9345);
nor U10262 (N_10262,N_9826,N_9059);
and U10263 (N_10263,N_9152,N_9554);
nor U10264 (N_10264,N_9476,N_9238);
nand U10265 (N_10265,N_9834,N_9637);
nand U10266 (N_10266,N_9892,N_9845);
or U10267 (N_10267,N_9986,N_9307);
nand U10268 (N_10268,N_9314,N_9855);
or U10269 (N_10269,N_9474,N_9419);
nor U10270 (N_10270,N_9912,N_9348);
or U10271 (N_10271,N_9854,N_9751);
nand U10272 (N_10272,N_9984,N_9416);
or U10273 (N_10273,N_9559,N_9620);
and U10274 (N_10274,N_9988,N_9297);
or U10275 (N_10275,N_9664,N_9461);
and U10276 (N_10276,N_9258,N_9041);
or U10277 (N_10277,N_9680,N_9527);
nor U10278 (N_10278,N_9363,N_9475);
or U10279 (N_10279,N_9937,N_9197);
or U10280 (N_10280,N_9585,N_9093);
nor U10281 (N_10281,N_9916,N_9165);
and U10282 (N_10282,N_9772,N_9549);
nor U10283 (N_10283,N_9898,N_9609);
or U10284 (N_10284,N_9633,N_9548);
nand U10285 (N_10285,N_9089,N_9389);
nor U10286 (N_10286,N_9582,N_9113);
and U10287 (N_10287,N_9052,N_9069);
xnor U10288 (N_10288,N_9364,N_9814);
xor U10289 (N_10289,N_9098,N_9767);
and U10290 (N_10290,N_9221,N_9129);
nand U10291 (N_10291,N_9874,N_9996);
and U10292 (N_10292,N_9862,N_9067);
nor U10293 (N_10293,N_9214,N_9632);
nor U10294 (N_10294,N_9645,N_9501);
or U10295 (N_10295,N_9119,N_9606);
xor U10296 (N_10296,N_9169,N_9195);
nor U10297 (N_10297,N_9715,N_9700);
xnor U10298 (N_10298,N_9009,N_9292);
nor U10299 (N_10299,N_9482,N_9815);
and U10300 (N_10300,N_9608,N_9983);
nand U10301 (N_10301,N_9338,N_9259);
nand U10302 (N_10302,N_9976,N_9293);
nor U10303 (N_10303,N_9954,N_9176);
nand U10304 (N_10304,N_9219,N_9848);
and U10305 (N_10305,N_9703,N_9747);
xnor U10306 (N_10306,N_9995,N_9042);
nand U10307 (N_10307,N_9653,N_9998);
and U10308 (N_10308,N_9144,N_9228);
xor U10309 (N_10309,N_9806,N_9717);
nand U10310 (N_10310,N_9121,N_9777);
xor U10311 (N_10311,N_9353,N_9434);
xor U10312 (N_10312,N_9087,N_9446);
and U10313 (N_10313,N_9902,N_9510);
nand U10314 (N_10314,N_9524,N_9698);
and U10315 (N_10315,N_9943,N_9979);
nand U10316 (N_10316,N_9448,N_9701);
nand U10317 (N_10317,N_9171,N_9222);
and U10318 (N_10318,N_9027,N_9711);
xor U10319 (N_10319,N_9316,N_9151);
nand U10320 (N_10320,N_9871,N_9395);
nor U10321 (N_10321,N_9202,N_9841);
nor U10322 (N_10322,N_9612,N_9498);
and U10323 (N_10323,N_9011,N_9960);
and U10324 (N_10324,N_9191,N_9469);
or U10325 (N_10325,N_9789,N_9738);
or U10326 (N_10326,N_9010,N_9891);
nand U10327 (N_10327,N_9393,N_9459);
xor U10328 (N_10328,N_9362,N_9120);
nor U10329 (N_10329,N_9284,N_9805);
nor U10330 (N_10330,N_9811,N_9750);
nor U10331 (N_10331,N_9427,N_9846);
nand U10332 (N_10332,N_9147,N_9247);
or U10333 (N_10333,N_9433,N_9595);
nand U10334 (N_10334,N_9866,N_9288);
nand U10335 (N_10335,N_9823,N_9159);
nand U10336 (N_10336,N_9959,N_9949);
or U10337 (N_10337,N_9201,N_9116);
nand U10338 (N_10338,N_9869,N_9079);
and U10339 (N_10339,N_9656,N_9904);
and U10340 (N_10340,N_9077,N_9798);
or U10341 (N_10341,N_9563,N_9156);
nor U10342 (N_10342,N_9287,N_9382);
nor U10343 (N_10343,N_9253,N_9868);
and U10344 (N_10344,N_9589,N_9504);
nand U10345 (N_10345,N_9861,N_9071);
nor U10346 (N_10346,N_9269,N_9405);
nor U10347 (N_10347,N_9901,N_9473);
nand U10348 (N_10348,N_9309,N_9350);
nand U10349 (N_10349,N_9844,N_9660);
and U10350 (N_10350,N_9181,N_9015);
and U10351 (N_10351,N_9813,N_9410);
xnor U10352 (N_10352,N_9163,N_9031);
nand U10353 (N_10353,N_9004,N_9392);
and U10354 (N_10354,N_9331,N_9699);
and U10355 (N_10355,N_9368,N_9824);
nor U10356 (N_10356,N_9387,N_9346);
nor U10357 (N_10357,N_9579,N_9239);
and U10358 (N_10358,N_9640,N_9143);
nor U10359 (N_10359,N_9766,N_9262);
nand U10360 (N_10360,N_9802,N_9929);
and U10361 (N_10361,N_9804,N_9592);
and U10362 (N_10362,N_9946,N_9489);
nor U10363 (N_10363,N_9333,N_9048);
and U10364 (N_10364,N_9111,N_9877);
nor U10365 (N_10365,N_9913,N_9054);
xnor U10366 (N_10366,N_9467,N_9423);
nand U10367 (N_10367,N_9496,N_9033);
or U10368 (N_10368,N_9370,N_9256);
or U10369 (N_10369,N_9535,N_9945);
and U10370 (N_10370,N_9280,N_9277);
nor U10371 (N_10371,N_9639,N_9403);
or U10372 (N_10372,N_9796,N_9677);
nand U10373 (N_10373,N_9829,N_9770);
or U10374 (N_10374,N_9135,N_9561);
nor U10375 (N_10375,N_9718,N_9068);
nand U10376 (N_10376,N_9884,N_9505);
and U10377 (N_10377,N_9614,N_9654);
xnor U10378 (N_10378,N_9727,N_9097);
nand U10379 (N_10379,N_9492,N_9942);
and U10380 (N_10380,N_9661,N_9146);
nor U10381 (N_10381,N_9542,N_9122);
nand U10382 (N_10382,N_9570,N_9255);
nor U10383 (N_10383,N_9819,N_9189);
nand U10384 (N_10384,N_9179,N_9206);
or U10385 (N_10385,N_9341,N_9971);
nor U10386 (N_10386,N_9682,N_9671);
and U10387 (N_10387,N_9018,N_9439);
nand U10388 (N_10388,N_9840,N_9310);
and U10389 (N_10389,N_9270,N_9786);
or U10390 (N_10390,N_9833,N_9462);
nand U10391 (N_10391,N_9056,N_9972);
and U10392 (N_10392,N_9430,N_9413);
and U10393 (N_10393,N_9038,N_9967);
and U10394 (N_10394,N_9604,N_9349);
nand U10395 (N_10395,N_9977,N_9792);
nor U10396 (N_10396,N_9357,N_9797);
or U10397 (N_10397,N_9573,N_9265);
and U10398 (N_10398,N_9001,N_9765);
and U10399 (N_10399,N_9086,N_9768);
or U10400 (N_10400,N_9105,N_9771);
nor U10401 (N_10401,N_9088,N_9300);
nand U10402 (N_10402,N_9759,N_9398);
nand U10403 (N_10403,N_9621,N_9026);
and U10404 (N_10404,N_9092,N_9985);
nand U10405 (N_10405,N_9101,N_9735);
and U10406 (N_10406,N_9479,N_9013);
or U10407 (N_10407,N_9354,N_9285);
and U10408 (N_10408,N_9673,N_9537);
and U10409 (N_10409,N_9888,N_9513);
nor U10410 (N_10410,N_9428,N_9885);
or U10411 (N_10411,N_9638,N_9352);
or U10412 (N_10412,N_9233,N_9503);
nand U10413 (N_10413,N_9076,N_9303);
and U10414 (N_10414,N_9666,N_9196);
nor U10415 (N_10415,N_9708,N_9066);
nand U10416 (N_10416,N_9291,N_9655);
or U10417 (N_10417,N_9742,N_9919);
or U10418 (N_10418,N_9319,N_9850);
or U10419 (N_10419,N_9294,N_9032);
and U10420 (N_10420,N_9359,N_9598);
and U10421 (N_10421,N_9157,N_9685);
or U10422 (N_10422,N_9571,N_9790);
nor U10423 (N_10423,N_9876,N_9947);
or U10424 (N_10424,N_9688,N_9679);
nor U10425 (N_10425,N_9966,N_9915);
and U10426 (N_10426,N_9545,N_9182);
nor U10427 (N_10427,N_9546,N_9689);
or U10428 (N_10428,N_9445,N_9136);
nor U10429 (N_10429,N_9969,N_9978);
nand U10430 (N_10430,N_9426,N_9511);
and U10431 (N_10431,N_9794,N_9417);
nand U10432 (N_10432,N_9822,N_9315);
or U10433 (N_10433,N_9252,N_9576);
or U10434 (N_10434,N_9207,N_9641);
or U10435 (N_10435,N_9375,N_9415);
nand U10436 (N_10436,N_9895,N_9541);
or U10437 (N_10437,N_9298,N_9675);
or U10438 (N_10438,N_9539,N_9520);
and U10439 (N_10439,N_9617,N_9493);
or U10440 (N_10440,N_9108,N_9973);
nor U10441 (N_10441,N_9274,N_9651);
nor U10442 (N_10442,N_9244,N_9167);
nand U10443 (N_10443,N_9502,N_9740);
xor U10444 (N_10444,N_9234,N_9441);
or U10445 (N_10445,N_9466,N_9499);
nor U10446 (N_10446,N_9644,N_9455);
nand U10447 (N_10447,N_9965,N_9443);
nand U10448 (N_10448,N_9090,N_9600);
and U10449 (N_10449,N_9204,N_9793);
and U10450 (N_10450,N_9373,N_9591);
and U10451 (N_10451,N_9431,N_9597);
or U10452 (N_10452,N_9133,N_9440);
and U10453 (N_10453,N_9248,N_9329);
and U10454 (N_10454,N_9016,N_9444);
xor U10455 (N_10455,N_9908,N_9783);
and U10456 (N_10456,N_9764,N_9421);
or U10457 (N_10457,N_9596,N_9557);
and U10458 (N_10458,N_9886,N_9005);
or U10459 (N_10459,N_9390,N_9982);
nand U10460 (N_10460,N_9081,N_9371);
or U10461 (N_10461,N_9857,N_9754);
nand U10462 (N_10462,N_9870,N_9361);
xor U10463 (N_10463,N_9642,N_9932);
nand U10464 (N_10464,N_9083,N_9843);
or U10465 (N_10465,N_9200,N_9325);
nand U10466 (N_10466,N_9453,N_9486);
or U10467 (N_10467,N_9615,N_9036);
nor U10468 (N_10468,N_9560,N_9468);
nor U10469 (N_10469,N_9924,N_9516);
and U10470 (N_10470,N_9435,N_9320);
nor U10471 (N_10471,N_9019,N_9029);
xnor U10472 (N_10472,N_9491,N_9184);
nand U10473 (N_10473,N_9531,N_9837);
or U10474 (N_10474,N_9131,N_9275);
or U10475 (N_10475,N_9534,N_9355);
nand U10476 (N_10476,N_9137,N_9471);
and U10477 (N_10477,N_9114,N_9590);
nor U10478 (N_10478,N_9663,N_9149);
nor U10479 (N_10479,N_9142,N_9607);
or U10480 (N_10480,N_9406,N_9211);
xnor U10481 (N_10481,N_9379,N_9926);
and U10482 (N_10482,N_9388,N_9939);
nand U10483 (N_10483,N_9956,N_9160);
and U10484 (N_10484,N_9518,N_9678);
or U10485 (N_10485,N_9745,N_9140);
xnor U10486 (N_10486,N_9903,N_9322);
nor U10487 (N_10487,N_9930,N_9334);
or U10488 (N_10488,N_9512,N_9611);
nand U10489 (N_10489,N_9251,N_9540);
nor U10490 (N_10490,N_9941,N_9425);
nand U10491 (N_10491,N_9102,N_9970);
nor U10492 (N_10492,N_9705,N_9117);
and U10493 (N_10493,N_9657,N_9414);
or U10494 (N_10494,N_9061,N_9192);
xor U10495 (N_10495,N_9264,N_9318);
nor U10496 (N_10496,N_9185,N_9324);
and U10497 (N_10497,N_9323,N_9075);
or U10498 (N_10498,N_9562,N_9991);
nand U10499 (N_10499,N_9810,N_9830);
nor U10500 (N_10500,N_9064,N_9609);
and U10501 (N_10501,N_9196,N_9129);
nand U10502 (N_10502,N_9682,N_9829);
nor U10503 (N_10503,N_9028,N_9925);
or U10504 (N_10504,N_9354,N_9764);
and U10505 (N_10505,N_9966,N_9994);
or U10506 (N_10506,N_9143,N_9319);
or U10507 (N_10507,N_9304,N_9267);
nand U10508 (N_10508,N_9497,N_9937);
nand U10509 (N_10509,N_9307,N_9472);
nand U10510 (N_10510,N_9928,N_9115);
nand U10511 (N_10511,N_9739,N_9324);
xor U10512 (N_10512,N_9675,N_9756);
nand U10513 (N_10513,N_9562,N_9760);
and U10514 (N_10514,N_9549,N_9824);
xor U10515 (N_10515,N_9798,N_9540);
xnor U10516 (N_10516,N_9132,N_9705);
and U10517 (N_10517,N_9725,N_9290);
and U10518 (N_10518,N_9698,N_9898);
and U10519 (N_10519,N_9435,N_9562);
nor U10520 (N_10520,N_9814,N_9940);
xnor U10521 (N_10521,N_9804,N_9715);
xnor U10522 (N_10522,N_9994,N_9667);
xnor U10523 (N_10523,N_9932,N_9724);
nor U10524 (N_10524,N_9583,N_9190);
nand U10525 (N_10525,N_9182,N_9223);
nand U10526 (N_10526,N_9582,N_9130);
and U10527 (N_10527,N_9486,N_9696);
and U10528 (N_10528,N_9217,N_9880);
or U10529 (N_10529,N_9274,N_9338);
nor U10530 (N_10530,N_9103,N_9115);
or U10531 (N_10531,N_9085,N_9077);
or U10532 (N_10532,N_9513,N_9781);
nor U10533 (N_10533,N_9210,N_9932);
or U10534 (N_10534,N_9465,N_9470);
or U10535 (N_10535,N_9885,N_9668);
xnor U10536 (N_10536,N_9559,N_9394);
nor U10537 (N_10537,N_9883,N_9851);
nand U10538 (N_10538,N_9224,N_9478);
nor U10539 (N_10539,N_9825,N_9684);
nand U10540 (N_10540,N_9806,N_9402);
nand U10541 (N_10541,N_9660,N_9148);
and U10542 (N_10542,N_9461,N_9745);
and U10543 (N_10543,N_9859,N_9474);
nand U10544 (N_10544,N_9426,N_9218);
nand U10545 (N_10545,N_9649,N_9610);
nand U10546 (N_10546,N_9355,N_9591);
or U10547 (N_10547,N_9711,N_9552);
nand U10548 (N_10548,N_9510,N_9434);
nand U10549 (N_10549,N_9278,N_9075);
nor U10550 (N_10550,N_9784,N_9609);
xor U10551 (N_10551,N_9439,N_9950);
and U10552 (N_10552,N_9903,N_9614);
and U10553 (N_10553,N_9034,N_9289);
and U10554 (N_10554,N_9733,N_9665);
and U10555 (N_10555,N_9266,N_9559);
xnor U10556 (N_10556,N_9164,N_9321);
nor U10557 (N_10557,N_9739,N_9941);
nor U10558 (N_10558,N_9831,N_9738);
nand U10559 (N_10559,N_9879,N_9065);
nand U10560 (N_10560,N_9120,N_9403);
nor U10561 (N_10561,N_9883,N_9064);
nor U10562 (N_10562,N_9331,N_9324);
or U10563 (N_10563,N_9378,N_9618);
nor U10564 (N_10564,N_9723,N_9141);
or U10565 (N_10565,N_9649,N_9152);
or U10566 (N_10566,N_9460,N_9871);
and U10567 (N_10567,N_9877,N_9888);
nor U10568 (N_10568,N_9674,N_9954);
nand U10569 (N_10569,N_9370,N_9714);
nor U10570 (N_10570,N_9816,N_9653);
or U10571 (N_10571,N_9383,N_9448);
and U10572 (N_10572,N_9012,N_9341);
nand U10573 (N_10573,N_9070,N_9575);
or U10574 (N_10574,N_9323,N_9544);
xnor U10575 (N_10575,N_9072,N_9905);
or U10576 (N_10576,N_9123,N_9902);
and U10577 (N_10577,N_9629,N_9401);
or U10578 (N_10578,N_9289,N_9119);
or U10579 (N_10579,N_9232,N_9738);
nor U10580 (N_10580,N_9545,N_9014);
or U10581 (N_10581,N_9689,N_9143);
and U10582 (N_10582,N_9979,N_9688);
or U10583 (N_10583,N_9909,N_9801);
or U10584 (N_10584,N_9309,N_9897);
xnor U10585 (N_10585,N_9117,N_9743);
or U10586 (N_10586,N_9532,N_9391);
and U10587 (N_10587,N_9186,N_9055);
nand U10588 (N_10588,N_9720,N_9102);
nand U10589 (N_10589,N_9299,N_9443);
and U10590 (N_10590,N_9442,N_9193);
and U10591 (N_10591,N_9592,N_9057);
nor U10592 (N_10592,N_9536,N_9612);
nand U10593 (N_10593,N_9692,N_9799);
and U10594 (N_10594,N_9665,N_9795);
xnor U10595 (N_10595,N_9460,N_9096);
nand U10596 (N_10596,N_9207,N_9114);
and U10597 (N_10597,N_9462,N_9250);
nor U10598 (N_10598,N_9600,N_9037);
nor U10599 (N_10599,N_9402,N_9211);
or U10600 (N_10600,N_9120,N_9921);
nor U10601 (N_10601,N_9106,N_9454);
nor U10602 (N_10602,N_9758,N_9573);
nand U10603 (N_10603,N_9207,N_9439);
or U10604 (N_10604,N_9940,N_9894);
or U10605 (N_10605,N_9884,N_9168);
nor U10606 (N_10606,N_9565,N_9772);
nand U10607 (N_10607,N_9032,N_9222);
or U10608 (N_10608,N_9776,N_9404);
nand U10609 (N_10609,N_9957,N_9434);
or U10610 (N_10610,N_9022,N_9139);
or U10611 (N_10611,N_9559,N_9500);
nand U10612 (N_10612,N_9863,N_9691);
or U10613 (N_10613,N_9782,N_9808);
and U10614 (N_10614,N_9178,N_9674);
xor U10615 (N_10615,N_9812,N_9027);
and U10616 (N_10616,N_9070,N_9194);
or U10617 (N_10617,N_9850,N_9603);
or U10618 (N_10618,N_9832,N_9082);
and U10619 (N_10619,N_9666,N_9066);
or U10620 (N_10620,N_9088,N_9588);
nand U10621 (N_10621,N_9963,N_9485);
nor U10622 (N_10622,N_9029,N_9537);
and U10623 (N_10623,N_9744,N_9251);
nand U10624 (N_10624,N_9154,N_9508);
and U10625 (N_10625,N_9031,N_9075);
or U10626 (N_10626,N_9333,N_9012);
and U10627 (N_10627,N_9288,N_9311);
nor U10628 (N_10628,N_9930,N_9201);
xor U10629 (N_10629,N_9961,N_9761);
and U10630 (N_10630,N_9407,N_9146);
or U10631 (N_10631,N_9679,N_9100);
and U10632 (N_10632,N_9792,N_9648);
or U10633 (N_10633,N_9741,N_9363);
or U10634 (N_10634,N_9571,N_9636);
or U10635 (N_10635,N_9381,N_9108);
or U10636 (N_10636,N_9321,N_9557);
nand U10637 (N_10637,N_9910,N_9834);
or U10638 (N_10638,N_9927,N_9573);
and U10639 (N_10639,N_9345,N_9208);
or U10640 (N_10640,N_9603,N_9458);
or U10641 (N_10641,N_9164,N_9044);
nor U10642 (N_10642,N_9016,N_9761);
nand U10643 (N_10643,N_9018,N_9919);
and U10644 (N_10644,N_9192,N_9281);
or U10645 (N_10645,N_9321,N_9666);
nor U10646 (N_10646,N_9841,N_9853);
nor U10647 (N_10647,N_9727,N_9064);
and U10648 (N_10648,N_9198,N_9138);
or U10649 (N_10649,N_9463,N_9291);
or U10650 (N_10650,N_9060,N_9163);
or U10651 (N_10651,N_9428,N_9860);
and U10652 (N_10652,N_9670,N_9792);
nand U10653 (N_10653,N_9363,N_9721);
nand U10654 (N_10654,N_9666,N_9505);
or U10655 (N_10655,N_9013,N_9791);
or U10656 (N_10656,N_9258,N_9338);
nor U10657 (N_10657,N_9291,N_9070);
nor U10658 (N_10658,N_9721,N_9289);
and U10659 (N_10659,N_9255,N_9525);
nand U10660 (N_10660,N_9404,N_9636);
and U10661 (N_10661,N_9524,N_9395);
and U10662 (N_10662,N_9099,N_9422);
and U10663 (N_10663,N_9452,N_9459);
and U10664 (N_10664,N_9053,N_9104);
or U10665 (N_10665,N_9212,N_9710);
nor U10666 (N_10666,N_9621,N_9123);
or U10667 (N_10667,N_9688,N_9310);
nand U10668 (N_10668,N_9510,N_9781);
nand U10669 (N_10669,N_9973,N_9638);
nand U10670 (N_10670,N_9608,N_9060);
nor U10671 (N_10671,N_9090,N_9073);
and U10672 (N_10672,N_9876,N_9173);
nand U10673 (N_10673,N_9864,N_9239);
or U10674 (N_10674,N_9360,N_9795);
and U10675 (N_10675,N_9800,N_9698);
or U10676 (N_10676,N_9440,N_9715);
or U10677 (N_10677,N_9364,N_9556);
nor U10678 (N_10678,N_9939,N_9904);
and U10679 (N_10679,N_9207,N_9623);
nor U10680 (N_10680,N_9320,N_9932);
nand U10681 (N_10681,N_9845,N_9429);
nor U10682 (N_10682,N_9943,N_9225);
and U10683 (N_10683,N_9248,N_9169);
nand U10684 (N_10684,N_9903,N_9641);
or U10685 (N_10685,N_9643,N_9900);
nor U10686 (N_10686,N_9357,N_9883);
nor U10687 (N_10687,N_9876,N_9321);
nand U10688 (N_10688,N_9124,N_9922);
or U10689 (N_10689,N_9764,N_9902);
nor U10690 (N_10690,N_9751,N_9248);
nand U10691 (N_10691,N_9905,N_9609);
and U10692 (N_10692,N_9452,N_9990);
nand U10693 (N_10693,N_9210,N_9043);
and U10694 (N_10694,N_9816,N_9096);
nand U10695 (N_10695,N_9465,N_9046);
or U10696 (N_10696,N_9658,N_9821);
nor U10697 (N_10697,N_9664,N_9502);
nand U10698 (N_10698,N_9933,N_9113);
nor U10699 (N_10699,N_9737,N_9409);
nand U10700 (N_10700,N_9384,N_9672);
or U10701 (N_10701,N_9903,N_9960);
or U10702 (N_10702,N_9266,N_9373);
xnor U10703 (N_10703,N_9748,N_9865);
xnor U10704 (N_10704,N_9059,N_9003);
or U10705 (N_10705,N_9478,N_9788);
and U10706 (N_10706,N_9785,N_9543);
and U10707 (N_10707,N_9903,N_9101);
nor U10708 (N_10708,N_9477,N_9723);
or U10709 (N_10709,N_9530,N_9087);
nand U10710 (N_10710,N_9299,N_9774);
nand U10711 (N_10711,N_9907,N_9418);
nand U10712 (N_10712,N_9696,N_9266);
or U10713 (N_10713,N_9971,N_9937);
nand U10714 (N_10714,N_9986,N_9171);
xor U10715 (N_10715,N_9626,N_9738);
xor U10716 (N_10716,N_9845,N_9838);
nand U10717 (N_10717,N_9017,N_9125);
and U10718 (N_10718,N_9492,N_9638);
and U10719 (N_10719,N_9800,N_9579);
nor U10720 (N_10720,N_9255,N_9440);
nand U10721 (N_10721,N_9503,N_9995);
nor U10722 (N_10722,N_9829,N_9732);
nand U10723 (N_10723,N_9096,N_9544);
or U10724 (N_10724,N_9681,N_9886);
xor U10725 (N_10725,N_9431,N_9345);
or U10726 (N_10726,N_9933,N_9508);
nor U10727 (N_10727,N_9501,N_9826);
nor U10728 (N_10728,N_9337,N_9255);
nand U10729 (N_10729,N_9676,N_9826);
or U10730 (N_10730,N_9252,N_9126);
and U10731 (N_10731,N_9595,N_9535);
and U10732 (N_10732,N_9642,N_9700);
nor U10733 (N_10733,N_9055,N_9516);
nand U10734 (N_10734,N_9577,N_9976);
and U10735 (N_10735,N_9275,N_9394);
or U10736 (N_10736,N_9205,N_9724);
nor U10737 (N_10737,N_9436,N_9057);
and U10738 (N_10738,N_9953,N_9763);
nand U10739 (N_10739,N_9690,N_9652);
and U10740 (N_10740,N_9794,N_9980);
nand U10741 (N_10741,N_9391,N_9182);
nor U10742 (N_10742,N_9501,N_9070);
or U10743 (N_10743,N_9653,N_9285);
nand U10744 (N_10744,N_9235,N_9502);
nor U10745 (N_10745,N_9192,N_9877);
and U10746 (N_10746,N_9174,N_9415);
nand U10747 (N_10747,N_9084,N_9373);
nor U10748 (N_10748,N_9517,N_9899);
nor U10749 (N_10749,N_9281,N_9909);
and U10750 (N_10750,N_9583,N_9959);
xnor U10751 (N_10751,N_9772,N_9502);
and U10752 (N_10752,N_9204,N_9869);
nand U10753 (N_10753,N_9844,N_9988);
nand U10754 (N_10754,N_9080,N_9684);
or U10755 (N_10755,N_9042,N_9893);
nand U10756 (N_10756,N_9839,N_9723);
nor U10757 (N_10757,N_9838,N_9918);
and U10758 (N_10758,N_9749,N_9207);
or U10759 (N_10759,N_9981,N_9012);
or U10760 (N_10760,N_9673,N_9224);
and U10761 (N_10761,N_9603,N_9559);
and U10762 (N_10762,N_9556,N_9974);
nand U10763 (N_10763,N_9590,N_9151);
nor U10764 (N_10764,N_9170,N_9195);
nor U10765 (N_10765,N_9866,N_9640);
nand U10766 (N_10766,N_9042,N_9287);
and U10767 (N_10767,N_9880,N_9288);
and U10768 (N_10768,N_9005,N_9465);
and U10769 (N_10769,N_9854,N_9889);
or U10770 (N_10770,N_9051,N_9429);
or U10771 (N_10771,N_9964,N_9030);
or U10772 (N_10772,N_9940,N_9767);
nand U10773 (N_10773,N_9708,N_9726);
and U10774 (N_10774,N_9352,N_9587);
and U10775 (N_10775,N_9637,N_9838);
and U10776 (N_10776,N_9992,N_9885);
nor U10777 (N_10777,N_9619,N_9066);
nand U10778 (N_10778,N_9774,N_9708);
and U10779 (N_10779,N_9243,N_9257);
or U10780 (N_10780,N_9463,N_9884);
and U10781 (N_10781,N_9863,N_9222);
xor U10782 (N_10782,N_9527,N_9115);
nor U10783 (N_10783,N_9171,N_9089);
nor U10784 (N_10784,N_9277,N_9766);
or U10785 (N_10785,N_9284,N_9866);
and U10786 (N_10786,N_9939,N_9041);
nor U10787 (N_10787,N_9094,N_9898);
and U10788 (N_10788,N_9208,N_9082);
nor U10789 (N_10789,N_9358,N_9004);
nand U10790 (N_10790,N_9065,N_9178);
nor U10791 (N_10791,N_9474,N_9359);
xnor U10792 (N_10792,N_9117,N_9463);
or U10793 (N_10793,N_9592,N_9987);
or U10794 (N_10794,N_9833,N_9489);
and U10795 (N_10795,N_9949,N_9967);
nand U10796 (N_10796,N_9127,N_9903);
or U10797 (N_10797,N_9169,N_9003);
and U10798 (N_10798,N_9536,N_9942);
or U10799 (N_10799,N_9121,N_9240);
and U10800 (N_10800,N_9977,N_9326);
xnor U10801 (N_10801,N_9689,N_9614);
nand U10802 (N_10802,N_9118,N_9222);
and U10803 (N_10803,N_9676,N_9344);
and U10804 (N_10804,N_9838,N_9294);
and U10805 (N_10805,N_9198,N_9102);
nand U10806 (N_10806,N_9489,N_9591);
and U10807 (N_10807,N_9704,N_9077);
nor U10808 (N_10808,N_9534,N_9612);
nor U10809 (N_10809,N_9998,N_9233);
nor U10810 (N_10810,N_9219,N_9429);
nand U10811 (N_10811,N_9521,N_9691);
nor U10812 (N_10812,N_9881,N_9011);
nand U10813 (N_10813,N_9842,N_9213);
nor U10814 (N_10814,N_9624,N_9501);
or U10815 (N_10815,N_9274,N_9109);
or U10816 (N_10816,N_9000,N_9707);
and U10817 (N_10817,N_9202,N_9054);
and U10818 (N_10818,N_9383,N_9036);
or U10819 (N_10819,N_9808,N_9389);
and U10820 (N_10820,N_9887,N_9601);
nand U10821 (N_10821,N_9428,N_9743);
nand U10822 (N_10822,N_9937,N_9131);
and U10823 (N_10823,N_9884,N_9826);
nand U10824 (N_10824,N_9617,N_9584);
or U10825 (N_10825,N_9195,N_9320);
and U10826 (N_10826,N_9218,N_9698);
and U10827 (N_10827,N_9478,N_9479);
or U10828 (N_10828,N_9278,N_9496);
or U10829 (N_10829,N_9618,N_9954);
nor U10830 (N_10830,N_9869,N_9454);
nor U10831 (N_10831,N_9273,N_9448);
or U10832 (N_10832,N_9325,N_9802);
or U10833 (N_10833,N_9269,N_9952);
or U10834 (N_10834,N_9026,N_9305);
nor U10835 (N_10835,N_9557,N_9230);
or U10836 (N_10836,N_9453,N_9653);
nor U10837 (N_10837,N_9078,N_9470);
or U10838 (N_10838,N_9345,N_9226);
and U10839 (N_10839,N_9746,N_9721);
nor U10840 (N_10840,N_9462,N_9488);
nor U10841 (N_10841,N_9806,N_9311);
and U10842 (N_10842,N_9174,N_9172);
nand U10843 (N_10843,N_9901,N_9035);
and U10844 (N_10844,N_9308,N_9210);
nor U10845 (N_10845,N_9115,N_9714);
or U10846 (N_10846,N_9827,N_9181);
nor U10847 (N_10847,N_9855,N_9363);
or U10848 (N_10848,N_9455,N_9656);
nor U10849 (N_10849,N_9020,N_9322);
nor U10850 (N_10850,N_9718,N_9549);
nand U10851 (N_10851,N_9015,N_9324);
nor U10852 (N_10852,N_9460,N_9004);
xnor U10853 (N_10853,N_9791,N_9878);
or U10854 (N_10854,N_9071,N_9181);
nor U10855 (N_10855,N_9297,N_9640);
and U10856 (N_10856,N_9119,N_9041);
or U10857 (N_10857,N_9823,N_9781);
nor U10858 (N_10858,N_9376,N_9941);
nor U10859 (N_10859,N_9262,N_9936);
nor U10860 (N_10860,N_9286,N_9525);
nor U10861 (N_10861,N_9303,N_9288);
or U10862 (N_10862,N_9966,N_9415);
nand U10863 (N_10863,N_9713,N_9402);
or U10864 (N_10864,N_9419,N_9953);
nor U10865 (N_10865,N_9617,N_9173);
nor U10866 (N_10866,N_9550,N_9025);
nor U10867 (N_10867,N_9774,N_9743);
xor U10868 (N_10868,N_9662,N_9744);
or U10869 (N_10869,N_9237,N_9249);
and U10870 (N_10870,N_9528,N_9460);
or U10871 (N_10871,N_9841,N_9185);
or U10872 (N_10872,N_9392,N_9441);
nand U10873 (N_10873,N_9074,N_9945);
and U10874 (N_10874,N_9917,N_9934);
nor U10875 (N_10875,N_9685,N_9110);
or U10876 (N_10876,N_9870,N_9132);
and U10877 (N_10877,N_9006,N_9372);
nand U10878 (N_10878,N_9791,N_9843);
and U10879 (N_10879,N_9336,N_9479);
nor U10880 (N_10880,N_9436,N_9286);
nand U10881 (N_10881,N_9476,N_9483);
nor U10882 (N_10882,N_9806,N_9262);
nand U10883 (N_10883,N_9041,N_9607);
nor U10884 (N_10884,N_9704,N_9630);
and U10885 (N_10885,N_9225,N_9343);
or U10886 (N_10886,N_9290,N_9149);
xnor U10887 (N_10887,N_9646,N_9664);
or U10888 (N_10888,N_9062,N_9121);
xnor U10889 (N_10889,N_9787,N_9306);
and U10890 (N_10890,N_9952,N_9346);
nor U10891 (N_10891,N_9930,N_9053);
and U10892 (N_10892,N_9496,N_9914);
xor U10893 (N_10893,N_9046,N_9718);
or U10894 (N_10894,N_9270,N_9011);
or U10895 (N_10895,N_9463,N_9316);
nor U10896 (N_10896,N_9417,N_9186);
nand U10897 (N_10897,N_9275,N_9831);
and U10898 (N_10898,N_9960,N_9235);
and U10899 (N_10899,N_9773,N_9913);
nand U10900 (N_10900,N_9477,N_9955);
nor U10901 (N_10901,N_9944,N_9795);
or U10902 (N_10902,N_9621,N_9303);
nor U10903 (N_10903,N_9600,N_9424);
or U10904 (N_10904,N_9087,N_9832);
and U10905 (N_10905,N_9552,N_9148);
or U10906 (N_10906,N_9497,N_9431);
and U10907 (N_10907,N_9197,N_9426);
nor U10908 (N_10908,N_9928,N_9463);
and U10909 (N_10909,N_9395,N_9557);
or U10910 (N_10910,N_9739,N_9144);
nand U10911 (N_10911,N_9550,N_9808);
nand U10912 (N_10912,N_9403,N_9506);
xor U10913 (N_10913,N_9398,N_9380);
and U10914 (N_10914,N_9361,N_9190);
and U10915 (N_10915,N_9188,N_9770);
xnor U10916 (N_10916,N_9199,N_9195);
or U10917 (N_10917,N_9222,N_9669);
nand U10918 (N_10918,N_9628,N_9776);
xnor U10919 (N_10919,N_9849,N_9627);
nor U10920 (N_10920,N_9270,N_9964);
nand U10921 (N_10921,N_9553,N_9742);
nor U10922 (N_10922,N_9772,N_9146);
xnor U10923 (N_10923,N_9472,N_9630);
and U10924 (N_10924,N_9641,N_9267);
or U10925 (N_10925,N_9590,N_9417);
xnor U10926 (N_10926,N_9298,N_9848);
nor U10927 (N_10927,N_9277,N_9186);
or U10928 (N_10928,N_9600,N_9170);
or U10929 (N_10929,N_9756,N_9149);
nor U10930 (N_10930,N_9950,N_9772);
or U10931 (N_10931,N_9733,N_9210);
or U10932 (N_10932,N_9422,N_9429);
and U10933 (N_10933,N_9301,N_9677);
nor U10934 (N_10934,N_9104,N_9623);
nor U10935 (N_10935,N_9193,N_9822);
nor U10936 (N_10936,N_9470,N_9885);
or U10937 (N_10937,N_9478,N_9390);
and U10938 (N_10938,N_9976,N_9768);
nor U10939 (N_10939,N_9567,N_9428);
or U10940 (N_10940,N_9051,N_9719);
or U10941 (N_10941,N_9116,N_9704);
nand U10942 (N_10942,N_9398,N_9992);
and U10943 (N_10943,N_9180,N_9464);
nand U10944 (N_10944,N_9332,N_9606);
nand U10945 (N_10945,N_9212,N_9480);
nor U10946 (N_10946,N_9482,N_9638);
nand U10947 (N_10947,N_9454,N_9239);
or U10948 (N_10948,N_9646,N_9556);
nand U10949 (N_10949,N_9385,N_9125);
or U10950 (N_10950,N_9052,N_9906);
or U10951 (N_10951,N_9391,N_9663);
nor U10952 (N_10952,N_9664,N_9823);
nor U10953 (N_10953,N_9913,N_9121);
nand U10954 (N_10954,N_9199,N_9601);
nor U10955 (N_10955,N_9411,N_9385);
and U10956 (N_10956,N_9282,N_9079);
nand U10957 (N_10957,N_9076,N_9407);
nor U10958 (N_10958,N_9808,N_9605);
or U10959 (N_10959,N_9812,N_9017);
nor U10960 (N_10960,N_9756,N_9666);
and U10961 (N_10961,N_9567,N_9665);
and U10962 (N_10962,N_9495,N_9869);
or U10963 (N_10963,N_9400,N_9975);
or U10964 (N_10964,N_9871,N_9711);
or U10965 (N_10965,N_9099,N_9666);
xor U10966 (N_10966,N_9133,N_9724);
and U10967 (N_10967,N_9532,N_9283);
or U10968 (N_10968,N_9616,N_9266);
and U10969 (N_10969,N_9183,N_9325);
nor U10970 (N_10970,N_9792,N_9120);
xnor U10971 (N_10971,N_9886,N_9641);
nor U10972 (N_10972,N_9609,N_9803);
or U10973 (N_10973,N_9486,N_9562);
nand U10974 (N_10974,N_9267,N_9061);
nand U10975 (N_10975,N_9251,N_9638);
and U10976 (N_10976,N_9293,N_9640);
nor U10977 (N_10977,N_9871,N_9927);
nor U10978 (N_10978,N_9865,N_9699);
and U10979 (N_10979,N_9437,N_9063);
xnor U10980 (N_10980,N_9513,N_9230);
or U10981 (N_10981,N_9981,N_9889);
or U10982 (N_10982,N_9969,N_9029);
nand U10983 (N_10983,N_9766,N_9116);
xor U10984 (N_10984,N_9518,N_9311);
nor U10985 (N_10985,N_9049,N_9540);
and U10986 (N_10986,N_9239,N_9169);
nand U10987 (N_10987,N_9601,N_9039);
nor U10988 (N_10988,N_9926,N_9415);
nor U10989 (N_10989,N_9946,N_9525);
and U10990 (N_10990,N_9058,N_9015);
and U10991 (N_10991,N_9018,N_9149);
or U10992 (N_10992,N_9670,N_9131);
or U10993 (N_10993,N_9378,N_9207);
and U10994 (N_10994,N_9035,N_9423);
and U10995 (N_10995,N_9753,N_9769);
and U10996 (N_10996,N_9600,N_9561);
and U10997 (N_10997,N_9925,N_9470);
and U10998 (N_10998,N_9003,N_9376);
nand U10999 (N_10999,N_9278,N_9706);
nor U11000 (N_11000,N_10107,N_10327);
nor U11001 (N_11001,N_10759,N_10893);
or U11002 (N_11002,N_10794,N_10095);
or U11003 (N_11003,N_10525,N_10684);
nor U11004 (N_11004,N_10260,N_10307);
and U11005 (N_11005,N_10408,N_10962);
and U11006 (N_11006,N_10083,N_10922);
nor U11007 (N_11007,N_10835,N_10057);
xor U11008 (N_11008,N_10556,N_10725);
xor U11009 (N_11009,N_10217,N_10886);
and U11010 (N_11010,N_10346,N_10477);
or U11011 (N_11011,N_10388,N_10843);
and U11012 (N_11012,N_10180,N_10741);
or U11013 (N_11013,N_10980,N_10324);
nor U11014 (N_11014,N_10310,N_10861);
or U11015 (N_11015,N_10281,N_10892);
nand U11016 (N_11016,N_10943,N_10485);
and U11017 (N_11017,N_10448,N_10969);
nor U11018 (N_11018,N_10793,N_10986);
xnor U11019 (N_11019,N_10070,N_10520);
nand U11020 (N_11020,N_10589,N_10784);
nand U11021 (N_11021,N_10930,N_10467);
nand U11022 (N_11022,N_10523,N_10912);
or U11023 (N_11023,N_10438,N_10689);
and U11024 (N_11024,N_10352,N_10361);
and U11025 (N_11025,N_10919,N_10472);
or U11026 (N_11026,N_10531,N_10109);
nor U11027 (N_11027,N_10380,N_10179);
nor U11028 (N_11028,N_10860,N_10096);
or U11029 (N_11029,N_10419,N_10123);
nor U11030 (N_11030,N_10937,N_10271);
and U11031 (N_11031,N_10965,N_10062);
xor U11032 (N_11032,N_10553,N_10368);
nand U11033 (N_11033,N_10124,N_10960);
or U11034 (N_11034,N_10133,N_10118);
or U11035 (N_11035,N_10596,N_10780);
and U11036 (N_11036,N_10158,N_10246);
and U11037 (N_11037,N_10293,N_10471);
or U11038 (N_11038,N_10239,N_10611);
nand U11039 (N_11039,N_10775,N_10480);
nor U11040 (N_11040,N_10474,N_10046);
xor U11041 (N_11041,N_10598,N_10848);
xor U11042 (N_11042,N_10989,N_10787);
xor U11043 (N_11043,N_10837,N_10898);
or U11044 (N_11044,N_10444,N_10134);
and U11045 (N_11045,N_10853,N_10103);
nor U11046 (N_11046,N_10509,N_10997);
nor U11047 (N_11047,N_10889,N_10156);
xor U11048 (N_11048,N_10636,N_10857);
or U11049 (N_11049,N_10617,N_10667);
or U11050 (N_11050,N_10334,N_10802);
nor U11051 (N_11051,N_10503,N_10573);
and U11052 (N_11052,N_10849,N_10588);
nand U11053 (N_11053,N_10265,N_10342);
nand U11054 (N_11054,N_10259,N_10884);
nor U11055 (N_11055,N_10097,N_10543);
or U11056 (N_11056,N_10079,N_10982);
nand U11057 (N_11057,N_10195,N_10401);
nand U11058 (N_11058,N_10882,N_10755);
or U11059 (N_11059,N_10938,N_10493);
nor U11060 (N_11060,N_10351,N_10619);
nand U11061 (N_11061,N_10582,N_10215);
nand U11062 (N_11062,N_10385,N_10516);
or U11063 (N_11063,N_10397,N_10491);
or U11064 (N_11064,N_10150,N_10717);
and U11065 (N_11065,N_10534,N_10439);
or U11066 (N_11066,N_10384,N_10470);
and U11067 (N_11067,N_10428,N_10077);
xor U11068 (N_11068,N_10946,N_10277);
and U11069 (N_11069,N_10216,N_10931);
or U11070 (N_11070,N_10068,N_10526);
nand U11071 (N_11071,N_10866,N_10869);
and U11072 (N_11072,N_10492,N_10443);
nor U11073 (N_11073,N_10942,N_10719);
nor U11074 (N_11074,N_10562,N_10569);
and U11075 (N_11075,N_10711,N_10877);
nand U11076 (N_11076,N_10159,N_10865);
or U11077 (N_11077,N_10666,N_10591);
and U11078 (N_11078,N_10669,N_10056);
and U11079 (N_11079,N_10744,N_10872);
xnor U11080 (N_11080,N_10161,N_10376);
or U11081 (N_11081,N_10303,N_10029);
or U11082 (N_11082,N_10813,N_10280);
and U11083 (N_11083,N_10597,N_10966);
and U11084 (N_11084,N_10404,N_10463);
nand U11085 (N_11085,N_10214,N_10776);
and U11086 (N_11086,N_10672,N_10445);
nand U11087 (N_11087,N_10567,N_10798);
xor U11088 (N_11088,N_10709,N_10829);
and U11089 (N_11089,N_10875,N_10757);
nand U11090 (N_11090,N_10483,N_10824);
or U11091 (N_11091,N_10082,N_10330);
or U11092 (N_11092,N_10940,N_10036);
or U11093 (N_11093,N_10906,N_10008);
or U11094 (N_11094,N_10763,N_10950);
or U11095 (N_11095,N_10733,N_10560);
nor U11096 (N_11096,N_10040,N_10706);
nor U11097 (N_11097,N_10718,N_10182);
nor U11098 (N_11098,N_10730,N_10498);
and U11099 (N_11099,N_10948,N_10681);
nand U11100 (N_11100,N_10031,N_10647);
nand U11101 (N_11101,N_10157,N_10178);
nand U11102 (N_11102,N_10344,N_10970);
nor U11103 (N_11103,N_10358,N_10081);
xnor U11104 (N_11104,N_10710,N_10137);
and U11105 (N_11105,N_10687,N_10292);
nor U11106 (N_11106,N_10957,N_10175);
and U11107 (N_11107,N_10519,N_10624);
and U11108 (N_11108,N_10742,N_10715);
nand U11109 (N_11109,N_10275,N_10985);
and U11110 (N_11110,N_10145,N_10633);
nor U11111 (N_11111,N_10231,N_10538);
and U11112 (N_11112,N_10536,N_10119);
and U11113 (N_11113,N_10440,N_10532);
nor U11114 (N_11114,N_10003,N_10171);
xor U11115 (N_11115,N_10041,N_10309);
nand U11116 (N_11116,N_10360,N_10786);
or U11117 (N_11117,N_10447,N_10566);
and U11118 (N_11118,N_10191,N_10457);
nor U11119 (N_11119,N_10166,N_10462);
nand U11120 (N_11120,N_10554,N_10874);
and U11121 (N_11121,N_10821,N_10100);
and U11122 (N_11122,N_10581,N_10690);
and U11123 (N_11123,N_10190,N_10839);
nand U11124 (N_11124,N_10055,N_10227);
xor U11125 (N_11125,N_10822,N_10076);
or U11126 (N_11126,N_10608,N_10010);
nor U11127 (N_11127,N_10499,N_10712);
or U11128 (N_11128,N_10832,N_10973);
nand U11129 (N_11129,N_10735,N_10495);
nand U11130 (N_11130,N_10936,N_10494);
and U11131 (N_11131,N_10748,N_10590);
and U11132 (N_11132,N_10308,N_10859);
and U11133 (N_11133,N_10521,N_10605);
nand U11134 (N_11134,N_10864,N_10306);
nor U11135 (N_11135,N_10508,N_10362);
xnor U11136 (N_11136,N_10071,N_10341);
or U11137 (N_11137,N_10431,N_10389);
nor U11138 (N_11138,N_10507,N_10571);
or U11139 (N_11139,N_10765,N_10354);
nand U11140 (N_11140,N_10585,N_10575);
or U11141 (N_11141,N_10305,N_10949);
nor U11142 (N_11142,N_10475,N_10593);
or U11143 (N_11143,N_10815,N_10628);
or U11144 (N_11144,N_10800,N_10623);
and U11145 (N_11145,N_10504,N_10760);
nand U11146 (N_11146,N_10952,N_10614);
nor U11147 (N_11147,N_10915,N_10085);
nand U11148 (N_11148,N_10000,N_10391);
and U11149 (N_11149,N_10325,N_10721);
nor U11150 (N_11150,N_10529,N_10541);
xor U11151 (N_11151,N_10203,N_10675);
or U11152 (N_11152,N_10991,N_10403);
and U11153 (N_11153,N_10651,N_10458);
nor U11154 (N_11154,N_10060,N_10226);
nor U11155 (N_11155,N_10382,N_10726);
or U11156 (N_11156,N_10032,N_10642);
nand U11157 (N_11157,N_10568,N_10916);
nor U11158 (N_11158,N_10602,N_10761);
nand U11159 (N_11159,N_10862,N_10048);
and U11160 (N_11160,N_10284,N_10580);
and U11161 (N_11161,N_10552,N_10393);
nand U11162 (N_11162,N_10871,N_10557);
and U11163 (N_11163,N_10563,N_10917);
nand U11164 (N_11164,N_10901,N_10170);
nand U11165 (N_11165,N_10319,N_10255);
nand U11166 (N_11166,N_10751,N_10790);
xnor U11167 (N_11167,N_10383,N_10935);
nor U11168 (N_11168,N_10063,N_10035);
nor U11169 (N_11169,N_10791,N_10181);
nor U11170 (N_11170,N_10204,N_10244);
or U11171 (N_11171,N_10782,N_10073);
nand U11172 (N_11172,N_10006,N_10959);
nand U11173 (N_11173,N_10732,N_10108);
or U11174 (N_11174,N_10080,N_10771);
nor U11175 (N_11175,N_10177,N_10264);
nor U11176 (N_11176,N_10551,N_10232);
or U11177 (N_11177,N_10599,N_10320);
and U11178 (N_11178,N_10198,N_10357);
xor U11179 (N_11179,N_10956,N_10331);
or U11180 (N_11180,N_10544,N_10479);
nand U11181 (N_11181,N_10924,N_10728);
nor U11182 (N_11182,N_10429,N_10466);
nand U11183 (N_11183,N_10828,N_10205);
or U11184 (N_11184,N_10117,N_10484);
and U11185 (N_11185,N_10631,N_10890);
nand U11186 (N_11186,N_10584,N_10564);
nor U11187 (N_11187,N_10896,N_10524);
or U11188 (N_11188,N_10643,N_10632);
nor U11189 (N_11189,N_10685,N_10435);
or U11190 (N_11190,N_10473,N_10128);
and U11191 (N_11191,N_10724,N_10703);
nand U11192 (N_11192,N_10367,N_10682);
and U11193 (N_11193,N_10064,N_10899);
nor U11194 (N_11194,N_10188,N_10372);
nor U11195 (N_11195,N_10767,N_10453);
and U11196 (N_11196,N_10356,N_10121);
and U11197 (N_11197,N_10678,N_10514);
xnor U11198 (N_11198,N_10530,N_10374);
nand U11199 (N_11199,N_10595,N_10752);
nor U11200 (N_11200,N_10967,N_10764);
or U11201 (N_11201,N_10015,N_10116);
nor U11202 (N_11202,N_10152,N_10990);
nor U11203 (N_11203,N_10847,N_10452);
or U11204 (N_11204,N_10299,N_10101);
or U11205 (N_11205,N_10753,N_10276);
nor U11206 (N_11206,N_10294,N_10148);
nand U11207 (N_11207,N_10572,N_10627);
or U11208 (N_11208,N_10207,N_10550);
nor U11209 (N_11209,N_10395,N_10009);
or U11210 (N_11210,N_10348,N_10511);
or U11211 (N_11211,N_10105,N_10799);
xor U11212 (N_11212,N_10897,N_10315);
nor U11213 (N_11213,N_10263,N_10515);
and U11214 (N_11214,N_10603,N_10069);
and U11215 (N_11215,N_10102,N_10045);
and U11216 (N_11216,N_10698,N_10424);
or U11217 (N_11217,N_10200,N_10225);
and U11218 (N_11218,N_10657,N_10285);
and U11219 (N_11219,N_10987,N_10257);
or U11220 (N_11220,N_10695,N_10378);
nor U11221 (N_11221,N_10547,N_10579);
xnor U11222 (N_11222,N_10594,N_10212);
or U11223 (N_11223,N_10891,N_10084);
and U11224 (N_11224,N_10363,N_10441);
nor U11225 (N_11225,N_10074,N_10038);
and U11226 (N_11226,N_10173,N_10456);
nor U11227 (N_11227,N_10149,N_10236);
nor U11228 (N_11228,N_10620,N_10674);
nand U11229 (N_11229,N_10845,N_10099);
nor U11230 (N_11230,N_10883,N_10988);
nor U11231 (N_11231,N_10196,N_10707);
and U11232 (N_11232,N_10072,N_10373);
and U11233 (N_11233,N_10012,N_10640);
nor U11234 (N_11234,N_10621,N_10201);
nand U11235 (N_11235,N_10037,N_10468);
nor U11236 (N_11236,N_10211,N_10638);
nor U11237 (N_11237,N_10774,N_10691);
or U11238 (N_11238,N_10039,N_10697);
nand U11239 (N_11239,N_10968,N_10664);
and U11240 (N_11240,N_10274,N_10876);
and U11241 (N_11241,N_10240,N_10827);
or U11242 (N_11242,N_10154,N_10731);
nand U11243 (N_11243,N_10164,N_10242);
or U11244 (N_11244,N_10298,N_10120);
and U11245 (N_11245,N_10779,N_10654);
nand U11246 (N_11246,N_10738,N_10954);
or U11247 (N_11247,N_10013,N_10381);
and U11248 (N_11248,N_10469,N_10688);
or U11249 (N_11249,N_10673,N_10720);
nor U11250 (N_11250,N_10464,N_10592);
and U11251 (N_11251,N_10737,N_10789);
nor U11252 (N_11252,N_10670,N_10676);
and U11253 (N_11253,N_10279,N_10364);
nor U11254 (N_11254,N_10696,N_10797);
xor U11255 (N_11255,N_10089,N_10411);
nand U11256 (N_11256,N_10729,N_10022);
and U11257 (N_11257,N_10151,N_10328);
or U11258 (N_11258,N_10481,N_10272);
and U11259 (N_11259,N_10951,N_10945);
nor U11260 (N_11260,N_10528,N_10020);
xnor U11261 (N_11261,N_10820,N_10850);
or U11262 (N_11262,N_10417,N_10863);
or U11263 (N_11263,N_10400,N_10768);
and U11264 (N_11264,N_10686,N_10256);
nand U11265 (N_11265,N_10808,N_10250);
or U11266 (N_11266,N_10539,N_10335);
xor U11267 (N_11267,N_10219,N_10518);
and U11268 (N_11268,N_10888,N_10488);
nor U11269 (N_11269,N_10088,N_10558);
or U11270 (N_11270,N_10313,N_10559);
nor U11271 (N_11271,N_10749,N_10542);
nor U11272 (N_11272,N_10977,N_10053);
nand U11273 (N_11273,N_10887,N_10144);
nor U11274 (N_11274,N_10296,N_10406);
xor U11275 (N_11275,N_10505,N_10833);
nand U11276 (N_11276,N_10693,N_10143);
and U11277 (N_11277,N_10206,N_10125);
nor U11278 (N_11278,N_10169,N_10834);
or U11279 (N_11279,N_10220,N_10996);
xor U11280 (N_11280,N_10911,N_10677);
and U11281 (N_11281,N_10909,N_10825);
or U11282 (N_11282,N_10014,N_10289);
xnor U11283 (N_11283,N_10366,N_10727);
and U11284 (N_11284,N_10933,N_10422);
xnor U11285 (N_11285,N_10816,N_10047);
and U11286 (N_11286,N_10634,N_10146);
and U11287 (N_11287,N_10365,N_10350);
or U11288 (N_11288,N_10482,N_10645);
and U11289 (N_11289,N_10881,N_10258);
nand U11290 (N_11290,N_10409,N_10830);
and U11291 (N_11291,N_10976,N_10024);
or U11292 (N_11292,N_10953,N_10455);
nand U11293 (N_11293,N_10734,N_10487);
and U11294 (N_11294,N_10241,N_10104);
xor U11295 (N_11295,N_10838,N_10016);
or U11296 (N_11296,N_10027,N_10185);
and U11297 (N_11297,N_10267,N_10322);
xor U11298 (N_11298,N_10772,N_10506);
nand U11299 (N_11299,N_10758,N_10437);
nor U11300 (N_11300,N_10921,N_10979);
xnor U11301 (N_11301,N_10692,N_10545);
nand U11302 (N_11302,N_10928,N_10637);
nand U11303 (N_11303,N_10460,N_10193);
nor U11304 (N_11304,N_10679,N_10394);
or U11305 (N_11305,N_10423,N_10927);
nor U11306 (N_11306,N_10172,N_10302);
and U11307 (N_11307,N_10972,N_10932);
or U11308 (N_11308,N_10223,N_10537);
xnor U11309 (N_11309,N_10754,N_10337);
nor U11310 (N_11310,N_10806,N_10489);
and U11311 (N_11311,N_10418,N_10746);
nand U11312 (N_11312,N_10221,N_10574);
nand U11313 (N_11313,N_10114,N_10333);
and U11314 (N_11314,N_10762,N_10336);
and U11315 (N_11315,N_10028,N_10873);
nand U11316 (N_11316,N_10926,N_10446);
nor U11317 (N_11317,N_10371,N_10249);
nand U11318 (N_11318,N_10338,N_10533);
nand U11319 (N_11319,N_10842,N_10208);
nand U11320 (N_11320,N_10043,N_10577);
nor U11321 (N_11321,N_10091,N_10270);
xnor U11322 (N_11322,N_10051,N_10370);
or U11323 (N_11323,N_10021,N_10421);
or U11324 (N_11324,N_10426,N_10176);
nand U11325 (N_11325,N_10803,N_10604);
and U11326 (N_11326,N_10609,N_10269);
and U11327 (N_11327,N_10412,N_10807);
and U11328 (N_11328,N_10318,N_10168);
nor U11329 (N_11329,N_10218,N_10766);
nor U11330 (N_11330,N_10998,N_10129);
nor U11331 (N_11331,N_10001,N_10167);
and U11332 (N_11332,N_10905,N_10958);
and U11333 (N_11333,N_10910,N_10110);
nor U11334 (N_11334,N_10809,N_10287);
and U11335 (N_11335,N_10785,N_10812);
or U11336 (N_11336,N_10377,N_10652);
and U11337 (N_11337,N_10653,N_10625);
or U11338 (N_11338,N_10846,N_10840);
nand U11339 (N_11339,N_10995,N_10549);
nor U11340 (N_11340,N_10407,N_10304);
nand U11341 (N_11341,N_10235,N_10778);
and U11342 (N_11342,N_10880,N_10914);
xnor U11343 (N_11343,N_10925,N_10399);
xor U11344 (N_11344,N_10601,N_10392);
nor U11345 (N_11345,N_10160,N_10610);
nor U11346 (N_11346,N_10034,N_10023);
or U11347 (N_11347,N_10713,N_10131);
nand U11348 (N_11348,N_10139,N_10290);
nor U11349 (N_11349,N_10345,N_10087);
and U11350 (N_11350,N_10955,N_10210);
or U11351 (N_11351,N_10359,N_10635);
nor U11352 (N_11352,N_10555,N_10369);
or U11353 (N_11353,N_10261,N_10405);
or U11354 (N_11354,N_10142,N_10823);
or U11355 (N_11355,N_10233,N_10750);
or U11356 (N_11356,N_10811,N_10092);
or U11357 (N_11357,N_10427,N_10213);
nand U11358 (N_11358,N_10900,N_10162);
xnor U11359 (N_11359,N_10098,N_10147);
nand U11360 (N_11360,N_10660,N_10075);
and U11361 (N_11361,N_10714,N_10964);
and U11362 (N_11362,N_10851,N_10723);
and U11363 (N_11363,N_10868,N_10184);
or U11364 (N_11364,N_10644,N_10756);
nand U11365 (N_11365,N_10273,N_10983);
nand U11366 (N_11366,N_10353,N_10540);
or U11367 (N_11367,N_10425,N_10415);
nand U11368 (N_11368,N_10894,N_10639);
nand U11369 (N_11369,N_10402,N_10316);
and U11370 (N_11370,N_10187,N_10646);
nand U11371 (N_11371,N_10326,N_10844);
or U11372 (N_11372,N_10093,N_10708);
xnor U11373 (N_11373,N_10814,N_10831);
nor U11374 (N_11374,N_10817,N_10517);
xor U11375 (N_11375,N_10512,N_10999);
nand U11376 (N_11376,N_10282,N_10449);
or U11377 (N_11377,N_10994,N_10459);
xor U11378 (N_11378,N_10049,N_10113);
nand U11379 (N_11379,N_10781,N_10317);
nand U11380 (N_11380,N_10238,N_10138);
or U11381 (N_11381,N_10130,N_10801);
nand U11382 (N_11382,N_10254,N_10078);
nor U11383 (N_11383,N_10243,N_10971);
and U11384 (N_11384,N_10658,N_10659);
nor U11385 (N_11385,N_10513,N_10583);
nand U11386 (N_11386,N_10153,N_10769);
and U11387 (N_11387,N_10115,N_10904);
nor U11388 (N_11388,N_10136,N_10339);
nor U11389 (N_11389,N_10224,N_10122);
nor U11390 (N_11390,N_10297,N_10026);
or U11391 (N_11391,N_10347,N_10135);
or U11392 (N_11392,N_10826,N_10410);
nand U11393 (N_11393,N_10094,N_10527);
and U11394 (N_11394,N_10312,N_10740);
nor U11395 (N_11395,N_10649,N_10655);
nor U11396 (N_11396,N_10112,N_10630);
nor U11397 (N_11397,N_10252,N_10434);
nand U11398 (N_11398,N_10663,N_10278);
nand U11399 (N_11399,N_10451,N_10854);
nor U11400 (N_11400,N_10615,N_10054);
nor U11401 (N_11401,N_10770,N_10189);
and U11402 (N_11402,N_10132,N_10268);
nand U11403 (N_11403,N_10939,N_10229);
or U11404 (N_11404,N_10461,N_10586);
nand U11405 (N_11405,N_10194,N_10548);
xnor U11406 (N_11406,N_10694,N_10661);
and U11407 (N_11407,N_10841,N_10668);
or U11408 (N_11408,N_10934,N_10902);
and U11409 (N_11409,N_10155,N_10052);
nand U11410 (N_11410,N_10701,N_10090);
nor U11411 (N_11411,N_10739,N_10502);
nand U11412 (N_11412,N_10974,N_10885);
or U11413 (N_11413,N_10126,N_10913);
and U11414 (N_11414,N_10736,N_10613);
xnor U11415 (N_11415,N_10648,N_10606);
nand U11416 (N_11416,N_10895,N_10030);
or U11417 (N_11417,N_10665,N_10650);
nand U11418 (N_11418,N_10745,N_10343);
nor U11419 (N_11419,N_10386,N_10490);
and U11420 (N_11420,N_10413,N_10903);
nor U11421 (N_11421,N_10918,N_10007);
xnor U11422 (N_11422,N_10127,N_10375);
nand U11423 (N_11423,N_10978,N_10332);
or U11424 (N_11424,N_10773,N_10183);
nor U11425 (N_11425,N_10981,N_10662);
and U11426 (N_11426,N_10819,N_10747);
and U11427 (N_11427,N_10199,N_10879);
nand U11428 (N_11428,N_10486,N_10283);
xnor U11429 (N_11429,N_10042,N_10044);
or U11430 (N_11430,N_10920,N_10396);
nor U11431 (N_11431,N_10025,N_10228);
xor U11432 (N_11432,N_10626,N_10059);
nor U11433 (N_11433,N_10416,N_10497);
nand U11434 (N_11434,N_10805,N_10465);
or U11435 (N_11435,N_10855,N_10033);
and U11436 (N_11436,N_10907,N_10222);
nor U11437 (N_11437,N_10011,N_10870);
or U11438 (N_11438,N_10420,N_10454);
nor U11439 (N_11439,N_10535,N_10963);
nand U11440 (N_11440,N_10795,N_10248);
xor U11441 (N_11441,N_10165,N_10783);
or U11442 (N_11442,N_10323,N_10565);
or U11443 (N_11443,N_10433,N_10852);
or U11444 (N_11444,N_10436,N_10355);
or U11445 (N_11445,N_10792,N_10600);
or U11446 (N_11446,N_10923,N_10578);
nand U11447 (N_11447,N_10607,N_10202);
or U11448 (N_11448,N_10671,N_10683);
nand U11449 (N_11449,N_10005,N_10140);
nand U11450 (N_11450,N_10329,N_10622);
or U11451 (N_11451,N_10186,N_10002);
and U11452 (N_11452,N_10111,N_10432);
or U11453 (N_11453,N_10941,N_10810);
xnor U11454 (N_11454,N_10546,N_10311);
or U11455 (N_11455,N_10629,N_10858);
nand U11456 (N_11456,N_10656,N_10018);
and U11457 (N_11457,N_10680,N_10251);
or U11458 (N_11458,N_10321,N_10017);
and U11459 (N_11459,N_10387,N_10300);
and U11460 (N_11460,N_10992,N_10262);
nor U11461 (N_11461,N_10174,N_10301);
xor U11462 (N_11462,N_10266,N_10478);
and U11463 (N_11463,N_10856,N_10442);
and U11464 (N_11464,N_10878,N_10209);
and U11465 (N_11465,N_10476,N_10796);
and U11466 (N_11466,N_10612,N_10340);
nand U11467 (N_11467,N_10237,N_10699);
nor U11468 (N_11468,N_10245,N_10961);
and U11469 (N_11469,N_10716,N_10230);
nand U11470 (N_11470,N_10561,N_10106);
xor U11471 (N_11471,N_10616,N_10501);
nand U11472 (N_11472,N_10050,N_10192);
or U11473 (N_11473,N_10295,N_10702);
or U11474 (N_11474,N_10743,N_10944);
and U11475 (N_11475,N_10993,N_10705);
nor U11476 (N_11476,N_10061,N_10641);
nor U11477 (N_11477,N_10947,N_10349);
nand U11478 (N_11478,N_10019,N_10700);
nand U11479 (N_11479,N_10500,N_10510);
or U11480 (N_11480,N_10398,N_10286);
nor U11481 (N_11481,N_10065,N_10984);
nand U11482 (N_11482,N_10197,N_10067);
and U11483 (N_11483,N_10496,N_10450);
or U11484 (N_11484,N_10975,N_10570);
or U11485 (N_11485,N_10818,N_10804);
nor U11486 (N_11486,N_10722,N_10086);
nor U11487 (N_11487,N_10576,N_10058);
xor U11488 (N_11488,N_10618,N_10163);
nor U11489 (N_11489,N_10004,N_10234);
nand U11490 (N_11490,N_10836,N_10288);
nand U11491 (N_11491,N_10704,N_10291);
or U11492 (N_11492,N_10379,N_10430);
or U11493 (N_11493,N_10390,N_10867);
nor U11494 (N_11494,N_10141,N_10522);
xor U11495 (N_11495,N_10253,N_10788);
or U11496 (N_11496,N_10247,N_10908);
xnor U11497 (N_11497,N_10414,N_10587);
or U11498 (N_11498,N_10929,N_10314);
and U11499 (N_11499,N_10777,N_10066);
xor U11500 (N_11500,N_10413,N_10802);
nand U11501 (N_11501,N_10574,N_10585);
xnor U11502 (N_11502,N_10188,N_10665);
nor U11503 (N_11503,N_10967,N_10573);
nor U11504 (N_11504,N_10930,N_10939);
or U11505 (N_11505,N_10099,N_10518);
nor U11506 (N_11506,N_10091,N_10958);
nor U11507 (N_11507,N_10291,N_10055);
or U11508 (N_11508,N_10101,N_10718);
or U11509 (N_11509,N_10068,N_10709);
and U11510 (N_11510,N_10802,N_10013);
xor U11511 (N_11511,N_10356,N_10506);
and U11512 (N_11512,N_10981,N_10715);
nor U11513 (N_11513,N_10619,N_10473);
xor U11514 (N_11514,N_10992,N_10903);
nor U11515 (N_11515,N_10278,N_10428);
and U11516 (N_11516,N_10363,N_10974);
or U11517 (N_11517,N_10233,N_10817);
nand U11518 (N_11518,N_10568,N_10277);
and U11519 (N_11519,N_10106,N_10045);
nor U11520 (N_11520,N_10913,N_10907);
nor U11521 (N_11521,N_10040,N_10220);
or U11522 (N_11522,N_10998,N_10020);
nor U11523 (N_11523,N_10009,N_10630);
and U11524 (N_11524,N_10663,N_10470);
nand U11525 (N_11525,N_10214,N_10377);
xnor U11526 (N_11526,N_10791,N_10034);
nand U11527 (N_11527,N_10448,N_10261);
nand U11528 (N_11528,N_10568,N_10820);
or U11529 (N_11529,N_10994,N_10752);
nor U11530 (N_11530,N_10472,N_10538);
and U11531 (N_11531,N_10794,N_10643);
or U11532 (N_11532,N_10873,N_10998);
nand U11533 (N_11533,N_10449,N_10656);
or U11534 (N_11534,N_10435,N_10509);
and U11535 (N_11535,N_10090,N_10255);
nand U11536 (N_11536,N_10782,N_10061);
or U11537 (N_11537,N_10285,N_10699);
and U11538 (N_11538,N_10547,N_10542);
and U11539 (N_11539,N_10434,N_10187);
or U11540 (N_11540,N_10713,N_10374);
nand U11541 (N_11541,N_10997,N_10724);
xnor U11542 (N_11542,N_10962,N_10451);
nand U11543 (N_11543,N_10945,N_10177);
nand U11544 (N_11544,N_10960,N_10812);
or U11545 (N_11545,N_10643,N_10333);
nor U11546 (N_11546,N_10336,N_10330);
nand U11547 (N_11547,N_10431,N_10271);
and U11548 (N_11548,N_10931,N_10669);
and U11549 (N_11549,N_10822,N_10090);
nor U11550 (N_11550,N_10418,N_10966);
nor U11551 (N_11551,N_10023,N_10401);
and U11552 (N_11552,N_10072,N_10609);
and U11553 (N_11553,N_10953,N_10479);
nor U11554 (N_11554,N_10409,N_10990);
or U11555 (N_11555,N_10170,N_10775);
or U11556 (N_11556,N_10252,N_10657);
xor U11557 (N_11557,N_10039,N_10931);
or U11558 (N_11558,N_10265,N_10762);
nor U11559 (N_11559,N_10058,N_10904);
nor U11560 (N_11560,N_10784,N_10586);
or U11561 (N_11561,N_10339,N_10352);
and U11562 (N_11562,N_10034,N_10698);
or U11563 (N_11563,N_10928,N_10251);
nor U11564 (N_11564,N_10339,N_10763);
or U11565 (N_11565,N_10194,N_10619);
or U11566 (N_11566,N_10030,N_10955);
and U11567 (N_11567,N_10784,N_10472);
xnor U11568 (N_11568,N_10603,N_10537);
or U11569 (N_11569,N_10651,N_10529);
xor U11570 (N_11570,N_10176,N_10372);
nand U11571 (N_11571,N_10043,N_10721);
xor U11572 (N_11572,N_10827,N_10274);
and U11573 (N_11573,N_10664,N_10972);
or U11574 (N_11574,N_10221,N_10771);
xor U11575 (N_11575,N_10069,N_10018);
or U11576 (N_11576,N_10074,N_10691);
or U11577 (N_11577,N_10342,N_10238);
and U11578 (N_11578,N_10943,N_10710);
or U11579 (N_11579,N_10503,N_10722);
nand U11580 (N_11580,N_10715,N_10676);
and U11581 (N_11581,N_10019,N_10028);
nor U11582 (N_11582,N_10392,N_10552);
nand U11583 (N_11583,N_10385,N_10623);
or U11584 (N_11584,N_10970,N_10243);
and U11585 (N_11585,N_10436,N_10897);
and U11586 (N_11586,N_10469,N_10838);
nor U11587 (N_11587,N_10655,N_10366);
nor U11588 (N_11588,N_10516,N_10210);
and U11589 (N_11589,N_10667,N_10020);
nor U11590 (N_11590,N_10700,N_10973);
nand U11591 (N_11591,N_10965,N_10186);
nor U11592 (N_11592,N_10867,N_10041);
nor U11593 (N_11593,N_10687,N_10507);
or U11594 (N_11594,N_10290,N_10724);
nor U11595 (N_11595,N_10948,N_10384);
and U11596 (N_11596,N_10973,N_10969);
xor U11597 (N_11597,N_10880,N_10222);
or U11598 (N_11598,N_10540,N_10903);
nand U11599 (N_11599,N_10173,N_10519);
nor U11600 (N_11600,N_10341,N_10369);
and U11601 (N_11601,N_10383,N_10602);
nor U11602 (N_11602,N_10167,N_10685);
xor U11603 (N_11603,N_10983,N_10405);
nor U11604 (N_11604,N_10883,N_10176);
and U11605 (N_11605,N_10488,N_10546);
or U11606 (N_11606,N_10972,N_10492);
and U11607 (N_11607,N_10155,N_10510);
nor U11608 (N_11608,N_10023,N_10935);
or U11609 (N_11609,N_10083,N_10024);
and U11610 (N_11610,N_10312,N_10016);
nand U11611 (N_11611,N_10853,N_10404);
nor U11612 (N_11612,N_10824,N_10321);
and U11613 (N_11613,N_10553,N_10208);
nor U11614 (N_11614,N_10637,N_10138);
nand U11615 (N_11615,N_10070,N_10282);
nand U11616 (N_11616,N_10510,N_10711);
and U11617 (N_11617,N_10645,N_10005);
and U11618 (N_11618,N_10165,N_10753);
or U11619 (N_11619,N_10123,N_10147);
and U11620 (N_11620,N_10541,N_10722);
and U11621 (N_11621,N_10714,N_10340);
xor U11622 (N_11622,N_10496,N_10615);
and U11623 (N_11623,N_10169,N_10203);
or U11624 (N_11624,N_10204,N_10224);
and U11625 (N_11625,N_10613,N_10851);
nand U11626 (N_11626,N_10412,N_10282);
or U11627 (N_11627,N_10156,N_10368);
or U11628 (N_11628,N_10016,N_10759);
nor U11629 (N_11629,N_10860,N_10505);
or U11630 (N_11630,N_10235,N_10813);
nand U11631 (N_11631,N_10260,N_10880);
nor U11632 (N_11632,N_10537,N_10810);
and U11633 (N_11633,N_10636,N_10049);
nor U11634 (N_11634,N_10089,N_10645);
and U11635 (N_11635,N_10190,N_10710);
or U11636 (N_11636,N_10195,N_10450);
nor U11637 (N_11637,N_10737,N_10093);
nor U11638 (N_11638,N_10783,N_10260);
nor U11639 (N_11639,N_10988,N_10717);
and U11640 (N_11640,N_10324,N_10985);
nor U11641 (N_11641,N_10718,N_10989);
xor U11642 (N_11642,N_10470,N_10197);
nor U11643 (N_11643,N_10911,N_10233);
or U11644 (N_11644,N_10502,N_10563);
nor U11645 (N_11645,N_10125,N_10751);
and U11646 (N_11646,N_10360,N_10173);
nor U11647 (N_11647,N_10452,N_10607);
nor U11648 (N_11648,N_10822,N_10577);
nor U11649 (N_11649,N_10984,N_10381);
nand U11650 (N_11650,N_10213,N_10368);
nand U11651 (N_11651,N_10961,N_10764);
or U11652 (N_11652,N_10228,N_10799);
or U11653 (N_11653,N_10796,N_10687);
and U11654 (N_11654,N_10923,N_10604);
or U11655 (N_11655,N_10221,N_10753);
nor U11656 (N_11656,N_10218,N_10337);
nor U11657 (N_11657,N_10804,N_10578);
xor U11658 (N_11658,N_10598,N_10555);
nor U11659 (N_11659,N_10045,N_10757);
nand U11660 (N_11660,N_10186,N_10500);
and U11661 (N_11661,N_10321,N_10514);
xnor U11662 (N_11662,N_10873,N_10634);
nor U11663 (N_11663,N_10640,N_10645);
or U11664 (N_11664,N_10411,N_10073);
nor U11665 (N_11665,N_10995,N_10111);
nor U11666 (N_11666,N_10549,N_10488);
nor U11667 (N_11667,N_10097,N_10322);
nand U11668 (N_11668,N_10852,N_10904);
and U11669 (N_11669,N_10071,N_10124);
nand U11670 (N_11670,N_10104,N_10722);
and U11671 (N_11671,N_10634,N_10446);
nor U11672 (N_11672,N_10780,N_10551);
nor U11673 (N_11673,N_10298,N_10752);
nand U11674 (N_11674,N_10582,N_10161);
nor U11675 (N_11675,N_10706,N_10068);
or U11676 (N_11676,N_10252,N_10255);
or U11677 (N_11677,N_10412,N_10327);
or U11678 (N_11678,N_10521,N_10451);
nor U11679 (N_11679,N_10477,N_10041);
or U11680 (N_11680,N_10329,N_10184);
nand U11681 (N_11681,N_10897,N_10959);
and U11682 (N_11682,N_10173,N_10777);
nor U11683 (N_11683,N_10230,N_10508);
xor U11684 (N_11684,N_10892,N_10046);
or U11685 (N_11685,N_10765,N_10934);
nand U11686 (N_11686,N_10359,N_10747);
or U11687 (N_11687,N_10399,N_10984);
nor U11688 (N_11688,N_10964,N_10136);
nor U11689 (N_11689,N_10967,N_10086);
xnor U11690 (N_11690,N_10454,N_10226);
and U11691 (N_11691,N_10344,N_10888);
xnor U11692 (N_11692,N_10955,N_10501);
nor U11693 (N_11693,N_10359,N_10935);
nand U11694 (N_11694,N_10227,N_10980);
nor U11695 (N_11695,N_10505,N_10016);
or U11696 (N_11696,N_10834,N_10242);
or U11697 (N_11697,N_10522,N_10471);
nor U11698 (N_11698,N_10124,N_10608);
or U11699 (N_11699,N_10103,N_10057);
nand U11700 (N_11700,N_10531,N_10791);
nor U11701 (N_11701,N_10808,N_10309);
nand U11702 (N_11702,N_10698,N_10233);
nand U11703 (N_11703,N_10282,N_10340);
nor U11704 (N_11704,N_10514,N_10242);
and U11705 (N_11705,N_10843,N_10441);
and U11706 (N_11706,N_10701,N_10945);
or U11707 (N_11707,N_10717,N_10562);
nand U11708 (N_11708,N_10918,N_10135);
or U11709 (N_11709,N_10337,N_10455);
or U11710 (N_11710,N_10126,N_10129);
nand U11711 (N_11711,N_10677,N_10327);
or U11712 (N_11712,N_10255,N_10699);
xnor U11713 (N_11713,N_10682,N_10375);
nor U11714 (N_11714,N_10547,N_10119);
nor U11715 (N_11715,N_10694,N_10466);
nand U11716 (N_11716,N_10874,N_10279);
and U11717 (N_11717,N_10927,N_10477);
and U11718 (N_11718,N_10197,N_10035);
nand U11719 (N_11719,N_10185,N_10988);
or U11720 (N_11720,N_10503,N_10328);
or U11721 (N_11721,N_10182,N_10821);
nand U11722 (N_11722,N_10251,N_10334);
nor U11723 (N_11723,N_10336,N_10539);
xor U11724 (N_11724,N_10852,N_10674);
and U11725 (N_11725,N_10881,N_10351);
or U11726 (N_11726,N_10551,N_10785);
or U11727 (N_11727,N_10733,N_10537);
or U11728 (N_11728,N_10383,N_10125);
and U11729 (N_11729,N_10359,N_10503);
and U11730 (N_11730,N_10835,N_10244);
or U11731 (N_11731,N_10589,N_10221);
nor U11732 (N_11732,N_10552,N_10205);
and U11733 (N_11733,N_10335,N_10659);
nand U11734 (N_11734,N_10675,N_10224);
xnor U11735 (N_11735,N_10183,N_10628);
nor U11736 (N_11736,N_10175,N_10196);
nor U11737 (N_11737,N_10626,N_10435);
and U11738 (N_11738,N_10342,N_10113);
and U11739 (N_11739,N_10468,N_10247);
nor U11740 (N_11740,N_10298,N_10816);
or U11741 (N_11741,N_10693,N_10402);
nand U11742 (N_11742,N_10374,N_10027);
xor U11743 (N_11743,N_10164,N_10670);
nand U11744 (N_11744,N_10354,N_10704);
nor U11745 (N_11745,N_10341,N_10303);
or U11746 (N_11746,N_10863,N_10634);
xnor U11747 (N_11747,N_10091,N_10329);
nor U11748 (N_11748,N_10726,N_10498);
xor U11749 (N_11749,N_10052,N_10185);
nand U11750 (N_11750,N_10008,N_10994);
or U11751 (N_11751,N_10820,N_10106);
or U11752 (N_11752,N_10947,N_10231);
and U11753 (N_11753,N_10413,N_10480);
and U11754 (N_11754,N_10548,N_10274);
and U11755 (N_11755,N_10729,N_10923);
nand U11756 (N_11756,N_10812,N_10863);
and U11757 (N_11757,N_10269,N_10479);
nand U11758 (N_11758,N_10507,N_10452);
or U11759 (N_11759,N_10908,N_10835);
and U11760 (N_11760,N_10549,N_10524);
and U11761 (N_11761,N_10365,N_10457);
and U11762 (N_11762,N_10908,N_10243);
nand U11763 (N_11763,N_10797,N_10852);
xor U11764 (N_11764,N_10832,N_10390);
and U11765 (N_11765,N_10671,N_10732);
nor U11766 (N_11766,N_10655,N_10149);
nor U11767 (N_11767,N_10415,N_10387);
nor U11768 (N_11768,N_10101,N_10758);
or U11769 (N_11769,N_10316,N_10876);
nand U11770 (N_11770,N_10323,N_10110);
xnor U11771 (N_11771,N_10191,N_10526);
nor U11772 (N_11772,N_10509,N_10184);
nor U11773 (N_11773,N_10947,N_10733);
nor U11774 (N_11774,N_10114,N_10558);
and U11775 (N_11775,N_10875,N_10161);
or U11776 (N_11776,N_10825,N_10109);
nor U11777 (N_11777,N_10037,N_10236);
and U11778 (N_11778,N_10505,N_10710);
or U11779 (N_11779,N_10098,N_10370);
and U11780 (N_11780,N_10259,N_10586);
nor U11781 (N_11781,N_10878,N_10339);
and U11782 (N_11782,N_10752,N_10103);
nor U11783 (N_11783,N_10635,N_10809);
xnor U11784 (N_11784,N_10747,N_10595);
nand U11785 (N_11785,N_10819,N_10961);
and U11786 (N_11786,N_10985,N_10194);
nand U11787 (N_11787,N_10700,N_10715);
or U11788 (N_11788,N_10984,N_10406);
nor U11789 (N_11789,N_10287,N_10828);
nand U11790 (N_11790,N_10913,N_10745);
xnor U11791 (N_11791,N_10608,N_10462);
or U11792 (N_11792,N_10148,N_10838);
or U11793 (N_11793,N_10326,N_10686);
or U11794 (N_11794,N_10806,N_10436);
and U11795 (N_11795,N_10831,N_10493);
nor U11796 (N_11796,N_10949,N_10433);
nor U11797 (N_11797,N_10981,N_10535);
nor U11798 (N_11798,N_10405,N_10356);
nand U11799 (N_11799,N_10987,N_10541);
nor U11800 (N_11800,N_10206,N_10655);
or U11801 (N_11801,N_10213,N_10016);
or U11802 (N_11802,N_10412,N_10512);
or U11803 (N_11803,N_10126,N_10396);
or U11804 (N_11804,N_10766,N_10376);
or U11805 (N_11805,N_10762,N_10125);
nand U11806 (N_11806,N_10058,N_10003);
nor U11807 (N_11807,N_10744,N_10580);
or U11808 (N_11808,N_10943,N_10933);
nor U11809 (N_11809,N_10303,N_10883);
nor U11810 (N_11810,N_10580,N_10931);
or U11811 (N_11811,N_10015,N_10297);
and U11812 (N_11812,N_10907,N_10901);
nand U11813 (N_11813,N_10301,N_10699);
nor U11814 (N_11814,N_10630,N_10223);
and U11815 (N_11815,N_10636,N_10130);
nor U11816 (N_11816,N_10001,N_10157);
nand U11817 (N_11817,N_10351,N_10883);
nor U11818 (N_11818,N_10388,N_10438);
xor U11819 (N_11819,N_10076,N_10519);
nand U11820 (N_11820,N_10453,N_10601);
or U11821 (N_11821,N_10067,N_10921);
or U11822 (N_11822,N_10369,N_10412);
nand U11823 (N_11823,N_10335,N_10826);
or U11824 (N_11824,N_10777,N_10054);
and U11825 (N_11825,N_10034,N_10676);
nand U11826 (N_11826,N_10377,N_10799);
or U11827 (N_11827,N_10170,N_10841);
and U11828 (N_11828,N_10623,N_10238);
or U11829 (N_11829,N_10446,N_10381);
and U11830 (N_11830,N_10300,N_10199);
nand U11831 (N_11831,N_10068,N_10315);
xor U11832 (N_11832,N_10304,N_10259);
nand U11833 (N_11833,N_10099,N_10407);
and U11834 (N_11834,N_10163,N_10280);
nor U11835 (N_11835,N_10529,N_10776);
nand U11836 (N_11836,N_10300,N_10379);
nor U11837 (N_11837,N_10320,N_10679);
and U11838 (N_11838,N_10557,N_10054);
or U11839 (N_11839,N_10225,N_10540);
and U11840 (N_11840,N_10054,N_10788);
nor U11841 (N_11841,N_10975,N_10206);
nor U11842 (N_11842,N_10288,N_10313);
and U11843 (N_11843,N_10123,N_10378);
nand U11844 (N_11844,N_10709,N_10592);
nand U11845 (N_11845,N_10734,N_10414);
or U11846 (N_11846,N_10311,N_10748);
xnor U11847 (N_11847,N_10435,N_10691);
and U11848 (N_11848,N_10066,N_10590);
nand U11849 (N_11849,N_10498,N_10359);
nand U11850 (N_11850,N_10078,N_10762);
or U11851 (N_11851,N_10212,N_10823);
nand U11852 (N_11852,N_10699,N_10307);
nor U11853 (N_11853,N_10494,N_10006);
or U11854 (N_11854,N_10284,N_10764);
and U11855 (N_11855,N_10253,N_10549);
and U11856 (N_11856,N_10368,N_10878);
or U11857 (N_11857,N_10359,N_10313);
nand U11858 (N_11858,N_10394,N_10122);
or U11859 (N_11859,N_10119,N_10418);
or U11860 (N_11860,N_10464,N_10905);
nor U11861 (N_11861,N_10379,N_10449);
nor U11862 (N_11862,N_10507,N_10175);
xnor U11863 (N_11863,N_10887,N_10208);
nand U11864 (N_11864,N_10637,N_10099);
xor U11865 (N_11865,N_10083,N_10649);
nor U11866 (N_11866,N_10840,N_10823);
or U11867 (N_11867,N_10979,N_10355);
and U11868 (N_11868,N_10892,N_10163);
nor U11869 (N_11869,N_10410,N_10489);
nand U11870 (N_11870,N_10709,N_10746);
or U11871 (N_11871,N_10276,N_10024);
and U11872 (N_11872,N_10649,N_10340);
nor U11873 (N_11873,N_10083,N_10739);
or U11874 (N_11874,N_10929,N_10432);
nand U11875 (N_11875,N_10922,N_10051);
nor U11876 (N_11876,N_10952,N_10376);
xor U11877 (N_11877,N_10360,N_10253);
nand U11878 (N_11878,N_10263,N_10137);
nand U11879 (N_11879,N_10817,N_10815);
nor U11880 (N_11880,N_10530,N_10556);
or U11881 (N_11881,N_10256,N_10360);
nand U11882 (N_11882,N_10021,N_10772);
nand U11883 (N_11883,N_10204,N_10337);
or U11884 (N_11884,N_10869,N_10150);
or U11885 (N_11885,N_10575,N_10795);
nor U11886 (N_11886,N_10817,N_10306);
and U11887 (N_11887,N_10021,N_10387);
nand U11888 (N_11888,N_10629,N_10527);
nor U11889 (N_11889,N_10208,N_10413);
nand U11890 (N_11890,N_10794,N_10862);
xor U11891 (N_11891,N_10248,N_10989);
and U11892 (N_11892,N_10493,N_10311);
and U11893 (N_11893,N_10764,N_10309);
and U11894 (N_11894,N_10404,N_10222);
or U11895 (N_11895,N_10314,N_10920);
or U11896 (N_11896,N_10542,N_10043);
nor U11897 (N_11897,N_10521,N_10374);
nand U11898 (N_11898,N_10977,N_10224);
and U11899 (N_11899,N_10482,N_10939);
and U11900 (N_11900,N_10144,N_10106);
nand U11901 (N_11901,N_10551,N_10248);
nand U11902 (N_11902,N_10228,N_10311);
and U11903 (N_11903,N_10176,N_10192);
nor U11904 (N_11904,N_10860,N_10635);
and U11905 (N_11905,N_10108,N_10418);
nand U11906 (N_11906,N_10548,N_10022);
xor U11907 (N_11907,N_10370,N_10661);
nand U11908 (N_11908,N_10454,N_10895);
nor U11909 (N_11909,N_10713,N_10757);
xor U11910 (N_11910,N_10390,N_10720);
nand U11911 (N_11911,N_10890,N_10585);
nor U11912 (N_11912,N_10959,N_10745);
and U11913 (N_11913,N_10219,N_10391);
nand U11914 (N_11914,N_10515,N_10281);
nand U11915 (N_11915,N_10632,N_10336);
and U11916 (N_11916,N_10078,N_10170);
nor U11917 (N_11917,N_10858,N_10437);
nor U11918 (N_11918,N_10443,N_10743);
nand U11919 (N_11919,N_10049,N_10411);
and U11920 (N_11920,N_10335,N_10294);
or U11921 (N_11921,N_10005,N_10042);
and U11922 (N_11922,N_10666,N_10413);
nand U11923 (N_11923,N_10204,N_10550);
and U11924 (N_11924,N_10182,N_10998);
nor U11925 (N_11925,N_10485,N_10053);
or U11926 (N_11926,N_10308,N_10675);
and U11927 (N_11927,N_10427,N_10718);
xor U11928 (N_11928,N_10910,N_10533);
nand U11929 (N_11929,N_10435,N_10361);
or U11930 (N_11930,N_10108,N_10376);
xor U11931 (N_11931,N_10149,N_10775);
and U11932 (N_11932,N_10966,N_10538);
and U11933 (N_11933,N_10798,N_10835);
and U11934 (N_11934,N_10363,N_10409);
nor U11935 (N_11935,N_10272,N_10915);
nand U11936 (N_11936,N_10448,N_10081);
nor U11937 (N_11937,N_10351,N_10938);
nand U11938 (N_11938,N_10577,N_10320);
and U11939 (N_11939,N_10082,N_10475);
and U11940 (N_11940,N_10681,N_10649);
and U11941 (N_11941,N_10067,N_10068);
and U11942 (N_11942,N_10150,N_10977);
or U11943 (N_11943,N_10560,N_10428);
xor U11944 (N_11944,N_10476,N_10121);
nor U11945 (N_11945,N_10247,N_10579);
nand U11946 (N_11946,N_10171,N_10014);
nor U11947 (N_11947,N_10514,N_10260);
or U11948 (N_11948,N_10038,N_10071);
xnor U11949 (N_11949,N_10100,N_10022);
nand U11950 (N_11950,N_10851,N_10429);
or U11951 (N_11951,N_10566,N_10058);
and U11952 (N_11952,N_10140,N_10319);
nand U11953 (N_11953,N_10296,N_10926);
nor U11954 (N_11954,N_10601,N_10765);
or U11955 (N_11955,N_10767,N_10871);
nor U11956 (N_11956,N_10469,N_10713);
and U11957 (N_11957,N_10354,N_10690);
nand U11958 (N_11958,N_10391,N_10469);
nor U11959 (N_11959,N_10044,N_10715);
or U11960 (N_11960,N_10503,N_10423);
nand U11961 (N_11961,N_10993,N_10679);
nand U11962 (N_11962,N_10099,N_10134);
nand U11963 (N_11963,N_10039,N_10005);
and U11964 (N_11964,N_10040,N_10913);
nor U11965 (N_11965,N_10061,N_10712);
or U11966 (N_11966,N_10211,N_10857);
or U11967 (N_11967,N_10543,N_10882);
nand U11968 (N_11968,N_10733,N_10357);
nor U11969 (N_11969,N_10677,N_10240);
nand U11970 (N_11970,N_10916,N_10982);
nor U11971 (N_11971,N_10463,N_10771);
and U11972 (N_11972,N_10529,N_10040);
or U11973 (N_11973,N_10737,N_10288);
nand U11974 (N_11974,N_10486,N_10828);
nand U11975 (N_11975,N_10896,N_10051);
nand U11976 (N_11976,N_10015,N_10775);
or U11977 (N_11977,N_10180,N_10309);
nand U11978 (N_11978,N_10432,N_10247);
or U11979 (N_11979,N_10288,N_10730);
and U11980 (N_11980,N_10175,N_10071);
and U11981 (N_11981,N_10951,N_10775);
nand U11982 (N_11982,N_10178,N_10302);
and U11983 (N_11983,N_10580,N_10574);
and U11984 (N_11984,N_10691,N_10405);
and U11985 (N_11985,N_10078,N_10169);
nand U11986 (N_11986,N_10340,N_10907);
nand U11987 (N_11987,N_10021,N_10426);
or U11988 (N_11988,N_10682,N_10566);
nand U11989 (N_11989,N_10584,N_10265);
nand U11990 (N_11990,N_10662,N_10103);
or U11991 (N_11991,N_10665,N_10558);
or U11992 (N_11992,N_10596,N_10527);
or U11993 (N_11993,N_10769,N_10981);
nor U11994 (N_11994,N_10883,N_10462);
nor U11995 (N_11995,N_10782,N_10075);
nand U11996 (N_11996,N_10049,N_10728);
and U11997 (N_11997,N_10946,N_10588);
nand U11998 (N_11998,N_10344,N_10864);
nand U11999 (N_11999,N_10873,N_10973);
and U12000 (N_12000,N_11418,N_11784);
nor U12001 (N_12001,N_11246,N_11605);
nor U12002 (N_12002,N_11009,N_11151);
xor U12003 (N_12003,N_11412,N_11919);
or U12004 (N_12004,N_11134,N_11245);
and U12005 (N_12005,N_11207,N_11724);
or U12006 (N_12006,N_11376,N_11046);
nor U12007 (N_12007,N_11800,N_11978);
and U12008 (N_12008,N_11008,N_11045);
or U12009 (N_12009,N_11544,N_11071);
or U12010 (N_12010,N_11692,N_11402);
or U12011 (N_12011,N_11860,N_11439);
and U12012 (N_12012,N_11503,N_11972);
and U12013 (N_12013,N_11483,N_11723);
or U12014 (N_12014,N_11881,N_11212);
and U12015 (N_12015,N_11489,N_11379);
nand U12016 (N_12016,N_11443,N_11598);
nor U12017 (N_12017,N_11691,N_11948);
xor U12018 (N_12018,N_11781,N_11345);
xor U12019 (N_12019,N_11844,N_11714);
nor U12020 (N_12020,N_11380,N_11421);
xor U12021 (N_12021,N_11417,N_11786);
and U12022 (N_12022,N_11119,N_11330);
and U12023 (N_12023,N_11419,N_11508);
and U12024 (N_12024,N_11658,N_11655);
xor U12025 (N_12025,N_11185,N_11387);
xor U12026 (N_12026,N_11196,N_11166);
or U12027 (N_12027,N_11879,N_11539);
xnor U12028 (N_12028,N_11877,N_11707);
or U12029 (N_12029,N_11610,N_11057);
nand U12030 (N_12030,N_11203,N_11636);
and U12031 (N_12031,N_11855,N_11322);
nor U12032 (N_12032,N_11302,N_11889);
or U12033 (N_12033,N_11351,N_11080);
and U12034 (N_12034,N_11159,N_11484);
or U12035 (N_12035,N_11911,N_11805);
and U12036 (N_12036,N_11609,N_11319);
or U12037 (N_12037,N_11431,N_11981);
nand U12038 (N_12038,N_11210,N_11390);
and U12039 (N_12039,N_11792,N_11353);
or U12040 (N_12040,N_11704,N_11482);
nor U12041 (N_12041,N_11359,N_11975);
nor U12042 (N_12042,N_11928,N_11654);
nor U12043 (N_12043,N_11006,N_11337);
nor U12044 (N_12044,N_11635,N_11278);
nand U12045 (N_12045,N_11634,N_11509);
nor U12046 (N_12046,N_11593,N_11410);
or U12047 (N_12047,N_11957,N_11361);
nor U12048 (N_12048,N_11478,N_11661);
nand U12049 (N_12049,N_11557,N_11721);
nand U12050 (N_12050,N_11644,N_11355);
or U12051 (N_12051,N_11317,N_11020);
and U12052 (N_12052,N_11730,N_11682);
nor U12053 (N_12053,N_11998,N_11833);
or U12054 (N_12054,N_11996,N_11727);
or U12055 (N_12055,N_11522,N_11687);
and U12056 (N_12056,N_11592,N_11165);
nor U12057 (N_12057,N_11914,N_11548);
and U12058 (N_12058,N_11876,N_11922);
and U12059 (N_12059,N_11095,N_11393);
and U12060 (N_12060,N_11872,N_11845);
nand U12061 (N_12061,N_11577,N_11912);
or U12062 (N_12062,N_11829,N_11125);
xor U12063 (N_12063,N_11683,N_11149);
or U12064 (N_12064,N_11686,N_11899);
nand U12065 (N_12065,N_11167,N_11816);
nor U12066 (N_12066,N_11329,N_11672);
xnor U12067 (N_12067,N_11910,N_11106);
nand U12068 (N_12068,N_11445,N_11733);
xor U12069 (N_12069,N_11316,N_11191);
nand U12070 (N_12070,N_11437,N_11334);
nand U12071 (N_12071,N_11465,N_11255);
nand U12072 (N_12072,N_11247,N_11959);
nor U12073 (N_12073,N_11513,N_11409);
nand U12074 (N_12074,N_11047,N_11012);
nand U12075 (N_12075,N_11271,N_11357);
nand U12076 (N_12076,N_11296,N_11123);
or U12077 (N_12077,N_11251,N_11115);
or U12078 (N_12078,N_11819,N_11164);
nand U12079 (N_12079,N_11101,N_11563);
nand U12080 (N_12080,N_11902,N_11462);
nor U12081 (N_12081,N_11734,N_11772);
nor U12082 (N_12082,N_11798,N_11823);
nand U12083 (N_12083,N_11146,N_11738);
nand U12084 (N_12084,N_11239,N_11973);
or U12085 (N_12085,N_11260,N_11556);
and U12086 (N_12086,N_11017,N_11270);
nor U12087 (N_12087,N_11339,N_11620);
nand U12088 (N_12088,N_11433,N_11003);
and U12089 (N_12089,N_11731,N_11524);
nand U12090 (N_12090,N_11931,N_11938);
and U12091 (N_12091,N_11184,N_11510);
nand U12092 (N_12092,N_11836,N_11237);
nor U12093 (N_12093,N_11920,N_11033);
nand U12094 (N_12094,N_11026,N_11214);
nand U12095 (N_12095,N_11621,N_11452);
or U12096 (N_12096,N_11340,N_11256);
nand U12097 (N_12097,N_11552,N_11386);
xnor U12098 (N_12098,N_11369,N_11954);
nand U12099 (N_12099,N_11362,N_11348);
or U12100 (N_12100,N_11579,N_11093);
nor U12101 (N_12101,N_11281,N_11516);
xnor U12102 (N_12102,N_11657,N_11092);
or U12103 (N_12103,N_11710,N_11016);
and U12104 (N_12104,N_11015,N_11314);
nor U12105 (N_12105,N_11793,N_11991);
and U12106 (N_12106,N_11666,N_11751);
and U12107 (N_12107,N_11542,N_11061);
or U12108 (N_12108,N_11013,N_11066);
nor U12109 (N_12109,N_11477,N_11964);
and U12110 (N_12110,N_11673,N_11364);
nand U12111 (N_12111,N_11486,N_11535);
nand U12112 (N_12112,N_11158,N_11933);
xor U12113 (N_12113,N_11985,N_11514);
xor U12114 (N_12114,N_11618,N_11269);
or U12115 (N_12115,N_11019,N_11900);
and U12116 (N_12116,N_11588,N_11617);
or U12117 (N_12117,N_11148,N_11089);
nand U12118 (N_12118,N_11528,N_11377);
nor U12119 (N_12119,N_11285,N_11648);
or U12120 (N_12120,N_11760,N_11541);
and U12121 (N_12121,N_11520,N_11966);
nand U12122 (N_12122,N_11077,N_11435);
and U12123 (N_12123,N_11001,N_11052);
and U12124 (N_12124,N_11534,N_11023);
and U12125 (N_12125,N_11096,N_11422);
and U12126 (N_12126,N_11315,N_11977);
and U12127 (N_12127,N_11457,N_11904);
nand U12128 (N_12128,N_11318,N_11383);
nand U12129 (N_12129,N_11109,N_11059);
nor U12130 (N_12130,N_11538,N_11062);
and U12131 (N_12131,N_11834,N_11397);
and U12132 (N_12132,N_11810,N_11058);
or U12133 (N_12133,N_11287,N_11613);
and U12134 (N_12134,N_11083,N_11408);
nand U12135 (N_12135,N_11328,N_11107);
nand U12136 (N_12136,N_11782,N_11822);
nand U12137 (N_12137,N_11669,N_11774);
or U12138 (N_12138,N_11471,N_11360);
nand U12139 (N_12139,N_11716,N_11965);
nor U12140 (N_12140,N_11138,N_11289);
nand U12141 (N_12141,N_11523,N_11627);
and U12142 (N_12142,N_11685,N_11086);
and U12143 (N_12143,N_11413,N_11982);
and U12144 (N_12144,N_11694,N_11124);
xor U12145 (N_12145,N_11916,N_11197);
or U12146 (N_12146,N_11229,N_11038);
and U12147 (N_12147,N_11582,N_11908);
nor U12148 (N_12148,N_11031,N_11030);
and U12149 (N_12149,N_11470,N_11349);
nand U12150 (N_12150,N_11127,N_11153);
xnor U12151 (N_12151,N_11495,N_11713);
nand U12152 (N_12152,N_11152,N_11945);
xor U12153 (N_12153,N_11332,N_11099);
or U12154 (N_12154,N_11652,N_11532);
nand U12155 (N_12155,N_11440,N_11554);
or U12156 (N_12156,N_11310,N_11097);
and U12157 (N_12157,N_11873,N_11612);
and U12158 (N_12158,N_11182,N_11788);
and U12159 (N_12159,N_11226,N_11280);
and U12160 (N_12160,N_11473,N_11250);
and U12161 (N_12161,N_11373,N_11479);
xnor U12162 (N_12162,N_11990,N_11924);
nor U12163 (N_12163,N_11449,N_11559);
and U12164 (N_12164,N_11626,N_11428);
and U12165 (N_12165,N_11915,N_11623);
and U12166 (N_12166,N_11041,N_11926);
or U12167 (N_12167,N_11335,N_11304);
nor U12168 (N_12168,N_11222,N_11370);
or U12169 (N_12169,N_11385,N_11519);
xnor U12170 (N_12170,N_11344,N_11223);
nor U12171 (N_12171,N_11909,N_11384);
or U12172 (N_12172,N_11728,N_11581);
and U12173 (N_12173,N_11117,N_11703);
or U12174 (N_12174,N_11027,N_11014);
nand U12175 (N_12175,N_11987,N_11290);
and U12176 (N_12176,N_11895,N_11211);
nand U12177 (N_12177,N_11841,N_11770);
or U12178 (N_12178,N_11679,N_11454);
xor U12179 (N_12179,N_11553,N_11120);
or U12180 (N_12180,N_11962,N_11804);
nor U12181 (N_12181,N_11814,N_11947);
and U12182 (N_12182,N_11111,N_11979);
nand U12183 (N_12183,N_11217,N_11791);
and U12184 (N_12184,N_11350,N_11546);
and U12185 (N_12185,N_11942,N_11264);
nor U12186 (N_12186,N_11491,N_11283);
nor U12187 (N_12187,N_11545,N_11358);
nand U12188 (N_12188,N_11901,N_11969);
and U12189 (N_12189,N_11244,N_11568);
xor U12190 (N_12190,N_11688,N_11154);
nor U12191 (N_12191,N_11789,N_11053);
nand U12192 (N_12192,N_11828,N_11464);
nand U12193 (N_12193,N_11684,N_11893);
nand U12194 (N_12194,N_11927,N_11840);
nor U12195 (N_12195,N_11416,N_11753);
nand U12196 (N_12196,N_11835,N_11411);
xnor U12197 (N_12197,N_11708,N_11320);
xor U12198 (N_12198,N_11859,N_11599);
nand U12199 (N_12199,N_11455,N_11637);
nand U12200 (N_12200,N_11653,N_11849);
or U12201 (N_12201,N_11073,N_11550);
nand U12202 (N_12202,N_11487,N_11311);
nor U12203 (N_12203,N_11032,N_11494);
nor U12204 (N_12204,N_11480,N_11997);
nand U12205 (N_12205,N_11596,N_11375);
xor U12206 (N_12206,N_11720,N_11143);
nand U12207 (N_12207,N_11586,N_11382);
and U12208 (N_12208,N_11907,N_11192);
nand U12209 (N_12209,N_11432,N_11923);
and U12210 (N_12210,N_11043,N_11286);
and U12211 (N_12211,N_11589,N_11137);
xor U12212 (N_12212,N_11299,N_11206);
xor U12213 (N_12213,N_11288,N_11021);
nor U12214 (N_12214,N_11434,N_11442);
nor U12215 (N_12215,N_11141,N_11160);
nor U12216 (N_12216,N_11850,N_11934);
or U12217 (N_12217,N_11263,N_11775);
or U12218 (N_12218,N_11749,N_11415);
nor U12219 (N_12219,N_11249,N_11324);
and U12220 (N_12220,N_11297,N_11960);
nand U12221 (N_12221,N_11401,N_11475);
or U12222 (N_12222,N_11807,N_11105);
xnor U12223 (N_12223,N_11614,N_11717);
nor U12224 (N_12224,N_11171,N_11305);
or U12225 (N_12225,N_11674,N_11762);
or U12226 (N_12226,N_11801,N_11374);
or U12227 (N_12227,N_11821,N_11170);
nand U12228 (N_12228,N_11967,N_11848);
nand U12229 (N_12229,N_11956,N_11750);
or U12230 (N_12230,N_11220,N_11885);
nand U12231 (N_12231,N_11949,N_11274);
nand U12232 (N_12232,N_11458,N_11221);
or U12233 (N_12233,N_11087,N_11248);
and U12234 (N_12234,N_11018,N_11129);
nor U12235 (N_12235,N_11268,N_11276);
nand U12236 (N_12236,N_11429,N_11500);
or U12237 (N_12237,N_11735,N_11701);
nand U12238 (N_12238,N_11980,N_11341);
and U12239 (N_12239,N_11547,N_11204);
nand U12240 (N_12240,N_11233,N_11321);
and U12241 (N_12241,N_11173,N_11729);
nand U12242 (N_12242,N_11347,N_11352);
nor U12243 (N_12243,N_11460,N_11748);
nand U12244 (N_12244,N_11961,N_11194);
and U12245 (N_12245,N_11504,N_11467);
nor U12246 (N_12246,N_11162,N_11183);
and U12247 (N_12247,N_11628,N_11543);
nor U12248 (N_12248,N_11871,N_11622);
nor U12249 (N_12249,N_11601,N_11651);
or U12250 (N_12250,N_11177,N_11608);
xor U12251 (N_12251,N_11533,N_11195);
or U12252 (N_12252,N_11824,N_11447);
nand U12253 (N_12253,N_11313,N_11414);
nand U12254 (N_12254,N_11604,N_11594);
or U12255 (N_12255,N_11832,N_11894);
nand U12256 (N_12256,N_11536,N_11726);
and U12257 (N_12257,N_11864,N_11968);
or U12258 (N_12258,N_11992,N_11744);
nand U12259 (N_12259,N_11079,N_11258);
and U12260 (N_12260,N_11279,N_11564);
nand U12261 (N_12261,N_11325,N_11048);
xor U12262 (N_12262,N_11036,N_11241);
or U12263 (N_12263,N_11875,N_11456);
xor U12264 (N_12264,N_11763,N_11575);
and U12265 (N_12265,N_11201,N_11827);
nor U12266 (N_12266,N_11126,N_11168);
nand U12267 (N_12267,N_11163,N_11140);
nand U12268 (N_12268,N_11863,N_11336);
nor U12269 (N_12269,N_11584,N_11113);
nand U12270 (N_12270,N_11198,N_11971);
xor U12271 (N_12271,N_11405,N_11112);
and U12272 (N_12272,N_11820,N_11631);
nor U12273 (N_12273,N_11852,N_11427);
nor U12274 (N_12274,N_11667,N_11797);
nor U12275 (N_12275,N_11441,N_11809);
nor U12276 (N_12276,N_11777,N_11783);
xnor U12277 (N_12277,N_11625,N_11022);
nand U12278 (N_12278,N_11224,N_11499);
nand U12279 (N_12279,N_11776,N_11696);
nor U12280 (N_12280,N_11769,N_11681);
or U12281 (N_12281,N_11024,N_11697);
and U12282 (N_12282,N_11282,N_11157);
nand U12283 (N_12283,N_11388,N_11817);
xnor U12284 (N_12284,N_11698,N_11606);
nor U12285 (N_12285,N_11799,N_11501);
nand U12286 (N_12286,N_11847,N_11139);
and U12287 (N_12287,N_11085,N_11231);
or U12288 (N_12288,N_11216,N_11913);
xor U12289 (N_12289,N_11110,N_11571);
xor U12290 (N_12290,N_11597,N_11144);
nor U12291 (N_12291,N_11267,N_11136);
nand U12292 (N_12292,N_11743,N_11010);
nor U12293 (N_12293,N_11147,N_11796);
nor U12294 (N_12294,N_11865,N_11378);
and U12295 (N_12295,N_11253,N_11754);
nor U12296 (N_12296,N_11172,N_11420);
xor U12297 (N_12297,N_11277,N_11940);
nand U12298 (N_12298,N_11272,N_11756);
nor U12299 (N_12299,N_11098,N_11150);
nor U12300 (N_12300,N_11044,N_11906);
nand U12301 (N_12301,N_11453,N_11853);
and U12302 (N_12302,N_11560,N_11936);
xor U12303 (N_12303,N_11179,N_11175);
xnor U12304 (N_12304,N_11890,N_11169);
or U12305 (N_12305,N_11642,N_11764);
nor U12306 (N_12306,N_11530,N_11525);
xnor U12307 (N_12307,N_11240,N_11825);
and U12308 (N_12308,N_11186,N_11752);
nor U12309 (N_12309,N_11811,N_11259);
nor U12310 (N_12310,N_11188,N_11448);
nor U12311 (N_12311,N_11338,N_11995);
and U12312 (N_12312,N_11787,N_11235);
nor U12313 (N_12313,N_11294,N_11831);
or U12314 (N_12314,N_11646,N_11578);
nor U12315 (N_12315,N_11426,N_11254);
or U12316 (N_12316,N_11367,N_11242);
or U12317 (N_12317,N_11573,N_11868);
xor U12318 (N_12318,N_11953,N_11747);
and U12319 (N_12319,N_11629,N_11404);
or U12320 (N_12320,N_11690,N_11490);
and U12321 (N_12321,N_11739,N_11502);
nor U12322 (N_12322,N_11903,N_11780);
and U12323 (N_12323,N_11131,N_11072);
nor U12324 (N_12324,N_11065,N_11069);
and U12325 (N_12325,N_11496,N_11549);
and U12326 (N_12326,N_11323,N_11883);
nand U12327 (N_12327,N_11689,N_11891);
or U12328 (N_12328,N_11371,N_11064);
or U12329 (N_12329,N_11630,N_11830);
nor U12330 (N_12330,N_11719,N_11736);
and U12331 (N_12331,N_11537,N_11759);
or U12332 (N_12332,N_11619,N_11857);
and U12333 (N_12333,N_11808,N_11795);
or U12334 (N_12334,N_11580,N_11063);
or U12335 (N_12335,N_11243,N_11213);
and U12336 (N_12336,N_11025,N_11540);
or U12337 (N_12337,N_11102,N_11624);
or U12338 (N_12338,N_11029,N_11342);
nor U12339 (N_12339,N_11989,N_11558);
nand U12340 (N_12340,N_11219,N_11647);
or U12341 (N_12341,N_11921,N_11943);
nor U12342 (N_12342,N_11988,N_11656);
or U12343 (N_12343,N_11918,N_11858);
or U12344 (N_12344,N_11257,N_11308);
and U12345 (N_12345,N_11035,N_11585);
nand U12346 (N_12346,N_11590,N_11293);
and U12347 (N_12347,N_11615,N_11051);
or U12348 (N_12348,N_11327,N_11711);
nand U12349 (N_12349,N_11189,N_11722);
nor U12350 (N_12350,N_11209,N_11765);
and U12351 (N_12351,N_11399,N_11952);
nor U12352 (N_12352,N_11768,N_11461);
nor U12353 (N_12353,N_11930,N_11699);
nor U12354 (N_12354,N_11794,N_11839);
xnor U12355 (N_12355,N_11517,N_11518);
nand U12356 (N_12356,N_11838,N_11778);
and U12357 (N_12357,N_11815,N_11870);
nor U12358 (N_12358,N_11643,N_11056);
nor U12359 (N_12359,N_11746,N_11664);
and U12360 (N_12360,N_11424,N_11826);
and U12361 (N_12361,N_11122,N_11551);
or U12362 (N_12362,N_11002,N_11156);
nor U12363 (N_12363,N_11205,N_11298);
nand U12364 (N_12364,N_11067,N_11676);
and U12365 (N_12365,N_11583,N_11265);
nand U12366 (N_12366,N_11854,N_11632);
nor U12367 (N_12367,N_11773,N_11639);
or U12368 (N_12368,N_11128,N_11463);
nor U12369 (N_12369,N_11202,N_11665);
and U12370 (N_12370,N_11130,N_11100);
nand U12371 (N_12371,N_11187,N_11042);
nor U12372 (N_12372,N_11935,N_11238);
and U12373 (N_12373,N_11074,N_11474);
nand U12374 (N_12374,N_11395,N_11236);
nand U12375 (N_12375,N_11104,N_11333);
nor U12376 (N_12376,N_11049,N_11252);
or U12377 (N_12377,N_11291,N_11331);
and U12378 (N_12378,N_11218,N_11561);
nand U12379 (N_12379,N_11572,N_11028);
nand U12380 (N_12380,N_11228,N_11090);
nand U12381 (N_12381,N_11084,N_11121);
and U12382 (N_12382,N_11176,N_11521);
and U12383 (N_12383,N_11529,N_11365);
xnor U12384 (N_12384,N_11755,N_11469);
nor U12385 (N_12385,N_11307,N_11869);
xor U12386 (N_12386,N_11430,N_11737);
and U12387 (N_12387,N_11234,N_11896);
xor U12388 (N_12388,N_11766,N_11929);
nor U12389 (N_12389,N_11668,N_11180);
and U12390 (N_12390,N_11312,N_11275);
and U12391 (N_12391,N_11999,N_11732);
nand U12392 (N_12392,N_11007,N_11459);
nor U12393 (N_12393,N_11273,N_11088);
nor U12394 (N_12394,N_11292,N_11649);
nand U12395 (N_12395,N_11472,N_11640);
or U12396 (N_12396,N_11555,N_11905);
and U12397 (N_12397,N_11812,N_11005);
nor U12398 (N_12398,N_11955,N_11142);
nor U12399 (N_12399,N_11497,N_11403);
nor U12400 (N_12400,N_11450,N_11803);
nor U12401 (N_12401,N_11000,N_11705);
or U12402 (N_12402,N_11937,N_11094);
xnor U12403 (N_12403,N_11963,N_11446);
nand U12404 (N_12404,N_11303,N_11193);
nand U12405 (N_12405,N_11946,N_11040);
nand U12406 (N_12406,N_11851,N_11468);
and U12407 (N_12407,N_11970,N_11660);
xnor U12408 (N_12408,N_11326,N_11343);
and U12409 (N_12409,N_11591,N_11114);
or U12410 (N_12410,N_11757,N_11381);
or U12411 (N_12411,N_11492,N_11986);
nand U12412 (N_12412,N_11266,N_11600);
or U12413 (N_12413,N_11715,N_11880);
or U12414 (N_12414,N_11761,N_11725);
nand U12415 (N_12415,N_11081,N_11897);
and U12416 (N_12416,N_11806,N_11145);
or U12417 (N_12417,N_11718,N_11438);
nand U12418 (N_12418,N_11227,N_11481);
nand U12419 (N_12419,N_11802,N_11082);
nor U12420 (N_12420,N_11225,N_11076);
and U12421 (N_12421,N_11230,N_11861);
and U12422 (N_12422,N_11118,N_11993);
xnor U12423 (N_12423,N_11565,N_11950);
and U12424 (N_12424,N_11133,N_11181);
nor U12425 (N_12425,N_11638,N_11466);
nor U12426 (N_12426,N_11569,N_11366);
xnor U12427 (N_12427,N_11994,N_11199);
and U12428 (N_12428,N_11862,N_11398);
nor U12429 (N_12429,N_11506,N_11132);
nand U12430 (N_12430,N_11842,N_11892);
nand U12431 (N_12431,N_11485,N_11675);
nor U12432 (N_12432,N_11958,N_11060);
or U12433 (N_12433,N_11531,N_11607);
nand U12434 (N_12434,N_11078,N_11741);
or U12435 (N_12435,N_11771,N_11785);
and U12436 (N_12436,N_11898,N_11451);
or U12437 (N_12437,N_11567,N_11846);
nand U12438 (N_12438,N_11611,N_11671);
or U12439 (N_12439,N_11011,N_11505);
nor U12440 (N_12440,N_11706,N_11702);
or U12441 (N_12441,N_11034,N_11300);
xor U12442 (N_12442,N_11301,N_11983);
or U12443 (N_12443,N_11917,N_11700);
and U12444 (N_12444,N_11867,N_11511);
nand U12445 (N_12445,N_11932,N_11488);
nor U12446 (N_12446,N_11354,N_11444);
nor U12447 (N_12447,N_11843,N_11306);
or U12448 (N_12448,N_11039,N_11155);
nor U12449 (N_12449,N_11887,N_11603);
xor U12450 (N_12450,N_11693,N_11562);
and U12451 (N_12451,N_11874,N_11709);
xor U12452 (N_12452,N_11570,N_11116);
nand U12453 (N_12453,N_11108,N_11392);
and U12454 (N_12454,N_11616,N_11944);
and U12455 (N_12455,N_11680,N_11262);
nor U12456 (N_12456,N_11866,N_11641);
and U12457 (N_12457,N_11678,N_11407);
nor U12458 (N_12458,N_11758,N_11574);
nor U12459 (N_12459,N_11507,N_11939);
or U12460 (N_12460,N_11368,N_11633);
nor U12461 (N_12461,N_11677,N_11161);
or U12462 (N_12462,N_11941,N_11178);
or U12463 (N_12463,N_11767,N_11576);
xnor U12464 (N_12464,N_11055,N_11695);
and U12465 (N_12465,N_11004,N_11745);
nor U12466 (N_12466,N_11396,N_11261);
nor U12467 (N_12467,N_11587,N_11595);
or U12468 (N_12468,N_11662,N_11493);
nor U12469 (N_12469,N_11951,N_11779);
and U12470 (N_12470,N_11645,N_11232);
and U12471 (N_12471,N_11068,N_11650);
or U12472 (N_12472,N_11309,N_11818);
xnor U12473 (N_12473,N_11356,N_11070);
or U12474 (N_12474,N_11406,N_11884);
xnor U12475 (N_12475,N_11790,N_11400);
nor U12476 (N_12476,N_11527,N_11200);
or U12477 (N_12477,N_11813,N_11856);
and U12478 (N_12478,N_11394,N_11174);
and U12479 (N_12479,N_11054,N_11050);
or U12480 (N_12480,N_11075,N_11037);
nand U12481 (N_12481,N_11389,N_11663);
or U12482 (N_12482,N_11423,N_11976);
nand U12483 (N_12483,N_11284,N_11295);
or U12484 (N_12484,N_11425,N_11526);
nor U12485 (N_12485,N_11363,N_11208);
or U12486 (N_12486,N_11476,N_11882);
nand U12487 (N_12487,N_11837,N_11740);
xnor U12488 (N_12488,N_11372,N_11515);
and U12489 (N_12489,N_11670,N_11436);
nand U12490 (N_12490,N_11712,N_11135);
and U12491 (N_12491,N_11886,N_11215);
or U12492 (N_12492,N_11498,N_11984);
xnor U12493 (N_12493,N_11566,N_11659);
nand U12494 (N_12494,N_11925,N_11742);
and U12495 (N_12495,N_11091,N_11602);
nor U12496 (N_12496,N_11190,N_11103);
nor U12497 (N_12497,N_11974,N_11346);
or U12498 (N_12498,N_11878,N_11391);
or U12499 (N_12499,N_11888,N_11512);
or U12500 (N_12500,N_11055,N_11399);
and U12501 (N_12501,N_11592,N_11125);
and U12502 (N_12502,N_11973,N_11610);
xor U12503 (N_12503,N_11630,N_11186);
or U12504 (N_12504,N_11228,N_11088);
and U12505 (N_12505,N_11776,N_11320);
nor U12506 (N_12506,N_11444,N_11050);
nor U12507 (N_12507,N_11804,N_11776);
or U12508 (N_12508,N_11490,N_11561);
or U12509 (N_12509,N_11617,N_11621);
and U12510 (N_12510,N_11872,N_11585);
nand U12511 (N_12511,N_11856,N_11118);
or U12512 (N_12512,N_11093,N_11462);
nand U12513 (N_12513,N_11946,N_11500);
nor U12514 (N_12514,N_11695,N_11440);
nor U12515 (N_12515,N_11827,N_11261);
xnor U12516 (N_12516,N_11813,N_11373);
nor U12517 (N_12517,N_11211,N_11425);
nand U12518 (N_12518,N_11664,N_11288);
or U12519 (N_12519,N_11013,N_11169);
nand U12520 (N_12520,N_11840,N_11427);
and U12521 (N_12521,N_11494,N_11436);
or U12522 (N_12522,N_11703,N_11673);
nand U12523 (N_12523,N_11976,N_11458);
nand U12524 (N_12524,N_11251,N_11667);
nand U12525 (N_12525,N_11727,N_11185);
or U12526 (N_12526,N_11317,N_11609);
or U12527 (N_12527,N_11996,N_11537);
and U12528 (N_12528,N_11306,N_11346);
or U12529 (N_12529,N_11468,N_11966);
nand U12530 (N_12530,N_11603,N_11948);
and U12531 (N_12531,N_11002,N_11241);
nand U12532 (N_12532,N_11576,N_11292);
nand U12533 (N_12533,N_11058,N_11384);
nand U12534 (N_12534,N_11844,N_11089);
xnor U12535 (N_12535,N_11731,N_11681);
or U12536 (N_12536,N_11905,N_11135);
or U12537 (N_12537,N_11750,N_11091);
nor U12538 (N_12538,N_11514,N_11539);
or U12539 (N_12539,N_11939,N_11664);
nand U12540 (N_12540,N_11296,N_11041);
and U12541 (N_12541,N_11274,N_11203);
nor U12542 (N_12542,N_11825,N_11553);
or U12543 (N_12543,N_11378,N_11505);
nand U12544 (N_12544,N_11874,N_11227);
or U12545 (N_12545,N_11187,N_11968);
nor U12546 (N_12546,N_11817,N_11673);
nor U12547 (N_12547,N_11642,N_11206);
and U12548 (N_12548,N_11211,N_11776);
nand U12549 (N_12549,N_11445,N_11731);
and U12550 (N_12550,N_11559,N_11614);
or U12551 (N_12551,N_11079,N_11321);
nand U12552 (N_12552,N_11765,N_11792);
nor U12553 (N_12553,N_11752,N_11119);
and U12554 (N_12554,N_11666,N_11245);
or U12555 (N_12555,N_11211,N_11812);
and U12556 (N_12556,N_11649,N_11965);
or U12557 (N_12557,N_11017,N_11798);
or U12558 (N_12558,N_11549,N_11229);
nand U12559 (N_12559,N_11417,N_11259);
and U12560 (N_12560,N_11071,N_11136);
nand U12561 (N_12561,N_11707,N_11234);
nand U12562 (N_12562,N_11172,N_11248);
and U12563 (N_12563,N_11418,N_11786);
nand U12564 (N_12564,N_11027,N_11009);
and U12565 (N_12565,N_11929,N_11079);
nor U12566 (N_12566,N_11161,N_11333);
nand U12567 (N_12567,N_11188,N_11036);
nor U12568 (N_12568,N_11217,N_11207);
or U12569 (N_12569,N_11680,N_11625);
or U12570 (N_12570,N_11499,N_11997);
nor U12571 (N_12571,N_11361,N_11619);
nand U12572 (N_12572,N_11344,N_11519);
nand U12573 (N_12573,N_11441,N_11221);
or U12574 (N_12574,N_11821,N_11055);
nand U12575 (N_12575,N_11666,N_11208);
xor U12576 (N_12576,N_11906,N_11784);
nor U12577 (N_12577,N_11837,N_11037);
or U12578 (N_12578,N_11721,N_11019);
nor U12579 (N_12579,N_11959,N_11189);
and U12580 (N_12580,N_11761,N_11460);
nand U12581 (N_12581,N_11727,N_11951);
or U12582 (N_12582,N_11257,N_11149);
nor U12583 (N_12583,N_11299,N_11950);
nor U12584 (N_12584,N_11435,N_11298);
nor U12585 (N_12585,N_11051,N_11044);
nand U12586 (N_12586,N_11759,N_11398);
xnor U12587 (N_12587,N_11867,N_11891);
and U12588 (N_12588,N_11184,N_11884);
nor U12589 (N_12589,N_11839,N_11457);
and U12590 (N_12590,N_11287,N_11875);
and U12591 (N_12591,N_11998,N_11949);
and U12592 (N_12592,N_11971,N_11896);
or U12593 (N_12593,N_11558,N_11953);
nand U12594 (N_12594,N_11733,N_11327);
or U12595 (N_12595,N_11706,N_11769);
and U12596 (N_12596,N_11144,N_11872);
or U12597 (N_12597,N_11954,N_11781);
or U12598 (N_12598,N_11462,N_11641);
nor U12599 (N_12599,N_11873,N_11839);
and U12600 (N_12600,N_11587,N_11870);
nand U12601 (N_12601,N_11537,N_11523);
nand U12602 (N_12602,N_11897,N_11014);
or U12603 (N_12603,N_11160,N_11130);
and U12604 (N_12604,N_11119,N_11464);
nor U12605 (N_12605,N_11535,N_11325);
nand U12606 (N_12606,N_11822,N_11761);
nand U12607 (N_12607,N_11690,N_11428);
and U12608 (N_12608,N_11953,N_11042);
nor U12609 (N_12609,N_11634,N_11358);
and U12610 (N_12610,N_11675,N_11583);
nor U12611 (N_12611,N_11879,N_11934);
and U12612 (N_12612,N_11770,N_11625);
nor U12613 (N_12613,N_11310,N_11171);
nor U12614 (N_12614,N_11766,N_11667);
nor U12615 (N_12615,N_11540,N_11138);
nor U12616 (N_12616,N_11929,N_11173);
xor U12617 (N_12617,N_11660,N_11005);
nor U12618 (N_12618,N_11623,N_11406);
nor U12619 (N_12619,N_11438,N_11406);
or U12620 (N_12620,N_11789,N_11308);
and U12621 (N_12621,N_11114,N_11108);
nand U12622 (N_12622,N_11204,N_11073);
or U12623 (N_12623,N_11876,N_11821);
and U12624 (N_12624,N_11010,N_11271);
and U12625 (N_12625,N_11850,N_11199);
and U12626 (N_12626,N_11609,N_11596);
xor U12627 (N_12627,N_11489,N_11729);
nand U12628 (N_12628,N_11418,N_11356);
nor U12629 (N_12629,N_11082,N_11839);
and U12630 (N_12630,N_11484,N_11306);
nand U12631 (N_12631,N_11020,N_11585);
and U12632 (N_12632,N_11925,N_11596);
nor U12633 (N_12633,N_11461,N_11531);
and U12634 (N_12634,N_11161,N_11928);
xor U12635 (N_12635,N_11117,N_11054);
xor U12636 (N_12636,N_11623,N_11807);
and U12637 (N_12637,N_11854,N_11417);
xnor U12638 (N_12638,N_11685,N_11798);
xnor U12639 (N_12639,N_11401,N_11755);
and U12640 (N_12640,N_11781,N_11960);
xor U12641 (N_12641,N_11292,N_11882);
or U12642 (N_12642,N_11628,N_11929);
or U12643 (N_12643,N_11231,N_11267);
nand U12644 (N_12644,N_11462,N_11938);
and U12645 (N_12645,N_11268,N_11684);
xnor U12646 (N_12646,N_11619,N_11858);
and U12647 (N_12647,N_11231,N_11708);
and U12648 (N_12648,N_11611,N_11306);
nor U12649 (N_12649,N_11723,N_11315);
xnor U12650 (N_12650,N_11262,N_11490);
xnor U12651 (N_12651,N_11621,N_11317);
nor U12652 (N_12652,N_11959,N_11595);
nor U12653 (N_12653,N_11994,N_11483);
nand U12654 (N_12654,N_11366,N_11673);
and U12655 (N_12655,N_11126,N_11428);
nand U12656 (N_12656,N_11832,N_11506);
nand U12657 (N_12657,N_11558,N_11904);
or U12658 (N_12658,N_11363,N_11501);
nand U12659 (N_12659,N_11250,N_11454);
nor U12660 (N_12660,N_11710,N_11078);
nor U12661 (N_12661,N_11456,N_11322);
or U12662 (N_12662,N_11250,N_11636);
or U12663 (N_12663,N_11178,N_11351);
and U12664 (N_12664,N_11997,N_11288);
or U12665 (N_12665,N_11949,N_11789);
nor U12666 (N_12666,N_11288,N_11701);
nand U12667 (N_12667,N_11265,N_11026);
nor U12668 (N_12668,N_11566,N_11046);
nand U12669 (N_12669,N_11997,N_11680);
nand U12670 (N_12670,N_11693,N_11424);
nor U12671 (N_12671,N_11382,N_11564);
nor U12672 (N_12672,N_11513,N_11924);
and U12673 (N_12673,N_11189,N_11341);
nor U12674 (N_12674,N_11961,N_11123);
and U12675 (N_12675,N_11169,N_11370);
and U12676 (N_12676,N_11581,N_11321);
or U12677 (N_12677,N_11438,N_11585);
nor U12678 (N_12678,N_11593,N_11308);
or U12679 (N_12679,N_11952,N_11829);
nand U12680 (N_12680,N_11330,N_11349);
xor U12681 (N_12681,N_11098,N_11220);
and U12682 (N_12682,N_11156,N_11501);
nor U12683 (N_12683,N_11467,N_11386);
or U12684 (N_12684,N_11950,N_11773);
xor U12685 (N_12685,N_11256,N_11084);
nand U12686 (N_12686,N_11491,N_11954);
and U12687 (N_12687,N_11235,N_11711);
nor U12688 (N_12688,N_11880,N_11081);
nand U12689 (N_12689,N_11575,N_11158);
xnor U12690 (N_12690,N_11631,N_11064);
or U12691 (N_12691,N_11707,N_11620);
and U12692 (N_12692,N_11780,N_11463);
and U12693 (N_12693,N_11659,N_11231);
and U12694 (N_12694,N_11659,N_11159);
or U12695 (N_12695,N_11494,N_11187);
and U12696 (N_12696,N_11103,N_11614);
nand U12697 (N_12697,N_11717,N_11520);
nand U12698 (N_12698,N_11313,N_11814);
nand U12699 (N_12699,N_11183,N_11870);
or U12700 (N_12700,N_11398,N_11619);
or U12701 (N_12701,N_11962,N_11734);
nor U12702 (N_12702,N_11848,N_11901);
nand U12703 (N_12703,N_11419,N_11512);
nor U12704 (N_12704,N_11161,N_11293);
nand U12705 (N_12705,N_11466,N_11137);
or U12706 (N_12706,N_11073,N_11072);
and U12707 (N_12707,N_11401,N_11528);
xor U12708 (N_12708,N_11520,N_11980);
or U12709 (N_12709,N_11094,N_11746);
and U12710 (N_12710,N_11617,N_11871);
xor U12711 (N_12711,N_11610,N_11183);
and U12712 (N_12712,N_11428,N_11508);
nor U12713 (N_12713,N_11517,N_11687);
or U12714 (N_12714,N_11773,N_11074);
nor U12715 (N_12715,N_11415,N_11750);
or U12716 (N_12716,N_11642,N_11355);
nor U12717 (N_12717,N_11188,N_11470);
nand U12718 (N_12718,N_11912,N_11725);
and U12719 (N_12719,N_11503,N_11880);
nand U12720 (N_12720,N_11791,N_11550);
or U12721 (N_12721,N_11287,N_11339);
nor U12722 (N_12722,N_11501,N_11234);
xnor U12723 (N_12723,N_11222,N_11862);
nor U12724 (N_12724,N_11493,N_11652);
xor U12725 (N_12725,N_11780,N_11484);
nor U12726 (N_12726,N_11834,N_11767);
or U12727 (N_12727,N_11457,N_11031);
nand U12728 (N_12728,N_11561,N_11854);
or U12729 (N_12729,N_11677,N_11952);
nand U12730 (N_12730,N_11508,N_11033);
nor U12731 (N_12731,N_11003,N_11551);
xnor U12732 (N_12732,N_11946,N_11959);
nand U12733 (N_12733,N_11531,N_11348);
nand U12734 (N_12734,N_11754,N_11821);
xnor U12735 (N_12735,N_11289,N_11496);
nand U12736 (N_12736,N_11220,N_11549);
xor U12737 (N_12737,N_11601,N_11117);
nor U12738 (N_12738,N_11891,N_11420);
nor U12739 (N_12739,N_11836,N_11785);
or U12740 (N_12740,N_11777,N_11668);
nand U12741 (N_12741,N_11761,N_11896);
xnor U12742 (N_12742,N_11510,N_11628);
nor U12743 (N_12743,N_11106,N_11498);
and U12744 (N_12744,N_11691,N_11132);
and U12745 (N_12745,N_11157,N_11881);
and U12746 (N_12746,N_11797,N_11176);
or U12747 (N_12747,N_11100,N_11506);
or U12748 (N_12748,N_11453,N_11289);
and U12749 (N_12749,N_11099,N_11908);
nand U12750 (N_12750,N_11859,N_11122);
and U12751 (N_12751,N_11368,N_11760);
nand U12752 (N_12752,N_11718,N_11213);
nor U12753 (N_12753,N_11480,N_11671);
xnor U12754 (N_12754,N_11088,N_11618);
nand U12755 (N_12755,N_11232,N_11892);
and U12756 (N_12756,N_11867,N_11044);
and U12757 (N_12757,N_11439,N_11639);
and U12758 (N_12758,N_11655,N_11066);
and U12759 (N_12759,N_11387,N_11440);
nor U12760 (N_12760,N_11665,N_11948);
nor U12761 (N_12761,N_11429,N_11016);
nor U12762 (N_12762,N_11982,N_11494);
and U12763 (N_12763,N_11665,N_11408);
nor U12764 (N_12764,N_11930,N_11738);
nand U12765 (N_12765,N_11567,N_11631);
or U12766 (N_12766,N_11452,N_11702);
nand U12767 (N_12767,N_11046,N_11932);
nand U12768 (N_12768,N_11683,N_11127);
or U12769 (N_12769,N_11045,N_11499);
nor U12770 (N_12770,N_11636,N_11169);
nor U12771 (N_12771,N_11679,N_11819);
nor U12772 (N_12772,N_11974,N_11255);
and U12773 (N_12773,N_11113,N_11496);
nand U12774 (N_12774,N_11944,N_11729);
and U12775 (N_12775,N_11608,N_11876);
xor U12776 (N_12776,N_11740,N_11536);
and U12777 (N_12777,N_11817,N_11423);
nor U12778 (N_12778,N_11087,N_11713);
nand U12779 (N_12779,N_11162,N_11194);
nor U12780 (N_12780,N_11879,N_11471);
and U12781 (N_12781,N_11704,N_11118);
nand U12782 (N_12782,N_11103,N_11350);
xor U12783 (N_12783,N_11813,N_11635);
or U12784 (N_12784,N_11905,N_11168);
nor U12785 (N_12785,N_11506,N_11766);
xnor U12786 (N_12786,N_11063,N_11372);
nor U12787 (N_12787,N_11267,N_11212);
and U12788 (N_12788,N_11889,N_11482);
xnor U12789 (N_12789,N_11485,N_11131);
and U12790 (N_12790,N_11888,N_11301);
nand U12791 (N_12791,N_11990,N_11725);
xor U12792 (N_12792,N_11925,N_11482);
and U12793 (N_12793,N_11554,N_11225);
and U12794 (N_12794,N_11188,N_11923);
xor U12795 (N_12795,N_11739,N_11900);
or U12796 (N_12796,N_11186,N_11853);
nor U12797 (N_12797,N_11736,N_11223);
or U12798 (N_12798,N_11187,N_11513);
and U12799 (N_12799,N_11874,N_11397);
nor U12800 (N_12800,N_11689,N_11543);
nand U12801 (N_12801,N_11757,N_11554);
xor U12802 (N_12802,N_11950,N_11442);
nor U12803 (N_12803,N_11556,N_11780);
xnor U12804 (N_12804,N_11748,N_11632);
nor U12805 (N_12805,N_11893,N_11170);
nand U12806 (N_12806,N_11154,N_11628);
and U12807 (N_12807,N_11329,N_11607);
or U12808 (N_12808,N_11406,N_11624);
nand U12809 (N_12809,N_11347,N_11807);
nor U12810 (N_12810,N_11019,N_11006);
nand U12811 (N_12811,N_11695,N_11091);
nor U12812 (N_12812,N_11415,N_11780);
or U12813 (N_12813,N_11815,N_11749);
or U12814 (N_12814,N_11894,N_11728);
nor U12815 (N_12815,N_11507,N_11161);
or U12816 (N_12816,N_11000,N_11069);
xor U12817 (N_12817,N_11190,N_11362);
or U12818 (N_12818,N_11009,N_11258);
nor U12819 (N_12819,N_11949,N_11460);
nand U12820 (N_12820,N_11741,N_11659);
or U12821 (N_12821,N_11703,N_11069);
or U12822 (N_12822,N_11648,N_11695);
or U12823 (N_12823,N_11842,N_11715);
nor U12824 (N_12824,N_11182,N_11064);
xnor U12825 (N_12825,N_11480,N_11052);
xor U12826 (N_12826,N_11693,N_11063);
nor U12827 (N_12827,N_11434,N_11395);
xnor U12828 (N_12828,N_11596,N_11470);
and U12829 (N_12829,N_11415,N_11571);
xor U12830 (N_12830,N_11718,N_11244);
nor U12831 (N_12831,N_11191,N_11212);
nand U12832 (N_12832,N_11984,N_11153);
nor U12833 (N_12833,N_11742,N_11468);
nand U12834 (N_12834,N_11286,N_11912);
and U12835 (N_12835,N_11342,N_11867);
nor U12836 (N_12836,N_11680,N_11947);
nor U12837 (N_12837,N_11177,N_11789);
nor U12838 (N_12838,N_11361,N_11176);
or U12839 (N_12839,N_11901,N_11150);
nand U12840 (N_12840,N_11550,N_11992);
or U12841 (N_12841,N_11823,N_11530);
nor U12842 (N_12842,N_11125,N_11286);
and U12843 (N_12843,N_11295,N_11494);
nand U12844 (N_12844,N_11345,N_11750);
and U12845 (N_12845,N_11369,N_11960);
nand U12846 (N_12846,N_11160,N_11496);
xnor U12847 (N_12847,N_11545,N_11909);
nor U12848 (N_12848,N_11126,N_11862);
or U12849 (N_12849,N_11681,N_11177);
and U12850 (N_12850,N_11102,N_11057);
or U12851 (N_12851,N_11975,N_11093);
and U12852 (N_12852,N_11029,N_11917);
nand U12853 (N_12853,N_11971,N_11183);
nor U12854 (N_12854,N_11525,N_11091);
or U12855 (N_12855,N_11485,N_11765);
nor U12856 (N_12856,N_11590,N_11268);
nor U12857 (N_12857,N_11940,N_11803);
nand U12858 (N_12858,N_11053,N_11362);
nand U12859 (N_12859,N_11035,N_11443);
and U12860 (N_12860,N_11725,N_11269);
nand U12861 (N_12861,N_11744,N_11690);
nor U12862 (N_12862,N_11480,N_11219);
nor U12863 (N_12863,N_11216,N_11211);
and U12864 (N_12864,N_11310,N_11320);
nor U12865 (N_12865,N_11844,N_11795);
xor U12866 (N_12866,N_11202,N_11369);
nor U12867 (N_12867,N_11278,N_11402);
or U12868 (N_12868,N_11168,N_11579);
xnor U12869 (N_12869,N_11075,N_11787);
nor U12870 (N_12870,N_11649,N_11157);
or U12871 (N_12871,N_11255,N_11626);
nor U12872 (N_12872,N_11350,N_11669);
nor U12873 (N_12873,N_11642,N_11671);
xnor U12874 (N_12874,N_11392,N_11735);
nor U12875 (N_12875,N_11776,N_11660);
and U12876 (N_12876,N_11878,N_11620);
and U12877 (N_12877,N_11797,N_11022);
nor U12878 (N_12878,N_11510,N_11114);
or U12879 (N_12879,N_11923,N_11131);
nor U12880 (N_12880,N_11575,N_11995);
and U12881 (N_12881,N_11713,N_11929);
or U12882 (N_12882,N_11691,N_11196);
xor U12883 (N_12883,N_11946,N_11828);
nand U12884 (N_12884,N_11443,N_11492);
nand U12885 (N_12885,N_11844,N_11826);
nand U12886 (N_12886,N_11535,N_11256);
nor U12887 (N_12887,N_11470,N_11579);
or U12888 (N_12888,N_11060,N_11280);
and U12889 (N_12889,N_11157,N_11593);
and U12890 (N_12890,N_11590,N_11107);
or U12891 (N_12891,N_11076,N_11944);
nand U12892 (N_12892,N_11903,N_11374);
or U12893 (N_12893,N_11219,N_11335);
and U12894 (N_12894,N_11909,N_11581);
xnor U12895 (N_12895,N_11189,N_11680);
or U12896 (N_12896,N_11622,N_11284);
xnor U12897 (N_12897,N_11424,N_11486);
and U12898 (N_12898,N_11893,N_11632);
nand U12899 (N_12899,N_11281,N_11088);
nand U12900 (N_12900,N_11810,N_11396);
and U12901 (N_12901,N_11430,N_11105);
or U12902 (N_12902,N_11102,N_11390);
and U12903 (N_12903,N_11478,N_11193);
nor U12904 (N_12904,N_11020,N_11920);
nand U12905 (N_12905,N_11791,N_11564);
nor U12906 (N_12906,N_11951,N_11494);
or U12907 (N_12907,N_11746,N_11104);
xnor U12908 (N_12908,N_11832,N_11400);
nor U12909 (N_12909,N_11091,N_11747);
nor U12910 (N_12910,N_11203,N_11659);
and U12911 (N_12911,N_11766,N_11273);
nand U12912 (N_12912,N_11981,N_11277);
and U12913 (N_12913,N_11133,N_11099);
and U12914 (N_12914,N_11744,N_11595);
nand U12915 (N_12915,N_11938,N_11075);
or U12916 (N_12916,N_11735,N_11558);
nand U12917 (N_12917,N_11122,N_11081);
nor U12918 (N_12918,N_11944,N_11286);
and U12919 (N_12919,N_11636,N_11455);
nand U12920 (N_12920,N_11011,N_11470);
nand U12921 (N_12921,N_11195,N_11630);
and U12922 (N_12922,N_11632,N_11365);
and U12923 (N_12923,N_11510,N_11671);
nor U12924 (N_12924,N_11246,N_11319);
nand U12925 (N_12925,N_11217,N_11512);
nand U12926 (N_12926,N_11633,N_11742);
nand U12927 (N_12927,N_11177,N_11386);
xnor U12928 (N_12928,N_11461,N_11710);
and U12929 (N_12929,N_11311,N_11235);
or U12930 (N_12930,N_11533,N_11718);
or U12931 (N_12931,N_11489,N_11712);
xor U12932 (N_12932,N_11477,N_11609);
xnor U12933 (N_12933,N_11823,N_11135);
nand U12934 (N_12934,N_11483,N_11811);
or U12935 (N_12935,N_11727,N_11430);
nor U12936 (N_12936,N_11165,N_11090);
nand U12937 (N_12937,N_11610,N_11526);
and U12938 (N_12938,N_11679,N_11736);
xor U12939 (N_12939,N_11049,N_11550);
nand U12940 (N_12940,N_11178,N_11871);
nand U12941 (N_12941,N_11548,N_11994);
and U12942 (N_12942,N_11477,N_11024);
nor U12943 (N_12943,N_11494,N_11670);
nand U12944 (N_12944,N_11713,N_11089);
and U12945 (N_12945,N_11460,N_11236);
and U12946 (N_12946,N_11612,N_11682);
nor U12947 (N_12947,N_11088,N_11380);
nand U12948 (N_12948,N_11560,N_11590);
and U12949 (N_12949,N_11594,N_11344);
nand U12950 (N_12950,N_11853,N_11335);
and U12951 (N_12951,N_11319,N_11595);
and U12952 (N_12952,N_11098,N_11807);
xnor U12953 (N_12953,N_11717,N_11481);
xor U12954 (N_12954,N_11923,N_11455);
nor U12955 (N_12955,N_11999,N_11069);
and U12956 (N_12956,N_11220,N_11374);
nor U12957 (N_12957,N_11679,N_11545);
and U12958 (N_12958,N_11076,N_11178);
nand U12959 (N_12959,N_11800,N_11461);
and U12960 (N_12960,N_11534,N_11886);
nand U12961 (N_12961,N_11473,N_11953);
xnor U12962 (N_12962,N_11363,N_11179);
or U12963 (N_12963,N_11392,N_11948);
nand U12964 (N_12964,N_11790,N_11373);
nand U12965 (N_12965,N_11635,N_11962);
xor U12966 (N_12966,N_11906,N_11690);
or U12967 (N_12967,N_11783,N_11170);
and U12968 (N_12968,N_11245,N_11774);
and U12969 (N_12969,N_11072,N_11917);
nand U12970 (N_12970,N_11384,N_11610);
nand U12971 (N_12971,N_11200,N_11374);
nor U12972 (N_12972,N_11436,N_11216);
or U12973 (N_12973,N_11641,N_11023);
nand U12974 (N_12974,N_11628,N_11481);
nor U12975 (N_12975,N_11804,N_11303);
or U12976 (N_12976,N_11491,N_11363);
nand U12977 (N_12977,N_11252,N_11918);
nor U12978 (N_12978,N_11883,N_11432);
nor U12979 (N_12979,N_11841,N_11666);
nor U12980 (N_12980,N_11351,N_11356);
or U12981 (N_12981,N_11128,N_11922);
xor U12982 (N_12982,N_11822,N_11053);
or U12983 (N_12983,N_11735,N_11496);
nand U12984 (N_12984,N_11452,N_11773);
and U12985 (N_12985,N_11887,N_11675);
xnor U12986 (N_12986,N_11180,N_11407);
nand U12987 (N_12987,N_11545,N_11590);
nor U12988 (N_12988,N_11597,N_11416);
nor U12989 (N_12989,N_11872,N_11094);
nand U12990 (N_12990,N_11377,N_11079);
nor U12991 (N_12991,N_11175,N_11734);
or U12992 (N_12992,N_11752,N_11600);
or U12993 (N_12993,N_11997,N_11242);
and U12994 (N_12994,N_11957,N_11422);
nand U12995 (N_12995,N_11201,N_11553);
nand U12996 (N_12996,N_11228,N_11021);
nand U12997 (N_12997,N_11781,N_11184);
and U12998 (N_12998,N_11490,N_11100);
nor U12999 (N_12999,N_11631,N_11950);
or U13000 (N_13000,N_12423,N_12325);
nand U13001 (N_13001,N_12228,N_12825);
nor U13002 (N_13002,N_12624,N_12638);
nor U13003 (N_13003,N_12412,N_12973);
nor U13004 (N_13004,N_12823,N_12506);
nor U13005 (N_13005,N_12579,N_12290);
nor U13006 (N_13006,N_12575,N_12968);
nor U13007 (N_13007,N_12830,N_12854);
or U13008 (N_13008,N_12381,N_12352);
xor U13009 (N_13009,N_12345,N_12684);
nor U13010 (N_13010,N_12033,N_12204);
or U13011 (N_13011,N_12330,N_12353);
and U13012 (N_13012,N_12809,N_12038);
and U13013 (N_13013,N_12976,N_12961);
and U13014 (N_13014,N_12131,N_12840);
nor U13015 (N_13015,N_12382,N_12877);
nand U13016 (N_13016,N_12483,N_12595);
or U13017 (N_13017,N_12135,N_12489);
nor U13018 (N_13018,N_12343,N_12675);
and U13019 (N_13019,N_12373,N_12372);
nor U13020 (N_13020,N_12570,N_12065);
and U13021 (N_13021,N_12704,N_12056);
or U13022 (N_13022,N_12517,N_12992);
or U13023 (N_13023,N_12113,N_12160);
xor U13024 (N_13024,N_12515,N_12660);
nor U13025 (N_13025,N_12256,N_12878);
nor U13026 (N_13026,N_12838,N_12199);
or U13027 (N_13027,N_12046,N_12607);
and U13028 (N_13028,N_12622,N_12773);
xnor U13029 (N_13029,N_12978,N_12647);
and U13030 (N_13030,N_12405,N_12875);
nor U13031 (N_13031,N_12498,N_12036);
and U13032 (N_13032,N_12674,N_12247);
and U13033 (N_13033,N_12406,N_12533);
and U13034 (N_13034,N_12841,N_12879);
xnor U13035 (N_13035,N_12260,N_12100);
or U13036 (N_13036,N_12418,N_12514);
xor U13037 (N_13037,N_12416,N_12503);
and U13038 (N_13038,N_12022,N_12829);
and U13039 (N_13039,N_12766,N_12760);
or U13040 (N_13040,N_12360,N_12990);
nand U13041 (N_13041,N_12756,N_12009);
xor U13042 (N_13042,N_12466,N_12654);
nand U13043 (N_13043,N_12478,N_12020);
nand U13044 (N_13044,N_12278,N_12114);
nand U13045 (N_13045,N_12634,N_12112);
nor U13046 (N_13046,N_12165,N_12185);
nor U13047 (N_13047,N_12720,N_12433);
nor U13048 (N_13048,N_12292,N_12035);
nor U13049 (N_13049,N_12813,N_12560);
or U13050 (N_13050,N_12557,N_12375);
and U13051 (N_13051,N_12715,N_12337);
and U13052 (N_13052,N_12884,N_12024);
nand U13053 (N_13053,N_12755,N_12816);
or U13054 (N_13054,N_12052,N_12497);
nor U13055 (N_13055,N_12665,N_12346);
or U13056 (N_13056,N_12846,N_12734);
nor U13057 (N_13057,N_12597,N_12267);
or U13058 (N_13058,N_12963,N_12989);
and U13059 (N_13059,N_12926,N_12856);
or U13060 (N_13060,N_12600,N_12094);
nand U13061 (N_13061,N_12646,N_12043);
nor U13062 (N_13062,N_12140,N_12243);
nor U13063 (N_13063,N_12312,N_12355);
or U13064 (N_13064,N_12387,N_12429);
nand U13065 (N_13065,N_12952,N_12127);
nand U13066 (N_13066,N_12724,N_12233);
nand U13067 (N_13067,N_12226,N_12297);
and U13068 (N_13068,N_12925,N_12504);
and U13069 (N_13069,N_12442,N_12837);
xnor U13070 (N_13070,N_12308,N_12408);
and U13071 (N_13071,N_12053,N_12222);
and U13072 (N_13072,N_12886,N_12998);
and U13073 (N_13073,N_12964,N_12251);
or U13074 (N_13074,N_12664,N_12893);
xnor U13075 (N_13075,N_12396,N_12142);
nand U13076 (N_13076,N_12379,N_12521);
and U13077 (N_13077,N_12640,N_12281);
and U13078 (N_13078,N_12527,N_12227);
nor U13079 (N_13079,N_12021,N_12883);
xnor U13080 (N_13080,N_12581,N_12249);
and U13081 (N_13081,N_12156,N_12628);
nand U13082 (N_13082,N_12459,N_12237);
nor U13083 (N_13083,N_12242,N_12802);
nor U13084 (N_13084,N_12592,N_12300);
or U13085 (N_13085,N_12780,N_12180);
and U13086 (N_13086,N_12136,N_12389);
or U13087 (N_13087,N_12351,N_12686);
and U13088 (N_13088,N_12655,N_12203);
or U13089 (N_13089,N_12073,N_12130);
and U13090 (N_13090,N_12842,N_12068);
and U13091 (N_13091,N_12186,N_12063);
nand U13092 (N_13092,N_12283,N_12455);
nor U13093 (N_13093,N_12688,N_12928);
nor U13094 (N_13094,N_12210,N_12190);
xnor U13095 (N_13095,N_12432,N_12800);
nand U13096 (N_13096,N_12635,N_12361);
or U13097 (N_13097,N_12093,N_12639);
xor U13098 (N_13098,N_12608,N_12195);
or U13099 (N_13099,N_12828,N_12157);
nand U13100 (N_13100,N_12604,N_12914);
nor U13101 (N_13101,N_12338,N_12170);
or U13102 (N_13102,N_12427,N_12534);
and U13103 (N_13103,N_12487,N_12370);
or U13104 (N_13104,N_12584,N_12531);
or U13105 (N_13105,N_12910,N_12788);
and U13106 (N_13106,N_12057,N_12008);
nand U13107 (N_13107,N_12995,N_12637);
nor U13108 (N_13108,N_12003,N_12398);
or U13109 (N_13109,N_12731,N_12894);
xnor U13110 (N_13110,N_12857,N_12431);
nor U13111 (N_13111,N_12150,N_12784);
nand U13112 (N_13112,N_12179,N_12123);
or U13113 (N_13113,N_12164,N_12316);
nand U13114 (N_13114,N_12519,N_12774);
and U13115 (N_13115,N_12806,N_12245);
and U13116 (N_13116,N_12318,N_12451);
nor U13117 (N_13117,N_12327,N_12400);
nand U13118 (N_13118,N_12148,N_12097);
nor U13119 (N_13119,N_12787,N_12781);
xnor U13120 (N_13120,N_12735,N_12512);
or U13121 (N_13121,N_12942,N_12306);
nand U13122 (N_13122,N_12540,N_12552);
xor U13123 (N_13123,N_12869,N_12023);
nand U13124 (N_13124,N_12469,N_12610);
nand U13125 (N_13125,N_12493,N_12444);
nor U13126 (N_13126,N_12144,N_12270);
nand U13127 (N_13127,N_12567,N_12409);
nand U13128 (N_13128,N_12633,N_12443);
nor U13129 (N_13129,N_12054,N_12101);
or U13130 (N_13130,N_12456,N_12916);
and U13131 (N_13131,N_12213,N_12103);
and U13132 (N_13132,N_12197,N_12693);
nor U13133 (N_13133,N_12191,N_12031);
nor U13134 (N_13134,N_12183,N_12808);
nor U13135 (N_13135,N_12717,N_12376);
and U13136 (N_13136,N_12804,N_12106);
or U13137 (N_13137,N_12859,N_12683);
nor U13138 (N_13138,N_12090,N_12701);
and U13139 (N_13139,N_12539,N_12757);
nand U13140 (N_13140,N_12865,N_12937);
nor U13141 (N_13141,N_12507,N_12803);
or U13142 (N_13142,N_12078,N_12137);
nor U13143 (N_13143,N_12726,N_12834);
nor U13144 (N_13144,N_12571,N_12898);
nor U13145 (N_13145,N_12027,N_12069);
and U13146 (N_13146,N_12870,N_12301);
nand U13147 (N_13147,N_12618,N_12430);
and U13148 (N_13148,N_12377,N_12189);
or U13149 (N_13149,N_12680,N_12289);
or U13150 (N_13150,N_12687,N_12783);
nor U13151 (N_13151,N_12000,N_12771);
and U13152 (N_13152,N_12836,N_12510);
nand U13153 (N_13153,N_12768,N_12039);
or U13154 (N_13154,N_12173,N_12366);
nand U13155 (N_13155,N_12643,N_12541);
nand U13156 (N_13156,N_12450,N_12881);
and U13157 (N_13157,N_12614,N_12873);
or U13158 (N_13158,N_12401,N_12263);
nor U13159 (N_13159,N_12254,N_12866);
nand U13160 (N_13160,N_12232,N_12088);
and U13161 (N_13161,N_12234,N_12542);
or U13162 (N_13162,N_12632,N_12590);
nor U13163 (N_13163,N_12616,N_12081);
nor U13164 (N_13164,N_12681,N_12511);
or U13165 (N_13165,N_12296,N_12485);
or U13166 (N_13166,N_12307,N_12229);
or U13167 (N_13167,N_12984,N_12520);
nor U13168 (N_13168,N_12922,N_12566);
xnor U13169 (N_13169,N_12721,N_12706);
nand U13170 (N_13170,N_12187,N_12761);
or U13171 (N_13171,N_12949,N_12257);
nor U13172 (N_13172,N_12547,N_12832);
and U13173 (N_13173,N_12315,N_12966);
nor U13174 (N_13174,N_12611,N_12246);
and U13175 (N_13175,N_12907,N_12132);
nor U13176 (N_13176,N_12819,N_12872);
nand U13177 (N_13177,N_12736,N_12240);
and U13178 (N_13178,N_12812,N_12653);
or U13179 (N_13179,N_12041,N_12115);
nor U13180 (N_13180,N_12967,N_12012);
or U13181 (N_13181,N_12748,N_12248);
nand U13182 (N_13182,N_12154,N_12900);
or U13183 (N_13183,N_12714,N_12320);
and U13184 (N_13184,N_12391,N_12287);
or U13185 (N_13185,N_12631,N_12758);
or U13186 (N_13186,N_12921,N_12261);
or U13187 (N_13187,N_12058,N_12770);
nor U13188 (N_13188,N_12850,N_12434);
nor U13189 (N_13189,N_12357,N_12750);
or U13190 (N_13190,N_12587,N_12801);
xnor U13191 (N_13191,N_12669,N_12550);
nor U13192 (N_13192,N_12906,N_12988);
or U13193 (N_13193,N_12956,N_12040);
and U13194 (N_13194,N_12076,N_12772);
or U13195 (N_13195,N_12847,N_12209);
nor U13196 (N_13196,N_12742,N_12790);
nor U13197 (N_13197,N_12577,N_12050);
nand U13198 (N_13198,N_12982,N_12075);
nand U13199 (N_13199,N_12013,N_12007);
and U13200 (N_13200,N_12957,N_12252);
and U13201 (N_13201,N_12933,N_12538);
and U13202 (N_13202,N_12079,N_12562);
nor U13203 (N_13203,N_12702,N_12713);
nand U13204 (N_13204,N_12960,N_12323);
nand U13205 (N_13205,N_12374,N_12733);
and U13206 (N_13206,N_12536,N_12282);
and U13207 (N_13207,N_12972,N_12798);
and U13208 (N_13208,N_12015,N_12211);
or U13209 (N_13209,N_12259,N_12668);
or U13210 (N_13210,N_12671,N_12491);
and U13211 (N_13211,N_12626,N_12439);
nor U13212 (N_13212,N_12285,N_12716);
xor U13213 (N_13213,N_12018,N_12965);
and U13214 (N_13214,N_12350,N_12134);
nor U13215 (N_13215,N_12580,N_12488);
nand U13216 (N_13216,N_12697,N_12386);
or U13217 (N_13217,N_12727,N_12913);
or U13218 (N_13218,N_12606,N_12014);
or U13219 (N_13219,N_12061,N_12392);
nand U13220 (N_13220,N_12365,N_12452);
and U13221 (N_13221,N_12464,N_12029);
nand U13222 (N_13222,N_12912,N_12977);
nand U13223 (N_13223,N_12426,N_12677);
or U13224 (N_13224,N_12095,N_12763);
and U13225 (N_13225,N_12358,N_12822);
or U13226 (N_13226,N_12482,N_12656);
nand U13227 (N_13227,N_12414,N_12786);
nand U13228 (N_13228,N_12291,N_12709);
xor U13229 (N_13229,N_12208,N_12744);
and U13230 (N_13230,N_12268,N_12133);
and U13231 (N_13231,N_12385,N_12126);
nor U13232 (N_13232,N_12932,N_12182);
nor U13233 (N_13233,N_12124,N_12331);
nand U13234 (N_13234,N_12642,N_12553);
and U13235 (N_13235,N_12349,N_12831);
xnor U13236 (N_13236,N_12099,N_12080);
nor U13237 (N_13237,N_12650,N_12994);
nor U13238 (N_13238,N_12419,N_12368);
xor U13239 (N_13239,N_12255,N_12192);
nand U13240 (N_13240,N_12609,N_12929);
and U13241 (N_13241,N_12629,N_12448);
and U13242 (N_13242,N_12162,N_12936);
nand U13243 (N_13243,N_12117,N_12923);
or U13244 (N_13244,N_12845,N_12207);
nor U13245 (N_13245,N_12169,N_12561);
or U13246 (N_13246,N_12924,N_12699);
nand U13247 (N_13247,N_12935,N_12411);
or U13248 (N_13248,N_12644,N_12084);
and U13249 (N_13249,N_12286,N_12746);
nand U13250 (N_13250,N_12805,N_12889);
xnor U13251 (N_13251,N_12593,N_12612);
or U13252 (N_13252,N_12779,N_12712);
nor U13253 (N_13253,N_12390,N_12447);
nand U13254 (N_13254,N_12722,N_12983);
or U13255 (N_13255,N_12118,N_12321);
or U13256 (N_13256,N_12522,N_12465);
or U13257 (N_13257,N_12970,N_12293);
nor U13258 (N_13258,N_12313,N_12996);
and U13259 (N_13259,N_12544,N_12902);
or U13260 (N_13260,N_12342,N_12911);
nand U13261 (N_13261,N_12892,N_12104);
nand U13262 (N_13262,N_12861,N_12867);
nand U13263 (N_13263,N_12725,N_12918);
nor U13264 (N_13264,N_12613,N_12676);
and U13265 (N_13265,N_12138,N_12317);
or U13266 (N_13266,N_12505,N_12258);
or U13267 (N_13267,N_12202,N_12563);
xor U13268 (N_13268,N_12602,N_12344);
nand U13269 (N_13269,N_12454,N_12905);
nor U13270 (N_13270,N_12383,N_12749);
or U13271 (N_13271,N_12303,N_12298);
nor U13272 (N_13272,N_12974,N_12874);
or U13273 (N_13273,N_12340,N_12876);
nor U13274 (N_13274,N_12166,N_12559);
nand U13275 (N_13275,N_12589,N_12472);
nand U13276 (N_13276,N_12045,N_12468);
nand U13277 (N_13277,N_12858,N_12890);
and U13278 (N_13278,N_12940,N_12436);
nor U13279 (N_13279,N_12230,N_12460);
and U13280 (N_13280,N_12105,N_12359);
xor U13281 (N_13281,N_12690,N_12767);
nand U13282 (N_13282,N_12215,N_12155);
nand U13283 (N_13283,N_12060,N_12621);
nand U13284 (N_13284,N_12049,N_12011);
or U13285 (N_13285,N_12367,N_12585);
nand U13286 (N_13286,N_12659,N_12122);
nand U13287 (N_13287,N_12754,N_12955);
or U13288 (N_13288,N_12369,N_12194);
nand U13289 (N_13289,N_12030,N_12474);
nand U13290 (N_13290,N_12703,N_12641);
or U13291 (N_13291,N_12818,N_12695);
nor U13292 (N_13292,N_12871,N_12214);
xnor U13293 (N_13293,N_12555,N_12266);
nor U13294 (N_13294,N_12732,N_12603);
nand U13295 (N_13295,N_12794,N_12143);
and U13296 (N_13296,N_12930,N_12931);
or U13297 (N_13297,N_12708,N_12775);
or U13298 (N_13298,N_12751,N_12212);
and U13299 (N_13299,N_12206,N_12388);
nor U13300 (N_13300,N_12591,N_12275);
nand U13301 (N_13301,N_12403,N_12471);
nand U13302 (N_13302,N_12778,N_12262);
and U13303 (N_13303,N_12384,N_12738);
or U13304 (N_13304,N_12513,N_12453);
or U13305 (N_13305,N_12324,N_12583);
or U13306 (N_13306,N_12161,N_12537);
and U13307 (N_13307,N_12225,N_12181);
and U13308 (N_13308,N_12530,N_12116);
or U13309 (N_13309,N_12371,N_12880);
nor U13310 (N_13310,N_12991,N_12002);
xor U13311 (N_13311,N_12380,N_12326);
nor U13312 (N_13312,N_12868,N_12605);
nor U13313 (N_13313,N_12274,N_12265);
and U13314 (N_13314,N_12091,N_12153);
nor U13315 (N_13315,N_12711,N_12919);
and U13316 (N_13316,N_12071,N_12554);
nor U13317 (N_13317,N_12168,N_12958);
nor U13318 (N_13318,N_12685,N_12250);
and U13319 (N_13319,N_12743,N_12198);
nand U13320 (N_13320,N_12066,N_12347);
nor U13321 (N_13321,N_12826,N_12666);
nand U13322 (N_13322,N_12363,N_12393);
or U13323 (N_13323,N_12565,N_12895);
or U13324 (N_13324,N_12810,N_12445);
and U13325 (N_13325,N_12329,N_12236);
and U13326 (N_13326,N_12499,N_12177);
or U13327 (N_13327,N_12305,N_12997);
nor U13328 (N_13328,N_12747,N_12903);
or U13329 (N_13329,N_12947,N_12026);
or U13330 (N_13330,N_12601,N_12814);
nand U13331 (N_13331,N_12146,N_12109);
nand U13332 (N_13332,N_12862,N_12938);
nand U13333 (N_13333,N_12835,N_12791);
nor U13334 (N_13334,N_12193,N_12620);
nand U13335 (N_13335,N_12863,N_12364);
nand U13336 (N_13336,N_12896,N_12897);
and U13337 (N_13337,N_12915,N_12855);
nor U13338 (N_13338,N_12969,N_12473);
and U13339 (N_13339,N_12435,N_12558);
nand U13340 (N_13340,N_12477,N_12572);
nand U13341 (N_13341,N_12904,N_12336);
or U13342 (N_13342,N_12110,N_12820);
or U13343 (N_13343,N_12718,N_12843);
or U13344 (N_13344,N_12086,N_12528);
nand U13345 (N_13345,N_12158,N_12524);
and U13346 (N_13346,N_12545,N_12944);
and U13347 (N_13347,N_12789,N_12615);
nor U13348 (N_13348,N_12529,N_12851);
or U13349 (N_13349,N_12980,N_12399);
nor U13350 (N_13350,N_12328,N_12993);
or U13351 (N_13351,N_12028,N_12220);
nand U13352 (N_13352,N_12920,N_12648);
and U13353 (N_13353,N_12516,N_12551);
and U13354 (N_13354,N_12070,N_12089);
nand U13355 (N_13355,N_12188,N_12707);
nand U13356 (N_13356,N_12304,N_12087);
nor U13357 (N_13357,N_12102,N_12753);
nor U13358 (N_13358,N_12999,N_12574);
or U13359 (N_13359,N_12273,N_12424);
and U13360 (N_13360,N_12421,N_12333);
and U13361 (N_13361,N_12217,N_12486);
nand U13362 (N_13362,N_12548,N_12692);
or U13363 (N_13363,N_12492,N_12034);
nand U13364 (N_13364,N_12378,N_12264);
and U13365 (N_13365,N_12532,N_12277);
and U13366 (N_13366,N_12864,N_12759);
and U13367 (N_13367,N_12568,N_12446);
nand U13368 (N_13368,N_12276,N_12064);
or U13369 (N_13369,N_12394,N_12059);
nand U13370 (N_13370,N_12025,N_12151);
nor U13371 (N_13371,N_12457,N_12407);
xnor U13372 (N_13372,N_12490,N_12844);
nand U13373 (N_13373,N_12279,N_12672);
nand U13374 (N_13374,N_12796,N_12792);
nor U13375 (N_13375,N_12397,N_12120);
or U13376 (N_13376,N_12037,N_12284);
and U13377 (N_13377,N_12096,N_12055);
and U13378 (N_13378,N_12067,N_12627);
and U13379 (N_13379,N_12987,N_12082);
and U13380 (N_13380,N_12174,N_12839);
xor U13381 (N_13381,N_12645,N_12909);
xor U13382 (N_13382,N_12167,N_12730);
or U13383 (N_13383,N_12549,N_12546);
xor U13384 (N_13384,N_12495,N_12218);
xnor U13385 (N_13385,N_12413,N_12111);
or U13386 (N_13386,N_12311,N_12848);
nand U13387 (N_13387,N_12543,N_12777);
nand U13388 (N_13388,N_12518,N_12852);
or U13389 (N_13389,N_12231,N_12171);
and U13390 (N_13390,N_12253,N_12971);
or U13391 (N_13391,N_12985,N_12223);
nor U13392 (N_13392,N_12619,N_12048);
xnor U13393 (N_13393,N_12623,N_12663);
nand U13394 (N_13394,N_12417,N_12885);
and U13395 (N_13395,N_12934,N_12649);
nand U13396 (N_13396,N_12462,N_12526);
or U13397 (N_13397,N_12481,N_12705);
and U13398 (N_13398,N_12441,N_12785);
nand U13399 (N_13399,N_12001,N_12484);
xor U13400 (N_13400,N_12765,N_12299);
and U13401 (N_13401,N_12004,N_12636);
and U13402 (N_13402,N_12428,N_12598);
or U13403 (N_13403,N_12362,N_12943);
nor U13404 (N_13404,N_12322,N_12032);
and U13405 (N_13405,N_12739,N_12425);
and U13406 (N_13406,N_12901,N_12216);
and U13407 (N_13407,N_12467,N_12047);
and U13408 (N_13408,N_12175,N_12288);
nand U13409 (N_13409,N_12596,N_12698);
nand U13410 (N_13410,N_12269,N_12420);
or U13411 (N_13411,N_12121,N_12582);
or U13412 (N_13412,N_12821,N_12051);
or U13413 (N_13413,N_12147,N_12927);
nor U13414 (N_13414,N_12334,N_12975);
nand U13415 (N_13415,N_12402,N_12630);
xor U13416 (N_13416,N_12849,N_12908);
or U13417 (N_13417,N_12332,N_12163);
or U13418 (N_13418,N_12271,N_12853);
nand U13419 (N_13419,N_12508,N_12016);
nand U13420 (N_13420,N_12815,N_12302);
nor U13421 (N_13421,N_12201,N_12824);
nand U13422 (N_13422,N_12776,N_12319);
nand U13423 (N_13423,N_12496,N_12083);
nand U13424 (N_13424,N_12556,N_12599);
nand U13425 (N_13425,N_12205,N_12440);
nor U13426 (N_13426,N_12107,N_12092);
and U13427 (N_13427,N_12573,N_12239);
nor U13428 (N_13428,N_12085,N_12017);
nor U13429 (N_13429,N_12617,N_12244);
nand U13430 (N_13430,N_12348,N_12238);
and U13431 (N_13431,N_12178,N_12042);
and U13432 (N_13432,N_12119,N_12335);
or U13433 (N_13433,N_12962,N_12172);
and U13434 (N_13434,N_12479,N_12679);
nand U13435 (N_13435,N_12691,N_12145);
and U13436 (N_13436,N_12948,N_12108);
nor U13437 (N_13437,N_12159,N_12764);
nor U13438 (N_13438,N_12807,N_12463);
nor U13439 (N_13439,N_12887,N_12694);
or U13440 (N_13440,N_12523,N_12811);
nand U13441 (N_13441,N_12625,N_12797);
xnor U13442 (N_13442,N_12354,N_12939);
or U13443 (N_13443,N_12728,N_12280);
nand U13444 (N_13444,N_12899,N_12795);
nor U13445 (N_13445,N_12072,N_12480);
nand U13446 (N_13446,N_12219,N_12986);
or U13447 (N_13447,N_12470,N_12509);
nor U13448 (N_13448,N_12494,N_12945);
and U13449 (N_13449,N_12745,N_12235);
and U13450 (N_13450,N_12652,N_12501);
nand U13451 (N_13451,N_12314,N_12141);
and U13452 (N_13452,N_12741,N_12010);
and U13453 (N_13453,N_12833,N_12586);
or U13454 (N_13454,N_12782,N_12710);
or U13455 (N_13455,N_12310,N_12395);
nand U13456 (N_13456,N_12661,N_12769);
and U13457 (N_13457,N_12077,N_12737);
nand U13458 (N_13458,N_12221,N_12128);
nor U13459 (N_13459,N_12272,N_12588);
nand U13460 (N_13460,N_12422,N_12098);
nand U13461 (N_13461,N_12651,N_12294);
nand U13462 (N_13462,N_12139,N_12438);
or U13463 (N_13463,N_12449,N_12979);
and U13464 (N_13464,N_12723,N_12535);
nand U13465 (N_13465,N_12196,N_12860);
and U13466 (N_13466,N_12569,N_12799);
or U13467 (N_13467,N_12594,N_12667);
nor U13468 (N_13468,N_12959,N_12941);
nor U13469 (N_13469,N_12125,N_12670);
nor U13470 (N_13470,N_12415,N_12475);
nor U13471 (N_13471,N_12176,N_12044);
nand U13472 (N_13472,N_12793,N_12662);
and U13473 (N_13473,N_12184,N_12019);
and U13474 (N_13474,N_12817,N_12224);
nor U13475 (N_13475,N_12951,N_12149);
nand U13476 (N_13476,N_12729,N_12005);
nand U13477 (N_13477,N_12200,N_12437);
nor U13478 (N_13478,N_12657,N_12682);
nor U13479 (N_13479,N_12476,N_12950);
and U13480 (N_13480,N_12762,N_12888);
nor U13481 (N_13481,N_12696,N_12954);
nor U13482 (N_13482,N_12410,N_12752);
nand U13483 (N_13483,N_12309,N_12062);
and U13484 (N_13484,N_12500,N_12525);
nand U13485 (N_13485,N_12564,N_12946);
nand U13486 (N_13486,N_12891,N_12673);
nor U13487 (N_13487,N_12689,N_12953);
nand U13488 (N_13488,N_12152,N_12719);
nor U13489 (N_13489,N_12295,N_12074);
and U13490 (N_13490,N_12578,N_12458);
nand U13491 (N_13491,N_12241,N_12341);
and U13492 (N_13492,N_12700,N_12502);
and U13493 (N_13493,N_12129,N_12006);
xor U13494 (N_13494,N_12576,N_12678);
nor U13495 (N_13495,N_12404,N_12827);
nand U13496 (N_13496,N_12339,N_12740);
nor U13497 (N_13497,N_12917,N_12981);
nor U13498 (N_13498,N_12658,N_12356);
or U13499 (N_13499,N_12882,N_12461);
or U13500 (N_13500,N_12602,N_12135);
xnor U13501 (N_13501,N_12284,N_12922);
nand U13502 (N_13502,N_12088,N_12731);
nor U13503 (N_13503,N_12714,N_12863);
and U13504 (N_13504,N_12175,N_12633);
and U13505 (N_13505,N_12323,N_12026);
and U13506 (N_13506,N_12945,N_12673);
nand U13507 (N_13507,N_12717,N_12054);
nand U13508 (N_13508,N_12213,N_12333);
nor U13509 (N_13509,N_12691,N_12194);
nor U13510 (N_13510,N_12857,N_12544);
or U13511 (N_13511,N_12693,N_12116);
or U13512 (N_13512,N_12646,N_12295);
nor U13513 (N_13513,N_12415,N_12516);
or U13514 (N_13514,N_12509,N_12646);
or U13515 (N_13515,N_12989,N_12923);
xnor U13516 (N_13516,N_12912,N_12587);
nor U13517 (N_13517,N_12980,N_12745);
or U13518 (N_13518,N_12369,N_12840);
or U13519 (N_13519,N_12977,N_12790);
or U13520 (N_13520,N_12004,N_12184);
nor U13521 (N_13521,N_12971,N_12012);
xor U13522 (N_13522,N_12223,N_12267);
nor U13523 (N_13523,N_12433,N_12910);
xor U13524 (N_13524,N_12178,N_12029);
and U13525 (N_13525,N_12501,N_12688);
and U13526 (N_13526,N_12523,N_12711);
or U13527 (N_13527,N_12550,N_12622);
nor U13528 (N_13528,N_12767,N_12762);
xnor U13529 (N_13529,N_12759,N_12595);
or U13530 (N_13530,N_12100,N_12346);
and U13531 (N_13531,N_12445,N_12400);
and U13532 (N_13532,N_12336,N_12555);
nor U13533 (N_13533,N_12451,N_12436);
nor U13534 (N_13534,N_12146,N_12154);
nand U13535 (N_13535,N_12060,N_12249);
nand U13536 (N_13536,N_12216,N_12130);
nand U13537 (N_13537,N_12769,N_12463);
nor U13538 (N_13538,N_12945,N_12805);
and U13539 (N_13539,N_12168,N_12617);
and U13540 (N_13540,N_12051,N_12918);
or U13541 (N_13541,N_12338,N_12824);
and U13542 (N_13542,N_12843,N_12091);
and U13543 (N_13543,N_12018,N_12270);
nand U13544 (N_13544,N_12771,N_12005);
or U13545 (N_13545,N_12342,N_12463);
nand U13546 (N_13546,N_12287,N_12710);
or U13547 (N_13547,N_12309,N_12014);
xor U13548 (N_13548,N_12917,N_12763);
nand U13549 (N_13549,N_12054,N_12637);
or U13550 (N_13550,N_12845,N_12786);
nand U13551 (N_13551,N_12206,N_12817);
or U13552 (N_13552,N_12487,N_12666);
nand U13553 (N_13553,N_12756,N_12276);
nand U13554 (N_13554,N_12360,N_12801);
nand U13555 (N_13555,N_12513,N_12529);
xor U13556 (N_13556,N_12338,N_12482);
and U13557 (N_13557,N_12574,N_12732);
nand U13558 (N_13558,N_12781,N_12058);
nand U13559 (N_13559,N_12595,N_12154);
nor U13560 (N_13560,N_12438,N_12241);
or U13561 (N_13561,N_12638,N_12062);
or U13562 (N_13562,N_12836,N_12077);
xor U13563 (N_13563,N_12474,N_12363);
nand U13564 (N_13564,N_12392,N_12434);
nand U13565 (N_13565,N_12632,N_12941);
xor U13566 (N_13566,N_12969,N_12863);
nor U13567 (N_13567,N_12948,N_12414);
nor U13568 (N_13568,N_12965,N_12285);
or U13569 (N_13569,N_12184,N_12756);
and U13570 (N_13570,N_12968,N_12298);
and U13571 (N_13571,N_12232,N_12338);
or U13572 (N_13572,N_12255,N_12570);
nor U13573 (N_13573,N_12325,N_12282);
and U13574 (N_13574,N_12760,N_12141);
nand U13575 (N_13575,N_12624,N_12856);
or U13576 (N_13576,N_12374,N_12031);
nor U13577 (N_13577,N_12219,N_12302);
nor U13578 (N_13578,N_12884,N_12478);
and U13579 (N_13579,N_12487,N_12315);
xor U13580 (N_13580,N_12449,N_12089);
nor U13581 (N_13581,N_12887,N_12643);
nand U13582 (N_13582,N_12446,N_12639);
or U13583 (N_13583,N_12083,N_12051);
and U13584 (N_13584,N_12030,N_12014);
nor U13585 (N_13585,N_12190,N_12887);
xor U13586 (N_13586,N_12138,N_12521);
nand U13587 (N_13587,N_12531,N_12605);
or U13588 (N_13588,N_12437,N_12964);
nand U13589 (N_13589,N_12407,N_12937);
xor U13590 (N_13590,N_12100,N_12661);
nand U13591 (N_13591,N_12374,N_12601);
or U13592 (N_13592,N_12043,N_12465);
or U13593 (N_13593,N_12595,N_12631);
nor U13594 (N_13594,N_12798,N_12065);
nor U13595 (N_13595,N_12942,N_12153);
or U13596 (N_13596,N_12122,N_12101);
nand U13597 (N_13597,N_12719,N_12889);
and U13598 (N_13598,N_12694,N_12285);
nand U13599 (N_13599,N_12261,N_12680);
or U13600 (N_13600,N_12009,N_12063);
nor U13601 (N_13601,N_12519,N_12907);
nor U13602 (N_13602,N_12669,N_12922);
or U13603 (N_13603,N_12429,N_12821);
xor U13604 (N_13604,N_12000,N_12220);
nand U13605 (N_13605,N_12359,N_12680);
or U13606 (N_13606,N_12647,N_12849);
nand U13607 (N_13607,N_12440,N_12312);
or U13608 (N_13608,N_12366,N_12933);
nor U13609 (N_13609,N_12819,N_12837);
and U13610 (N_13610,N_12042,N_12627);
nand U13611 (N_13611,N_12897,N_12204);
nand U13612 (N_13612,N_12007,N_12212);
xor U13613 (N_13613,N_12987,N_12360);
and U13614 (N_13614,N_12944,N_12758);
and U13615 (N_13615,N_12802,N_12006);
and U13616 (N_13616,N_12878,N_12251);
nor U13617 (N_13617,N_12312,N_12894);
nand U13618 (N_13618,N_12109,N_12470);
nor U13619 (N_13619,N_12484,N_12397);
xnor U13620 (N_13620,N_12467,N_12864);
and U13621 (N_13621,N_12311,N_12303);
nand U13622 (N_13622,N_12895,N_12222);
xor U13623 (N_13623,N_12497,N_12564);
and U13624 (N_13624,N_12144,N_12640);
or U13625 (N_13625,N_12548,N_12292);
nor U13626 (N_13626,N_12939,N_12719);
xnor U13627 (N_13627,N_12168,N_12062);
and U13628 (N_13628,N_12239,N_12990);
or U13629 (N_13629,N_12680,N_12034);
and U13630 (N_13630,N_12514,N_12105);
nor U13631 (N_13631,N_12010,N_12736);
nor U13632 (N_13632,N_12880,N_12925);
or U13633 (N_13633,N_12488,N_12161);
and U13634 (N_13634,N_12954,N_12852);
nand U13635 (N_13635,N_12263,N_12918);
nor U13636 (N_13636,N_12887,N_12253);
and U13637 (N_13637,N_12454,N_12058);
and U13638 (N_13638,N_12021,N_12198);
nand U13639 (N_13639,N_12179,N_12830);
nor U13640 (N_13640,N_12099,N_12442);
nand U13641 (N_13641,N_12995,N_12319);
nand U13642 (N_13642,N_12830,N_12533);
and U13643 (N_13643,N_12786,N_12631);
nor U13644 (N_13644,N_12550,N_12485);
nor U13645 (N_13645,N_12490,N_12026);
or U13646 (N_13646,N_12475,N_12758);
or U13647 (N_13647,N_12463,N_12114);
or U13648 (N_13648,N_12164,N_12333);
or U13649 (N_13649,N_12184,N_12481);
and U13650 (N_13650,N_12158,N_12791);
or U13651 (N_13651,N_12674,N_12678);
or U13652 (N_13652,N_12876,N_12459);
and U13653 (N_13653,N_12446,N_12550);
nor U13654 (N_13654,N_12703,N_12086);
nand U13655 (N_13655,N_12835,N_12691);
and U13656 (N_13656,N_12867,N_12282);
nand U13657 (N_13657,N_12097,N_12453);
xor U13658 (N_13658,N_12775,N_12522);
nand U13659 (N_13659,N_12934,N_12251);
xnor U13660 (N_13660,N_12452,N_12811);
nand U13661 (N_13661,N_12223,N_12711);
or U13662 (N_13662,N_12628,N_12020);
nand U13663 (N_13663,N_12430,N_12820);
xnor U13664 (N_13664,N_12518,N_12748);
and U13665 (N_13665,N_12462,N_12004);
and U13666 (N_13666,N_12787,N_12874);
nor U13667 (N_13667,N_12625,N_12913);
nand U13668 (N_13668,N_12601,N_12796);
nor U13669 (N_13669,N_12303,N_12338);
nand U13670 (N_13670,N_12192,N_12797);
or U13671 (N_13671,N_12645,N_12376);
and U13672 (N_13672,N_12470,N_12687);
nand U13673 (N_13673,N_12308,N_12852);
or U13674 (N_13674,N_12286,N_12004);
or U13675 (N_13675,N_12087,N_12670);
nand U13676 (N_13676,N_12025,N_12618);
xor U13677 (N_13677,N_12077,N_12040);
nand U13678 (N_13678,N_12350,N_12925);
nor U13679 (N_13679,N_12496,N_12911);
or U13680 (N_13680,N_12404,N_12430);
xnor U13681 (N_13681,N_12602,N_12163);
or U13682 (N_13682,N_12330,N_12495);
or U13683 (N_13683,N_12830,N_12695);
and U13684 (N_13684,N_12035,N_12338);
and U13685 (N_13685,N_12638,N_12906);
nor U13686 (N_13686,N_12586,N_12446);
or U13687 (N_13687,N_12280,N_12823);
xnor U13688 (N_13688,N_12289,N_12179);
nor U13689 (N_13689,N_12638,N_12386);
and U13690 (N_13690,N_12255,N_12612);
nand U13691 (N_13691,N_12321,N_12962);
nand U13692 (N_13692,N_12181,N_12485);
or U13693 (N_13693,N_12131,N_12746);
or U13694 (N_13694,N_12703,N_12915);
and U13695 (N_13695,N_12007,N_12796);
and U13696 (N_13696,N_12925,N_12929);
or U13697 (N_13697,N_12839,N_12355);
or U13698 (N_13698,N_12540,N_12863);
nor U13699 (N_13699,N_12035,N_12024);
nand U13700 (N_13700,N_12625,N_12242);
or U13701 (N_13701,N_12372,N_12181);
nor U13702 (N_13702,N_12512,N_12000);
nor U13703 (N_13703,N_12010,N_12783);
nor U13704 (N_13704,N_12465,N_12797);
and U13705 (N_13705,N_12556,N_12716);
or U13706 (N_13706,N_12005,N_12829);
and U13707 (N_13707,N_12010,N_12213);
nand U13708 (N_13708,N_12055,N_12747);
nand U13709 (N_13709,N_12371,N_12790);
nor U13710 (N_13710,N_12852,N_12563);
xor U13711 (N_13711,N_12429,N_12965);
xnor U13712 (N_13712,N_12840,N_12215);
nand U13713 (N_13713,N_12491,N_12224);
and U13714 (N_13714,N_12785,N_12983);
nor U13715 (N_13715,N_12535,N_12048);
xor U13716 (N_13716,N_12893,N_12929);
nor U13717 (N_13717,N_12124,N_12600);
or U13718 (N_13718,N_12635,N_12661);
nand U13719 (N_13719,N_12637,N_12715);
and U13720 (N_13720,N_12413,N_12846);
nand U13721 (N_13721,N_12683,N_12942);
or U13722 (N_13722,N_12488,N_12674);
nand U13723 (N_13723,N_12447,N_12499);
nor U13724 (N_13724,N_12376,N_12027);
nor U13725 (N_13725,N_12975,N_12713);
and U13726 (N_13726,N_12645,N_12044);
nand U13727 (N_13727,N_12943,N_12098);
and U13728 (N_13728,N_12284,N_12156);
nand U13729 (N_13729,N_12050,N_12043);
and U13730 (N_13730,N_12629,N_12094);
and U13731 (N_13731,N_12625,N_12755);
and U13732 (N_13732,N_12967,N_12391);
nand U13733 (N_13733,N_12608,N_12924);
or U13734 (N_13734,N_12854,N_12674);
or U13735 (N_13735,N_12374,N_12589);
nor U13736 (N_13736,N_12019,N_12944);
xor U13737 (N_13737,N_12378,N_12889);
and U13738 (N_13738,N_12774,N_12133);
and U13739 (N_13739,N_12056,N_12699);
and U13740 (N_13740,N_12651,N_12122);
nand U13741 (N_13741,N_12236,N_12215);
or U13742 (N_13742,N_12862,N_12868);
nor U13743 (N_13743,N_12340,N_12001);
nor U13744 (N_13744,N_12417,N_12842);
or U13745 (N_13745,N_12345,N_12571);
and U13746 (N_13746,N_12235,N_12443);
nor U13747 (N_13747,N_12848,N_12068);
xor U13748 (N_13748,N_12003,N_12442);
nand U13749 (N_13749,N_12621,N_12894);
and U13750 (N_13750,N_12729,N_12647);
nor U13751 (N_13751,N_12933,N_12162);
nor U13752 (N_13752,N_12809,N_12337);
nor U13753 (N_13753,N_12330,N_12076);
nor U13754 (N_13754,N_12285,N_12687);
xnor U13755 (N_13755,N_12026,N_12107);
and U13756 (N_13756,N_12884,N_12745);
nor U13757 (N_13757,N_12011,N_12785);
and U13758 (N_13758,N_12924,N_12950);
or U13759 (N_13759,N_12465,N_12601);
or U13760 (N_13760,N_12313,N_12135);
nor U13761 (N_13761,N_12596,N_12548);
nand U13762 (N_13762,N_12595,N_12600);
or U13763 (N_13763,N_12400,N_12984);
nor U13764 (N_13764,N_12786,N_12815);
and U13765 (N_13765,N_12591,N_12236);
nor U13766 (N_13766,N_12048,N_12746);
nor U13767 (N_13767,N_12186,N_12244);
nor U13768 (N_13768,N_12582,N_12100);
or U13769 (N_13769,N_12202,N_12978);
nand U13770 (N_13770,N_12781,N_12355);
nor U13771 (N_13771,N_12304,N_12565);
or U13772 (N_13772,N_12647,N_12029);
or U13773 (N_13773,N_12138,N_12018);
xor U13774 (N_13774,N_12937,N_12593);
and U13775 (N_13775,N_12649,N_12048);
nor U13776 (N_13776,N_12887,N_12063);
and U13777 (N_13777,N_12485,N_12412);
nor U13778 (N_13778,N_12421,N_12968);
nand U13779 (N_13779,N_12967,N_12929);
nand U13780 (N_13780,N_12497,N_12649);
or U13781 (N_13781,N_12916,N_12705);
and U13782 (N_13782,N_12448,N_12013);
xor U13783 (N_13783,N_12344,N_12234);
nor U13784 (N_13784,N_12576,N_12515);
xnor U13785 (N_13785,N_12415,N_12321);
nand U13786 (N_13786,N_12605,N_12990);
nor U13787 (N_13787,N_12234,N_12389);
and U13788 (N_13788,N_12716,N_12034);
and U13789 (N_13789,N_12862,N_12779);
xor U13790 (N_13790,N_12398,N_12862);
and U13791 (N_13791,N_12677,N_12531);
nand U13792 (N_13792,N_12213,N_12221);
nor U13793 (N_13793,N_12811,N_12045);
xnor U13794 (N_13794,N_12401,N_12713);
and U13795 (N_13795,N_12961,N_12906);
and U13796 (N_13796,N_12661,N_12250);
xor U13797 (N_13797,N_12212,N_12320);
xor U13798 (N_13798,N_12481,N_12850);
or U13799 (N_13799,N_12320,N_12648);
nand U13800 (N_13800,N_12458,N_12779);
and U13801 (N_13801,N_12335,N_12218);
nor U13802 (N_13802,N_12735,N_12647);
nand U13803 (N_13803,N_12099,N_12955);
nor U13804 (N_13804,N_12191,N_12337);
and U13805 (N_13805,N_12283,N_12493);
nor U13806 (N_13806,N_12198,N_12142);
or U13807 (N_13807,N_12486,N_12990);
nand U13808 (N_13808,N_12339,N_12826);
or U13809 (N_13809,N_12615,N_12037);
and U13810 (N_13810,N_12520,N_12717);
or U13811 (N_13811,N_12133,N_12325);
nand U13812 (N_13812,N_12742,N_12021);
nor U13813 (N_13813,N_12949,N_12324);
nor U13814 (N_13814,N_12650,N_12136);
or U13815 (N_13815,N_12088,N_12746);
nand U13816 (N_13816,N_12051,N_12398);
nand U13817 (N_13817,N_12849,N_12617);
nand U13818 (N_13818,N_12559,N_12478);
xnor U13819 (N_13819,N_12842,N_12339);
nand U13820 (N_13820,N_12822,N_12728);
nand U13821 (N_13821,N_12724,N_12521);
and U13822 (N_13822,N_12032,N_12551);
xnor U13823 (N_13823,N_12000,N_12404);
nand U13824 (N_13824,N_12668,N_12252);
nand U13825 (N_13825,N_12397,N_12302);
and U13826 (N_13826,N_12628,N_12168);
or U13827 (N_13827,N_12199,N_12583);
nor U13828 (N_13828,N_12817,N_12871);
nor U13829 (N_13829,N_12879,N_12589);
nor U13830 (N_13830,N_12035,N_12067);
nor U13831 (N_13831,N_12296,N_12499);
nor U13832 (N_13832,N_12188,N_12026);
nand U13833 (N_13833,N_12072,N_12999);
or U13834 (N_13834,N_12717,N_12339);
nor U13835 (N_13835,N_12171,N_12229);
xor U13836 (N_13836,N_12804,N_12526);
nand U13837 (N_13837,N_12530,N_12234);
and U13838 (N_13838,N_12713,N_12131);
and U13839 (N_13839,N_12952,N_12733);
and U13840 (N_13840,N_12169,N_12660);
or U13841 (N_13841,N_12822,N_12960);
or U13842 (N_13842,N_12994,N_12524);
xor U13843 (N_13843,N_12250,N_12397);
xnor U13844 (N_13844,N_12902,N_12932);
or U13845 (N_13845,N_12093,N_12054);
xor U13846 (N_13846,N_12829,N_12625);
or U13847 (N_13847,N_12135,N_12218);
xnor U13848 (N_13848,N_12323,N_12169);
nor U13849 (N_13849,N_12779,N_12686);
nor U13850 (N_13850,N_12008,N_12271);
nor U13851 (N_13851,N_12106,N_12244);
or U13852 (N_13852,N_12841,N_12796);
nor U13853 (N_13853,N_12070,N_12530);
nand U13854 (N_13854,N_12414,N_12077);
or U13855 (N_13855,N_12307,N_12931);
or U13856 (N_13856,N_12440,N_12043);
or U13857 (N_13857,N_12867,N_12615);
nor U13858 (N_13858,N_12022,N_12312);
xor U13859 (N_13859,N_12629,N_12164);
nand U13860 (N_13860,N_12666,N_12347);
or U13861 (N_13861,N_12708,N_12020);
nor U13862 (N_13862,N_12825,N_12070);
nor U13863 (N_13863,N_12487,N_12883);
or U13864 (N_13864,N_12713,N_12324);
xor U13865 (N_13865,N_12381,N_12601);
nor U13866 (N_13866,N_12205,N_12341);
nor U13867 (N_13867,N_12384,N_12367);
or U13868 (N_13868,N_12652,N_12621);
and U13869 (N_13869,N_12747,N_12821);
and U13870 (N_13870,N_12239,N_12610);
and U13871 (N_13871,N_12238,N_12279);
and U13872 (N_13872,N_12820,N_12271);
or U13873 (N_13873,N_12844,N_12784);
or U13874 (N_13874,N_12196,N_12606);
and U13875 (N_13875,N_12622,N_12504);
and U13876 (N_13876,N_12945,N_12405);
and U13877 (N_13877,N_12147,N_12649);
nand U13878 (N_13878,N_12834,N_12590);
nand U13879 (N_13879,N_12892,N_12225);
and U13880 (N_13880,N_12142,N_12693);
nor U13881 (N_13881,N_12844,N_12804);
or U13882 (N_13882,N_12891,N_12684);
nand U13883 (N_13883,N_12933,N_12922);
and U13884 (N_13884,N_12468,N_12775);
nor U13885 (N_13885,N_12999,N_12729);
nor U13886 (N_13886,N_12852,N_12583);
xnor U13887 (N_13887,N_12879,N_12309);
nor U13888 (N_13888,N_12336,N_12996);
or U13889 (N_13889,N_12340,N_12096);
nor U13890 (N_13890,N_12148,N_12267);
or U13891 (N_13891,N_12817,N_12427);
nand U13892 (N_13892,N_12564,N_12513);
nor U13893 (N_13893,N_12521,N_12626);
and U13894 (N_13894,N_12224,N_12150);
nand U13895 (N_13895,N_12592,N_12660);
and U13896 (N_13896,N_12618,N_12549);
or U13897 (N_13897,N_12193,N_12386);
or U13898 (N_13898,N_12597,N_12579);
or U13899 (N_13899,N_12414,N_12967);
nand U13900 (N_13900,N_12194,N_12346);
nor U13901 (N_13901,N_12766,N_12313);
nand U13902 (N_13902,N_12304,N_12463);
nor U13903 (N_13903,N_12543,N_12610);
nor U13904 (N_13904,N_12686,N_12089);
nand U13905 (N_13905,N_12980,N_12145);
xor U13906 (N_13906,N_12735,N_12107);
nor U13907 (N_13907,N_12601,N_12265);
nor U13908 (N_13908,N_12168,N_12738);
xor U13909 (N_13909,N_12892,N_12720);
or U13910 (N_13910,N_12415,N_12904);
or U13911 (N_13911,N_12188,N_12233);
nand U13912 (N_13912,N_12977,N_12090);
nand U13913 (N_13913,N_12573,N_12765);
or U13914 (N_13914,N_12207,N_12960);
nor U13915 (N_13915,N_12888,N_12791);
nand U13916 (N_13916,N_12986,N_12033);
and U13917 (N_13917,N_12850,N_12798);
nor U13918 (N_13918,N_12739,N_12305);
or U13919 (N_13919,N_12759,N_12039);
nor U13920 (N_13920,N_12702,N_12789);
nand U13921 (N_13921,N_12343,N_12979);
xnor U13922 (N_13922,N_12623,N_12179);
and U13923 (N_13923,N_12368,N_12860);
or U13924 (N_13924,N_12392,N_12118);
and U13925 (N_13925,N_12613,N_12573);
xnor U13926 (N_13926,N_12680,N_12450);
or U13927 (N_13927,N_12209,N_12829);
nand U13928 (N_13928,N_12751,N_12098);
nand U13929 (N_13929,N_12225,N_12497);
nand U13930 (N_13930,N_12269,N_12976);
or U13931 (N_13931,N_12398,N_12087);
nor U13932 (N_13932,N_12994,N_12838);
nor U13933 (N_13933,N_12920,N_12197);
or U13934 (N_13934,N_12550,N_12667);
or U13935 (N_13935,N_12218,N_12972);
or U13936 (N_13936,N_12157,N_12218);
or U13937 (N_13937,N_12645,N_12726);
nor U13938 (N_13938,N_12609,N_12498);
nand U13939 (N_13939,N_12949,N_12095);
nand U13940 (N_13940,N_12640,N_12717);
nor U13941 (N_13941,N_12328,N_12421);
or U13942 (N_13942,N_12697,N_12118);
nand U13943 (N_13943,N_12966,N_12120);
and U13944 (N_13944,N_12699,N_12381);
or U13945 (N_13945,N_12707,N_12217);
nand U13946 (N_13946,N_12209,N_12589);
and U13947 (N_13947,N_12709,N_12889);
nor U13948 (N_13948,N_12213,N_12212);
nor U13949 (N_13949,N_12450,N_12034);
nand U13950 (N_13950,N_12448,N_12560);
nand U13951 (N_13951,N_12223,N_12997);
xor U13952 (N_13952,N_12163,N_12323);
nand U13953 (N_13953,N_12856,N_12371);
or U13954 (N_13954,N_12488,N_12496);
and U13955 (N_13955,N_12180,N_12322);
and U13956 (N_13956,N_12304,N_12134);
or U13957 (N_13957,N_12388,N_12565);
and U13958 (N_13958,N_12614,N_12793);
nand U13959 (N_13959,N_12111,N_12185);
nor U13960 (N_13960,N_12327,N_12676);
xor U13961 (N_13961,N_12433,N_12044);
and U13962 (N_13962,N_12332,N_12944);
nor U13963 (N_13963,N_12197,N_12051);
nor U13964 (N_13964,N_12786,N_12990);
nor U13965 (N_13965,N_12090,N_12718);
or U13966 (N_13966,N_12920,N_12866);
nand U13967 (N_13967,N_12793,N_12253);
xnor U13968 (N_13968,N_12946,N_12166);
nand U13969 (N_13969,N_12653,N_12254);
and U13970 (N_13970,N_12764,N_12174);
nand U13971 (N_13971,N_12119,N_12943);
and U13972 (N_13972,N_12148,N_12184);
nand U13973 (N_13973,N_12374,N_12432);
or U13974 (N_13974,N_12938,N_12298);
nor U13975 (N_13975,N_12643,N_12681);
xor U13976 (N_13976,N_12353,N_12029);
and U13977 (N_13977,N_12070,N_12744);
nor U13978 (N_13978,N_12629,N_12333);
nor U13979 (N_13979,N_12739,N_12355);
xor U13980 (N_13980,N_12366,N_12197);
nor U13981 (N_13981,N_12590,N_12023);
nand U13982 (N_13982,N_12754,N_12165);
nor U13983 (N_13983,N_12127,N_12441);
or U13984 (N_13984,N_12869,N_12134);
and U13985 (N_13985,N_12233,N_12471);
or U13986 (N_13986,N_12729,N_12340);
nor U13987 (N_13987,N_12926,N_12317);
and U13988 (N_13988,N_12336,N_12757);
nand U13989 (N_13989,N_12689,N_12414);
or U13990 (N_13990,N_12463,N_12095);
and U13991 (N_13991,N_12804,N_12735);
nor U13992 (N_13992,N_12452,N_12893);
nand U13993 (N_13993,N_12452,N_12096);
nor U13994 (N_13994,N_12357,N_12401);
or U13995 (N_13995,N_12375,N_12437);
xnor U13996 (N_13996,N_12637,N_12419);
nand U13997 (N_13997,N_12558,N_12678);
and U13998 (N_13998,N_12935,N_12969);
xnor U13999 (N_13999,N_12106,N_12201);
or U14000 (N_14000,N_13913,N_13814);
nand U14001 (N_14001,N_13616,N_13447);
xor U14002 (N_14002,N_13816,N_13439);
nor U14003 (N_14003,N_13080,N_13842);
and U14004 (N_14004,N_13098,N_13507);
nor U14005 (N_14005,N_13602,N_13810);
nand U14006 (N_14006,N_13496,N_13627);
nor U14007 (N_14007,N_13015,N_13948);
and U14008 (N_14008,N_13401,N_13093);
or U14009 (N_14009,N_13916,N_13407);
and U14010 (N_14010,N_13506,N_13620);
xnor U14011 (N_14011,N_13514,N_13185);
nor U14012 (N_14012,N_13357,N_13873);
nor U14013 (N_14013,N_13706,N_13188);
nand U14014 (N_14014,N_13542,N_13809);
nor U14015 (N_14015,N_13333,N_13575);
nor U14016 (N_14016,N_13885,N_13690);
or U14017 (N_14017,N_13298,N_13902);
or U14018 (N_14018,N_13246,N_13515);
and U14019 (N_14019,N_13009,N_13905);
nand U14020 (N_14020,N_13911,N_13623);
or U14021 (N_14021,N_13284,N_13405);
or U14022 (N_14022,N_13541,N_13451);
nor U14023 (N_14023,N_13326,N_13003);
xnor U14024 (N_14024,N_13356,N_13556);
xor U14025 (N_14025,N_13440,N_13625);
nor U14026 (N_14026,N_13638,N_13520);
nand U14027 (N_14027,N_13586,N_13239);
or U14028 (N_14028,N_13686,N_13685);
and U14029 (N_14029,N_13202,N_13938);
xnor U14030 (N_14030,N_13752,N_13632);
nor U14031 (N_14031,N_13151,N_13508);
and U14032 (N_14032,N_13473,N_13875);
or U14033 (N_14033,N_13497,N_13976);
nor U14034 (N_14034,N_13593,N_13245);
and U14035 (N_14035,N_13987,N_13466);
nand U14036 (N_14036,N_13846,N_13636);
nand U14037 (N_14037,N_13692,N_13789);
nand U14038 (N_14038,N_13524,N_13642);
and U14039 (N_14039,N_13805,N_13995);
nand U14040 (N_14040,N_13844,N_13768);
nand U14041 (N_14041,N_13989,N_13621);
nand U14042 (N_14042,N_13014,N_13582);
and U14043 (N_14043,N_13088,N_13445);
nor U14044 (N_14044,N_13662,N_13584);
nand U14045 (N_14045,N_13763,N_13571);
nor U14046 (N_14046,N_13229,N_13078);
or U14047 (N_14047,N_13269,N_13173);
and U14048 (N_14048,N_13598,N_13589);
and U14049 (N_14049,N_13489,N_13937);
nor U14050 (N_14050,N_13635,N_13176);
and U14051 (N_14051,N_13831,N_13566);
or U14052 (N_14052,N_13106,N_13544);
and U14053 (N_14053,N_13626,N_13950);
nor U14054 (N_14054,N_13067,N_13784);
nor U14055 (N_14055,N_13209,N_13683);
nor U14056 (N_14056,N_13069,N_13155);
nor U14057 (N_14057,N_13214,N_13211);
or U14058 (N_14058,N_13167,N_13526);
nand U14059 (N_14059,N_13231,N_13296);
nor U14060 (N_14060,N_13047,N_13083);
and U14061 (N_14061,N_13787,N_13999);
xor U14062 (N_14062,N_13591,N_13415);
or U14063 (N_14063,N_13222,N_13745);
or U14064 (N_14064,N_13827,N_13652);
nand U14065 (N_14065,N_13131,N_13878);
or U14066 (N_14066,N_13534,N_13278);
nand U14067 (N_14067,N_13917,N_13133);
and U14068 (N_14068,N_13693,N_13302);
nor U14069 (N_14069,N_13578,N_13321);
and U14070 (N_14070,N_13247,N_13882);
nor U14071 (N_14071,N_13871,N_13852);
xor U14072 (N_14072,N_13157,N_13117);
nand U14073 (N_14073,N_13528,N_13741);
or U14074 (N_14074,N_13703,N_13694);
or U14075 (N_14075,N_13747,N_13709);
nand U14076 (N_14076,N_13596,N_13316);
and U14077 (N_14077,N_13114,N_13656);
nor U14078 (N_14078,N_13863,N_13272);
nand U14079 (N_14079,N_13590,N_13144);
nand U14080 (N_14080,N_13370,N_13314);
and U14081 (N_14081,N_13287,N_13251);
xnor U14082 (N_14082,N_13695,N_13874);
or U14083 (N_14083,N_13998,N_13957);
nand U14084 (N_14084,N_13647,N_13881);
nand U14085 (N_14085,N_13261,N_13471);
nand U14086 (N_14086,N_13487,N_13563);
and U14087 (N_14087,N_13672,N_13033);
or U14088 (N_14088,N_13315,N_13353);
or U14089 (N_14089,N_13066,N_13048);
nand U14090 (N_14090,N_13644,N_13630);
or U14091 (N_14091,N_13103,N_13944);
xnor U14092 (N_14092,N_13488,N_13348);
nor U14093 (N_14093,N_13062,N_13412);
nand U14094 (N_14094,N_13354,N_13901);
or U14095 (N_14095,N_13076,N_13979);
and U14096 (N_14096,N_13678,N_13132);
and U14097 (N_14097,N_13404,N_13297);
nand U14098 (N_14098,N_13539,N_13158);
nor U14099 (N_14099,N_13500,N_13702);
or U14100 (N_14100,N_13442,N_13855);
nand U14101 (N_14101,N_13565,N_13713);
nor U14102 (N_14102,N_13474,N_13007);
nand U14103 (N_14103,N_13603,N_13365);
nand U14104 (N_14104,N_13559,N_13380);
nand U14105 (N_14105,N_13955,N_13966);
nor U14106 (N_14106,N_13569,N_13854);
and U14107 (N_14107,N_13336,N_13414);
nor U14108 (N_14108,N_13910,N_13480);
nand U14109 (N_14109,N_13241,N_13537);
nor U14110 (N_14110,N_13026,N_13041);
or U14111 (N_14111,N_13772,N_13425);
nand U14112 (N_14112,N_13079,N_13084);
or U14113 (N_14113,N_13605,N_13096);
nor U14114 (N_14114,N_13051,N_13243);
nand U14115 (N_14115,N_13043,N_13344);
xnor U14116 (N_14116,N_13734,N_13729);
and U14117 (N_14117,N_13207,N_13866);
nand U14118 (N_14118,N_13481,N_13583);
and U14119 (N_14119,N_13639,N_13149);
nand U14120 (N_14120,N_13485,N_13705);
and U14121 (N_14121,N_13651,N_13509);
and U14122 (N_14122,N_13483,N_13351);
xor U14123 (N_14123,N_13720,N_13056);
nand U14124 (N_14124,N_13749,N_13286);
or U14125 (N_14125,N_13118,N_13794);
and U14126 (N_14126,N_13002,N_13965);
xor U14127 (N_14127,N_13939,N_13545);
or U14128 (N_14128,N_13894,N_13925);
and U14129 (N_14129,N_13028,N_13889);
nand U14130 (N_14130,N_13199,N_13535);
and U14131 (N_14131,N_13073,N_13850);
nor U14132 (N_14132,N_13654,N_13463);
nor U14133 (N_14133,N_13250,N_13550);
nor U14134 (N_14134,N_13477,N_13232);
nor U14135 (N_14135,N_13862,N_13663);
nand U14136 (N_14136,N_13266,N_13484);
or U14137 (N_14137,N_13162,N_13853);
or U14138 (N_14138,N_13601,N_13869);
nor U14139 (N_14139,N_13826,N_13576);
nand U14140 (N_14140,N_13494,N_13818);
nand U14141 (N_14141,N_13519,N_13137);
or U14142 (N_14142,N_13588,N_13505);
xor U14143 (N_14143,N_13437,N_13270);
nor U14144 (N_14144,N_13413,N_13371);
and U14145 (N_14145,N_13152,N_13666);
and U14146 (N_14146,N_13472,N_13930);
nand U14147 (N_14147,N_13951,N_13529);
nand U14148 (N_14148,N_13574,N_13629);
nand U14149 (N_14149,N_13070,N_13547);
nor U14150 (N_14150,N_13608,N_13912);
and U14151 (N_14151,N_13641,N_13971);
and U14152 (N_14152,N_13019,N_13216);
or U14153 (N_14153,N_13521,N_13455);
xor U14154 (N_14154,N_13517,N_13097);
xnor U14155 (N_14155,N_13113,N_13184);
and U14156 (N_14156,N_13478,N_13935);
nand U14157 (N_14157,N_13461,N_13735);
nand U14158 (N_14158,N_13962,N_13397);
nand U14159 (N_14159,N_13991,N_13345);
nor U14160 (N_14160,N_13701,N_13774);
or U14161 (N_14161,N_13819,N_13967);
nor U14162 (N_14162,N_13154,N_13392);
nand U14163 (N_14163,N_13503,N_13631);
nand U14164 (N_14164,N_13587,N_13406);
and U14165 (N_14165,N_13281,N_13125);
nor U14166 (N_14166,N_13884,N_13408);
nor U14167 (N_14167,N_13646,N_13218);
or U14168 (N_14168,N_13004,N_13759);
and U14169 (N_14169,N_13420,N_13432);
nor U14170 (N_14170,N_13227,N_13904);
xor U14171 (N_14171,N_13023,N_13769);
nand U14172 (N_14172,N_13259,N_13754);
nor U14173 (N_14173,N_13704,N_13822);
nor U14174 (N_14174,N_13021,N_13548);
or U14175 (N_14175,N_13361,N_13201);
xor U14176 (N_14176,N_13757,N_13148);
nor U14177 (N_14177,N_13766,N_13712);
nand U14178 (N_14178,N_13134,N_13783);
nand U14179 (N_14179,N_13640,N_13867);
nor U14180 (N_14180,N_13311,N_13553);
xor U14181 (N_14181,N_13358,N_13612);
and U14182 (N_14182,N_13419,N_13391);
or U14183 (N_14183,N_13244,N_13659);
nand U14184 (N_14184,N_13436,N_13318);
and U14185 (N_14185,N_13428,N_13441);
nor U14186 (N_14186,N_13776,N_13551);
and U14187 (N_14187,N_13755,N_13087);
or U14188 (N_14188,N_13613,N_13464);
nand U14189 (N_14189,N_13057,N_13614);
xnor U14190 (N_14190,N_13561,N_13634);
nor U14191 (N_14191,N_13619,N_13332);
and U14192 (N_14192,N_13168,N_13674);
nor U14193 (N_14193,N_13249,N_13238);
nand U14194 (N_14194,N_13011,N_13200);
nand U14195 (N_14195,N_13458,N_13327);
or U14196 (N_14196,N_13914,N_13271);
nor U14197 (N_14197,N_13624,N_13510);
and U14198 (N_14198,N_13949,N_13960);
and U14199 (N_14199,N_13372,N_13929);
nor U14200 (N_14200,N_13411,N_13276);
nand U14201 (N_14201,N_13970,N_13123);
and U14202 (N_14202,N_13675,N_13525);
and U14203 (N_14203,N_13511,N_13398);
nand U14204 (N_14204,N_13549,N_13851);
nand U14205 (N_14205,N_13434,N_13174);
nand U14206 (N_14206,N_13217,N_13920);
nand U14207 (N_14207,N_13126,N_13068);
nand U14208 (N_14208,N_13600,N_13710);
or U14209 (N_14209,N_13277,N_13400);
nand U14210 (N_14210,N_13812,N_13791);
or U14211 (N_14211,N_13191,N_13359);
and U14212 (N_14212,N_13845,N_13963);
xor U14213 (N_14213,N_13403,N_13116);
nor U14214 (N_14214,N_13758,N_13292);
nand U14215 (N_14215,N_13653,N_13060);
and U14216 (N_14216,N_13982,N_13182);
and U14217 (N_14217,N_13807,N_13504);
nor U14218 (N_14218,N_13546,N_13981);
or U14219 (N_14219,N_13773,N_13921);
or U14220 (N_14220,N_13954,N_13252);
nand U14221 (N_14221,N_13990,N_13648);
nand U14222 (N_14222,N_13145,N_13977);
nor U14223 (N_14223,N_13804,N_13102);
or U14224 (N_14224,N_13823,N_13645);
xor U14225 (N_14225,N_13039,N_13595);
or U14226 (N_14226,N_13150,N_13908);
and U14227 (N_14227,N_13670,N_13604);
and U14228 (N_14228,N_13376,N_13760);
xnor U14229 (N_14229,N_13291,N_13307);
or U14230 (N_14230,N_13597,N_13175);
nor U14231 (N_14231,N_13898,N_13988);
or U14232 (N_14232,N_13147,N_13491);
nor U14233 (N_14233,N_13196,N_13897);
or U14234 (N_14234,N_13101,N_13020);
or U14235 (N_14235,N_13085,N_13045);
xor U14236 (N_14236,N_13655,N_13649);
nor U14237 (N_14237,N_13708,N_13585);
nand U14238 (N_14238,N_13936,N_13718);
or U14239 (N_14239,N_13953,N_13499);
nand U14240 (N_14240,N_13219,N_13817);
xnor U14241 (N_14241,N_13793,N_13426);
nand U14242 (N_14242,N_13091,N_13857);
xor U14243 (N_14243,N_13849,N_13082);
xnor U14244 (N_14244,N_13355,N_13205);
nand U14245 (N_14245,N_13049,N_13985);
nor U14246 (N_14246,N_13388,N_13288);
and U14247 (N_14247,N_13622,N_13443);
nor U14248 (N_14248,N_13864,N_13927);
and U14249 (N_14249,N_13731,N_13036);
xor U14250 (N_14250,N_13055,N_13334);
and U14251 (N_14251,N_13206,N_13115);
and U14252 (N_14252,N_13204,N_13417);
and U14253 (N_14253,N_13470,N_13740);
and U14254 (N_14254,N_13153,N_13861);
or U14255 (N_14255,N_13267,N_13340);
nand U14256 (N_14256,N_13299,N_13254);
nand U14257 (N_14257,N_13761,N_13260);
nand U14258 (N_14258,N_13637,N_13012);
nand U14259 (N_14259,N_13446,N_13808);
or U14260 (N_14260,N_13468,N_13942);
nor U14261 (N_14261,N_13300,N_13554);
nor U14262 (N_14262,N_13431,N_13959);
and U14263 (N_14263,N_13138,N_13492);
nor U14264 (N_14264,N_13567,N_13194);
nor U14265 (N_14265,N_13592,N_13657);
or U14266 (N_14266,N_13847,N_13617);
xor U14267 (N_14267,N_13746,N_13786);
or U14268 (N_14268,N_13696,N_13453);
nor U14269 (N_14269,N_13972,N_13337);
and U14270 (N_14270,N_13378,N_13285);
and U14271 (N_14271,N_13581,N_13189);
nor U14272 (N_14272,N_13280,N_13715);
nor U14273 (N_14273,N_13975,N_13399);
nor U14274 (N_14274,N_13161,N_13226);
and U14275 (N_14275,N_13518,N_13555);
nand U14276 (N_14276,N_13890,N_13486);
nor U14277 (N_14277,N_13723,N_13865);
and U14278 (N_14278,N_13628,N_13532);
and U14279 (N_14279,N_13140,N_13738);
nand U14280 (N_14280,N_13177,N_13046);
or U14281 (N_14281,N_13329,N_13389);
nand U14282 (N_14282,N_13658,N_13018);
nand U14283 (N_14283,N_13516,N_13611);
nand U14284 (N_14284,N_13859,N_13006);
nand U14285 (N_14285,N_13824,N_13368);
nand U14286 (N_14286,N_13512,N_13751);
or U14287 (N_14287,N_13108,N_13557);
and U14288 (N_14288,N_13034,N_13837);
nor U14289 (N_14289,N_13562,N_13689);
nor U14290 (N_14290,N_13171,N_13893);
or U14291 (N_14291,N_13700,N_13390);
and U14292 (N_14292,N_13086,N_13536);
nor U14293 (N_14293,N_13213,N_13843);
or U14294 (N_14294,N_13900,N_13811);
nand U14295 (N_14295,N_13796,N_13730);
nor U14296 (N_14296,N_13792,N_13531);
and U14297 (N_14297,N_13952,N_13465);
or U14298 (N_14298,N_13107,N_13430);
or U14299 (N_14299,N_13899,N_13170);
or U14300 (N_14300,N_13264,N_13120);
or U14301 (N_14301,N_13552,N_13779);
nand U14302 (N_14302,N_13139,N_13956);
nor U14303 (N_14303,N_13221,N_13934);
and U14304 (N_14304,N_13215,N_13037);
xnor U14305 (N_14305,N_13384,N_13253);
nor U14306 (N_14306,N_13172,N_13691);
nor U14307 (N_14307,N_13416,N_13886);
nand U14308 (N_14308,N_13328,N_13178);
and U14309 (N_14309,N_13360,N_13887);
nor U14310 (N_14310,N_13423,N_13347);
xor U14311 (N_14311,N_13947,N_13858);
nand U14312 (N_14312,N_13223,N_13829);
nand U14313 (N_14313,N_13274,N_13909);
and U14314 (N_14314,N_13788,N_13748);
and U14315 (N_14315,N_13984,N_13742);
nand U14316 (N_14316,N_13257,N_13717);
nand U14317 (N_14317,N_13522,N_13782);
nand U14318 (N_14318,N_13928,N_13072);
nand U14319 (N_14319,N_13462,N_13933);
and U14320 (N_14320,N_13109,N_13444);
nor U14321 (N_14321,N_13615,N_13836);
nor U14322 (N_14322,N_13094,N_13313);
or U14323 (N_14323,N_13127,N_13838);
and U14324 (N_14324,N_13183,N_13737);
or U14325 (N_14325,N_13719,N_13306);
and U14326 (N_14326,N_13000,N_13090);
and U14327 (N_14327,N_13130,N_13310);
and U14328 (N_14328,N_13821,N_13568);
nor U14329 (N_14329,N_13833,N_13100);
xor U14330 (N_14330,N_13242,N_13181);
nand U14331 (N_14331,N_13490,N_13476);
nor U14332 (N_14332,N_13095,N_13338);
or U14333 (N_14333,N_13017,N_13262);
or U14334 (N_14334,N_13643,N_13008);
and U14335 (N_14335,N_13771,N_13876);
nand U14336 (N_14336,N_13610,N_13753);
nor U14337 (N_14337,N_13452,N_13053);
and U14338 (N_14338,N_13165,N_13235);
and U14339 (N_14339,N_13688,N_13739);
nor U14340 (N_14340,N_13743,N_13558);
or U14341 (N_14341,N_13770,N_13330);
and U14342 (N_14342,N_13728,N_13427);
or U14343 (N_14343,N_13190,N_13606);
xnor U14344 (N_14344,N_13350,N_13124);
nor U14345 (N_14345,N_13295,N_13732);
nor U14346 (N_14346,N_13042,N_13467);
nand U14347 (N_14347,N_13092,N_13830);
nor U14348 (N_14348,N_13958,N_13377);
nor U14349 (N_14349,N_13156,N_13099);
and U14350 (N_14350,N_13393,N_13044);
and U14351 (N_14351,N_13832,N_13931);
and U14352 (N_14352,N_13339,N_13025);
nor U14353 (N_14353,N_13744,N_13128);
nand U14354 (N_14354,N_13993,N_13322);
or U14355 (N_14355,N_13454,N_13650);
or U14356 (N_14356,N_13104,N_13841);
nor U14357 (N_14357,N_13698,N_13924);
nand U14358 (N_14358,N_13711,N_13785);
nor U14359 (N_14359,N_13860,N_13422);
or U14360 (N_14360,N_13580,N_13164);
nor U14361 (N_14361,N_13179,N_13594);
nor U14362 (N_14362,N_13840,N_13237);
nor U14363 (N_14363,N_13325,N_13892);
nand U14364 (N_14364,N_13077,N_13800);
and U14365 (N_14365,N_13736,N_13290);
and U14366 (N_14366,N_13402,N_13362);
nor U14367 (N_14367,N_13880,N_13180);
or U14368 (N_14368,N_13667,N_13081);
nor U14369 (N_14369,N_13320,N_13996);
xnor U14370 (N_14370,N_13828,N_13501);
nor U14371 (N_14371,N_13727,N_13224);
or U14372 (N_14372,N_13961,N_13112);
nand U14373 (N_14373,N_13677,N_13721);
and U14374 (N_14374,N_13697,N_13105);
or U14375 (N_14375,N_13110,N_13054);
and U14376 (N_14376,N_13803,N_13543);
and U14377 (N_14377,N_13038,N_13294);
xor U14378 (N_14378,N_13946,N_13386);
nor U14379 (N_14379,N_13383,N_13756);
nor U14380 (N_14380,N_13680,N_13834);
or U14381 (N_14381,N_13983,N_13456);
or U14382 (N_14382,N_13293,N_13230);
nor U14383 (N_14383,N_13074,N_13136);
or U14384 (N_14384,N_13312,N_13573);
or U14385 (N_14385,N_13363,N_13027);
xor U14386 (N_14386,N_13208,N_13064);
and U14387 (N_14387,N_13795,N_13579);
or U14388 (N_14388,N_13806,N_13121);
and U14389 (N_14389,N_13160,N_13319);
or U14390 (N_14390,N_13513,N_13323);
nand U14391 (N_14391,N_13815,N_13945);
or U14392 (N_14392,N_13040,N_13324);
or U14393 (N_14393,N_13052,N_13146);
nand U14394 (N_14394,N_13379,N_13716);
or U14395 (N_14395,N_13063,N_13781);
xnor U14396 (N_14396,N_13263,N_13331);
nand U14397 (N_14397,N_13410,N_13289);
nor U14398 (N_14398,N_13367,N_13777);
nand U14399 (N_14399,N_13059,N_13891);
nor U14400 (N_14400,N_13801,N_13335);
or U14401 (N_14401,N_13964,N_13304);
and U14402 (N_14402,N_13203,N_13381);
nor U14403 (N_14403,N_13024,N_13013);
nor U14404 (N_14404,N_13778,N_13839);
or U14405 (N_14405,N_13031,N_13725);
nand U14406 (N_14406,N_13256,N_13618);
or U14407 (N_14407,N_13058,N_13065);
and U14408 (N_14408,N_13016,N_13450);
and U14409 (N_14409,N_13119,N_13906);
or U14410 (N_14410,N_13926,N_13883);
xnor U14411 (N_14411,N_13978,N_13980);
or U14412 (N_14412,N_13868,N_13479);
or U14413 (N_14413,N_13343,N_13714);
and U14414 (N_14414,N_13540,N_13560);
xor U14415 (N_14415,N_13309,N_13679);
nand U14416 (N_14416,N_13767,N_13341);
and U14417 (N_14417,N_13820,N_13159);
and U14418 (N_14418,N_13699,N_13502);
or U14419 (N_14419,N_13915,N_13475);
and U14420 (N_14420,N_13240,N_13660);
xnor U14421 (N_14421,N_13438,N_13283);
nand U14422 (N_14422,N_13969,N_13523);
nand U14423 (N_14423,N_13308,N_13364);
and U14424 (N_14424,N_13918,N_13071);
nor U14425 (N_14425,N_13448,N_13870);
nor U14426 (N_14426,N_13802,N_13396);
and U14427 (N_14427,N_13236,N_13141);
and U14428 (N_14428,N_13225,N_13061);
and U14429 (N_14429,N_13197,N_13193);
and U14430 (N_14430,N_13366,N_13352);
nor U14431 (N_14431,N_13301,N_13907);
xor U14432 (N_14432,N_13192,N_13564);
nor U14433 (N_14433,N_13668,N_13879);
nor U14434 (N_14434,N_13922,N_13687);
nor U14435 (N_14435,N_13848,N_13421);
xor U14436 (N_14436,N_13813,N_13665);
nor U14437 (N_14437,N_13780,N_13943);
or U14438 (N_14438,N_13233,N_13268);
nor U14439 (N_14439,N_13111,N_13382);
and U14440 (N_14440,N_13765,N_13375);
nor U14441 (N_14441,N_13273,N_13527);
nand U14442 (N_14442,N_13409,N_13533);
nand U14443 (N_14443,N_13135,N_13373);
nand U14444 (N_14444,N_13530,N_13258);
xnor U14445 (N_14445,N_13633,N_13968);
or U14446 (N_14446,N_13129,N_13460);
nand U14447 (N_14447,N_13986,N_13495);
nand U14448 (N_14448,N_13387,N_13493);
nand U14449 (N_14449,N_13724,N_13895);
xor U14450 (N_14450,N_13940,N_13248);
nand U14451 (N_14451,N_13609,N_13143);
nor U14452 (N_14452,N_13265,N_13877);
xor U14453 (N_14453,N_13825,N_13570);
or U14454 (N_14454,N_13349,N_13255);
or U14455 (N_14455,N_13676,N_13435);
and U14456 (N_14456,N_13195,N_13210);
nor U14457 (N_14457,N_13305,N_13682);
nand U14458 (N_14458,N_13346,N_13684);
or U14459 (N_14459,N_13459,N_13726);
nor U14460 (N_14460,N_13166,N_13722);
and U14461 (N_14461,N_13992,N_13856);
nor U14462 (N_14462,N_13664,N_13790);
and U14463 (N_14463,N_13764,N_13029);
nand U14464 (N_14464,N_13835,N_13896);
or U14465 (N_14465,N_13799,N_13449);
xor U14466 (N_14466,N_13941,N_13394);
nand U14467 (N_14467,N_13498,N_13279);
nor U14468 (N_14468,N_13457,N_13607);
and U14469 (N_14469,N_13903,N_13212);
xnor U14470 (N_14470,N_13797,N_13282);
nor U14471 (N_14471,N_13035,N_13923);
nor U14472 (N_14472,N_13198,N_13385);
or U14473 (N_14473,N_13186,N_13707);
or U14474 (N_14474,N_13775,N_13997);
nand U14475 (N_14475,N_13163,N_13872);
or U14476 (N_14476,N_13994,N_13001);
nand U14477 (N_14477,N_13469,N_13973);
and U14478 (N_14478,N_13673,N_13228);
xnor U14479 (N_14479,N_13538,N_13418);
nand U14480 (N_14480,N_13932,N_13169);
or U14481 (N_14481,N_13220,N_13888);
xnor U14482 (N_14482,N_13661,N_13681);
or U14483 (N_14483,N_13733,N_13303);
nand U14484 (N_14484,N_13374,N_13599);
and U14485 (N_14485,N_13142,N_13433);
nor U14486 (N_14486,N_13750,N_13030);
nor U14487 (N_14487,N_13075,N_13424);
and U14488 (N_14488,N_13234,N_13317);
or U14489 (N_14489,N_13010,N_13572);
nand U14490 (N_14490,N_13395,N_13050);
and U14491 (N_14491,N_13577,N_13369);
or U14492 (N_14492,N_13005,N_13187);
xor U14493 (N_14493,N_13429,N_13669);
nand U14494 (N_14494,N_13762,N_13974);
nand U14495 (N_14495,N_13089,N_13671);
nor U14496 (N_14496,N_13022,N_13919);
and U14497 (N_14497,N_13798,N_13275);
or U14498 (N_14498,N_13482,N_13032);
or U14499 (N_14499,N_13342,N_13122);
nor U14500 (N_14500,N_13542,N_13165);
nor U14501 (N_14501,N_13013,N_13915);
nor U14502 (N_14502,N_13432,N_13684);
nor U14503 (N_14503,N_13106,N_13172);
nand U14504 (N_14504,N_13673,N_13250);
xnor U14505 (N_14505,N_13084,N_13729);
or U14506 (N_14506,N_13162,N_13303);
nand U14507 (N_14507,N_13586,N_13871);
xor U14508 (N_14508,N_13886,N_13191);
nand U14509 (N_14509,N_13515,N_13731);
nor U14510 (N_14510,N_13967,N_13629);
nor U14511 (N_14511,N_13824,N_13700);
or U14512 (N_14512,N_13928,N_13198);
and U14513 (N_14513,N_13860,N_13754);
xnor U14514 (N_14514,N_13150,N_13210);
xor U14515 (N_14515,N_13093,N_13431);
xnor U14516 (N_14516,N_13193,N_13669);
nand U14517 (N_14517,N_13813,N_13364);
and U14518 (N_14518,N_13602,N_13249);
nand U14519 (N_14519,N_13223,N_13290);
nor U14520 (N_14520,N_13897,N_13465);
and U14521 (N_14521,N_13688,N_13231);
nor U14522 (N_14522,N_13098,N_13031);
or U14523 (N_14523,N_13758,N_13013);
and U14524 (N_14524,N_13132,N_13083);
nor U14525 (N_14525,N_13382,N_13739);
xor U14526 (N_14526,N_13210,N_13207);
or U14527 (N_14527,N_13085,N_13433);
or U14528 (N_14528,N_13755,N_13100);
nor U14529 (N_14529,N_13951,N_13566);
or U14530 (N_14530,N_13297,N_13102);
nor U14531 (N_14531,N_13738,N_13563);
nand U14532 (N_14532,N_13845,N_13383);
nor U14533 (N_14533,N_13350,N_13964);
nor U14534 (N_14534,N_13022,N_13491);
xor U14535 (N_14535,N_13677,N_13060);
nand U14536 (N_14536,N_13619,N_13309);
xor U14537 (N_14537,N_13683,N_13300);
nor U14538 (N_14538,N_13844,N_13132);
or U14539 (N_14539,N_13537,N_13904);
xnor U14540 (N_14540,N_13820,N_13841);
and U14541 (N_14541,N_13108,N_13798);
nand U14542 (N_14542,N_13078,N_13642);
or U14543 (N_14543,N_13312,N_13252);
nor U14544 (N_14544,N_13090,N_13258);
nor U14545 (N_14545,N_13463,N_13798);
xor U14546 (N_14546,N_13190,N_13944);
or U14547 (N_14547,N_13928,N_13377);
nor U14548 (N_14548,N_13297,N_13812);
nor U14549 (N_14549,N_13678,N_13039);
xnor U14550 (N_14550,N_13605,N_13645);
nor U14551 (N_14551,N_13286,N_13499);
or U14552 (N_14552,N_13799,N_13549);
or U14553 (N_14553,N_13448,N_13135);
nand U14554 (N_14554,N_13922,N_13495);
nand U14555 (N_14555,N_13630,N_13223);
xor U14556 (N_14556,N_13297,N_13020);
and U14557 (N_14557,N_13788,N_13669);
xor U14558 (N_14558,N_13916,N_13708);
nor U14559 (N_14559,N_13078,N_13784);
or U14560 (N_14560,N_13916,N_13238);
nor U14561 (N_14561,N_13295,N_13975);
xnor U14562 (N_14562,N_13460,N_13049);
and U14563 (N_14563,N_13105,N_13643);
and U14564 (N_14564,N_13004,N_13983);
or U14565 (N_14565,N_13907,N_13009);
xor U14566 (N_14566,N_13003,N_13030);
nor U14567 (N_14567,N_13165,N_13026);
and U14568 (N_14568,N_13293,N_13167);
nand U14569 (N_14569,N_13261,N_13832);
xnor U14570 (N_14570,N_13842,N_13988);
xor U14571 (N_14571,N_13281,N_13089);
xor U14572 (N_14572,N_13475,N_13298);
or U14573 (N_14573,N_13097,N_13406);
nor U14574 (N_14574,N_13234,N_13643);
or U14575 (N_14575,N_13446,N_13529);
and U14576 (N_14576,N_13530,N_13818);
nand U14577 (N_14577,N_13008,N_13266);
and U14578 (N_14578,N_13402,N_13819);
and U14579 (N_14579,N_13690,N_13482);
or U14580 (N_14580,N_13298,N_13628);
nand U14581 (N_14581,N_13584,N_13235);
or U14582 (N_14582,N_13866,N_13780);
or U14583 (N_14583,N_13299,N_13195);
nor U14584 (N_14584,N_13346,N_13833);
and U14585 (N_14585,N_13690,N_13558);
or U14586 (N_14586,N_13187,N_13926);
and U14587 (N_14587,N_13308,N_13340);
or U14588 (N_14588,N_13988,N_13607);
nand U14589 (N_14589,N_13031,N_13741);
nand U14590 (N_14590,N_13877,N_13393);
nand U14591 (N_14591,N_13499,N_13574);
nor U14592 (N_14592,N_13750,N_13754);
or U14593 (N_14593,N_13550,N_13229);
and U14594 (N_14594,N_13848,N_13553);
and U14595 (N_14595,N_13187,N_13810);
nor U14596 (N_14596,N_13901,N_13895);
nand U14597 (N_14597,N_13528,N_13493);
and U14598 (N_14598,N_13943,N_13480);
xor U14599 (N_14599,N_13028,N_13185);
xor U14600 (N_14600,N_13584,N_13402);
nand U14601 (N_14601,N_13076,N_13483);
or U14602 (N_14602,N_13999,N_13703);
or U14603 (N_14603,N_13837,N_13656);
and U14604 (N_14604,N_13364,N_13880);
or U14605 (N_14605,N_13807,N_13399);
and U14606 (N_14606,N_13595,N_13644);
or U14607 (N_14607,N_13350,N_13574);
nor U14608 (N_14608,N_13255,N_13109);
nor U14609 (N_14609,N_13161,N_13723);
nor U14610 (N_14610,N_13094,N_13333);
or U14611 (N_14611,N_13543,N_13577);
nor U14612 (N_14612,N_13119,N_13778);
and U14613 (N_14613,N_13080,N_13965);
nor U14614 (N_14614,N_13478,N_13884);
nor U14615 (N_14615,N_13807,N_13321);
and U14616 (N_14616,N_13221,N_13309);
or U14617 (N_14617,N_13720,N_13803);
or U14618 (N_14618,N_13467,N_13830);
or U14619 (N_14619,N_13843,N_13018);
xnor U14620 (N_14620,N_13370,N_13231);
nor U14621 (N_14621,N_13884,N_13033);
and U14622 (N_14622,N_13527,N_13579);
nand U14623 (N_14623,N_13017,N_13135);
xor U14624 (N_14624,N_13260,N_13056);
xor U14625 (N_14625,N_13771,N_13808);
and U14626 (N_14626,N_13741,N_13180);
nor U14627 (N_14627,N_13431,N_13399);
nor U14628 (N_14628,N_13159,N_13897);
and U14629 (N_14629,N_13086,N_13927);
and U14630 (N_14630,N_13171,N_13232);
nor U14631 (N_14631,N_13390,N_13358);
and U14632 (N_14632,N_13947,N_13641);
or U14633 (N_14633,N_13707,N_13496);
nand U14634 (N_14634,N_13035,N_13075);
nor U14635 (N_14635,N_13386,N_13882);
xor U14636 (N_14636,N_13340,N_13874);
nand U14637 (N_14637,N_13819,N_13266);
nor U14638 (N_14638,N_13327,N_13985);
nor U14639 (N_14639,N_13045,N_13243);
or U14640 (N_14640,N_13910,N_13328);
nand U14641 (N_14641,N_13063,N_13534);
nand U14642 (N_14642,N_13923,N_13585);
or U14643 (N_14643,N_13092,N_13014);
nor U14644 (N_14644,N_13829,N_13001);
nor U14645 (N_14645,N_13164,N_13625);
or U14646 (N_14646,N_13775,N_13166);
nand U14647 (N_14647,N_13510,N_13426);
nor U14648 (N_14648,N_13932,N_13217);
and U14649 (N_14649,N_13508,N_13423);
nand U14650 (N_14650,N_13425,N_13537);
nor U14651 (N_14651,N_13570,N_13203);
nor U14652 (N_14652,N_13567,N_13020);
xor U14653 (N_14653,N_13673,N_13909);
nand U14654 (N_14654,N_13427,N_13248);
nand U14655 (N_14655,N_13555,N_13638);
nor U14656 (N_14656,N_13585,N_13501);
or U14657 (N_14657,N_13001,N_13159);
or U14658 (N_14658,N_13418,N_13938);
and U14659 (N_14659,N_13028,N_13503);
nand U14660 (N_14660,N_13454,N_13806);
and U14661 (N_14661,N_13074,N_13155);
xor U14662 (N_14662,N_13961,N_13998);
or U14663 (N_14663,N_13592,N_13617);
nand U14664 (N_14664,N_13230,N_13060);
nor U14665 (N_14665,N_13742,N_13904);
or U14666 (N_14666,N_13626,N_13253);
and U14667 (N_14667,N_13375,N_13150);
nand U14668 (N_14668,N_13686,N_13951);
or U14669 (N_14669,N_13037,N_13521);
nor U14670 (N_14670,N_13949,N_13516);
nor U14671 (N_14671,N_13943,N_13276);
nor U14672 (N_14672,N_13278,N_13989);
or U14673 (N_14673,N_13915,N_13230);
or U14674 (N_14674,N_13120,N_13898);
nor U14675 (N_14675,N_13615,N_13763);
nand U14676 (N_14676,N_13427,N_13704);
and U14677 (N_14677,N_13335,N_13247);
or U14678 (N_14678,N_13560,N_13941);
nand U14679 (N_14679,N_13335,N_13134);
or U14680 (N_14680,N_13861,N_13978);
xnor U14681 (N_14681,N_13285,N_13360);
and U14682 (N_14682,N_13698,N_13409);
nand U14683 (N_14683,N_13979,N_13227);
or U14684 (N_14684,N_13064,N_13102);
nand U14685 (N_14685,N_13650,N_13784);
xor U14686 (N_14686,N_13051,N_13904);
or U14687 (N_14687,N_13783,N_13999);
nor U14688 (N_14688,N_13581,N_13406);
or U14689 (N_14689,N_13724,N_13003);
nor U14690 (N_14690,N_13941,N_13315);
xnor U14691 (N_14691,N_13457,N_13700);
nand U14692 (N_14692,N_13532,N_13857);
nand U14693 (N_14693,N_13414,N_13850);
and U14694 (N_14694,N_13742,N_13911);
nor U14695 (N_14695,N_13506,N_13915);
or U14696 (N_14696,N_13109,N_13058);
and U14697 (N_14697,N_13789,N_13061);
or U14698 (N_14698,N_13528,N_13549);
nor U14699 (N_14699,N_13992,N_13082);
and U14700 (N_14700,N_13835,N_13082);
and U14701 (N_14701,N_13678,N_13604);
and U14702 (N_14702,N_13564,N_13710);
nand U14703 (N_14703,N_13021,N_13372);
or U14704 (N_14704,N_13941,N_13475);
nand U14705 (N_14705,N_13566,N_13531);
nor U14706 (N_14706,N_13014,N_13643);
nor U14707 (N_14707,N_13554,N_13297);
and U14708 (N_14708,N_13855,N_13069);
xnor U14709 (N_14709,N_13241,N_13340);
or U14710 (N_14710,N_13314,N_13921);
nand U14711 (N_14711,N_13933,N_13454);
nor U14712 (N_14712,N_13830,N_13887);
and U14713 (N_14713,N_13748,N_13113);
nor U14714 (N_14714,N_13747,N_13488);
nor U14715 (N_14715,N_13034,N_13863);
and U14716 (N_14716,N_13460,N_13656);
nor U14717 (N_14717,N_13579,N_13802);
xnor U14718 (N_14718,N_13106,N_13996);
or U14719 (N_14719,N_13694,N_13990);
nor U14720 (N_14720,N_13507,N_13693);
xnor U14721 (N_14721,N_13319,N_13905);
or U14722 (N_14722,N_13798,N_13332);
or U14723 (N_14723,N_13718,N_13986);
or U14724 (N_14724,N_13458,N_13273);
nor U14725 (N_14725,N_13886,N_13649);
and U14726 (N_14726,N_13247,N_13704);
nor U14727 (N_14727,N_13294,N_13422);
and U14728 (N_14728,N_13878,N_13830);
nor U14729 (N_14729,N_13364,N_13594);
or U14730 (N_14730,N_13365,N_13882);
and U14731 (N_14731,N_13268,N_13440);
nand U14732 (N_14732,N_13994,N_13740);
or U14733 (N_14733,N_13700,N_13714);
nor U14734 (N_14734,N_13297,N_13031);
and U14735 (N_14735,N_13340,N_13251);
and U14736 (N_14736,N_13588,N_13414);
or U14737 (N_14737,N_13071,N_13688);
or U14738 (N_14738,N_13308,N_13404);
and U14739 (N_14739,N_13861,N_13860);
or U14740 (N_14740,N_13692,N_13728);
and U14741 (N_14741,N_13568,N_13880);
or U14742 (N_14742,N_13235,N_13109);
or U14743 (N_14743,N_13998,N_13769);
xor U14744 (N_14744,N_13235,N_13287);
nand U14745 (N_14745,N_13124,N_13333);
and U14746 (N_14746,N_13485,N_13164);
or U14747 (N_14747,N_13859,N_13933);
nor U14748 (N_14748,N_13229,N_13541);
or U14749 (N_14749,N_13183,N_13808);
nor U14750 (N_14750,N_13307,N_13863);
xor U14751 (N_14751,N_13416,N_13587);
nand U14752 (N_14752,N_13245,N_13763);
or U14753 (N_14753,N_13852,N_13625);
nor U14754 (N_14754,N_13796,N_13146);
or U14755 (N_14755,N_13874,N_13640);
xnor U14756 (N_14756,N_13899,N_13255);
nand U14757 (N_14757,N_13328,N_13731);
and U14758 (N_14758,N_13812,N_13942);
nor U14759 (N_14759,N_13102,N_13858);
xor U14760 (N_14760,N_13164,N_13612);
or U14761 (N_14761,N_13430,N_13052);
and U14762 (N_14762,N_13584,N_13356);
and U14763 (N_14763,N_13290,N_13596);
nand U14764 (N_14764,N_13733,N_13656);
nor U14765 (N_14765,N_13362,N_13266);
xor U14766 (N_14766,N_13801,N_13437);
and U14767 (N_14767,N_13976,N_13427);
or U14768 (N_14768,N_13334,N_13142);
and U14769 (N_14769,N_13078,N_13552);
and U14770 (N_14770,N_13692,N_13060);
nand U14771 (N_14771,N_13726,N_13298);
nor U14772 (N_14772,N_13528,N_13449);
and U14773 (N_14773,N_13251,N_13586);
xor U14774 (N_14774,N_13265,N_13498);
or U14775 (N_14775,N_13053,N_13930);
nor U14776 (N_14776,N_13306,N_13996);
nor U14777 (N_14777,N_13266,N_13621);
or U14778 (N_14778,N_13895,N_13161);
or U14779 (N_14779,N_13030,N_13805);
and U14780 (N_14780,N_13134,N_13912);
or U14781 (N_14781,N_13589,N_13922);
nor U14782 (N_14782,N_13837,N_13375);
and U14783 (N_14783,N_13900,N_13036);
and U14784 (N_14784,N_13963,N_13324);
and U14785 (N_14785,N_13525,N_13959);
and U14786 (N_14786,N_13704,N_13223);
xor U14787 (N_14787,N_13267,N_13619);
and U14788 (N_14788,N_13183,N_13241);
nor U14789 (N_14789,N_13653,N_13083);
or U14790 (N_14790,N_13412,N_13487);
or U14791 (N_14791,N_13399,N_13386);
nand U14792 (N_14792,N_13216,N_13672);
xor U14793 (N_14793,N_13041,N_13803);
or U14794 (N_14794,N_13752,N_13218);
nand U14795 (N_14795,N_13431,N_13081);
nor U14796 (N_14796,N_13417,N_13515);
nor U14797 (N_14797,N_13329,N_13558);
xnor U14798 (N_14798,N_13531,N_13298);
nor U14799 (N_14799,N_13089,N_13963);
and U14800 (N_14800,N_13947,N_13737);
and U14801 (N_14801,N_13719,N_13090);
and U14802 (N_14802,N_13562,N_13093);
nand U14803 (N_14803,N_13489,N_13660);
and U14804 (N_14804,N_13807,N_13732);
nor U14805 (N_14805,N_13056,N_13377);
and U14806 (N_14806,N_13814,N_13860);
nand U14807 (N_14807,N_13539,N_13571);
or U14808 (N_14808,N_13449,N_13358);
nor U14809 (N_14809,N_13642,N_13052);
nor U14810 (N_14810,N_13313,N_13462);
nand U14811 (N_14811,N_13966,N_13705);
nor U14812 (N_14812,N_13235,N_13711);
xor U14813 (N_14813,N_13667,N_13530);
nor U14814 (N_14814,N_13962,N_13566);
or U14815 (N_14815,N_13984,N_13520);
nand U14816 (N_14816,N_13278,N_13347);
nand U14817 (N_14817,N_13457,N_13743);
nor U14818 (N_14818,N_13469,N_13784);
or U14819 (N_14819,N_13062,N_13967);
or U14820 (N_14820,N_13575,N_13895);
nor U14821 (N_14821,N_13657,N_13631);
nor U14822 (N_14822,N_13323,N_13941);
xor U14823 (N_14823,N_13438,N_13849);
or U14824 (N_14824,N_13632,N_13485);
nor U14825 (N_14825,N_13936,N_13300);
nor U14826 (N_14826,N_13544,N_13964);
nand U14827 (N_14827,N_13224,N_13770);
or U14828 (N_14828,N_13228,N_13482);
and U14829 (N_14829,N_13766,N_13601);
xnor U14830 (N_14830,N_13040,N_13058);
nor U14831 (N_14831,N_13356,N_13623);
xnor U14832 (N_14832,N_13455,N_13624);
and U14833 (N_14833,N_13230,N_13111);
or U14834 (N_14834,N_13508,N_13359);
or U14835 (N_14835,N_13677,N_13749);
xnor U14836 (N_14836,N_13029,N_13467);
xor U14837 (N_14837,N_13661,N_13740);
nand U14838 (N_14838,N_13978,N_13886);
or U14839 (N_14839,N_13692,N_13561);
nor U14840 (N_14840,N_13978,N_13998);
or U14841 (N_14841,N_13888,N_13831);
nor U14842 (N_14842,N_13352,N_13552);
and U14843 (N_14843,N_13291,N_13356);
and U14844 (N_14844,N_13475,N_13520);
or U14845 (N_14845,N_13322,N_13220);
nor U14846 (N_14846,N_13072,N_13480);
nor U14847 (N_14847,N_13845,N_13375);
or U14848 (N_14848,N_13672,N_13157);
or U14849 (N_14849,N_13355,N_13018);
and U14850 (N_14850,N_13676,N_13202);
nand U14851 (N_14851,N_13431,N_13282);
nor U14852 (N_14852,N_13054,N_13674);
nand U14853 (N_14853,N_13719,N_13163);
or U14854 (N_14854,N_13768,N_13472);
nor U14855 (N_14855,N_13290,N_13522);
and U14856 (N_14856,N_13258,N_13375);
or U14857 (N_14857,N_13795,N_13958);
and U14858 (N_14858,N_13036,N_13457);
nand U14859 (N_14859,N_13959,N_13400);
xnor U14860 (N_14860,N_13578,N_13277);
nor U14861 (N_14861,N_13518,N_13548);
nor U14862 (N_14862,N_13653,N_13527);
and U14863 (N_14863,N_13074,N_13849);
xor U14864 (N_14864,N_13548,N_13760);
nand U14865 (N_14865,N_13357,N_13392);
or U14866 (N_14866,N_13292,N_13162);
and U14867 (N_14867,N_13256,N_13411);
and U14868 (N_14868,N_13131,N_13254);
nor U14869 (N_14869,N_13064,N_13585);
nand U14870 (N_14870,N_13271,N_13438);
nor U14871 (N_14871,N_13556,N_13694);
xnor U14872 (N_14872,N_13137,N_13912);
or U14873 (N_14873,N_13785,N_13240);
or U14874 (N_14874,N_13948,N_13464);
xor U14875 (N_14875,N_13706,N_13189);
nor U14876 (N_14876,N_13484,N_13124);
and U14877 (N_14877,N_13333,N_13222);
or U14878 (N_14878,N_13019,N_13127);
nand U14879 (N_14879,N_13143,N_13941);
nor U14880 (N_14880,N_13982,N_13338);
nor U14881 (N_14881,N_13860,N_13314);
nand U14882 (N_14882,N_13628,N_13971);
and U14883 (N_14883,N_13241,N_13778);
and U14884 (N_14884,N_13120,N_13689);
xor U14885 (N_14885,N_13270,N_13247);
and U14886 (N_14886,N_13404,N_13723);
or U14887 (N_14887,N_13706,N_13125);
nand U14888 (N_14888,N_13732,N_13497);
or U14889 (N_14889,N_13180,N_13535);
xor U14890 (N_14890,N_13011,N_13450);
xor U14891 (N_14891,N_13015,N_13866);
and U14892 (N_14892,N_13527,N_13194);
xnor U14893 (N_14893,N_13361,N_13930);
nand U14894 (N_14894,N_13079,N_13843);
or U14895 (N_14895,N_13710,N_13080);
and U14896 (N_14896,N_13253,N_13825);
nor U14897 (N_14897,N_13837,N_13099);
xor U14898 (N_14898,N_13855,N_13014);
xnor U14899 (N_14899,N_13493,N_13123);
nor U14900 (N_14900,N_13619,N_13221);
or U14901 (N_14901,N_13661,N_13316);
nor U14902 (N_14902,N_13469,N_13565);
and U14903 (N_14903,N_13240,N_13299);
and U14904 (N_14904,N_13495,N_13045);
or U14905 (N_14905,N_13319,N_13975);
and U14906 (N_14906,N_13897,N_13175);
or U14907 (N_14907,N_13255,N_13713);
nand U14908 (N_14908,N_13569,N_13702);
nand U14909 (N_14909,N_13494,N_13571);
nor U14910 (N_14910,N_13603,N_13925);
nor U14911 (N_14911,N_13805,N_13570);
and U14912 (N_14912,N_13742,N_13045);
and U14913 (N_14913,N_13149,N_13942);
nand U14914 (N_14914,N_13526,N_13316);
and U14915 (N_14915,N_13718,N_13908);
xnor U14916 (N_14916,N_13456,N_13695);
or U14917 (N_14917,N_13408,N_13357);
nor U14918 (N_14918,N_13311,N_13559);
or U14919 (N_14919,N_13812,N_13138);
and U14920 (N_14920,N_13982,N_13110);
or U14921 (N_14921,N_13468,N_13332);
and U14922 (N_14922,N_13448,N_13942);
nor U14923 (N_14923,N_13754,N_13380);
or U14924 (N_14924,N_13543,N_13270);
nand U14925 (N_14925,N_13180,N_13665);
or U14926 (N_14926,N_13355,N_13861);
or U14927 (N_14927,N_13647,N_13009);
nor U14928 (N_14928,N_13482,N_13701);
nor U14929 (N_14929,N_13235,N_13278);
or U14930 (N_14930,N_13906,N_13358);
or U14931 (N_14931,N_13931,N_13643);
nand U14932 (N_14932,N_13640,N_13404);
and U14933 (N_14933,N_13878,N_13487);
nand U14934 (N_14934,N_13144,N_13549);
nand U14935 (N_14935,N_13624,N_13843);
nor U14936 (N_14936,N_13582,N_13025);
nor U14937 (N_14937,N_13504,N_13565);
nand U14938 (N_14938,N_13050,N_13138);
and U14939 (N_14939,N_13059,N_13523);
and U14940 (N_14940,N_13662,N_13086);
nor U14941 (N_14941,N_13580,N_13545);
and U14942 (N_14942,N_13736,N_13616);
and U14943 (N_14943,N_13936,N_13896);
nand U14944 (N_14944,N_13248,N_13657);
xor U14945 (N_14945,N_13757,N_13807);
and U14946 (N_14946,N_13892,N_13093);
and U14947 (N_14947,N_13615,N_13256);
xnor U14948 (N_14948,N_13061,N_13355);
or U14949 (N_14949,N_13346,N_13635);
nor U14950 (N_14950,N_13641,N_13108);
nor U14951 (N_14951,N_13237,N_13065);
nor U14952 (N_14952,N_13857,N_13713);
nand U14953 (N_14953,N_13764,N_13790);
nor U14954 (N_14954,N_13423,N_13326);
or U14955 (N_14955,N_13481,N_13346);
nor U14956 (N_14956,N_13572,N_13301);
nand U14957 (N_14957,N_13945,N_13183);
nor U14958 (N_14958,N_13499,N_13946);
or U14959 (N_14959,N_13659,N_13612);
or U14960 (N_14960,N_13420,N_13213);
nand U14961 (N_14961,N_13433,N_13706);
xor U14962 (N_14962,N_13173,N_13796);
xor U14963 (N_14963,N_13058,N_13326);
and U14964 (N_14964,N_13004,N_13027);
or U14965 (N_14965,N_13641,N_13848);
nand U14966 (N_14966,N_13426,N_13140);
and U14967 (N_14967,N_13919,N_13867);
and U14968 (N_14968,N_13552,N_13047);
and U14969 (N_14969,N_13258,N_13656);
and U14970 (N_14970,N_13885,N_13353);
nor U14971 (N_14971,N_13501,N_13703);
nor U14972 (N_14972,N_13106,N_13934);
nand U14973 (N_14973,N_13748,N_13776);
nor U14974 (N_14974,N_13848,N_13861);
nand U14975 (N_14975,N_13461,N_13628);
nor U14976 (N_14976,N_13983,N_13478);
or U14977 (N_14977,N_13342,N_13785);
or U14978 (N_14978,N_13554,N_13095);
and U14979 (N_14979,N_13571,N_13350);
and U14980 (N_14980,N_13763,N_13094);
nand U14981 (N_14981,N_13395,N_13788);
xnor U14982 (N_14982,N_13972,N_13019);
nand U14983 (N_14983,N_13289,N_13578);
and U14984 (N_14984,N_13748,N_13720);
nand U14985 (N_14985,N_13362,N_13201);
and U14986 (N_14986,N_13800,N_13140);
or U14987 (N_14987,N_13731,N_13804);
nand U14988 (N_14988,N_13750,N_13165);
nand U14989 (N_14989,N_13090,N_13493);
and U14990 (N_14990,N_13839,N_13050);
and U14991 (N_14991,N_13131,N_13574);
nand U14992 (N_14992,N_13447,N_13379);
or U14993 (N_14993,N_13092,N_13157);
nor U14994 (N_14994,N_13675,N_13238);
or U14995 (N_14995,N_13734,N_13458);
or U14996 (N_14996,N_13361,N_13670);
xnor U14997 (N_14997,N_13047,N_13890);
or U14998 (N_14998,N_13812,N_13914);
and U14999 (N_14999,N_13765,N_13797);
nor UO_0 (O_0,N_14587,N_14810);
or UO_1 (O_1,N_14839,N_14772);
nor UO_2 (O_2,N_14061,N_14570);
nor UO_3 (O_3,N_14196,N_14649);
or UO_4 (O_4,N_14966,N_14999);
or UO_5 (O_5,N_14412,N_14174);
nor UO_6 (O_6,N_14064,N_14493);
or UO_7 (O_7,N_14115,N_14343);
or UO_8 (O_8,N_14494,N_14199);
and UO_9 (O_9,N_14325,N_14243);
and UO_10 (O_10,N_14331,N_14079);
nand UO_11 (O_11,N_14785,N_14101);
nand UO_12 (O_12,N_14751,N_14367);
or UO_13 (O_13,N_14216,N_14789);
or UO_14 (O_14,N_14022,N_14204);
nor UO_15 (O_15,N_14518,N_14226);
nor UO_16 (O_16,N_14597,N_14076);
nor UO_17 (O_17,N_14956,N_14608);
or UO_18 (O_18,N_14060,N_14313);
nand UO_19 (O_19,N_14055,N_14417);
nand UO_20 (O_20,N_14705,N_14276);
nor UO_21 (O_21,N_14534,N_14780);
or UO_22 (O_22,N_14007,N_14891);
nor UO_23 (O_23,N_14162,N_14663);
and UO_24 (O_24,N_14519,N_14644);
nand UO_25 (O_25,N_14855,N_14748);
nand UO_26 (O_26,N_14821,N_14374);
nand UO_27 (O_27,N_14660,N_14320);
or UO_28 (O_28,N_14967,N_14184);
nand UO_29 (O_29,N_14119,N_14275);
or UO_30 (O_30,N_14652,N_14048);
and UO_31 (O_31,N_14526,N_14292);
and UO_32 (O_32,N_14269,N_14582);
nor UO_33 (O_33,N_14865,N_14172);
nor UO_34 (O_34,N_14816,N_14293);
and UO_35 (O_35,N_14573,N_14026);
nor UO_36 (O_36,N_14131,N_14757);
and UO_37 (O_37,N_14797,N_14399);
xnor UO_38 (O_38,N_14223,N_14837);
xnor UO_39 (O_39,N_14423,N_14273);
and UO_40 (O_40,N_14856,N_14181);
nor UO_41 (O_41,N_14539,N_14592);
nand UO_42 (O_42,N_14874,N_14274);
and UO_43 (O_43,N_14200,N_14237);
nand UO_44 (O_44,N_14585,N_14943);
nand UO_45 (O_45,N_14169,N_14998);
xnor UO_46 (O_46,N_14686,N_14375);
and UO_47 (O_47,N_14572,N_14233);
nand UO_48 (O_48,N_14287,N_14762);
nand UO_49 (O_49,N_14366,N_14257);
or UO_50 (O_50,N_14121,N_14405);
or UO_51 (O_51,N_14791,N_14471);
or UO_52 (O_52,N_14890,N_14372);
and UO_53 (O_53,N_14160,N_14738);
nor UO_54 (O_54,N_14279,N_14744);
or UO_55 (O_55,N_14349,N_14787);
or UO_56 (O_56,N_14595,N_14345);
or UO_57 (O_57,N_14522,N_14511);
and UO_58 (O_58,N_14490,N_14838);
nor UO_59 (O_59,N_14932,N_14866);
nand UO_60 (O_60,N_14496,N_14877);
nor UO_61 (O_61,N_14189,N_14662);
nand UO_62 (O_62,N_14393,N_14538);
nor UO_63 (O_63,N_14616,N_14224);
nand UO_64 (O_64,N_14763,N_14182);
or UO_65 (O_65,N_14097,N_14438);
xor UO_66 (O_66,N_14642,N_14802);
nand UO_67 (O_67,N_14152,N_14042);
nor UO_68 (O_68,N_14986,N_14485);
nand UO_69 (O_69,N_14626,N_14256);
or UO_70 (O_70,N_14926,N_14533);
and UO_71 (O_71,N_14911,N_14825);
or UO_72 (O_72,N_14148,N_14197);
nand UO_73 (O_73,N_14103,N_14795);
and UO_74 (O_74,N_14057,N_14672);
and UO_75 (O_75,N_14283,N_14841);
xor UO_76 (O_76,N_14435,N_14898);
or UO_77 (O_77,N_14150,N_14428);
nor UO_78 (O_78,N_14736,N_14901);
and UO_79 (O_79,N_14019,N_14715);
nor UO_80 (O_80,N_14873,N_14422);
and UO_81 (O_81,N_14457,N_14832);
or UO_82 (O_82,N_14770,N_14537);
nor UO_83 (O_83,N_14447,N_14563);
nand UO_84 (O_84,N_14364,N_14786);
nor UO_85 (O_85,N_14136,N_14588);
or UO_86 (O_86,N_14981,N_14408);
nand UO_87 (O_87,N_14957,N_14657);
nor UO_88 (O_88,N_14694,N_14466);
or UO_89 (O_89,N_14098,N_14056);
nand UO_90 (O_90,N_14779,N_14149);
xor UO_91 (O_91,N_14730,N_14888);
xor UO_92 (O_92,N_14215,N_14488);
nor UO_93 (O_93,N_14454,N_14727);
nand UO_94 (O_94,N_14213,N_14960);
nor UO_95 (O_95,N_14432,N_14555);
and UO_96 (O_96,N_14604,N_14589);
or UO_97 (O_97,N_14872,N_14909);
nor UO_98 (O_98,N_14979,N_14851);
and UO_99 (O_99,N_14147,N_14983);
and UO_100 (O_100,N_14191,N_14869);
nand UO_101 (O_101,N_14504,N_14370);
nor UO_102 (O_102,N_14940,N_14567);
and UO_103 (O_103,N_14426,N_14247);
nand UO_104 (O_104,N_14497,N_14424);
and UO_105 (O_105,N_14985,N_14557);
or UO_106 (O_106,N_14348,N_14452);
nand UO_107 (O_107,N_14655,N_14951);
nor UO_108 (O_108,N_14982,N_14716);
nor UO_109 (O_109,N_14719,N_14826);
and UO_110 (O_110,N_14993,N_14962);
nand UO_111 (O_111,N_14380,N_14709);
or UO_112 (O_112,N_14352,N_14677);
or UO_113 (O_113,N_14938,N_14599);
nor UO_114 (O_114,N_14868,N_14092);
nor UO_115 (O_115,N_14397,N_14445);
nand UO_116 (O_116,N_14384,N_14137);
nand UO_117 (O_117,N_14858,N_14790);
or UO_118 (O_118,N_14344,N_14516);
and UO_119 (O_119,N_14603,N_14508);
or UO_120 (O_120,N_14116,N_14914);
or UO_121 (O_121,N_14971,N_14921);
nor UO_122 (O_122,N_14812,N_14126);
nor UO_123 (O_123,N_14823,N_14469);
and UO_124 (O_124,N_14842,N_14752);
nand UO_125 (O_125,N_14562,N_14910);
nor UO_126 (O_126,N_14300,N_14388);
and UO_127 (O_127,N_14402,N_14613);
nand UO_128 (O_128,N_14928,N_14646);
nand UO_129 (O_129,N_14864,N_14569);
xnor UO_130 (O_130,N_14647,N_14578);
nand UO_131 (O_131,N_14581,N_14666);
or UO_132 (O_132,N_14483,N_14086);
nand UO_133 (O_133,N_14122,N_14777);
nor UO_134 (O_134,N_14693,N_14704);
nand UO_135 (O_135,N_14210,N_14029);
and UO_136 (O_136,N_14846,N_14706);
and UO_137 (O_137,N_14106,N_14164);
and UO_138 (O_138,N_14617,N_14318);
or UO_139 (O_139,N_14536,N_14753);
or UO_140 (O_140,N_14593,N_14404);
and UO_141 (O_141,N_14749,N_14586);
or UO_142 (O_142,N_14299,N_14782);
nor UO_143 (O_143,N_14840,N_14886);
xnor UO_144 (O_144,N_14958,N_14282);
or UO_145 (O_145,N_14072,N_14000);
nand UO_146 (O_146,N_14711,N_14168);
nor UO_147 (O_147,N_14110,N_14355);
or UO_148 (O_148,N_14140,N_14338);
and UO_149 (O_149,N_14176,N_14077);
and UO_150 (O_150,N_14734,N_14661);
and UO_151 (O_151,N_14643,N_14442);
nor UO_152 (O_152,N_14698,N_14193);
and UO_153 (O_153,N_14255,N_14378);
or UO_154 (O_154,N_14512,N_14259);
xnor UO_155 (O_155,N_14684,N_14188);
nor UO_156 (O_156,N_14712,N_14532);
nand UO_157 (O_157,N_14852,N_14212);
nor UO_158 (O_158,N_14130,N_14612);
nand UO_159 (O_159,N_14605,N_14429);
and UO_160 (O_160,N_14623,N_14031);
nand UO_161 (O_161,N_14545,N_14175);
nor UO_162 (O_162,N_14362,N_14792);
xnor UO_163 (O_163,N_14847,N_14203);
nand UO_164 (O_164,N_14850,N_14479);
or UO_165 (O_165,N_14687,N_14472);
nand UO_166 (O_166,N_14069,N_14540);
and UO_167 (O_167,N_14067,N_14844);
nand UO_168 (O_168,N_14195,N_14547);
nand UO_169 (O_169,N_14087,N_14333);
or UO_170 (O_170,N_14930,N_14509);
and UO_171 (O_171,N_14924,N_14353);
nand UO_172 (O_172,N_14024,N_14946);
and UO_173 (O_173,N_14571,N_14037);
nor UO_174 (O_174,N_14499,N_14436);
nand UO_175 (O_175,N_14099,N_14440);
nand UO_176 (O_176,N_14641,N_14228);
nor UO_177 (O_177,N_14120,N_14030);
nor UO_178 (O_178,N_14095,N_14574);
nor UO_179 (O_179,N_14679,N_14936);
nor UO_180 (O_180,N_14317,N_14633);
and UO_181 (O_181,N_14968,N_14773);
and UO_182 (O_182,N_14887,N_14740);
xnor UO_183 (O_183,N_14339,N_14066);
nor UO_184 (O_184,N_14922,N_14398);
and UO_185 (O_185,N_14093,N_14674);
nand UO_186 (O_186,N_14668,N_14034);
nand UO_187 (O_187,N_14368,N_14141);
nor UO_188 (O_188,N_14123,N_14225);
xor UO_189 (O_189,N_14453,N_14735);
and UO_190 (O_190,N_14319,N_14265);
nor UO_191 (O_191,N_14996,N_14281);
and UO_192 (O_192,N_14251,N_14023);
nor UO_193 (O_193,N_14854,N_14052);
nor UO_194 (O_194,N_14403,N_14607);
or UO_195 (O_195,N_14879,N_14796);
or UO_196 (O_196,N_14845,N_14503);
nor UO_197 (O_197,N_14009,N_14420);
xnor UO_198 (O_198,N_14272,N_14733);
nor UO_199 (O_199,N_14492,N_14878);
and UO_200 (O_200,N_14920,N_14827);
nand UO_201 (O_201,N_14918,N_14018);
and UO_202 (O_202,N_14202,N_14798);
or UO_203 (O_203,N_14699,N_14171);
xor UO_204 (O_204,N_14448,N_14462);
or UO_205 (O_205,N_14290,N_14482);
nor UO_206 (O_206,N_14044,N_14238);
and UO_207 (O_207,N_14811,N_14289);
or UO_208 (O_208,N_14903,N_14336);
and UO_209 (O_209,N_14531,N_14696);
and UO_210 (O_210,N_14543,N_14041);
and UO_211 (O_211,N_14082,N_14630);
and UO_212 (O_212,N_14559,N_14080);
and UO_213 (O_213,N_14594,N_14470);
nor UO_214 (O_214,N_14477,N_14973);
and UO_215 (O_215,N_14818,N_14863);
and UO_216 (O_216,N_14411,N_14908);
and UO_217 (O_217,N_14640,N_14419);
nor UO_218 (O_218,N_14558,N_14520);
nor UO_219 (O_219,N_14484,N_14389);
and UO_220 (O_220,N_14305,N_14745);
xor UO_221 (O_221,N_14142,N_14400);
nand UO_222 (O_222,N_14964,N_14965);
nand UO_223 (O_223,N_14510,N_14710);
or UO_224 (O_224,N_14486,N_14070);
nor UO_225 (O_225,N_14312,N_14241);
and UO_226 (O_226,N_14675,N_14871);
nor UO_227 (O_227,N_14135,N_14867);
nand UO_228 (O_228,N_14244,N_14737);
xnor UO_229 (O_229,N_14764,N_14671);
nor UO_230 (O_230,N_14058,N_14731);
xor UO_231 (O_231,N_14288,N_14134);
nor UO_232 (O_232,N_14309,N_14154);
nand UO_233 (O_233,N_14383,N_14377);
nor UO_234 (O_234,N_14434,N_14253);
nand UO_235 (O_235,N_14584,N_14109);
nand UO_236 (O_236,N_14491,N_14459);
nor UO_237 (O_237,N_14021,N_14340);
and UO_238 (O_238,N_14885,N_14893);
or UO_239 (O_239,N_14799,N_14915);
nand UO_240 (O_240,N_14307,N_14218);
and UO_241 (O_241,N_14899,N_14304);
xnor UO_242 (O_242,N_14028,N_14853);
xnor UO_243 (O_243,N_14664,N_14989);
and UO_244 (O_244,N_14033,N_14179);
xor UO_245 (O_245,N_14451,N_14342);
nor UO_246 (O_246,N_14718,N_14027);
nand UO_247 (O_247,N_14895,N_14732);
nor UO_248 (O_248,N_14270,N_14187);
xnor UO_249 (O_249,N_14465,N_14180);
and UO_250 (O_250,N_14321,N_14173);
nor UO_251 (O_251,N_14954,N_14970);
and UO_252 (O_252,N_14258,N_14689);
and UO_253 (O_253,N_14760,N_14074);
or UO_254 (O_254,N_14326,N_14291);
and UO_255 (O_255,N_14206,N_14328);
nor UO_256 (O_256,N_14260,N_14278);
and UO_257 (O_257,N_14564,N_14468);
and UO_258 (O_258,N_14622,N_14580);
and UO_259 (O_259,N_14513,N_14722);
nor UO_260 (O_260,N_14955,N_14783);
nand UO_261 (O_261,N_14357,N_14314);
nor UO_262 (O_262,N_14221,N_14334);
nor UO_263 (O_263,N_14591,N_14747);
xnor UO_264 (O_264,N_14062,N_14254);
xnor UO_265 (O_265,N_14190,N_14804);
nor UO_266 (O_266,N_14145,N_14359);
nand UO_267 (O_267,N_14517,N_14553);
nand UO_268 (O_268,N_14682,N_14112);
and UO_269 (O_269,N_14455,N_14515);
nor UO_270 (O_270,N_14183,N_14984);
nand UO_271 (O_271,N_14941,N_14988);
and UO_272 (O_272,N_14807,N_14390);
nor UO_273 (O_273,N_14945,N_14209);
nor UO_274 (O_274,N_14670,N_14146);
or UO_275 (O_275,N_14083,N_14952);
nand UO_276 (O_276,N_14950,N_14648);
and UO_277 (O_277,N_14600,N_14781);
and UO_278 (O_278,N_14409,N_14401);
xnor UO_279 (O_279,N_14113,N_14102);
nor UO_280 (O_280,N_14156,N_14096);
and UO_281 (O_281,N_14415,N_14161);
nor UO_282 (O_282,N_14038,N_14576);
and UO_283 (O_283,N_14788,N_14794);
nand UO_284 (O_284,N_14151,N_14046);
nor UO_285 (O_285,N_14870,N_14916);
or UO_286 (O_286,N_14327,N_14669);
nor UO_287 (O_287,N_14656,N_14658);
nand UO_288 (O_288,N_14242,N_14163);
and UO_289 (O_289,N_14262,N_14111);
nor UO_290 (O_290,N_14094,N_14506);
nor UO_291 (O_291,N_14475,N_14778);
nor UO_292 (O_292,N_14008,N_14128);
and UO_293 (O_293,N_14386,N_14020);
nand UO_294 (O_294,N_14373,N_14606);
nand UO_295 (O_295,N_14117,N_14654);
and UO_296 (O_296,N_14329,N_14155);
and UO_297 (O_297,N_14741,N_14820);
and UO_298 (O_298,N_14430,N_14725);
and UO_299 (O_299,N_14546,N_14628);
nor UO_300 (O_300,N_14263,N_14896);
nand UO_301 (O_301,N_14925,N_14396);
nand UO_302 (O_302,N_14014,N_14073);
xor UO_303 (O_303,N_14615,N_14529);
and UO_304 (O_304,N_14489,N_14474);
nor UO_305 (O_305,N_14205,N_14054);
and UO_306 (O_306,N_14157,N_14166);
nor UO_307 (O_307,N_14219,N_14676);
nor UO_308 (O_308,N_14894,N_14602);
nand UO_309 (O_309,N_14691,N_14892);
nand UO_310 (O_310,N_14857,N_14651);
nor UO_311 (O_311,N_14011,N_14801);
nor UO_312 (O_312,N_14421,N_14460);
and UO_313 (O_313,N_14449,N_14158);
xnor UO_314 (O_314,N_14977,N_14583);
and UO_315 (O_315,N_14088,N_14045);
or UO_316 (O_316,N_14379,N_14542);
nor UO_317 (O_317,N_14084,N_14905);
or UO_318 (O_318,N_14929,N_14467);
and UO_319 (O_319,N_14234,N_14815);
and UO_320 (O_320,N_14053,N_14685);
and UO_321 (O_321,N_14443,N_14501);
nand UO_322 (O_322,N_14860,N_14198);
or UO_323 (O_323,N_14805,N_14025);
or UO_324 (O_324,N_14036,N_14723);
or UO_325 (O_325,N_14978,N_14264);
and UO_326 (O_326,N_14391,N_14268);
or UO_327 (O_327,N_14627,N_14793);
and UO_328 (O_328,N_14549,N_14541);
or UO_329 (O_329,N_14902,N_14828);
and UO_330 (O_330,N_14575,N_14039);
nand UO_331 (O_331,N_14610,N_14322);
nor UO_332 (O_332,N_14624,N_14523);
and UO_333 (O_333,N_14476,N_14129);
or UO_334 (O_334,N_14972,N_14285);
nand UO_335 (O_335,N_14301,N_14458);
or UO_336 (O_336,N_14806,N_14439);
or UO_337 (O_337,N_14566,N_14769);
and UO_338 (O_338,N_14132,N_14310);
and UO_339 (O_339,N_14100,N_14267);
xor UO_340 (O_340,N_14337,N_14765);
nor UO_341 (O_341,N_14713,N_14834);
or UO_342 (O_342,N_14880,N_14948);
and UO_343 (O_343,N_14414,N_14207);
or UO_344 (O_344,N_14833,N_14211);
or UO_345 (O_345,N_14843,N_14114);
nand UO_346 (O_346,N_14848,N_14824);
nand UO_347 (O_347,N_14923,N_14323);
nand UO_348 (O_348,N_14835,N_14561);
or UO_349 (O_349,N_14961,N_14728);
nor UO_350 (O_350,N_14360,N_14487);
or UO_351 (O_351,N_14876,N_14002);
nor UO_352 (O_352,N_14683,N_14280);
nand UO_353 (O_353,N_14013,N_14629);
and UO_354 (O_354,N_14695,N_14665);
and UO_355 (O_355,N_14105,N_14230);
nor UO_356 (O_356,N_14358,N_14369);
nor UO_357 (O_357,N_14995,N_14758);
or UO_358 (O_358,N_14217,N_14724);
or UO_359 (O_359,N_14784,N_14708);
or UO_360 (O_360,N_14406,N_14601);
nand UO_361 (O_361,N_14530,N_14963);
or UO_362 (O_362,N_14814,N_14809);
or UO_363 (O_363,N_14089,N_14227);
and UO_364 (O_364,N_14756,N_14277);
nor UO_365 (O_365,N_14882,N_14005);
nor UO_366 (O_366,N_14296,N_14376);
or UO_367 (O_367,N_14551,N_14808);
nor UO_368 (O_368,N_14186,N_14165);
nand UO_369 (O_369,N_14208,N_14768);
or UO_370 (O_370,N_14248,N_14987);
nand UO_371 (O_371,N_14904,N_14767);
and UO_372 (O_372,N_14441,N_14939);
xor UO_373 (O_373,N_14521,N_14418);
nor UO_374 (O_374,N_14498,N_14650);
and UO_375 (O_375,N_14912,N_14621);
nor UO_376 (O_376,N_14473,N_14680);
or UO_377 (O_377,N_14681,N_14632);
nand UO_378 (O_378,N_14803,N_14298);
or UO_379 (O_379,N_14720,N_14346);
nor UO_380 (O_380,N_14619,N_14565);
nand UO_381 (O_381,N_14351,N_14836);
or UO_382 (O_382,N_14638,N_14266);
and UO_383 (O_383,N_14246,N_14742);
or UO_384 (O_384,N_14104,N_14068);
and UO_385 (O_385,N_14554,N_14245);
nor UO_386 (O_386,N_14461,N_14759);
xnor UO_387 (O_387,N_14625,N_14059);
nor UO_388 (O_388,N_14636,N_14697);
and UO_389 (O_389,N_14556,N_14611);
nand UO_390 (O_390,N_14639,N_14075);
nand UO_391 (O_391,N_14678,N_14222);
and UO_392 (O_392,N_14437,N_14250);
or UO_393 (O_393,N_14303,N_14232);
and UO_394 (O_394,N_14618,N_14634);
xnor UO_395 (O_395,N_14385,N_14933);
or UO_396 (O_396,N_14813,N_14528);
nor UO_397 (O_397,N_14822,N_14849);
nand UO_398 (O_398,N_14953,N_14381);
or UO_399 (O_399,N_14975,N_14235);
or UO_400 (O_400,N_14495,N_14286);
nor UO_401 (O_401,N_14177,N_14577);
or UO_402 (O_402,N_14444,N_14315);
nor UO_403 (O_403,N_14347,N_14047);
nand UO_404 (O_404,N_14051,N_14862);
nand UO_405 (O_405,N_14078,N_14308);
xnor UO_406 (O_406,N_14249,N_14776);
or UO_407 (O_407,N_14252,N_14167);
and UO_408 (O_408,N_14108,N_14771);
nand UO_409 (O_409,N_14387,N_14271);
nor UO_410 (O_410,N_14294,N_14937);
and UO_411 (O_411,N_14341,N_14478);
nor UO_412 (O_412,N_14133,N_14917);
nand UO_413 (O_413,N_14049,N_14579);
or UO_414 (O_414,N_14284,N_14859);
xor UO_415 (O_415,N_14500,N_14947);
nor UO_416 (O_416,N_14090,N_14091);
nor UO_417 (O_417,N_14897,N_14707);
nor UO_418 (O_418,N_14139,N_14138);
nand UO_419 (O_419,N_14702,N_14544);
or UO_420 (O_420,N_14560,N_14050);
xnor UO_421 (O_421,N_14118,N_14889);
nor UO_422 (O_422,N_14124,N_14861);
xor UO_423 (O_423,N_14035,N_14356);
nor UO_424 (O_424,N_14598,N_14201);
or UO_425 (O_425,N_14906,N_14800);
or UO_426 (O_426,N_14775,N_14297);
and UO_427 (O_427,N_14302,N_14726);
or UO_428 (O_428,N_14729,N_14407);
or UO_429 (O_429,N_14739,N_14332);
nand UO_430 (O_430,N_14363,N_14015);
or UO_431 (O_431,N_14919,N_14959);
and UO_432 (O_432,N_14692,N_14017);
nor UO_433 (O_433,N_14596,N_14976);
nor UO_434 (O_434,N_14178,N_14214);
nor UO_435 (O_435,N_14907,N_14395);
or UO_436 (O_436,N_14875,N_14830);
and UO_437 (O_437,N_14324,N_14829);
or UO_438 (O_438,N_14365,N_14690);
nor UO_439 (O_439,N_14653,N_14010);
nand UO_440 (O_440,N_14431,N_14330);
or UO_441 (O_441,N_14761,N_14502);
and UO_442 (O_442,N_14754,N_14703);
and UO_443 (O_443,N_14980,N_14934);
or UO_444 (O_444,N_14394,N_14153);
or UO_445 (O_445,N_14645,N_14371);
nor UO_446 (O_446,N_14416,N_14992);
and UO_447 (O_447,N_14819,N_14306);
and UO_448 (O_448,N_14354,N_14942);
nor UO_449 (O_449,N_14991,N_14614);
nand UO_450 (O_450,N_14659,N_14548);
nor UO_451 (O_451,N_14170,N_14032);
nor UO_452 (O_452,N_14755,N_14714);
nand UO_453 (O_453,N_14935,N_14673);
nor UO_454 (O_454,N_14446,N_14231);
nor UO_455 (O_455,N_14392,N_14480);
or UO_456 (O_456,N_14817,N_14456);
xor UO_457 (O_457,N_14900,N_14413);
nor UO_458 (O_458,N_14144,N_14743);
nand UO_459 (O_459,N_14524,N_14944);
nand UO_460 (O_460,N_14295,N_14990);
and UO_461 (O_461,N_14609,N_14004);
nand UO_462 (O_462,N_14335,N_14717);
or UO_463 (O_463,N_14746,N_14550);
xnor UO_464 (O_464,N_14127,N_14040);
nand UO_465 (O_465,N_14464,N_14236);
and UO_466 (O_466,N_14316,N_14107);
or UO_467 (O_467,N_14159,N_14974);
xnor UO_468 (O_468,N_14700,N_14590);
nand UO_469 (O_469,N_14003,N_14514);
and UO_470 (O_470,N_14881,N_14507);
xnor UO_471 (O_471,N_14997,N_14085);
nor UO_472 (O_472,N_14535,N_14631);
and UO_473 (O_473,N_14505,N_14552);
nand UO_474 (O_474,N_14143,N_14194);
nor UO_475 (O_475,N_14927,N_14125);
and UO_476 (O_476,N_14001,N_14261);
nand UO_477 (O_477,N_14361,N_14410);
xnor UO_478 (O_478,N_14568,N_14774);
or UO_479 (O_479,N_14065,N_14433);
xnor UO_480 (O_480,N_14525,N_14481);
nor UO_481 (O_481,N_14701,N_14071);
nor UO_482 (O_482,N_14425,N_14750);
or UO_483 (O_483,N_14931,N_14949);
nand UO_484 (O_484,N_14450,N_14884);
or UO_485 (O_485,N_14883,N_14463);
nand UO_486 (O_486,N_14081,N_14192);
and UO_487 (O_487,N_14239,N_14620);
nor UO_488 (O_488,N_14350,N_14240);
nand UO_489 (O_489,N_14229,N_14637);
nand UO_490 (O_490,N_14311,N_14012);
xnor UO_491 (O_491,N_14831,N_14969);
and UO_492 (O_492,N_14043,N_14913);
or UO_493 (O_493,N_14382,N_14667);
or UO_494 (O_494,N_14006,N_14766);
nand UO_495 (O_495,N_14427,N_14185);
nand UO_496 (O_496,N_14635,N_14688);
nand UO_497 (O_497,N_14016,N_14527);
nor UO_498 (O_498,N_14220,N_14063);
nor UO_499 (O_499,N_14721,N_14994);
nand UO_500 (O_500,N_14993,N_14893);
or UO_501 (O_501,N_14867,N_14802);
nand UO_502 (O_502,N_14066,N_14996);
nand UO_503 (O_503,N_14851,N_14405);
xor UO_504 (O_504,N_14905,N_14951);
nor UO_505 (O_505,N_14174,N_14385);
or UO_506 (O_506,N_14114,N_14712);
nor UO_507 (O_507,N_14721,N_14776);
nor UO_508 (O_508,N_14015,N_14904);
nor UO_509 (O_509,N_14539,N_14687);
nor UO_510 (O_510,N_14025,N_14966);
or UO_511 (O_511,N_14110,N_14580);
xnor UO_512 (O_512,N_14598,N_14345);
nand UO_513 (O_513,N_14293,N_14773);
and UO_514 (O_514,N_14088,N_14564);
or UO_515 (O_515,N_14886,N_14610);
nand UO_516 (O_516,N_14239,N_14971);
and UO_517 (O_517,N_14780,N_14475);
and UO_518 (O_518,N_14372,N_14159);
nand UO_519 (O_519,N_14762,N_14719);
and UO_520 (O_520,N_14384,N_14054);
nand UO_521 (O_521,N_14362,N_14742);
nor UO_522 (O_522,N_14250,N_14640);
and UO_523 (O_523,N_14683,N_14313);
nor UO_524 (O_524,N_14075,N_14191);
or UO_525 (O_525,N_14351,N_14434);
nand UO_526 (O_526,N_14073,N_14693);
and UO_527 (O_527,N_14652,N_14204);
nand UO_528 (O_528,N_14822,N_14140);
nor UO_529 (O_529,N_14068,N_14557);
and UO_530 (O_530,N_14200,N_14314);
nor UO_531 (O_531,N_14642,N_14369);
nor UO_532 (O_532,N_14624,N_14287);
nor UO_533 (O_533,N_14013,N_14767);
and UO_534 (O_534,N_14425,N_14942);
or UO_535 (O_535,N_14215,N_14721);
nor UO_536 (O_536,N_14683,N_14080);
nand UO_537 (O_537,N_14505,N_14376);
and UO_538 (O_538,N_14217,N_14494);
nor UO_539 (O_539,N_14550,N_14626);
xnor UO_540 (O_540,N_14511,N_14397);
and UO_541 (O_541,N_14670,N_14317);
nand UO_542 (O_542,N_14218,N_14006);
or UO_543 (O_543,N_14963,N_14375);
and UO_544 (O_544,N_14251,N_14925);
xnor UO_545 (O_545,N_14815,N_14991);
nand UO_546 (O_546,N_14778,N_14730);
nor UO_547 (O_547,N_14774,N_14250);
or UO_548 (O_548,N_14614,N_14628);
and UO_549 (O_549,N_14162,N_14090);
nor UO_550 (O_550,N_14325,N_14324);
nand UO_551 (O_551,N_14992,N_14515);
nor UO_552 (O_552,N_14323,N_14156);
nand UO_553 (O_553,N_14185,N_14400);
nand UO_554 (O_554,N_14941,N_14104);
nor UO_555 (O_555,N_14265,N_14353);
and UO_556 (O_556,N_14484,N_14527);
or UO_557 (O_557,N_14136,N_14862);
and UO_558 (O_558,N_14591,N_14472);
nand UO_559 (O_559,N_14572,N_14796);
or UO_560 (O_560,N_14028,N_14953);
and UO_561 (O_561,N_14169,N_14849);
and UO_562 (O_562,N_14515,N_14983);
and UO_563 (O_563,N_14170,N_14104);
or UO_564 (O_564,N_14134,N_14727);
nand UO_565 (O_565,N_14761,N_14034);
nor UO_566 (O_566,N_14408,N_14552);
nand UO_567 (O_567,N_14208,N_14107);
nand UO_568 (O_568,N_14942,N_14064);
nand UO_569 (O_569,N_14179,N_14238);
nor UO_570 (O_570,N_14798,N_14046);
nor UO_571 (O_571,N_14524,N_14336);
or UO_572 (O_572,N_14786,N_14238);
xnor UO_573 (O_573,N_14791,N_14216);
or UO_574 (O_574,N_14748,N_14820);
nor UO_575 (O_575,N_14113,N_14138);
and UO_576 (O_576,N_14320,N_14758);
xnor UO_577 (O_577,N_14557,N_14719);
nand UO_578 (O_578,N_14917,N_14533);
nand UO_579 (O_579,N_14795,N_14992);
or UO_580 (O_580,N_14940,N_14486);
nor UO_581 (O_581,N_14509,N_14984);
nor UO_582 (O_582,N_14046,N_14915);
and UO_583 (O_583,N_14714,N_14185);
and UO_584 (O_584,N_14295,N_14889);
xor UO_585 (O_585,N_14505,N_14922);
nand UO_586 (O_586,N_14641,N_14068);
nand UO_587 (O_587,N_14777,N_14898);
and UO_588 (O_588,N_14702,N_14976);
xor UO_589 (O_589,N_14914,N_14121);
or UO_590 (O_590,N_14696,N_14457);
or UO_591 (O_591,N_14645,N_14227);
and UO_592 (O_592,N_14254,N_14500);
nand UO_593 (O_593,N_14931,N_14658);
or UO_594 (O_594,N_14772,N_14557);
nand UO_595 (O_595,N_14450,N_14828);
and UO_596 (O_596,N_14791,N_14770);
xor UO_597 (O_597,N_14844,N_14247);
and UO_598 (O_598,N_14223,N_14085);
nand UO_599 (O_599,N_14581,N_14892);
nand UO_600 (O_600,N_14895,N_14483);
or UO_601 (O_601,N_14067,N_14371);
or UO_602 (O_602,N_14849,N_14906);
nand UO_603 (O_603,N_14825,N_14708);
and UO_604 (O_604,N_14247,N_14051);
nor UO_605 (O_605,N_14719,N_14732);
or UO_606 (O_606,N_14073,N_14623);
and UO_607 (O_607,N_14685,N_14442);
nor UO_608 (O_608,N_14354,N_14521);
nor UO_609 (O_609,N_14797,N_14497);
nor UO_610 (O_610,N_14284,N_14444);
or UO_611 (O_611,N_14243,N_14458);
and UO_612 (O_612,N_14220,N_14362);
nor UO_613 (O_613,N_14672,N_14079);
and UO_614 (O_614,N_14065,N_14577);
and UO_615 (O_615,N_14718,N_14880);
nor UO_616 (O_616,N_14604,N_14017);
xor UO_617 (O_617,N_14698,N_14399);
nand UO_618 (O_618,N_14244,N_14566);
nand UO_619 (O_619,N_14621,N_14335);
or UO_620 (O_620,N_14382,N_14072);
nor UO_621 (O_621,N_14170,N_14405);
nor UO_622 (O_622,N_14516,N_14401);
nand UO_623 (O_623,N_14960,N_14411);
or UO_624 (O_624,N_14595,N_14216);
nor UO_625 (O_625,N_14624,N_14833);
or UO_626 (O_626,N_14225,N_14272);
nor UO_627 (O_627,N_14744,N_14242);
nor UO_628 (O_628,N_14019,N_14255);
nor UO_629 (O_629,N_14932,N_14869);
xnor UO_630 (O_630,N_14996,N_14515);
or UO_631 (O_631,N_14316,N_14056);
nand UO_632 (O_632,N_14405,N_14763);
nor UO_633 (O_633,N_14919,N_14072);
nand UO_634 (O_634,N_14369,N_14629);
and UO_635 (O_635,N_14036,N_14061);
nand UO_636 (O_636,N_14703,N_14430);
and UO_637 (O_637,N_14496,N_14762);
and UO_638 (O_638,N_14455,N_14078);
or UO_639 (O_639,N_14690,N_14310);
nand UO_640 (O_640,N_14371,N_14843);
and UO_641 (O_641,N_14116,N_14478);
xnor UO_642 (O_642,N_14131,N_14182);
or UO_643 (O_643,N_14626,N_14304);
nand UO_644 (O_644,N_14123,N_14318);
nand UO_645 (O_645,N_14408,N_14901);
or UO_646 (O_646,N_14590,N_14324);
or UO_647 (O_647,N_14926,N_14584);
nor UO_648 (O_648,N_14735,N_14612);
xnor UO_649 (O_649,N_14120,N_14313);
nor UO_650 (O_650,N_14146,N_14620);
or UO_651 (O_651,N_14277,N_14039);
or UO_652 (O_652,N_14951,N_14044);
and UO_653 (O_653,N_14808,N_14519);
and UO_654 (O_654,N_14661,N_14453);
xor UO_655 (O_655,N_14626,N_14371);
and UO_656 (O_656,N_14344,N_14623);
nor UO_657 (O_657,N_14427,N_14504);
nand UO_658 (O_658,N_14357,N_14918);
nor UO_659 (O_659,N_14419,N_14664);
or UO_660 (O_660,N_14076,N_14939);
nor UO_661 (O_661,N_14325,N_14024);
and UO_662 (O_662,N_14171,N_14553);
or UO_663 (O_663,N_14767,N_14711);
nor UO_664 (O_664,N_14376,N_14507);
nor UO_665 (O_665,N_14927,N_14299);
nor UO_666 (O_666,N_14225,N_14943);
xnor UO_667 (O_667,N_14396,N_14449);
xor UO_668 (O_668,N_14147,N_14080);
and UO_669 (O_669,N_14697,N_14545);
or UO_670 (O_670,N_14914,N_14202);
nand UO_671 (O_671,N_14354,N_14127);
or UO_672 (O_672,N_14323,N_14130);
or UO_673 (O_673,N_14174,N_14031);
nand UO_674 (O_674,N_14073,N_14219);
and UO_675 (O_675,N_14908,N_14869);
or UO_676 (O_676,N_14839,N_14512);
and UO_677 (O_677,N_14007,N_14726);
nor UO_678 (O_678,N_14402,N_14154);
nor UO_679 (O_679,N_14008,N_14310);
nor UO_680 (O_680,N_14501,N_14953);
and UO_681 (O_681,N_14229,N_14803);
xor UO_682 (O_682,N_14242,N_14573);
nand UO_683 (O_683,N_14549,N_14644);
and UO_684 (O_684,N_14490,N_14547);
or UO_685 (O_685,N_14682,N_14443);
nand UO_686 (O_686,N_14553,N_14025);
and UO_687 (O_687,N_14012,N_14948);
or UO_688 (O_688,N_14789,N_14615);
xor UO_689 (O_689,N_14430,N_14520);
and UO_690 (O_690,N_14381,N_14872);
or UO_691 (O_691,N_14075,N_14085);
or UO_692 (O_692,N_14370,N_14762);
nor UO_693 (O_693,N_14448,N_14123);
or UO_694 (O_694,N_14518,N_14609);
nand UO_695 (O_695,N_14469,N_14027);
nor UO_696 (O_696,N_14095,N_14603);
and UO_697 (O_697,N_14036,N_14697);
or UO_698 (O_698,N_14017,N_14021);
and UO_699 (O_699,N_14678,N_14475);
or UO_700 (O_700,N_14198,N_14386);
or UO_701 (O_701,N_14956,N_14759);
nor UO_702 (O_702,N_14983,N_14735);
xor UO_703 (O_703,N_14765,N_14984);
nor UO_704 (O_704,N_14283,N_14008);
or UO_705 (O_705,N_14494,N_14210);
or UO_706 (O_706,N_14947,N_14807);
xor UO_707 (O_707,N_14920,N_14509);
nand UO_708 (O_708,N_14993,N_14939);
xor UO_709 (O_709,N_14235,N_14678);
or UO_710 (O_710,N_14850,N_14145);
nor UO_711 (O_711,N_14962,N_14890);
nor UO_712 (O_712,N_14080,N_14415);
and UO_713 (O_713,N_14362,N_14880);
and UO_714 (O_714,N_14528,N_14853);
and UO_715 (O_715,N_14645,N_14085);
and UO_716 (O_716,N_14934,N_14899);
nand UO_717 (O_717,N_14793,N_14239);
nor UO_718 (O_718,N_14912,N_14469);
nand UO_719 (O_719,N_14888,N_14369);
and UO_720 (O_720,N_14053,N_14728);
and UO_721 (O_721,N_14075,N_14528);
or UO_722 (O_722,N_14756,N_14064);
xnor UO_723 (O_723,N_14241,N_14159);
nor UO_724 (O_724,N_14588,N_14491);
nand UO_725 (O_725,N_14639,N_14311);
nor UO_726 (O_726,N_14921,N_14757);
nand UO_727 (O_727,N_14825,N_14466);
nand UO_728 (O_728,N_14502,N_14394);
and UO_729 (O_729,N_14653,N_14173);
nand UO_730 (O_730,N_14249,N_14913);
nand UO_731 (O_731,N_14861,N_14867);
nor UO_732 (O_732,N_14274,N_14332);
or UO_733 (O_733,N_14491,N_14297);
nor UO_734 (O_734,N_14663,N_14448);
and UO_735 (O_735,N_14156,N_14547);
nor UO_736 (O_736,N_14572,N_14552);
nand UO_737 (O_737,N_14818,N_14822);
nor UO_738 (O_738,N_14451,N_14562);
or UO_739 (O_739,N_14771,N_14587);
and UO_740 (O_740,N_14041,N_14063);
nand UO_741 (O_741,N_14008,N_14850);
xor UO_742 (O_742,N_14574,N_14749);
and UO_743 (O_743,N_14479,N_14620);
nor UO_744 (O_744,N_14221,N_14144);
nor UO_745 (O_745,N_14233,N_14917);
nor UO_746 (O_746,N_14346,N_14911);
nor UO_747 (O_747,N_14757,N_14232);
nor UO_748 (O_748,N_14121,N_14979);
or UO_749 (O_749,N_14427,N_14021);
xnor UO_750 (O_750,N_14224,N_14473);
and UO_751 (O_751,N_14032,N_14008);
nor UO_752 (O_752,N_14368,N_14629);
nand UO_753 (O_753,N_14938,N_14078);
xnor UO_754 (O_754,N_14497,N_14945);
nand UO_755 (O_755,N_14467,N_14105);
xnor UO_756 (O_756,N_14101,N_14635);
or UO_757 (O_757,N_14643,N_14038);
or UO_758 (O_758,N_14969,N_14214);
nor UO_759 (O_759,N_14851,N_14199);
nand UO_760 (O_760,N_14270,N_14463);
or UO_761 (O_761,N_14583,N_14460);
nor UO_762 (O_762,N_14228,N_14653);
xor UO_763 (O_763,N_14430,N_14835);
xnor UO_764 (O_764,N_14772,N_14381);
nor UO_765 (O_765,N_14057,N_14247);
nand UO_766 (O_766,N_14813,N_14737);
or UO_767 (O_767,N_14073,N_14715);
and UO_768 (O_768,N_14082,N_14739);
nor UO_769 (O_769,N_14149,N_14964);
or UO_770 (O_770,N_14685,N_14839);
and UO_771 (O_771,N_14660,N_14567);
or UO_772 (O_772,N_14256,N_14734);
or UO_773 (O_773,N_14378,N_14751);
and UO_774 (O_774,N_14683,N_14239);
xor UO_775 (O_775,N_14664,N_14000);
nor UO_776 (O_776,N_14298,N_14029);
xnor UO_777 (O_777,N_14617,N_14555);
or UO_778 (O_778,N_14737,N_14336);
and UO_779 (O_779,N_14515,N_14304);
nor UO_780 (O_780,N_14526,N_14344);
or UO_781 (O_781,N_14855,N_14084);
xor UO_782 (O_782,N_14770,N_14004);
or UO_783 (O_783,N_14002,N_14654);
nand UO_784 (O_784,N_14542,N_14221);
or UO_785 (O_785,N_14343,N_14322);
xnor UO_786 (O_786,N_14991,N_14411);
and UO_787 (O_787,N_14273,N_14521);
and UO_788 (O_788,N_14222,N_14645);
nand UO_789 (O_789,N_14999,N_14822);
or UO_790 (O_790,N_14299,N_14283);
and UO_791 (O_791,N_14236,N_14303);
or UO_792 (O_792,N_14474,N_14426);
nor UO_793 (O_793,N_14037,N_14320);
nor UO_794 (O_794,N_14483,N_14644);
nor UO_795 (O_795,N_14359,N_14028);
nand UO_796 (O_796,N_14572,N_14805);
nand UO_797 (O_797,N_14078,N_14287);
nor UO_798 (O_798,N_14511,N_14572);
and UO_799 (O_799,N_14478,N_14804);
nor UO_800 (O_800,N_14369,N_14174);
and UO_801 (O_801,N_14693,N_14356);
or UO_802 (O_802,N_14498,N_14547);
or UO_803 (O_803,N_14604,N_14028);
nand UO_804 (O_804,N_14409,N_14823);
or UO_805 (O_805,N_14688,N_14658);
or UO_806 (O_806,N_14322,N_14903);
or UO_807 (O_807,N_14835,N_14745);
nand UO_808 (O_808,N_14344,N_14546);
or UO_809 (O_809,N_14609,N_14338);
or UO_810 (O_810,N_14763,N_14963);
and UO_811 (O_811,N_14911,N_14521);
and UO_812 (O_812,N_14916,N_14657);
nand UO_813 (O_813,N_14276,N_14494);
nor UO_814 (O_814,N_14635,N_14444);
nor UO_815 (O_815,N_14714,N_14912);
or UO_816 (O_816,N_14423,N_14633);
and UO_817 (O_817,N_14378,N_14439);
nand UO_818 (O_818,N_14964,N_14809);
nand UO_819 (O_819,N_14567,N_14600);
and UO_820 (O_820,N_14761,N_14155);
and UO_821 (O_821,N_14525,N_14603);
or UO_822 (O_822,N_14820,N_14182);
or UO_823 (O_823,N_14314,N_14172);
and UO_824 (O_824,N_14154,N_14842);
and UO_825 (O_825,N_14113,N_14812);
xor UO_826 (O_826,N_14677,N_14345);
nor UO_827 (O_827,N_14508,N_14208);
and UO_828 (O_828,N_14424,N_14470);
or UO_829 (O_829,N_14805,N_14315);
and UO_830 (O_830,N_14001,N_14407);
xnor UO_831 (O_831,N_14426,N_14260);
and UO_832 (O_832,N_14154,N_14713);
and UO_833 (O_833,N_14436,N_14676);
nand UO_834 (O_834,N_14237,N_14933);
nor UO_835 (O_835,N_14520,N_14248);
nand UO_836 (O_836,N_14067,N_14002);
nand UO_837 (O_837,N_14749,N_14742);
or UO_838 (O_838,N_14182,N_14064);
nor UO_839 (O_839,N_14199,N_14945);
or UO_840 (O_840,N_14502,N_14039);
nor UO_841 (O_841,N_14350,N_14883);
or UO_842 (O_842,N_14017,N_14970);
or UO_843 (O_843,N_14776,N_14691);
and UO_844 (O_844,N_14227,N_14925);
nor UO_845 (O_845,N_14291,N_14105);
nor UO_846 (O_846,N_14513,N_14944);
xor UO_847 (O_847,N_14090,N_14243);
nand UO_848 (O_848,N_14877,N_14357);
nand UO_849 (O_849,N_14552,N_14507);
or UO_850 (O_850,N_14663,N_14804);
nor UO_851 (O_851,N_14482,N_14643);
nand UO_852 (O_852,N_14123,N_14558);
nor UO_853 (O_853,N_14496,N_14466);
and UO_854 (O_854,N_14139,N_14801);
and UO_855 (O_855,N_14929,N_14232);
nand UO_856 (O_856,N_14374,N_14071);
nand UO_857 (O_857,N_14591,N_14300);
xor UO_858 (O_858,N_14337,N_14307);
nand UO_859 (O_859,N_14935,N_14890);
nor UO_860 (O_860,N_14804,N_14047);
nand UO_861 (O_861,N_14369,N_14727);
nor UO_862 (O_862,N_14805,N_14124);
nand UO_863 (O_863,N_14447,N_14560);
nor UO_864 (O_864,N_14235,N_14752);
nand UO_865 (O_865,N_14673,N_14624);
or UO_866 (O_866,N_14057,N_14543);
or UO_867 (O_867,N_14509,N_14302);
and UO_868 (O_868,N_14034,N_14422);
nor UO_869 (O_869,N_14172,N_14037);
or UO_870 (O_870,N_14141,N_14518);
and UO_871 (O_871,N_14560,N_14720);
or UO_872 (O_872,N_14238,N_14950);
or UO_873 (O_873,N_14065,N_14774);
and UO_874 (O_874,N_14893,N_14688);
and UO_875 (O_875,N_14947,N_14605);
and UO_876 (O_876,N_14751,N_14810);
or UO_877 (O_877,N_14275,N_14893);
nor UO_878 (O_878,N_14429,N_14261);
xnor UO_879 (O_879,N_14009,N_14658);
nand UO_880 (O_880,N_14397,N_14007);
xnor UO_881 (O_881,N_14516,N_14864);
nor UO_882 (O_882,N_14986,N_14439);
and UO_883 (O_883,N_14293,N_14475);
nor UO_884 (O_884,N_14171,N_14492);
or UO_885 (O_885,N_14432,N_14419);
nor UO_886 (O_886,N_14644,N_14726);
xnor UO_887 (O_887,N_14341,N_14650);
nand UO_888 (O_888,N_14993,N_14808);
or UO_889 (O_889,N_14777,N_14238);
or UO_890 (O_890,N_14468,N_14429);
nor UO_891 (O_891,N_14769,N_14534);
nand UO_892 (O_892,N_14883,N_14492);
xor UO_893 (O_893,N_14990,N_14123);
xnor UO_894 (O_894,N_14999,N_14481);
and UO_895 (O_895,N_14889,N_14061);
and UO_896 (O_896,N_14591,N_14169);
nand UO_897 (O_897,N_14549,N_14372);
nor UO_898 (O_898,N_14889,N_14005);
xnor UO_899 (O_899,N_14768,N_14224);
and UO_900 (O_900,N_14875,N_14693);
nor UO_901 (O_901,N_14386,N_14123);
nor UO_902 (O_902,N_14591,N_14164);
or UO_903 (O_903,N_14045,N_14435);
nand UO_904 (O_904,N_14537,N_14664);
nand UO_905 (O_905,N_14500,N_14613);
or UO_906 (O_906,N_14508,N_14108);
and UO_907 (O_907,N_14085,N_14312);
nor UO_908 (O_908,N_14322,N_14719);
nor UO_909 (O_909,N_14228,N_14789);
nand UO_910 (O_910,N_14854,N_14149);
or UO_911 (O_911,N_14297,N_14133);
nand UO_912 (O_912,N_14539,N_14682);
nor UO_913 (O_913,N_14995,N_14704);
nand UO_914 (O_914,N_14766,N_14031);
and UO_915 (O_915,N_14538,N_14617);
or UO_916 (O_916,N_14238,N_14410);
and UO_917 (O_917,N_14656,N_14158);
and UO_918 (O_918,N_14335,N_14366);
xor UO_919 (O_919,N_14258,N_14274);
xnor UO_920 (O_920,N_14132,N_14923);
nand UO_921 (O_921,N_14865,N_14488);
nand UO_922 (O_922,N_14935,N_14543);
nor UO_923 (O_923,N_14008,N_14950);
nor UO_924 (O_924,N_14743,N_14250);
nand UO_925 (O_925,N_14254,N_14304);
nor UO_926 (O_926,N_14882,N_14122);
nor UO_927 (O_927,N_14623,N_14151);
nand UO_928 (O_928,N_14562,N_14495);
xor UO_929 (O_929,N_14794,N_14077);
and UO_930 (O_930,N_14447,N_14845);
or UO_931 (O_931,N_14924,N_14957);
xor UO_932 (O_932,N_14689,N_14184);
nand UO_933 (O_933,N_14996,N_14628);
and UO_934 (O_934,N_14630,N_14389);
and UO_935 (O_935,N_14297,N_14748);
and UO_936 (O_936,N_14086,N_14153);
or UO_937 (O_937,N_14568,N_14239);
and UO_938 (O_938,N_14666,N_14087);
nand UO_939 (O_939,N_14220,N_14606);
nand UO_940 (O_940,N_14181,N_14163);
or UO_941 (O_941,N_14699,N_14417);
and UO_942 (O_942,N_14412,N_14193);
nor UO_943 (O_943,N_14045,N_14224);
or UO_944 (O_944,N_14851,N_14599);
nor UO_945 (O_945,N_14637,N_14488);
nand UO_946 (O_946,N_14593,N_14862);
or UO_947 (O_947,N_14694,N_14026);
and UO_948 (O_948,N_14823,N_14499);
and UO_949 (O_949,N_14857,N_14989);
and UO_950 (O_950,N_14292,N_14093);
nor UO_951 (O_951,N_14431,N_14838);
nor UO_952 (O_952,N_14794,N_14471);
nand UO_953 (O_953,N_14354,N_14599);
or UO_954 (O_954,N_14889,N_14743);
nand UO_955 (O_955,N_14405,N_14849);
xor UO_956 (O_956,N_14548,N_14349);
nand UO_957 (O_957,N_14046,N_14543);
and UO_958 (O_958,N_14847,N_14791);
xor UO_959 (O_959,N_14715,N_14565);
nor UO_960 (O_960,N_14844,N_14240);
nand UO_961 (O_961,N_14459,N_14244);
nor UO_962 (O_962,N_14196,N_14018);
nand UO_963 (O_963,N_14692,N_14025);
and UO_964 (O_964,N_14566,N_14255);
nand UO_965 (O_965,N_14366,N_14615);
and UO_966 (O_966,N_14678,N_14446);
nand UO_967 (O_967,N_14390,N_14247);
nor UO_968 (O_968,N_14284,N_14934);
and UO_969 (O_969,N_14514,N_14319);
nand UO_970 (O_970,N_14965,N_14147);
nor UO_971 (O_971,N_14567,N_14658);
or UO_972 (O_972,N_14519,N_14521);
nand UO_973 (O_973,N_14524,N_14096);
or UO_974 (O_974,N_14399,N_14691);
nand UO_975 (O_975,N_14141,N_14049);
nor UO_976 (O_976,N_14599,N_14227);
and UO_977 (O_977,N_14133,N_14193);
or UO_978 (O_978,N_14077,N_14448);
and UO_979 (O_979,N_14280,N_14471);
nand UO_980 (O_980,N_14758,N_14154);
xor UO_981 (O_981,N_14538,N_14892);
nand UO_982 (O_982,N_14630,N_14102);
and UO_983 (O_983,N_14266,N_14623);
or UO_984 (O_984,N_14494,N_14693);
nor UO_985 (O_985,N_14995,N_14541);
or UO_986 (O_986,N_14730,N_14555);
and UO_987 (O_987,N_14117,N_14299);
nor UO_988 (O_988,N_14062,N_14429);
nor UO_989 (O_989,N_14118,N_14371);
nand UO_990 (O_990,N_14950,N_14901);
nor UO_991 (O_991,N_14312,N_14170);
nand UO_992 (O_992,N_14066,N_14801);
and UO_993 (O_993,N_14109,N_14030);
nor UO_994 (O_994,N_14305,N_14259);
or UO_995 (O_995,N_14185,N_14700);
and UO_996 (O_996,N_14185,N_14097);
nand UO_997 (O_997,N_14455,N_14444);
or UO_998 (O_998,N_14366,N_14735);
and UO_999 (O_999,N_14943,N_14466);
nand UO_1000 (O_1000,N_14591,N_14718);
nor UO_1001 (O_1001,N_14544,N_14216);
nand UO_1002 (O_1002,N_14316,N_14129);
or UO_1003 (O_1003,N_14474,N_14690);
nand UO_1004 (O_1004,N_14404,N_14377);
or UO_1005 (O_1005,N_14337,N_14396);
nor UO_1006 (O_1006,N_14140,N_14799);
or UO_1007 (O_1007,N_14496,N_14134);
or UO_1008 (O_1008,N_14060,N_14339);
nand UO_1009 (O_1009,N_14058,N_14756);
nand UO_1010 (O_1010,N_14979,N_14399);
and UO_1011 (O_1011,N_14234,N_14061);
and UO_1012 (O_1012,N_14857,N_14302);
and UO_1013 (O_1013,N_14591,N_14379);
and UO_1014 (O_1014,N_14068,N_14089);
or UO_1015 (O_1015,N_14399,N_14044);
nand UO_1016 (O_1016,N_14796,N_14533);
nand UO_1017 (O_1017,N_14630,N_14022);
nor UO_1018 (O_1018,N_14898,N_14082);
xnor UO_1019 (O_1019,N_14952,N_14698);
nor UO_1020 (O_1020,N_14534,N_14795);
nand UO_1021 (O_1021,N_14602,N_14174);
nand UO_1022 (O_1022,N_14836,N_14932);
nor UO_1023 (O_1023,N_14469,N_14596);
and UO_1024 (O_1024,N_14374,N_14128);
nand UO_1025 (O_1025,N_14817,N_14302);
xnor UO_1026 (O_1026,N_14983,N_14111);
or UO_1027 (O_1027,N_14349,N_14168);
nand UO_1028 (O_1028,N_14300,N_14846);
nor UO_1029 (O_1029,N_14808,N_14566);
nor UO_1030 (O_1030,N_14811,N_14528);
xnor UO_1031 (O_1031,N_14235,N_14930);
nor UO_1032 (O_1032,N_14953,N_14608);
or UO_1033 (O_1033,N_14040,N_14599);
xnor UO_1034 (O_1034,N_14193,N_14445);
nand UO_1035 (O_1035,N_14300,N_14480);
xor UO_1036 (O_1036,N_14559,N_14648);
xnor UO_1037 (O_1037,N_14850,N_14951);
nand UO_1038 (O_1038,N_14975,N_14325);
and UO_1039 (O_1039,N_14030,N_14457);
nand UO_1040 (O_1040,N_14026,N_14317);
nand UO_1041 (O_1041,N_14047,N_14464);
or UO_1042 (O_1042,N_14078,N_14143);
xor UO_1043 (O_1043,N_14163,N_14982);
or UO_1044 (O_1044,N_14204,N_14733);
nand UO_1045 (O_1045,N_14778,N_14092);
or UO_1046 (O_1046,N_14992,N_14772);
nor UO_1047 (O_1047,N_14091,N_14733);
and UO_1048 (O_1048,N_14311,N_14871);
nand UO_1049 (O_1049,N_14404,N_14748);
or UO_1050 (O_1050,N_14469,N_14735);
nand UO_1051 (O_1051,N_14919,N_14221);
nand UO_1052 (O_1052,N_14676,N_14802);
nand UO_1053 (O_1053,N_14641,N_14820);
and UO_1054 (O_1054,N_14022,N_14032);
nor UO_1055 (O_1055,N_14473,N_14078);
nor UO_1056 (O_1056,N_14502,N_14454);
nand UO_1057 (O_1057,N_14198,N_14253);
and UO_1058 (O_1058,N_14549,N_14718);
nor UO_1059 (O_1059,N_14388,N_14566);
nor UO_1060 (O_1060,N_14749,N_14955);
xor UO_1061 (O_1061,N_14368,N_14308);
nand UO_1062 (O_1062,N_14101,N_14172);
and UO_1063 (O_1063,N_14226,N_14277);
and UO_1064 (O_1064,N_14971,N_14335);
and UO_1065 (O_1065,N_14276,N_14001);
nor UO_1066 (O_1066,N_14690,N_14563);
and UO_1067 (O_1067,N_14849,N_14528);
nor UO_1068 (O_1068,N_14707,N_14991);
and UO_1069 (O_1069,N_14106,N_14946);
nand UO_1070 (O_1070,N_14478,N_14865);
nand UO_1071 (O_1071,N_14807,N_14239);
and UO_1072 (O_1072,N_14198,N_14577);
and UO_1073 (O_1073,N_14481,N_14565);
and UO_1074 (O_1074,N_14709,N_14208);
nand UO_1075 (O_1075,N_14500,N_14035);
and UO_1076 (O_1076,N_14777,N_14727);
nor UO_1077 (O_1077,N_14614,N_14056);
nor UO_1078 (O_1078,N_14321,N_14790);
nor UO_1079 (O_1079,N_14237,N_14814);
nor UO_1080 (O_1080,N_14186,N_14143);
nand UO_1081 (O_1081,N_14517,N_14398);
nand UO_1082 (O_1082,N_14397,N_14278);
and UO_1083 (O_1083,N_14019,N_14446);
or UO_1084 (O_1084,N_14459,N_14060);
xor UO_1085 (O_1085,N_14111,N_14384);
nand UO_1086 (O_1086,N_14658,N_14806);
nand UO_1087 (O_1087,N_14802,N_14052);
and UO_1088 (O_1088,N_14180,N_14428);
or UO_1089 (O_1089,N_14963,N_14300);
xor UO_1090 (O_1090,N_14513,N_14036);
or UO_1091 (O_1091,N_14838,N_14267);
nand UO_1092 (O_1092,N_14353,N_14036);
xnor UO_1093 (O_1093,N_14634,N_14037);
nand UO_1094 (O_1094,N_14620,N_14573);
nor UO_1095 (O_1095,N_14566,N_14452);
nand UO_1096 (O_1096,N_14554,N_14015);
and UO_1097 (O_1097,N_14745,N_14583);
nor UO_1098 (O_1098,N_14641,N_14211);
and UO_1099 (O_1099,N_14172,N_14356);
nor UO_1100 (O_1100,N_14724,N_14872);
nor UO_1101 (O_1101,N_14626,N_14507);
nor UO_1102 (O_1102,N_14473,N_14701);
nor UO_1103 (O_1103,N_14326,N_14766);
or UO_1104 (O_1104,N_14807,N_14203);
or UO_1105 (O_1105,N_14278,N_14189);
or UO_1106 (O_1106,N_14449,N_14320);
nor UO_1107 (O_1107,N_14950,N_14104);
nand UO_1108 (O_1108,N_14035,N_14334);
or UO_1109 (O_1109,N_14860,N_14251);
nor UO_1110 (O_1110,N_14079,N_14099);
xnor UO_1111 (O_1111,N_14765,N_14078);
and UO_1112 (O_1112,N_14712,N_14496);
nand UO_1113 (O_1113,N_14716,N_14809);
and UO_1114 (O_1114,N_14707,N_14410);
or UO_1115 (O_1115,N_14615,N_14129);
and UO_1116 (O_1116,N_14705,N_14768);
and UO_1117 (O_1117,N_14933,N_14702);
nor UO_1118 (O_1118,N_14365,N_14459);
xor UO_1119 (O_1119,N_14109,N_14520);
or UO_1120 (O_1120,N_14736,N_14891);
or UO_1121 (O_1121,N_14676,N_14950);
or UO_1122 (O_1122,N_14896,N_14354);
and UO_1123 (O_1123,N_14784,N_14810);
and UO_1124 (O_1124,N_14666,N_14936);
and UO_1125 (O_1125,N_14956,N_14930);
or UO_1126 (O_1126,N_14832,N_14174);
nor UO_1127 (O_1127,N_14262,N_14645);
nand UO_1128 (O_1128,N_14249,N_14170);
nor UO_1129 (O_1129,N_14770,N_14778);
nor UO_1130 (O_1130,N_14324,N_14179);
and UO_1131 (O_1131,N_14329,N_14421);
and UO_1132 (O_1132,N_14313,N_14808);
or UO_1133 (O_1133,N_14974,N_14342);
nand UO_1134 (O_1134,N_14755,N_14831);
or UO_1135 (O_1135,N_14973,N_14506);
nor UO_1136 (O_1136,N_14732,N_14950);
nor UO_1137 (O_1137,N_14806,N_14561);
nor UO_1138 (O_1138,N_14332,N_14912);
nor UO_1139 (O_1139,N_14028,N_14693);
nand UO_1140 (O_1140,N_14218,N_14687);
or UO_1141 (O_1141,N_14600,N_14353);
nand UO_1142 (O_1142,N_14470,N_14103);
nand UO_1143 (O_1143,N_14302,N_14917);
xor UO_1144 (O_1144,N_14609,N_14457);
nand UO_1145 (O_1145,N_14472,N_14384);
or UO_1146 (O_1146,N_14168,N_14741);
nor UO_1147 (O_1147,N_14479,N_14169);
nor UO_1148 (O_1148,N_14561,N_14623);
and UO_1149 (O_1149,N_14676,N_14224);
or UO_1150 (O_1150,N_14801,N_14569);
xnor UO_1151 (O_1151,N_14695,N_14875);
or UO_1152 (O_1152,N_14849,N_14026);
and UO_1153 (O_1153,N_14566,N_14007);
nor UO_1154 (O_1154,N_14387,N_14976);
nor UO_1155 (O_1155,N_14174,N_14667);
xnor UO_1156 (O_1156,N_14130,N_14458);
nand UO_1157 (O_1157,N_14247,N_14925);
and UO_1158 (O_1158,N_14586,N_14688);
nand UO_1159 (O_1159,N_14880,N_14716);
and UO_1160 (O_1160,N_14853,N_14728);
nor UO_1161 (O_1161,N_14049,N_14586);
or UO_1162 (O_1162,N_14027,N_14208);
and UO_1163 (O_1163,N_14803,N_14943);
or UO_1164 (O_1164,N_14436,N_14274);
nor UO_1165 (O_1165,N_14253,N_14392);
or UO_1166 (O_1166,N_14662,N_14088);
nand UO_1167 (O_1167,N_14987,N_14752);
nand UO_1168 (O_1168,N_14075,N_14602);
nand UO_1169 (O_1169,N_14792,N_14254);
nand UO_1170 (O_1170,N_14066,N_14468);
xor UO_1171 (O_1171,N_14587,N_14677);
xnor UO_1172 (O_1172,N_14580,N_14397);
nor UO_1173 (O_1173,N_14307,N_14920);
nor UO_1174 (O_1174,N_14769,N_14684);
nand UO_1175 (O_1175,N_14010,N_14673);
nand UO_1176 (O_1176,N_14857,N_14320);
or UO_1177 (O_1177,N_14520,N_14698);
and UO_1178 (O_1178,N_14565,N_14222);
nor UO_1179 (O_1179,N_14355,N_14984);
nand UO_1180 (O_1180,N_14814,N_14895);
or UO_1181 (O_1181,N_14588,N_14598);
nand UO_1182 (O_1182,N_14498,N_14857);
or UO_1183 (O_1183,N_14146,N_14634);
nand UO_1184 (O_1184,N_14410,N_14715);
and UO_1185 (O_1185,N_14922,N_14247);
nand UO_1186 (O_1186,N_14754,N_14451);
or UO_1187 (O_1187,N_14250,N_14749);
nor UO_1188 (O_1188,N_14368,N_14431);
nand UO_1189 (O_1189,N_14441,N_14982);
or UO_1190 (O_1190,N_14947,N_14037);
nand UO_1191 (O_1191,N_14856,N_14656);
nand UO_1192 (O_1192,N_14308,N_14161);
or UO_1193 (O_1193,N_14613,N_14705);
nor UO_1194 (O_1194,N_14869,N_14446);
xor UO_1195 (O_1195,N_14985,N_14652);
nor UO_1196 (O_1196,N_14558,N_14706);
or UO_1197 (O_1197,N_14884,N_14482);
or UO_1198 (O_1198,N_14529,N_14964);
xnor UO_1199 (O_1199,N_14688,N_14945);
or UO_1200 (O_1200,N_14641,N_14141);
xnor UO_1201 (O_1201,N_14956,N_14965);
and UO_1202 (O_1202,N_14766,N_14224);
nand UO_1203 (O_1203,N_14732,N_14835);
and UO_1204 (O_1204,N_14580,N_14347);
nor UO_1205 (O_1205,N_14670,N_14373);
nand UO_1206 (O_1206,N_14748,N_14266);
and UO_1207 (O_1207,N_14370,N_14357);
and UO_1208 (O_1208,N_14688,N_14433);
xnor UO_1209 (O_1209,N_14509,N_14655);
nand UO_1210 (O_1210,N_14890,N_14568);
nor UO_1211 (O_1211,N_14076,N_14657);
nor UO_1212 (O_1212,N_14334,N_14770);
nand UO_1213 (O_1213,N_14609,N_14069);
or UO_1214 (O_1214,N_14674,N_14971);
nor UO_1215 (O_1215,N_14208,N_14016);
nand UO_1216 (O_1216,N_14712,N_14529);
or UO_1217 (O_1217,N_14244,N_14048);
nor UO_1218 (O_1218,N_14822,N_14311);
or UO_1219 (O_1219,N_14623,N_14843);
and UO_1220 (O_1220,N_14414,N_14887);
nand UO_1221 (O_1221,N_14808,N_14030);
nand UO_1222 (O_1222,N_14266,N_14364);
xnor UO_1223 (O_1223,N_14675,N_14002);
and UO_1224 (O_1224,N_14414,N_14137);
or UO_1225 (O_1225,N_14781,N_14686);
and UO_1226 (O_1226,N_14770,N_14316);
and UO_1227 (O_1227,N_14968,N_14181);
nor UO_1228 (O_1228,N_14552,N_14089);
xnor UO_1229 (O_1229,N_14406,N_14183);
or UO_1230 (O_1230,N_14994,N_14939);
and UO_1231 (O_1231,N_14208,N_14991);
nor UO_1232 (O_1232,N_14506,N_14488);
nand UO_1233 (O_1233,N_14047,N_14482);
xnor UO_1234 (O_1234,N_14293,N_14250);
nor UO_1235 (O_1235,N_14599,N_14044);
and UO_1236 (O_1236,N_14361,N_14826);
and UO_1237 (O_1237,N_14760,N_14293);
nand UO_1238 (O_1238,N_14354,N_14164);
nand UO_1239 (O_1239,N_14542,N_14508);
or UO_1240 (O_1240,N_14297,N_14093);
xnor UO_1241 (O_1241,N_14659,N_14592);
xor UO_1242 (O_1242,N_14411,N_14260);
or UO_1243 (O_1243,N_14650,N_14742);
nand UO_1244 (O_1244,N_14900,N_14078);
or UO_1245 (O_1245,N_14858,N_14955);
and UO_1246 (O_1246,N_14772,N_14375);
nor UO_1247 (O_1247,N_14175,N_14306);
and UO_1248 (O_1248,N_14995,N_14345);
or UO_1249 (O_1249,N_14295,N_14683);
nand UO_1250 (O_1250,N_14098,N_14770);
nor UO_1251 (O_1251,N_14876,N_14094);
and UO_1252 (O_1252,N_14687,N_14455);
and UO_1253 (O_1253,N_14693,N_14308);
nor UO_1254 (O_1254,N_14828,N_14835);
and UO_1255 (O_1255,N_14351,N_14432);
nand UO_1256 (O_1256,N_14848,N_14492);
and UO_1257 (O_1257,N_14770,N_14982);
nor UO_1258 (O_1258,N_14564,N_14370);
or UO_1259 (O_1259,N_14735,N_14674);
nor UO_1260 (O_1260,N_14303,N_14150);
and UO_1261 (O_1261,N_14652,N_14647);
xor UO_1262 (O_1262,N_14733,N_14130);
and UO_1263 (O_1263,N_14383,N_14712);
nand UO_1264 (O_1264,N_14019,N_14644);
and UO_1265 (O_1265,N_14685,N_14719);
nor UO_1266 (O_1266,N_14178,N_14825);
nand UO_1267 (O_1267,N_14198,N_14686);
nor UO_1268 (O_1268,N_14767,N_14827);
and UO_1269 (O_1269,N_14506,N_14589);
and UO_1270 (O_1270,N_14875,N_14906);
and UO_1271 (O_1271,N_14138,N_14620);
nor UO_1272 (O_1272,N_14484,N_14784);
or UO_1273 (O_1273,N_14220,N_14041);
and UO_1274 (O_1274,N_14208,N_14053);
and UO_1275 (O_1275,N_14196,N_14240);
nor UO_1276 (O_1276,N_14580,N_14162);
or UO_1277 (O_1277,N_14238,N_14426);
nor UO_1278 (O_1278,N_14801,N_14947);
and UO_1279 (O_1279,N_14614,N_14446);
nand UO_1280 (O_1280,N_14455,N_14778);
nand UO_1281 (O_1281,N_14376,N_14576);
nand UO_1282 (O_1282,N_14365,N_14444);
nor UO_1283 (O_1283,N_14655,N_14244);
nand UO_1284 (O_1284,N_14206,N_14426);
and UO_1285 (O_1285,N_14389,N_14231);
nor UO_1286 (O_1286,N_14400,N_14416);
nor UO_1287 (O_1287,N_14559,N_14967);
or UO_1288 (O_1288,N_14682,N_14491);
or UO_1289 (O_1289,N_14254,N_14771);
nand UO_1290 (O_1290,N_14457,N_14079);
nand UO_1291 (O_1291,N_14334,N_14730);
nand UO_1292 (O_1292,N_14401,N_14437);
nor UO_1293 (O_1293,N_14574,N_14321);
and UO_1294 (O_1294,N_14845,N_14858);
xnor UO_1295 (O_1295,N_14466,N_14864);
xnor UO_1296 (O_1296,N_14534,N_14407);
or UO_1297 (O_1297,N_14591,N_14867);
and UO_1298 (O_1298,N_14234,N_14999);
nand UO_1299 (O_1299,N_14594,N_14648);
and UO_1300 (O_1300,N_14277,N_14930);
and UO_1301 (O_1301,N_14134,N_14221);
or UO_1302 (O_1302,N_14357,N_14909);
and UO_1303 (O_1303,N_14099,N_14758);
or UO_1304 (O_1304,N_14906,N_14919);
or UO_1305 (O_1305,N_14024,N_14920);
and UO_1306 (O_1306,N_14848,N_14085);
xor UO_1307 (O_1307,N_14780,N_14775);
xor UO_1308 (O_1308,N_14205,N_14954);
nand UO_1309 (O_1309,N_14291,N_14388);
or UO_1310 (O_1310,N_14352,N_14395);
and UO_1311 (O_1311,N_14779,N_14542);
nor UO_1312 (O_1312,N_14178,N_14526);
or UO_1313 (O_1313,N_14562,N_14977);
xor UO_1314 (O_1314,N_14809,N_14738);
nor UO_1315 (O_1315,N_14980,N_14799);
or UO_1316 (O_1316,N_14549,N_14565);
and UO_1317 (O_1317,N_14506,N_14676);
nor UO_1318 (O_1318,N_14855,N_14628);
or UO_1319 (O_1319,N_14086,N_14973);
nand UO_1320 (O_1320,N_14265,N_14808);
and UO_1321 (O_1321,N_14989,N_14227);
and UO_1322 (O_1322,N_14218,N_14339);
and UO_1323 (O_1323,N_14385,N_14553);
xor UO_1324 (O_1324,N_14562,N_14882);
or UO_1325 (O_1325,N_14590,N_14832);
or UO_1326 (O_1326,N_14951,N_14276);
nor UO_1327 (O_1327,N_14100,N_14495);
nand UO_1328 (O_1328,N_14704,N_14932);
or UO_1329 (O_1329,N_14879,N_14442);
nor UO_1330 (O_1330,N_14723,N_14298);
nor UO_1331 (O_1331,N_14253,N_14638);
nor UO_1332 (O_1332,N_14948,N_14858);
or UO_1333 (O_1333,N_14638,N_14622);
or UO_1334 (O_1334,N_14097,N_14258);
or UO_1335 (O_1335,N_14767,N_14077);
nor UO_1336 (O_1336,N_14766,N_14064);
nand UO_1337 (O_1337,N_14230,N_14369);
and UO_1338 (O_1338,N_14270,N_14325);
or UO_1339 (O_1339,N_14111,N_14578);
and UO_1340 (O_1340,N_14734,N_14654);
or UO_1341 (O_1341,N_14013,N_14746);
nor UO_1342 (O_1342,N_14140,N_14648);
nand UO_1343 (O_1343,N_14882,N_14845);
or UO_1344 (O_1344,N_14671,N_14818);
nor UO_1345 (O_1345,N_14826,N_14174);
or UO_1346 (O_1346,N_14955,N_14286);
nor UO_1347 (O_1347,N_14120,N_14119);
and UO_1348 (O_1348,N_14852,N_14950);
nand UO_1349 (O_1349,N_14052,N_14786);
or UO_1350 (O_1350,N_14507,N_14317);
or UO_1351 (O_1351,N_14691,N_14532);
and UO_1352 (O_1352,N_14415,N_14595);
or UO_1353 (O_1353,N_14109,N_14969);
nor UO_1354 (O_1354,N_14995,N_14160);
xnor UO_1355 (O_1355,N_14762,N_14790);
nor UO_1356 (O_1356,N_14368,N_14115);
nor UO_1357 (O_1357,N_14435,N_14073);
xor UO_1358 (O_1358,N_14539,N_14102);
nand UO_1359 (O_1359,N_14073,N_14674);
and UO_1360 (O_1360,N_14669,N_14568);
or UO_1361 (O_1361,N_14909,N_14292);
or UO_1362 (O_1362,N_14451,N_14538);
nand UO_1363 (O_1363,N_14231,N_14705);
and UO_1364 (O_1364,N_14935,N_14761);
nor UO_1365 (O_1365,N_14510,N_14019);
and UO_1366 (O_1366,N_14570,N_14993);
and UO_1367 (O_1367,N_14249,N_14882);
nand UO_1368 (O_1368,N_14965,N_14693);
or UO_1369 (O_1369,N_14098,N_14663);
or UO_1370 (O_1370,N_14928,N_14066);
and UO_1371 (O_1371,N_14631,N_14019);
xor UO_1372 (O_1372,N_14444,N_14845);
nand UO_1373 (O_1373,N_14026,N_14214);
and UO_1374 (O_1374,N_14929,N_14984);
nand UO_1375 (O_1375,N_14228,N_14748);
and UO_1376 (O_1376,N_14656,N_14298);
or UO_1377 (O_1377,N_14018,N_14256);
or UO_1378 (O_1378,N_14200,N_14832);
or UO_1379 (O_1379,N_14746,N_14441);
xor UO_1380 (O_1380,N_14714,N_14510);
nor UO_1381 (O_1381,N_14598,N_14238);
nor UO_1382 (O_1382,N_14945,N_14980);
nand UO_1383 (O_1383,N_14319,N_14478);
and UO_1384 (O_1384,N_14377,N_14250);
or UO_1385 (O_1385,N_14565,N_14037);
xor UO_1386 (O_1386,N_14588,N_14846);
nor UO_1387 (O_1387,N_14481,N_14310);
nand UO_1388 (O_1388,N_14767,N_14247);
nand UO_1389 (O_1389,N_14113,N_14908);
nand UO_1390 (O_1390,N_14962,N_14238);
nor UO_1391 (O_1391,N_14057,N_14503);
and UO_1392 (O_1392,N_14510,N_14067);
nand UO_1393 (O_1393,N_14845,N_14048);
xor UO_1394 (O_1394,N_14341,N_14829);
nand UO_1395 (O_1395,N_14770,N_14270);
nand UO_1396 (O_1396,N_14549,N_14339);
nor UO_1397 (O_1397,N_14029,N_14173);
nor UO_1398 (O_1398,N_14922,N_14777);
or UO_1399 (O_1399,N_14817,N_14916);
nand UO_1400 (O_1400,N_14214,N_14848);
nand UO_1401 (O_1401,N_14540,N_14876);
xor UO_1402 (O_1402,N_14369,N_14899);
and UO_1403 (O_1403,N_14982,N_14587);
nand UO_1404 (O_1404,N_14470,N_14809);
nand UO_1405 (O_1405,N_14226,N_14527);
and UO_1406 (O_1406,N_14534,N_14857);
or UO_1407 (O_1407,N_14140,N_14144);
nor UO_1408 (O_1408,N_14092,N_14723);
or UO_1409 (O_1409,N_14374,N_14651);
and UO_1410 (O_1410,N_14659,N_14536);
nor UO_1411 (O_1411,N_14910,N_14324);
and UO_1412 (O_1412,N_14221,N_14748);
or UO_1413 (O_1413,N_14053,N_14172);
and UO_1414 (O_1414,N_14862,N_14211);
or UO_1415 (O_1415,N_14377,N_14986);
and UO_1416 (O_1416,N_14811,N_14149);
nor UO_1417 (O_1417,N_14629,N_14207);
nand UO_1418 (O_1418,N_14270,N_14792);
nor UO_1419 (O_1419,N_14224,N_14755);
or UO_1420 (O_1420,N_14979,N_14420);
and UO_1421 (O_1421,N_14849,N_14647);
nand UO_1422 (O_1422,N_14814,N_14025);
and UO_1423 (O_1423,N_14933,N_14973);
nand UO_1424 (O_1424,N_14307,N_14459);
or UO_1425 (O_1425,N_14947,N_14067);
and UO_1426 (O_1426,N_14054,N_14529);
nor UO_1427 (O_1427,N_14446,N_14259);
xor UO_1428 (O_1428,N_14101,N_14189);
nand UO_1429 (O_1429,N_14098,N_14812);
and UO_1430 (O_1430,N_14702,N_14780);
xnor UO_1431 (O_1431,N_14383,N_14366);
and UO_1432 (O_1432,N_14411,N_14483);
nor UO_1433 (O_1433,N_14330,N_14506);
nand UO_1434 (O_1434,N_14737,N_14414);
nand UO_1435 (O_1435,N_14366,N_14707);
or UO_1436 (O_1436,N_14210,N_14647);
and UO_1437 (O_1437,N_14751,N_14763);
or UO_1438 (O_1438,N_14821,N_14756);
xor UO_1439 (O_1439,N_14854,N_14977);
or UO_1440 (O_1440,N_14234,N_14572);
nand UO_1441 (O_1441,N_14966,N_14147);
nor UO_1442 (O_1442,N_14282,N_14342);
nor UO_1443 (O_1443,N_14084,N_14615);
or UO_1444 (O_1444,N_14904,N_14011);
nand UO_1445 (O_1445,N_14030,N_14226);
or UO_1446 (O_1446,N_14103,N_14624);
or UO_1447 (O_1447,N_14572,N_14035);
nand UO_1448 (O_1448,N_14577,N_14541);
xor UO_1449 (O_1449,N_14838,N_14732);
xnor UO_1450 (O_1450,N_14141,N_14455);
or UO_1451 (O_1451,N_14221,N_14304);
and UO_1452 (O_1452,N_14728,N_14635);
and UO_1453 (O_1453,N_14084,N_14078);
nand UO_1454 (O_1454,N_14167,N_14986);
xnor UO_1455 (O_1455,N_14476,N_14638);
and UO_1456 (O_1456,N_14748,N_14539);
nor UO_1457 (O_1457,N_14273,N_14898);
or UO_1458 (O_1458,N_14086,N_14525);
and UO_1459 (O_1459,N_14417,N_14725);
nor UO_1460 (O_1460,N_14049,N_14286);
xor UO_1461 (O_1461,N_14936,N_14226);
nand UO_1462 (O_1462,N_14119,N_14215);
nand UO_1463 (O_1463,N_14794,N_14745);
xor UO_1464 (O_1464,N_14782,N_14606);
or UO_1465 (O_1465,N_14048,N_14499);
or UO_1466 (O_1466,N_14248,N_14380);
nor UO_1467 (O_1467,N_14116,N_14485);
or UO_1468 (O_1468,N_14528,N_14765);
or UO_1469 (O_1469,N_14912,N_14354);
nand UO_1470 (O_1470,N_14870,N_14953);
and UO_1471 (O_1471,N_14856,N_14017);
and UO_1472 (O_1472,N_14195,N_14001);
and UO_1473 (O_1473,N_14080,N_14667);
nor UO_1474 (O_1474,N_14463,N_14335);
nor UO_1475 (O_1475,N_14519,N_14483);
nand UO_1476 (O_1476,N_14433,N_14997);
xnor UO_1477 (O_1477,N_14489,N_14895);
and UO_1478 (O_1478,N_14568,N_14595);
xnor UO_1479 (O_1479,N_14260,N_14207);
and UO_1480 (O_1480,N_14489,N_14613);
nor UO_1481 (O_1481,N_14700,N_14045);
xor UO_1482 (O_1482,N_14046,N_14396);
or UO_1483 (O_1483,N_14094,N_14080);
nor UO_1484 (O_1484,N_14246,N_14339);
nand UO_1485 (O_1485,N_14055,N_14309);
nand UO_1486 (O_1486,N_14089,N_14235);
and UO_1487 (O_1487,N_14480,N_14997);
or UO_1488 (O_1488,N_14063,N_14064);
and UO_1489 (O_1489,N_14735,N_14889);
xnor UO_1490 (O_1490,N_14783,N_14171);
and UO_1491 (O_1491,N_14762,N_14173);
nand UO_1492 (O_1492,N_14867,N_14678);
nor UO_1493 (O_1493,N_14672,N_14622);
or UO_1494 (O_1494,N_14104,N_14120);
nand UO_1495 (O_1495,N_14128,N_14404);
and UO_1496 (O_1496,N_14492,N_14055);
nor UO_1497 (O_1497,N_14307,N_14870);
xnor UO_1498 (O_1498,N_14475,N_14565);
and UO_1499 (O_1499,N_14921,N_14833);
and UO_1500 (O_1500,N_14781,N_14488);
nor UO_1501 (O_1501,N_14501,N_14101);
nor UO_1502 (O_1502,N_14454,N_14752);
nor UO_1503 (O_1503,N_14015,N_14076);
xnor UO_1504 (O_1504,N_14677,N_14213);
or UO_1505 (O_1505,N_14406,N_14122);
nor UO_1506 (O_1506,N_14103,N_14059);
nor UO_1507 (O_1507,N_14649,N_14893);
nand UO_1508 (O_1508,N_14059,N_14375);
nor UO_1509 (O_1509,N_14508,N_14178);
nand UO_1510 (O_1510,N_14035,N_14382);
and UO_1511 (O_1511,N_14565,N_14911);
nand UO_1512 (O_1512,N_14838,N_14161);
nand UO_1513 (O_1513,N_14949,N_14234);
and UO_1514 (O_1514,N_14792,N_14358);
and UO_1515 (O_1515,N_14989,N_14022);
nor UO_1516 (O_1516,N_14665,N_14674);
nor UO_1517 (O_1517,N_14144,N_14865);
and UO_1518 (O_1518,N_14029,N_14628);
nor UO_1519 (O_1519,N_14699,N_14176);
or UO_1520 (O_1520,N_14206,N_14222);
and UO_1521 (O_1521,N_14016,N_14458);
nand UO_1522 (O_1522,N_14652,N_14077);
and UO_1523 (O_1523,N_14949,N_14792);
nor UO_1524 (O_1524,N_14559,N_14963);
or UO_1525 (O_1525,N_14747,N_14709);
nor UO_1526 (O_1526,N_14916,N_14060);
or UO_1527 (O_1527,N_14657,N_14138);
or UO_1528 (O_1528,N_14442,N_14983);
nand UO_1529 (O_1529,N_14710,N_14854);
and UO_1530 (O_1530,N_14812,N_14722);
or UO_1531 (O_1531,N_14570,N_14433);
nand UO_1532 (O_1532,N_14672,N_14615);
nand UO_1533 (O_1533,N_14937,N_14545);
nor UO_1534 (O_1534,N_14734,N_14561);
or UO_1535 (O_1535,N_14544,N_14908);
or UO_1536 (O_1536,N_14392,N_14050);
nor UO_1537 (O_1537,N_14895,N_14407);
nand UO_1538 (O_1538,N_14052,N_14625);
nand UO_1539 (O_1539,N_14636,N_14541);
nor UO_1540 (O_1540,N_14988,N_14590);
or UO_1541 (O_1541,N_14886,N_14697);
xor UO_1542 (O_1542,N_14171,N_14169);
xnor UO_1543 (O_1543,N_14594,N_14695);
or UO_1544 (O_1544,N_14051,N_14948);
nand UO_1545 (O_1545,N_14603,N_14974);
or UO_1546 (O_1546,N_14441,N_14260);
nor UO_1547 (O_1547,N_14095,N_14354);
or UO_1548 (O_1548,N_14015,N_14483);
or UO_1549 (O_1549,N_14502,N_14597);
nand UO_1550 (O_1550,N_14132,N_14283);
and UO_1551 (O_1551,N_14185,N_14312);
xor UO_1552 (O_1552,N_14032,N_14761);
xnor UO_1553 (O_1553,N_14194,N_14063);
and UO_1554 (O_1554,N_14532,N_14177);
xor UO_1555 (O_1555,N_14758,N_14299);
nor UO_1556 (O_1556,N_14653,N_14313);
or UO_1557 (O_1557,N_14093,N_14207);
xor UO_1558 (O_1558,N_14978,N_14737);
and UO_1559 (O_1559,N_14330,N_14301);
and UO_1560 (O_1560,N_14552,N_14709);
nand UO_1561 (O_1561,N_14288,N_14342);
nand UO_1562 (O_1562,N_14511,N_14757);
or UO_1563 (O_1563,N_14581,N_14994);
and UO_1564 (O_1564,N_14527,N_14474);
nand UO_1565 (O_1565,N_14589,N_14127);
nor UO_1566 (O_1566,N_14139,N_14044);
nand UO_1567 (O_1567,N_14507,N_14791);
or UO_1568 (O_1568,N_14087,N_14733);
and UO_1569 (O_1569,N_14317,N_14103);
or UO_1570 (O_1570,N_14748,N_14254);
nor UO_1571 (O_1571,N_14532,N_14892);
nand UO_1572 (O_1572,N_14173,N_14880);
nor UO_1573 (O_1573,N_14108,N_14069);
or UO_1574 (O_1574,N_14984,N_14386);
and UO_1575 (O_1575,N_14017,N_14382);
xor UO_1576 (O_1576,N_14523,N_14024);
or UO_1577 (O_1577,N_14389,N_14938);
or UO_1578 (O_1578,N_14098,N_14425);
or UO_1579 (O_1579,N_14974,N_14254);
or UO_1580 (O_1580,N_14810,N_14756);
xnor UO_1581 (O_1581,N_14371,N_14488);
or UO_1582 (O_1582,N_14516,N_14253);
nor UO_1583 (O_1583,N_14626,N_14328);
or UO_1584 (O_1584,N_14966,N_14101);
nor UO_1585 (O_1585,N_14388,N_14620);
or UO_1586 (O_1586,N_14482,N_14447);
nor UO_1587 (O_1587,N_14854,N_14457);
and UO_1588 (O_1588,N_14352,N_14164);
nand UO_1589 (O_1589,N_14335,N_14837);
nand UO_1590 (O_1590,N_14716,N_14285);
nor UO_1591 (O_1591,N_14847,N_14693);
nand UO_1592 (O_1592,N_14540,N_14418);
and UO_1593 (O_1593,N_14032,N_14682);
nand UO_1594 (O_1594,N_14791,N_14844);
nor UO_1595 (O_1595,N_14557,N_14276);
or UO_1596 (O_1596,N_14584,N_14515);
nand UO_1597 (O_1597,N_14989,N_14763);
nor UO_1598 (O_1598,N_14581,N_14991);
nor UO_1599 (O_1599,N_14099,N_14017);
nand UO_1600 (O_1600,N_14185,N_14972);
nor UO_1601 (O_1601,N_14973,N_14799);
or UO_1602 (O_1602,N_14202,N_14241);
or UO_1603 (O_1603,N_14116,N_14095);
or UO_1604 (O_1604,N_14886,N_14138);
nand UO_1605 (O_1605,N_14871,N_14113);
nor UO_1606 (O_1606,N_14016,N_14738);
nand UO_1607 (O_1607,N_14500,N_14875);
nand UO_1608 (O_1608,N_14331,N_14375);
and UO_1609 (O_1609,N_14616,N_14398);
and UO_1610 (O_1610,N_14273,N_14818);
nor UO_1611 (O_1611,N_14536,N_14746);
or UO_1612 (O_1612,N_14183,N_14148);
nor UO_1613 (O_1613,N_14525,N_14387);
xor UO_1614 (O_1614,N_14687,N_14810);
nand UO_1615 (O_1615,N_14662,N_14485);
or UO_1616 (O_1616,N_14557,N_14213);
or UO_1617 (O_1617,N_14271,N_14772);
xor UO_1618 (O_1618,N_14506,N_14982);
nand UO_1619 (O_1619,N_14149,N_14039);
nor UO_1620 (O_1620,N_14744,N_14509);
nand UO_1621 (O_1621,N_14931,N_14231);
nand UO_1622 (O_1622,N_14049,N_14926);
nand UO_1623 (O_1623,N_14505,N_14420);
and UO_1624 (O_1624,N_14809,N_14923);
xor UO_1625 (O_1625,N_14280,N_14001);
or UO_1626 (O_1626,N_14727,N_14138);
xor UO_1627 (O_1627,N_14053,N_14244);
nor UO_1628 (O_1628,N_14137,N_14479);
or UO_1629 (O_1629,N_14594,N_14712);
and UO_1630 (O_1630,N_14020,N_14546);
or UO_1631 (O_1631,N_14982,N_14205);
and UO_1632 (O_1632,N_14985,N_14961);
and UO_1633 (O_1633,N_14648,N_14986);
and UO_1634 (O_1634,N_14392,N_14701);
and UO_1635 (O_1635,N_14207,N_14691);
or UO_1636 (O_1636,N_14257,N_14896);
nor UO_1637 (O_1637,N_14635,N_14322);
or UO_1638 (O_1638,N_14034,N_14206);
or UO_1639 (O_1639,N_14225,N_14139);
or UO_1640 (O_1640,N_14996,N_14157);
and UO_1641 (O_1641,N_14229,N_14903);
and UO_1642 (O_1642,N_14801,N_14351);
and UO_1643 (O_1643,N_14098,N_14349);
nor UO_1644 (O_1644,N_14258,N_14641);
and UO_1645 (O_1645,N_14516,N_14098);
nand UO_1646 (O_1646,N_14301,N_14267);
nand UO_1647 (O_1647,N_14200,N_14932);
and UO_1648 (O_1648,N_14917,N_14920);
or UO_1649 (O_1649,N_14755,N_14291);
nor UO_1650 (O_1650,N_14822,N_14688);
nand UO_1651 (O_1651,N_14767,N_14068);
and UO_1652 (O_1652,N_14397,N_14069);
or UO_1653 (O_1653,N_14485,N_14435);
nand UO_1654 (O_1654,N_14437,N_14218);
or UO_1655 (O_1655,N_14297,N_14167);
or UO_1656 (O_1656,N_14213,N_14446);
nand UO_1657 (O_1657,N_14129,N_14772);
and UO_1658 (O_1658,N_14680,N_14499);
xor UO_1659 (O_1659,N_14408,N_14887);
and UO_1660 (O_1660,N_14649,N_14708);
and UO_1661 (O_1661,N_14921,N_14918);
nor UO_1662 (O_1662,N_14964,N_14064);
and UO_1663 (O_1663,N_14986,N_14348);
nand UO_1664 (O_1664,N_14682,N_14430);
or UO_1665 (O_1665,N_14879,N_14699);
xnor UO_1666 (O_1666,N_14806,N_14380);
nand UO_1667 (O_1667,N_14966,N_14544);
nor UO_1668 (O_1668,N_14521,N_14135);
and UO_1669 (O_1669,N_14313,N_14826);
and UO_1670 (O_1670,N_14885,N_14148);
nor UO_1671 (O_1671,N_14487,N_14972);
nand UO_1672 (O_1672,N_14914,N_14219);
or UO_1673 (O_1673,N_14614,N_14766);
nand UO_1674 (O_1674,N_14237,N_14793);
or UO_1675 (O_1675,N_14150,N_14513);
nand UO_1676 (O_1676,N_14321,N_14814);
xor UO_1677 (O_1677,N_14515,N_14071);
or UO_1678 (O_1678,N_14702,N_14973);
nand UO_1679 (O_1679,N_14481,N_14473);
nand UO_1680 (O_1680,N_14899,N_14946);
and UO_1681 (O_1681,N_14452,N_14834);
nand UO_1682 (O_1682,N_14990,N_14683);
nor UO_1683 (O_1683,N_14127,N_14096);
or UO_1684 (O_1684,N_14785,N_14473);
and UO_1685 (O_1685,N_14975,N_14473);
nand UO_1686 (O_1686,N_14635,N_14392);
and UO_1687 (O_1687,N_14965,N_14605);
nor UO_1688 (O_1688,N_14966,N_14371);
xor UO_1689 (O_1689,N_14013,N_14169);
and UO_1690 (O_1690,N_14737,N_14899);
or UO_1691 (O_1691,N_14920,N_14419);
xnor UO_1692 (O_1692,N_14068,N_14332);
xnor UO_1693 (O_1693,N_14036,N_14313);
nor UO_1694 (O_1694,N_14741,N_14653);
or UO_1695 (O_1695,N_14567,N_14472);
nor UO_1696 (O_1696,N_14999,N_14396);
or UO_1697 (O_1697,N_14829,N_14490);
and UO_1698 (O_1698,N_14561,N_14299);
nand UO_1699 (O_1699,N_14338,N_14268);
nor UO_1700 (O_1700,N_14337,N_14273);
and UO_1701 (O_1701,N_14006,N_14818);
and UO_1702 (O_1702,N_14929,N_14512);
nand UO_1703 (O_1703,N_14736,N_14940);
and UO_1704 (O_1704,N_14440,N_14416);
xor UO_1705 (O_1705,N_14818,N_14587);
nand UO_1706 (O_1706,N_14251,N_14881);
nand UO_1707 (O_1707,N_14938,N_14479);
nor UO_1708 (O_1708,N_14001,N_14851);
and UO_1709 (O_1709,N_14825,N_14056);
nor UO_1710 (O_1710,N_14404,N_14747);
and UO_1711 (O_1711,N_14218,N_14330);
nand UO_1712 (O_1712,N_14212,N_14720);
nor UO_1713 (O_1713,N_14145,N_14535);
nand UO_1714 (O_1714,N_14931,N_14758);
or UO_1715 (O_1715,N_14613,N_14988);
nor UO_1716 (O_1716,N_14771,N_14426);
and UO_1717 (O_1717,N_14024,N_14787);
nand UO_1718 (O_1718,N_14011,N_14772);
or UO_1719 (O_1719,N_14445,N_14442);
nand UO_1720 (O_1720,N_14836,N_14517);
nand UO_1721 (O_1721,N_14531,N_14636);
or UO_1722 (O_1722,N_14207,N_14317);
nand UO_1723 (O_1723,N_14789,N_14889);
nand UO_1724 (O_1724,N_14679,N_14722);
or UO_1725 (O_1725,N_14139,N_14748);
nor UO_1726 (O_1726,N_14017,N_14585);
and UO_1727 (O_1727,N_14571,N_14259);
or UO_1728 (O_1728,N_14285,N_14028);
or UO_1729 (O_1729,N_14157,N_14643);
nand UO_1730 (O_1730,N_14219,N_14407);
xnor UO_1731 (O_1731,N_14157,N_14380);
nor UO_1732 (O_1732,N_14718,N_14165);
nand UO_1733 (O_1733,N_14060,N_14875);
nor UO_1734 (O_1734,N_14619,N_14169);
and UO_1735 (O_1735,N_14494,N_14698);
xor UO_1736 (O_1736,N_14476,N_14119);
and UO_1737 (O_1737,N_14603,N_14329);
and UO_1738 (O_1738,N_14531,N_14395);
or UO_1739 (O_1739,N_14024,N_14271);
and UO_1740 (O_1740,N_14302,N_14376);
nor UO_1741 (O_1741,N_14309,N_14773);
nand UO_1742 (O_1742,N_14764,N_14385);
nor UO_1743 (O_1743,N_14645,N_14814);
nand UO_1744 (O_1744,N_14197,N_14371);
and UO_1745 (O_1745,N_14086,N_14392);
nor UO_1746 (O_1746,N_14674,N_14731);
nand UO_1747 (O_1747,N_14529,N_14617);
or UO_1748 (O_1748,N_14686,N_14758);
nand UO_1749 (O_1749,N_14247,N_14465);
and UO_1750 (O_1750,N_14223,N_14911);
or UO_1751 (O_1751,N_14821,N_14509);
nand UO_1752 (O_1752,N_14830,N_14050);
and UO_1753 (O_1753,N_14444,N_14165);
and UO_1754 (O_1754,N_14240,N_14158);
or UO_1755 (O_1755,N_14883,N_14517);
xor UO_1756 (O_1756,N_14074,N_14102);
nand UO_1757 (O_1757,N_14609,N_14567);
nand UO_1758 (O_1758,N_14579,N_14074);
and UO_1759 (O_1759,N_14522,N_14799);
and UO_1760 (O_1760,N_14237,N_14614);
nor UO_1761 (O_1761,N_14213,N_14425);
nand UO_1762 (O_1762,N_14787,N_14259);
xor UO_1763 (O_1763,N_14388,N_14837);
and UO_1764 (O_1764,N_14114,N_14568);
nand UO_1765 (O_1765,N_14372,N_14884);
nor UO_1766 (O_1766,N_14459,N_14135);
nor UO_1767 (O_1767,N_14945,N_14443);
or UO_1768 (O_1768,N_14433,N_14307);
nor UO_1769 (O_1769,N_14718,N_14138);
or UO_1770 (O_1770,N_14708,N_14546);
and UO_1771 (O_1771,N_14424,N_14895);
or UO_1772 (O_1772,N_14056,N_14756);
nor UO_1773 (O_1773,N_14923,N_14442);
nor UO_1774 (O_1774,N_14765,N_14141);
nand UO_1775 (O_1775,N_14103,N_14751);
or UO_1776 (O_1776,N_14106,N_14668);
nor UO_1777 (O_1777,N_14210,N_14872);
nor UO_1778 (O_1778,N_14443,N_14738);
and UO_1779 (O_1779,N_14608,N_14429);
or UO_1780 (O_1780,N_14017,N_14232);
xor UO_1781 (O_1781,N_14426,N_14947);
nor UO_1782 (O_1782,N_14531,N_14035);
nand UO_1783 (O_1783,N_14466,N_14652);
nand UO_1784 (O_1784,N_14416,N_14641);
nor UO_1785 (O_1785,N_14284,N_14222);
nand UO_1786 (O_1786,N_14800,N_14746);
and UO_1787 (O_1787,N_14830,N_14915);
xor UO_1788 (O_1788,N_14974,N_14984);
nor UO_1789 (O_1789,N_14183,N_14439);
and UO_1790 (O_1790,N_14051,N_14404);
or UO_1791 (O_1791,N_14400,N_14808);
nor UO_1792 (O_1792,N_14499,N_14691);
xor UO_1793 (O_1793,N_14323,N_14982);
nor UO_1794 (O_1794,N_14548,N_14361);
nor UO_1795 (O_1795,N_14918,N_14177);
nor UO_1796 (O_1796,N_14003,N_14361);
and UO_1797 (O_1797,N_14600,N_14877);
or UO_1798 (O_1798,N_14432,N_14318);
nor UO_1799 (O_1799,N_14902,N_14892);
or UO_1800 (O_1800,N_14792,N_14170);
nor UO_1801 (O_1801,N_14849,N_14675);
or UO_1802 (O_1802,N_14840,N_14395);
or UO_1803 (O_1803,N_14930,N_14496);
nor UO_1804 (O_1804,N_14789,N_14002);
or UO_1805 (O_1805,N_14071,N_14596);
and UO_1806 (O_1806,N_14375,N_14847);
nor UO_1807 (O_1807,N_14359,N_14713);
nor UO_1808 (O_1808,N_14728,N_14223);
or UO_1809 (O_1809,N_14051,N_14947);
and UO_1810 (O_1810,N_14706,N_14191);
xor UO_1811 (O_1811,N_14504,N_14242);
and UO_1812 (O_1812,N_14769,N_14081);
xor UO_1813 (O_1813,N_14002,N_14412);
xnor UO_1814 (O_1814,N_14722,N_14685);
and UO_1815 (O_1815,N_14276,N_14040);
or UO_1816 (O_1816,N_14402,N_14033);
or UO_1817 (O_1817,N_14554,N_14976);
nand UO_1818 (O_1818,N_14171,N_14020);
xor UO_1819 (O_1819,N_14198,N_14115);
xnor UO_1820 (O_1820,N_14611,N_14797);
nor UO_1821 (O_1821,N_14283,N_14055);
and UO_1822 (O_1822,N_14562,N_14862);
nand UO_1823 (O_1823,N_14995,N_14308);
nor UO_1824 (O_1824,N_14994,N_14690);
nor UO_1825 (O_1825,N_14915,N_14998);
nor UO_1826 (O_1826,N_14256,N_14127);
nand UO_1827 (O_1827,N_14620,N_14695);
and UO_1828 (O_1828,N_14953,N_14599);
or UO_1829 (O_1829,N_14544,N_14018);
and UO_1830 (O_1830,N_14987,N_14492);
xor UO_1831 (O_1831,N_14619,N_14536);
and UO_1832 (O_1832,N_14190,N_14923);
nand UO_1833 (O_1833,N_14946,N_14760);
nand UO_1834 (O_1834,N_14642,N_14680);
nand UO_1835 (O_1835,N_14537,N_14727);
nor UO_1836 (O_1836,N_14445,N_14791);
nor UO_1837 (O_1837,N_14754,N_14134);
nand UO_1838 (O_1838,N_14899,N_14172);
xor UO_1839 (O_1839,N_14337,N_14145);
nor UO_1840 (O_1840,N_14579,N_14025);
nor UO_1841 (O_1841,N_14582,N_14627);
nor UO_1842 (O_1842,N_14147,N_14833);
nor UO_1843 (O_1843,N_14716,N_14815);
or UO_1844 (O_1844,N_14227,N_14094);
and UO_1845 (O_1845,N_14515,N_14755);
nand UO_1846 (O_1846,N_14912,N_14414);
or UO_1847 (O_1847,N_14287,N_14221);
and UO_1848 (O_1848,N_14563,N_14772);
or UO_1849 (O_1849,N_14918,N_14602);
nor UO_1850 (O_1850,N_14174,N_14819);
xnor UO_1851 (O_1851,N_14922,N_14587);
nand UO_1852 (O_1852,N_14035,N_14768);
nor UO_1853 (O_1853,N_14080,N_14502);
nor UO_1854 (O_1854,N_14751,N_14140);
nor UO_1855 (O_1855,N_14052,N_14024);
and UO_1856 (O_1856,N_14127,N_14465);
or UO_1857 (O_1857,N_14489,N_14099);
nor UO_1858 (O_1858,N_14160,N_14422);
or UO_1859 (O_1859,N_14831,N_14229);
nand UO_1860 (O_1860,N_14203,N_14169);
nand UO_1861 (O_1861,N_14141,N_14500);
or UO_1862 (O_1862,N_14161,N_14295);
or UO_1863 (O_1863,N_14225,N_14241);
or UO_1864 (O_1864,N_14728,N_14696);
or UO_1865 (O_1865,N_14271,N_14091);
nor UO_1866 (O_1866,N_14798,N_14538);
nor UO_1867 (O_1867,N_14566,N_14298);
xnor UO_1868 (O_1868,N_14715,N_14543);
and UO_1869 (O_1869,N_14722,N_14262);
nor UO_1870 (O_1870,N_14593,N_14483);
nand UO_1871 (O_1871,N_14067,N_14963);
xnor UO_1872 (O_1872,N_14469,N_14013);
xnor UO_1873 (O_1873,N_14102,N_14012);
and UO_1874 (O_1874,N_14232,N_14365);
and UO_1875 (O_1875,N_14341,N_14256);
and UO_1876 (O_1876,N_14206,N_14444);
or UO_1877 (O_1877,N_14820,N_14930);
and UO_1878 (O_1878,N_14917,N_14679);
or UO_1879 (O_1879,N_14379,N_14928);
xor UO_1880 (O_1880,N_14938,N_14981);
nand UO_1881 (O_1881,N_14067,N_14390);
nor UO_1882 (O_1882,N_14535,N_14171);
nand UO_1883 (O_1883,N_14408,N_14776);
nor UO_1884 (O_1884,N_14548,N_14358);
or UO_1885 (O_1885,N_14520,N_14695);
xor UO_1886 (O_1886,N_14802,N_14471);
xnor UO_1887 (O_1887,N_14894,N_14511);
and UO_1888 (O_1888,N_14192,N_14579);
nor UO_1889 (O_1889,N_14325,N_14246);
and UO_1890 (O_1890,N_14954,N_14017);
nand UO_1891 (O_1891,N_14791,N_14702);
or UO_1892 (O_1892,N_14615,N_14232);
nor UO_1893 (O_1893,N_14864,N_14891);
or UO_1894 (O_1894,N_14940,N_14706);
nand UO_1895 (O_1895,N_14830,N_14590);
or UO_1896 (O_1896,N_14538,N_14351);
or UO_1897 (O_1897,N_14250,N_14602);
or UO_1898 (O_1898,N_14690,N_14958);
xor UO_1899 (O_1899,N_14142,N_14815);
or UO_1900 (O_1900,N_14816,N_14443);
nand UO_1901 (O_1901,N_14578,N_14133);
and UO_1902 (O_1902,N_14064,N_14320);
nand UO_1903 (O_1903,N_14606,N_14276);
nor UO_1904 (O_1904,N_14483,N_14410);
xnor UO_1905 (O_1905,N_14942,N_14710);
and UO_1906 (O_1906,N_14444,N_14172);
or UO_1907 (O_1907,N_14555,N_14238);
and UO_1908 (O_1908,N_14976,N_14257);
or UO_1909 (O_1909,N_14529,N_14771);
and UO_1910 (O_1910,N_14101,N_14401);
nand UO_1911 (O_1911,N_14310,N_14355);
or UO_1912 (O_1912,N_14246,N_14798);
or UO_1913 (O_1913,N_14563,N_14197);
or UO_1914 (O_1914,N_14302,N_14443);
and UO_1915 (O_1915,N_14606,N_14931);
nand UO_1916 (O_1916,N_14593,N_14006);
and UO_1917 (O_1917,N_14185,N_14158);
nor UO_1918 (O_1918,N_14262,N_14057);
and UO_1919 (O_1919,N_14383,N_14733);
nand UO_1920 (O_1920,N_14641,N_14596);
xnor UO_1921 (O_1921,N_14561,N_14678);
or UO_1922 (O_1922,N_14880,N_14987);
and UO_1923 (O_1923,N_14368,N_14379);
or UO_1924 (O_1924,N_14298,N_14130);
xor UO_1925 (O_1925,N_14970,N_14410);
xor UO_1926 (O_1926,N_14913,N_14091);
nor UO_1927 (O_1927,N_14535,N_14648);
xnor UO_1928 (O_1928,N_14340,N_14243);
nor UO_1929 (O_1929,N_14524,N_14491);
nor UO_1930 (O_1930,N_14760,N_14906);
or UO_1931 (O_1931,N_14038,N_14444);
nor UO_1932 (O_1932,N_14353,N_14298);
or UO_1933 (O_1933,N_14217,N_14718);
nor UO_1934 (O_1934,N_14443,N_14775);
nand UO_1935 (O_1935,N_14868,N_14630);
nand UO_1936 (O_1936,N_14276,N_14469);
xnor UO_1937 (O_1937,N_14515,N_14253);
nand UO_1938 (O_1938,N_14841,N_14951);
or UO_1939 (O_1939,N_14189,N_14624);
nand UO_1940 (O_1940,N_14576,N_14167);
xnor UO_1941 (O_1941,N_14906,N_14005);
and UO_1942 (O_1942,N_14126,N_14100);
or UO_1943 (O_1943,N_14200,N_14817);
or UO_1944 (O_1944,N_14668,N_14182);
or UO_1945 (O_1945,N_14331,N_14420);
or UO_1946 (O_1946,N_14430,N_14717);
and UO_1947 (O_1947,N_14852,N_14099);
nand UO_1948 (O_1948,N_14791,N_14736);
nor UO_1949 (O_1949,N_14702,N_14140);
and UO_1950 (O_1950,N_14173,N_14958);
nand UO_1951 (O_1951,N_14730,N_14048);
nand UO_1952 (O_1952,N_14127,N_14850);
nor UO_1953 (O_1953,N_14949,N_14744);
and UO_1954 (O_1954,N_14619,N_14447);
and UO_1955 (O_1955,N_14048,N_14202);
xnor UO_1956 (O_1956,N_14226,N_14152);
nand UO_1957 (O_1957,N_14137,N_14863);
nor UO_1958 (O_1958,N_14589,N_14051);
or UO_1959 (O_1959,N_14236,N_14309);
nand UO_1960 (O_1960,N_14314,N_14583);
and UO_1961 (O_1961,N_14192,N_14858);
or UO_1962 (O_1962,N_14043,N_14094);
nor UO_1963 (O_1963,N_14849,N_14904);
nor UO_1964 (O_1964,N_14972,N_14849);
nor UO_1965 (O_1965,N_14475,N_14137);
nor UO_1966 (O_1966,N_14032,N_14843);
or UO_1967 (O_1967,N_14563,N_14267);
or UO_1968 (O_1968,N_14475,N_14320);
or UO_1969 (O_1969,N_14188,N_14795);
or UO_1970 (O_1970,N_14373,N_14684);
and UO_1971 (O_1971,N_14142,N_14644);
xnor UO_1972 (O_1972,N_14496,N_14091);
nor UO_1973 (O_1973,N_14994,N_14824);
nor UO_1974 (O_1974,N_14694,N_14259);
and UO_1975 (O_1975,N_14193,N_14466);
or UO_1976 (O_1976,N_14640,N_14655);
or UO_1977 (O_1977,N_14651,N_14887);
nand UO_1978 (O_1978,N_14359,N_14618);
or UO_1979 (O_1979,N_14233,N_14530);
or UO_1980 (O_1980,N_14641,N_14590);
nand UO_1981 (O_1981,N_14489,N_14788);
nor UO_1982 (O_1982,N_14544,N_14384);
nand UO_1983 (O_1983,N_14123,N_14884);
and UO_1984 (O_1984,N_14972,N_14035);
nand UO_1985 (O_1985,N_14867,N_14610);
and UO_1986 (O_1986,N_14595,N_14864);
and UO_1987 (O_1987,N_14992,N_14761);
or UO_1988 (O_1988,N_14844,N_14824);
or UO_1989 (O_1989,N_14261,N_14456);
nand UO_1990 (O_1990,N_14216,N_14240);
nor UO_1991 (O_1991,N_14232,N_14884);
and UO_1992 (O_1992,N_14022,N_14848);
and UO_1993 (O_1993,N_14042,N_14716);
or UO_1994 (O_1994,N_14813,N_14398);
and UO_1995 (O_1995,N_14744,N_14327);
and UO_1996 (O_1996,N_14141,N_14739);
and UO_1997 (O_1997,N_14601,N_14025);
nor UO_1998 (O_1998,N_14052,N_14083);
or UO_1999 (O_1999,N_14314,N_14608);
endmodule