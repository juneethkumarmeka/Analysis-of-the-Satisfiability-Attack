module basic_3000_30000_3500_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_626,In_2237);
xnor U1 (N_1,In_1654,In_38);
xnor U2 (N_2,In_1597,In_2297);
and U3 (N_3,In_248,In_2374);
nor U4 (N_4,In_2325,In_160);
or U5 (N_5,In_530,In_387);
and U6 (N_6,In_399,In_1175);
xor U7 (N_7,In_1603,In_2951);
and U8 (N_8,In_2306,In_1650);
nor U9 (N_9,In_1489,In_1524);
or U10 (N_10,In_2668,In_260);
nand U11 (N_11,In_1308,In_481);
nor U12 (N_12,In_491,In_2858);
nand U13 (N_13,In_2528,In_1341);
nor U14 (N_14,In_2447,In_2546);
and U15 (N_15,In_2885,In_236);
xor U16 (N_16,In_1004,In_2746);
xor U17 (N_17,In_2415,In_2018);
xnor U18 (N_18,In_2023,In_91);
nand U19 (N_19,In_360,In_2117);
nor U20 (N_20,In_1198,In_613);
nor U21 (N_21,In_1362,In_2379);
nand U22 (N_22,In_737,In_2848);
nand U23 (N_23,In_1759,In_134);
nor U24 (N_24,In_1275,In_805);
and U25 (N_25,In_704,In_982);
nand U26 (N_26,In_129,In_1557);
nand U27 (N_27,In_1699,In_510);
nand U28 (N_28,In_2655,In_81);
or U29 (N_29,In_1564,In_2884);
and U30 (N_30,In_2006,In_786);
nor U31 (N_31,In_1156,In_1955);
and U32 (N_32,In_1586,In_2915);
xnor U33 (N_33,In_2444,In_2749);
nor U34 (N_34,In_65,In_2847);
nor U35 (N_35,In_1648,In_2068);
nor U36 (N_36,In_1686,In_482);
nor U37 (N_37,In_426,In_705);
and U38 (N_38,In_215,In_1729);
or U39 (N_39,In_213,In_2716);
or U40 (N_40,In_1492,In_2796);
or U41 (N_41,In_2417,In_524);
and U42 (N_42,In_128,In_2673);
or U43 (N_43,In_2704,In_87);
xnor U44 (N_44,In_2132,In_2083);
nor U45 (N_45,In_1528,In_1688);
nor U46 (N_46,In_942,In_504);
nor U47 (N_47,In_1851,In_2369);
xnor U48 (N_48,In_2700,In_1862);
or U49 (N_49,In_365,In_1289);
and U50 (N_50,In_1947,In_1779);
or U51 (N_51,In_2330,In_1908);
or U52 (N_52,In_1962,In_2945);
or U53 (N_53,In_2190,In_560);
nand U54 (N_54,In_1230,In_1536);
nand U55 (N_55,In_232,In_846);
or U56 (N_56,In_781,In_1457);
nand U57 (N_57,In_1878,In_2544);
nand U58 (N_58,In_1605,In_108);
nor U59 (N_59,In_2515,In_2824);
nor U60 (N_60,In_1455,In_2855);
nor U61 (N_61,In_442,In_1055);
nand U62 (N_62,In_540,In_1741);
nor U63 (N_63,In_1241,In_1112);
nand U64 (N_64,In_66,In_2652);
nand U65 (N_65,In_1364,In_1935);
xnor U66 (N_66,In_2961,In_340);
and U67 (N_67,In_1824,In_2856);
or U68 (N_68,In_881,In_2118);
and U69 (N_69,In_515,In_1745);
nor U70 (N_70,In_642,In_800);
or U71 (N_71,In_2553,In_2833);
or U72 (N_72,In_1171,In_1332);
or U73 (N_73,In_276,In_988);
xor U74 (N_74,In_1306,In_1937);
or U75 (N_75,In_1222,In_2743);
nor U76 (N_76,In_1003,In_2284);
and U77 (N_77,In_975,In_614);
xor U78 (N_78,In_1304,In_1563);
nand U79 (N_79,In_1429,In_559);
and U80 (N_80,In_961,In_1969);
or U81 (N_81,In_1982,In_2274);
xor U82 (N_82,In_1452,In_2577);
nand U83 (N_83,In_870,In_2108);
nand U84 (N_84,In_2597,In_840);
and U85 (N_85,In_1746,In_1555);
or U86 (N_86,In_683,In_2060);
or U87 (N_87,In_2627,In_2305);
xor U88 (N_88,In_716,In_752);
xnor U89 (N_89,In_2817,In_2794);
nand U90 (N_90,In_2017,In_674);
nor U91 (N_91,In_1122,In_1626);
nor U92 (N_92,In_845,In_563);
nor U93 (N_93,In_1981,In_2908);
and U94 (N_94,In_258,In_1795);
and U95 (N_95,In_523,In_2932);
nand U96 (N_96,In_450,In_720);
nor U97 (N_97,In_2022,In_2482);
or U98 (N_98,In_499,In_1166);
and U99 (N_99,In_83,In_1469);
nand U100 (N_100,In_2499,In_2137);
nor U101 (N_101,In_2697,In_1617);
and U102 (N_102,In_464,In_312);
or U103 (N_103,In_463,In_2027);
nand U104 (N_104,In_2396,In_2950);
or U105 (N_105,In_521,In_2557);
xnor U106 (N_106,In_2598,In_241);
and U107 (N_107,In_1726,In_132);
nor U108 (N_108,In_2150,In_1761);
nor U109 (N_109,In_2625,In_1121);
and U110 (N_110,In_1623,In_1403);
xnor U111 (N_111,In_2635,In_996);
or U112 (N_112,In_631,In_649);
xor U113 (N_113,In_2208,In_1641);
and U114 (N_114,In_2798,In_1008);
and U115 (N_115,In_2787,In_896);
or U116 (N_116,In_1702,In_1879);
and U117 (N_117,In_2064,In_832);
or U118 (N_118,In_1394,In_1507);
or U119 (N_119,In_644,In_1352);
nand U120 (N_120,In_1044,In_1393);
nand U121 (N_121,In_1372,In_2620);
xor U122 (N_122,In_410,In_591);
xnor U123 (N_123,In_147,In_2596);
nand U124 (N_124,In_174,In_2730);
nor U125 (N_125,In_130,In_1985);
or U126 (N_126,In_1833,In_1110);
xor U127 (N_127,In_956,In_133);
nor U128 (N_128,In_121,In_1900);
xnor U129 (N_129,In_18,In_2923);
or U130 (N_130,In_2383,In_778);
and U131 (N_131,In_2247,In_2760);
xnor U132 (N_132,In_884,In_583);
or U133 (N_133,In_1984,In_2633);
or U134 (N_134,In_2819,In_2203);
nor U135 (N_135,In_490,In_1343);
or U136 (N_136,In_1771,In_2810);
nand U137 (N_137,In_2928,In_952);
or U138 (N_138,In_651,In_2822);
xor U139 (N_139,In_577,In_1310);
and U140 (N_140,In_62,In_1784);
xnor U141 (N_141,In_2727,In_1443);
and U142 (N_142,In_688,In_1252);
xor U143 (N_143,In_268,In_1825);
nand U144 (N_144,In_1285,In_1178);
or U145 (N_145,In_592,In_1484);
nor U146 (N_146,In_2339,In_2636);
nor U147 (N_147,In_467,In_971);
xor U148 (N_148,In_327,In_1594);
and U149 (N_149,In_335,In_445);
and U150 (N_150,In_2734,In_873);
xnor U151 (N_151,In_1644,In_2510);
nor U152 (N_152,In_2562,In_1126);
and U153 (N_153,In_2789,In_1268);
and U154 (N_154,In_1000,In_1490);
nor U155 (N_155,In_2509,In_2493);
nor U156 (N_156,In_757,In_1047);
xor U157 (N_157,In_113,In_1711);
xnor U158 (N_158,In_461,In_1762);
or U159 (N_159,In_1899,In_2114);
nand U160 (N_160,In_97,In_2109);
and U161 (N_161,In_1284,In_2556);
nand U162 (N_162,In_615,In_1062);
and U163 (N_163,In_125,In_2438);
or U164 (N_164,In_519,In_1621);
nor U165 (N_165,In_1078,In_337);
and U166 (N_166,In_444,In_1646);
or U167 (N_167,In_1181,In_2019);
nand U168 (N_168,In_42,In_1048);
nor U169 (N_169,In_1090,In_2210);
and U170 (N_170,In_2576,In_139);
nand U171 (N_171,In_2995,In_1486);
xor U172 (N_172,In_2926,In_124);
nand U173 (N_173,In_1913,In_2702);
nand U174 (N_174,In_1829,In_2663);
xnor U175 (N_175,In_2611,In_1315);
xor U176 (N_176,In_963,In_1113);
nand U177 (N_177,In_989,In_526);
xnor U178 (N_178,In_529,In_1189);
and U179 (N_179,In_2041,In_2194);
nor U180 (N_180,In_2537,In_2260);
and U181 (N_181,In_839,In_1926);
xnor U182 (N_182,In_1465,In_842);
nor U183 (N_183,In_2497,In_2236);
xor U184 (N_184,In_403,In_1499);
or U185 (N_185,In_440,In_1141);
nand U186 (N_186,In_2650,In_1147);
nor U187 (N_187,In_566,In_2690);
xnor U188 (N_188,In_2289,In_314);
nor U189 (N_189,In_1119,In_1018);
and U190 (N_190,In_2914,In_1533);
nand U191 (N_191,In_822,In_929);
nand U192 (N_192,In_962,In_2154);
xnor U193 (N_193,In_2595,In_1590);
nand U194 (N_194,In_1059,In_2165);
or U195 (N_195,In_681,In_1625);
nand U196 (N_196,In_1517,In_935);
xor U197 (N_197,In_111,In_162);
nand U198 (N_198,In_2474,In_2197);
xor U199 (N_199,In_1250,In_2823);
and U200 (N_200,In_1948,In_2192);
nor U201 (N_201,In_2138,In_696);
and U202 (N_202,In_1753,In_2917);
and U203 (N_203,In_1389,In_907);
or U204 (N_204,In_2622,In_1548);
or U205 (N_205,In_1973,In_1397);
nor U206 (N_206,In_386,In_2464);
nor U207 (N_207,In_1838,In_2178);
nor U208 (N_208,In_34,In_1731);
nand U209 (N_209,In_1087,In_1693);
nor U210 (N_210,In_1440,In_2678);
nand U211 (N_211,In_188,In_738);
or U212 (N_212,In_345,In_1763);
and U213 (N_213,In_787,In_1260);
and U214 (N_214,In_1420,In_2573);
and U215 (N_215,In_2454,In_921);
nand U216 (N_216,In_293,In_1127);
xor U217 (N_217,In_1464,In_578);
nor U218 (N_218,In_2968,In_2451);
or U219 (N_219,In_671,In_905);
or U220 (N_220,In_430,In_2840);
xnor U221 (N_221,In_1886,In_2616);
xnor U222 (N_222,In_2922,In_1842);
nor U223 (N_223,In_1167,In_2147);
nor U224 (N_224,In_2867,In_2412);
or U225 (N_225,In_2722,In_2095);
and U226 (N_226,In_2773,In_2066);
or U227 (N_227,In_718,In_1019);
nand U228 (N_228,In_1498,In_1082);
or U229 (N_229,In_2039,In_930);
and U230 (N_230,In_900,In_1506);
xor U231 (N_231,In_2176,In_92);
and U232 (N_232,In_2987,In_1521);
and U233 (N_233,In_2632,In_173);
nor U234 (N_234,In_1334,In_2930);
xnor U235 (N_235,In_2093,In_1470);
nand U236 (N_236,In_2389,In_295);
nand U237 (N_237,In_2301,In_137);
xor U238 (N_238,In_1054,In_2313);
or U239 (N_239,In_2771,In_175);
xor U240 (N_240,In_1211,In_191);
and U241 (N_241,In_2708,In_497);
and U242 (N_242,In_1321,In_2029);
xnor U243 (N_243,In_35,In_707);
and U244 (N_244,In_1559,In_1724);
nor U245 (N_245,In_1925,In_1337);
or U246 (N_246,In_2335,In_808);
nand U247 (N_247,In_747,In_19);
or U248 (N_248,In_182,In_2872);
nor U249 (N_249,In_909,In_2554);
nor U250 (N_250,In_1235,In_2326);
xor U251 (N_251,In_1581,In_1800);
xnor U252 (N_252,In_1149,In_2278);
nor U253 (N_253,In_1298,In_872);
nor U254 (N_254,In_885,In_2988);
or U255 (N_255,In_2759,In_294);
or U256 (N_256,In_1927,In_120);
nor U257 (N_257,In_2549,In_1379);
nor U258 (N_258,In_2900,In_927);
xor U259 (N_259,In_2607,In_648);
and U260 (N_260,In_149,In_2662);
nor U261 (N_261,In_831,In_94);
nand U262 (N_262,In_486,In_2624);
and U263 (N_263,In_730,In_2099);
or U264 (N_264,In_2223,In_1497);
nor U265 (N_265,In_1042,In_939);
nor U266 (N_266,In_2048,In_871);
xnor U267 (N_267,In_1382,In_46);
or U268 (N_268,In_910,In_2879);
xnor U269 (N_269,In_2707,In_355);
xnor U270 (N_270,In_1238,In_922);
nor U271 (N_271,In_1953,In_409);
nor U272 (N_272,In_1173,In_1084);
nor U273 (N_273,In_902,In_416);
nor U274 (N_274,In_1651,In_154);
nand U275 (N_275,In_257,In_1154);
xnor U276 (N_276,In_2986,In_1602);
and U277 (N_277,In_1125,In_2906);
nand U278 (N_278,In_1013,In_1116);
nor U279 (N_279,In_633,In_2084);
nor U280 (N_280,In_2449,In_2929);
nor U281 (N_281,In_2242,In_1647);
or U282 (N_282,In_261,In_2845);
xnor U283 (N_283,In_632,In_955);
or U284 (N_284,In_1229,In_965);
xnor U285 (N_285,In_1271,In_1277);
nand U286 (N_286,In_2251,In_702);
nor U287 (N_287,In_1854,In_520);
or U288 (N_288,In_2256,In_1278);
nor U289 (N_289,In_2529,In_2762);
nand U290 (N_290,In_472,In_447);
and U291 (N_291,In_793,In_1653);
nor U292 (N_292,In_677,In_1295);
and U293 (N_293,In_2641,In_1200);
xnor U294 (N_294,In_1801,In_2228);
nand U295 (N_295,In_1424,In_2680);
or U296 (N_296,In_2045,In_433);
or U297 (N_297,In_2846,In_2955);
xor U298 (N_298,In_685,In_675);
xor U299 (N_299,In_1155,In_1613);
nor U300 (N_300,In_2784,In_1012);
or U301 (N_301,In_682,In_2857);
nand U302 (N_302,In_1328,In_1205);
xor U303 (N_303,In_1709,In_1259);
xnor U304 (N_304,In_2631,In_1704);
nand U305 (N_305,In_2752,In_2468);
nor U306 (N_306,In_724,In_2455);
xnor U307 (N_307,In_1811,In_251);
or U308 (N_308,In_2070,In_1441);
nor U309 (N_309,In_2937,In_2429);
nor U310 (N_310,In_2504,In_383);
xnor U311 (N_311,In_1462,In_572);
or U312 (N_312,In_513,In_2999);
nor U313 (N_313,In_1212,In_739);
nor U314 (N_314,In_2737,In_1137);
nor U315 (N_315,In_1978,In_663);
xnor U316 (N_316,In_2604,In_1512);
and U317 (N_317,In_573,In_2550);
xor U318 (N_318,In_2956,In_402);
or U319 (N_319,In_2268,In_1115);
nand U320 (N_320,In_745,In_1550);
xor U321 (N_321,In_2523,In_1383);
nor U322 (N_322,In_2698,In_226);
nor U323 (N_323,In_732,In_2740);
nand U324 (N_324,In_296,In_79);
xor U325 (N_325,In_790,In_535);
or U326 (N_326,In_1875,In_1177);
or U327 (N_327,In_1946,In_864);
nor U328 (N_328,In_2465,In_1570);
and U329 (N_329,In_369,In_2841);
nand U330 (N_330,In_1816,In_2320);
nand U331 (N_331,In_725,In_380);
or U332 (N_332,In_1301,In_629);
nor U333 (N_333,In_794,In_1952);
xnor U334 (N_334,In_2691,In_155);
xor U335 (N_335,In_378,In_2500);
xor U336 (N_336,In_1596,In_2225);
and U337 (N_337,In_1448,In_1708);
or U338 (N_338,In_2940,In_2938);
or U339 (N_339,In_813,In_1544);
or U340 (N_340,In_1808,In_2842);
nand U341 (N_341,In_2074,In_2234);
or U342 (N_342,In_51,In_1031);
nand U343 (N_343,In_2891,In_1575);
nor U344 (N_344,In_1216,In_824);
xor U345 (N_345,In_1002,In_2993);
xor U346 (N_346,In_1942,In_1234);
or U347 (N_347,In_2984,In_356);
nand U348 (N_348,In_61,In_1244);
nor U349 (N_349,In_2912,In_2100);
and U350 (N_350,In_2839,In_1355);
nor U351 (N_351,In_2209,In_503);
nand U352 (N_352,In_2222,In_1138);
nor U353 (N_353,In_1302,In_1923);
and U354 (N_354,In_853,In_7);
or U355 (N_355,In_934,In_986);
nor U356 (N_356,In_1583,In_2016);
nand U357 (N_357,In_2484,In_2411);
nand U358 (N_358,In_1860,In_2795);
xor U359 (N_359,In_1805,In_2457);
xor U360 (N_360,In_2925,In_2776);
or U361 (N_361,In_1695,In_1773);
nor U362 (N_362,In_2766,In_286);
nor U363 (N_363,In_695,In_2426);
or U364 (N_364,In_1066,In_1209);
nor U365 (N_365,In_2127,In_1676);
nand U366 (N_366,In_1399,In_2913);
nand U367 (N_367,In_2719,In_2931);
nor U368 (N_368,In_1100,In_1416);
xor U369 (N_369,In_1819,In_1427);
nand U370 (N_370,In_1672,In_575);
and U371 (N_371,In_653,In_557);
and U372 (N_372,In_377,In_814);
xnor U373 (N_373,In_1485,In_2807);
nor U374 (N_374,In_2187,In_2407);
xnor U375 (N_375,In_917,In_1656);
xor U376 (N_376,In_301,In_799);
nand U377 (N_377,In_954,In_1894);
xor U378 (N_378,In_1188,In_471);
xor U379 (N_379,In_165,In_2543);
or U380 (N_380,In_2312,In_668);
or U381 (N_381,In_2646,In_2303);
nor U382 (N_382,In_2958,In_366);
xnor U383 (N_383,In_1351,In_2976);
nand U384 (N_384,In_2503,In_820);
or U385 (N_385,In_1917,In_2207);
xor U386 (N_386,In_1589,In_782);
xnor U387 (N_387,In_2978,In_1451);
and U388 (N_388,In_2753,In_553);
nor U389 (N_389,In_1700,In_1560);
or U390 (N_390,In_999,In_1273);
or U391 (N_391,In_2801,In_2649);
and U392 (N_392,In_2825,In_2448);
nor U393 (N_393,In_2878,In_874);
or U394 (N_394,In_2123,In_2460);
or U395 (N_395,In_652,In_539);
nand U396 (N_396,In_906,In_1823);
or U397 (N_397,In_266,In_1099);
nor U398 (N_398,In_2096,In_2140);
and U399 (N_399,In_2952,In_2894);
nand U400 (N_400,In_285,In_744);
and U401 (N_401,In_1515,In_496);
nor U402 (N_402,In_1233,In_607);
nand U403 (N_403,In_546,In_895);
and U404 (N_404,In_1245,In_21);
xnor U405 (N_405,In_2648,In_2381);
xnor U406 (N_406,In_765,In_1006);
nand U407 (N_407,In_2443,In_396);
and U408 (N_408,In_2145,In_1929);
and U409 (N_409,In_847,In_897);
and U410 (N_410,In_2059,In_280);
and U411 (N_411,In_2693,In_2670);
xor U412 (N_412,In_536,In_2715);
xnor U413 (N_413,In_1297,In_1776);
or U414 (N_414,In_2015,In_2469);
or U415 (N_415,In_1627,In_2805);
and U416 (N_416,In_1170,In_2399);
xnor U417 (N_417,In_2416,In_1785);
or U418 (N_418,In_2397,In_379);
nand U419 (N_419,In_2488,In_689);
nand U420 (N_420,In_142,In_2492);
nand U421 (N_421,In_415,In_1293);
and U422 (N_422,In_2600,In_2370);
xnor U423 (N_423,In_2647,In_2072);
xor U424 (N_424,In_1701,In_2115);
nand U425 (N_425,In_586,In_525);
nor U426 (N_426,In_1069,In_1354);
and U427 (N_427,In_918,In_2821);
nand U428 (N_428,In_1941,In_100);
nor U429 (N_429,In_2861,In_2);
and U430 (N_430,In_1643,In_508);
or U431 (N_431,In_405,In_1531);
or U432 (N_432,In_1760,In_1057);
xnor U433 (N_433,In_1685,In_723);
nand U434 (N_434,In_2220,In_2037);
nand U435 (N_435,In_1798,In_1208);
or U436 (N_436,In_1777,In_2706);
or U437 (N_437,In_1479,In_784);
nor U438 (N_438,In_2248,In_584);
nand U439 (N_439,In_1096,In_1949);
or U440 (N_440,In_2479,In_623);
xor U441 (N_441,In_1148,In_2713);
xnor U442 (N_442,In_1659,In_197);
or U443 (N_443,In_2161,In_2677);
nand U444 (N_444,In_987,In_2402);
and U445 (N_445,In_1938,In_1494);
nand U446 (N_446,In_1979,In_1053);
and U447 (N_447,In_889,In_2263);
nor U448 (N_448,In_1599,In_522);
nand U449 (N_449,In_341,In_2026);
or U450 (N_450,In_1015,In_1669);
nand U451 (N_451,In_391,In_1320);
xor U452 (N_452,In_579,In_818);
nand U453 (N_453,In_1791,In_2347);
nand U454 (N_454,In_227,In_562);
xnor U455 (N_455,In_2282,In_2036);
nor U456 (N_456,In_2215,In_158);
or U457 (N_457,In_1718,In_2896);
xnor U458 (N_458,In_2491,In_284);
xnor U459 (N_459,In_1614,In_710);
nor U460 (N_460,In_736,In_1050);
nand U461 (N_461,In_2486,In_145);
nand U462 (N_462,In_2583,In_899);
nor U463 (N_463,In_1906,In_2615);
or U464 (N_464,In_587,In_1963);
nand U465 (N_465,In_231,In_45);
xor U466 (N_466,In_1561,In_1265);
xor U467 (N_467,In_2097,In_1770);
or U468 (N_468,In_1580,In_1142);
nor U469 (N_469,In_2395,In_833);
xor U470 (N_470,In_2404,In_2349);
xnor U471 (N_471,In_1638,In_2078);
xnor U472 (N_472,In_2466,In_979);
nor U473 (N_473,In_518,In_1687);
or U474 (N_474,In_502,In_1950);
nor U475 (N_475,In_2139,In_2360);
nand U476 (N_476,In_1020,In_2131);
xor U477 (N_477,In_2832,In_1859);
nor U478 (N_478,In_2869,In_753);
xnor U479 (N_479,In_2392,In_2254);
and U480 (N_480,In_1989,In_2934);
xor U481 (N_481,In_119,In_662);
nor U482 (N_482,In_2315,In_1312);
or U483 (N_483,In_235,In_382);
nor U484 (N_484,In_1966,In_126);
or U485 (N_485,In_49,In_347);
or U486 (N_486,In_828,In_1442);
or U487 (N_487,In_2262,In_679);
xnor U488 (N_488,In_2258,In_2136);
xor U489 (N_489,In_2024,In_1324);
nor U490 (N_490,In_1192,In_2590);
nand U491 (N_491,In_2920,In_620);
and U492 (N_492,In_1483,In_2643);
nor U493 (N_493,In_2324,In_362);
nand U494 (N_494,In_2329,In_2195);
or U495 (N_495,In_2902,In_2682);
or U496 (N_496,In_2889,In_2681);
and U497 (N_497,In_2566,In_1505);
and U498 (N_498,In_621,In_931);
and U499 (N_499,In_10,In_1475);
nor U500 (N_500,In_2560,In_63);
nand U501 (N_501,In_1794,In_1153);
or U502 (N_502,In_229,In_1123);
nand U503 (N_503,In_2198,In_390);
or U504 (N_504,In_1056,In_1677);
nand U505 (N_505,In_1689,In_2782);
nor U506 (N_506,In_1080,In_460);
xor U507 (N_507,In_2882,In_2877);
nor U508 (N_508,In_945,In_2501);
nor U509 (N_509,In_2113,In_1288);
xnor U510 (N_510,In_2703,In_1679);
or U511 (N_511,In_977,In_1832);
and U512 (N_512,In_2744,In_849);
xor U513 (N_513,In_1,In_2992);
or U514 (N_514,In_2799,In_2695);
nand U515 (N_515,In_740,In_2375);
or U516 (N_516,In_206,In_748);
nor U517 (N_517,In_1916,In_2935);
and U518 (N_518,In_1025,In_2300);
xnor U519 (N_519,In_135,In_427);
xor U520 (N_520,In_1114,In_1573);
and U521 (N_521,In_1678,In_1311);
or U522 (N_522,In_2101,In_1458);
nor U523 (N_523,In_207,In_2519);
nand U524 (N_524,In_2255,In_1487);
nand U525 (N_525,In_2480,In_2812);
xor U526 (N_526,In_2572,In_2711);
and U527 (N_527,In_2494,In_507);
xor U528 (N_528,In_703,In_2831);
nor U529 (N_529,In_264,In_255);
or U530 (N_530,In_2747,In_1028);
or U531 (N_531,In_24,In_2838);
and U532 (N_532,In_1749,In_1620);
or U533 (N_533,In_532,In_2818);
or U534 (N_534,In_1390,In_1522);
or U535 (N_535,In_452,In_2605);
or U536 (N_536,In_2151,In_2149);
nor U537 (N_537,In_2327,In_1782);
or U538 (N_538,In_2265,In_289);
nor U539 (N_539,In_1045,In_2963);
nor U540 (N_540,In_1697,In_1595);
nand U541 (N_541,In_1291,In_1450);
xor U542 (N_542,In_2343,In_43);
nor U543 (N_543,In_1977,In_319);
or U544 (N_544,In_205,In_2126);
or U545 (N_545,In_1437,In_2267);
xnor U546 (N_546,In_346,In_2245);
and U547 (N_547,In_856,In_333);
nand U548 (N_548,In_1616,In_1772);
or U549 (N_549,In_271,In_250);
xnor U550 (N_550,In_997,In_2754);
and U551 (N_551,In_23,In_2458);
nor U552 (N_552,In_302,In_252);
and U553 (N_553,In_883,In_1592);
xor U554 (N_554,In_2110,In_1796);
and U555 (N_555,In_434,In_136);
nand U556 (N_556,In_422,In_2204);
nor U557 (N_557,In_2828,In_1511);
or U558 (N_558,In_300,In_1500);
nor U559 (N_559,In_1593,In_2233);
nor U560 (N_560,In_1675,In_680);
nand U561 (N_561,In_804,In_843);
xnor U562 (N_562,In_2621,In_2792);
xnor U563 (N_563,In_1435,In_2240);
nand U564 (N_564,In_2384,In_2299);
or U565 (N_565,In_1109,In_2013);
xnor U566 (N_566,In_763,In_2954);
or U567 (N_567,In_454,In_2973);
xnor U568 (N_568,In_352,In_1107);
nand U569 (N_569,In_2445,In_322);
nand U570 (N_570,In_2167,In_1662);
or U571 (N_571,In_2053,In_969);
nand U572 (N_572,In_116,In_1964);
and U573 (N_573,In_363,In_2852);
or U574 (N_574,In_400,In_2400);
and U575 (N_575,In_699,In_2946);
and U576 (N_576,In_990,In_1806);
or U577 (N_577,In_200,In_411);
xor U578 (N_578,In_789,In_611);
or U579 (N_579,In_2319,In_2196);
and U580 (N_580,In_2579,In_265);
and U581 (N_581,In_1388,In_890);
xnor U582 (N_582,In_1279,In_2541);
nand U583 (N_583,In_2073,In_2067);
xor U584 (N_584,In_2378,In_978);
xnor U585 (N_585,In_938,In_1566);
nor U586 (N_586,In_1921,In_476);
and U587 (N_587,In_2345,In_2214);
or U588 (N_588,In_1344,In_194);
or U589 (N_589,In_983,In_1992);
nor U590 (N_590,In_2134,In_2058);
and U591 (N_591,In_1579,In_2243);
xor U592 (N_592,In_1889,In_169);
nand U593 (N_593,In_2974,In_801);
and U594 (N_594,In_2962,In_2285);
nor U595 (N_595,In_774,In_2475);
xor U596 (N_596,In_329,In_2811);
xnor U597 (N_597,In_2296,In_1108);
nor U598 (N_598,In_1185,In_1671);
and U599 (N_599,In_2564,In_1079);
xor U600 (N_600,In_1890,In_2337);
and U601 (N_601,In_1748,In_798);
nand U602 (N_602,In_2069,In_1360);
nor U603 (N_603,In_1095,In_273);
xor U604 (N_604,In_1775,In_1914);
xor U605 (N_605,In_17,In_1706);
nand U606 (N_606,In_2336,In_221);
xnor U607 (N_607,In_1674,In_1714);
xor U608 (N_608,In_1282,In_531);
and U609 (N_609,In_545,In_2169);
or U610 (N_610,In_604,In_1600);
nor U611 (N_611,In_2390,In_1404);
xnor U612 (N_612,In_1491,In_1545);
or U613 (N_613,In_1228,In_179);
or U614 (N_614,In_1719,In_880);
nor U615 (N_615,In_2205,In_1024);
nor U616 (N_616,In_1329,In_59);
and U617 (N_617,In_2413,In_555);
or U618 (N_618,In_2514,In_1601);
nor U619 (N_619,In_937,In_2009);
nand U620 (N_620,In_1117,In_2183);
and U621 (N_621,In_1051,In_1132);
xor U622 (N_622,In_941,In_2410);
or U623 (N_623,In_2216,In_719);
and U624 (N_624,In_2362,In_1027);
and U625 (N_625,In_166,In_107);
xnor U626 (N_626,In_1172,In_1454);
nand U627 (N_627,In_2614,In_1248);
and U628 (N_628,In_807,In_1530);
nand U629 (N_629,In_157,In_1033);
and U630 (N_630,In_1961,In_146);
or U631 (N_631,In_755,In_1349);
nand U632 (N_632,In_2774,In_636);
nor U633 (N_633,In_2808,In_423);
xor U634 (N_634,In_1131,In_949);
nor U635 (N_635,In_244,In_2526);
or U636 (N_636,In_1920,In_1904);
and U637 (N_637,In_278,In_1182);
and U638 (N_638,In_60,In_1303);
and U639 (N_639,In_771,In_542);
xor U640 (N_640,In_2212,In_2664);
nand U641 (N_641,In_180,In_2323);
and U642 (N_642,In_1384,In_1335);
xor U643 (N_643,In_438,In_2477);
xor U644 (N_644,In_878,In_1857);
nand U645 (N_645,In_96,In_71);
or U646 (N_646,In_2534,In_773);
and U647 (N_647,In_2143,In_1846);
nand U648 (N_648,In_1813,In_767);
or U649 (N_649,In_2440,In_1827);
or U650 (N_650,In_1867,In_1480);
nand U651 (N_651,In_2542,In_1036);
or U652 (N_652,In_893,In_105);
xor U653 (N_653,In_1826,In_246);
nor U654 (N_654,In_851,In_2219);
or U655 (N_655,In_1543,In_2276);
or U656 (N_656,In_1294,In_1309);
nand U657 (N_657,In_211,In_164);
and U658 (N_658,In_331,In_14);
xor U659 (N_659,In_2102,In_2116);
nand U660 (N_660,In_2269,In_2660);
nor U661 (N_661,In_354,In_1016);
and U662 (N_662,In_230,In_2314);
nand U663 (N_663,In_2133,In_612);
or U664 (N_664,In_1135,In_2121);
nor U665 (N_665,In_691,In_2436);
and U666 (N_666,In_484,In_2521);
and U667 (N_667,In_1227,In_676);
or U668 (N_668,In_1598,In_2406);
nor U669 (N_669,In_694,In_1348);
or U670 (N_670,In_2270,In_2424);
xor U671 (N_671,In_2899,In_2351);
and U672 (N_672,In_1307,In_358);
xnor U673 (N_673,In_817,In_1768);
nor U674 (N_674,In_2859,In_1873);
nor U675 (N_675,In_1258,In_2283);
nor U676 (N_676,In_1007,In_1196);
nor U677 (N_677,In_1658,In_2683);
nor U678 (N_678,In_2569,In_721);
or U679 (N_679,In_2666,In_1591);
nor U680 (N_680,In_2651,In_1068);
xnor U681 (N_681,In_877,In_2348);
nand U682 (N_682,In_574,In_1128);
nor U683 (N_683,In_2478,In_2062);
and U684 (N_684,In_210,In_2777);
or U685 (N_685,In_1254,In_1280);
and U686 (N_686,In_1206,In_48);
and U687 (N_687,In_446,In_1738);
and U688 (N_688,In_1060,In_228);
or U689 (N_689,In_1326,In_1035);
nand U690 (N_690,In_441,In_1852);
nand U691 (N_691,In_974,In_728);
xnor U692 (N_692,In_666,In_2786);
nand U693 (N_693,In_2441,In_2403);
or U694 (N_694,In_534,In_1692);
xor U695 (N_695,In_2189,In_1990);
or U696 (N_696,In_332,In_1632);
nand U697 (N_697,In_2342,In_2586);
and U698 (N_698,In_2174,In_1014);
or U699 (N_699,In_1267,In_2830);
nor U700 (N_700,In_1997,In_810);
nor U701 (N_701,In_879,In_1615);
nor U702 (N_702,In_759,In_686);
and U703 (N_703,In_1144,In_2532);
nor U704 (N_704,In_1504,In_2603);
nand U705 (N_705,In_2368,In_1569);
and U706 (N_706,In_550,In_2050);
or U707 (N_707,In_1408,In_406);
nand U708 (N_708,In_2046,In_104);
and U709 (N_709,In_684,In_894);
xor U710 (N_710,In_225,In_152);
and U711 (N_711,In_2538,In_234);
xor U712 (N_712,In_970,In_1664);
and U713 (N_713,In_2476,In_1224);
nor U714 (N_714,In_859,In_30);
nor U715 (N_715,In_1363,In_109);
or U716 (N_716,In_928,In_1882);
xnor U717 (N_717,In_1263,In_1970);
xnor U718 (N_718,In_898,In_960);
nor U719 (N_719,In_548,In_891);
nand U720 (N_720,In_1568,In_2990);
nand U721 (N_721,In_2814,In_404);
or U722 (N_722,In_1866,In_1912);
nor U723 (N_723,In_1089,In_2675);
nand U724 (N_724,In_1169,In_2281);
and U725 (N_725,In_1778,In_2177);
nor U726 (N_726,In_2077,In_1370);
and U727 (N_727,In_2977,In_1939);
and U728 (N_728,In_599,In_1077);
nor U729 (N_729,In_1553,In_588);
or U730 (N_730,In_2261,In_754);
nor U731 (N_731,In_1323,In_2338);
nand U732 (N_732,In_2609,In_2439);
nand U733 (N_733,In_758,In_1377);
nor U734 (N_734,In_2040,In_361);
nor U735 (N_735,In_597,In_1965);
xor U736 (N_736,In_1657,In_2235);
nand U737 (N_737,In_1835,In_1769);
nand U738 (N_738,In_1988,In_514);
nand U739 (N_739,In_217,In_2629);
nand U740 (N_740,In_1163,In_2640);
nand U741 (N_741,In_1831,In_1136);
xnor U742 (N_742,In_1502,In_313);
nor U743 (N_743,In_2409,In_2302);
nor U744 (N_744,In_1915,In_1338);
xor U745 (N_745,In_2667,In_1735);
nor U746 (N_746,In_2051,In_1532);
and U747 (N_747,In_1237,In_1634);
nand U748 (N_748,In_625,In_2052);
nor U749 (N_749,In_2989,In_1839);
or U750 (N_750,In_141,In_2244);
or U751 (N_751,In_1176,In_857);
xor U752 (N_752,In_1604,In_2853);
xor U753 (N_753,In_2718,In_1426);
and U754 (N_754,In_1733,In_373);
or U755 (N_755,In_186,In_2739);
nor U756 (N_756,In_488,In_1804);
nand U757 (N_757,In_2525,In_590);
or U758 (N_758,In_1742,In_1877);
nor U759 (N_759,In_2393,In_1821);
nor U760 (N_760,In_700,In_1305);
nor U761 (N_761,In_2813,In_985);
xor U762 (N_762,In_2405,In_2571);
or U763 (N_763,In_1339,In_1174);
and U764 (N_764,In_123,In_1752);
nand U765 (N_765,In_1064,In_2211);
or U766 (N_766,In_1681,In_1204);
nor U767 (N_767,In_1898,In_2639);
nand U768 (N_768,In_2717,In_1134);
or U769 (N_769,In_469,In_2071);
or U770 (N_770,In_2008,In_1052);
nand U771 (N_771,In_1909,In_2981);
and U772 (N_772,In_627,In_2307);
nand U773 (N_773,In_2456,In_2076);
nand U774 (N_774,In_722,In_6);
or U775 (N_775,In_2094,In_209);
and U776 (N_776,In_2608,In_742);
xnor U777 (N_777,In_1928,In_1191);
xnor U778 (N_778,In_1865,In_2991);
or U779 (N_779,In_1931,In_2876);
or U780 (N_780,In_2275,In_1510);
nand U781 (N_781,In_85,In_2788);
and U782 (N_782,In_1802,In_1286);
nor U783 (N_783,In_1300,In_1814);
and U784 (N_784,In_1509,In_2103);
or U785 (N_785,In_315,In_2522);
or U786 (N_786,In_1438,In_1070);
and U787 (N_787,In_310,In_1612);
or U788 (N_788,In_1385,In_1145);
xor U789 (N_789,In_1959,In_171);
nand U790 (N_790,In_192,In_852);
xor U791 (N_791,In_769,In_2295);
xnor U792 (N_792,In_20,In_1151);
nand U793 (N_793,In_2536,In_1870);
and U794 (N_794,In_2129,In_1133);
nor U795 (N_795,In_498,In_2088);
xor U796 (N_796,In_561,In_281);
and U797 (N_797,In_993,In_53);
nand U798 (N_798,In_2567,In_2893);
xor U799 (N_799,In_622,In_1986);
xor U800 (N_800,In_2202,In_101);
xnor U801 (N_801,In_678,In_645);
xor U802 (N_802,In_1327,In_1951);
or U803 (N_803,In_1546,In_2696);
or U804 (N_804,In_1905,In_33);
nor U805 (N_805,In_2184,In_1812);
or U806 (N_806,In_630,In_1974);
xor U807 (N_807,In_2751,In_1140);
nor U808 (N_808,In_56,In_1392);
or U809 (N_809,In_1030,In_2701);
and U810 (N_810,In_2328,In_397);
xor U811 (N_811,In_0,In_1097);
xor U812 (N_812,In_492,In_2755);
nand U813 (N_813,In_2430,In_2548);
nand U814 (N_814,In_981,In_2511);
or U815 (N_815,In_1264,In_825);
nand U816 (N_816,In_2224,In_2943);
and U817 (N_817,In_199,In_2687);
nor U818 (N_818,In_1508,In_2520);
nor U819 (N_819,In_2152,In_1368);
and U820 (N_820,In_1933,In_635);
xnor U821 (N_821,In_2286,In_2552);
or U822 (N_822,In_2835,In_1887);
and U823 (N_823,In_1797,In_2487);
nor U824 (N_824,In_1628,In_1428);
xnor U825 (N_825,In_138,In_2002);
nand U826 (N_826,In_1043,In_1611);
nand U827 (N_827,In_2768,In_2162);
nand U828 (N_828,In_2851,In_2331);
and U829 (N_829,In_1574,In_272);
nand U830 (N_830,In_541,In_270);
xnor U831 (N_831,In_715,In_2909);
nand U832 (N_832,In_1764,In_2495);
xnor U833 (N_833,In_357,In_1609);
or U834 (N_834,In_654,In_892);
xnor U835 (N_835,In_1436,In_2619);
nor U836 (N_836,In_2054,In_220);
or U837 (N_837,In_551,In_2155);
nand U838 (N_838,In_1101,In_2180);
or U839 (N_839,In_368,In_608);
xnor U840 (N_840,In_903,In_1317);
nand U841 (N_841,In_298,In_552);
nand U842 (N_842,In_375,In_282);
nor U843 (N_843,In_2120,In_2271);
and U844 (N_844,In_1565,In_1539);
nand U845 (N_845,In_2352,In_944);
xnor U846 (N_846,In_436,In_2756);
or U847 (N_847,In_1622,In_913);
nand U848 (N_848,In_2642,In_1715);
xor U849 (N_849,In_2505,In_2874);
nor U850 (N_850,In_1331,In_2481);
nor U851 (N_851,In_1400,In_1371);
nor U852 (N_852,In_866,In_638);
nand U853 (N_853,In_2736,In_2112);
or U854 (N_854,In_1619,In_2181);
and U855 (N_855,In_1098,In_1076);
and U856 (N_856,In_1270,In_1283);
nor U857 (N_857,In_1266,In_1269);
nor U858 (N_858,In_64,In_1956);
xor U859 (N_859,In_2049,In_93);
and U860 (N_860,In_1074,In_371);
nor U861 (N_861,In_920,In_1734);
or U862 (N_862,In_320,In_1415);
or U863 (N_863,In_600,In_1158);
or U864 (N_864,In_1365,In_967);
or U865 (N_865,In_2865,In_2728);
or U866 (N_866,In_634,In_1542);
nor U867 (N_867,In_1029,In_2997);
or U868 (N_868,In_687,In_2130);
or U869 (N_869,In_1830,In_1717);
nand U870 (N_870,In_2942,In_2311);
and U871 (N_871,In_2547,In_1071);
or U872 (N_872,In_1472,In_2365);
nor U873 (N_873,In_1010,In_908);
or U874 (N_874,In_2720,In_398);
and U875 (N_875,In_487,In_1810);
xnor U876 (N_876,In_1840,In_697);
or U877 (N_877,In_2578,In_1290);
xor U878 (N_878,In_803,In_57);
xor U879 (N_879,In_2725,In_713);
nor U880 (N_880,In_172,In_1350);
or U881 (N_881,In_672,In_943);
or U882 (N_882,In_505,In_330);
xnor U883 (N_883,In_283,In_932);
xnor U884 (N_884,In_819,In_2723);
or U885 (N_885,In_1468,In_1446);
and U886 (N_886,In_2344,In_1356);
xnor U887 (N_887,In_1549,In_1380);
or U888 (N_888,In_2779,In_1065);
xnor U889 (N_889,In_495,In_1874);
nor U890 (N_890,In_304,In_760);
xor U891 (N_891,In_1316,In_923);
and U892 (N_892,In_2091,In_479);
xor U893 (N_893,In_1026,In_2775);
and U894 (N_894,In_1608,In_2081);
nand U895 (N_895,In_1246,In_2637);
or U896 (N_896,In_947,In_2570);
and U897 (N_897,In_746,In_517);
nor U898 (N_898,In_2745,In_2082);
and U899 (N_899,In_564,In_13);
nor U900 (N_900,In_1727,In_750);
xor U901 (N_901,In_238,In_1481);
and U902 (N_902,In_2257,In_1861);
and U903 (N_903,In_2031,In_1179);
or U904 (N_904,In_984,In_2014);
nand U905 (N_905,In_1124,In_1629);
xor U906 (N_906,In_1635,In_919);
or U907 (N_907,In_11,In_1432);
xnor U908 (N_908,In_198,In_1747);
nor U909 (N_909,In_384,In_483);
and U910 (N_910,In_609,In_2160);
nor U911 (N_911,In_749,In_1554);
xor U912 (N_912,In_605,In_1361);
xor U913 (N_913,In_565,In_161);
nor U914 (N_914,In_1197,In_2452);
and U915 (N_915,In_788,In_216);
and U916 (N_916,In_2781,In_106);
nor U917 (N_917,In_459,In_1256);
or U918 (N_918,In_2582,In_364);
nor U919 (N_919,In_2386,In_1325);
xor U920 (N_920,In_1240,In_1991);
and U921 (N_921,In_1187,In_770);
nand U922 (N_922,In_2229,In_661);
and U923 (N_923,In_1243,In_1022);
xor U924 (N_924,In_233,In_2689);
xor U925 (N_925,In_1847,In_1213);
nor U926 (N_926,In_177,In_570);
and U927 (N_927,In_2063,In_2437);
nand U928 (N_928,In_973,In_1527);
nor U929 (N_929,In_2250,In_2472);
nor U930 (N_930,In_1703,In_924);
nand U931 (N_931,In_1165,In_1720);
nor U932 (N_932,In_1046,In_381);
or U933 (N_933,In_708,In_2540);
and U934 (N_934,In_1571,In_2163);
and U935 (N_935,In_420,In_1111);
nand U936 (N_936,In_2653,In_964);
nor U937 (N_937,In_2959,In_2654);
or U938 (N_938,In_2030,In_2790);
xor U939 (N_939,In_2421,In_1444);
nand U940 (N_940,In_2927,In_796);
or U941 (N_941,In_1447,In_2601);
xnor U942 (N_942,In_1226,In_968);
or U943 (N_943,In_1757,In_308);
and U944 (N_944,In_1958,In_1975);
nand U945 (N_945,In_1037,In_1231);
nor U946 (N_946,In_616,In_1930);
or U947 (N_947,In_1535,In_1421);
xor U948 (N_948,In_659,In_1023);
nor U949 (N_949,In_2450,In_2422);
xnor U950 (N_950,In_465,In_88);
and U951 (N_951,In_2979,In_1094);
or U952 (N_952,In_2007,In_506);
xor U953 (N_953,In_1980,In_1844);
xor U954 (N_954,In_2433,In_2804);
xnor U955 (N_955,In_348,In_297);
nor U956 (N_956,In_589,In_1640);
and U957 (N_957,In_1017,In_2738);
nand U958 (N_958,In_1292,In_1402);
nand U959 (N_959,In_2883,In_2467);
nor U960 (N_960,In_26,In_664);
nand U961 (N_961,In_2075,In_1221);
xnor U962 (N_962,In_2965,In_291);
xnor U963 (N_963,In_2610,In_2427);
nand U964 (N_964,In_1668,In_2034);
nor U965 (N_965,In_2316,In_1691);
nor U966 (N_966,In_435,In_657);
nor U967 (N_967,In_122,In_594);
or U968 (N_968,In_1386,In_1159);
nor U969 (N_969,In_2512,In_1129);
nor U970 (N_970,In_2425,In_72);
or U971 (N_971,In_669,In_1072);
or U972 (N_972,In_82,In_527);
nor U973 (N_973,In_2135,In_1445);
and U974 (N_974,In_2969,In_243);
xor U975 (N_975,In_263,In_78);
or U976 (N_976,In_2559,In_2431);
xnor U977 (N_977,In_2288,In_1670);
or U978 (N_978,In_756,In_439);
nor U979 (N_979,In_417,In_1667);
or U980 (N_980,In_994,In_2530);
or U981 (N_981,In_279,In_946);
and U982 (N_982,In_741,In_1631);
or U983 (N_983,In_2408,In_834);
nand U984 (N_984,In_1105,In_1461);
nor U985 (N_985,In_453,In_196);
nand U986 (N_986,In_299,In_2057);
and U987 (N_987,In_2124,In_190);
xnor U988 (N_988,In_1075,In_1287);
nor U989 (N_989,In_1410,In_2699);
and U990 (N_990,In_2924,In_27);
xnor U991 (N_991,In_1918,In_292);
and U992 (N_992,In_815,In_1786);
nor U993 (N_993,In_2461,In_2854);
nor U994 (N_994,In_2800,In_876);
nand U995 (N_995,In_980,In_2533);
nand U996 (N_996,In_2785,In_2809);
and U997 (N_997,In_528,In_150);
xnor U998 (N_998,In_655,In_2936);
nor U999 (N_999,In_2568,In_2757);
nor U1000 (N_1000,In_547,In_1968);
or U1001 (N_1001,In_2104,In_2516);
nand U1002 (N_1002,In_2964,In_1567);
and U1003 (N_1003,In_394,In_1423);
nor U1004 (N_1004,In_610,In_140);
or U1005 (N_1005,In_2918,In_665);
and U1006 (N_1006,In_458,In_1716);
or U1007 (N_1007,In_2356,In_1799);
or U1008 (N_1008,In_1848,In_2517);
and U1009 (N_1009,In_2960,In_1157);
nand U1010 (N_1010,In_2733,In_2626);
xnor U1011 (N_1011,In_1551,In_569);
xnor U1012 (N_1012,In_2750,In_602);
and U1013 (N_1013,In_1493,In_1407);
or U1014 (N_1014,In_1663,In_1885);
nor U1015 (N_1015,In_2011,In_1251);
and U1016 (N_1016,In_1496,In_44);
nand U1017 (N_1017,In_1525,In_2592);
nand U1018 (N_1018,In_2574,In_656);
xnor U1019 (N_1019,In_1281,In_2047);
and U1020 (N_1020,In_867,In_2166);
nand U1021 (N_1021,In_112,In_350);
nand U1022 (N_1022,In_425,In_2527);
and U1023 (N_1023,In_762,In_861);
nand U1024 (N_1024,In_159,In_901);
xor U1025 (N_1025,In_1787,In_2679);
and U1026 (N_1026,In_2588,In_2658);
and U1027 (N_1027,In_2157,In_1093);
and U1028 (N_1028,In_2086,In_84);
or U1029 (N_1029,In_1460,In_1822);
nand U1030 (N_1030,In_418,In_887);
xor U1031 (N_1031,In_509,In_203);
or U1032 (N_1032,In_1431,In_837);
xnor U1033 (N_1033,In_170,In_2044);
or U1034 (N_1034,In_886,In_317);
and U1035 (N_1035,In_2020,In_2148);
or U1036 (N_1036,In_1518,In_1932);
nor U1037 (N_1037,In_1552,In_751);
xor U1038 (N_1038,In_1253,In_1322);
nor U1039 (N_1039,In_2558,In_2231);
xor U1040 (N_1040,In_2767,In_1807);
xor U1041 (N_1041,In_1750,In_958);
and U1042 (N_1042,In_1425,In_2453);
xnor U1043 (N_1043,In_2042,In_1152);
nand U1044 (N_1044,In_1683,In_812);
nand U1045 (N_1045,In_1537,In_2227);
nor U1046 (N_1046,In_2038,In_2172);
nand U1047 (N_1047,In_326,In_1330);
and U1048 (N_1048,In_2815,In_1897);
nand U1049 (N_1049,In_288,In_307);
nor U1050 (N_1050,In_475,In_1743);
or U1051 (N_1051,In_2394,In_1976);
nand U1052 (N_1052,In_1834,In_339);
and U1053 (N_1053,In_2957,In_2518);
nor U1054 (N_1054,In_2033,In_118);
nor U1055 (N_1055,In_2159,In_114);
and U1056 (N_1056,In_68,In_848);
nor U1057 (N_1057,In_1998,In_948);
and U1058 (N_1058,In_2589,In_1576);
nand U1059 (N_1059,In_1417,In_2141);
nor U1060 (N_1060,In_2764,In_1387);
and U1061 (N_1061,In_151,In_2471);
nand U1062 (N_1062,In_1406,In_690);
nor U1063 (N_1063,In_1843,In_1585);
nand U1064 (N_1064,In_2498,In_421);
or U1065 (N_1065,In_617,In_1710);
nand U1066 (N_1066,In_882,In_593);
nor U1067 (N_1067,In_86,In_1562);
nor U1068 (N_1068,In_392,In_2778);
and U1069 (N_1069,In_2612,In_239);
and U1070 (N_1070,In_1520,In_549);
and U1071 (N_1071,In_253,In_334);
and U1072 (N_1072,In_437,In_195);
or U1073 (N_1073,In_2322,In_2171);
xnor U1074 (N_1074,In_933,In_457);
nand U1075 (N_1075,In_1705,In_338);
or U1076 (N_1076,In_2377,In_311);
nand U1077 (N_1077,In_776,In_1652);
or U1078 (N_1078,In_1526,In_89);
xnor U1079 (N_1079,In_218,In_2001);
xnor U1080 (N_1080,In_473,In_2318);
or U1081 (N_1081,In_926,In_2186);
and U1082 (N_1082,In_1633,In_494);
nand U1083 (N_1083,In_780,In_2551);
or U1084 (N_1084,In_2142,In_2661);
nor U1085 (N_1085,In_324,In_2061);
xnor U1086 (N_1086,In_1993,In_309);
nand U1087 (N_1087,In_1817,In_1381);
or U1088 (N_1088,In_2911,In_1684);
xnor U1089 (N_1089,In_2153,In_2866);
nor U1090 (N_1090,In_2252,In_544);
or U1091 (N_1091,In_554,In_2606);
or U1092 (N_1092,In_1405,In_2903);
or U1093 (N_1093,In_1501,In_4);
nand U1094 (N_1094,In_2916,In_2232);
and U1095 (N_1095,In_658,In_259);
nor U1096 (N_1096,In_2264,In_2731);
nand U1097 (N_1097,In_1118,In_2005);
or U1098 (N_1098,In_1744,In_841);
or U1099 (N_1099,In_388,In_1881);
or U1100 (N_1100,In_2724,In_1453);
nor U1101 (N_1101,In_2688,In_568);
and U1102 (N_1102,In_2657,In_328);
xor U1103 (N_1103,In_2334,In_2239);
nor U1104 (N_1104,In_802,In_245);
nand U1105 (N_1105,In_2353,In_2164);
xnor U1106 (N_1106,In_2901,In_1896);
nand U1107 (N_1107,In_1645,In_809);
and U1108 (N_1108,In_2179,In_2864);
or U1109 (N_1109,In_73,In_2206);
or U1110 (N_1110,In_1430,In_2545);
nor U1111 (N_1111,In_603,In_1739);
xnor U1112 (N_1112,In_660,In_1073);
nor U1113 (N_1113,In_1523,In_1476);
nand U1114 (N_1114,In_1299,In_1503);
nand U1115 (N_1115,In_1983,In_2732);
nand U1116 (N_1116,In_1766,In_1624);
nand U1117 (N_1117,In_2982,In_1803);
xnor U1118 (N_1118,In_667,In_1987);
or U1119 (N_1119,In_316,In_726);
xnor U1120 (N_1120,In_2217,In_606);
or U1121 (N_1121,In_1195,In_2185);
xor U1122 (N_1122,In_2618,In_456);
and U1123 (N_1123,In_595,In_2665);
and U1124 (N_1124,In_2686,In_734);
nand U1125 (N_1125,In_1934,In_2373);
or U1126 (N_1126,In_995,In_2249);
nor U1127 (N_1127,In_1618,In_1314);
nor U1128 (N_1128,In_359,In_2826);
and U1129 (N_1129,In_2111,In_693);
xor U1130 (N_1130,In_1895,In_2594);
and U1131 (N_1131,In_2432,In_2107);
nand U1132 (N_1132,In_2246,In_1183);
xnor U1133 (N_1133,In_1011,In_2905);
xor U1134 (N_1134,In_287,In_1818);
and U1135 (N_1135,In_1255,In_1841);
xnor U1136 (N_1136,In_2721,In_277);
xnor U1137 (N_1137,In_618,In_1789);
nor U1138 (N_1138,In_854,In_791);
nor U1139 (N_1139,In_1061,In_429);
nand U1140 (N_1140,In_2355,In_2028);
nand U1141 (N_1141,In_2423,In_777);
or U1142 (N_1142,In_1730,In_1083);
and U1143 (N_1143,In_639,In_1220);
nor U1144 (N_1144,In_176,In_2346);
nor U1145 (N_1145,In_2098,In_2765);
or U1146 (N_1146,In_936,In_601);
or U1147 (N_1147,In_58,In_1936);
xnor U1148 (N_1148,In_2191,In_143);
nor U1149 (N_1149,In_1639,In_571);
or U1150 (N_1150,In_1767,In_2613);
nor U1151 (N_1151,In_1737,In_2200);
and U1152 (N_1152,In_2881,In_585);
and U1153 (N_1153,In_827,In_1610);
and U1154 (N_1154,In_485,In_2321);
nor U1155 (N_1155,In_792,In_1891);
nor U1156 (N_1156,In_144,In_2849);
xor U1157 (N_1157,In_2628,In_925);
nor U1158 (N_1158,In_1199,In_451);
xnor U1159 (N_1159,In_1868,In_1202);
and U1160 (N_1160,In_1850,In_2391);
or U1161 (N_1161,In_2354,In_915);
nor U1162 (N_1162,In_1106,In_372);
xor U1163 (N_1163,In_1391,In_2904);
xor U1164 (N_1164,In_2382,In_1788);
xnor U1165 (N_1165,In_219,In_1893);
xnor U1166 (N_1166,In_247,In_2226);
and U1167 (N_1167,In_2875,In_1038);
xor U1168 (N_1168,In_1774,In_516);
nor U1169 (N_1169,In_2599,In_2726);
xor U1170 (N_1170,In_2280,In_222);
nor U1171 (N_1171,In_1673,In_1375);
nor U1172 (N_1172,In_1723,In_1347);
and U1173 (N_1173,In_2998,In_2065);
and U1174 (N_1174,In_2003,In_1409);
nand U1175 (N_1175,In_2298,In_953);
nor U1176 (N_1176,In_1021,In_2671);
or U1177 (N_1177,In_1863,In_1488);
nand U1178 (N_1178,In_1463,In_2714);
or U1179 (N_1179,In_353,In_2820);
and U1180 (N_1180,In_1139,In_1495);
or U1181 (N_1181,In_262,In_2090);
xnor U1182 (N_1182,In_1910,In_1698);
nand U1183 (N_1183,In_184,In_2308);
nor U1184 (N_1184,In_1902,In_2398);
nand U1185 (N_1185,In_2971,In_1751);
xor U1186 (N_1186,In_2895,In_2770);
xor U1187 (N_1187,In_2507,In_2277);
nor U1188 (N_1188,In_1449,In_254);
nor U1189 (N_1189,In_1081,In_1707);
nor U1190 (N_1190,In_2079,In_115);
xor U1191 (N_1191,In_1146,In_2146);
nand U1192 (N_1192,In_2531,In_1722);
or U1193 (N_1193,In_624,In_419);
or U1194 (N_1194,In_916,In_37);
or U1195 (N_1195,In_2873,In_224);
xor U1196 (N_1196,In_1225,In_202);
nand U1197 (N_1197,In_1242,In_1869);
and U1198 (N_1198,In_2010,In_336);
nor U1199 (N_1199,In_2290,In_2742);
nand U1200 (N_1200,In_558,In_2201);
xor U1201 (N_1201,In_826,In_2634);
and U1202 (N_1202,In_1901,In_1396);
xnor U1203 (N_1203,In_2949,In_2581);
nor U1204 (N_1204,In_2446,In_712);
nand U1205 (N_1205,In_127,In_1972);
nand U1206 (N_1206,In_389,In_80);
and U1207 (N_1207,In_256,In_1728);
or U1208 (N_1208,In_959,In_477);
nor U1209 (N_1209,In_761,In_1207);
nand U1210 (N_1210,In_766,In_2434);
nand U1211 (N_1211,In_775,In_432);
nor U1212 (N_1212,In_2056,In_395);
nor U1213 (N_1213,In_729,In_407);
and U1214 (N_1214,In_2170,In_1398);
nor U1215 (N_1215,In_2508,In_2367);
or U1216 (N_1216,In_1519,In_1655);
or U1217 (N_1217,In_768,In_2144);
xor U1218 (N_1218,In_1247,In_2887);
nand U1219 (N_1219,In_2414,In_1630);
and U1220 (N_1220,In_349,In_1418);
and U1221 (N_1221,In_2193,In_670);
xor U1222 (N_1222,In_2156,In_1419);
nand U1223 (N_1223,In_2897,In_1232);
nor U1224 (N_1224,In_1547,In_868);
nor U1225 (N_1225,In_1578,In_2372);
nand U1226 (N_1226,In_2376,In_2602);
and U1227 (N_1227,In_2593,In_1783);
nor U1228 (N_1228,In_1085,In_214);
nand U1229 (N_1229,In_619,In_413);
and U1230 (N_1230,In_1849,In_70);
nor U1231 (N_1231,In_830,In_2783);
or U1232 (N_1232,In_376,In_318);
or U1233 (N_1233,In_2287,In_914);
or U1234 (N_1234,In_2797,In_511);
and U1235 (N_1235,In_2419,In_1210);
xor U1236 (N_1236,In_275,In_1376);
or U1237 (N_1237,In_2975,In_1434);
nor U1238 (N_1238,In_1809,In_117);
and U1239 (N_1239,In_1682,In_1649);
xnor U1240 (N_1240,In_1088,In_2862);
xor U1241 (N_1241,In_835,In_1143);
and U1242 (N_1242,In_1478,In_1346);
and U1243 (N_1243,In_2333,In_2359);
or U1244 (N_1244,In_576,In_596);
xnor U1245 (N_1245,In_1374,In_428);
or U1246 (N_1246,In_2401,In_2442);
nor U1247 (N_1247,In_385,In_2638);
or U1248 (N_1248,In_468,In_2575);
nor U1249 (N_1249,In_1032,In_1086);
xnor U1250 (N_1250,In_1058,In_1690);
nand U1251 (N_1251,In_2980,In_1049);
xnor U1252 (N_1252,In_2463,In_2892);
or U1253 (N_1253,In_2371,In_1856);
nand U1254 (N_1254,In_2188,In_2748);
or U1255 (N_1255,In_2119,In_41);
or U1256 (N_1256,In_2043,In_698);
nand U1257 (N_1257,In_2630,In_733);
xnor U1258 (N_1258,In_1855,In_2933);
nor U1259 (N_1259,In_1236,In_1957);
and U1260 (N_1260,In_183,In_178);
or U1261 (N_1261,In_992,In_2886);
xor U1262 (N_1262,In_1756,In_240);
nor U1263 (N_1263,In_2266,In_1665);
nor U1264 (N_1264,In_76,In_1845);
nand U1265 (N_1265,In_90,In_2985);
xor U1266 (N_1266,In_1102,In_2580);
nor U1267 (N_1267,In_1366,In_1067);
and U1268 (N_1268,In_2898,In_2953);
nor U1269 (N_1269,In_1911,In_2907);
and U1270 (N_1270,In_2880,In_1001);
xor U1271 (N_1271,In_1996,In_1395);
nand U1272 (N_1272,In_567,In_717);
nor U1273 (N_1273,In_1666,In_1713);
or U1274 (N_1274,In_2080,In_36);
and U1275 (N_1275,In_2341,In_1876);
xor U1276 (N_1276,In_1960,In_2837);
and U1277 (N_1277,In_2459,In_74);
xnor U1278 (N_1278,In_991,In_727);
or U1279 (N_1279,In_40,In_1336);
xnor U1280 (N_1280,In_709,In_1945);
nand U1281 (N_1281,In_2669,In_1276);
xnor U1282 (N_1282,In_1883,In_1201);
or U1283 (N_1283,In_1780,In_1063);
and U1284 (N_1284,In_2863,In_1333);
nand U1285 (N_1285,In_2983,In_2829);
or U1286 (N_1286,In_1516,In_806);
xor U1287 (N_1287,In_77,In_1864);
or U1288 (N_1288,In_2387,In_836);
or U1289 (N_1289,In_1892,In_201);
xor U1290 (N_1290,In_855,In_2584);
nand U1291 (N_1291,In_2539,In_1858);
nor U1292 (N_1292,In_1249,In_2238);
nor U1293 (N_1293,In_448,In_701);
or U1294 (N_1294,In_2684,In_16);
xnor U1295 (N_1295,In_29,In_2350);
xnor U1296 (N_1296,In_2173,In_1971);
nor U1297 (N_1297,In_2672,In_1513);
nor U1298 (N_1298,In_412,In_2435);
or U1299 (N_1299,In_829,In_2868);
xor U1300 (N_1300,In_2860,In_2656);
xnor U1301 (N_1301,In_1340,In_957);
nor U1302 (N_1302,In_2122,In_1272);
nand U1303 (N_1303,In_2055,In_2366);
nor U1304 (N_1304,In_1473,In_512);
nand U1305 (N_1305,In_2158,In_2850);
nand U1306 (N_1306,In_25,In_2310);
and U1307 (N_1307,In_1607,In_2473);
nor U1308 (N_1308,In_1223,In_274);
and U1309 (N_1309,In_1318,In_306);
nand U1310 (N_1310,In_637,In_470);
nor U1311 (N_1311,In_2340,In_414);
nand U1312 (N_1312,In_2843,In_1637);
nand U1313 (N_1313,In_267,In_543);
nand U1314 (N_1314,In_1943,In_2948);
nor U1315 (N_1315,In_1828,In_12);
and U1316 (N_1316,In_582,In_189);
nor U1317 (N_1317,In_1888,In_110);
or U1318 (N_1318,In_647,In_1944);
nand U1319 (N_1319,In_2705,In_1660);
xnor U1320 (N_1320,In_863,In_2524);
nand U1321 (N_1321,In_821,In_2021);
xnor U1322 (N_1322,In_1754,In_1103);
and U1323 (N_1323,In_474,In_2012);
xnor U1324 (N_1324,In_2182,In_646);
and U1325 (N_1325,In_2175,In_1034);
xnor U1326 (N_1326,In_2694,In_1120);
nor U1327 (N_1327,In_2230,In_2085);
nand U1328 (N_1328,In_2420,In_1239);
xor U1329 (N_1329,In_1150,In_1529);
xor U1330 (N_1330,In_2803,In_480);
and U1331 (N_1331,In_1218,In_1853);
nand U1332 (N_1332,In_1792,In_1967);
xnor U1333 (N_1333,In_823,In_1274);
nor U1334 (N_1334,In_5,In_99);
nor U1335 (N_1335,In_1369,In_1466);
or U1336 (N_1336,In_1296,In_2470);
nor U1337 (N_1337,In_181,In_860);
nand U1338 (N_1338,In_911,In_2490);
and U1339 (N_1339,In_344,In_2591);
nand U1340 (N_1340,In_2919,In_393);
xor U1341 (N_1341,In_1161,In_714);
nand U1342 (N_1342,In_269,In_1005);
or U1343 (N_1343,In_2259,In_2513);
xnor U1344 (N_1344,In_2836,In_1471);
or U1345 (N_1345,In_2168,In_131);
nor U1346 (N_1346,In_47,In_772);
nand U1347 (N_1347,In_598,In_797);
xor U1348 (N_1348,In_1587,In_783);
or U1349 (N_1349,In_1160,In_2994);
nand U1350 (N_1350,In_2939,In_1836);
nand U1351 (N_1351,In_850,In_2947);
and U1352 (N_1352,In_208,In_478);
nor U1353 (N_1353,In_1414,In_69);
nand U1354 (N_1354,In_1219,In_2585);
nor U1355 (N_1355,In_816,In_1790);
or U1356 (N_1356,In_2834,In_2357);
and U1357 (N_1357,In_1217,In_1541);
xor U1358 (N_1358,In_998,In_1214);
and U1359 (N_1359,In_2944,In_692);
nand U1360 (N_1360,In_2506,In_1482);
and U1361 (N_1361,In_2218,In_1837);
and U1362 (N_1362,In_342,In_1712);
and U1363 (N_1363,In_3,In_556);
xor U1364 (N_1364,In_370,In_580);
and U1365 (N_1365,In_2292,In_2890);
nor U1366 (N_1366,In_1680,In_2358);
nand U1367 (N_1367,In_493,In_187);
nand U1368 (N_1368,In_1184,In_2561);
xnor U1369 (N_1369,In_103,In_1534);
and U1370 (N_1370,In_1765,In_1514);
xnor U1371 (N_1371,In_2791,In_2888);
nor U1372 (N_1372,In_673,In_1924);
nand U1373 (N_1373,In_1661,In_869);
xor U1374 (N_1374,In_2617,In_1582);
nand U1375 (N_1375,In_1262,In_764);
nor U1376 (N_1376,In_858,In_1696);
and U1377 (N_1377,In_972,In_31);
or U1378 (N_1378,In_904,In_538);
nand U1379 (N_1379,In_1358,In_1359);
and U1380 (N_1380,In_2587,In_290);
nand U1381 (N_1381,In_343,In_237);
xor U1382 (N_1382,In_2496,In_2793);
nand U1383 (N_1383,In_2769,In_1884);
and U1384 (N_1384,In_2967,In_650);
or U1385 (N_1385,In_2644,In_1721);
nor U1386 (N_1386,In_2710,In_163);
and U1387 (N_1387,In_1606,In_2970);
nor U1388 (N_1388,In_706,In_2388);
nor U1389 (N_1389,In_1091,In_401);
xnor U1390 (N_1390,In_1880,In_1009);
nor U1391 (N_1391,In_2772,In_1588);
and U1392 (N_1392,In_2870,In_1725);
nand U1393 (N_1393,In_2709,In_249);
nand U1394 (N_1394,In_844,In_1130);
or U1395 (N_1395,In_52,In_1194);
and U1396 (N_1396,In_1732,In_2910);
and U1397 (N_1397,In_1433,In_408);
and U1398 (N_1398,In_2489,In_641);
and U1399 (N_1399,In_98,In_1477);
nand U1400 (N_1400,In_1793,In_2780);
and U1401 (N_1401,In_2941,In_223);
or U1402 (N_1402,In_1203,In_1995);
and U1403 (N_1403,In_1922,In_323);
xor U1404 (N_1404,In_2032,In_2659);
and U1405 (N_1405,In_2125,In_455);
and U1406 (N_1406,In_2806,In_1474);
and U1407 (N_1407,In_374,In_640);
or U1408 (N_1408,In_2623,In_367);
and U1409 (N_1409,In_951,In_1357);
and U1410 (N_1410,In_2921,In_966);
xnor U1411 (N_1411,In_2364,In_168);
and U1412 (N_1412,In_1736,In_1215);
nor U1413 (N_1413,In_1439,In_9);
and U1414 (N_1414,In_1994,In_1186);
and U1415 (N_1415,In_1190,In_67);
nand U1416 (N_1416,In_1353,In_2380);
nand U1417 (N_1417,In_2092,In_1168);
nor U1418 (N_1418,In_501,In_50);
xnor U1419 (N_1419,In_2735,In_862);
nor U1420 (N_1420,In_431,In_1871);
xor U1421 (N_1421,In_351,In_22);
nand U1422 (N_1422,In_15,In_1907);
and U1423 (N_1423,In_1558,In_1540);
xor U1424 (N_1424,In_54,In_976);
and U1425 (N_1425,In_1467,In_1180);
nor U1426 (N_1426,In_2363,In_102);
and U1427 (N_1427,In_1584,In_212);
nand U1428 (N_1428,In_2332,In_1954);
nor U1429 (N_1429,In_1092,In_743);
and U1430 (N_1430,In_2035,In_2816);
nor U1431 (N_1431,In_2087,In_1919);
nand U1432 (N_1432,In_1999,In_2645);
nand U1433 (N_1433,In_466,In_2241);
and U1434 (N_1434,In_2000,In_731);
nand U1435 (N_1435,In_2761,In_581);
or U1436 (N_1436,In_2105,In_2676);
nor U1437 (N_1437,In_1411,In_795);
and U1438 (N_1438,In_1257,In_193);
or U1439 (N_1439,In_628,In_2485);
nor U1440 (N_1440,In_1538,In_711);
nor U1441 (N_1441,In_1413,In_940);
nor U1442 (N_1442,In_1781,In_2741);
or U1443 (N_1443,In_785,In_1940);
nand U1444 (N_1444,In_865,In_2966);
nand U1445 (N_1445,In_28,In_2106);
or U1446 (N_1446,In_1694,In_1755);
xor U1447 (N_1447,In_1345,In_75);
xnor U1448 (N_1448,In_2871,In_2563);
xor U1449 (N_1449,In_888,In_875);
nand U1450 (N_1450,In_1367,In_1459);
nor U1451 (N_1451,In_2309,In_2972);
and U1452 (N_1452,In_2272,In_2844);
or U1453 (N_1453,In_735,In_153);
nor U1454 (N_1454,In_2128,In_1758);
or U1455 (N_1455,In_1041,In_2428);
xor U1456 (N_1456,In_1373,In_1572);
nand U1457 (N_1457,In_2535,In_2213);
or U1458 (N_1458,In_1162,In_1164);
nand U1459 (N_1459,In_2802,In_2004);
xnor U1460 (N_1460,In_1642,In_8);
nor U1461 (N_1461,In_1378,In_2674);
nor U1462 (N_1462,In_1313,In_2729);
nor U1463 (N_1463,In_449,In_643);
or U1464 (N_1464,In_912,In_1872);
nor U1465 (N_1465,In_2418,In_2253);
nand U1466 (N_1466,In_2089,In_2293);
and U1467 (N_1467,In_1342,In_1577);
nand U1468 (N_1468,In_1422,In_148);
nand U1469 (N_1469,In_156,In_2685);
or U1470 (N_1470,In_2291,In_1820);
xnor U1471 (N_1471,In_489,In_443);
nand U1472 (N_1472,In_242,In_2692);
nand U1473 (N_1473,In_424,In_305);
or U1474 (N_1474,In_838,In_1456);
nand U1475 (N_1475,In_32,In_2221);
nand U1476 (N_1476,In_811,In_537);
or U1477 (N_1477,In_325,In_1412);
and U1478 (N_1478,In_1261,In_950);
nor U1479 (N_1479,In_2462,In_2279);
nand U1480 (N_1480,In_2483,In_2827);
and U1481 (N_1481,In_2025,In_204);
xor U1482 (N_1482,In_95,In_1319);
nor U1483 (N_1483,In_39,In_2385);
xnor U1484 (N_1484,In_1040,In_2763);
and U1485 (N_1485,In_2758,In_2273);
nor U1486 (N_1486,In_2294,In_1903);
xnor U1487 (N_1487,In_2565,In_1193);
xnor U1488 (N_1488,In_167,In_2502);
nand U1489 (N_1489,In_1556,In_303);
nand U1490 (N_1490,In_2361,In_2996);
and U1491 (N_1491,In_1740,In_1104);
xnor U1492 (N_1492,In_185,In_2555);
nor U1493 (N_1493,In_2317,In_1815);
nand U1494 (N_1494,In_321,In_2199);
xor U1495 (N_1495,In_2304,In_1636);
nand U1496 (N_1496,In_779,In_462);
nor U1497 (N_1497,In_55,In_500);
xor U1498 (N_1498,In_2712,In_533);
xnor U1499 (N_1499,In_1039,In_1401);
xnor U1500 (N_1500,In_2528,In_2903);
nor U1501 (N_1501,In_2717,In_2900);
nand U1502 (N_1502,In_1254,In_245);
or U1503 (N_1503,In_2481,In_315);
xor U1504 (N_1504,In_1597,In_2433);
xnor U1505 (N_1505,In_630,In_1053);
nand U1506 (N_1506,In_2663,In_2433);
and U1507 (N_1507,In_611,In_984);
nand U1508 (N_1508,In_332,In_2671);
or U1509 (N_1509,In_1154,In_404);
nand U1510 (N_1510,In_1623,In_1478);
nand U1511 (N_1511,In_1661,In_1973);
nor U1512 (N_1512,In_1397,In_2952);
nor U1513 (N_1513,In_528,In_2486);
and U1514 (N_1514,In_614,In_2136);
nand U1515 (N_1515,In_1392,In_879);
or U1516 (N_1516,In_2940,In_2086);
nand U1517 (N_1517,In_2835,In_1442);
xnor U1518 (N_1518,In_1521,In_2175);
nand U1519 (N_1519,In_2059,In_117);
nor U1520 (N_1520,In_1671,In_883);
nor U1521 (N_1521,In_1862,In_2480);
nor U1522 (N_1522,In_1571,In_1248);
xor U1523 (N_1523,In_1703,In_2107);
xnor U1524 (N_1524,In_33,In_1717);
nand U1525 (N_1525,In_1686,In_2588);
nor U1526 (N_1526,In_375,In_1545);
or U1527 (N_1527,In_2610,In_745);
nor U1528 (N_1528,In_1547,In_286);
nor U1529 (N_1529,In_716,In_2677);
nand U1530 (N_1530,In_1586,In_1614);
or U1531 (N_1531,In_1505,In_1602);
nand U1532 (N_1532,In_1417,In_1036);
nor U1533 (N_1533,In_489,In_2708);
and U1534 (N_1534,In_2367,In_994);
nor U1535 (N_1535,In_1328,In_708);
xnor U1536 (N_1536,In_2957,In_2042);
and U1537 (N_1537,In_130,In_1281);
or U1538 (N_1538,In_1679,In_1637);
or U1539 (N_1539,In_976,In_607);
nand U1540 (N_1540,In_394,In_2115);
nor U1541 (N_1541,In_2548,In_2340);
and U1542 (N_1542,In_2899,In_2728);
xnor U1543 (N_1543,In_2802,In_2847);
or U1544 (N_1544,In_791,In_511);
nand U1545 (N_1545,In_1269,In_741);
xnor U1546 (N_1546,In_864,In_349);
or U1547 (N_1547,In_696,In_541);
xnor U1548 (N_1548,In_1594,In_2689);
or U1549 (N_1549,In_689,In_2175);
nor U1550 (N_1550,In_1963,In_2877);
nand U1551 (N_1551,In_551,In_287);
and U1552 (N_1552,In_324,In_262);
nand U1553 (N_1553,In_1535,In_305);
xor U1554 (N_1554,In_1852,In_1559);
and U1555 (N_1555,In_2705,In_1923);
or U1556 (N_1556,In_356,In_392);
nand U1557 (N_1557,In_713,In_1124);
nand U1558 (N_1558,In_2435,In_929);
nand U1559 (N_1559,In_1795,In_1115);
xnor U1560 (N_1560,In_611,In_1499);
and U1561 (N_1561,In_1210,In_506);
nand U1562 (N_1562,In_1469,In_2092);
or U1563 (N_1563,In_2976,In_2302);
or U1564 (N_1564,In_317,In_1577);
nand U1565 (N_1565,In_2154,In_749);
xnor U1566 (N_1566,In_683,In_2874);
nor U1567 (N_1567,In_2299,In_501);
and U1568 (N_1568,In_2192,In_1747);
and U1569 (N_1569,In_557,In_1066);
or U1570 (N_1570,In_1205,In_2742);
or U1571 (N_1571,In_2635,In_2469);
or U1572 (N_1572,In_763,In_252);
nand U1573 (N_1573,In_1442,In_1780);
nor U1574 (N_1574,In_38,In_2287);
nand U1575 (N_1575,In_1785,In_2310);
or U1576 (N_1576,In_912,In_156);
xnor U1577 (N_1577,In_685,In_387);
nand U1578 (N_1578,In_535,In_1650);
and U1579 (N_1579,In_2539,In_1435);
and U1580 (N_1580,In_1888,In_1632);
and U1581 (N_1581,In_1622,In_2350);
nand U1582 (N_1582,In_1338,In_1191);
nor U1583 (N_1583,In_2414,In_1210);
and U1584 (N_1584,In_2671,In_1164);
and U1585 (N_1585,In_2134,In_1621);
and U1586 (N_1586,In_2313,In_255);
and U1587 (N_1587,In_2761,In_557);
xnor U1588 (N_1588,In_1489,In_466);
nor U1589 (N_1589,In_2740,In_2404);
and U1590 (N_1590,In_1993,In_1590);
and U1591 (N_1591,In_318,In_1899);
or U1592 (N_1592,In_2915,In_583);
nand U1593 (N_1593,In_1638,In_1760);
xnor U1594 (N_1594,In_2054,In_737);
nor U1595 (N_1595,In_1843,In_2083);
nand U1596 (N_1596,In_1639,In_532);
xnor U1597 (N_1597,In_524,In_1163);
nor U1598 (N_1598,In_2785,In_2331);
nand U1599 (N_1599,In_1458,In_864);
xnor U1600 (N_1600,In_60,In_588);
and U1601 (N_1601,In_2915,In_2871);
nand U1602 (N_1602,In_597,In_2362);
nand U1603 (N_1603,In_1332,In_1742);
nand U1604 (N_1604,In_368,In_2720);
or U1605 (N_1605,In_1394,In_2397);
nand U1606 (N_1606,In_1420,In_1407);
xor U1607 (N_1607,In_1044,In_769);
nor U1608 (N_1608,In_2059,In_979);
nand U1609 (N_1609,In_567,In_2286);
nor U1610 (N_1610,In_2461,In_2172);
and U1611 (N_1611,In_1475,In_2208);
nand U1612 (N_1612,In_1107,In_1702);
nor U1613 (N_1613,In_1892,In_249);
xor U1614 (N_1614,In_1613,In_1784);
and U1615 (N_1615,In_4,In_2902);
nor U1616 (N_1616,In_703,In_1211);
xnor U1617 (N_1617,In_290,In_951);
or U1618 (N_1618,In_2812,In_1242);
or U1619 (N_1619,In_800,In_836);
xor U1620 (N_1620,In_160,In_880);
and U1621 (N_1621,In_2522,In_2176);
or U1622 (N_1622,In_168,In_2360);
nor U1623 (N_1623,In_2636,In_930);
and U1624 (N_1624,In_811,In_804);
nor U1625 (N_1625,In_1780,In_2806);
and U1626 (N_1626,In_2318,In_908);
xnor U1627 (N_1627,In_647,In_339);
xor U1628 (N_1628,In_1202,In_1590);
xor U1629 (N_1629,In_1692,In_2399);
xnor U1630 (N_1630,In_154,In_758);
or U1631 (N_1631,In_1126,In_1800);
nand U1632 (N_1632,In_1550,In_472);
nand U1633 (N_1633,In_1991,In_795);
xor U1634 (N_1634,In_798,In_1763);
and U1635 (N_1635,In_2608,In_322);
nor U1636 (N_1636,In_2940,In_2233);
and U1637 (N_1637,In_1953,In_1134);
nand U1638 (N_1638,In_230,In_131);
xnor U1639 (N_1639,In_1686,In_590);
xor U1640 (N_1640,In_1666,In_725);
and U1641 (N_1641,In_402,In_1588);
nor U1642 (N_1642,In_2180,In_1130);
or U1643 (N_1643,In_2971,In_2951);
xor U1644 (N_1644,In_2121,In_27);
nor U1645 (N_1645,In_2295,In_2217);
and U1646 (N_1646,In_2056,In_2786);
and U1647 (N_1647,In_2511,In_293);
nor U1648 (N_1648,In_917,In_461);
or U1649 (N_1649,In_1704,In_472);
xnor U1650 (N_1650,In_2426,In_953);
nand U1651 (N_1651,In_2672,In_2495);
xor U1652 (N_1652,In_67,In_2513);
or U1653 (N_1653,In_2855,In_370);
nor U1654 (N_1654,In_607,In_123);
nor U1655 (N_1655,In_2787,In_2322);
or U1656 (N_1656,In_162,In_889);
or U1657 (N_1657,In_255,In_1647);
xnor U1658 (N_1658,In_441,In_521);
or U1659 (N_1659,In_1732,In_2479);
nor U1660 (N_1660,In_1282,In_458);
or U1661 (N_1661,In_1196,In_1015);
xnor U1662 (N_1662,In_2493,In_2476);
or U1663 (N_1663,In_624,In_2728);
xnor U1664 (N_1664,In_1085,In_983);
xor U1665 (N_1665,In_2325,In_2618);
nor U1666 (N_1666,In_2045,In_394);
nand U1667 (N_1667,In_1059,In_169);
nand U1668 (N_1668,In_1944,In_1492);
nand U1669 (N_1669,In_2678,In_449);
nor U1670 (N_1670,In_746,In_1633);
nand U1671 (N_1671,In_612,In_2416);
nand U1672 (N_1672,In_1264,In_1806);
nand U1673 (N_1673,In_551,In_2611);
and U1674 (N_1674,In_773,In_2159);
xor U1675 (N_1675,In_441,In_468);
and U1676 (N_1676,In_1705,In_1373);
nor U1677 (N_1677,In_514,In_2366);
or U1678 (N_1678,In_1815,In_293);
or U1679 (N_1679,In_2092,In_2607);
or U1680 (N_1680,In_1545,In_1997);
nand U1681 (N_1681,In_1949,In_679);
or U1682 (N_1682,In_8,In_482);
and U1683 (N_1683,In_109,In_1371);
xnor U1684 (N_1684,In_2645,In_1458);
nand U1685 (N_1685,In_2535,In_2061);
and U1686 (N_1686,In_2830,In_147);
xor U1687 (N_1687,In_1937,In_682);
nor U1688 (N_1688,In_1224,In_1637);
nor U1689 (N_1689,In_188,In_1227);
nand U1690 (N_1690,In_1931,In_137);
nand U1691 (N_1691,In_931,In_1188);
and U1692 (N_1692,In_2002,In_1559);
nand U1693 (N_1693,In_1479,In_2976);
nand U1694 (N_1694,In_2202,In_2702);
and U1695 (N_1695,In_1881,In_421);
nand U1696 (N_1696,In_1254,In_113);
nand U1697 (N_1697,In_2358,In_2522);
nand U1698 (N_1698,In_1745,In_2379);
or U1699 (N_1699,In_1768,In_2823);
and U1700 (N_1700,In_1387,In_1525);
or U1701 (N_1701,In_1728,In_2233);
nor U1702 (N_1702,In_819,In_442);
nand U1703 (N_1703,In_1409,In_2903);
nand U1704 (N_1704,In_873,In_1131);
or U1705 (N_1705,In_1169,In_2096);
nor U1706 (N_1706,In_2343,In_641);
xor U1707 (N_1707,In_2293,In_1857);
and U1708 (N_1708,In_2304,In_1869);
nor U1709 (N_1709,In_2207,In_804);
xor U1710 (N_1710,In_2017,In_1494);
nand U1711 (N_1711,In_2437,In_923);
nor U1712 (N_1712,In_2228,In_1285);
nor U1713 (N_1713,In_1213,In_690);
nand U1714 (N_1714,In_578,In_2424);
or U1715 (N_1715,In_2272,In_205);
or U1716 (N_1716,In_1933,In_1422);
nand U1717 (N_1717,In_2266,In_690);
and U1718 (N_1718,In_2505,In_853);
nor U1719 (N_1719,In_1689,In_1353);
nand U1720 (N_1720,In_1647,In_615);
and U1721 (N_1721,In_1524,In_2386);
xor U1722 (N_1722,In_51,In_670);
nand U1723 (N_1723,In_2048,In_2368);
xor U1724 (N_1724,In_253,In_2935);
or U1725 (N_1725,In_73,In_2780);
or U1726 (N_1726,In_984,In_44);
nor U1727 (N_1727,In_1288,In_2236);
xor U1728 (N_1728,In_1558,In_510);
and U1729 (N_1729,In_669,In_823);
or U1730 (N_1730,In_2362,In_876);
and U1731 (N_1731,In_2110,In_1688);
nor U1732 (N_1732,In_1004,In_2341);
xor U1733 (N_1733,In_913,In_1634);
or U1734 (N_1734,In_997,In_1680);
and U1735 (N_1735,In_2304,In_1555);
or U1736 (N_1736,In_2564,In_2249);
nor U1737 (N_1737,In_1107,In_295);
nand U1738 (N_1738,In_1804,In_1959);
or U1739 (N_1739,In_1626,In_2231);
and U1740 (N_1740,In_409,In_1000);
or U1741 (N_1741,In_1213,In_259);
nand U1742 (N_1742,In_2318,In_1240);
nand U1743 (N_1743,In_474,In_2698);
xnor U1744 (N_1744,In_3,In_893);
and U1745 (N_1745,In_1494,In_2802);
xor U1746 (N_1746,In_803,In_854);
nand U1747 (N_1747,In_2278,In_196);
or U1748 (N_1748,In_2357,In_1713);
nor U1749 (N_1749,In_1804,In_392);
nor U1750 (N_1750,In_1221,In_1481);
and U1751 (N_1751,In_1825,In_744);
and U1752 (N_1752,In_1351,In_1374);
xnor U1753 (N_1753,In_1307,In_968);
or U1754 (N_1754,In_875,In_2063);
nand U1755 (N_1755,In_1664,In_367);
nor U1756 (N_1756,In_1511,In_2778);
or U1757 (N_1757,In_2421,In_1699);
and U1758 (N_1758,In_2043,In_2799);
or U1759 (N_1759,In_1495,In_2142);
nor U1760 (N_1760,In_2788,In_1815);
nand U1761 (N_1761,In_1089,In_1025);
or U1762 (N_1762,In_1484,In_731);
xnor U1763 (N_1763,In_2062,In_226);
and U1764 (N_1764,In_1887,In_85);
nand U1765 (N_1765,In_617,In_1370);
or U1766 (N_1766,In_1234,In_2939);
nand U1767 (N_1767,In_1710,In_1539);
nor U1768 (N_1768,In_2944,In_2046);
nand U1769 (N_1769,In_2286,In_2104);
or U1770 (N_1770,In_1357,In_1127);
or U1771 (N_1771,In_398,In_1757);
xnor U1772 (N_1772,In_2055,In_1212);
or U1773 (N_1773,In_108,In_2199);
and U1774 (N_1774,In_2732,In_1672);
xor U1775 (N_1775,In_1752,In_2555);
and U1776 (N_1776,In_90,In_2042);
and U1777 (N_1777,In_2685,In_1672);
and U1778 (N_1778,In_2004,In_1793);
nor U1779 (N_1779,In_1428,In_2048);
xor U1780 (N_1780,In_374,In_2813);
nor U1781 (N_1781,In_1741,In_2164);
and U1782 (N_1782,In_1819,In_2093);
or U1783 (N_1783,In_2806,In_2638);
xnor U1784 (N_1784,In_1470,In_16);
and U1785 (N_1785,In_637,In_2428);
and U1786 (N_1786,In_478,In_2946);
xnor U1787 (N_1787,In_862,In_2473);
and U1788 (N_1788,In_1297,In_243);
and U1789 (N_1789,In_2608,In_101);
nand U1790 (N_1790,In_1879,In_131);
xnor U1791 (N_1791,In_34,In_1247);
nand U1792 (N_1792,In_1831,In_901);
nand U1793 (N_1793,In_2602,In_1403);
and U1794 (N_1794,In_1764,In_732);
nand U1795 (N_1795,In_390,In_1627);
nand U1796 (N_1796,In_1191,In_2538);
xnor U1797 (N_1797,In_2171,In_1366);
and U1798 (N_1798,In_1514,In_1773);
xnor U1799 (N_1799,In_1437,In_664);
nor U1800 (N_1800,In_892,In_1698);
nor U1801 (N_1801,In_2122,In_775);
or U1802 (N_1802,In_2649,In_139);
nand U1803 (N_1803,In_1105,In_1222);
or U1804 (N_1804,In_1005,In_1973);
and U1805 (N_1805,In_2983,In_671);
and U1806 (N_1806,In_1358,In_187);
nor U1807 (N_1807,In_64,In_1776);
nor U1808 (N_1808,In_2841,In_2517);
or U1809 (N_1809,In_2630,In_1036);
or U1810 (N_1810,In_2582,In_1570);
or U1811 (N_1811,In_739,In_2117);
nand U1812 (N_1812,In_1407,In_2279);
and U1813 (N_1813,In_2298,In_74);
nor U1814 (N_1814,In_788,In_2498);
nor U1815 (N_1815,In_2822,In_903);
and U1816 (N_1816,In_494,In_1272);
and U1817 (N_1817,In_155,In_2116);
nor U1818 (N_1818,In_1961,In_2821);
or U1819 (N_1819,In_147,In_2919);
or U1820 (N_1820,In_1464,In_652);
or U1821 (N_1821,In_2989,In_783);
nand U1822 (N_1822,In_1846,In_716);
and U1823 (N_1823,In_2139,In_1963);
and U1824 (N_1824,In_1106,In_1703);
xnor U1825 (N_1825,In_1963,In_1716);
and U1826 (N_1826,In_457,In_2136);
nor U1827 (N_1827,In_528,In_1232);
nand U1828 (N_1828,In_655,In_1784);
nand U1829 (N_1829,In_1673,In_2466);
xnor U1830 (N_1830,In_2236,In_2328);
nor U1831 (N_1831,In_204,In_176);
nand U1832 (N_1832,In_970,In_2902);
nor U1833 (N_1833,In_2727,In_2150);
nand U1834 (N_1834,In_2095,In_2466);
nand U1835 (N_1835,In_2046,In_2487);
nor U1836 (N_1836,In_658,In_233);
xor U1837 (N_1837,In_2755,In_1366);
or U1838 (N_1838,In_2149,In_2539);
xnor U1839 (N_1839,In_909,In_1677);
nand U1840 (N_1840,In_555,In_2966);
and U1841 (N_1841,In_2932,In_1973);
nor U1842 (N_1842,In_2799,In_1872);
or U1843 (N_1843,In_954,In_940);
and U1844 (N_1844,In_480,In_1635);
or U1845 (N_1845,In_1543,In_1955);
and U1846 (N_1846,In_399,In_2226);
or U1847 (N_1847,In_1388,In_1908);
and U1848 (N_1848,In_227,In_954);
xnor U1849 (N_1849,In_2667,In_817);
nor U1850 (N_1850,In_1741,In_1494);
nor U1851 (N_1851,In_1811,In_1078);
nor U1852 (N_1852,In_1829,In_567);
nor U1853 (N_1853,In_187,In_1288);
xnor U1854 (N_1854,In_2751,In_1427);
or U1855 (N_1855,In_2704,In_749);
or U1856 (N_1856,In_357,In_1343);
or U1857 (N_1857,In_2675,In_1468);
and U1858 (N_1858,In_569,In_100);
or U1859 (N_1859,In_1255,In_2766);
or U1860 (N_1860,In_2552,In_1011);
nor U1861 (N_1861,In_1601,In_2312);
nand U1862 (N_1862,In_1631,In_1135);
nand U1863 (N_1863,In_940,In_1468);
and U1864 (N_1864,In_2718,In_284);
xnor U1865 (N_1865,In_698,In_1719);
xor U1866 (N_1866,In_909,In_1590);
nand U1867 (N_1867,In_2710,In_1011);
nor U1868 (N_1868,In_2950,In_2844);
or U1869 (N_1869,In_374,In_740);
and U1870 (N_1870,In_507,In_1473);
nand U1871 (N_1871,In_1305,In_1777);
and U1872 (N_1872,In_593,In_989);
nor U1873 (N_1873,In_1524,In_629);
nor U1874 (N_1874,In_2372,In_2906);
nand U1875 (N_1875,In_2782,In_1446);
and U1876 (N_1876,In_1754,In_436);
or U1877 (N_1877,In_747,In_859);
xnor U1878 (N_1878,In_807,In_2033);
or U1879 (N_1879,In_2525,In_1725);
xor U1880 (N_1880,In_672,In_2614);
xnor U1881 (N_1881,In_2561,In_474);
and U1882 (N_1882,In_149,In_2128);
nor U1883 (N_1883,In_1639,In_2387);
xnor U1884 (N_1884,In_1701,In_1427);
xnor U1885 (N_1885,In_1176,In_2727);
xor U1886 (N_1886,In_919,In_2809);
or U1887 (N_1887,In_1555,In_2634);
xor U1888 (N_1888,In_2309,In_1679);
or U1889 (N_1889,In_2632,In_887);
nand U1890 (N_1890,In_2517,In_1759);
and U1891 (N_1891,In_1207,In_1025);
and U1892 (N_1892,In_1689,In_1844);
nand U1893 (N_1893,In_1368,In_2459);
nand U1894 (N_1894,In_294,In_1888);
nor U1895 (N_1895,In_2267,In_1050);
and U1896 (N_1896,In_81,In_817);
or U1897 (N_1897,In_1799,In_2502);
xor U1898 (N_1898,In_2356,In_2162);
and U1899 (N_1899,In_2957,In_1089);
nor U1900 (N_1900,In_1097,In_129);
nor U1901 (N_1901,In_2460,In_1580);
or U1902 (N_1902,In_1955,In_1826);
nand U1903 (N_1903,In_2067,In_2639);
nor U1904 (N_1904,In_304,In_2113);
nand U1905 (N_1905,In_1641,In_1036);
and U1906 (N_1906,In_2386,In_2043);
nand U1907 (N_1907,In_1806,In_226);
nand U1908 (N_1908,In_2973,In_1416);
xor U1909 (N_1909,In_680,In_450);
and U1910 (N_1910,In_2836,In_2509);
xnor U1911 (N_1911,In_1138,In_381);
nor U1912 (N_1912,In_298,In_236);
nor U1913 (N_1913,In_2720,In_1259);
nand U1914 (N_1914,In_2328,In_2307);
nor U1915 (N_1915,In_2135,In_1123);
nand U1916 (N_1916,In_2750,In_344);
and U1917 (N_1917,In_2284,In_2715);
nor U1918 (N_1918,In_1810,In_1281);
or U1919 (N_1919,In_1998,In_1304);
and U1920 (N_1920,In_2189,In_428);
and U1921 (N_1921,In_2655,In_220);
xnor U1922 (N_1922,In_1938,In_1508);
nor U1923 (N_1923,In_542,In_2377);
nor U1924 (N_1924,In_1638,In_2940);
nor U1925 (N_1925,In_2954,In_1485);
and U1926 (N_1926,In_2220,In_1884);
nand U1927 (N_1927,In_858,In_716);
and U1928 (N_1928,In_244,In_1527);
nand U1929 (N_1929,In_894,In_2922);
and U1930 (N_1930,In_2991,In_1138);
or U1931 (N_1931,In_2460,In_2964);
nand U1932 (N_1932,In_2313,In_472);
and U1933 (N_1933,In_2698,In_1134);
or U1934 (N_1934,In_827,In_2234);
or U1935 (N_1935,In_2216,In_621);
nand U1936 (N_1936,In_2947,In_2531);
and U1937 (N_1937,In_2067,In_2452);
nand U1938 (N_1938,In_2977,In_2783);
xnor U1939 (N_1939,In_112,In_1234);
nor U1940 (N_1940,In_2686,In_1185);
xor U1941 (N_1941,In_1465,In_844);
or U1942 (N_1942,In_1148,In_174);
nor U1943 (N_1943,In_2004,In_2637);
xnor U1944 (N_1944,In_1479,In_2118);
xnor U1945 (N_1945,In_1187,In_1476);
and U1946 (N_1946,In_2488,In_997);
nor U1947 (N_1947,In_475,In_826);
and U1948 (N_1948,In_1383,In_1344);
and U1949 (N_1949,In_1215,In_2009);
xor U1950 (N_1950,In_2836,In_684);
nand U1951 (N_1951,In_2237,In_2376);
or U1952 (N_1952,In_583,In_2141);
xor U1953 (N_1953,In_1143,In_2784);
and U1954 (N_1954,In_2490,In_1824);
or U1955 (N_1955,In_2170,In_2977);
nor U1956 (N_1956,In_690,In_1128);
nand U1957 (N_1957,In_2747,In_2061);
nor U1958 (N_1958,In_1856,In_208);
or U1959 (N_1959,In_468,In_1787);
xor U1960 (N_1960,In_1840,In_1208);
nor U1961 (N_1961,In_902,In_1560);
xor U1962 (N_1962,In_1674,In_456);
xor U1963 (N_1963,In_2762,In_1898);
xor U1964 (N_1964,In_1000,In_1339);
or U1965 (N_1965,In_2183,In_2234);
xnor U1966 (N_1966,In_4,In_2484);
xnor U1967 (N_1967,In_352,In_2925);
and U1968 (N_1968,In_1568,In_927);
and U1969 (N_1969,In_1715,In_7);
and U1970 (N_1970,In_978,In_2891);
xnor U1971 (N_1971,In_1417,In_2810);
nor U1972 (N_1972,In_2017,In_461);
or U1973 (N_1973,In_2402,In_670);
or U1974 (N_1974,In_2060,In_1036);
or U1975 (N_1975,In_522,In_2124);
xor U1976 (N_1976,In_1860,In_13);
nand U1977 (N_1977,In_577,In_728);
xnor U1978 (N_1978,In_2872,In_557);
and U1979 (N_1979,In_1963,In_1223);
nor U1980 (N_1980,In_2207,In_2005);
xor U1981 (N_1981,In_978,In_1071);
xor U1982 (N_1982,In_2062,In_552);
xor U1983 (N_1983,In_2541,In_1836);
or U1984 (N_1984,In_2000,In_328);
and U1985 (N_1985,In_625,In_753);
nor U1986 (N_1986,In_2553,In_2720);
xor U1987 (N_1987,In_914,In_2860);
nor U1988 (N_1988,In_2784,In_2841);
or U1989 (N_1989,In_1167,In_2279);
or U1990 (N_1990,In_2793,In_1942);
or U1991 (N_1991,In_1876,In_1074);
or U1992 (N_1992,In_471,In_827);
or U1993 (N_1993,In_2651,In_26);
or U1994 (N_1994,In_2141,In_991);
nand U1995 (N_1995,In_610,In_2986);
nand U1996 (N_1996,In_2696,In_2908);
nand U1997 (N_1997,In_1046,In_2638);
or U1998 (N_1998,In_2235,In_589);
or U1999 (N_1999,In_704,In_1786);
or U2000 (N_2000,In_2814,In_2076);
nand U2001 (N_2001,In_171,In_547);
nor U2002 (N_2002,In_1314,In_1533);
nor U2003 (N_2003,In_732,In_350);
nand U2004 (N_2004,In_2502,In_763);
and U2005 (N_2005,In_1036,In_2637);
and U2006 (N_2006,In_836,In_1288);
and U2007 (N_2007,In_1300,In_2010);
and U2008 (N_2008,In_2364,In_232);
and U2009 (N_2009,In_1568,In_1208);
and U2010 (N_2010,In_841,In_2540);
xor U2011 (N_2011,In_146,In_1834);
nand U2012 (N_2012,In_607,In_447);
nor U2013 (N_2013,In_1623,In_1666);
nand U2014 (N_2014,In_1984,In_2062);
and U2015 (N_2015,In_2145,In_2896);
xor U2016 (N_2016,In_1530,In_2662);
or U2017 (N_2017,In_136,In_2065);
nor U2018 (N_2018,In_1633,In_1640);
nor U2019 (N_2019,In_2532,In_243);
and U2020 (N_2020,In_1062,In_1362);
nand U2021 (N_2021,In_2022,In_1674);
or U2022 (N_2022,In_372,In_359);
nand U2023 (N_2023,In_622,In_2367);
nand U2024 (N_2024,In_2066,In_2704);
nor U2025 (N_2025,In_1164,In_1582);
nor U2026 (N_2026,In_2320,In_2804);
and U2027 (N_2027,In_425,In_2423);
nand U2028 (N_2028,In_2719,In_2475);
or U2029 (N_2029,In_606,In_689);
nand U2030 (N_2030,In_498,In_1542);
and U2031 (N_2031,In_1043,In_1343);
nor U2032 (N_2032,In_1893,In_2049);
or U2033 (N_2033,In_96,In_812);
and U2034 (N_2034,In_884,In_1807);
or U2035 (N_2035,In_835,In_2685);
or U2036 (N_2036,In_1080,In_2413);
xor U2037 (N_2037,In_21,In_2406);
nand U2038 (N_2038,In_512,In_719);
xor U2039 (N_2039,In_1051,In_2520);
xnor U2040 (N_2040,In_1740,In_1820);
nand U2041 (N_2041,In_149,In_346);
xor U2042 (N_2042,In_151,In_1836);
nor U2043 (N_2043,In_237,In_1713);
nor U2044 (N_2044,In_2117,In_1835);
xor U2045 (N_2045,In_2306,In_1015);
xor U2046 (N_2046,In_1314,In_1008);
nor U2047 (N_2047,In_2537,In_983);
nor U2048 (N_2048,In_1515,In_2851);
and U2049 (N_2049,In_2062,In_1853);
and U2050 (N_2050,In_1423,In_2335);
and U2051 (N_2051,In_476,In_938);
and U2052 (N_2052,In_2523,In_1120);
and U2053 (N_2053,In_1990,In_649);
and U2054 (N_2054,In_1243,In_658);
xnor U2055 (N_2055,In_1840,In_1058);
nor U2056 (N_2056,In_884,In_895);
or U2057 (N_2057,In_738,In_1752);
xnor U2058 (N_2058,In_476,In_679);
nor U2059 (N_2059,In_2016,In_361);
and U2060 (N_2060,In_1121,In_1256);
xor U2061 (N_2061,In_2277,In_1103);
xor U2062 (N_2062,In_2086,In_453);
xnor U2063 (N_2063,In_145,In_2802);
and U2064 (N_2064,In_952,In_2131);
nand U2065 (N_2065,In_1956,In_2670);
and U2066 (N_2066,In_1567,In_47);
xnor U2067 (N_2067,In_790,In_658);
nor U2068 (N_2068,In_165,In_280);
and U2069 (N_2069,In_28,In_2269);
or U2070 (N_2070,In_1006,In_2749);
and U2071 (N_2071,In_1488,In_2586);
or U2072 (N_2072,In_1622,In_1992);
and U2073 (N_2073,In_2095,In_2090);
and U2074 (N_2074,In_547,In_1283);
or U2075 (N_2075,In_1862,In_636);
xor U2076 (N_2076,In_341,In_1695);
xnor U2077 (N_2077,In_760,In_1185);
xnor U2078 (N_2078,In_880,In_1359);
or U2079 (N_2079,In_1380,In_236);
or U2080 (N_2080,In_2932,In_2965);
nand U2081 (N_2081,In_667,In_2496);
nor U2082 (N_2082,In_696,In_2148);
or U2083 (N_2083,In_2047,In_947);
or U2084 (N_2084,In_1380,In_471);
xor U2085 (N_2085,In_1665,In_2441);
or U2086 (N_2086,In_786,In_2804);
and U2087 (N_2087,In_1067,In_561);
or U2088 (N_2088,In_2422,In_803);
nor U2089 (N_2089,In_1954,In_682);
nor U2090 (N_2090,In_1380,In_1553);
or U2091 (N_2091,In_2549,In_2983);
nor U2092 (N_2092,In_2718,In_2231);
and U2093 (N_2093,In_1873,In_2341);
and U2094 (N_2094,In_2391,In_2180);
and U2095 (N_2095,In_1863,In_250);
and U2096 (N_2096,In_475,In_1284);
xor U2097 (N_2097,In_167,In_2595);
nor U2098 (N_2098,In_1813,In_33);
or U2099 (N_2099,In_342,In_2437);
xor U2100 (N_2100,In_2878,In_291);
or U2101 (N_2101,In_1524,In_1627);
nor U2102 (N_2102,In_1553,In_228);
nand U2103 (N_2103,In_2556,In_2037);
and U2104 (N_2104,In_2697,In_351);
and U2105 (N_2105,In_2527,In_1920);
nor U2106 (N_2106,In_425,In_341);
and U2107 (N_2107,In_2639,In_2419);
xnor U2108 (N_2108,In_2084,In_1305);
nor U2109 (N_2109,In_2863,In_2325);
nor U2110 (N_2110,In_2990,In_1343);
nand U2111 (N_2111,In_270,In_2553);
or U2112 (N_2112,In_203,In_2734);
nand U2113 (N_2113,In_2545,In_1630);
xor U2114 (N_2114,In_2524,In_2267);
and U2115 (N_2115,In_834,In_2021);
and U2116 (N_2116,In_1805,In_1963);
nor U2117 (N_2117,In_764,In_2696);
xnor U2118 (N_2118,In_1879,In_2290);
or U2119 (N_2119,In_1809,In_536);
nor U2120 (N_2120,In_196,In_527);
or U2121 (N_2121,In_2116,In_1202);
and U2122 (N_2122,In_469,In_1450);
and U2123 (N_2123,In_2965,In_2545);
nand U2124 (N_2124,In_2099,In_1805);
xor U2125 (N_2125,In_1280,In_131);
and U2126 (N_2126,In_2058,In_2512);
xnor U2127 (N_2127,In_934,In_1566);
and U2128 (N_2128,In_1525,In_2862);
or U2129 (N_2129,In_1866,In_1414);
nand U2130 (N_2130,In_1379,In_2265);
and U2131 (N_2131,In_809,In_2459);
nand U2132 (N_2132,In_2158,In_2460);
and U2133 (N_2133,In_32,In_330);
xnor U2134 (N_2134,In_396,In_1592);
xnor U2135 (N_2135,In_430,In_287);
nand U2136 (N_2136,In_2339,In_695);
or U2137 (N_2137,In_694,In_1944);
nand U2138 (N_2138,In_1245,In_2384);
and U2139 (N_2139,In_928,In_2290);
nand U2140 (N_2140,In_1292,In_1188);
nand U2141 (N_2141,In_2159,In_1258);
and U2142 (N_2142,In_2397,In_662);
and U2143 (N_2143,In_1312,In_2277);
and U2144 (N_2144,In_1513,In_893);
nor U2145 (N_2145,In_188,In_5);
or U2146 (N_2146,In_2822,In_1837);
or U2147 (N_2147,In_2087,In_1436);
nor U2148 (N_2148,In_1945,In_1347);
nor U2149 (N_2149,In_996,In_1053);
nor U2150 (N_2150,In_85,In_1745);
xor U2151 (N_2151,In_2442,In_1006);
and U2152 (N_2152,In_95,In_2059);
or U2153 (N_2153,In_2148,In_186);
nor U2154 (N_2154,In_34,In_1088);
and U2155 (N_2155,In_1137,In_867);
xor U2156 (N_2156,In_2244,In_1604);
or U2157 (N_2157,In_2624,In_772);
xor U2158 (N_2158,In_467,In_423);
nand U2159 (N_2159,In_2902,In_2102);
and U2160 (N_2160,In_1489,In_1166);
and U2161 (N_2161,In_583,In_597);
nor U2162 (N_2162,In_2542,In_1620);
and U2163 (N_2163,In_2631,In_2119);
and U2164 (N_2164,In_258,In_2048);
nand U2165 (N_2165,In_2495,In_1393);
nor U2166 (N_2166,In_1904,In_124);
nor U2167 (N_2167,In_2679,In_1825);
nand U2168 (N_2168,In_1605,In_2422);
xnor U2169 (N_2169,In_2190,In_104);
nand U2170 (N_2170,In_1722,In_2711);
xnor U2171 (N_2171,In_1890,In_2464);
xor U2172 (N_2172,In_1043,In_64);
and U2173 (N_2173,In_1625,In_593);
nor U2174 (N_2174,In_323,In_1703);
nor U2175 (N_2175,In_1841,In_2123);
nand U2176 (N_2176,In_1703,In_856);
nand U2177 (N_2177,In_1143,In_1330);
nor U2178 (N_2178,In_2684,In_692);
nor U2179 (N_2179,In_781,In_190);
nand U2180 (N_2180,In_1887,In_488);
xnor U2181 (N_2181,In_2001,In_2795);
or U2182 (N_2182,In_774,In_1305);
nor U2183 (N_2183,In_1914,In_562);
and U2184 (N_2184,In_630,In_738);
nand U2185 (N_2185,In_441,In_45);
and U2186 (N_2186,In_2637,In_2499);
nor U2187 (N_2187,In_333,In_2575);
xnor U2188 (N_2188,In_250,In_1257);
and U2189 (N_2189,In_1307,In_639);
nor U2190 (N_2190,In_1657,In_2203);
xnor U2191 (N_2191,In_988,In_2491);
nand U2192 (N_2192,In_1615,In_166);
nand U2193 (N_2193,In_2023,In_2016);
xor U2194 (N_2194,In_2695,In_633);
nor U2195 (N_2195,In_894,In_661);
xnor U2196 (N_2196,In_711,In_2760);
or U2197 (N_2197,In_745,In_2721);
nand U2198 (N_2198,In_1833,In_1595);
xor U2199 (N_2199,In_2727,In_1555);
nand U2200 (N_2200,In_1335,In_2328);
or U2201 (N_2201,In_1296,In_1510);
or U2202 (N_2202,In_2873,In_1031);
xor U2203 (N_2203,In_2196,In_2166);
or U2204 (N_2204,In_1235,In_1766);
nand U2205 (N_2205,In_1005,In_2504);
xnor U2206 (N_2206,In_1663,In_981);
and U2207 (N_2207,In_2186,In_63);
or U2208 (N_2208,In_794,In_1679);
xor U2209 (N_2209,In_2327,In_2106);
nor U2210 (N_2210,In_652,In_2563);
or U2211 (N_2211,In_1541,In_2992);
and U2212 (N_2212,In_2777,In_2518);
xor U2213 (N_2213,In_118,In_515);
and U2214 (N_2214,In_2602,In_488);
xor U2215 (N_2215,In_411,In_2540);
or U2216 (N_2216,In_1482,In_2454);
nand U2217 (N_2217,In_954,In_2350);
nand U2218 (N_2218,In_1822,In_865);
or U2219 (N_2219,In_2063,In_768);
and U2220 (N_2220,In_1015,In_362);
xnor U2221 (N_2221,In_1847,In_591);
xnor U2222 (N_2222,In_798,In_383);
nand U2223 (N_2223,In_2857,In_1265);
xor U2224 (N_2224,In_402,In_2341);
nor U2225 (N_2225,In_811,In_2103);
nand U2226 (N_2226,In_558,In_767);
xor U2227 (N_2227,In_1378,In_285);
xnor U2228 (N_2228,In_1615,In_2844);
or U2229 (N_2229,In_2498,In_781);
xor U2230 (N_2230,In_1245,In_1158);
xor U2231 (N_2231,In_1807,In_1936);
nand U2232 (N_2232,In_7,In_2163);
and U2233 (N_2233,In_1756,In_635);
and U2234 (N_2234,In_529,In_544);
and U2235 (N_2235,In_339,In_1605);
and U2236 (N_2236,In_778,In_500);
xnor U2237 (N_2237,In_1472,In_2558);
and U2238 (N_2238,In_2849,In_997);
nand U2239 (N_2239,In_2618,In_787);
nand U2240 (N_2240,In_2384,In_2434);
and U2241 (N_2241,In_878,In_2496);
xnor U2242 (N_2242,In_2864,In_1699);
nand U2243 (N_2243,In_1995,In_2970);
or U2244 (N_2244,In_1102,In_469);
nor U2245 (N_2245,In_894,In_104);
xor U2246 (N_2246,In_2815,In_2392);
xnor U2247 (N_2247,In_1063,In_1642);
nor U2248 (N_2248,In_2107,In_675);
nand U2249 (N_2249,In_2271,In_1950);
or U2250 (N_2250,In_1003,In_1270);
xor U2251 (N_2251,In_93,In_2375);
or U2252 (N_2252,In_1357,In_1301);
nand U2253 (N_2253,In_925,In_2550);
nand U2254 (N_2254,In_2871,In_1547);
nor U2255 (N_2255,In_1633,In_2809);
or U2256 (N_2256,In_1198,In_1581);
and U2257 (N_2257,In_2791,In_233);
and U2258 (N_2258,In_1621,In_1044);
nor U2259 (N_2259,In_2698,In_1740);
xnor U2260 (N_2260,In_806,In_2946);
xor U2261 (N_2261,In_2484,In_1755);
xor U2262 (N_2262,In_2132,In_2326);
xnor U2263 (N_2263,In_1387,In_2571);
xnor U2264 (N_2264,In_472,In_2080);
xor U2265 (N_2265,In_2405,In_2096);
and U2266 (N_2266,In_666,In_2818);
and U2267 (N_2267,In_2179,In_1586);
nor U2268 (N_2268,In_2029,In_397);
xor U2269 (N_2269,In_537,In_1394);
or U2270 (N_2270,In_2214,In_1113);
and U2271 (N_2271,In_2974,In_2786);
nand U2272 (N_2272,In_2434,In_1729);
and U2273 (N_2273,In_668,In_699);
nand U2274 (N_2274,In_1140,In_1710);
xnor U2275 (N_2275,In_908,In_1217);
and U2276 (N_2276,In_1996,In_1572);
or U2277 (N_2277,In_1020,In_361);
xor U2278 (N_2278,In_706,In_2675);
nor U2279 (N_2279,In_87,In_101);
nor U2280 (N_2280,In_2022,In_1595);
xor U2281 (N_2281,In_2770,In_2588);
nand U2282 (N_2282,In_494,In_1743);
nand U2283 (N_2283,In_1097,In_2363);
or U2284 (N_2284,In_2345,In_1884);
or U2285 (N_2285,In_2736,In_2767);
and U2286 (N_2286,In_1102,In_1026);
nand U2287 (N_2287,In_2866,In_2102);
xor U2288 (N_2288,In_2348,In_1080);
nand U2289 (N_2289,In_276,In_1049);
or U2290 (N_2290,In_1944,In_1774);
nand U2291 (N_2291,In_2802,In_1794);
xnor U2292 (N_2292,In_2411,In_1773);
nand U2293 (N_2293,In_2280,In_2986);
nand U2294 (N_2294,In_2417,In_326);
nand U2295 (N_2295,In_1341,In_1511);
nor U2296 (N_2296,In_2580,In_1714);
or U2297 (N_2297,In_2235,In_2745);
nand U2298 (N_2298,In_2836,In_446);
and U2299 (N_2299,In_2079,In_167);
nor U2300 (N_2300,In_2040,In_2042);
nand U2301 (N_2301,In_589,In_1420);
nand U2302 (N_2302,In_259,In_2874);
and U2303 (N_2303,In_581,In_1523);
xnor U2304 (N_2304,In_11,In_774);
xnor U2305 (N_2305,In_2489,In_1701);
xnor U2306 (N_2306,In_442,In_2528);
nand U2307 (N_2307,In_1072,In_741);
nand U2308 (N_2308,In_2978,In_759);
and U2309 (N_2309,In_1432,In_1925);
nand U2310 (N_2310,In_2819,In_549);
or U2311 (N_2311,In_208,In_4);
or U2312 (N_2312,In_466,In_204);
nand U2313 (N_2313,In_1495,In_431);
xor U2314 (N_2314,In_1932,In_381);
nand U2315 (N_2315,In_2758,In_428);
or U2316 (N_2316,In_194,In_1606);
or U2317 (N_2317,In_1257,In_2045);
and U2318 (N_2318,In_891,In_1103);
and U2319 (N_2319,In_485,In_1641);
and U2320 (N_2320,In_1381,In_362);
and U2321 (N_2321,In_2222,In_2522);
xnor U2322 (N_2322,In_1304,In_706);
xor U2323 (N_2323,In_2091,In_484);
or U2324 (N_2324,In_120,In_1763);
or U2325 (N_2325,In_2767,In_854);
and U2326 (N_2326,In_1559,In_2135);
or U2327 (N_2327,In_2543,In_2451);
xor U2328 (N_2328,In_1329,In_2096);
xor U2329 (N_2329,In_2803,In_1640);
nor U2330 (N_2330,In_1031,In_2222);
xor U2331 (N_2331,In_1329,In_1663);
xnor U2332 (N_2332,In_1820,In_2016);
nor U2333 (N_2333,In_2493,In_236);
and U2334 (N_2334,In_2244,In_1731);
nand U2335 (N_2335,In_1595,In_2720);
or U2336 (N_2336,In_2631,In_2580);
nor U2337 (N_2337,In_2632,In_2766);
and U2338 (N_2338,In_1604,In_647);
or U2339 (N_2339,In_1212,In_1241);
nand U2340 (N_2340,In_1946,In_48);
or U2341 (N_2341,In_1553,In_1233);
or U2342 (N_2342,In_1796,In_2173);
and U2343 (N_2343,In_1709,In_2422);
or U2344 (N_2344,In_1662,In_1899);
or U2345 (N_2345,In_157,In_2563);
nand U2346 (N_2346,In_271,In_2955);
nand U2347 (N_2347,In_2035,In_2851);
xnor U2348 (N_2348,In_1110,In_690);
xnor U2349 (N_2349,In_2417,In_1520);
and U2350 (N_2350,In_563,In_433);
or U2351 (N_2351,In_2178,In_1179);
or U2352 (N_2352,In_414,In_2164);
nand U2353 (N_2353,In_2467,In_1009);
and U2354 (N_2354,In_500,In_1619);
xnor U2355 (N_2355,In_592,In_332);
xor U2356 (N_2356,In_356,In_2897);
nor U2357 (N_2357,In_2014,In_2502);
xnor U2358 (N_2358,In_272,In_2480);
and U2359 (N_2359,In_364,In_1661);
or U2360 (N_2360,In_1540,In_2419);
nand U2361 (N_2361,In_604,In_1535);
xnor U2362 (N_2362,In_831,In_2816);
or U2363 (N_2363,In_1773,In_2520);
and U2364 (N_2364,In_1248,In_1928);
nand U2365 (N_2365,In_1158,In_2211);
and U2366 (N_2366,In_2835,In_2134);
or U2367 (N_2367,In_1392,In_1254);
xnor U2368 (N_2368,In_481,In_224);
xnor U2369 (N_2369,In_467,In_1421);
xor U2370 (N_2370,In_2528,In_1573);
xnor U2371 (N_2371,In_2695,In_2381);
nand U2372 (N_2372,In_2408,In_1325);
xnor U2373 (N_2373,In_2057,In_2080);
and U2374 (N_2374,In_246,In_1318);
xor U2375 (N_2375,In_301,In_1168);
nor U2376 (N_2376,In_1805,In_101);
nand U2377 (N_2377,In_1547,In_2379);
nor U2378 (N_2378,In_2267,In_703);
and U2379 (N_2379,In_1552,In_927);
and U2380 (N_2380,In_274,In_2945);
nor U2381 (N_2381,In_1679,In_2499);
and U2382 (N_2382,In_1456,In_611);
xnor U2383 (N_2383,In_2376,In_490);
or U2384 (N_2384,In_2917,In_525);
nand U2385 (N_2385,In_2462,In_1462);
nand U2386 (N_2386,In_744,In_1722);
nor U2387 (N_2387,In_2747,In_314);
nand U2388 (N_2388,In_2045,In_352);
nand U2389 (N_2389,In_1700,In_63);
or U2390 (N_2390,In_1681,In_197);
xor U2391 (N_2391,In_1290,In_2127);
nor U2392 (N_2392,In_2735,In_2320);
nand U2393 (N_2393,In_675,In_2964);
nor U2394 (N_2394,In_125,In_2208);
xor U2395 (N_2395,In_1718,In_2772);
and U2396 (N_2396,In_2043,In_1001);
xor U2397 (N_2397,In_2083,In_2171);
and U2398 (N_2398,In_932,In_992);
nor U2399 (N_2399,In_1309,In_1027);
xor U2400 (N_2400,In_425,In_637);
xnor U2401 (N_2401,In_2816,In_2018);
xor U2402 (N_2402,In_56,In_351);
or U2403 (N_2403,In_1773,In_1062);
nand U2404 (N_2404,In_713,In_2197);
or U2405 (N_2405,In_2039,In_2845);
or U2406 (N_2406,In_1572,In_2139);
xnor U2407 (N_2407,In_2910,In_1878);
and U2408 (N_2408,In_2018,In_2481);
nor U2409 (N_2409,In_2839,In_2237);
nand U2410 (N_2410,In_2209,In_893);
and U2411 (N_2411,In_2030,In_2529);
nand U2412 (N_2412,In_2316,In_1622);
or U2413 (N_2413,In_2857,In_1686);
and U2414 (N_2414,In_2104,In_1275);
nor U2415 (N_2415,In_1464,In_1100);
xor U2416 (N_2416,In_1561,In_1223);
xnor U2417 (N_2417,In_217,In_267);
nor U2418 (N_2418,In_1038,In_324);
xor U2419 (N_2419,In_2603,In_1132);
and U2420 (N_2420,In_1451,In_2419);
xnor U2421 (N_2421,In_2130,In_413);
xnor U2422 (N_2422,In_2774,In_1863);
nor U2423 (N_2423,In_260,In_342);
nand U2424 (N_2424,In_2325,In_1070);
xnor U2425 (N_2425,In_731,In_2254);
or U2426 (N_2426,In_1344,In_2530);
or U2427 (N_2427,In_357,In_1409);
nor U2428 (N_2428,In_2840,In_1814);
and U2429 (N_2429,In_2544,In_618);
nor U2430 (N_2430,In_560,In_387);
nand U2431 (N_2431,In_2188,In_2673);
xnor U2432 (N_2432,In_1230,In_66);
nor U2433 (N_2433,In_1382,In_247);
xor U2434 (N_2434,In_475,In_2926);
or U2435 (N_2435,In_1289,In_2326);
nor U2436 (N_2436,In_404,In_336);
or U2437 (N_2437,In_657,In_2137);
nor U2438 (N_2438,In_559,In_1210);
nor U2439 (N_2439,In_2985,In_1634);
nor U2440 (N_2440,In_776,In_35);
xnor U2441 (N_2441,In_1902,In_107);
xnor U2442 (N_2442,In_2639,In_2666);
nand U2443 (N_2443,In_196,In_1830);
or U2444 (N_2444,In_2351,In_1051);
xor U2445 (N_2445,In_1688,In_1433);
nor U2446 (N_2446,In_2485,In_1687);
nor U2447 (N_2447,In_2200,In_1242);
nand U2448 (N_2448,In_86,In_447);
xnor U2449 (N_2449,In_63,In_2515);
nor U2450 (N_2450,In_2615,In_1473);
nor U2451 (N_2451,In_2768,In_346);
nor U2452 (N_2452,In_59,In_2805);
nor U2453 (N_2453,In_261,In_2566);
and U2454 (N_2454,In_973,In_2998);
nand U2455 (N_2455,In_2423,In_831);
nand U2456 (N_2456,In_558,In_1785);
or U2457 (N_2457,In_1739,In_167);
and U2458 (N_2458,In_1036,In_2329);
nand U2459 (N_2459,In_1186,In_1535);
nand U2460 (N_2460,In_2015,In_2800);
and U2461 (N_2461,In_1121,In_354);
nor U2462 (N_2462,In_2207,In_2349);
nand U2463 (N_2463,In_2089,In_1587);
nand U2464 (N_2464,In_1143,In_221);
xor U2465 (N_2465,In_2105,In_885);
nand U2466 (N_2466,In_2415,In_2101);
nand U2467 (N_2467,In_22,In_922);
and U2468 (N_2468,In_2816,In_2594);
and U2469 (N_2469,In_320,In_1241);
or U2470 (N_2470,In_2089,In_1262);
nand U2471 (N_2471,In_2481,In_2046);
and U2472 (N_2472,In_1710,In_1993);
nand U2473 (N_2473,In_2755,In_2349);
nand U2474 (N_2474,In_998,In_2191);
and U2475 (N_2475,In_1083,In_205);
or U2476 (N_2476,In_2951,In_2803);
xor U2477 (N_2477,In_1923,In_1571);
nor U2478 (N_2478,In_1174,In_692);
nor U2479 (N_2479,In_2641,In_201);
and U2480 (N_2480,In_994,In_151);
nor U2481 (N_2481,In_1427,In_292);
nor U2482 (N_2482,In_2369,In_1974);
nor U2483 (N_2483,In_678,In_722);
or U2484 (N_2484,In_1897,In_2827);
or U2485 (N_2485,In_2419,In_2060);
nor U2486 (N_2486,In_1288,In_2010);
nand U2487 (N_2487,In_1373,In_79);
nand U2488 (N_2488,In_555,In_1217);
nor U2489 (N_2489,In_1523,In_1839);
nor U2490 (N_2490,In_266,In_1102);
and U2491 (N_2491,In_2272,In_2073);
nand U2492 (N_2492,In_2563,In_820);
xor U2493 (N_2493,In_2386,In_525);
nand U2494 (N_2494,In_80,In_271);
xnor U2495 (N_2495,In_2575,In_244);
nand U2496 (N_2496,In_2688,In_1986);
or U2497 (N_2497,In_615,In_2949);
nand U2498 (N_2498,In_1425,In_2837);
nand U2499 (N_2499,In_2138,In_716);
and U2500 (N_2500,In_2234,In_116);
xor U2501 (N_2501,In_1162,In_486);
and U2502 (N_2502,In_807,In_2770);
nor U2503 (N_2503,In_1147,In_2991);
nor U2504 (N_2504,In_412,In_397);
and U2505 (N_2505,In_2825,In_708);
nand U2506 (N_2506,In_2371,In_1867);
and U2507 (N_2507,In_579,In_235);
xor U2508 (N_2508,In_1482,In_2199);
nor U2509 (N_2509,In_456,In_467);
xnor U2510 (N_2510,In_1502,In_2694);
and U2511 (N_2511,In_1686,In_45);
xnor U2512 (N_2512,In_125,In_1592);
and U2513 (N_2513,In_1391,In_2422);
xor U2514 (N_2514,In_1268,In_2767);
nor U2515 (N_2515,In_1272,In_101);
nand U2516 (N_2516,In_347,In_135);
xnor U2517 (N_2517,In_2941,In_289);
nand U2518 (N_2518,In_36,In_2504);
nand U2519 (N_2519,In_1343,In_1397);
and U2520 (N_2520,In_185,In_838);
nor U2521 (N_2521,In_1927,In_1021);
nand U2522 (N_2522,In_894,In_995);
or U2523 (N_2523,In_1837,In_969);
and U2524 (N_2524,In_310,In_607);
nand U2525 (N_2525,In_1628,In_2167);
and U2526 (N_2526,In_2555,In_1963);
and U2527 (N_2527,In_2652,In_1343);
xor U2528 (N_2528,In_1272,In_1242);
and U2529 (N_2529,In_832,In_329);
and U2530 (N_2530,In_2758,In_265);
or U2531 (N_2531,In_2809,In_2043);
and U2532 (N_2532,In_2768,In_1684);
xor U2533 (N_2533,In_2158,In_783);
nor U2534 (N_2534,In_101,In_1840);
and U2535 (N_2535,In_1610,In_2210);
nand U2536 (N_2536,In_2644,In_1829);
nand U2537 (N_2537,In_282,In_1175);
nor U2538 (N_2538,In_2311,In_1495);
nand U2539 (N_2539,In_2519,In_1861);
and U2540 (N_2540,In_1289,In_2635);
nor U2541 (N_2541,In_2616,In_617);
nor U2542 (N_2542,In_2480,In_757);
xnor U2543 (N_2543,In_2625,In_822);
xnor U2544 (N_2544,In_2142,In_2296);
and U2545 (N_2545,In_2056,In_2964);
nor U2546 (N_2546,In_2273,In_488);
xnor U2547 (N_2547,In_1032,In_1909);
nand U2548 (N_2548,In_2452,In_1570);
nor U2549 (N_2549,In_183,In_792);
or U2550 (N_2550,In_1297,In_134);
and U2551 (N_2551,In_735,In_1474);
or U2552 (N_2552,In_2830,In_2298);
xor U2553 (N_2553,In_2343,In_1292);
nand U2554 (N_2554,In_827,In_394);
nand U2555 (N_2555,In_480,In_2999);
nand U2556 (N_2556,In_22,In_2827);
nor U2557 (N_2557,In_420,In_1298);
and U2558 (N_2558,In_2915,In_729);
nor U2559 (N_2559,In_605,In_1159);
nand U2560 (N_2560,In_1735,In_44);
xor U2561 (N_2561,In_1185,In_781);
nor U2562 (N_2562,In_1901,In_20);
nor U2563 (N_2563,In_875,In_1505);
xnor U2564 (N_2564,In_2812,In_1813);
nand U2565 (N_2565,In_419,In_339);
nor U2566 (N_2566,In_2141,In_2112);
nand U2567 (N_2567,In_2096,In_2419);
nand U2568 (N_2568,In_844,In_2355);
or U2569 (N_2569,In_503,In_432);
nor U2570 (N_2570,In_390,In_1699);
nand U2571 (N_2571,In_90,In_1171);
nand U2572 (N_2572,In_650,In_2851);
nand U2573 (N_2573,In_2652,In_1717);
and U2574 (N_2574,In_1089,In_1101);
nand U2575 (N_2575,In_2100,In_2979);
and U2576 (N_2576,In_2054,In_2604);
or U2577 (N_2577,In_126,In_309);
or U2578 (N_2578,In_2956,In_1866);
nor U2579 (N_2579,In_1752,In_1363);
nor U2580 (N_2580,In_1294,In_2504);
nand U2581 (N_2581,In_1764,In_2624);
nand U2582 (N_2582,In_2780,In_543);
or U2583 (N_2583,In_2053,In_2845);
and U2584 (N_2584,In_734,In_1815);
or U2585 (N_2585,In_698,In_780);
or U2586 (N_2586,In_1047,In_1719);
nand U2587 (N_2587,In_2183,In_2908);
nand U2588 (N_2588,In_1752,In_2874);
and U2589 (N_2589,In_73,In_2791);
nand U2590 (N_2590,In_2596,In_656);
nor U2591 (N_2591,In_547,In_650);
and U2592 (N_2592,In_137,In_1811);
xor U2593 (N_2593,In_2806,In_230);
and U2594 (N_2594,In_1366,In_150);
xnor U2595 (N_2595,In_432,In_2662);
and U2596 (N_2596,In_2818,In_2923);
and U2597 (N_2597,In_1560,In_1410);
nand U2598 (N_2598,In_2551,In_2301);
xor U2599 (N_2599,In_2349,In_1186);
nor U2600 (N_2600,In_290,In_548);
nand U2601 (N_2601,In_2575,In_256);
and U2602 (N_2602,In_2034,In_2675);
nand U2603 (N_2603,In_133,In_1783);
nand U2604 (N_2604,In_271,In_2416);
xnor U2605 (N_2605,In_8,In_1559);
xnor U2606 (N_2606,In_1986,In_2621);
xnor U2607 (N_2607,In_2687,In_2972);
nand U2608 (N_2608,In_1135,In_717);
nand U2609 (N_2609,In_2845,In_1483);
and U2610 (N_2610,In_652,In_2196);
xnor U2611 (N_2611,In_1965,In_1243);
and U2612 (N_2612,In_2347,In_890);
or U2613 (N_2613,In_114,In_2109);
and U2614 (N_2614,In_1638,In_1855);
xor U2615 (N_2615,In_625,In_2662);
and U2616 (N_2616,In_1642,In_432);
nor U2617 (N_2617,In_2546,In_126);
and U2618 (N_2618,In_2437,In_1089);
xnor U2619 (N_2619,In_2495,In_1548);
and U2620 (N_2620,In_1809,In_1864);
or U2621 (N_2621,In_130,In_389);
nand U2622 (N_2622,In_49,In_59);
xor U2623 (N_2623,In_1093,In_2740);
nor U2624 (N_2624,In_1179,In_1497);
and U2625 (N_2625,In_230,In_1003);
nand U2626 (N_2626,In_1196,In_986);
xnor U2627 (N_2627,In_216,In_2107);
xor U2628 (N_2628,In_859,In_683);
or U2629 (N_2629,In_1002,In_1792);
xnor U2630 (N_2630,In_1972,In_2676);
xnor U2631 (N_2631,In_2167,In_1235);
nand U2632 (N_2632,In_2281,In_619);
nor U2633 (N_2633,In_1531,In_699);
xor U2634 (N_2634,In_512,In_400);
and U2635 (N_2635,In_2787,In_1913);
or U2636 (N_2636,In_29,In_1088);
nor U2637 (N_2637,In_929,In_2091);
and U2638 (N_2638,In_2588,In_1343);
and U2639 (N_2639,In_1188,In_1070);
and U2640 (N_2640,In_2786,In_759);
nand U2641 (N_2641,In_497,In_751);
nor U2642 (N_2642,In_1101,In_610);
xnor U2643 (N_2643,In_420,In_2611);
nor U2644 (N_2644,In_1095,In_2724);
nand U2645 (N_2645,In_2169,In_2664);
nand U2646 (N_2646,In_367,In_454);
or U2647 (N_2647,In_1403,In_2804);
and U2648 (N_2648,In_495,In_1795);
nor U2649 (N_2649,In_2014,In_2898);
nand U2650 (N_2650,In_1337,In_1511);
xor U2651 (N_2651,In_2466,In_327);
xor U2652 (N_2652,In_774,In_2754);
or U2653 (N_2653,In_2758,In_2252);
nand U2654 (N_2654,In_1343,In_700);
nor U2655 (N_2655,In_1507,In_1102);
or U2656 (N_2656,In_517,In_2550);
xor U2657 (N_2657,In_629,In_1125);
or U2658 (N_2658,In_1994,In_532);
nor U2659 (N_2659,In_581,In_2926);
or U2660 (N_2660,In_233,In_1435);
and U2661 (N_2661,In_811,In_530);
or U2662 (N_2662,In_2300,In_1060);
nand U2663 (N_2663,In_240,In_827);
nor U2664 (N_2664,In_1440,In_2096);
or U2665 (N_2665,In_2150,In_1934);
xnor U2666 (N_2666,In_799,In_2115);
and U2667 (N_2667,In_641,In_974);
and U2668 (N_2668,In_222,In_60);
xnor U2669 (N_2669,In_1123,In_934);
xor U2670 (N_2670,In_2940,In_1685);
nand U2671 (N_2671,In_488,In_1546);
nor U2672 (N_2672,In_1909,In_2577);
nand U2673 (N_2673,In_518,In_2085);
xor U2674 (N_2674,In_1354,In_1540);
or U2675 (N_2675,In_1063,In_306);
or U2676 (N_2676,In_2981,In_2054);
and U2677 (N_2677,In_1211,In_2281);
xor U2678 (N_2678,In_943,In_2719);
xnor U2679 (N_2679,In_212,In_2823);
or U2680 (N_2680,In_364,In_1755);
xnor U2681 (N_2681,In_1960,In_347);
xor U2682 (N_2682,In_2625,In_747);
nand U2683 (N_2683,In_1486,In_410);
xnor U2684 (N_2684,In_1898,In_537);
or U2685 (N_2685,In_2134,In_853);
and U2686 (N_2686,In_433,In_1549);
and U2687 (N_2687,In_1972,In_1331);
and U2688 (N_2688,In_1290,In_213);
nor U2689 (N_2689,In_1353,In_2261);
xor U2690 (N_2690,In_1287,In_1631);
and U2691 (N_2691,In_2613,In_1711);
or U2692 (N_2692,In_1688,In_2097);
or U2693 (N_2693,In_667,In_1695);
nand U2694 (N_2694,In_176,In_1069);
nor U2695 (N_2695,In_1279,In_1557);
and U2696 (N_2696,In_1823,In_1262);
nand U2697 (N_2697,In_1699,In_2949);
or U2698 (N_2698,In_416,In_1582);
nor U2699 (N_2699,In_2044,In_2957);
and U2700 (N_2700,In_1524,In_2642);
and U2701 (N_2701,In_2773,In_2892);
or U2702 (N_2702,In_1785,In_176);
or U2703 (N_2703,In_2508,In_161);
or U2704 (N_2704,In_1454,In_1242);
or U2705 (N_2705,In_1329,In_1165);
or U2706 (N_2706,In_2586,In_2646);
or U2707 (N_2707,In_2058,In_1942);
nor U2708 (N_2708,In_2601,In_2771);
xnor U2709 (N_2709,In_768,In_2023);
nor U2710 (N_2710,In_2474,In_1630);
nand U2711 (N_2711,In_1731,In_2185);
nand U2712 (N_2712,In_555,In_2435);
or U2713 (N_2713,In_395,In_1045);
or U2714 (N_2714,In_1788,In_2202);
and U2715 (N_2715,In_157,In_1095);
or U2716 (N_2716,In_1523,In_464);
xnor U2717 (N_2717,In_1107,In_1121);
xnor U2718 (N_2718,In_2368,In_2444);
xnor U2719 (N_2719,In_178,In_659);
nand U2720 (N_2720,In_1173,In_794);
nand U2721 (N_2721,In_82,In_622);
nand U2722 (N_2722,In_1132,In_235);
and U2723 (N_2723,In_890,In_2463);
and U2724 (N_2724,In_1593,In_1396);
xnor U2725 (N_2725,In_1527,In_1872);
nor U2726 (N_2726,In_612,In_1829);
nand U2727 (N_2727,In_1334,In_1184);
or U2728 (N_2728,In_1579,In_2439);
nor U2729 (N_2729,In_1108,In_1631);
or U2730 (N_2730,In_1698,In_1741);
nor U2731 (N_2731,In_1525,In_1919);
nor U2732 (N_2732,In_373,In_1617);
nor U2733 (N_2733,In_112,In_663);
or U2734 (N_2734,In_530,In_860);
nor U2735 (N_2735,In_1008,In_1371);
or U2736 (N_2736,In_2898,In_2439);
xor U2737 (N_2737,In_97,In_1574);
xor U2738 (N_2738,In_2587,In_2456);
or U2739 (N_2739,In_1299,In_557);
or U2740 (N_2740,In_1808,In_234);
and U2741 (N_2741,In_521,In_2435);
or U2742 (N_2742,In_1589,In_1660);
nand U2743 (N_2743,In_997,In_328);
nor U2744 (N_2744,In_2441,In_883);
xor U2745 (N_2745,In_185,In_2846);
xor U2746 (N_2746,In_2268,In_128);
nor U2747 (N_2747,In_1948,In_656);
or U2748 (N_2748,In_1745,In_1338);
xor U2749 (N_2749,In_1463,In_2451);
nor U2750 (N_2750,In_1583,In_1272);
xnor U2751 (N_2751,In_66,In_2508);
nor U2752 (N_2752,In_340,In_952);
nand U2753 (N_2753,In_707,In_1151);
or U2754 (N_2754,In_1285,In_2436);
xnor U2755 (N_2755,In_2623,In_1814);
nor U2756 (N_2756,In_242,In_73);
xnor U2757 (N_2757,In_1925,In_1888);
nor U2758 (N_2758,In_440,In_2780);
xor U2759 (N_2759,In_1093,In_2923);
or U2760 (N_2760,In_587,In_1514);
or U2761 (N_2761,In_2946,In_1623);
nor U2762 (N_2762,In_2910,In_64);
and U2763 (N_2763,In_2289,In_1579);
nand U2764 (N_2764,In_1112,In_1919);
and U2765 (N_2765,In_21,In_1555);
xor U2766 (N_2766,In_2476,In_1259);
or U2767 (N_2767,In_1554,In_1291);
nor U2768 (N_2768,In_2648,In_751);
xnor U2769 (N_2769,In_235,In_2223);
nor U2770 (N_2770,In_158,In_2829);
xnor U2771 (N_2771,In_2764,In_2658);
nand U2772 (N_2772,In_84,In_2614);
nor U2773 (N_2773,In_2759,In_2949);
nor U2774 (N_2774,In_2256,In_2728);
nand U2775 (N_2775,In_559,In_369);
nor U2776 (N_2776,In_506,In_410);
nor U2777 (N_2777,In_2572,In_1277);
nor U2778 (N_2778,In_1131,In_2112);
nand U2779 (N_2779,In_1027,In_2415);
xor U2780 (N_2780,In_2437,In_2101);
nand U2781 (N_2781,In_1868,In_129);
or U2782 (N_2782,In_2414,In_1201);
xor U2783 (N_2783,In_545,In_2062);
xnor U2784 (N_2784,In_2495,In_319);
nand U2785 (N_2785,In_2946,In_1444);
or U2786 (N_2786,In_1190,In_564);
or U2787 (N_2787,In_2735,In_1427);
or U2788 (N_2788,In_2269,In_1003);
nand U2789 (N_2789,In_853,In_1821);
xor U2790 (N_2790,In_29,In_1885);
nand U2791 (N_2791,In_2978,In_1207);
xnor U2792 (N_2792,In_696,In_1093);
nand U2793 (N_2793,In_1991,In_1851);
nor U2794 (N_2794,In_2066,In_1194);
xnor U2795 (N_2795,In_106,In_1756);
nand U2796 (N_2796,In_2127,In_2375);
and U2797 (N_2797,In_2451,In_1106);
or U2798 (N_2798,In_1252,In_459);
xnor U2799 (N_2799,In_1500,In_2870);
and U2800 (N_2800,In_293,In_2322);
nand U2801 (N_2801,In_2661,In_1593);
nor U2802 (N_2802,In_907,In_1165);
xnor U2803 (N_2803,In_874,In_2862);
and U2804 (N_2804,In_56,In_2171);
xnor U2805 (N_2805,In_2318,In_2782);
nor U2806 (N_2806,In_1868,In_1648);
or U2807 (N_2807,In_1249,In_313);
nand U2808 (N_2808,In_663,In_13);
nor U2809 (N_2809,In_969,In_2072);
nand U2810 (N_2810,In_1721,In_129);
nand U2811 (N_2811,In_2596,In_375);
nand U2812 (N_2812,In_2660,In_399);
nand U2813 (N_2813,In_1052,In_2780);
xor U2814 (N_2814,In_1215,In_646);
and U2815 (N_2815,In_1979,In_2156);
nand U2816 (N_2816,In_351,In_2694);
nor U2817 (N_2817,In_2141,In_885);
nand U2818 (N_2818,In_1077,In_1964);
or U2819 (N_2819,In_2764,In_1549);
nand U2820 (N_2820,In_470,In_1837);
xnor U2821 (N_2821,In_1532,In_1310);
nor U2822 (N_2822,In_2683,In_2944);
nor U2823 (N_2823,In_1911,In_2786);
or U2824 (N_2824,In_2907,In_562);
or U2825 (N_2825,In_2248,In_1928);
xor U2826 (N_2826,In_1777,In_1442);
nor U2827 (N_2827,In_1984,In_297);
xnor U2828 (N_2828,In_181,In_1626);
and U2829 (N_2829,In_1826,In_2458);
nor U2830 (N_2830,In_1663,In_584);
nor U2831 (N_2831,In_2660,In_1834);
nand U2832 (N_2832,In_935,In_2722);
or U2833 (N_2833,In_2561,In_614);
xnor U2834 (N_2834,In_1663,In_104);
nand U2835 (N_2835,In_2866,In_1472);
and U2836 (N_2836,In_80,In_115);
and U2837 (N_2837,In_2602,In_786);
and U2838 (N_2838,In_2463,In_60);
nand U2839 (N_2839,In_2551,In_2773);
nand U2840 (N_2840,In_1156,In_246);
or U2841 (N_2841,In_1450,In_2130);
nor U2842 (N_2842,In_845,In_1583);
and U2843 (N_2843,In_766,In_1326);
and U2844 (N_2844,In_2694,In_1520);
nor U2845 (N_2845,In_1339,In_1251);
nor U2846 (N_2846,In_2899,In_2842);
nor U2847 (N_2847,In_2852,In_1992);
xnor U2848 (N_2848,In_2465,In_1766);
or U2849 (N_2849,In_19,In_1201);
or U2850 (N_2850,In_2017,In_1800);
nand U2851 (N_2851,In_1745,In_332);
or U2852 (N_2852,In_1637,In_1137);
xnor U2853 (N_2853,In_1619,In_907);
xnor U2854 (N_2854,In_346,In_2517);
nor U2855 (N_2855,In_1585,In_860);
nor U2856 (N_2856,In_326,In_2098);
xor U2857 (N_2857,In_16,In_2132);
and U2858 (N_2858,In_2853,In_2328);
or U2859 (N_2859,In_1636,In_2855);
nand U2860 (N_2860,In_985,In_515);
nor U2861 (N_2861,In_666,In_2931);
xor U2862 (N_2862,In_320,In_495);
nor U2863 (N_2863,In_1162,In_1923);
nand U2864 (N_2864,In_694,In_833);
or U2865 (N_2865,In_2367,In_432);
nand U2866 (N_2866,In_2565,In_1095);
nand U2867 (N_2867,In_1430,In_2757);
or U2868 (N_2868,In_1780,In_279);
and U2869 (N_2869,In_2740,In_1985);
and U2870 (N_2870,In_1296,In_312);
xor U2871 (N_2871,In_852,In_528);
xor U2872 (N_2872,In_2444,In_1886);
nand U2873 (N_2873,In_1542,In_2760);
xor U2874 (N_2874,In_600,In_1065);
nor U2875 (N_2875,In_19,In_2441);
xor U2876 (N_2876,In_2445,In_378);
or U2877 (N_2877,In_126,In_1777);
nor U2878 (N_2878,In_2287,In_747);
and U2879 (N_2879,In_1682,In_131);
nand U2880 (N_2880,In_1207,In_231);
xor U2881 (N_2881,In_1783,In_1560);
nor U2882 (N_2882,In_241,In_1054);
and U2883 (N_2883,In_1277,In_2959);
or U2884 (N_2884,In_2495,In_2138);
xnor U2885 (N_2885,In_1326,In_1531);
or U2886 (N_2886,In_1727,In_337);
or U2887 (N_2887,In_1609,In_1982);
or U2888 (N_2888,In_2681,In_56);
xor U2889 (N_2889,In_2241,In_2328);
nor U2890 (N_2890,In_441,In_2368);
nand U2891 (N_2891,In_2521,In_64);
nor U2892 (N_2892,In_2221,In_2906);
nand U2893 (N_2893,In_436,In_339);
xor U2894 (N_2894,In_2888,In_2541);
or U2895 (N_2895,In_462,In_1788);
nand U2896 (N_2896,In_676,In_304);
nand U2897 (N_2897,In_2219,In_2606);
and U2898 (N_2898,In_76,In_1017);
nand U2899 (N_2899,In_1065,In_506);
nor U2900 (N_2900,In_170,In_91);
xnor U2901 (N_2901,In_458,In_2470);
nor U2902 (N_2902,In_2720,In_2231);
nand U2903 (N_2903,In_1364,In_1830);
and U2904 (N_2904,In_1990,In_2115);
or U2905 (N_2905,In_1537,In_700);
nor U2906 (N_2906,In_1323,In_1996);
or U2907 (N_2907,In_1492,In_1981);
or U2908 (N_2908,In_2397,In_1965);
and U2909 (N_2909,In_1457,In_1353);
and U2910 (N_2910,In_618,In_2691);
and U2911 (N_2911,In_2015,In_2756);
nor U2912 (N_2912,In_1488,In_2393);
xor U2913 (N_2913,In_1772,In_2134);
and U2914 (N_2914,In_1100,In_790);
or U2915 (N_2915,In_1590,In_221);
xnor U2916 (N_2916,In_2215,In_2765);
nor U2917 (N_2917,In_640,In_2117);
and U2918 (N_2918,In_574,In_191);
nand U2919 (N_2919,In_2289,In_259);
or U2920 (N_2920,In_1967,In_1000);
nor U2921 (N_2921,In_1331,In_2647);
and U2922 (N_2922,In_2179,In_2699);
xnor U2923 (N_2923,In_2033,In_2368);
nor U2924 (N_2924,In_2993,In_1929);
xnor U2925 (N_2925,In_634,In_772);
nor U2926 (N_2926,In_258,In_674);
xor U2927 (N_2927,In_704,In_2762);
and U2928 (N_2928,In_1046,In_131);
nor U2929 (N_2929,In_1226,In_2459);
nand U2930 (N_2930,In_1377,In_1650);
nand U2931 (N_2931,In_1732,In_1977);
and U2932 (N_2932,In_394,In_1300);
and U2933 (N_2933,In_1655,In_2443);
xnor U2934 (N_2934,In_1710,In_868);
xnor U2935 (N_2935,In_2621,In_1242);
nor U2936 (N_2936,In_2579,In_2900);
nand U2937 (N_2937,In_915,In_1264);
or U2938 (N_2938,In_276,In_2444);
nor U2939 (N_2939,In_382,In_1282);
and U2940 (N_2940,In_2342,In_2769);
and U2941 (N_2941,In_2418,In_367);
nand U2942 (N_2942,In_382,In_256);
xor U2943 (N_2943,In_2932,In_31);
or U2944 (N_2944,In_2570,In_1384);
and U2945 (N_2945,In_2294,In_2043);
or U2946 (N_2946,In_1116,In_1570);
xnor U2947 (N_2947,In_698,In_2904);
nand U2948 (N_2948,In_1384,In_755);
nand U2949 (N_2949,In_23,In_2883);
nand U2950 (N_2950,In_854,In_1696);
xor U2951 (N_2951,In_182,In_566);
and U2952 (N_2952,In_415,In_1619);
nand U2953 (N_2953,In_66,In_586);
and U2954 (N_2954,In_1999,In_1066);
nand U2955 (N_2955,In_316,In_1567);
or U2956 (N_2956,In_30,In_530);
or U2957 (N_2957,In_936,In_1728);
or U2958 (N_2958,In_2020,In_684);
nor U2959 (N_2959,In_333,In_591);
nor U2960 (N_2960,In_1247,In_833);
or U2961 (N_2961,In_1124,In_719);
xnor U2962 (N_2962,In_1397,In_72);
and U2963 (N_2963,In_1632,In_314);
nand U2964 (N_2964,In_204,In_131);
or U2965 (N_2965,In_259,In_1202);
nor U2966 (N_2966,In_1168,In_1616);
xnor U2967 (N_2967,In_16,In_2187);
nor U2968 (N_2968,In_1127,In_1607);
nor U2969 (N_2969,In_1000,In_2860);
xnor U2970 (N_2970,In_872,In_187);
nand U2971 (N_2971,In_2649,In_2308);
and U2972 (N_2972,In_1899,In_2270);
or U2973 (N_2973,In_1271,In_1726);
and U2974 (N_2974,In_1401,In_360);
or U2975 (N_2975,In_1203,In_1974);
nor U2976 (N_2976,In_2961,In_2444);
nor U2977 (N_2977,In_2548,In_881);
xor U2978 (N_2978,In_204,In_2575);
or U2979 (N_2979,In_1332,In_2385);
and U2980 (N_2980,In_2827,In_2856);
nand U2981 (N_2981,In_998,In_1202);
xor U2982 (N_2982,In_1438,In_1573);
nand U2983 (N_2983,In_1445,In_128);
nor U2984 (N_2984,In_1388,In_2887);
xnor U2985 (N_2985,In_2261,In_2970);
xor U2986 (N_2986,In_1725,In_345);
nor U2987 (N_2987,In_814,In_539);
nor U2988 (N_2988,In_2875,In_2350);
or U2989 (N_2989,In_2376,In_1398);
nor U2990 (N_2990,In_1093,In_1930);
nor U2991 (N_2991,In_1229,In_1943);
nand U2992 (N_2992,In_2191,In_144);
xor U2993 (N_2993,In_2554,In_1607);
nor U2994 (N_2994,In_1285,In_2238);
xor U2995 (N_2995,In_884,In_2012);
nor U2996 (N_2996,In_1360,In_2452);
and U2997 (N_2997,In_1976,In_424);
xor U2998 (N_2998,In_1432,In_1292);
or U2999 (N_2999,In_902,In_2503);
xnor U3000 (N_3000,N_1010,N_2832);
or U3001 (N_3001,N_2815,N_1158);
nand U3002 (N_3002,N_2376,N_2227);
and U3003 (N_3003,N_1812,N_1904);
xnor U3004 (N_3004,N_2858,N_1244);
nand U3005 (N_3005,N_1971,N_1004);
and U3006 (N_3006,N_764,N_357);
nand U3007 (N_3007,N_457,N_467);
or U3008 (N_3008,N_1151,N_2439);
and U3009 (N_3009,N_1930,N_1814);
or U3010 (N_3010,N_780,N_1515);
nand U3011 (N_3011,N_2324,N_2842);
or U3012 (N_3012,N_1332,N_117);
or U3013 (N_3013,N_113,N_1961);
or U3014 (N_3014,N_417,N_2702);
nor U3015 (N_3015,N_456,N_1622);
and U3016 (N_3016,N_2345,N_2387);
or U3017 (N_3017,N_1299,N_1140);
xnor U3018 (N_3018,N_801,N_1389);
or U3019 (N_3019,N_2887,N_1231);
xnor U3020 (N_3020,N_2169,N_2148);
or U3021 (N_3021,N_572,N_2817);
and U3022 (N_3022,N_950,N_2233);
xnor U3023 (N_3023,N_2911,N_2728);
and U3024 (N_3024,N_2602,N_628);
xor U3025 (N_3025,N_1734,N_2415);
nor U3026 (N_3026,N_1426,N_591);
or U3027 (N_3027,N_74,N_1078);
xnor U3028 (N_3028,N_2119,N_1890);
and U3029 (N_3029,N_161,N_488);
or U3030 (N_3030,N_2133,N_778);
or U3031 (N_3031,N_364,N_2459);
and U3032 (N_3032,N_2481,N_404);
nor U3033 (N_3033,N_1459,N_2562);
nand U3034 (N_3034,N_694,N_605);
nor U3035 (N_3035,N_2897,N_2218);
and U3036 (N_3036,N_1778,N_2098);
or U3037 (N_3037,N_2157,N_14);
xnor U3038 (N_3038,N_552,N_1540);
nor U3039 (N_3039,N_1434,N_284);
nand U3040 (N_3040,N_2733,N_1940);
and U3041 (N_3041,N_1290,N_2834);
nor U3042 (N_3042,N_1900,N_2927);
or U3043 (N_3043,N_2706,N_843);
nor U3044 (N_3044,N_2285,N_2339);
and U3045 (N_3045,N_2498,N_750);
nand U3046 (N_3046,N_2045,N_2076);
nand U3047 (N_3047,N_351,N_1929);
nand U3048 (N_3048,N_1356,N_1935);
nor U3049 (N_3049,N_899,N_783);
nor U3050 (N_3050,N_2759,N_2618);
and U3051 (N_3051,N_1797,N_127);
or U3052 (N_3052,N_2021,N_964);
nor U3053 (N_3053,N_390,N_1892);
and U3054 (N_3054,N_2626,N_1784);
nand U3055 (N_3055,N_2305,N_641);
or U3056 (N_3056,N_312,N_1427);
xor U3057 (N_3057,N_2968,N_1988);
nand U3058 (N_3058,N_2757,N_1313);
nor U3059 (N_3059,N_1106,N_805);
and U3060 (N_3060,N_2752,N_1191);
and U3061 (N_3061,N_294,N_1746);
nand U3062 (N_3062,N_1287,N_2585);
xnor U3063 (N_3063,N_111,N_724);
or U3064 (N_3064,N_2252,N_333);
nor U3065 (N_3065,N_68,N_558);
xnor U3066 (N_3066,N_1508,N_2317);
nand U3067 (N_3067,N_665,N_1333);
or U3068 (N_3068,N_1410,N_2939);
and U3069 (N_3069,N_278,N_1517);
nor U3070 (N_3070,N_388,N_1009);
nand U3071 (N_3071,N_1700,N_658);
nand U3072 (N_3072,N_1314,N_1268);
nand U3073 (N_3073,N_1882,N_37);
xor U3074 (N_3074,N_2994,N_1371);
or U3075 (N_3075,N_2126,N_2782);
and U3076 (N_3076,N_1589,N_2807);
and U3077 (N_3077,N_2427,N_2686);
nand U3078 (N_3078,N_2494,N_151);
nand U3079 (N_3079,N_561,N_2957);
or U3080 (N_3080,N_1302,N_148);
or U3081 (N_3081,N_2643,N_249);
xnor U3082 (N_3082,N_2599,N_2668);
nand U3083 (N_3083,N_2596,N_1458);
nand U3084 (N_3084,N_1196,N_2783);
or U3085 (N_3085,N_2322,N_1130);
nor U3086 (N_3086,N_2223,N_2767);
nand U3087 (N_3087,N_2907,N_2342);
and U3088 (N_3088,N_1505,N_1876);
nor U3089 (N_3089,N_2992,N_2377);
nor U3090 (N_3090,N_675,N_2306);
nand U3091 (N_3091,N_2117,N_1174);
and U3092 (N_3092,N_2298,N_671);
nor U3093 (N_3093,N_474,N_2120);
nor U3094 (N_3094,N_2823,N_316);
nor U3095 (N_3095,N_1133,N_1858);
nor U3096 (N_3096,N_2205,N_2676);
nand U3097 (N_3097,N_216,N_1147);
nand U3098 (N_3098,N_2959,N_1249);
and U3099 (N_3099,N_159,N_1412);
xnor U3100 (N_3100,N_1295,N_989);
xnor U3101 (N_3101,N_859,N_2932);
and U3102 (N_3102,N_2154,N_551);
xnor U3103 (N_3103,N_1834,N_189);
nand U3104 (N_3104,N_2809,N_708);
nand U3105 (N_3105,N_1733,N_996);
nand U3106 (N_3106,N_1730,N_512);
and U3107 (N_3107,N_459,N_2040);
and U3108 (N_3108,N_1316,N_2244);
xnor U3109 (N_3109,N_358,N_570);
and U3110 (N_3110,N_1280,N_1217);
and U3111 (N_3111,N_2852,N_2193);
or U3112 (N_3112,N_1139,N_2988);
or U3113 (N_3113,N_877,N_1388);
and U3114 (N_3114,N_1861,N_2810);
and U3115 (N_3115,N_98,N_777);
or U3116 (N_3116,N_637,N_1568);
or U3117 (N_3117,N_2636,N_2138);
and U3118 (N_3118,N_257,N_1799);
and U3119 (N_3119,N_1918,N_2411);
and U3120 (N_3120,N_543,N_355);
or U3121 (N_3121,N_422,N_1845);
nor U3122 (N_3122,N_2447,N_1786);
and U3123 (N_3123,N_218,N_1126);
and U3124 (N_3124,N_639,N_28);
xor U3125 (N_3125,N_1436,N_1398);
nand U3126 (N_3126,N_2836,N_46);
xor U3127 (N_3127,N_2627,N_2066);
nand U3128 (N_3128,N_2987,N_2026);
or U3129 (N_3129,N_2956,N_2257);
and U3130 (N_3130,N_1770,N_2129);
xnor U3131 (N_3131,N_2850,N_581);
and U3132 (N_3132,N_2487,N_1857);
nor U3133 (N_3133,N_1723,N_2327);
and U3134 (N_3134,N_1198,N_1652);
and U3135 (N_3135,N_2267,N_2990);
or U3136 (N_3136,N_2640,N_1941);
nand U3137 (N_3137,N_391,N_880);
and U3138 (N_3138,N_2450,N_1162);
and U3139 (N_3139,N_1645,N_541);
or U3140 (N_3140,N_2632,N_1600);
or U3141 (N_3141,N_2480,N_2028);
and U3142 (N_3142,N_1190,N_85);
nand U3143 (N_3143,N_1493,N_405);
nand U3144 (N_3144,N_933,N_1632);
and U3145 (N_3145,N_2680,N_1362);
nor U3146 (N_3146,N_436,N_505);
and U3147 (N_3147,N_2540,N_2857);
nand U3148 (N_3148,N_657,N_553);
or U3149 (N_3149,N_1115,N_2399);
xor U3150 (N_3150,N_872,N_1704);
xnor U3151 (N_3151,N_1644,N_2710);
or U3152 (N_3152,N_1418,N_1141);
nor U3153 (N_3153,N_825,N_1509);
nand U3154 (N_3154,N_210,N_1895);
nand U3155 (N_3155,N_282,N_279);
nor U3156 (N_3156,N_2916,N_2266);
and U3157 (N_3157,N_64,N_1794);
nor U3158 (N_3158,N_1820,N_2280);
or U3159 (N_3159,N_2406,N_2435);
nand U3160 (N_3160,N_994,N_112);
or U3161 (N_3161,N_1576,N_237);
and U3162 (N_3162,N_1283,N_2981);
and U3163 (N_3163,N_2657,N_269);
nor U3164 (N_3164,N_2228,N_584);
nand U3165 (N_3165,N_1286,N_1042);
and U3166 (N_3166,N_302,N_696);
xnor U3167 (N_3167,N_2938,N_555);
xor U3168 (N_3168,N_1604,N_1945);
xor U3169 (N_3169,N_475,N_2732);
nand U3170 (N_3170,N_1226,N_2433);
nor U3171 (N_3171,N_753,N_244);
and U3172 (N_3172,N_430,N_2371);
nand U3173 (N_3173,N_710,N_582);
nor U3174 (N_3174,N_612,N_2763);
xor U3175 (N_3175,N_2720,N_485);
and U3176 (N_3176,N_530,N_854);
and U3177 (N_3177,N_2388,N_450);
nor U3178 (N_3178,N_1021,N_17);
and U3179 (N_3179,N_377,N_2774);
nor U3180 (N_3180,N_147,N_35);
xor U3181 (N_3181,N_1178,N_2110);
nand U3182 (N_3182,N_2895,N_1579);
nand U3183 (N_3183,N_349,N_2695);
and U3184 (N_3184,N_2806,N_1229);
nor U3185 (N_3185,N_1346,N_1052);
nor U3186 (N_3186,N_1179,N_803);
xor U3187 (N_3187,N_1536,N_2422);
and U3188 (N_3188,N_517,N_2569);
and U3189 (N_3189,N_863,N_874);
nand U3190 (N_3190,N_744,N_1938);
xnor U3191 (N_3191,N_400,N_2063);
xor U3192 (N_3192,N_451,N_2017);
or U3193 (N_3193,N_1109,N_2923);
nor U3194 (N_3194,N_2242,N_1867);
nor U3195 (N_3195,N_1987,N_1699);
nand U3196 (N_3196,N_1888,N_701);
or U3197 (N_3197,N_2854,N_1233);
nand U3198 (N_3198,N_22,N_48);
and U3199 (N_3199,N_908,N_2265);
and U3200 (N_3200,N_84,N_1532);
nor U3201 (N_3201,N_2699,N_2264);
xnor U3202 (N_3202,N_290,N_1897);
nand U3203 (N_3203,N_674,N_407);
or U3204 (N_3204,N_856,N_170);
and U3205 (N_3205,N_1447,N_2697);
and U3206 (N_3206,N_67,N_368);
nand U3207 (N_3207,N_2163,N_215);
nand U3208 (N_3208,N_493,N_2894);
nor U3209 (N_3209,N_1815,N_981);
xor U3210 (N_3210,N_336,N_2115);
nor U3211 (N_3211,N_1970,N_2507);
xor U3212 (N_3212,N_238,N_2600);
or U3213 (N_3213,N_2597,N_108);
nor U3214 (N_3214,N_449,N_2598);
and U3215 (N_3215,N_1791,N_894);
or U3216 (N_3216,N_2917,N_668);
xnor U3217 (N_3217,N_1007,N_609);
xnor U3218 (N_3218,N_326,N_1658);
xor U3219 (N_3219,N_259,N_1457);
xnor U3220 (N_3220,N_2593,N_2079);
nand U3221 (N_3221,N_2928,N_1949);
or U3222 (N_3222,N_596,N_2455);
or U3223 (N_3223,N_2194,N_321);
or U3224 (N_3224,N_2426,N_522);
and U3225 (N_3225,N_939,N_1461);
xnor U3226 (N_3226,N_1683,N_2364);
nor U3227 (N_3227,N_1850,N_2178);
nor U3228 (N_3228,N_506,N_2440);
xnor U3229 (N_3229,N_478,N_63);
xor U3230 (N_3230,N_49,N_2226);
or U3231 (N_3231,N_1762,N_2344);
or U3232 (N_3232,N_871,N_1027);
and U3233 (N_3233,N_2742,N_2261);
nand U3234 (N_3234,N_763,N_1610);
nor U3235 (N_3235,N_1101,N_1959);
xor U3236 (N_3236,N_633,N_2294);
or U3237 (N_3237,N_115,N_2681);
and U3238 (N_3238,N_589,N_2508);
nor U3239 (N_3239,N_2064,N_311);
nand U3240 (N_3240,N_2013,N_1011);
or U3241 (N_3241,N_1006,N_1967);
nor U3242 (N_3242,N_2660,N_2086);
or U3243 (N_3243,N_2696,N_2007);
and U3244 (N_3244,N_1430,N_2047);
xnor U3245 (N_3245,N_2308,N_739);
nand U3246 (N_3246,N_145,N_546);
nand U3247 (N_3247,N_268,N_1124);
and U3248 (N_3248,N_2184,N_1686);
nand U3249 (N_3249,N_2675,N_2984);
xor U3250 (N_3250,N_443,N_1752);
and U3251 (N_3251,N_901,N_673);
nor U3252 (N_3252,N_43,N_2151);
nor U3253 (N_3253,N_1891,N_150);
and U3254 (N_3254,N_464,N_389);
and U3255 (N_3255,N_1444,N_2094);
xnor U3256 (N_3256,N_274,N_1616);
xor U3257 (N_3257,N_2551,N_1975);
or U3258 (N_3258,N_2030,N_1466);
nor U3259 (N_3259,N_2029,N_2878);
or U3260 (N_3260,N_1617,N_2531);
or U3261 (N_3261,N_1340,N_525);
xor U3262 (N_3262,N_2396,N_1423);
xor U3263 (N_3263,N_1860,N_926);
nor U3264 (N_3264,N_57,N_1926);
nor U3265 (N_3265,N_500,N_1354);
and U3266 (N_3266,N_1511,N_2018);
nor U3267 (N_3267,N_1728,N_1747);
nor U3268 (N_3268,N_1634,N_1761);
or U3269 (N_3269,N_1074,N_394);
or U3270 (N_3270,N_1460,N_1152);
nand U3271 (N_3271,N_1881,N_1242);
and U3272 (N_3272,N_53,N_2457);
nor U3273 (N_3273,N_1467,N_1199);
nor U3274 (N_3274,N_2526,N_1836);
nand U3275 (N_3275,N_2830,N_1090);
nor U3276 (N_3276,N_1525,N_2088);
nor U3277 (N_3277,N_1702,N_1574);
xnor U3278 (N_3278,N_1779,N_782);
or U3279 (N_3279,N_2413,N_2870);
and U3280 (N_3280,N_415,N_942);
nor U3281 (N_3281,N_1558,N_1781);
nand U3282 (N_3282,N_71,N_82);
or U3283 (N_3283,N_2141,N_1489);
and U3284 (N_3284,N_1901,N_2853);
nand U3285 (N_3285,N_1394,N_2645);
and U3286 (N_3286,N_1972,N_2886);
or U3287 (N_3287,N_684,N_692);
xor U3288 (N_3288,N_1353,N_1565);
nand U3289 (N_3289,N_1392,N_1232);
and U3290 (N_3290,N_1985,N_2448);
xor U3291 (N_3291,N_2725,N_126);
xor U3292 (N_3292,N_2014,N_1326);
nand U3293 (N_3293,N_1017,N_1735);
and U3294 (N_3294,N_306,N_2472);
or U3295 (N_3295,N_1303,N_1486);
and U3296 (N_3296,N_2271,N_1800);
nand U3297 (N_3297,N_2882,N_2880);
xor U3298 (N_3298,N_2254,N_109);
nand U3299 (N_3299,N_1393,N_130);
xor U3300 (N_3300,N_2476,N_2682);
and U3301 (N_3301,N_1107,N_1218);
xnor U3302 (N_3302,N_102,N_212);
nand U3303 (N_3303,N_1189,N_1056);
nor U3304 (N_3304,N_2665,N_1468);
nor U3305 (N_3305,N_826,N_164);
and U3306 (N_3306,N_2292,N_2691);
nor U3307 (N_3307,N_2779,N_2952);
nand U3308 (N_3308,N_2397,N_2370);
and U3309 (N_3309,N_1663,N_667);
xor U3310 (N_3310,N_2859,N_413);
xnor U3311 (N_3311,N_559,N_2719);
and U3312 (N_3312,N_402,N_2515);
nor U3313 (N_3313,N_95,N_1349);
or U3314 (N_3314,N_1990,N_932);
nand U3315 (N_3315,N_2042,N_1494);
nor U3316 (N_3316,N_1059,N_1086);
and U3317 (N_3317,N_1539,N_1236);
and U3318 (N_3318,N_700,N_2136);
or U3319 (N_3319,N_2239,N_534);
nand U3320 (N_3320,N_1611,N_1046);
nand U3321 (N_3321,N_2062,N_1753);
and U3322 (N_3322,N_554,N_354);
xor U3323 (N_3323,N_757,N_75);
and U3324 (N_3324,N_248,N_2855);
xor U3325 (N_3325,N_1265,N_2052);
nand U3326 (N_3326,N_850,N_393);
xnor U3327 (N_3327,N_1002,N_2466);
and U3328 (N_3328,N_1998,N_233);
xnor U3329 (N_3329,N_1035,N_904);
or U3330 (N_3330,N_317,N_1308);
xor U3331 (N_3331,N_718,N_2482);
and U3332 (N_3332,N_1832,N_47);
nor U3333 (N_3333,N_878,N_2824);
nor U3334 (N_3334,N_273,N_2847);
nor U3335 (N_3335,N_549,N_599);
and U3336 (N_3336,N_1586,N_1089);
nor U3337 (N_3337,N_1275,N_1562);
nor U3338 (N_3338,N_1813,N_1448);
and U3339 (N_3339,N_2024,N_177);
nor U3340 (N_3340,N_751,N_2049);
or U3341 (N_3341,N_2612,N_742);
or U3342 (N_3342,N_137,N_460);
nor U3343 (N_3343,N_1722,N_66);
or U3344 (N_3344,N_2549,N_1245);
nand U3345 (N_3345,N_1592,N_2412);
nand U3346 (N_3346,N_1903,N_479);
xor U3347 (N_3347,N_2838,N_2423);
xnor U3348 (N_3348,N_1479,N_2799);
nand U3349 (N_3349,N_535,N_2142);
xor U3350 (N_3350,N_2320,N_2579);
xor U3351 (N_3351,N_240,N_624);
xor U3352 (N_3352,N_1053,N_828);
or U3353 (N_3353,N_1667,N_1931);
xnor U3354 (N_3354,N_473,N_9);
nand U3355 (N_3355,N_296,N_1624);
xnor U3356 (N_3356,N_1880,N_12);
xor U3357 (N_3357,N_518,N_1519);
nand U3358 (N_3358,N_371,N_1962);
xor U3359 (N_3359,N_2666,N_2189);
nor U3360 (N_3360,N_2789,N_2528);
nor U3361 (N_3361,N_2970,N_977);
or U3362 (N_3362,N_96,N_45);
or U3363 (N_3363,N_494,N_951);
or U3364 (N_3364,N_1289,N_288);
xnor U3365 (N_3365,N_2827,N_144);
and U3366 (N_3366,N_2492,N_2524);
nand U3367 (N_3367,N_136,N_2761);
or U3368 (N_3368,N_1057,N_666);
nor U3369 (N_3369,N_2467,N_1391);
and U3370 (N_3370,N_2404,N_1964);
and U3371 (N_3371,N_1177,N_2619);
and U3372 (N_3372,N_1194,N_1201);
or U3373 (N_3373,N_250,N_2654);
xnor U3374 (N_3374,N_135,N_2560);
nand U3375 (N_3375,N_1811,N_110);
nor U3376 (N_3376,N_1269,N_2253);
nand U3377 (N_3377,N_123,N_196);
nor U3378 (N_3378,N_2283,N_1122);
nor U3379 (N_3379,N_2912,N_2776);
or U3380 (N_3380,N_1965,N_2837);
xnor U3381 (N_3381,N_142,N_1409);
and U3382 (N_3382,N_676,N_2653);
and U3383 (N_3383,N_532,N_2888);
nand U3384 (N_3384,N_1749,N_209);
or U3385 (N_3385,N_313,N_719);
nor U3386 (N_3386,N_563,N_1015);
nand U3387 (N_3387,N_1739,N_2158);
or U3388 (N_3388,N_2209,N_806);
or U3389 (N_3389,N_1476,N_1344);
and U3390 (N_3390,N_2258,N_1403);
nor U3391 (N_3391,N_1503,N_1069);
nor U3392 (N_3392,N_2519,N_1756);
and U3393 (N_3393,N_601,N_2249);
and U3394 (N_3394,N_2769,N_426);
nor U3395 (N_3395,N_414,N_2937);
or U3396 (N_3396,N_2896,N_2785);
nor U3397 (N_3397,N_1318,N_1358);
xnor U3398 (N_3398,N_1480,N_1963);
xnor U3399 (N_3399,N_1243,N_2892);
nand U3400 (N_3400,N_1094,N_89);
nor U3401 (N_3401,N_2875,N_1270);
and U3402 (N_3402,N_2590,N_2445);
nand U3403 (N_3403,N_925,N_2478);
xnor U3404 (N_3404,N_481,N_1615);
xor U3405 (N_3405,N_2991,N_1135);
and U3406 (N_3406,N_2944,N_1414);
xnor U3407 (N_3407,N_1530,N_2974);
nor U3408 (N_3408,N_2514,N_1385);
or U3409 (N_3409,N_1682,N_2967);
nor U3410 (N_3410,N_2260,N_162);
nand U3411 (N_3411,N_2068,N_1185);
xor U3412 (N_3412,N_2424,N_1014);
nor U3413 (N_3413,N_616,N_2846);
or U3414 (N_3414,N_403,N_2576);
and U3415 (N_3415,N_2051,N_194);
nor U3416 (N_3416,N_2350,N_1060);
or U3417 (N_3417,N_303,N_425);
nand U3418 (N_3418,N_2337,N_1446);
and U3419 (N_3419,N_2224,N_527);
nand U3420 (N_3420,N_2452,N_1087);
and U3421 (N_3421,N_2667,N_575);
or U3422 (N_3422,N_1347,N_2070);
xnor U3423 (N_3423,N_469,N_1228);
or U3424 (N_3424,N_513,N_2711);
xor U3425 (N_3425,N_1205,N_957);
nand U3426 (N_3426,N_491,N_1743);
nand U3427 (N_3427,N_1137,N_2085);
and U3428 (N_3428,N_1100,N_401);
or U3429 (N_3429,N_341,N_2281);
nand U3430 (N_3430,N_738,N_804);
nand U3431 (N_3431,N_770,N_1116);
nor U3432 (N_3432,N_1348,N_1870);
nor U3433 (N_3433,N_1977,N_1950);
xnor U3434 (N_3434,N_2,N_677);
or U3435 (N_3435,N_93,N_1176);
or U3436 (N_3436,N_823,N_997);
nand U3437 (N_3437,N_315,N_384);
nor U3438 (N_3438,N_1569,N_2207);
and U3439 (N_3439,N_699,N_726);
nor U3440 (N_3440,N_246,N_1921);
or U3441 (N_3441,N_1363,N_116);
or U3442 (N_3442,N_956,N_1309);
and U3443 (N_3443,N_155,N_647);
xor U3444 (N_3444,N_1550,N_2962);
nand U3445 (N_3445,N_669,N_56);
and U3446 (N_3446,N_1361,N_608);
and U3447 (N_3447,N_2997,N_2659);
nand U3448 (N_3448,N_1750,N_2383);
and U3449 (N_3449,N_2693,N_2831);
nand U3450 (N_3450,N_329,N_1104);
nor U3451 (N_3451,N_2794,N_490);
xnor U3452 (N_3452,N_2278,N_911);
and U3453 (N_3453,N_953,N_2468);
nand U3454 (N_3454,N_2731,N_2536);
xnor U3455 (N_3455,N_1922,N_510);
or U3456 (N_3456,N_2269,N_1654);
and U3457 (N_3457,N_2754,N_2945);
nand U3458 (N_3458,N_2357,N_1148);
nor U3459 (N_3459,N_2712,N_1885);
nor U3460 (N_3460,N_1470,N_1830);
nand U3461 (N_3461,N_1334,N_2958);
nand U3462 (N_3462,N_2301,N_1986);
and U3463 (N_3463,N_2474,N_2999);
nor U3464 (N_3464,N_2434,N_234);
or U3465 (N_3465,N_511,N_205);
nor U3466 (N_3466,N_1475,N_598);
or U3467 (N_3467,N_2035,N_670);
xor U3468 (N_3468,N_245,N_2716);
nor U3469 (N_3469,N_1518,N_1720);
xor U3470 (N_3470,N_2865,N_445);
or U3471 (N_3471,N_2669,N_755);
and U3472 (N_3472,N_928,N_704);
nand U3473 (N_3473,N_1108,N_1821);
nor U3474 (N_3474,N_815,N_2311);
nand U3475 (N_3475,N_2493,N_2122);
xnor U3476 (N_3476,N_2781,N_1301);
and U3477 (N_3477,N_1715,N_2012);
or U3478 (N_3478,N_1570,N_2362);
nor U3479 (N_3479,N_2134,N_1311);
nand U3480 (N_3480,N_1635,N_2438);
nor U3481 (N_3481,N_499,N_740);
nand U3482 (N_3482,N_44,N_2905);
nand U3483 (N_3483,N_2486,N_231);
xor U3484 (N_3484,N_1771,N_1835);
nor U3485 (N_3485,N_2644,N_2707);
or U3486 (N_3486,N_2067,N_416);
or U3487 (N_3487,N_1671,N_2661);
nor U3488 (N_3488,N_736,N_2348);
nand U3489 (N_3489,N_1048,N_1968);
or U3490 (N_3490,N_36,N_746);
nand U3491 (N_3491,N_2340,N_258);
and U3492 (N_3492,N_1372,N_2622);
nor U3493 (N_3493,N_2787,N_2023);
and U3494 (N_3494,N_2704,N_802);
xor U3495 (N_3495,N_2369,N_421);
and U3496 (N_3496,N_1050,N_2537);
or U3497 (N_3497,N_936,N_962);
nor U3498 (N_3498,N_2768,N_756);
and U3499 (N_3499,N_2521,N_1071);
and U3500 (N_3500,N_2061,N_262);
nand U3501 (N_3501,N_687,N_2499);
or U3502 (N_3502,N_1404,N_2276);
or U3503 (N_3503,N_2198,N_484);
nor U3504 (N_3504,N_340,N_1441);
or U3505 (N_3505,N_27,N_165);
or U3506 (N_3506,N_1648,N_2747);
nor U3507 (N_3507,N_885,N_260);
and U3508 (N_3508,N_2309,N_2186);
and U3509 (N_3509,N_1293,N_1481);
or U3510 (N_3510,N_1974,N_344);
nor U3511 (N_3511,N_995,N_1642);
xor U3512 (N_3512,N_367,N_1034);
nand U3513 (N_3513,N_1693,N_2456);
or U3514 (N_3514,N_884,N_252);
or U3515 (N_3515,N_2812,N_1673);
nor U3516 (N_3516,N_2950,N_1978);
or U3517 (N_3517,N_1923,N_2147);
or U3518 (N_3518,N_565,N_2248);
xnor U3519 (N_3519,N_2420,N_540);
nand U3520 (N_3520,N_1375,N_2611);
and U3521 (N_3521,N_2821,N_2353);
or U3522 (N_3522,N_1553,N_454);
or U3523 (N_3523,N_1442,N_92);
nand U3524 (N_3524,N_1960,N_2743);
or U3525 (N_3525,N_2453,N_810);
or U3526 (N_3526,N_2299,N_304);
xnor U3527 (N_3527,N_381,N_2307);
and U3528 (N_3528,N_848,N_385);
or U3529 (N_3529,N_2744,N_2568);
nand U3530 (N_3530,N_1111,N_835);
or U3531 (N_3531,N_935,N_2001);
and U3532 (N_3532,N_519,N_1806);
xnor U3533 (N_3533,N_25,N_1328);
or U3534 (N_3534,N_978,N_1542);
and U3535 (N_3535,N_1044,N_1408);
nor U3536 (N_3536,N_2312,N_597);
nand U3537 (N_3537,N_2145,N_1405);
nor U3538 (N_3538,N_749,N_526);
nor U3539 (N_3539,N_2215,N_768);
or U3540 (N_3540,N_1956,N_1001);
nor U3541 (N_3541,N_1760,N_418);
and U3542 (N_3542,N_214,N_1437);
or U3543 (N_3543,N_1737,N_1273);
xor U3544 (N_3544,N_2436,N_1763);
nand U3545 (N_3545,N_382,N_737);
nor U3546 (N_3546,N_577,N_106);
or U3547 (N_3547,N_1337,N_1927);
nand U3548 (N_3548,N_651,N_2361);
nor U3549 (N_3549,N_1597,N_1879);
and U3550 (N_3550,N_266,N_225);
and U3551 (N_3551,N_547,N_1321);
or U3552 (N_3552,N_1810,N_1157);
nand U3553 (N_3553,N_2167,N_2000);
and U3554 (N_3554,N_219,N_1701);
xnor U3555 (N_3555,N_587,N_1887);
nor U3556 (N_3556,N_2400,N_2038);
or U3557 (N_3557,N_774,N_2036);
or U3558 (N_3558,N_934,N_2405);
nand U3559 (N_3559,N_2277,N_761);
nor U3560 (N_3560,N_1944,N_1203);
nor U3561 (N_3561,N_2670,N_2554);
xnor U3562 (N_3562,N_646,N_293);
nand U3563 (N_3563,N_1783,N_787);
nand U3564 (N_3564,N_1613,N_2727);
nand U3565 (N_3565,N_1523,N_1402);
xor U3566 (N_3566,N_626,N_999);
nor U3567 (N_3567,N_759,N_2922);
nand U3568 (N_3568,N_1877,N_397);
or U3569 (N_3569,N_78,N_1501);
nand U3570 (N_3570,N_735,N_1917);
or U3571 (N_3571,N_2784,N_1675);
nor U3572 (N_3572,N_411,N_2246);
nor U3573 (N_3573,N_270,N_2188);
and U3574 (N_3574,N_1227,N_1655);
or U3575 (N_3575,N_1384,N_378);
nand U3576 (N_3576,N_808,N_919);
nor U3577 (N_3577,N_1999,N_640);
nand U3578 (N_3578,N_1966,N_2709);
nor U3579 (N_3579,N_1992,N_1036);
nor U3580 (N_3580,N_4,N_486);
nor U3581 (N_3581,N_2918,N_1370);
xor U3582 (N_3582,N_960,N_471);
xnor U3583 (N_3583,N_650,N_760);
nand U3584 (N_3584,N_980,N_1452);
xnor U3585 (N_3585,N_1716,N_2583);
nor U3586 (N_3586,N_2208,N_2845);
or U3587 (N_3587,N_2176,N_286);
nor U3588 (N_3588,N_2385,N_337);
nor U3589 (N_3589,N_1317,N_2473);
nand U3590 (N_3590,N_291,N_396);
nand U3591 (N_3591,N_1304,N_2256);
xor U3592 (N_3592,N_949,N_1981);
and U3593 (N_3593,N_1112,N_2152);
xor U3594 (N_3594,N_2532,N_662);
nor U3595 (N_3595,N_1288,N_1136);
xor U3596 (N_3596,N_2721,N_2060);
nor U3597 (N_3597,N_1726,N_1484);
nor U3598 (N_3598,N_2980,N_1947);
and U3599 (N_3599,N_346,N_2303);
nor U3600 (N_3600,N_1808,N_100);
or U3601 (N_3601,N_2658,N_153);
nand U3602 (N_3602,N_2591,N_1315);
and U3603 (N_3603,N_1016,N_2690);
or U3604 (N_3604,N_544,N_1825);
and U3605 (N_3605,N_2724,N_2685);
nand U3606 (N_3606,N_1502,N_1544);
and U3607 (N_3607,N_182,N_2616);
nand U3608 (N_3608,N_732,N_2801);
nand U3609 (N_3609,N_1368,N_983);
and U3610 (N_3610,N_858,N_2915);
or U3611 (N_3611,N_2213,N_2976);
and U3612 (N_3612,N_2171,N_2391);
nand U3613 (N_3613,N_2241,N_138);
or U3614 (N_3614,N_1732,N_1554);
xor U3615 (N_3615,N_2941,N_2737);
or U3616 (N_3616,N_1496,N_362);
and U3617 (N_3617,N_2656,N_2867);
nand U3618 (N_3618,N_2965,N_410);
or U3619 (N_3619,N_2139,N_2243);
or U3620 (N_3620,N_495,N_2935);
xnor U3621 (N_3621,N_178,N_1522);
and U3622 (N_3622,N_615,N_1512);
nand U3623 (N_3623,N_2072,N_2639);
xor U3624 (N_3624,N_267,N_419);
nand U3625 (N_3625,N_166,N_567);
xor U3626 (N_3626,N_6,N_1804);
nor U3627 (N_3627,N_247,N_287);
or U3628 (N_3628,N_1455,N_548);
nand U3629 (N_3629,N_2803,N_176);
or U3630 (N_3630,N_263,N_2300);
or U3631 (N_3631,N_890,N_1742);
xnor U3632 (N_3632,N_1848,N_1246);
nor U3633 (N_3633,N_2883,N_1224);
nor U3634 (N_3634,N_1755,N_2975);
or U3635 (N_3635,N_898,N_2032);
xnor U3636 (N_3636,N_472,N_930);
nor U3637 (N_3637,N_2563,N_2212);
nor U3638 (N_3638,N_864,N_1110);
nand U3639 (N_3639,N_32,N_566);
and U3640 (N_3640,N_1795,N_1951);
and U3641 (N_3641,N_2633,N_322);
xnor U3642 (N_3642,N_2221,N_2586);
and U3643 (N_3643,N_2082,N_154);
nand U3644 (N_3644,N_2103,N_188);
or U3645 (N_3645,N_785,N_86);
xnor U3646 (N_3646,N_101,N_656);
or U3647 (N_3647,N_2758,N_91);
nand U3648 (N_3648,N_283,N_1593);
and U3649 (N_3649,N_487,N_1678);
xor U3650 (N_3650,N_2963,N_839);
nor U3651 (N_3651,N_593,N_2715);
and U3652 (N_3652,N_2534,N_1058);
nand U3653 (N_3653,N_2410,N_1664);
and U3654 (N_3654,N_2084,N_1432);
xnor U3655 (N_3655,N_1443,N_2077);
and U3656 (N_3656,N_946,N_1661);
or U3657 (N_3657,N_2272,N_893);
nor U3658 (N_3658,N_8,N_398);
or U3659 (N_3659,N_2355,N_2200);
nand U3660 (N_3660,N_945,N_2700);
xnor U3661 (N_3661,N_1989,N_158);
or U3662 (N_3662,N_2123,N_1092);
xor U3663 (N_3663,N_265,N_77);
xor U3664 (N_3664,N_2753,N_2245);
xor U3665 (N_3665,N_23,N_251);
nand U3666 (N_3666,N_793,N_1260);
and U3667 (N_3667,N_2366,N_1449);
nand U3668 (N_3668,N_498,N_1777);
and U3669 (N_3669,N_1012,N_631);
or U3670 (N_3670,N_2512,N_2839);
nand U3671 (N_3671,N_2347,N_976);
nand U3672 (N_3672,N_2321,N_1253);
nor U3673 (N_3673,N_1906,N_2949);
xnor U3674 (N_3674,N_622,N_2726);
xnor U3675 (N_3675,N_634,N_2401);
and U3676 (N_3676,N_1849,N_503);
and U3677 (N_3677,N_974,N_15);
xnor U3678 (N_3678,N_128,N_681);
xnor U3679 (N_3679,N_2705,N_2331);
xnor U3680 (N_3680,N_2247,N_987);
nor U3681 (N_3681,N_979,N_1473);
and U3682 (N_3682,N_1787,N_2629);
or U3683 (N_3683,N_420,N_2985);
and U3684 (N_3684,N_437,N_876);
xor U3685 (N_3685,N_882,N_1520);
xor U3686 (N_3686,N_62,N_2637);
and U3687 (N_3687,N_2849,N_2954);
nand U3688 (N_3688,N_702,N_2713);
nand U3689 (N_3689,N_2802,N_1271);
or U3690 (N_3690,N_583,N_2190);
and U3691 (N_3691,N_1324,N_2446);
or U3692 (N_3692,N_2140,N_298);
xor U3693 (N_3693,N_816,N_2835);
and U3694 (N_3694,N_1219,N_1894);
or U3695 (N_3695,N_715,N_2648);
nand U3696 (N_3696,N_2587,N_1669);
nand U3697 (N_3697,N_2960,N_2177);
and U3698 (N_3698,N_2408,N_2010);
or U3699 (N_3699,N_2651,N_2874);
nor U3700 (N_3700,N_1210,N_492);
and U3701 (N_3701,N_982,N_2511);
or U3702 (N_3702,N_799,N_392);
and U3703 (N_3703,N_444,N_927);
and U3704 (N_3704,N_1792,N_838);
xor U3705 (N_3705,N_538,N_2161);
nor U3706 (N_3706,N_1188,N_1666);
nand U3707 (N_3707,N_1093,N_620);
nand U3708 (N_3708,N_941,N_603);
and U3709 (N_3709,N_842,N_2441);
xnor U3710 (N_3710,N_2268,N_2930);
or U3711 (N_3711,N_406,N_502);
or U3712 (N_3712,N_990,N_1223);
nor U3713 (N_3713,N_2741,N_2594);
and U3714 (N_3714,N_1721,N_16);
nor U3715 (N_3715,N_1859,N_1852);
nor U3716 (N_3716,N_2748,N_1545);
nor U3717 (N_3717,N_1504,N_65);
nand U3718 (N_3718,N_2663,N_827);
nand U3719 (N_3719,N_2230,N_2287);
or U3720 (N_3720,N_2800,N_191);
nand U3721 (N_3721,N_1541,N_1213);
nor U3722 (N_3722,N_623,N_2326);
nor U3723 (N_3723,N_1128,N_2196);
or U3724 (N_3724,N_1327,N_703);
xnor U3725 (N_3725,N_1230,N_690);
and U3726 (N_3726,N_2323,N_2964);
xor U3727 (N_3727,N_2497,N_427);
nor U3728 (N_3728,N_1908,N_1695);
xnor U3729 (N_3729,N_496,N_531);
nor U3730 (N_3730,N_1957,N_2869);
nor U3731 (N_3731,N_361,N_1428);
and U3732 (N_3732,N_2793,N_2646);
nand U3733 (N_3733,N_2352,N_2961);
or U3734 (N_3734,N_1707,N_1084);
nor U3735 (N_3735,N_347,N_664);
nor U3736 (N_3736,N_470,N_31);
nand U3737 (N_3737,N_1123,N_2195);
nor U3738 (N_3738,N_2003,N_2947);
xor U3739 (N_3739,N_1928,N_2943);
xnor U3740 (N_3740,N_1234,N_447);
nand U3741 (N_3741,N_2701,N_1214);
and U3742 (N_3742,N_1608,N_2159);
xnor U3743 (N_3743,N_1623,N_1440);
and U3744 (N_3744,N_2955,N_1352);
or U3745 (N_3745,N_2328,N_271);
or U3746 (N_3746,N_1823,N_1319);
xor U3747 (N_3747,N_1381,N_428);
nand U3748 (N_3748,N_1662,N_206);
xnor U3749 (N_3749,N_1433,N_2108);
and U3750 (N_3750,N_2510,N_2876);
nand U3751 (N_3751,N_1982,N_2503);
and U3752 (N_3752,N_2529,N_2649);
and U3753 (N_3753,N_955,N_2259);
xnor U3754 (N_3754,N_173,N_2601);
nand U3755 (N_3755,N_2861,N_308);
nor U3756 (N_3756,N_2764,N_199);
nor U3757 (N_3757,N_1153,N_1156);
or U3758 (N_3758,N_1953,N_1383);
and U3759 (N_3759,N_1325,N_1008);
nor U3760 (N_3760,N_1621,N_379);
nor U3761 (N_3761,N_921,N_728);
nor U3762 (N_3762,N_912,N_213);
and U3763 (N_3763,N_211,N_1166);
nor U3764 (N_3764,N_1769,N_1099);
nand U3765 (N_3765,N_2495,N_870);
and U3766 (N_3766,N_2458,N_2522);
or U3767 (N_3767,N_1039,N_2181);
nor U3768 (N_3768,N_2797,N_1898);
and U3769 (N_3769,N_1790,N_2983);
nor U3770 (N_3770,N_2635,N_462);
nand U3771 (N_3771,N_2775,N_2015);
nand U3772 (N_3772,N_1516,N_1983);
nor U3773 (N_3773,N_125,N_1765);
and U3774 (N_3774,N_2316,N_2058);
nor U3775 (N_3775,N_2872,N_1883);
xnor U3776 (N_3776,N_2217,N_289);
or U3777 (N_3777,N_2153,N_226);
nor U3778 (N_3778,N_1833,N_1864);
and U3779 (N_3779,N_1132,N_747);
xnor U3780 (N_3780,N_2232,N_776);
and U3781 (N_3781,N_2571,N_2820);
and U3782 (N_3782,N_1320,N_1839);
nand U3783 (N_3783,N_973,N_1495);
or U3784 (N_3784,N_873,N_1365);
nand U3785 (N_3785,N_2509,N_1438);
or U3786 (N_3786,N_592,N_594);
or U3787 (N_3787,N_600,N_2595);
nor U3788 (N_3788,N_21,N_922);
nor U3789 (N_3789,N_2813,N_1469);
nor U3790 (N_3790,N_1711,N_168);
xor U3791 (N_3791,N_301,N_2929);
and U3792 (N_3792,N_1129,N_1889);
xor U3793 (N_3793,N_2936,N_2034);
nor U3794 (N_3794,N_2580,N_1647);
xor U3795 (N_3795,N_1359,N_223);
nand U3796 (N_3796,N_971,N_1170);
nand U3797 (N_3797,N_1033,N_931);
nand U3798 (N_3798,N_1207,N_607);
or U3799 (N_3799,N_1942,N_2547);
xor U3800 (N_3800,N_1019,N_468);
nand U3801 (N_3801,N_2903,N_1905);
xnor U3802 (N_3802,N_2652,N_254);
nand U3803 (N_3803,N_1143,N_2027);
nand U3804 (N_3804,N_1200,N_2402);
or U3805 (N_3805,N_423,N_2919);
nand U3806 (N_3806,N_798,N_1413);
and U3807 (N_3807,N_2973,N_1548);
nand U3808 (N_3808,N_2150,N_1866);
nand U3809 (N_3809,N_1279,N_222);
xor U3810 (N_3810,N_2933,N_300);
nor U3811 (N_3811,N_2389,N_2165);
nor U3812 (N_3812,N_645,N_2860);
nor U3813 (N_3813,N_2137,N_865);
and U3814 (N_3814,N_1712,N_2229);
xnor U3815 (N_3815,N_180,N_353);
and U3816 (N_3816,N_910,N_2608);
nor U3817 (N_3817,N_2628,N_564);
and U3818 (N_3818,N_1256,N_542);
xnor U3819 (N_3819,N_814,N_992);
xor U3820 (N_3820,N_845,N_1692);
or U3821 (N_3821,N_947,N_2251);
and U3822 (N_3822,N_2107,N_1809);
and U3823 (N_3823,N_157,N_463);
nor U3824 (N_3824,N_847,N_2610);
or U3825 (N_3825,N_706,N_331);
xor U3826 (N_3826,N_1638,N_2128);
or U3827 (N_3827,N_359,N_52);
and U3828 (N_3828,N_1150,N_175);
nor U3829 (N_3829,N_458,N_1387);
nand U3830 (N_3830,N_2469,N_1225);
nand U3831 (N_3831,N_2343,N_1994);
or U3832 (N_3832,N_2506,N_1424);
nand U3833 (N_3833,N_2977,N_834);
xor U3834 (N_3834,N_2334,N_2851);
nand U3835 (N_3835,N_1577,N_1248);
or U3836 (N_3836,N_1948,N_2517);
and U3837 (N_3837,N_2124,N_343);
nor U3838 (N_3838,N_966,N_1165);
and U3839 (N_3839,N_1182,N_2630);
xnor U3840 (N_3840,N_627,N_539);
nand U3841 (N_3841,N_879,N_2745);
nand U3842 (N_3842,N_1801,N_383);
nand U3843 (N_3843,N_1294,N_2351);
nor U3844 (N_3844,N_1582,N_2097);
xor U3845 (N_3845,N_2884,N_1997);
or U3846 (N_3846,N_2313,N_2255);
and U3847 (N_3847,N_1181,N_1220);
nor U3848 (N_3848,N_72,N_1274);
nor U3849 (N_3849,N_434,N_788);
nor U3850 (N_3850,N_1513,N_374);
nand U3851 (N_3851,N_2557,N_228);
or U3852 (N_3852,N_2624,N_2819);
or U3853 (N_3853,N_2548,N_197);
xnor U3854 (N_3854,N_2780,N_1650);
xnor U3855 (N_3855,N_784,N_1263);
xnor U3856 (N_3856,N_2948,N_968);
xor U3857 (N_3857,N_916,N_2155);
xnor U3858 (N_3858,N_2900,N_648);
nand U3859 (N_3859,N_2048,N_1488);
nand U3860 (N_3860,N_2735,N_2214);
nor U3861 (N_3861,N_556,N_1453);
nor U3862 (N_3862,N_2315,N_1788);
xor U3863 (N_3863,N_1341,N_2856);
nor U3864 (N_3864,N_208,N_924);
xnor U3865 (N_3865,N_1607,N_60);
xor U3866 (N_3866,N_1146,N_2460);
nor U3867 (N_3867,N_606,N_1844);
and U3868 (N_3868,N_1113,N_2734);
or U3869 (N_3869,N_771,N_2083);
and U3870 (N_3870,N_1764,N_986);
or U3871 (N_3871,N_370,N_943);
and U3872 (N_3872,N_621,N_991);
nor U3873 (N_3873,N_334,N_387);
nor U3874 (N_3874,N_1485,N_220);
and U3875 (N_3875,N_143,N_1696);
and U3876 (N_3876,N_1454,N_1215);
nor U3877 (N_3877,N_2736,N_235);
and U3878 (N_3878,N_515,N_2044);
and U3879 (N_3879,N_1478,N_87);
nand U3880 (N_3880,N_993,N_2384);
and U3881 (N_3881,N_1639,N_1252);
xor U3882 (N_3882,N_2056,N_1121);
or U3883 (N_3883,N_752,N_2879);
or U3884 (N_3884,N_1656,N_1875);
nor U3885 (N_3885,N_1037,N_190);
nand U3886 (N_3886,N_958,N_1719);
nor U3887 (N_3887,N_1703,N_169);
or U3888 (N_3888,N_276,N_2979);
and U3889 (N_3889,N_2913,N_2443);
nor U3890 (N_3890,N_2262,N_1024);
and U3891 (N_3891,N_2118,N_2105);
and U3892 (N_3892,N_489,N_779);
xor U3893 (N_3893,N_99,N_2934);
xnor U3894 (N_3894,N_2471,N_2527);
nor U3895 (N_3895,N_1091,N_195);
xnor U3896 (N_3896,N_2899,N_1587);
nor U3897 (N_3897,N_889,N_2926);
and U3898 (N_3898,N_2104,N_1973);
xnor U3899 (N_3899,N_2496,N_1296);
and U3900 (N_3900,N_2057,N_1307);
nor U3901 (N_3901,N_2558,N_442);
or U3902 (N_3902,N_2555,N_1625);
nand U3903 (N_3903,N_2430,N_19);
nor U3904 (N_3904,N_831,N_1401);
nand U3905 (N_3905,N_1838,N_2101);
and U3906 (N_3906,N_2805,N_2019);
nor U3907 (N_3907,N_121,N_2127);
or U3908 (N_3908,N_1386,N_1920);
xor U3909 (N_3909,N_2451,N_2286);
or U3910 (N_3910,N_2004,N_2314);
or U3911 (N_3911,N_2380,N_844);
or U3912 (N_3912,N_2046,N_2168);
and U3913 (N_3913,N_497,N_1780);
xor U3914 (N_3914,N_1710,N_1872);
and U3915 (N_3915,N_2677,N_2885);
nand U3916 (N_3916,N_1874,N_118);
nand U3917 (N_3917,N_243,N_1893);
nand U3918 (N_3918,N_1557,N_1896);
or U3919 (N_3919,N_2841,N_1070);
nand U3920 (N_3920,N_714,N_789);
nand U3921 (N_3921,N_412,N_2333);
or U3922 (N_3922,N_2539,N_773);
nor U3923 (N_3923,N_1980,N_1377);
or U3924 (N_3924,N_1629,N_914);
nand U3925 (N_3925,N_2786,N_1420);
nand U3926 (N_3926,N_2795,N_2284);
nand U3927 (N_3927,N_1911,N_1679);
and U3928 (N_3928,N_1125,N_2421);
xnor U3929 (N_3929,N_1924,N_1514);
nand U3930 (N_3930,N_2518,N_81);
or U3931 (N_3931,N_2588,N_192);
or U3932 (N_3932,N_661,N_891);
xor U3933 (N_3933,N_725,N_2814);
or U3934 (N_3934,N_1080,N_323);
and U3935 (N_3935,N_2796,N_1878);
xor U3936 (N_3936,N_765,N_217);
nor U3937 (N_3937,N_2095,N_482);
nand U3938 (N_3938,N_2638,N_2106);
or U3939 (N_3939,N_227,N_1127);
xor U3940 (N_3940,N_2025,N_1312);
nor U3941 (N_3941,N_514,N_1373);
or U3942 (N_3942,N_184,N_1837);
nor U3943 (N_3943,N_2092,N_1668);
nor U3944 (N_3944,N_688,N_314);
or U3945 (N_3945,N_969,N_2822);
nand U3946 (N_3946,N_580,N_2113);
or U3947 (N_3947,N_2358,N_319);
nor U3948 (N_3948,N_1677,N_179);
xnor U3949 (N_3949,N_1429,N_2953);
or U3950 (N_3950,N_2225,N_2516);
nor U3951 (N_3951,N_2792,N_2889);
nand U3952 (N_3952,N_1026,N_1697);
nand U3953 (N_3953,N_7,N_1376);
nor U3954 (N_3954,N_2206,N_1843);
xor U3955 (N_3955,N_1899,N_1868);
nand U3956 (N_3956,N_79,N_2179);
or U3957 (N_3957,N_295,N_2080);
and U3958 (N_3958,N_797,N_452);
xor U3959 (N_3959,N_1258,N_69);
or U3960 (N_3960,N_809,N_611);
xnor U3961 (N_3961,N_2031,N_2100);
nand U3962 (N_3962,N_1709,N_2089);
and U3963 (N_3963,N_1641,N_1571);
xor U3964 (N_3964,N_2671,N_1118);
or U3965 (N_3965,N_2942,N_277);
and U3966 (N_3966,N_2993,N_1435);
nand U3967 (N_3967,N_2204,N_1117);
nand U3968 (N_3968,N_70,N_1556);
nor U3969 (N_3969,N_181,N_395);
xnor U3970 (N_3970,N_141,N_1789);
xor U3971 (N_3971,N_204,N_1000);
and U3972 (N_3972,N_2289,N_1105);
or U3973 (N_3973,N_574,N_2565);
and U3974 (N_3974,N_2544,N_2891);
and U3975 (N_3975,N_2621,N_1144);
xnor U3976 (N_3976,N_2263,N_2904);
nor U3977 (N_3977,N_1088,N_2373);
xnor U3978 (N_3978,N_1581,N_103);
and U3979 (N_3979,N_2788,N_167);
and U3980 (N_3980,N_790,N_2055);
or U3981 (N_3981,N_1714,N_2201);
xnor U3982 (N_3982,N_2282,N_1406);
and U3983 (N_3983,N_1272,N_698);
nor U3984 (N_3984,N_480,N_654);
nor U3985 (N_3985,N_1276,N_1551);
or U3986 (N_3986,N_2202,N_1247);
or U3987 (N_3987,N_97,N_1842);
and U3988 (N_3988,N_1916,N_2297);
and U3989 (N_3989,N_1097,N_1681);
nor U3990 (N_3990,N_1119,N_465);
nand U3991 (N_3991,N_2605,N_1098);
xor U3992 (N_3992,N_1725,N_2372);
nor U3993 (N_3993,N_1564,N_2059);
xor U3994 (N_3994,N_1351,N_1694);
and U3995 (N_3995,N_1445,N_1772);
nor U3996 (N_3996,N_1082,N_1306);
nor U3997 (N_3997,N_1758,N_1345);
nor U3998 (N_3998,N_2504,N_1909);
xor U3999 (N_3999,N_2109,N_731);
or U4000 (N_4000,N_1267,N_1023);
or U4001 (N_4001,N_508,N_2483);
and U4002 (N_4002,N_1946,N_1531);
nand U4003 (N_4003,N_280,N_2381);
nand U4004 (N_4004,N_2662,N_325);
or U4005 (N_4005,N_576,N_1528);
nand U4006 (N_4006,N_38,N_697);
nand U4007 (N_4007,N_723,N_1025);
xor U4008 (N_4008,N_972,N_711);
and U4009 (N_4009,N_41,N_2575);
nor U4010 (N_4010,N_2946,N_1416);
nand U4011 (N_4011,N_813,N_10);
nand U4012 (N_4012,N_2462,N_352);
and U4013 (N_4013,N_915,N_2183);
nor U4014 (N_4014,N_1886,N_1740);
and U4015 (N_4015,N_1005,N_1633);
nor U4016 (N_4016,N_2488,N_131);
and U4017 (N_4017,N_2808,N_439);
or U4018 (N_4018,N_533,N_733);
nand U4019 (N_4019,N_883,N_73);
or U4020 (N_4020,N_1096,N_1237);
nand U4021 (N_4021,N_869,N_792);
xnor U4022 (N_4022,N_2075,N_1072);
nor U4023 (N_4023,N_1853,N_2581);
and U4024 (N_4024,N_832,N_2766);
and U4025 (N_4025,N_1222,N_2310);
xor U4026 (N_4026,N_717,N_2143);
nand U4027 (N_4027,N_1934,N_2050);
nor U4028 (N_4028,N_653,N_887);
and U4029 (N_4029,N_363,N_2604);
or U4030 (N_4030,N_1472,N_1251);
nor U4031 (N_4031,N_2081,N_432);
xnor U4032 (N_4032,N_1180,N_1793);
or U4033 (N_4033,N_1186,N_1095);
and U4034 (N_4034,N_680,N_1490);
and U4035 (N_4035,N_1239,N_2718);
nor U4036 (N_4036,N_975,N_2647);
and U4037 (N_4037,N_2335,N_18);
nand U4038 (N_4038,N_2125,N_1706);
nor U4039 (N_4039,N_1840,N_1724);
nor U4040 (N_4040,N_1546,N_2185);
and U4041 (N_4041,N_1759,N_2382);
or U4042 (N_4042,N_501,N_281);
or U4043 (N_4043,N_1450,N_629);
nor U4044 (N_4044,N_1831,N_2398);
and U4045 (N_4045,N_1163,N_2564);
nand U4046 (N_4046,N_2749,N_2773);
or U4047 (N_4047,N_1369,N_743);
nand U4048 (N_4048,N_2545,N_2135);
and U4049 (N_4049,N_1915,N_1407);
and U4050 (N_4050,N_345,N_156);
and U4051 (N_4051,N_830,N_2755);
xnor U4052 (N_4052,N_1689,N_1798);
xor U4053 (N_4053,N_1996,N_2099);
xnor U4054 (N_4054,N_1259,N_2187);
xor U4055 (N_4055,N_1718,N_2546);
and U4056 (N_4056,N_896,N_965);
nand U4057 (N_4057,N_2523,N_2093);
nand U4058 (N_4058,N_2156,N_683);
or U4059 (N_4059,N_1979,N_1184);
xnor U4060 (N_4060,N_2477,N_1628);
nand U4061 (N_4061,N_2750,N_590);
nand U4062 (N_4062,N_507,N_918);
nor U4063 (N_4063,N_2689,N_2386);
or U4064 (N_4064,N_636,N_297);
xor U4065 (N_4065,N_1043,N_1149);
and U4066 (N_4066,N_1040,N_409);
nand U4067 (N_4067,N_727,N_1003);
nor U4068 (N_4068,N_630,N_2698);
xnor U4069 (N_4069,N_1601,N_795);
nor U4070 (N_4070,N_523,N_1465);
xor U4071 (N_4071,N_1626,N_2291);
and U4072 (N_4072,N_1168,N_1585);
xnor U4073 (N_4073,N_888,N_1754);
and U4074 (N_4074,N_920,N_253);
or U4075 (N_4075,N_2160,N_1415);
nand U4076 (N_4076,N_2008,N_2553);
nand U4077 (N_4077,N_1884,N_691);
and U4078 (N_4078,N_2073,N_1566);
or U4079 (N_4079,N_1499,N_1120);
and U4080 (N_4080,N_2777,N_1068);
nand U4081 (N_4081,N_2678,N_875);
nand U4082 (N_4082,N_578,N_2890);
nand U4083 (N_4083,N_2087,N_1041);
nor U4084 (N_4084,N_846,N_2346);
and U4085 (N_4085,N_2418,N_2054);
nand U4086 (N_4086,N_2561,N_2978);
nand U4087 (N_4087,N_1651,N_903);
and U4088 (N_4088,N_61,N_1487);
or U4089 (N_4089,N_2290,N_961);
nor U4090 (N_4090,N_529,N_712);
or U4091 (N_4091,N_2367,N_200);
nor U4092 (N_4092,N_852,N_2240);
nand U4093 (N_4093,N_917,N_504);
nor U4094 (N_4094,N_682,N_1439);
or U4095 (N_4095,N_2375,N_2893);
nor U4096 (N_4096,N_229,N_1175);
nand U4097 (N_4097,N_348,N_1171);
nand U4098 (N_4098,N_1329,N_183);
and U4099 (N_4099,N_860,N_959);
and U4100 (N_4100,N_2770,N_1155);
or U4101 (N_4101,N_655,N_264);
xnor U4102 (N_4102,N_2844,N_424);
nand U4103 (N_4103,N_1687,N_455);
or U4104 (N_4104,N_2833,N_1029);
and U4105 (N_4105,N_2219,N_1646);
xor U4106 (N_4106,N_520,N_54);
nor U4107 (N_4107,N_2765,N_24);
nand U4108 (N_4108,N_2275,N_310);
and U4109 (N_4109,N_55,N_305);
xnor U4110 (N_4110,N_2390,N_812);
nor U4111 (N_4111,N_1653,N_350);
nand U4112 (N_4112,N_1936,N_2009);
and U4113 (N_4113,N_2940,N_59);
nor U4114 (N_4114,N_2329,N_652);
and U4115 (N_4115,N_1775,N_2931);
or U4116 (N_4116,N_2182,N_1083);
xor U4117 (N_4117,N_1665,N_1952);
and U4118 (N_4118,N_2220,N_1708);
and U4119 (N_4119,N_1277,N_2368);
xor U4120 (N_4120,N_2920,N_174);
xor U4121 (N_4121,N_791,N_767);
and U4122 (N_4122,N_307,N_1828);
and U4123 (N_4123,N_1537,N_2871);
nand U4124 (N_4124,N_1049,N_748);
or U4125 (N_4125,N_855,N_2778);
and U4126 (N_4126,N_299,N_892);
or U4127 (N_4127,N_230,N_822);
nand U4128 (N_4128,N_1018,N_1609);
nand U4129 (N_4129,N_275,N_1527);
nor U4130 (N_4130,N_2578,N_1578);
nor U4131 (N_4131,N_272,N_2714);
nand U4132 (N_4132,N_324,N_2325);
xnor U4133 (N_4133,N_1841,N_172);
and U4134 (N_4134,N_1066,N_2829);
and U4135 (N_4135,N_1431,N_1079);
nor U4136 (N_4136,N_1768,N_1081);
and U4137 (N_4137,N_365,N_446);
nor U4138 (N_4138,N_2192,N_907);
xnor U4139 (N_4139,N_1856,N_2664);
and U4140 (N_4140,N_2533,N_2102);
or U4141 (N_4141,N_2210,N_1670);
nand U4142 (N_4142,N_745,N_758);
xor U4143 (N_4143,N_107,N_1285);
or U4144 (N_4144,N_1969,N_114);
nor U4145 (N_4145,N_2738,N_1463);
xnor U4146 (N_4146,N_569,N_937);
nand U4147 (N_4147,N_2465,N_2746);
nor U4148 (N_4148,N_2111,N_1355);
nand U4149 (N_4149,N_2790,N_134);
nand U4150 (N_4150,N_638,N_42);
nand U4151 (N_4151,N_1534,N_2864);
and U4152 (N_4152,N_1183,N_617);
xor U4153 (N_4153,N_1204,N_938);
nand U4154 (N_4154,N_5,N_1907);
xor U4155 (N_4155,N_2002,N_2552);
nor U4156 (N_4156,N_895,N_2349);
nand U4157 (N_4157,N_2525,N_338);
nand U4158 (N_4158,N_2655,N_356);
xor U4159 (N_4159,N_2513,N_2772);
nand U4160 (N_4160,N_1631,N_1266);
nor U4161 (N_4161,N_1382,N_2170);
or U4162 (N_4162,N_1736,N_1038);
or U4163 (N_4163,N_3,N_2403);
nor U4164 (N_4164,N_1206,N_1241);
or U4165 (N_4165,N_998,N_1264);
and U4166 (N_4166,N_618,N_2791);
xor U4167 (N_4167,N_2199,N_2567);
xnor U4168 (N_4168,N_868,N_1744);
and U4169 (N_4169,N_2631,N_713);
and U4170 (N_4170,N_2485,N_2843);
xor U4171 (N_4171,N_2041,N_1727);
nor U4172 (N_4172,N_1169,N_1939);
and U4173 (N_4173,N_33,N_1343);
and U4174 (N_4174,N_2751,N_2613);
nand U4175 (N_4175,N_2722,N_2692);
and U4176 (N_4176,N_1659,N_139);
xnor U4177 (N_4177,N_775,N_1561);
and U4178 (N_4178,N_58,N_2416);
nand U4179 (N_4179,N_1657,N_2174);
xnor U4180 (N_4180,N_441,N_1560);
xor U4181 (N_4181,N_80,N_335);
or U4182 (N_4182,N_2804,N_1255);
xor U4183 (N_4183,N_1031,N_2356);
or U4184 (N_4184,N_221,N_2541);
nor U4185 (N_4185,N_1278,N_20);
xor U4186 (N_4186,N_881,N_2392);
and U4187 (N_4187,N_660,N_2694);
or U4188 (N_4188,N_796,N_261);
and U4189 (N_4189,N_1559,N_2180);
and U4190 (N_4190,N_1691,N_1154);
xnor U4191 (N_4191,N_2428,N_2442);
or U4192 (N_4192,N_285,N_39);
nand U4193 (N_4193,N_619,N_342);
and U4194 (N_4194,N_2914,N_824);
or U4195 (N_4195,N_1854,N_537);
or U4196 (N_4196,N_1030,N_985);
xor U4197 (N_4197,N_693,N_0);
nor U4198 (N_4198,N_1871,N_1933);
nor U4199 (N_4199,N_1212,N_1943);
or U4200 (N_4200,N_83,N_242);
xor U4201 (N_4201,N_1932,N_1065);
nor U4202 (N_4202,N_90,N_2505);
xnor U4203 (N_4203,N_1643,N_1471);
xor U4204 (N_4204,N_2197,N_2811);
nor U4205 (N_4205,N_1464,N_105);
xnor U4206 (N_4206,N_255,N_435);
nor U4207 (N_4207,N_807,N_861);
xor U4208 (N_4208,N_2868,N_149);
nor U4209 (N_4209,N_2969,N_2449);
or U4210 (N_4210,N_829,N_2166);
nor U4211 (N_4211,N_2530,N_1672);
and U4212 (N_4212,N_1390,N_2378);
or U4213 (N_4213,N_1397,N_2683);
xor U4214 (N_4214,N_509,N_1627);
nor U4215 (N_4215,N_678,N_2222);
xnor U4216 (N_4216,N_372,N_1549);
and U4217 (N_4217,N_1028,N_967);
and U4218 (N_4218,N_2250,N_2828);
and U4219 (N_4219,N_1262,N_1805);
nor U4220 (N_4220,N_2862,N_897);
nor U4221 (N_4221,N_1211,N_2898);
and U4222 (N_4222,N_2572,N_602);
or U4223 (N_4223,N_1937,N_2490);
or U4224 (N_4224,N_1159,N_900);
or U4225 (N_4225,N_1167,N_586);
xor U4226 (N_4226,N_2394,N_2556);
nor U4227 (N_4227,N_476,N_2464);
or U4228 (N_4228,N_923,N_2078);
nand U4229 (N_4229,N_1417,N_1776);
and U4230 (N_4230,N_2234,N_1552);
nor U4231 (N_4231,N_30,N_614);
xor U4232 (N_4232,N_13,N_51);
nand U4233 (N_4233,N_729,N_320);
or U4234 (N_4234,N_309,N_1131);
xnor U4235 (N_4235,N_1114,N_2818);
xor U4236 (N_4236,N_140,N_1984);
or U4237 (N_4237,N_2501,N_2363);
and U4238 (N_4238,N_1338,N_1250);
xor U4239 (N_4239,N_625,N_328);
or U4240 (N_4240,N_171,N_1807);
and U4241 (N_4241,N_1379,N_2432);
xor U4242 (N_4242,N_1142,N_902);
or U4243 (N_4243,N_707,N_2989);
or U4244 (N_4244,N_2982,N_2617);
nand U4245 (N_4245,N_2520,N_1757);
and U4246 (N_4246,N_1567,N_1063);
or U4247 (N_4247,N_2175,N_2338);
xnor U4248 (N_4248,N_1164,N_241);
nor U4249 (N_4249,N_819,N_146);
xor U4250 (N_4250,N_1958,N_672);
and U4251 (N_4251,N_1605,N_571);
and U4252 (N_4252,N_2577,N_1717);
nor U4253 (N_4253,N_88,N_1187);
nor U4254 (N_4254,N_1563,N_1526);
and U4255 (N_4255,N_448,N_466);
or U4256 (N_4256,N_2365,N_1766);
and U4257 (N_4257,N_2131,N_1816);
nand U4258 (N_4258,N_2273,N_929);
nor U4259 (N_4259,N_2729,N_198);
nor U4260 (N_4260,N_1497,N_2235);
nor U4261 (N_4261,N_1591,N_1619);
or U4262 (N_4262,N_659,N_1323);
nor U4263 (N_4263,N_232,N_2114);
and U4264 (N_4264,N_1538,N_1738);
nor U4265 (N_4265,N_1221,N_1533);
nand U4266 (N_4266,N_332,N_2033);
or U4267 (N_4267,N_2304,N_2112);
nor U4268 (N_4268,N_1912,N_2006);
or U4269 (N_4269,N_1785,N_1618);
and U4270 (N_4270,N_1674,N_2172);
nor U4271 (N_4271,N_1862,N_2542);
and U4272 (N_4272,N_1474,N_1913);
or U4273 (N_4273,N_524,N_1378);
nor U4274 (N_4274,N_2069,N_2739);
or U4275 (N_4275,N_2479,N_1851);
nand U4276 (N_4276,N_1195,N_431);
nor U4277 (N_4277,N_1047,N_1062);
nand U4278 (N_4278,N_124,N_104);
nand U4279 (N_4279,N_2570,N_644);
nor U4280 (N_4280,N_1575,N_2559);
and U4281 (N_4281,N_1803,N_2908);
and U4282 (N_4282,N_122,N_649);
or U4283 (N_4283,N_1818,N_1197);
xnor U4284 (N_4284,N_1422,N_786);
nor U4285 (N_4285,N_26,N_841);
or U4286 (N_4286,N_2673,N_1055);
or U4287 (N_4287,N_2074,N_2798);
and U4288 (N_4288,N_2463,N_1282);
nor U4289 (N_4289,N_2996,N_721);
xnor U4290 (N_4290,N_1817,N_1995);
xnor U4291 (N_4291,N_2096,N_689);
xor U4292 (N_4292,N_2461,N_794);
xor U4293 (N_4293,N_2902,N_1506);
nor U4294 (N_4294,N_840,N_433);
nor U4295 (N_4295,N_1336,N_1298);
xor U4296 (N_4296,N_2071,N_2065);
xnor U4297 (N_4297,N_1032,N_2502);
nand U4298 (N_4298,N_952,N_1583);
and U4299 (N_4299,N_1955,N_2625);
or U4300 (N_4300,N_766,N_579);
nor U4301 (N_4301,N_2771,N_2762);
and U4302 (N_4302,N_1819,N_857);
nand U4303 (N_4303,N_2417,N_610);
nor U4304 (N_4304,N_1134,N_2592);
nand U4305 (N_4305,N_1284,N_1462);
nand U4306 (N_4306,N_1873,N_1395);
xnor U4307 (N_4307,N_327,N_339);
and U4308 (N_4308,N_1524,N_2425);
or U4309 (N_4309,N_2925,N_2816);
or U4310 (N_4310,N_50,N_821);
nor U4311 (N_4311,N_1713,N_1630);
nand U4312 (N_4312,N_1061,N_2005);
and U4313 (N_4313,N_438,N_1993);
or U4314 (N_4314,N_2848,N_1535);
and U4315 (N_4315,N_2437,N_239);
nor U4316 (N_4316,N_1064,N_1013);
and U4317 (N_4317,N_1731,N_2475);
or U4318 (N_4318,N_1257,N_2419);
xor U4319 (N_4319,N_1919,N_2429);
and U4320 (N_4320,N_2609,N_1543);
and U4321 (N_4321,N_585,N_1400);
nand U4322 (N_4322,N_663,N_1020);
and U4323 (N_4323,N_1521,N_2374);
xnor U4324 (N_4324,N_2620,N_201);
nor U4325 (N_4325,N_613,N_1482);
nor U4326 (N_4326,N_2825,N_940);
and U4327 (N_4327,N_2760,N_2409);
or U4328 (N_4328,N_1297,N_1547);
or U4329 (N_4329,N_186,N_1824);
or U4330 (N_4330,N_2146,N_2043);
nand U4331 (N_4331,N_386,N_1698);
or U4332 (N_4332,N_913,N_1491);
nand U4333 (N_4333,N_1555,N_1865);
nand U4334 (N_4334,N_1705,N_800);
or U4335 (N_4335,N_2393,N_2130);
and U4336 (N_4336,N_2203,N_2684);
or U4337 (N_4337,N_318,N_373);
or U4338 (N_4338,N_1846,N_1822);
xnor U4339 (N_4339,N_2863,N_2826);
nor U4340 (N_4340,N_2121,N_560);
nor U4341 (N_4341,N_120,N_375);
xnor U4342 (N_4342,N_1073,N_906);
xnor U4343 (N_4343,N_2924,N_2951);
or U4344 (N_4344,N_1281,N_1573);
xor U4345 (N_4345,N_2039,N_1741);
and U4346 (N_4346,N_1826,N_2614);
or U4347 (N_4347,N_2708,N_781);
nand U4348 (N_4348,N_1172,N_1364);
and U4349 (N_4349,N_1745,N_2395);
nand U4350 (N_4350,N_1492,N_2535);
nand U4351 (N_4351,N_1193,N_2341);
xnor U4352 (N_4352,N_2986,N_1507);
or U4353 (N_4353,N_2489,N_2238);
and U4354 (N_4354,N_1202,N_1477);
or U4355 (N_4355,N_1366,N_360);
nor U4356 (N_4356,N_132,N_2274);
xnor U4357 (N_4357,N_1054,N_477);
xor U4358 (N_4358,N_862,N_1075);
or U4359 (N_4359,N_685,N_772);
or U4360 (N_4360,N_1529,N_1684);
xnor U4361 (N_4361,N_11,N_2332);
nand U4362 (N_4362,N_2971,N_2379);
or U4363 (N_4363,N_1602,N_1500);
nor U4364 (N_4364,N_1782,N_836);
nor U4365 (N_4365,N_2116,N_1902);
or U4366 (N_4366,N_2589,N_1261);
or U4367 (N_4367,N_954,N_1173);
nand U4368 (N_4368,N_867,N_380);
xnor U4369 (N_4369,N_2634,N_2360);
nand U4370 (N_4370,N_1331,N_1335);
or U4371 (N_4371,N_1240,N_29);
xnor U4372 (N_4372,N_1802,N_851);
or U4373 (N_4373,N_1572,N_160);
nand U4374 (N_4374,N_2687,N_545);
nor U4375 (N_4375,N_2756,N_2688);
xor U4376 (N_4376,N_1380,N_2995);
nor U4377 (N_4377,N_2703,N_632);
nand U4378 (N_4378,N_2500,N_909);
xor U4379 (N_4379,N_1160,N_366);
nand U4380 (N_4380,N_453,N_1051);
or U4381 (N_4381,N_2288,N_207);
nand U4382 (N_4382,N_1411,N_1925);
nor U4383 (N_4383,N_521,N_679);
nor U4384 (N_4384,N_330,N_1350);
or U4385 (N_4385,N_2011,N_133);
nor U4386 (N_4386,N_741,N_2674);
nand U4387 (N_4387,N_604,N_970);
xor U4388 (N_4388,N_2881,N_720);
and U4389 (N_4389,N_1690,N_1829);
nor U4390 (N_4390,N_1606,N_1594);
nor U4391 (N_4391,N_817,N_557);
nand U4392 (N_4392,N_1342,N_833);
nor U4393 (N_4393,N_1102,N_2336);
nor U4394 (N_4394,N_1751,N_1596);
nor U4395 (N_4395,N_818,N_1419);
nor U4396 (N_4396,N_2607,N_1729);
xnor U4397 (N_4397,N_1076,N_2910);
xor U4398 (N_4398,N_94,N_1360);
nor U4399 (N_4399,N_1396,N_1680);
nand U4400 (N_4400,N_129,N_2470);
nor U4401 (N_4401,N_2022,N_203);
xor U4402 (N_4402,N_2730,N_528);
and U4403 (N_4403,N_2966,N_2319);
nor U4404 (N_4404,N_1483,N_2236);
and U4405 (N_4405,N_754,N_1330);
or U4406 (N_4406,N_2538,N_185);
nand U4407 (N_4407,N_119,N_2998);
or U4408 (N_4408,N_2484,N_1676);
and U4409 (N_4409,N_1292,N_2164);
nor U4410 (N_4410,N_2550,N_2144);
nand U4411 (N_4411,N_2302,N_1339);
and U4412 (N_4412,N_642,N_762);
or U4413 (N_4413,N_256,N_944);
or U4414 (N_4414,N_461,N_1637);
nand U4415 (N_4415,N_2877,N_1399);
nor U4416 (N_4416,N_905,N_1584);
and U4417 (N_4417,N_1685,N_635);
xor U4418 (N_4418,N_399,N_853);
nor U4419 (N_4419,N_1603,N_536);
and U4420 (N_4420,N_1767,N_1138);
nor U4421 (N_4421,N_1456,N_1357);
nand U4422 (N_4422,N_705,N_963);
xnor U4423 (N_4423,N_1595,N_2723);
or U4424 (N_4424,N_2641,N_292);
or U4425 (N_4425,N_716,N_1291);
and U4426 (N_4426,N_2615,N_516);
or U4427 (N_4427,N_1254,N_2866);
and U4428 (N_4428,N_2606,N_2444);
or U4429 (N_4429,N_152,N_2584);
nor U4430 (N_4430,N_1498,N_1614);
nor U4431 (N_4431,N_2642,N_722);
or U4432 (N_4432,N_2679,N_2582);
nand U4433 (N_4433,N_1910,N_2740);
nand U4434 (N_4434,N_1421,N_2016);
or U4435 (N_4435,N_1847,N_1796);
nand U4436 (N_4436,N_811,N_2231);
or U4437 (N_4437,N_2237,N_1216);
nand U4438 (N_4438,N_769,N_2279);
nor U4439 (N_4439,N_1322,N_1300);
or U4440 (N_4440,N_1773,N_837);
and U4441 (N_4441,N_948,N_1209);
nor U4442 (N_4442,N_550,N_2623);
xnor U4443 (N_4443,N_1855,N_2717);
and U4444 (N_4444,N_595,N_866);
xor U4445 (N_4445,N_2901,N_2020);
and U4446 (N_4446,N_429,N_2162);
or U4447 (N_4447,N_76,N_1636);
and U4448 (N_4448,N_1045,N_1451);
and U4449 (N_4449,N_193,N_34);
nand U4450 (N_4450,N_1235,N_1510);
or U4451 (N_4451,N_562,N_236);
or U4452 (N_4452,N_1954,N_1598);
or U4453 (N_4453,N_1580,N_2906);
and U4454 (N_4454,N_1649,N_2330);
and U4455 (N_4455,N_2149,N_2873);
and U4456 (N_4456,N_1620,N_2296);
xnor U4457 (N_4457,N_1238,N_2293);
nor U4458 (N_4458,N_1161,N_1374);
xnor U4459 (N_4459,N_1914,N_820);
xor U4460 (N_4460,N_2454,N_1688);
xnor U4461 (N_4461,N_1,N_1208);
nor U4462 (N_4462,N_734,N_2431);
and U4463 (N_4463,N_2840,N_2650);
and U4464 (N_4464,N_1077,N_2191);
nor U4465 (N_4465,N_1310,N_695);
and U4466 (N_4466,N_2295,N_2037);
and U4467 (N_4467,N_2603,N_1991);
xor U4468 (N_4468,N_187,N_573);
or U4469 (N_4469,N_2921,N_686);
nand U4470 (N_4470,N_588,N_1774);
nand U4471 (N_4471,N_2090,N_40);
or U4472 (N_4472,N_483,N_1827);
or U4473 (N_4473,N_1863,N_2270);
nor U4474 (N_4474,N_408,N_730);
and U4475 (N_4475,N_376,N_1660);
and U4476 (N_4476,N_886,N_2211);
nand U4477 (N_4477,N_1192,N_2173);
nor U4478 (N_4478,N_1425,N_984);
nor U4479 (N_4479,N_2566,N_1748);
nand U4480 (N_4480,N_2091,N_2672);
nand U4481 (N_4481,N_1640,N_2359);
and U4482 (N_4482,N_1067,N_1305);
nor U4483 (N_4483,N_849,N_224);
nor U4484 (N_4484,N_2909,N_1590);
and U4485 (N_4485,N_2407,N_1085);
nor U4486 (N_4486,N_1599,N_2414);
xor U4487 (N_4487,N_1022,N_1976);
or U4488 (N_4488,N_2132,N_2053);
xnor U4489 (N_4489,N_369,N_643);
and U4490 (N_4490,N_2543,N_988);
xor U4491 (N_4491,N_1367,N_2972);
or U4492 (N_4492,N_2573,N_1103);
nand U4493 (N_4493,N_163,N_1612);
xnor U4494 (N_4494,N_440,N_2216);
or U4495 (N_4495,N_1145,N_2491);
xnor U4496 (N_4496,N_202,N_568);
nor U4497 (N_4497,N_709,N_1588);
nor U4498 (N_4498,N_2318,N_1869);
and U4499 (N_4499,N_2574,N_2354);
nand U4500 (N_4500,N_2121,N_2592);
nor U4501 (N_4501,N_2655,N_1597);
nor U4502 (N_4502,N_1317,N_1883);
or U4503 (N_4503,N_2372,N_1027);
and U4504 (N_4504,N_2222,N_2694);
xor U4505 (N_4505,N_647,N_2253);
or U4506 (N_4506,N_2433,N_1562);
nor U4507 (N_4507,N_2756,N_1223);
xnor U4508 (N_4508,N_1995,N_2964);
xor U4509 (N_4509,N_1833,N_1202);
nor U4510 (N_4510,N_2776,N_1106);
nor U4511 (N_4511,N_256,N_2886);
xnor U4512 (N_4512,N_1815,N_2439);
nor U4513 (N_4513,N_1992,N_1833);
and U4514 (N_4514,N_2002,N_2612);
nor U4515 (N_4515,N_1098,N_762);
xnor U4516 (N_4516,N_305,N_1403);
and U4517 (N_4517,N_410,N_2069);
xnor U4518 (N_4518,N_168,N_1574);
or U4519 (N_4519,N_533,N_1169);
nor U4520 (N_4520,N_822,N_1565);
xnor U4521 (N_4521,N_1609,N_494);
or U4522 (N_4522,N_216,N_2142);
and U4523 (N_4523,N_2591,N_874);
and U4524 (N_4524,N_2092,N_1408);
xnor U4525 (N_4525,N_82,N_2774);
nor U4526 (N_4526,N_2139,N_1803);
nor U4527 (N_4527,N_1694,N_2799);
and U4528 (N_4528,N_558,N_2543);
nand U4529 (N_4529,N_1271,N_2842);
nor U4530 (N_4530,N_509,N_1702);
nor U4531 (N_4531,N_163,N_2366);
and U4532 (N_4532,N_2169,N_878);
or U4533 (N_4533,N_2002,N_2986);
and U4534 (N_4534,N_2524,N_1816);
and U4535 (N_4535,N_2080,N_1567);
xor U4536 (N_4536,N_647,N_2052);
or U4537 (N_4537,N_690,N_2304);
and U4538 (N_4538,N_1529,N_1464);
xor U4539 (N_4539,N_2018,N_440);
and U4540 (N_4540,N_340,N_2297);
nor U4541 (N_4541,N_502,N_0);
and U4542 (N_4542,N_2867,N_638);
nand U4543 (N_4543,N_853,N_1168);
or U4544 (N_4544,N_892,N_2197);
nor U4545 (N_4545,N_13,N_2077);
or U4546 (N_4546,N_2705,N_714);
and U4547 (N_4547,N_2758,N_2656);
nor U4548 (N_4548,N_1547,N_396);
and U4549 (N_4549,N_2238,N_1376);
and U4550 (N_4550,N_779,N_2499);
nand U4551 (N_4551,N_2204,N_593);
nand U4552 (N_4552,N_109,N_1689);
or U4553 (N_4553,N_1738,N_1427);
nor U4554 (N_4554,N_1626,N_1546);
xnor U4555 (N_4555,N_305,N_552);
xor U4556 (N_4556,N_730,N_1472);
nor U4557 (N_4557,N_909,N_677);
xnor U4558 (N_4558,N_1419,N_2690);
or U4559 (N_4559,N_1392,N_2921);
or U4560 (N_4560,N_2285,N_2500);
and U4561 (N_4561,N_1764,N_1004);
xor U4562 (N_4562,N_236,N_2927);
nand U4563 (N_4563,N_1530,N_2624);
nor U4564 (N_4564,N_1377,N_2527);
nor U4565 (N_4565,N_299,N_1815);
nand U4566 (N_4566,N_2850,N_1532);
and U4567 (N_4567,N_619,N_1853);
nand U4568 (N_4568,N_2472,N_1374);
xor U4569 (N_4569,N_1108,N_1465);
nor U4570 (N_4570,N_1073,N_631);
and U4571 (N_4571,N_2680,N_2608);
nor U4572 (N_4572,N_2911,N_2883);
or U4573 (N_4573,N_1264,N_629);
nand U4574 (N_4574,N_1170,N_187);
and U4575 (N_4575,N_1683,N_871);
xnor U4576 (N_4576,N_1908,N_2766);
nand U4577 (N_4577,N_1628,N_2976);
nand U4578 (N_4578,N_2724,N_2737);
nand U4579 (N_4579,N_2780,N_1734);
or U4580 (N_4580,N_1141,N_2795);
xnor U4581 (N_4581,N_1118,N_1419);
nor U4582 (N_4582,N_834,N_2812);
and U4583 (N_4583,N_748,N_1746);
xor U4584 (N_4584,N_1273,N_2248);
nor U4585 (N_4585,N_895,N_2724);
xnor U4586 (N_4586,N_2668,N_830);
nand U4587 (N_4587,N_567,N_1019);
xor U4588 (N_4588,N_2305,N_1662);
nor U4589 (N_4589,N_1485,N_519);
and U4590 (N_4590,N_2531,N_2612);
xor U4591 (N_4591,N_1466,N_1686);
nor U4592 (N_4592,N_1882,N_815);
nand U4593 (N_4593,N_2972,N_2520);
or U4594 (N_4594,N_897,N_2024);
and U4595 (N_4595,N_2739,N_500);
nor U4596 (N_4596,N_1649,N_2918);
xor U4597 (N_4597,N_2212,N_2260);
or U4598 (N_4598,N_1671,N_1090);
nand U4599 (N_4599,N_2189,N_1671);
nand U4600 (N_4600,N_1353,N_1357);
or U4601 (N_4601,N_598,N_737);
or U4602 (N_4602,N_2606,N_1595);
nor U4603 (N_4603,N_1456,N_1441);
nor U4604 (N_4604,N_1062,N_2988);
or U4605 (N_4605,N_1303,N_2220);
nand U4606 (N_4606,N_2598,N_1216);
xnor U4607 (N_4607,N_1316,N_1902);
or U4608 (N_4608,N_2568,N_219);
and U4609 (N_4609,N_2166,N_752);
and U4610 (N_4610,N_1849,N_1461);
or U4611 (N_4611,N_1647,N_1269);
nor U4612 (N_4612,N_2143,N_1761);
or U4613 (N_4613,N_275,N_2658);
or U4614 (N_4614,N_186,N_782);
and U4615 (N_4615,N_2881,N_2339);
nand U4616 (N_4616,N_347,N_2267);
nor U4617 (N_4617,N_933,N_965);
xor U4618 (N_4618,N_2041,N_677);
and U4619 (N_4619,N_299,N_579);
or U4620 (N_4620,N_994,N_1589);
or U4621 (N_4621,N_1698,N_427);
nand U4622 (N_4622,N_1678,N_1475);
xnor U4623 (N_4623,N_699,N_947);
nand U4624 (N_4624,N_2325,N_32);
or U4625 (N_4625,N_1804,N_1108);
xnor U4626 (N_4626,N_1051,N_2772);
and U4627 (N_4627,N_1357,N_2627);
nand U4628 (N_4628,N_1919,N_27);
and U4629 (N_4629,N_1871,N_1578);
xor U4630 (N_4630,N_1473,N_1592);
nand U4631 (N_4631,N_1211,N_156);
nor U4632 (N_4632,N_183,N_2896);
nand U4633 (N_4633,N_90,N_923);
or U4634 (N_4634,N_254,N_931);
nand U4635 (N_4635,N_2754,N_2492);
nor U4636 (N_4636,N_59,N_237);
xor U4637 (N_4637,N_2286,N_2360);
and U4638 (N_4638,N_1967,N_1430);
xnor U4639 (N_4639,N_1217,N_970);
nor U4640 (N_4640,N_511,N_351);
and U4641 (N_4641,N_1940,N_752);
nor U4642 (N_4642,N_1951,N_2844);
xnor U4643 (N_4643,N_513,N_2977);
and U4644 (N_4644,N_1356,N_1280);
xnor U4645 (N_4645,N_2603,N_699);
nor U4646 (N_4646,N_880,N_1099);
or U4647 (N_4647,N_2409,N_567);
and U4648 (N_4648,N_442,N_2175);
and U4649 (N_4649,N_1674,N_1805);
or U4650 (N_4650,N_1255,N_2726);
or U4651 (N_4651,N_2955,N_343);
xor U4652 (N_4652,N_218,N_316);
xor U4653 (N_4653,N_607,N_888);
nor U4654 (N_4654,N_1887,N_1488);
xnor U4655 (N_4655,N_2069,N_1868);
nand U4656 (N_4656,N_254,N_1899);
nor U4657 (N_4657,N_2820,N_848);
nand U4658 (N_4658,N_2408,N_976);
or U4659 (N_4659,N_1574,N_708);
and U4660 (N_4660,N_1396,N_2072);
xnor U4661 (N_4661,N_593,N_2542);
or U4662 (N_4662,N_1004,N_2185);
xor U4663 (N_4663,N_1704,N_1606);
nor U4664 (N_4664,N_2117,N_272);
xor U4665 (N_4665,N_1221,N_2472);
or U4666 (N_4666,N_2765,N_2079);
nand U4667 (N_4667,N_546,N_148);
nor U4668 (N_4668,N_1694,N_2548);
and U4669 (N_4669,N_2582,N_85);
or U4670 (N_4670,N_2336,N_2440);
xnor U4671 (N_4671,N_2276,N_2940);
xnor U4672 (N_4672,N_1912,N_1380);
nand U4673 (N_4673,N_498,N_849);
xnor U4674 (N_4674,N_2814,N_2014);
nand U4675 (N_4675,N_979,N_1701);
nor U4676 (N_4676,N_2403,N_2026);
nor U4677 (N_4677,N_1391,N_408);
xnor U4678 (N_4678,N_2289,N_974);
nand U4679 (N_4679,N_1192,N_1914);
nand U4680 (N_4680,N_1642,N_2192);
or U4681 (N_4681,N_2499,N_1332);
xor U4682 (N_4682,N_2402,N_1013);
or U4683 (N_4683,N_1898,N_832);
or U4684 (N_4684,N_1902,N_1253);
xnor U4685 (N_4685,N_2898,N_2416);
nand U4686 (N_4686,N_1225,N_2688);
nor U4687 (N_4687,N_2197,N_575);
or U4688 (N_4688,N_892,N_2897);
and U4689 (N_4689,N_359,N_2410);
and U4690 (N_4690,N_2207,N_2);
nand U4691 (N_4691,N_2322,N_2890);
nand U4692 (N_4692,N_1406,N_2828);
and U4693 (N_4693,N_2512,N_2429);
nor U4694 (N_4694,N_575,N_2632);
xor U4695 (N_4695,N_1780,N_187);
nand U4696 (N_4696,N_1364,N_1137);
or U4697 (N_4697,N_619,N_2396);
nand U4698 (N_4698,N_2129,N_2733);
nand U4699 (N_4699,N_2954,N_2829);
xor U4700 (N_4700,N_883,N_1062);
and U4701 (N_4701,N_1137,N_1636);
nor U4702 (N_4702,N_2779,N_2471);
nand U4703 (N_4703,N_606,N_2976);
and U4704 (N_4704,N_389,N_842);
nor U4705 (N_4705,N_2971,N_1091);
or U4706 (N_4706,N_2051,N_1770);
or U4707 (N_4707,N_1732,N_2343);
xnor U4708 (N_4708,N_825,N_365);
and U4709 (N_4709,N_325,N_2836);
or U4710 (N_4710,N_2886,N_1413);
or U4711 (N_4711,N_870,N_972);
nand U4712 (N_4712,N_1559,N_2654);
and U4713 (N_4713,N_1243,N_729);
or U4714 (N_4714,N_2329,N_2134);
and U4715 (N_4715,N_875,N_862);
nor U4716 (N_4716,N_333,N_1605);
nor U4717 (N_4717,N_2844,N_171);
nand U4718 (N_4718,N_506,N_2979);
or U4719 (N_4719,N_2107,N_178);
nand U4720 (N_4720,N_2334,N_1668);
nor U4721 (N_4721,N_9,N_1834);
xnor U4722 (N_4722,N_2039,N_2753);
xor U4723 (N_4723,N_2640,N_2213);
nor U4724 (N_4724,N_79,N_443);
nand U4725 (N_4725,N_1519,N_2485);
xnor U4726 (N_4726,N_1828,N_1887);
xor U4727 (N_4727,N_1747,N_823);
nand U4728 (N_4728,N_1490,N_2744);
nor U4729 (N_4729,N_1156,N_2765);
nand U4730 (N_4730,N_948,N_2036);
xor U4731 (N_4731,N_2854,N_1437);
and U4732 (N_4732,N_1391,N_466);
xnor U4733 (N_4733,N_893,N_641);
nand U4734 (N_4734,N_223,N_2648);
xnor U4735 (N_4735,N_2618,N_2593);
or U4736 (N_4736,N_2651,N_336);
nor U4737 (N_4737,N_941,N_1723);
nor U4738 (N_4738,N_2413,N_1329);
xnor U4739 (N_4739,N_308,N_637);
and U4740 (N_4740,N_1298,N_1717);
nand U4741 (N_4741,N_2534,N_2420);
nand U4742 (N_4742,N_411,N_2155);
xnor U4743 (N_4743,N_681,N_753);
and U4744 (N_4744,N_1076,N_835);
nand U4745 (N_4745,N_1732,N_2416);
nor U4746 (N_4746,N_374,N_808);
nor U4747 (N_4747,N_479,N_2569);
and U4748 (N_4748,N_530,N_2409);
xnor U4749 (N_4749,N_1039,N_1984);
nand U4750 (N_4750,N_1792,N_1411);
nor U4751 (N_4751,N_2611,N_1847);
nand U4752 (N_4752,N_1335,N_2642);
nand U4753 (N_4753,N_102,N_1004);
xor U4754 (N_4754,N_413,N_148);
or U4755 (N_4755,N_2258,N_1359);
nor U4756 (N_4756,N_2527,N_2340);
xnor U4757 (N_4757,N_1271,N_2720);
nor U4758 (N_4758,N_2436,N_1561);
nor U4759 (N_4759,N_1942,N_2139);
and U4760 (N_4760,N_658,N_34);
nand U4761 (N_4761,N_2701,N_2396);
or U4762 (N_4762,N_2036,N_2129);
nor U4763 (N_4763,N_957,N_286);
nand U4764 (N_4764,N_1754,N_1020);
and U4765 (N_4765,N_2275,N_632);
nor U4766 (N_4766,N_330,N_1380);
xor U4767 (N_4767,N_1813,N_1492);
xnor U4768 (N_4768,N_2862,N_479);
nand U4769 (N_4769,N_2876,N_2068);
nor U4770 (N_4770,N_1654,N_371);
or U4771 (N_4771,N_2258,N_605);
and U4772 (N_4772,N_2493,N_957);
and U4773 (N_4773,N_1092,N_2114);
and U4774 (N_4774,N_146,N_2873);
or U4775 (N_4775,N_56,N_1720);
nor U4776 (N_4776,N_2438,N_2857);
and U4777 (N_4777,N_930,N_1053);
nand U4778 (N_4778,N_2091,N_603);
or U4779 (N_4779,N_193,N_426);
or U4780 (N_4780,N_802,N_140);
and U4781 (N_4781,N_1495,N_1662);
and U4782 (N_4782,N_1074,N_733);
nand U4783 (N_4783,N_2224,N_1122);
nand U4784 (N_4784,N_2191,N_1927);
nor U4785 (N_4785,N_2444,N_450);
or U4786 (N_4786,N_145,N_1912);
nand U4787 (N_4787,N_191,N_1454);
and U4788 (N_4788,N_1961,N_107);
and U4789 (N_4789,N_342,N_439);
xor U4790 (N_4790,N_640,N_839);
xnor U4791 (N_4791,N_1299,N_2214);
nor U4792 (N_4792,N_905,N_1414);
and U4793 (N_4793,N_2798,N_899);
xor U4794 (N_4794,N_379,N_2342);
and U4795 (N_4795,N_2618,N_2241);
nand U4796 (N_4796,N_22,N_19);
and U4797 (N_4797,N_267,N_958);
or U4798 (N_4798,N_1586,N_1312);
or U4799 (N_4799,N_1981,N_907);
and U4800 (N_4800,N_1139,N_644);
nor U4801 (N_4801,N_468,N_2612);
and U4802 (N_4802,N_737,N_1567);
or U4803 (N_4803,N_340,N_2558);
nor U4804 (N_4804,N_630,N_961);
or U4805 (N_4805,N_2500,N_514);
and U4806 (N_4806,N_2435,N_494);
nor U4807 (N_4807,N_2469,N_325);
xnor U4808 (N_4808,N_1975,N_2812);
or U4809 (N_4809,N_2891,N_2233);
xnor U4810 (N_4810,N_2741,N_2712);
nor U4811 (N_4811,N_2411,N_1514);
or U4812 (N_4812,N_1320,N_1918);
xor U4813 (N_4813,N_1822,N_2044);
xor U4814 (N_4814,N_971,N_1839);
xor U4815 (N_4815,N_2796,N_529);
and U4816 (N_4816,N_1604,N_528);
or U4817 (N_4817,N_219,N_204);
nand U4818 (N_4818,N_1738,N_1785);
nand U4819 (N_4819,N_1086,N_2057);
nor U4820 (N_4820,N_1162,N_2572);
nand U4821 (N_4821,N_2316,N_1927);
xor U4822 (N_4822,N_1036,N_2059);
and U4823 (N_4823,N_2867,N_2754);
nand U4824 (N_4824,N_2450,N_2096);
nor U4825 (N_4825,N_750,N_1568);
xor U4826 (N_4826,N_2363,N_2528);
and U4827 (N_4827,N_2743,N_2237);
xor U4828 (N_4828,N_2905,N_1962);
or U4829 (N_4829,N_476,N_34);
or U4830 (N_4830,N_2447,N_650);
and U4831 (N_4831,N_2156,N_1756);
or U4832 (N_4832,N_395,N_762);
nand U4833 (N_4833,N_196,N_476);
xnor U4834 (N_4834,N_1604,N_584);
nand U4835 (N_4835,N_2385,N_1939);
or U4836 (N_4836,N_2456,N_2172);
nor U4837 (N_4837,N_7,N_1012);
xnor U4838 (N_4838,N_2684,N_2380);
nor U4839 (N_4839,N_1719,N_974);
nand U4840 (N_4840,N_1796,N_2001);
and U4841 (N_4841,N_344,N_2884);
nand U4842 (N_4842,N_284,N_2005);
and U4843 (N_4843,N_2386,N_1919);
or U4844 (N_4844,N_1847,N_2671);
or U4845 (N_4845,N_221,N_2767);
and U4846 (N_4846,N_33,N_1811);
nand U4847 (N_4847,N_2039,N_2451);
and U4848 (N_4848,N_867,N_1767);
and U4849 (N_4849,N_544,N_279);
nor U4850 (N_4850,N_1872,N_644);
and U4851 (N_4851,N_1108,N_553);
or U4852 (N_4852,N_871,N_2024);
nor U4853 (N_4853,N_2827,N_440);
xnor U4854 (N_4854,N_344,N_2603);
or U4855 (N_4855,N_105,N_167);
xnor U4856 (N_4856,N_447,N_1055);
or U4857 (N_4857,N_1202,N_2113);
or U4858 (N_4858,N_1583,N_2775);
nor U4859 (N_4859,N_192,N_2921);
and U4860 (N_4860,N_1568,N_2199);
and U4861 (N_4861,N_42,N_800);
xnor U4862 (N_4862,N_116,N_1568);
xor U4863 (N_4863,N_854,N_466);
or U4864 (N_4864,N_1875,N_4);
nor U4865 (N_4865,N_1078,N_190);
or U4866 (N_4866,N_2518,N_1410);
or U4867 (N_4867,N_2180,N_19);
and U4868 (N_4868,N_2602,N_991);
nand U4869 (N_4869,N_566,N_630);
nor U4870 (N_4870,N_300,N_1353);
xnor U4871 (N_4871,N_2464,N_2428);
xnor U4872 (N_4872,N_836,N_931);
nor U4873 (N_4873,N_2300,N_2251);
nand U4874 (N_4874,N_1605,N_173);
or U4875 (N_4875,N_2857,N_1729);
xnor U4876 (N_4876,N_1942,N_988);
nand U4877 (N_4877,N_2443,N_267);
and U4878 (N_4878,N_2095,N_1545);
nand U4879 (N_4879,N_2638,N_1743);
or U4880 (N_4880,N_2066,N_1850);
xor U4881 (N_4881,N_2645,N_1937);
and U4882 (N_4882,N_539,N_149);
and U4883 (N_4883,N_893,N_698);
or U4884 (N_4884,N_158,N_2231);
xor U4885 (N_4885,N_815,N_245);
xnor U4886 (N_4886,N_680,N_2323);
or U4887 (N_4887,N_1074,N_2886);
xor U4888 (N_4888,N_318,N_37);
nor U4889 (N_4889,N_2080,N_2974);
nand U4890 (N_4890,N_1862,N_512);
nor U4891 (N_4891,N_19,N_1923);
nor U4892 (N_4892,N_1384,N_1845);
xnor U4893 (N_4893,N_2112,N_2309);
or U4894 (N_4894,N_2850,N_2361);
and U4895 (N_4895,N_2468,N_216);
nor U4896 (N_4896,N_98,N_2074);
or U4897 (N_4897,N_969,N_2873);
nand U4898 (N_4898,N_1589,N_2709);
and U4899 (N_4899,N_600,N_1007);
nand U4900 (N_4900,N_1360,N_2598);
or U4901 (N_4901,N_1545,N_1515);
and U4902 (N_4902,N_711,N_2059);
or U4903 (N_4903,N_1514,N_2611);
nor U4904 (N_4904,N_1445,N_1501);
and U4905 (N_4905,N_2045,N_668);
nand U4906 (N_4906,N_1926,N_2653);
or U4907 (N_4907,N_715,N_1921);
xor U4908 (N_4908,N_98,N_20);
nand U4909 (N_4909,N_1482,N_2401);
and U4910 (N_4910,N_1929,N_2279);
xor U4911 (N_4911,N_113,N_104);
xnor U4912 (N_4912,N_252,N_1633);
nand U4913 (N_4913,N_8,N_1998);
and U4914 (N_4914,N_2576,N_1543);
and U4915 (N_4915,N_2999,N_437);
xor U4916 (N_4916,N_1539,N_967);
or U4917 (N_4917,N_41,N_1412);
nand U4918 (N_4918,N_721,N_1393);
or U4919 (N_4919,N_1481,N_273);
nor U4920 (N_4920,N_711,N_1950);
and U4921 (N_4921,N_702,N_1378);
nand U4922 (N_4922,N_2374,N_807);
nor U4923 (N_4923,N_753,N_2014);
or U4924 (N_4924,N_2481,N_1005);
or U4925 (N_4925,N_946,N_1470);
nor U4926 (N_4926,N_970,N_2758);
xnor U4927 (N_4927,N_1569,N_27);
and U4928 (N_4928,N_745,N_544);
nor U4929 (N_4929,N_1873,N_1643);
or U4930 (N_4930,N_1350,N_657);
nand U4931 (N_4931,N_1890,N_1341);
and U4932 (N_4932,N_2162,N_1910);
nand U4933 (N_4933,N_614,N_2865);
xor U4934 (N_4934,N_2278,N_41);
or U4935 (N_4935,N_2595,N_2238);
or U4936 (N_4936,N_2126,N_706);
xor U4937 (N_4937,N_1648,N_2973);
or U4938 (N_4938,N_767,N_2206);
xnor U4939 (N_4939,N_1643,N_1942);
nor U4940 (N_4940,N_2971,N_2304);
or U4941 (N_4941,N_2193,N_485);
xor U4942 (N_4942,N_2814,N_1954);
or U4943 (N_4943,N_2588,N_2845);
and U4944 (N_4944,N_89,N_1031);
nand U4945 (N_4945,N_2142,N_1297);
xor U4946 (N_4946,N_1,N_644);
nor U4947 (N_4947,N_2990,N_619);
or U4948 (N_4948,N_2324,N_1590);
nor U4949 (N_4949,N_2265,N_301);
and U4950 (N_4950,N_2040,N_1237);
nand U4951 (N_4951,N_876,N_1148);
nand U4952 (N_4952,N_2382,N_687);
and U4953 (N_4953,N_1892,N_775);
nand U4954 (N_4954,N_1048,N_2754);
or U4955 (N_4955,N_1330,N_14);
nand U4956 (N_4956,N_912,N_2365);
nand U4957 (N_4957,N_2322,N_1143);
and U4958 (N_4958,N_1493,N_2741);
nand U4959 (N_4959,N_1956,N_2793);
nor U4960 (N_4960,N_1952,N_1604);
or U4961 (N_4961,N_1060,N_2100);
xnor U4962 (N_4962,N_798,N_1473);
or U4963 (N_4963,N_260,N_2550);
nand U4964 (N_4964,N_1531,N_484);
nand U4965 (N_4965,N_2034,N_2792);
nor U4966 (N_4966,N_2103,N_1279);
nand U4967 (N_4967,N_169,N_1474);
nand U4968 (N_4968,N_2916,N_1087);
or U4969 (N_4969,N_1454,N_1990);
or U4970 (N_4970,N_1344,N_2368);
or U4971 (N_4971,N_2288,N_2819);
xnor U4972 (N_4972,N_190,N_2925);
and U4973 (N_4973,N_2098,N_825);
and U4974 (N_4974,N_1412,N_2853);
nor U4975 (N_4975,N_572,N_2379);
or U4976 (N_4976,N_1796,N_2665);
xor U4977 (N_4977,N_1514,N_2768);
or U4978 (N_4978,N_129,N_2342);
or U4979 (N_4979,N_531,N_1574);
nor U4980 (N_4980,N_1487,N_1532);
nor U4981 (N_4981,N_1162,N_690);
or U4982 (N_4982,N_2404,N_1628);
and U4983 (N_4983,N_93,N_2877);
nand U4984 (N_4984,N_259,N_2561);
or U4985 (N_4985,N_646,N_1492);
and U4986 (N_4986,N_1412,N_2340);
and U4987 (N_4987,N_802,N_590);
xnor U4988 (N_4988,N_2710,N_209);
xor U4989 (N_4989,N_2426,N_830);
or U4990 (N_4990,N_2393,N_1781);
nand U4991 (N_4991,N_1786,N_1493);
nor U4992 (N_4992,N_2505,N_272);
nand U4993 (N_4993,N_887,N_2771);
and U4994 (N_4994,N_2386,N_2172);
nand U4995 (N_4995,N_2046,N_960);
and U4996 (N_4996,N_969,N_1328);
or U4997 (N_4997,N_230,N_1085);
nand U4998 (N_4998,N_2052,N_1651);
nand U4999 (N_4999,N_1523,N_130);
nand U5000 (N_5000,N_2324,N_2217);
nor U5001 (N_5001,N_2138,N_1306);
xor U5002 (N_5002,N_436,N_934);
nor U5003 (N_5003,N_358,N_768);
nand U5004 (N_5004,N_558,N_1222);
and U5005 (N_5005,N_836,N_2955);
nor U5006 (N_5006,N_107,N_2791);
xnor U5007 (N_5007,N_1992,N_1446);
xor U5008 (N_5008,N_2471,N_486);
or U5009 (N_5009,N_752,N_2493);
and U5010 (N_5010,N_951,N_971);
nand U5011 (N_5011,N_296,N_2822);
or U5012 (N_5012,N_1020,N_2999);
and U5013 (N_5013,N_2325,N_1090);
nand U5014 (N_5014,N_1551,N_2937);
or U5015 (N_5015,N_744,N_192);
and U5016 (N_5016,N_101,N_1865);
and U5017 (N_5017,N_1386,N_1034);
nand U5018 (N_5018,N_26,N_631);
xor U5019 (N_5019,N_1386,N_1128);
or U5020 (N_5020,N_2752,N_335);
nand U5021 (N_5021,N_1591,N_2130);
and U5022 (N_5022,N_1433,N_1193);
nor U5023 (N_5023,N_603,N_2061);
or U5024 (N_5024,N_239,N_1811);
nor U5025 (N_5025,N_2886,N_1271);
nor U5026 (N_5026,N_61,N_2682);
nand U5027 (N_5027,N_2534,N_359);
or U5028 (N_5028,N_2016,N_2083);
nor U5029 (N_5029,N_821,N_2051);
and U5030 (N_5030,N_430,N_1027);
nor U5031 (N_5031,N_845,N_2372);
or U5032 (N_5032,N_1252,N_1770);
nor U5033 (N_5033,N_2762,N_1841);
nor U5034 (N_5034,N_266,N_495);
xor U5035 (N_5035,N_964,N_2204);
or U5036 (N_5036,N_1472,N_2109);
or U5037 (N_5037,N_1494,N_1819);
nand U5038 (N_5038,N_2339,N_91);
nand U5039 (N_5039,N_890,N_1951);
nand U5040 (N_5040,N_2313,N_869);
xor U5041 (N_5041,N_1890,N_354);
xnor U5042 (N_5042,N_1786,N_878);
and U5043 (N_5043,N_836,N_2591);
and U5044 (N_5044,N_595,N_1635);
xnor U5045 (N_5045,N_2300,N_695);
xnor U5046 (N_5046,N_748,N_971);
xnor U5047 (N_5047,N_1984,N_1094);
nand U5048 (N_5048,N_622,N_2063);
or U5049 (N_5049,N_1721,N_2610);
xor U5050 (N_5050,N_2740,N_494);
or U5051 (N_5051,N_1844,N_667);
and U5052 (N_5052,N_1491,N_2117);
nand U5053 (N_5053,N_160,N_1833);
xnor U5054 (N_5054,N_2214,N_2878);
or U5055 (N_5055,N_2229,N_2939);
nor U5056 (N_5056,N_2932,N_205);
or U5057 (N_5057,N_598,N_2338);
and U5058 (N_5058,N_1347,N_2516);
xor U5059 (N_5059,N_1000,N_890);
and U5060 (N_5060,N_1611,N_32);
nor U5061 (N_5061,N_430,N_2604);
xor U5062 (N_5062,N_1356,N_2082);
nor U5063 (N_5063,N_1562,N_2645);
or U5064 (N_5064,N_2719,N_2974);
or U5065 (N_5065,N_1082,N_1568);
nor U5066 (N_5066,N_781,N_2766);
or U5067 (N_5067,N_2600,N_95);
or U5068 (N_5068,N_1246,N_1937);
and U5069 (N_5069,N_610,N_2723);
or U5070 (N_5070,N_1557,N_800);
nand U5071 (N_5071,N_2607,N_2996);
nor U5072 (N_5072,N_2592,N_1042);
nor U5073 (N_5073,N_2334,N_810);
nand U5074 (N_5074,N_2145,N_314);
or U5075 (N_5075,N_1027,N_996);
nor U5076 (N_5076,N_1735,N_2463);
nor U5077 (N_5077,N_19,N_1154);
nor U5078 (N_5078,N_1492,N_2332);
nand U5079 (N_5079,N_2508,N_2315);
and U5080 (N_5080,N_1762,N_1247);
or U5081 (N_5081,N_153,N_2923);
nand U5082 (N_5082,N_2869,N_1469);
and U5083 (N_5083,N_1150,N_1180);
nor U5084 (N_5084,N_1149,N_1442);
nand U5085 (N_5085,N_605,N_2771);
xnor U5086 (N_5086,N_897,N_2359);
xnor U5087 (N_5087,N_798,N_2383);
or U5088 (N_5088,N_926,N_678);
xnor U5089 (N_5089,N_1102,N_2452);
xor U5090 (N_5090,N_297,N_1374);
and U5091 (N_5091,N_2116,N_158);
and U5092 (N_5092,N_1711,N_2733);
nand U5093 (N_5093,N_1297,N_764);
or U5094 (N_5094,N_132,N_1875);
xnor U5095 (N_5095,N_314,N_1007);
or U5096 (N_5096,N_1428,N_584);
or U5097 (N_5097,N_560,N_2549);
or U5098 (N_5098,N_1090,N_2177);
nor U5099 (N_5099,N_459,N_1818);
nand U5100 (N_5100,N_819,N_2357);
xnor U5101 (N_5101,N_1179,N_1218);
nand U5102 (N_5102,N_417,N_1514);
and U5103 (N_5103,N_1871,N_2648);
xor U5104 (N_5104,N_2091,N_321);
nor U5105 (N_5105,N_2504,N_2439);
xnor U5106 (N_5106,N_806,N_1541);
and U5107 (N_5107,N_163,N_1676);
nor U5108 (N_5108,N_669,N_308);
and U5109 (N_5109,N_2649,N_1020);
nor U5110 (N_5110,N_1083,N_526);
or U5111 (N_5111,N_2566,N_634);
and U5112 (N_5112,N_1634,N_1326);
or U5113 (N_5113,N_581,N_2905);
xor U5114 (N_5114,N_929,N_2563);
nor U5115 (N_5115,N_1999,N_2873);
xor U5116 (N_5116,N_455,N_2843);
nand U5117 (N_5117,N_1552,N_2593);
and U5118 (N_5118,N_2377,N_204);
or U5119 (N_5119,N_951,N_773);
and U5120 (N_5120,N_1435,N_1429);
or U5121 (N_5121,N_508,N_387);
or U5122 (N_5122,N_398,N_2011);
nor U5123 (N_5123,N_1817,N_2062);
xnor U5124 (N_5124,N_440,N_530);
xnor U5125 (N_5125,N_882,N_1391);
xor U5126 (N_5126,N_2196,N_429);
and U5127 (N_5127,N_2886,N_559);
and U5128 (N_5128,N_2888,N_2952);
xor U5129 (N_5129,N_554,N_2072);
and U5130 (N_5130,N_2259,N_1400);
nand U5131 (N_5131,N_1496,N_826);
nor U5132 (N_5132,N_631,N_2009);
and U5133 (N_5133,N_1124,N_1728);
nor U5134 (N_5134,N_868,N_219);
nand U5135 (N_5135,N_2385,N_1203);
and U5136 (N_5136,N_388,N_692);
xor U5137 (N_5137,N_1736,N_1359);
or U5138 (N_5138,N_2962,N_1162);
nand U5139 (N_5139,N_2024,N_1709);
or U5140 (N_5140,N_1208,N_813);
xor U5141 (N_5141,N_2925,N_2415);
and U5142 (N_5142,N_525,N_2989);
nor U5143 (N_5143,N_1993,N_2487);
xor U5144 (N_5144,N_1368,N_1241);
and U5145 (N_5145,N_1492,N_2995);
and U5146 (N_5146,N_630,N_2372);
nand U5147 (N_5147,N_357,N_1863);
nor U5148 (N_5148,N_241,N_1524);
or U5149 (N_5149,N_323,N_349);
xnor U5150 (N_5150,N_2649,N_2270);
and U5151 (N_5151,N_486,N_1369);
nand U5152 (N_5152,N_87,N_1070);
nor U5153 (N_5153,N_79,N_2220);
nor U5154 (N_5154,N_868,N_1676);
and U5155 (N_5155,N_1315,N_1361);
xor U5156 (N_5156,N_1433,N_292);
and U5157 (N_5157,N_1586,N_671);
or U5158 (N_5158,N_910,N_1541);
xnor U5159 (N_5159,N_2188,N_857);
nand U5160 (N_5160,N_663,N_2457);
nand U5161 (N_5161,N_1737,N_803);
and U5162 (N_5162,N_1957,N_1655);
xor U5163 (N_5163,N_1551,N_2240);
and U5164 (N_5164,N_2179,N_1826);
nand U5165 (N_5165,N_1702,N_2677);
nand U5166 (N_5166,N_621,N_2124);
or U5167 (N_5167,N_143,N_2933);
nand U5168 (N_5168,N_1125,N_693);
or U5169 (N_5169,N_326,N_1996);
nor U5170 (N_5170,N_1539,N_1472);
and U5171 (N_5171,N_1251,N_1261);
nand U5172 (N_5172,N_90,N_186);
or U5173 (N_5173,N_1868,N_1382);
and U5174 (N_5174,N_1448,N_97);
or U5175 (N_5175,N_2116,N_1388);
and U5176 (N_5176,N_1111,N_2741);
or U5177 (N_5177,N_459,N_2463);
and U5178 (N_5178,N_1332,N_1421);
xnor U5179 (N_5179,N_2389,N_2577);
nand U5180 (N_5180,N_1011,N_2432);
xor U5181 (N_5181,N_1107,N_1046);
and U5182 (N_5182,N_2018,N_2433);
and U5183 (N_5183,N_1035,N_1482);
and U5184 (N_5184,N_1229,N_1463);
xnor U5185 (N_5185,N_2682,N_2328);
or U5186 (N_5186,N_1033,N_2022);
nor U5187 (N_5187,N_1724,N_477);
nand U5188 (N_5188,N_2822,N_2763);
nand U5189 (N_5189,N_1685,N_1977);
nor U5190 (N_5190,N_1973,N_92);
nor U5191 (N_5191,N_615,N_1884);
xor U5192 (N_5192,N_1487,N_200);
and U5193 (N_5193,N_929,N_2027);
and U5194 (N_5194,N_1644,N_1586);
nand U5195 (N_5195,N_1507,N_1546);
xor U5196 (N_5196,N_1266,N_2184);
or U5197 (N_5197,N_1463,N_1068);
xnor U5198 (N_5198,N_2442,N_212);
or U5199 (N_5199,N_194,N_146);
and U5200 (N_5200,N_351,N_451);
nor U5201 (N_5201,N_1732,N_721);
nand U5202 (N_5202,N_1144,N_1442);
nand U5203 (N_5203,N_303,N_539);
and U5204 (N_5204,N_181,N_491);
or U5205 (N_5205,N_2866,N_818);
xnor U5206 (N_5206,N_1418,N_846);
xor U5207 (N_5207,N_875,N_276);
xor U5208 (N_5208,N_197,N_1068);
nand U5209 (N_5209,N_1814,N_2699);
or U5210 (N_5210,N_205,N_2747);
xnor U5211 (N_5211,N_1288,N_1921);
xor U5212 (N_5212,N_1680,N_1115);
nor U5213 (N_5213,N_1358,N_1762);
nand U5214 (N_5214,N_976,N_2604);
nand U5215 (N_5215,N_773,N_1267);
and U5216 (N_5216,N_2986,N_2713);
nand U5217 (N_5217,N_838,N_984);
xnor U5218 (N_5218,N_788,N_346);
nand U5219 (N_5219,N_1630,N_608);
and U5220 (N_5220,N_1697,N_2580);
nand U5221 (N_5221,N_839,N_830);
nor U5222 (N_5222,N_1785,N_1271);
or U5223 (N_5223,N_2811,N_2740);
nor U5224 (N_5224,N_2035,N_832);
nor U5225 (N_5225,N_582,N_1221);
nor U5226 (N_5226,N_182,N_286);
xor U5227 (N_5227,N_2132,N_1168);
and U5228 (N_5228,N_576,N_2860);
or U5229 (N_5229,N_2997,N_991);
nor U5230 (N_5230,N_1951,N_244);
and U5231 (N_5231,N_1574,N_456);
nand U5232 (N_5232,N_123,N_2536);
nand U5233 (N_5233,N_1825,N_1021);
nor U5234 (N_5234,N_2576,N_1261);
or U5235 (N_5235,N_964,N_570);
nand U5236 (N_5236,N_1428,N_1139);
nand U5237 (N_5237,N_2193,N_1569);
nand U5238 (N_5238,N_2038,N_1697);
or U5239 (N_5239,N_2078,N_730);
or U5240 (N_5240,N_1567,N_2734);
nand U5241 (N_5241,N_404,N_1254);
or U5242 (N_5242,N_1392,N_2995);
or U5243 (N_5243,N_2876,N_2883);
xnor U5244 (N_5244,N_199,N_2780);
nand U5245 (N_5245,N_1573,N_1628);
nand U5246 (N_5246,N_988,N_1212);
nand U5247 (N_5247,N_2722,N_659);
or U5248 (N_5248,N_134,N_1991);
xnor U5249 (N_5249,N_929,N_522);
nand U5250 (N_5250,N_1908,N_1673);
nand U5251 (N_5251,N_2413,N_2284);
nand U5252 (N_5252,N_2590,N_2928);
xnor U5253 (N_5253,N_2440,N_2448);
xnor U5254 (N_5254,N_549,N_1014);
or U5255 (N_5255,N_500,N_2971);
or U5256 (N_5256,N_1415,N_621);
or U5257 (N_5257,N_2849,N_2795);
or U5258 (N_5258,N_1639,N_561);
and U5259 (N_5259,N_128,N_891);
xor U5260 (N_5260,N_1544,N_858);
nor U5261 (N_5261,N_2007,N_1376);
nand U5262 (N_5262,N_2287,N_2844);
nor U5263 (N_5263,N_2104,N_96);
nor U5264 (N_5264,N_2173,N_1798);
or U5265 (N_5265,N_2807,N_2264);
nand U5266 (N_5266,N_2406,N_245);
nor U5267 (N_5267,N_1135,N_2150);
nand U5268 (N_5268,N_874,N_2924);
nor U5269 (N_5269,N_1887,N_325);
and U5270 (N_5270,N_1489,N_813);
and U5271 (N_5271,N_2083,N_2674);
or U5272 (N_5272,N_2709,N_16);
xnor U5273 (N_5273,N_2586,N_2205);
and U5274 (N_5274,N_1255,N_473);
and U5275 (N_5275,N_207,N_987);
nor U5276 (N_5276,N_1515,N_1159);
xnor U5277 (N_5277,N_555,N_1103);
or U5278 (N_5278,N_2350,N_1343);
nor U5279 (N_5279,N_587,N_2624);
and U5280 (N_5280,N_314,N_1432);
nor U5281 (N_5281,N_348,N_28);
xor U5282 (N_5282,N_2857,N_72);
nor U5283 (N_5283,N_458,N_753);
nor U5284 (N_5284,N_489,N_2431);
and U5285 (N_5285,N_414,N_1780);
or U5286 (N_5286,N_2313,N_694);
nand U5287 (N_5287,N_148,N_1829);
or U5288 (N_5288,N_146,N_783);
or U5289 (N_5289,N_2805,N_1666);
xnor U5290 (N_5290,N_2489,N_919);
xor U5291 (N_5291,N_226,N_2518);
or U5292 (N_5292,N_2575,N_2509);
or U5293 (N_5293,N_290,N_2458);
or U5294 (N_5294,N_1485,N_254);
nor U5295 (N_5295,N_291,N_2837);
or U5296 (N_5296,N_526,N_2470);
and U5297 (N_5297,N_868,N_1029);
xnor U5298 (N_5298,N_878,N_2124);
nand U5299 (N_5299,N_682,N_2068);
xor U5300 (N_5300,N_1192,N_2740);
and U5301 (N_5301,N_2354,N_2013);
and U5302 (N_5302,N_2436,N_298);
nor U5303 (N_5303,N_1066,N_590);
xor U5304 (N_5304,N_1881,N_1001);
nand U5305 (N_5305,N_1436,N_255);
nand U5306 (N_5306,N_140,N_173);
or U5307 (N_5307,N_1874,N_410);
nor U5308 (N_5308,N_2795,N_2777);
xor U5309 (N_5309,N_1030,N_2513);
or U5310 (N_5310,N_2315,N_2789);
nand U5311 (N_5311,N_2282,N_2172);
or U5312 (N_5312,N_1686,N_2719);
nand U5313 (N_5313,N_1785,N_2616);
or U5314 (N_5314,N_1319,N_1115);
or U5315 (N_5315,N_22,N_1342);
nor U5316 (N_5316,N_2090,N_2706);
nand U5317 (N_5317,N_740,N_46);
and U5318 (N_5318,N_1588,N_2016);
xnor U5319 (N_5319,N_1335,N_194);
and U5320 (N_5320,N_1180,N_2481);
or U5321 (N_5321,N_2491,N_1466);
and U5322 (N_5322,N_1635,N_345);
nand U5323 (N_5323,N_467,N_2035);
xnor U5324 (N_5324,N_198,N_1597);
xnor U5325 (N_5325,N_940,N_1839);
or U5326 (N_5326,N_1259,N_1861);
nand U5327 (N_5327,N_2454,N_1267);
nand U5328 (N_5328,N_1163,N_1243);
or U5329 (N_5329,N_1381,N_547);
nand U5330 (N_5330,N_1886,N_1911);
and U5331 (N_5331,N_2696,N_2810);
nand U5332 (N_5332,N_898,N_2361);
nor U5333 (N_5333,N_2649,N_829);
xnor U5334 (N_5334,N_2362,N_775);
nand U5335 (N_5335,N_819,N_2037);
nor U5336 (N_5336,N_316,N_662);
nor U5337 (N_5337,N_449,N_566);
or U5338 (N_5338,N_1715,N_2161);
xor U5339 (N_5339,N_21,N_431);
nand U5340 (N_5340,N_2647,N_1094);
nand U5341 (N_5341,N_2517,N_2672);
nor U5342 (N_5342,N_2127,N_148);
xor U5343 (N_5343,N_589,N_2888);
nand U5344 (N_5344,N_646,N_2423);
nor U5345 (N_5345,N_2670,N_663);
nor U5346 (N_5346,N_504,N_1306);
nand U5347 (N_5347,N_2070,N_1096);
xnor U5348 (N_5348,N_1737,N_2595);
nand U5349 (N_5349,N_880,N_2041);
or U5350 (N_5350,N_1064,N_2993);
nand U5351 (N_5351,N_2301,N_1105);
or U5352 (N_5352,N_1046,N_747);
nor U5353 (N_5353,N_2787,N_2855);
xnor U5354 (N_5354,N_248,N_466);
or U5355 (N_5355,N_282,N_2243);
or U5356 (N_5356,N_964,N_756);
or U5357 (N_5357,N_261,N_1782);
nand U5358 (N_5358,N_2620,N_148);
nor U5359 (N_5359,N_954,N_2404);
nand U5360 (N_5360,N_1426,N_1559);
xnor U5361 (N_5361,N_100,N_739);
nand U5362 (N_5362,N_652,N_2122);
xor U5363 (N_5363,N_2984,N_1545);
and U5364 (N_5364,N_972,N_2380);
nor U5365 (N_5365,N_2560,N_1532);
or U5366 (N_5366,N_2001,N_1680);
nand U5367 (N_5367,N_2598,N_1234);
xnor U5368 (N_5368,N_1476,N_2387);
nor U5369 (N_5369,N_1621,N_2136);
or U5370 (N_5370,N_592,N_1234);
or U5371 (N_5371,N_639,N_2006);
xor U5372 (N_5372,N_89,N_725);
and U5373 (N_5373,N_2243,N_2831);
nor U5374 (N_5374,N_1447,N_2303);
or U5375 (N_5375,N_1193,N_1104);
nand U5376 (N_5376,N_67,N_1056);
nand U5377 (N_5377,N_302,N_1126);
or U5378 (N_5378,N_2255,N_2590);
nand U5379 (N_5379,N_490,N_2530);
or U5380 (N_5380,N_795,N_2456);
nor U5381 (N_5381,N_112,N_143);
xnor U5382 (N_5382,N_2221,N_1494);
nand U5383 (N_5383,N_2243,N_345);
xor U5384 (N_5384,N_2856,N_2484);
nand U5385 (N_5385,N_1118,N_2127);
xnor U5386 (N_5386,N_1724,N_554);
xor U5387 (N_5387,N_2491,N_426);
xnor U5388 (N_5388,N_1193,N_2200);
xnor U5389 (N_5389,N_648,N_1893);
nand U5390 (N_5390,N_1699,N_247);
nand U5391 (N_5391,N_1613,N_457);
or U5392 (N_5392,N_548,N_2952);
or U5393 (N_5393,N_1638,N_1683);
or U5394 (N_5394,N_417,N_1813);
nor U5395 (N_5395,N_1549,N_233);
nand U5396 (N_5396,N_2985,N_2457);
nor U5397 (N_5397,N_970,N_1271);
nand U5398 (N_5398,N_2539,N_2279);
or U5399 (N_5399,N_1697,N_2346);
nand U5400 (N_5400,N_2853,N_1478);
nor U5401 (N_5401,N_933,N_1414);
xnor U5402 (N_5402,N_2244,N_2257);
or U5403 (N_5403,N_206,N_2254);
nand U5404 (N_5404,N_113,N_1138);
nor U5405 (N_5405,N_2685,N_1479);
and U5406 (N_5406,N_1439,N_191);
and U5407 (N_5407,N_2812,N_209);
nor U5408 (N_5408,N_1941,N_2977);
xor U5409 (N_5409,N_432,N_972);
xnor U5410 (N_5410,N_1580,N_2510);
xor U5411 (N_5411,N_2942,N_2455);
nor U5412 (N_5412,N_410,N_2887);
and U5413 (N_5413,N_1858,N_390);
nor U5414 (N_5414,N_2999,N_18);
nand U5415 (N_5415,N_2513,N_1476);
xor U5416 (N_5416,N_1701,N_843);
and U5417 (N_5417,N_829,N_862);
xor U5418 (N_5418,N_280,N_2635);
nand U5419 (N_5419,N_976,N_1777);
or U5420 (N_5420,N_1359,N_249);
nand U5421 (N_5421,N_2246,N_241);
and U5422 (N_5422,N_2445,N_700);
nand U5423 (N_5423,N_395,N_348);
and U5424 (N_5424,N_1483,N_2975);
nand U5425 (N_5425,N_2132,N_294);
and U5426 (N_5426,N_2141,N_949);
nand U5427 (N_5427,N_1660,N_2139);
xnor U5428 (N_5428,N_611,N_2093);
nand U5429 (N_5429,N_2649,N_213);
nand U5430 (N_5430,N_1767,N_1846);
nand U5431 (N_5431,N_1620,N_1290);
xor U5432 (N_5432,N_2294,N_182);
and U5433 (N_5433,N_1632,N_468);
nand U5434 (N_5434,N_2286,N_2400);
nand U5435 (N_5435,N_455,N_660);
or U5436 (N_5436,N_1812,N_2519);
nand U5437 (N_5437,N_150,N_1442);
or U5438 (N_5438,N_1893,N_2366);
nand U5439 (N_5439,N_788,N_2619);
or U5440 (N_5440,N_2536,N_2508);
nor U5441 (N_5441,N_249,N_2499);
or U5442 (N_5442,N_2204,N_1396);
nor U5443 (N_5443,N_1176,N_645);
nor U5444 (N_5444,N_82,N_1608);
nand U5445 (N_5445,N_130,N_832);
nand U5446 (N_5446,N_2215,N_1849);
or U5447 (N_5447,N_2151,N_870);
xor U5448 (N_5448,N_1593,N_404);
and U5449 (N_5449,N_757,N_2903);
nand U5450 (N_5450,N_551,N_1798);
or U5451 (N_5451,N_721,N_1273);
or U5452 (N_5452,N_73,N_41);
nand U5453 (N_5453,N_2779,N_2534);
nor U5454 (N_5454,N_1440,N_2004);
or U5455 (N_5455,N_2284,N_680);
or U5456 (N_5456,N_2690,N_912);
nor U5457 (N_5457,N_435,N_2209);
nand U5458 (N_5458,N_2366,N_1998);
nand U5459 (N_5459,N_2169,N_1880);
xor U5460 (N_5460,N_1268,N_277);
xnor U5461 (N_5461,N_1185,N_2498);
xnor U5462 (N_5462,N_675,N_2935);
and U5463 (N_5463,N_234,N_258);
and U5464 (N_5464,N_812,N_521);
and U5465 (N_5465,N_610,N_1149);
xnor U5466 (N_5466,N_2755,N_224);
nand U5467 (N_5467,N_1182,N_2784);
nor U5468 (N_5468,N_1582,N_923);
or U5469 (N_5469,N_2428,N_2320);
and U5470 (N_5470,N_1334,N_1654);
and U5471 (N_5471,N_2710,N_525);
and U5472 (N_5472,N_2588,N_2055);
and U5473 (N_5473,N_1125,N_2640);
nor U5474 (N_5474,N_522,N_460);
nand U5475 (N_5475,N_2251,N_496);
and U5476 (N_5476,N_957,N_2803);
nor U5477 (N_5477,N_2248,N_291);
nand U5478 (N_5478,N_2066,N_1650);
xor U5479 (N_5479,N_2835,N_23);
nor U5480 (N_5480,N_2837,N_2807);
nand U5481 (N_5481,N_894,N_2601);
or U5482 (N_5482,N_1581,N_193);
and U5483 (N_5483,N_2658,N_1099);
nand U5484 (N_5484,N_2248,N_2086);
nor U5485 (N_5485,N_1774,N_250);
xnor U5486 (N_5486,N_403,N_1318);
nor U5487 (N_5487,N_1095,N_2605);
nand U5488 (N_5488,N_699,N_1069);
or U5489 (N_5489,N_2251,N_135);
and U5490 (N_5490,N_1712,N_718);
nand U5491 (N_5491,N_2614,N_2494);
nand U5492 (N_5492,N_1624,N_2082);
nor U5493 (N_5493,N_2225,N_1673);
and U5494 (N_5494,N_1702,N_2354);
or U5495 (N_5495,N_1862,N_870);
xor U5496 (N_5496,N_1800,N_1428);
nand U5497 (N_5497,N_1221,N_646);
or U5498 (N_5498,N_966,N_1301);
nor U5499 (N_5499,N_441,N_258);
xnor U5500 (N_5500,N_2825,N_2399);
or U5501 (N_5501,N_1677,N_1801);
or U5502 (N_5502,N_860,N_2221);
nor U5503 (N_5503,N_1927,N_363);
xnor U5504 (N_5504,N_1358,N_258);
nand U5505 (N_5505,N_1524,N_573);
and U5506 (N_5506,N_2571,N_1436);
xor U5507 (N_5507,N_2049,N_1176);
xor U5508 (N_5508,N_1803,N_2141);
xnor U5509 (N_5509,N_1975,N_2343);
xnor U5510 (N_5510,N_327,N_608);
or U5511 (N_5511,N_959,N_10);
xnor U5512 (N_5512,N_153,N_2609);
and U5513 (N_5513,N_1604,N_1341);
nor U5514 (N_5514,N_560,N_2280);
and U5515 (N_5515,N_577,N_1683);
xnor U5516 (N_5516,N_2208,N_14);
or U5517 (N_5517,N_1874,N_1778);
and U5518 (N_5518,N_2509,N_1304);
or U5519 (N_5519,N_2665,N_1623);
and U5520 (N_5520,N_2668,N_22);
and U5521 (N_5521,N_471,N_653);
nand U5522 (N_5522,N_608,N_2114);
or U5523 (N_5523,N_1619,N_2226);
or U5524 (N_5524,N_2794,N_1546);
and U5525 (N_5525,N_554,N_2920);
nand U5526 (N_5526,N_2957,N_368);
and U5527 (N_5527,N_626,N_1151);
nand U5528 (N_5528,N_1592,N_2018);
or U5529 (N_5529,N_2646,N_123);
and U5530 (N_5530,N_1568,N_1026);
and U5531 (N_5531,N_47,N_1000);
nand U5532 (N_5532,N_707,N_1124);
xnor U5533 (N_5533,N_994,N_1854);
and U5534 (N_5534,N_733,N_2805);
or U5535 (N_5535,N_364,N_288);
nor U5536 (N_5536,N_2271,N_2689);
or U5537 (N_5537,N_497,N_1681);
or U5538 (N_5538,N_1353,N_1604);
nor U5539 (N_5539,N_846,N_2394);
xor U5540 (N_5540,N_2053,N_692);
nand U5541 (N_5541,N_640,N_1951);
and U5542 (N_5542,N_696,N_2398);
xor U5543 (N_5543,N_1153,N_134);
nand U5544 (N_5544,N_2848,N_952);
xor U5545 (N_5545,N_128,N_28);
nor U5546 (N_5546,N_2495,N_2700);
or U5547 (N_5547,N_2387,N_390);
nand U5548 (N_5548,N_1871,N_1851);
or U5549 (N_5549,N_998,N_1043);
xnor U5550 (N_5550,N_18,N_1539);
or U5551 (N_5551,N_2528,N_2501);
or U5552 (N_5552,N_2820,N_1380);
nand U5553 (N_5553,N_1076,N_2482);
and U5554 (N_5554,N_2050,N_870);
xor U5555 (N_5555,N_1581,N_53);
and U5556 (N_5556,N_2187,N_1510);
and U5557 (N_5557,N_2412,N_1303);
nand U5558 (N_5558,N_2033,N_324);
xor U5559 (N_5559,N_1107,N_2638);
nand U5560 (N_5560,N_1103,N_2035);
or U5561 (N_5561,N_2246,N_1080);
nor U5562 (N_5562,N_1682,N_1817);
and U5563 (N_5563,N_304,N_528);
xnor U5564 (N_5564,N_931,N_1966);
nand U5565 (N_5565,N_1119,N_125);
or U5566 (N_5566,N_980,N_1581);
xnor U5567 (N_5567,N_1757,N_643);
nand U5568 (N_5568,N_2363,N_1704);
xor U5569 (N_5569,N_1141,N_2912);
nor U5570 (N_5570,N_1286,N_2000);
xor U5571 (N_5571,N_1162,N_1253);
and U5572 (N_5572,N_567,N_2183);
nor U5573 (N_5573,N_282,N_1790);
xor U5574 (N_5574,N_2644,N_913);
xor U5575 (N_5575,N_1780,N_729);
xor U5576 (N_5576,N_306,N_1954);
nand U5577 (N_5577,N_2819,N_880);
nor U5578 (N_5578,N_1769,N_679);
or U5579 (N_5579,N_241,N_880);
and U5580 (N_5580,N_2029,N_1704);
nor U5581 (N_5581,N_2453,N_1872);
nand U5582 (N_5582,N_857,N_1274);
xnor U5583 (N_5583,N_448,N_2915);
or U5584 (N_5584,N_1781,N_1650);
or U5585 (N_5585,N_853,N_1950);
or U5586 (N_5586,N_395,N_1240);
nand U5587 (N_5587,N_1062,N_892);
and U5588 (N_5588,N_221,N_248);
xnor U5589 (N_5589,N_1970,N_2091);
xor U5590 (N_5590,N_2364,N_1006);
or U5591 (N_5591,N_1170,N_99);
nand U5592 (N_5592,N_1447,N_2984);
or U5593 (N_5593,N_2415,N_1796);
nor U5594 (N_5594,N_1906,N_757);
nand U5595 (N_5595,N_467,N_2461);
and U5596 (N_5596,N_2174,N_650);
and U5597 (N_5597,N_881,N_595);
and U5598 (N_5598,N_905,N_353);
and U5599 (N_5599,N_502,N_1855);
or U5600 (N_5600,N_265,N_1977);
nand U5601 (N_5601,N_1933,N_1931);
and U5602 (N_5602,N_39,N_2411);
and U5603 (N_5603,N_2242,N_2257);
and U5604 (N_5604,N_2522,N_1116);
xor U5605 (N_5605,N_2112,N_2220);
nor U5606 (N_5606,N_1717,N_1748);
and U5607 (N_5607,N_102,N_2782);
and U5608 (N_5608,N_384,N_2504);
and U5609 (N_5609,N_2766,N_2971);
nor U5610 (N_5610,N_2487,N_1332);
nand U5611 (N_5611,N_1649,N_1016);
and U5612 (N_5612,N_775,N_1895);
xnor U5613 (N_5613,N_2678,N_2234);
xor U5614 (N_5614,N_775,N_1016);
and U5615 (N_5615,N_2890,N_1782);
nand U5616 (N_5616,N_1217,N_2890);
or U5617 (N_5617,N_1543,N_1026);
nand U5618 (N_5618,N_2826,N_1371);
xnor U5619 (N_5619,N_200,N_1318);
nor U5620 (N_5620,N_625,N_245);
xnor U5621 (N_5621,N_86,N_147);
xor U5622 (N_5622,N_1293,N_2610);
xor U5623 (N_5623,N_1214,N_1);
and U5624 (N_5624,N_1319,N_1555);
and U5625 (N_5625,N_269,N_1148);
and U5626 (N_5626,N_2294,N_1835);
xor U5627 (N_5627,N_1426,N_1154);
nand U5628 (N_5628,N_679,N_1457);
xnor U5629 (N_5629,N_1244,N_630);
xor U5630 (N_5630,N_2287,N_451);
nor U5631 (N_5631,N_432,N_2228);
or U5632 (N_5632,N_547,N_613);
nor U5633 (N_5633,N_2280,N_2792);
xnor U5634 (N_5634,N_2977,N_1729);
or U5635 (N_5635,N_2683,N_264);
or U5636 (N_5636,N_586,N_166);
nor U5637 (N_5637,N_772,N_2535);
and U5638 (N_5638,N_1716,N_2956);
nor U5639 (N_5639,N_2227,N_1647);
xnor U5640 (N_5640,N_851,N_1965);
or U5641 (N_5641,N_234,N_1323);
and U5642 (N_5642,N_796,N_899);
or U5643 (N_5643,N_1091,N_1755);
or U5644 (N_5644,N_2294,N_1796);
nor U5645 (N_5645,N_632,N_377);
nor U5646 (N_5646,N_1752,N_1112);
and U5647 (N_5647,N_1865,N_2271);
and U5648 (N_5648,N_1560,N_201);
or U5649 (N_5649,N_2400,N_8);
nor U5650 (N_5650,N_1455,N_1777);
xnor U5651 (N_5651,N_1964,N_46);
and U5652 (N_5652,N_977,N_2327);
or U5653 (N_5653,N_1835,N_2168);
xnor U5654 (N_5654,N_2738,N_2148);
xor U5655 (N_5655,N_1635,N_2705);
xor U5656 (N_5656,N_433,N_2023);
nand U5657 (N_5657,N_310,N_715);
nor U5658 (N_5658,N_2537,N_2478);
and U5659 (N_5659,N_992,N_2454);
nand U5660 (N_5660,N_2440,N_652);
nand U5661 (N_5661,N_73,N_2522);
and U5662 (N_5662,N_2419,N_76);
or U5663 (N_5663,N_2256,N_324);
xor U5664 (N_5664,N_241,N_1580);
nor U5665 (N_5665,N_2981,N_1530);
and U5666 (N_5666,N_2484,N_1984);
or U5667 (N_5667,N_2053,N_72);
nand U5668 (N_5668,N_1689,N_2566);
and U5669 (N_5669,N_1005,N_762);
nand U5670 (N_5670,N_2311,N_2220);
nor U5671 (N_5671,N_1184,N_571);
xor U5672 (N_5672,N_2644,N_356);
xor U5673 (N_5673,N_1202,N_2362);
xnor U5674 (N_5674,N_2557,N_431);
and U5675 (N_5675,N_1908,N_646);
xnor U5676 (N_5676,N_706,N_1731);
nand U5677 (N_5677,N_1973,N_1980);
nor U5678 (N_5678,N_733,N_1446);
nand U5679 (N_5679,N_2732,N_486);
nor U5680 (N_5680,N_2322,N_197);
nor U5681 (N_5681,N_120,N_1048);
xnor U5682 (N_5682,N_2077,N_2440);
nor U5683 (N_5683,N_592,N_757);
nor U5684 (N_5684,N_1539,N_860);
and U5685 (N_5685,N_2951,N_352);
and U5686 (N_5686,N_1100,N_988);
xor U5687 (N_5687,N_319,N_2508);
or U5688 (N_5688,N_679,N_1417);
nor U5689 (N_5689,N_1369,N_1105);
and U5690 (N_5690,N_764,N_979);
and U5691 (N_5691,N_1565,N_2025);
and U5692 (N_5692,N_2804,N_2460);
and U5693 (N_5693,N_690,N_2614);
xor U5694 (N_5694,N_1901,N_1522);
nor U5695 (N_5695,N_2475,N_1431);
nor U5696 (N_5696,N_2081,N_1852);
nand U5697 (N_5697,N_2108,N_695);
or U5698 (N_5698,N_2101,N_1639);
and U5699 (N_5699,N_303,N_2884);
xnor U5700 (N_5700,N_2761,N_1511);
or U5701 (N_5701,N_2658,N_2397);
and U5702 (N_5702,N_2711,N_430);
xnor U5703 (N_5703,N_2165,N_500);
nand U5704 (N_5704,N_2913,N_688);
or U5705 (N_5705,N_1541,N_274);
nand U5706 (N_5706,N_2757,N_329);
or U5707 (N_5707,N_2850,N_834);
nand U5708 (N_5708,N_2380,N_1581);
or U5709 (N_5709,N_2624,N_1169);
xor U5710 (N_5710,N_2665,N_1885);
or U5711 (N_5711,N_2565,N_2897);
nand U5712 (N_5712,N_1667,N_111);
nor U5713 (N_5713,N_319,N_1356);
xnor U5714 (N_5714,N_2770,N_2261);
or U5715 (N_5715,N_2819,N_2426);
xnor U5716 (N_5716,N_2539,N_2583);
xnor U5717 (N_5717,N_234,N_565);
xnor U5718 (N_5718,N_1801,N_596);
nor U5719 (N_5719,N_28,N_1858);
nor U5720 (N_5720,N_2746,N_168);
or U5721 (N_5721,N_1022,N_1772);
or U5722 (N_5722,N_182,N_1457);
xor U5723 (N_5723,N_1895,N_315);
or U5724 (N_5724,N_785,N_1339);
xnor U5725 (N_5725,N_90,N_1985);
and U5726 (N_5726,N_2611,N_451);
and U5727 (N_5727,N_1525,N_1603);
xnor U5728 (N_5728,N_1245,N_1584);
nor U5729 (N_5729,N_1356,N_370);
and U5730 (N_5730,N_564,N_1306);
or U5731 (N_5731,N_1082,N_1281);
xnor U5732 (N_5732,N_483,N_2724);
nor U5733 (N_5733,N_2725,N_1657);
and U5734 (N_5734,N_1173,N_2959);
and U5735 (N_5735,N_715,N_641);
or U5736 (N_5736,N_2813,N_107);
and U5737 (N_5737,N_485,N_2438);
or U5738 (N_5738,N_2261,N_673);
and U5739 (N_5739,N_140,N_1071);
or U5740 (N_5740,N_783,N_2860);
nor U5741 (N_5741,N_145,N_2357);
or U5742 (N_5742,N_2733,N_1128);
nand U5743 (N_5743,N_2817,N_1012);
and U5744 (N_5744,N_782,N_1092);
nor U5745 (N_5745,N_776,N_1201);
and U5746 (N_5746,N_440,N_509);
nand U5747 (N_5747,N_429,N_2557);
xor U5748 (N_5748,N_663,N_1363);
nor U5749 (N_5749,N_2745,N_2870);
nor U5750 (N_5750,N_1252,N_1769);
xor U5751 (N_5751,N_1514,N_1691);
and U5752 (N_5752,N_28,N_2190);
and U5753 (N_5753,N_1184,N_955);
or U5754 (N_5754,N_1340,N_2385);
nor U5755 (N_5755,N_2522,N_1849);
or U5756 (N_5756,N_572,N_146);
xor U5757 (N_5757,N_704,N_658);
nor U5758 (N_5758,N_440,N_638);
xor U5759 (N_5759,N_217,N_2877);
nand U5760 (N_5760,N_2537,N_1399);
or U5761 (N_5761,N_889,N_49);
nor U5762 (N_5762,N_2198,N_429);
xnor U5763 (N_5763,N_222,N_2557);
and U5764 (N_5764,N_1809,N_1256);
nor U5765 (N_5765,N_467,N_2682);
and U5766 (N_5766,N_1604,N_1586);
and U5767 (N_5767,N_1426,N_2990);
xor U5768 (N_5768,N_46,N_2438);
nor U5769 (N_5769,N_2699,N_1963);
nor U5770 (N_5770,N_1340,N_2461);
and U5771 (N_5771,N_2918,N_797);
xor U5772 (N_5772,N_1970,N_739);
and U5773 (N_5773,N_515,N_1934);
nor U5774 (N_5774,N_2067,N_2670);
or U5775 (N_5775,N_2779,N_413);
or U5776 (N_5776,N_754,N_1924);
and U5777 (N_5777,N_2825,N_1645);
nand U5778 (N_5778,N_47,N_798);
or U5779 (N_5779,N_595,N_924);
and U5780 (N_5780,N_952,N_1367);
nor U5781 (N_5781,N_2041,N_695);
nor U5782 (N_5782,N_2639,N_785);
nor U5783 (N_5783,N_2706,N_2582);
nor U5784 (N_5784,N_21,N_680);
xor U5785 (N_5785,N_494,N_1700);
or U5786 (N_5786,N_2304,N_2531);
and U5787 (N_5787,N_1098,N_1910);
nand U5788 (N_5788,N_593,N_185);
or U5789 (N_5789,N_363,N_2082);
nand U5790 (N_5790,N_1076,N_2545);
and U5791 (N_5791,N_456,N_1006);
nor U5792 (N_5792,N_561,N_658);
xor U5793 (N_5793,N_1425,N_2783);
nand U5794 (N_5794,N_1473,N_2321);
and U5795 (N_5795,N_571,N_2661);
nand U5796 (N_5796,N_1462,N_831);
nor U5797 (N_5797,N_1826,N_493);
nor U5798 (N_5798,N_2821,N_126);
nand U5799 (N_5799,N_156,N_1931);
or U5800 (N_5800,N_913,N_1391);
xnor U5801 (N_5801,N_1342,N_1750);
nand U5802 (N_5802,N_2874,N_2435);
and U5803 (N_5803,N_2612,N_1408);
nor U5804 (N_5804,N_487,N_801);
nand U5805 (N_5805,N_392,N_1246);
or U5806 (N_5806,N_596,N_1131);
and U5807 (N_5807,N_2276,N_2722);
nor U5808 (N_5808,N_1722,N_503);
nand U5809 (N_5809,N_1266,N_98);
nor U5810 (N_5810,N_2882,N_1586);
nand U5811 (N_5811,N_2181,N_1411);
and U5812 (N_5812,N_758,N_2122);
or U5813 (N_5813,N_1063,N_2937);
nand U5814 (N_5814,N_2324,N_2147);
and U5815 (N_5815,N_2717,N_2150);
or U5816 (N_5816,N_1794,N_25);
xnor U5817 (N_5817,N_441,N_1049);
xnor U5818 (N_5818,N_897,N_147);
nor U5819 (N_5819,N_1037,N_59);
and U5820 (N_5820,N_1834,N_2818);
or U5821 (N_5821,N_208,N_1244);
nand U5822 (N_5822,N_2970,N_2533);
and U5823 (N_5823,N_931,N_2084);
nand U5824 (N_5824,N_127,N_977);
or U5825 (N_5825,N_383,N_2722);
xnor U5826 (N_5826,N_2728,N_1183);
and U5827 (N_5827,N_150,N_1832);
and U5828 (N_5828,N_152,N_2032);
xnor U5829 (N_5829,N_1978,N_2056);
nand U5830 (N_5830,N_2398,N_422);
or U5831 (N_5831,N_1976,N_1176);
xnor U5832 (N_5832,N_1041,N_302);
nand U5833 (N_5833,N_2330,N_2921);
or U5834 (N_5834,N_2624,N_929);
nand U5835 (N_5835,N_2150,N_1288);
nand U5836 (N_5836,N_1975,N_2680);
nand U5837 (N_5837,N_2883,N_526);
nand U5838 (N_5838,N_837,N_434);
nor U5839 (N_5839,N_969,N_712);
nand U5840 (N_5840,N_2975,N_1347);
nand U5841 (N_5841,N_2500,N_2370);
and U5842 (N_5842,N_1304,N_855);
or U5843 (N_5843,N_1087,N_2097);
xor U5844 (N_5844,N_44,N_15);
and U5845 (N_5845,N_1117,N_2181);
nand U5846 (N_5846,N_2935,N_612);
nand U5847 (N_5847,N_1750,N_564);
nand U5848 (N_5848,N_1953,N_1562);
or U5849 (N_5849,N_1502,N_233);
xnor U5850 (N_5850,N_149,N_1005);
nor U5851 (N_5851,N_499,N_2741);
xnor U5852 (N_5852,N_2565,N_736);
and U5853 (N_5853,N_455,N_2381);
xnor U5854 (N_5854,N_2229,N_2899);
or U5855 (N_5855,N_2157,N_925);
or U5856 (N_5856,N_1987,N_2659);
nand U5857 (N_5857,N_209,N_1225);
or U5858 (N_5858,N_1858,N_183);
and U5859 (N_5859,N_1997,N_925);
or U5860 (N_5860,N_1357,N_2898);
and U5861 (N_5861,N_373,N_2327);
nor U5862 (N_5862,N_1162,N_196);
xor U5863 (N_5863,N_1568,N_440);
nor U5864 (N_5864,N_1668,N_2548);
and U5865 (N_5865,N_1635,N_712);
and U5866 (N_5866,N_545,N_2600);
nand U5867 (N_5867,N_2387,N_1530);
xor U5868 (N_5868,N_944,N_2562);
xnor U5869 (N_5869,N_1872,N_352);
and U5870 (N_5870,N_1654,N_577);
xor U5871 (N_5871,N_2972,N_1371);
xnor U5872 (N_5872,N_184,N_1979);
nor U5873 (N_5873,N_178,N_2034);
or U5874 (N_5874,N_1934,N_763);
and U5875 (N_5875,N_939,N_465);
xnor U5876 (N_5876,N_1678,N_1831);
nor U5877 (N_5877,N_1838,N_363);
or U5878 (N_5878,N_1677,N_2435);
nand U5879 (N_5879,N_135,N_1128);
or U5880 (N_5880,N_2241,N_74);
xnor U5881 (N_5881,N_2503,N_2415);
nand U5882 (N_5882,N_35,N_1559);
or U5883 (N_5883,N_2579,N_64);
nand U5884 (N_5884,N_205,N_1091);
and U5885 (N_5885,N_2678,N_2849);
nor U5886 (N_5886,N_502,N_1457);
nand U5887 (N_5887,N_1240,N_1443);
nand U5888 (N_5888,N_1321,N_901);
xnor U5889 (N_5889,N_867,N_2468);
or U5890 (N_5890,N_709,N_2606);
xor U5891 (N_5891,N_784,N_1186);
nor U5892 (N_5892,N_2585,N_1015);
and U5893 (N_5893,N_2704,N_1113);
nor U5894 (N_5894,N_1353,N_52);
nor U5895 (N_5895,N_110,N_1109);
nand U5896 (N_5896,N_2763,N_2910);
and U5897 (N_5897,N_1113,N_2514);
and U5898 (N_5898,N_181,N_2961);
nand U5899 (N_5899,N_636,N_858);
nor U5900 (N_5900,N_870,N_1897);
xnor U5901 (N_5901,N_2568,N_700);
nand U5902 (N_5902,N_2970,N_2603);
xor U5903 (N_5903,N_347,N_2005);
xor U5904 (N_5904,N_1667,N_2536);
xnor U5905 (N_5905,N_818,N_2173);
or U5906 (N_5906,N_2044,N_574);
and U5907 (N_5907,N_2912,N_2020);
nor U5908 (N_5908,N_1386,N_1309);
and U5909 (N_5909,N_1965,N_2926);
xnor U5910 (N_5910,N_821,N_2688);
xor U5911 (N_5911,N_2910,N_2315);
nor U5912 (N_5912,N_2154,N_495);
nand U5913 (N_5913,N_1044,N_2557);
nor U5914 (N_5914,N_1069,N_89);
xnor U5915 (N_5915,N_363,N_1561);
xnor U5916 (N_5916,N_747,N_2221);
xnor U5917 (N_5917,N_112,N_403);
nor U5918 (N_5918,N_168,N_2393);
xnor U5919 (N_5919,N_1422,N_2029);
xnor U5920 (N_5920,N_1764,N_568);
or U5921 (N_5921,N_893,N_1370);
nor U5922 (N_5922,N_2075,N_1454);
xor U5923 (N_5923,N_2772,N_2579);
nand U5924 (N_5924,N_713,N_235);
xor U5925 (N_5925,N_2624,N_706);
nand U5926 (N_5926,N_921,N_1067);
nor U5927 (N_5927,N_936,N_147);
nand U5928 (N_5928,N_1958,N_407);
nand U5929 (N_5929,N_289,N_2008);
xor U5930 (N_5930,N_1326,N_702);
or U5931 (N_5931,N_133,N_2852);
and U5932 (N_5932,N_88,N_2976);
or U5933 (N_5933,N_1478,N_543);
and U5934 (N_5934,N_519,N_1229);
xor U5935 (N_5935,N_968,N_1824);
xor U5936 (N_5936,N_1166,N_2913);
or U5937 (N_5937,N_2051,N_2583);
nor U5938 (N_5938,N_1868,N_2541);
nand U5939 (N_5939,N_150,N_642);
and U5940 (N_5940,N_2579,N_2716);
and U5941 (N_5941,N_614,N_546);
or U5942 (N_5942,N_2217,N_879);
xor U5943 (N_5943,N_130,N_1184);
nor U5944 (N_5944,N_1987,N_1923);
xor U5945 (N_5945,N_1714,N_1431);
or U5946 (N_5946,N_1095,N_2741);
and U5947 (N_5947,N_2792,N_573);
and U5948 (N_5948,N_2026,N_1691);
and U5949 (N_5949,N_2813,N_2434);
or U5950 (N_5950,N_989,N_1181);
or U5951 (N_5951,N_2732,N_2570);
or U5952 (N_5952,N_1819,N_2163);
and U5953 (N_5953,N_122,N_2962);
nor U5954 (N_5954,N_1397,N_1608);
and U5955 (N_5955,N_1812,N_2777);
nand U5956 (N_5956,N_1853,N_81);
and U5957 (N_5957,N_78,N_2221);
and U5958 (N_5958,N_756,N_1072);
nor U5959 (N_5959,N_1778,N_796);
xor U5960 (N_5960,N_1199,N_2997);
or U5961 (N_5961,N_83,N_247);
and U5962 (N_5962,N_1766,N_2064);
and U5963 (N_5963,N_1752,N_1024);
nand U5964 (N_5964,N_944,N_1191);
nor U5965 (N_5965,N_829,N_2300);
xnor U5966 (N_5966,N_2040,N_269);
nor U5967 (N_5967,N_890,N_2615);
and U5968 (N_5968,N_1804,N_1886);
or U5969 (N_5969,N_1053,N_1471);
nand U5970 (N_5970,N_1078,N_1752);
and U5971 (N_5971,N_278,N_1693);
or U5972 (N_5972,N_518,N_2729);
nor U5973 (N_5973,N_2882,N_529);
nor U5974 (N_5974,N_2868,N_2768);
and U5975 (N_5975,N_2501,N_320);
xor U5976 (N_5976,N_2989,N_637);
xor U5977 (N_5977,N_1540,N_1521);
xor U5978 (N_5978,N_224,N_1764);
nand U5979 (N_5979,N_1424,N_470);
nor U5980 (N_5980,N_1917,N_1167);
xnor U5981 (N_5981,N_2620,N_639);
or U5982 (N_5982,N_2825,N_2600);
and U5983 (N_5983,N_2255,N_2983);
nor U5984 (N_5984,N_1066,N_656);
nand U5985 (N_5985,N_2351,N_792);
xor U5986 (N_5986,N_295,N_806);
or U5987 (N_5987,N_2748,N_109);
nor U5988 (N_5988,N_2730,N_2636);
nor U5989 (N_5989,N_2826,N_1309);
nand U5990 (N_5990,N_2489,N_2017);
xnor U5991 (N_5991,N_1455,N_1892);
or U5992 (N_5992,N_1786,N_1823);
nor U5993 (N_5993,N_2776,N_1847);
nor U5994 (N_5994,N_954,N_1208);
and U5995 (N_5995,N_461,N_2968);
nor U5996 (N_5996,N_2068,N_1320);
nand U5997 (N_5997,N_2382,N_2517);
nor U5998 (N_5998,N_1565,N_2052);
and U5999 (N_5999,N_2551,N_1267);
nand U6000 (N_6000,N_5924,N_4976);
nand U6001 (N_6001,N_4050,N_3884);
xor U6002 (N_6002,N_4618,N_3926);
and U6003 (N_6003,N_5237,N_4583);
or U6004 (N_6004,N_3063,N_3402);
nor U6005 (N_6005,N_5517,N_5164);
or U6006 (N_6006,N_5484,N_4448);
xor U6007 (N_6007,N_4750,N_4310);
nor U6008 (N_6008,N_4646,N_3578);
and U6009 (N_6009,N_3454,N_3825);
or U6010 (N_6010,N_5615,N_4185);
xor U6011 (N_6011,N_4862,N_4198);
or U6012 (N_6012,N_3896,N_4298);
and U6013 (N_6013,N_5243,N_3904);
or U6014 (N_6014,N_5144,N_4777);
and U6015 (N_6015,N_4598,N_4799);
nor U6016 (N_6016,N_5651,N_4032);
xnor U6017 (N_6017,N_5664,N_3324);
xor U6018 (N_6018,N_4007,N_4359);
xor U6019 (N_6019,N_3134,N_5897);
nand U6020 (N_6020,N_3009,N_4140);
nand U6021 (N_6021,N_5832,N_4278);
nand U6022 (N_6022,N_4654,N_5327);
and U6023 (N_6023,N_3546,N_5479);
nor U6024 (N_6024,N_4605,N_5362);
and U6025 (N_6025,N_4116,N_5351);
xor U6026 (N_6026,N_3483,N_5815);
nand U6027 (N_6027,N_4016,N_4131);
xor U6028 (N_6028,N_5223,N_4866);
nand U6029 (N_6029,N_3087,N_4308);
nand U6030 (N_6030,N_5538,N_4912);
nand U6031 (N_6031,N_3777,N_3301);
or U6032 (N_6032,N_3507,N_5563);
or U6033 (N_6033,N_3580,N_3760);
and U6034 (N_6034,N_4699,N_5839);
nand U6035 (N_6035,N_5930,N_3560);
nand U6036 (N_6036,N_5017,N_5512);
nand U6037 (N_6037,N_5444,N_5738);
and U6038 (N_6038,N_3733,N_3433);
nor U6039 (N_6039,N_5572,N_4965);
or U6040 (N_6040,N_3807,N_5697);
xnor U6041 (N_6041,N_5357,N_3321);
nand U6042 (N_6042,N_5993,N_5313);
xnor U6043 (N_6043,N_5483,N_5730);
nand U6044 (N_6044,N_3533,N_4571);
nor U6045 (N_6045,N_5957,N_5435);
and U6046 (N_6046,N_5079,N_3119);
nor U6047 (N_6047,N_4877,N_3252);
and U6048 (N_6048,N_5946,N_4405);
and U6049 (N_6049,N_4521,N_4462);
nand U6050 (N_6050,N_3864,N_3923);
nand U6051 (N_6051,N_4668,N_5699);
xnor U6052 (N_6052,N_4361,N_4392);
and U6053 (N_6053,N_4441,N_4080);
nand U6054 (N_6054,N_5727,N_3334);
xor U6055 (N_6055,N_5352,N_4005);
xnor U6056 (N_6056,N_4536,N_4388);
and U6057 (N_6057,N_3770,N_5658);
nand U6058 (N_6058,N_5912,N_5662);
xnor U6059 (N_6059,N_4487,N_3136);
nor U6060 (N_6060,N_3144,N_5659);
xor U6061 (N_6061,N_4286,N_4369);
xor U6062 (N_6062,N_5457,N_5918);
nand U6063 (N_6063,N_5093,N_4404);
xor U6064 (N_6064,N_5272,N_4009);
and U6065 (N_6065,N_4692,N_4003);
nand U6066 (N_6066,N_4440,N_3853);
xor U6067 (N_6067,N_3818,N_4088);
and U6068 (N_6068,N_4191,N_3885);
or U6069 (N_6069,N_3690,N_3429);
nand U6070 (N_6070,N_3931,N_3431);
xor U6071 (N_6071,N_4432,N_4568);
and U6072 (N_6072,N_4613,N_4320);
xnor U6073 (N_6073,N_5940,N_5758);
and U6074 (N_6074,N_3695,N_5577);
nand U6075 (N_6075,N_4386,N_4220);
nor U6076 (N_6076,N_4381,N_5835);
nor U6077 (N_6077,N_4752,N_4218);
nor U6078 (N_6078,N_4451,N_4987);
nor U6079 (N_6079,N_4751,N_3508);
xor U6080 (N_6080,N_3559,N_4450);
or U6081 (N_6081,N_5082,N_3849);
and U6082 (N_6082,N_3435,N_4720);
and U6083 (N_6083,N_4611,N_5455);
nor U6084 (N_6084,N_3499,N_5436);
xnor U6085 (N_6085,N_5083,N_4172);
nor U6086 (N_6086,N_3484,N_4409);
xor U6087 (N_6087,N_4306,N_5129);
and U6088 (N_6088,N_5437,N_3459);
or U6089 (N_6089,N_5076,N_3889);
nand U6090 (N_6090,N_5383,N_4160);
or U6091 (N_6091,N_4921,N_5152);
nand U6092 (N_6092,N_3363,N_3198);
xor U6093 (N_6093,N_4681,N_5911);
xor U6094 (N_6094,N_4721,N_5130);
or U6095 (N_6095,N_5163,N_3469);
nor U6096 (N_6096,N_3290,N_5988);
xnor U6097 (N_6097,N_5258,N_5225);
xnor U6098 (N_6098,N_3295,N_3640);
or U6099 (N_6099,N_4367,N_3018);
or U6100 (N_6100,N_3306,N_4057);
and U6101 (N_6101,N_4424,N_3960);
nand U6102 (N_6102,N_5096,N_5695);
and U6103 (N_6103,N_5778,N_3743);
or U6104 (N_6104,N_4667,N_4727);
nand U6105 (N_6105,N_5863,N_4397);
xor U6106 (N_6106,N_5294,N_5604);
nor U6107 (N_6107,N_4765,N_5330);
nor U6108 (N_6108,N_3123,N_3995);
xnor U6109 (N_6109,N_5286,N_3422);
nand U6110 (N_6110,N_4280,N_5817);
nor U6111 (N_6111,N_3831,N_4798);
and U6112 (N_6112,N_3792,N_3667);
xor U6113 (N_6113,N_5683,N_3031);
and U6114 (N_6114,N_4433,N_3449);
nor U6115 (N_6115,N_3066,N_4851);
and U6116 (N_6116,N_3978,N_3491);
nand U6117 (N_6117,N_4118,N_5112);
or U6118 (N_6118,N_3268,N_4573);
xor U6119 (N_6119,N_4484,N_3922);
and U6120 (N_6120,N_3397,N_4947);
xnor U6121 (N_6121,N_4588,N_4077);
or U6122 (N_6122,N_3972,N_4575);
or U6123 (N_6123,N_5197,N_4844);
and U6124 (N_6124,N_4565,N_4456);
nand U6125 (N_6125,N_5055,N_3901);
or U6126 (N_6126,N_4993,N_4151);
nor U6127 (N_6127,N_5598,N_3999);
or U6128 (N_6128,N_3407,N_5895);
and U6129 (N_6129,N_3586,N_4012);
and U6130 (N_6130,N_4437,N_4744);
xor U6131 (N_6131,N_3045,N_4128);
xnor U6132 (N_6132,N_3079,N_4070);
xor U6133 (N_6133,N_5419,N_4015);
nand U6134 (N_6134,N_3907,N_4674);
or U6135 (N_6135,N_5776,N_5505);
nor U6136 (N_6136,N_4971,N_5760);
xor U6137 (N_6137,N_5767,N_3118);
or U6138 (N_6138,N_5668,N_3065);
xor U6139 (N_6139,N_3364,N_3163);
xnor U6140 (N_6140,N_5217,N_4081);
or U6141 (N_6141,N_4193,N_3354);
nand U6142 (N_6142,N_5627,N_5689);
or U6143 (N_6143,N_5247,N_4855);
nand U6144 (N_6144,N_4497,N_5049);
and U6145 (N_6145,N_5648,N_3406);
nor U6146 (N_6146,N_5004,N_4793);
nor U6147 (N_6147,N_3619,N_3215);
nor U6148 (N_6148,N_5447,N_5690);
or U6149 (N_6149,N_3120,N_4302);
or U6150 (N_6150,N_5291,N_3353);
nor U6151 (N_6151,N_4978,N_3446);
or U6152 (N_6152,N_5820,N_5273);
xnor U6153 (N_6153,N_3730,N_5792);
nand U6154 (N_6154,N_3426,N_4210);
nand U6155 (N_6155,N_5393,N_4443);
or U6156 (N_6156,N_3893,N_4387);
xnor U6157 (N_6157,N_3838,N_3713);
or U6158 (N_6158,N_5931,N_3073);
nand U6159 (N_6159,N_5169,N_3387);
nand U6160 (N_6160,N_4885,N_3418);
nand U6161 (N_6161,N_4600,N_5100);
and U6162 (N_6162,N_3585,N_5873);
nand U6163 (N_6163,N_4335,N_3724);
xnor U6164 (N_6164,N_4835,N_5857);
or U6165 (N_6165,N_5982,N_3094);
nand U6166 (N_6166,N_4147,N_5955);
xor U6167 (N_6167,N_4871,N_3748);
and U6168 (N_6168,N_5408,N_3538);
xor U6169 (N_6169,N_4103,N_5781);
and U6170 (N_6170,N_3764,N_3859);
and U6171 (N_6171,N_4027,N_4511);
xor U6172 (N_6172,N_5644,N_5274);
and U6173 (N_6173,N_5544,N_5080);
or U6174 (N_6174,N_3845,N_4545);
nor U6175 (N_6175,N_4104,N_4828);
and U6176 (N_6176,N_4800,N_5132);
or U6177 (N_6177,N_3808,N_3034);
nand U6178 (N_6178,N_5915,N_4876);
nand U6179 (N_6179,N_5248,N_4966);
xnor U6180 (N_6180,N_5926,N_4469);
nor U6181 (N_6181,N_4833,N_3942);
xor U6182 (N_6182,N_4256,N_5746);
xnor U6183 (N_6183,N_3276,N_5656);
nand U6184 (N_6184,N_3501,N_5963);
and U6185 (N_6185,N_5595,N_4934);
nand U6186 (N_6186,N_4223,N_5747);
nand U6187 (N_6187,N_5711,N_3248);
nand U6188 (N_6188,N_4804,N_3330);
and U6189 (N_6189,N_5126,N_5414);
and U6190 (N_6190,N_5222,N_4636);
xor U6191 (N_6191,N_3027,N_3647);
xnor U6192 (N_6192,N_3361,N_4084);
and U6193 (N_6193,N_3753,N_4709);
xor U6194 (N_6194,N_5947,N_3882);
and U6195 (N_6195,N_4023,N_5710);
nor U6196 (N_6196,N_3540,N_3957);
or U6197 (N_6197,N_3138,N_4235);
nor U6198 (N_6198,N_3490,N_5310);
xnor U6199 (N_6199,N_4132,N_3750);
or U6200 (N_6200,N_3858,N_5023);
or U6201 (N_6201,N_4505,N_4334);
or U6202 (N_6202,N_4465,N_3012);
nand U6203 (N_6203,N_4498,N_3570);
nand U6204 (N_6204,N_5680,N_3661);
xor U6205 (N_6205,N_3379,N_4974);
and U6206 (N_6206,N_5904,N_5087);
xnor U6207 (N_6207,N_5220,N_4282);
or U6208 (N_6208,N_5340,N_5858);
and U6209 (N_6209,N_5501,N_4069);
nand U6210 (N_6210,N_4741,N_3167);
nor U6211 (N_6211,N_3384,N_3180);
and U6212 (N_6212,N_3515,N_3537);
or U6213 (N_6213,N_4449,N_3061);
or U6214 (N_6214,N_3032,N_3178);
or U6215 (N_6215,N_5761,N_4933);
or U6216 (N_6216,N_5521,N_3544);
nor U6217 (N_6217,N_4812,N_5876);
or U6218 (N_6218,N_3480,N_3104);
nor U6219 (N_6219,N_5188,N_5388);
nand U6220 (N_6220,N_3427,N_5688);
xor U6221 (N_6221,N_3679,N_3680);
xor U6222 (N_6222,N_3795,N_5390);
nor U6223 (N_6223,N_4805,N_4427);
nand U6224 (N_6224,N_4346,N_4330);
nor U6225 (N_6225,N_5703,N_5753);
nor U6226 (N_6226,N_3817,N_3157);
nor U6227 (N_6227,N_5072,N_3605);
nand U6228 (N_6228,N_5670,N_4706);
and U6229 (N_6229,N_4595,N_5092);
nand U6230 (N_6230,N_4688,N_4478);
nor U6231 (N_6231,N_5459,N_5614);
nand U6232 (N_6232,N_5938,N_3294);
nand U6233 (N_6233,N_5283,N_3133);
nor U6234 (N_6234,N_5307,N_3039);
xor U6235 (N_6235,N_3368,N_4211);
xor U6236 (N_6236,N_5246,N_5255);
or U6237 (N_6237,N_4466,N_5523);
and U6238 (N_6238,N_5552,N_3323);
and U6239 (N_6239,N_5492,N_3511);
and U6240 (N_6240,N_5431,N_4406);
nor U6241 (N_6241,N_3358,N_5321);
nand U6242 (N_6242,N_3698,N_5530);
or U6243 (N_6243,N_5650,N_5181);
and U6244 (N_6244,N_3708,N_5201);
nand U6245 (N_6245,N_5125,N_5573);
nor U6246 (N_6246,N_5951,N_3542);
xnor U6247 (N_6247,N_4480,N_5516);
nand U6248 (N_6248,N_3500,N_4019);
or U6249 (N_6249,N_5145,N_4593);
or U6250 (N_6250,N_4888,N_3297);
xor U6251 (N_6251,N_3651,N_3359);
and U6252 (N_6252,N_3488,N_3600);
nor U6253 (N_6253,N_4614,N_4953);
xnor U6254 (N_6254,N_5421,N_4420);
xnor U6255 (N_6255,N_3279,N_4893);
nor U6256 (N_6256,N_4663,N_3374);
xor U6257 (N_6257,N_3909,N_5156);
nor U6258 (N_6258,N_5382,N_4470);
and U6259 (N_6259,N_5328,N_4638);
nor U6260 (N_6260,N_4643,N_3865);
xnor U6261 (N_6261,N_3776,N_3932);
nor U6262 (N_6262,N_3399,N_5406);
or U6263 (N_6263,N_4803,N_4790);
xor U6264 (N_6264,N_5852,N_5821);
xor U6265 (N_6265,N_3329,N_3541);
nor U6266 (N_6266,N_3876,N_5187);
or U6267 (N_6267,N_4718,N_4021);
or U6268 (N_6268,N_3934,N_4701);
nand U6269 (N_6269,N_5102,N_3221);
and U6270 (N_6270,N_5645,N_5033);
nand U6271 (N_6271,N_5840,N_5941);
and U6272 (N_6272,N_4990,N_3964);
xor U6273 (N_6273,N_4246,N_4189);
nand U6274 (N_6274,N_3269,N_5039);
nor U6275 (N_6275,N_5816,N_5259);
and U6276 (N_6276,N_5547,N_4891);
and U6277 (N_6277,N_4178,N_4120);
nor U6278 (N_6278,N_3924,N_4779);
and U6279 (N_6279,N_3809,N_4184);
nor U6280 (N_6280,N_3262,N_5734);
xor U6281 (N_6281,N_3420,N_4930);
nand U6282 (N_6282,N_3263,N_3260);
xnor U6283 (N_6283,N_5041,N_4243);
nand U6284 (N_6284,N_5365,N_3883);
or U6285 (N_6285,N_5950,N_3176);
nand U6286 (N_6286,N_5811,N_5115);
or U6287 (N_6287,N_4033,N_5477);
nor U6288 (N_6288,N_3911,N_3028);
xnor U6289 (N_6289,N_5496,N_3556);
and U6290 (N_6290,N_4730,N_3416);
xor U6291 (N_6291,N_3506,N_3342);
nor U6292 (N_6292,N_5589,N_5473);
or U6293 (N_6293,N_5966,N_5822);
xnor U6294 (N_6294,N_3906,N_5846);
xnor U6295 (N_6295,N_4578,N_5588);
nand U6296 (N_6296,N_3971,N_4678);
xnor U6297 (N_6297,N_4053,N_3191);
nand U6298 (N_6298,N_4529,N_3196);
xnor U6299 (N_6299,N_4471,N_4152);
nand U6300 (N_6300,N_4354,N_3746);
xor U6301 (N_6301,N_3707,N_3240);
nor U6302 (N_6302,N_4922,N_5312);
xor U6303 (N_6303,N_5612,N_5134);
xnor U6304 (N_6304,N_5174,N_3436);
or U6305 (N_6305,N_3417,N_3389);
or U6306 (N_6306,N_3203,N_3111);
nor U6307 (N_6307,N_5452,N_4943);
nand U6308 (N_6308,N_4616,N_4687);
nor U6309 (N_6309,N_4910,N_5474);
nor U6310 (N_6310,N_3627,N_5090);
xor U6311 (N_6311,N_4905,N_5366);
or U6312 (N_6312,N_4245,N_4783);
nand U6313 (N_6313,N_5865,N_3947);
nand U6314 (N_6314,N_3109,N_5336);
xor U6315 (N_6315,N_4747,N_3002);
or U6316 (N_6316,N_5642,N_5284);
or U6317 (N_6317,N_5003,N_5551);
xnor U6318 (N_6318,N_4507,N_3970);
nand U6319 (N_6319,N_5304,N_4928);
and U6320 (N_6320,N_3813,N_4055);
and U6321 (N_6321,N_5883,N_5179);
nand U6322 (N_6322,N_3021,N_3386);
xor U6323 (N_6323,N_5341,N_3632);
nor U6324 (N_6324,N_5101,N_3516);
or U6325 (N_6325,N_4807,N_5239);
or U6326 (N_6326,N_3617,N_4683);
nor U6327 (N_6327,N_3582,N_3550);
nor U6328 (N_6328,N_4279,N_3700);
or U6329 (N_6329,N_4760,N_4626);
or U6330 (N_6330,N_5095,N_5277);
nand U6331 (N_6331,N_5066,N_3185);
or U6332 (N_6332,N_5244,N_5303);
or U6333 (N_6333,N_4061,N_5416);
xor U6334 (N_6334,N_4394,N_4766);
xnor U6335 (N_6335,N_4195,N_3315);
nor U6336 (N_6336,N_4827,N_4666);
nor U6337 (N_6337,N_5339,N_4168);
xor U6338 (N_6338,N_5016,N_4272);
or U6339 (N_6339,N_4964,N_5789);
and U6340 (N_6340,N_5649,N_4938);
or U6341 (N_6341,N_3356,N_3505);
nand U6342 (N_6342,N_3930,N_3997);
and U6343 (N_6343,N_4742,N_4731);
xnor U6344 (N_6344,N_5800,N_4292);
and U6345 (N_6345,N_5482,N_4379);
nor U6346 (N_6346,N_4102,N_3232);
nand U6347 (N_6347,N_3567,N_3602);
nand U6348 (N_6348,N_3634,N_3694);
and U6349 (N_6349,N_3638,N_5906);
nor U6350 (N_6350,N_5808,N_4506);
or U6351 (N_6351,N_3457,N_3655);
xnor U6352 (N_6352,N_5995,N_4501);
and U6353 (N_6353,N_3820,N_5866);
and U6354 (N_6354,N_4241,N_3826);
or U6355 (N_6355,N_4517,N_3812);
or U6356 (N_6356,N_5774,N_4148);
nor U6357 (N_6357,N_4818,N_3571);
or U6358 (N_6358,N_3444,N_5043);
xor U6359 (N_6359,N_3986,N_5186);
nand U6360 (N_6360,N_5985,N_4201);
nor U6361 (N_6361,N_5769,N_5685);
xor U6362 (N_6362,N_3058,N_5878);
xor U6363 (N_6363,N_5190,N_4117);
nand U6364 (N_6364,N_4457,N_3141);
xnor U6365 (N_6365,N_4530,N_4299);
or U6366 (N_6366,N_3522,N_4254);
and U6367 (N_6367,N_4360,N_3453);
and U6368 (N_6368,N_3839,N_5133);
nand U6369 (N_6369,N_5607,N_3340);
xnor U6370 (N_6370,N_4740,N_3209);
nor U6371 (N_6371,N_4340,N_5374);
or U6372 (N_6372,N_5917,N_5508);
or U6373 (N_6373,N_5999,N_5624);
nor U6374 (N_6374,N_5293,N_4253);
and U6375 (N_6375,N_5089,N_3662);
or U6376 (N_6376,N_4762,N_4821);
xnor U6377 (N_6377,N_3794,N_3112);
nand U6378 (N_6378,N_5019,N_3769);
or U6379 (N_6379,N_3352,N_3096);
or U6380 (N_6380,N_4635,N_5849);
xnor U6381 (N_6381,N_3313,N_4205);
nor U6382 (N_6382,N_4173,N_3834);
nor U6383 (N_6383,N_4628,N_3062);
or U6384 (N_6384,N_4935,N_4485);
nor U6385 (N_6385,N_5919,N_4436);
nand U6386 (N_6386,N_3390,N_3266);
or U6387 (N_6387,N_5571,N_3071);
xor U6388 (N_6388,N_4534,N_5086);
nor U6389 (N_6389,N_3738,N_5721);
or U6390 (N_6390,N_5661,N_3720);
xor U6391 (N_6391,N_4648,N_4199);
nand U6392 (N_6392,N_5251,N_4587);
and U6393 (N_6393,N_5813,N_5833);
and U6394 (N_6394,N_4854,N_5491);
and U6395 (N_6395,N_3517,N_3519);
nor U6396 (N_6396,N_3304,N_4400);
xor U6397 (N_6397,N_3478,N_3692);
or U6398 (N_6398,N_5135,N_4590);
nor U6399 (N_6399,N_4823,N_4028);
and U6400 (N_6400,N_3015,N_5990);
nor U6401 (N_6401,N_3686,N_5602);
and U6402 (N_6402,N_5018,N_4402);
and U6403 (N_6403,N_3190,N_4244);
nand U6404 (N_6404,N_3347,N_5907);
nor U6405 (N_6405,N_5078,N_3202);
nand U6406 (N_6406,N_4999,N_4474);
nor U6407 (N_6407,N_5226,N_4515);
nand U6408 (N_6408,N_5640,N_3958);
or U6409 (N_6409,N_3524,N_4761);
nor U6410 (N_6410,N_5410,N_3967);
nand U6411 (N_6411,N_3950,N_3333);
xnor U6412 (N_6412,N_5285,N_4916);
nor U6413 (N_6413,N_4035,N_3837);
nand U6414 (N_6414,N_4042,N_5094);
xnor U6415 (N_6415,N_4895,N_5302);
nand U6416 (N_6416,N_4995,N_3588);
nor U6417 (N_6417,N_3056,N_4412);
nor U6418 (N_6418,N_4169,N_5387);
nor U6419 (N_6419,N_4200,N_3914);
or U6420 (N_6420,N_4925,N_5241);
nor U6421 (N_6421,N_3860,N_4094);
or U6422 (N_6422,N_3241,N_4775);
and U6423 (N_6423,N_4984,N_4531);
nor U6424 (N_6424,N_3114,N_5887);
and U6425 (N_6425,N_3534,N_5983);
nor U6426 (N_6426,N_5044,N_5743);
nand U6427 (N_6427,N_3900,N_5507);
or U6428 (N_6428,N_3082,N_4528);
nand U6429 (N_6429,N_5889,N_4736);
xnor U6430 (N_6430,N_4242,N_3216);
nor U6431 (N_6431,N_3367,N_4137);
xor U6432 (N_6432,N_3678,N_3529);
and U6433 (N_6433,N_4870,N_5210);
nand U6434 (N_6434,N_5349,N_5515);
nand U6435 (N_6435,N_5430,N_4525);
nor U6436 (N_6436,N_4228,N_3668);
and U6437 (N_6437,N_3755,N_3395);
or U6438 (N_6438,N_5456,N_3335);
or U6439 (N_6439,N_4945,N_4384);
nor U6440 (N_6440,N_3287,N_4608);
nor U6441 (N_6441,N_3919,N_5830);
xnor U6442 (N_6442,N_3493,N_5757);
nor U6443 (N_6443,N_5218,N_3916);
nand U6444 (N_6444,N_4390,N_5194);
and U6445 (N_6445,N_3767,N_3635);
xor U6446 (N_6446,N_4333,N_5065);
or U6447 (N_6447,N_5981,N_3715);
and U6448 (N_6448,N_3721,N_3803);
or U6449 (N_6449,N_5038,N_3129);
and U6450 (N_6450,N_4060,N_3629);
nand U6451 (N_6451,N_3208,N_4257);
or U6452 (N_6452,N_5289,N_3195);
nand U6453 (N_6453,N_5550,N_4671);
xor U6454 (N_6454,N_3010,N_3380);
nor U6455 (N_6455,N_4723,N_4046);
or U6456 (N_6456,N_4499,N_5070);
or U6457 (N_6457,N_5189,N_3917);
nor U6458 (N_6458,N_5868,N_3394);
or U6459 (N_6459,N_5793,N_5841);
and U6460 (N_6460,N_5411,N_4255);
or U6461 (N_6461,N_4154,N_3574);
nand U6462 (N_6462,N_4038,N_5600);
and U6463 (N_6463,N_5371,N_3348);
xnor U6464 (N_6464,N_4227,N_3150);
nand U6465 (N_6465,N_4261,N_5370);
nor U6466 (N_6466,N_5969,N_3458);
or U6467 (N_6467,N_5593,N_4770);
nand U6468 (N_6468,N_4493,N_4669);
nand U6469 (N_6469,N_5765,N_4323);
nand U6470 (N_6470,N_3025,N_5296);
xor U6471 (N_6471,N_4956,N_3612);
xnor U6472 (N_6472,N_3477,N_5718);
xor U6473 (N_6473,N_4090,N_3944);
nor U6474 (N_6474,N_5057,N_4715);
nor U6475 (N_6475,N_5203,N_3665);
or U6476 (N_6476,N_5796,N_3165);
nor U6477 (N_6477,N_3171,N_4724);
xnor U6478 (N_6478,N_4874,N_4836);
or U6479 (N_6479,N_5991,N_3412);
nand U6480 (N_6480,N_5617,N_3460);
nand U6481 (N_6481,N_4431,N_5827);
nand U6482 (N_6482,N_5570,N_5048);
and U6483 (N_6483,N_4848,N_3110);
or U6484 (N_6484,N_3649,N_4708);
nand U6485 (N_6485,N_5204,N_5771);
nor U6486 (N_6486,N_5696,N_5537);
and U6487 (N_6487,N_4024,N_5104);
and U6488 (N_6488,N_5006,N_5678);
nor U6489 (N_6489,N_5433,N_3193);
nand U6490 (N_6490,N_3965,N_5657);
and U6491 (N_6491,N_5489,N_4358);
and U6492 (N_6492,N_3822,N_3465);
nor U6493 (N_6493,N_3059,N_4625);
or U6494 (N_6494,N_3169,N_4732);
xor U6495 (N_6495,N_4276,N_3789);
and U6496 (N_6496,N_3877,N_5305);
nor U6497 (N_6497,N_4232,N_3331);
nor U6498 (N_6498,N_4725,N_3691);
xor U6499 (N_6499,N_3464,N_5462);
or U6500 (N_6500,N_3681,N_4262);
nor U6501 (N_6501,N_4083,N_3148);
or U6502 (N_6502,N_4759,N_4229);
xnor U6503 (N_6503,N_3797,N_4434);
and U6504 (N_6504,N_3552,N_4087);
and U6505 (N_6505,N_3194,N_4074);
nor U6506 (N_6506,N_4939,N_4789);
nor U6507 (N_6507,N_3953,N_4410);
nand U6508 (N_6508,N_5005,N_3731);
xnor U6509 (N_6509,N_3630,N_4142);
xor U6510 (N_6510,N_5116,N_3131);
nand U6511 (N_6511,N_4351,N_5438);
xor U6512 (N_6512,N_4542,N_3030);
nand U6513 (N_6513,N_4591,N_3577);
or U6514 (N_6514,N_5238,N_4859);
nand U6515 (N_6515,N_5329,N_5785);
or U6516 (N_6516,N_5347,N_4037);
nand U6517 (N_6517,N_4236,N_4651);
nor U6518 (N_6518,N_4632,N_3805);
and U6519 (N_6519,N_3787,N_3174);
nor U6520 (N_6520,N_4543,N_5783);
nand U6521 (N_6521,N_3494,N_3549);
nand U6522 (N_6522,N_5500,N_5001);
nand U6523 (N_6523,N_3286,N_5603);
and U6524 (N_6524,N_4746,N_4603);
or U6525 (N_6525,N_4502,N_3563);
or U6526 (N_6526,N_3564,N_3309);
nand U6527 (N_6527,N_3915,N_5613);
xor U6528 (N_6528,N_5564,N_3020);
and U6529 (N_6529,N_4010,N_3067);
or U6530 (N_6530,N_5219,N_4479);
or U6531 (N_6531,N_4537,N_3962);
and U6532 (N_6532,N_3725,N_5788);
and U6533 (N_6533,N_4890,N_5316);
xor U6534 (N_6534,N_4305,N_5042);
xor U6535 (N_6535,N_3963,N_4064);
xor U6536 (N_6536,N_3992,N_5892);
nand U6537 (N_6537,N_3362,N_5638);
xnor U6538 (N_6538,N_3565,N_5242);
or U6539 (N_6539,N_4670,N_3891);
and U6540 (N_6540,N_5837,N_3413);
nand U6541 (N_6541,N_5844,N_5514);
xor U6542 (N_6542,N_5355,N_5497);
nor U6543 (N_6543,N_4277,N_4264);
xor U6544 (N_6544,N_4810,N_5335);
nand U6545 (N_6545,N_4872,N_4641);
or U6546 (N_6546,N_3461,N_4774);
xor U6547 (N_6547,N_5709,N_4396);
nor U6548 (N_6548,N_3682,N_5937);
xnor U6549 (N_6549,N_4576,N_4086);
or U6550 (N_6550,N_3128,N_4129);
and U6551 (N_6551,N_5441,N_5677);
nand U6552 (N_6552,N_3870,N_4619);
nand U6553 (N_6553,N_3867,N_5737);
xnor U6554 (N_6554,N_4597,N_3637);
or U6555 (N_6555,N_4365,N_5026);
nand U6556 (N_6556,N_5510,N_5494);
xor U6557 (N_6557,N_4353,N_5527);
xnor U6558 (N_6558,N_3130,N_5056);
nor U6559 (N_6559,N_3591,N_5454);
nor U6560 (N_6560,N_3149,N_4689);
xor U6561 (N_6561,N_3227,N_4962);
nor U6562 (N_6562,N_4389,N_4123);
nand U6563 (N_6563,N_3403,N_4979);
or U6564 (N_6564,N_4378,N_5834);
xor U6565 (N_6565,N_3022,N_5900);
and U6566 (N_6566,N_5701,N_5583);
and U6567 (N_6567,N_5403,N_5392);
nand U6568 (N_6568,N_3751,N_5601);
or U6569 (N_6569,N_5319,N_3233);
nand U6570 (N_6570,N_4696,N_5401);
or U6571 (N_6571,N_3863,N_4271);
or U6572 (N_6572,N_4514,N_4284);
and U6573 (N_6573,N_3369,N_3747);
xor U6574 (N_6574,N_3437,N_4644);
xnor U6575 (N_6575,N_5554,N_4882);
xor U6576 (N_6576,N_5625,N_4806);
nor U6577 (N_6577,N_4951,N_3456);
nor U6578 (N_6578,N_5175,N_4426);
xor U6579 (N_6579,N_4937,N_4577);
xor U6580 (N_6580,N_4383,N_5524);
xnor U6581 (N_6581,N_3688,N_5845);
or U6582 (N_6582,N_3595,N_5014);
or U6583 (N_6583,N_5939,N_3675);
nand U6584 (N_6584,N_5205,N_5733);
xor U6585 (N_6585,N_5278,N_3938);
xnor U6586 (N_6586,N_5943,N_3177);
nand U6587 (N_6587,N_4564,N_3523);
xnor U6588 (N_6588,N_4395,N_4138);
xor U6589 (N_6589,N_5252,N_3804);
or U6590 (N_6590,N_3044,N_5030);
nand U6591 (N_6591,N_4940,N_3762);
and U6592 (N_6592,N_5035,N_4461);
or U6593 (N_6593,N_4036,N_3497);
nand U6594 (N_6594,N_5807,N_4734);
xnor U6595 (N_6595,N_4630,N_4749);
and U6596 (N_6596,N_3162,N_5045);
xor U6597 (N_6597,N_4908,N_5348);
and U6598 (N_6598,N_3514,N_3674);
or U6599 (N_6599,N_5215,N_3154);
nor U6600 (N_6600,N_5397,N_5987);
or U6601 (N_6601,N_4980,N_4192);
xnor U6602 (N_6602,N_3443,N_5360);
nor U6603 (N_6603,N_5749,N_3756);
xor U6604 (N_6604,N_5691,N_4071);
or U6605 (N_6605,N_4216,N_4983);
nor U6606 (N_6606,N_3246,N_5605);
nand U6607 (N_6607,N_3543,N_3802);
or U6608 (N_6608,N_5914,N_5575);
or U6609 (N_6609,N_3902,N_5728);
nor U6610 (N_6610,N_4834,N_4658);
nor U6611 (N_6611,N_5493,N_3758);
xor U6612 (N_6612,N_5831,N_5768);
nand U6613 (N_6613,N_3439,N_4541);
and U6614 (N_6614,N_5585,N_5967);
and U6615 (N_6615,N_4230,N_3868);
and U6616 (N_6616,N_5234,N_3055);
or U6617 (N_6617,N_3836,N_4655);
nor U6618 (N_6618,N_4134,N_3928);
nor U6619 (N_6619,N_3083,N_5269);
or U6620 (N_6620,N_4547,N_3685);
or U6621 (N_6621,N_3645,N_5472);
nor U6622 (N_6622,N_4768,N_3869);
xnor U6623 (N_6623,N_4342,N_3146);
xnor U6624 (N_6624,N_5117,N_3894);
xnor U6625 (N_6625,N_3676,N_3985);
xnor U6626 (N_6626,N_5686,N_3466);
and U6627 (N_6627,N_3401,N_4758);
nor U6628 (N_6628,N_3899,N_3937);
xor U6629 (N_6629,N_3790,N_5608);
nor U6630 (N_6630,N_3503,N_4839);
nand U6631 (N_6631,N_4713,N_5470);
nand U6632 (N_6632,N_4554,N_3064);
nor U6633 (N_6633,N_4099,N_4313);
xor U6634 (N_6634,N_4532,N_3013);
or U6635 (N_6635,N_4796,N_3814);
nand U6636 (N_6636,N_5942,N_5535);
nand U6637 (N_6637,N_3145,N_4029);
and U6638 (N_6638,N_5923,N_5182);
xnor U6639 (N_6639,N_3393,N_4550);
nand U6640 (N_6640,N_3448,N_3314);
xnor U6641 (N_6641,N_4300,N_3322);
nor U6642 (N_6642,N_4685,N_4878);
xor U6643 (N_6643,N_5712,N_4837);
and U6644 (N_6644,N_4303,N_4975);
xor U6645 (N_6645,N_4398,N_5268);
nor U6646 (N_6646,N_4902,N_5978);
nor U6647 (N_6647,N_3495,N_5467);
xor U6648 (N_6648,N_5754,N_5693);
nor U6649 (N_6649,N_3719,N_3360);
and U6650 (N_6650,N_4991,N_5287);
nand U6651 (N_6651,N_4321,N_4082);
nor U6652 (N_6652,N_4911,N_3850);
and U6653 (N_6653,N_4156,N_4247);
nor U6654 (N_6654,N_5324,N_4495);
nor U6655 (N_6655,N_5899,N_3918);
nand U6656 (N_6656,N_3656,N_5173);
or U6657 (N_6657,N_5451,N_3801);
and U6658 (N_6658,N_4722,N_3569);
or U6659 (N_6659,N_5980,N_4260);
xor U6660 (N_6660,N_5427,N_3851);
xor U6661 (N_6661,N_3729,N_3613);
nor U6662 (N_6662,N_5464,N_4222);
nor U6663 (N_6663,N_3616,N_3349);
nor U6664 (N_6664,N_5108,N_3788);
nand U6665 (N_6665,N_5097,N_4813);
nand U6666 (N_6666,N_3017,N_5000);
and U6667 (N_6667,N_4920,N_3468);
nand U6668 (N_6668,N_4363,N_4250);
nor U6669 (N_6669,N_3378,N_4560);
or U6670 (N_6670,N_5763,N_3217);
nor U6671 (N_6671,N_3303,N_4336);
or U6672 (N_6672,N_4665,N_3424);
and U6673 (N_6673,N_4091,N_4884);
nor U6674 (N_6674,N_3122,N_5020);
or U6675 (N_6675,N_5128,N_4994);
or U6676 (N_6676,N_5198,N_3626);
or U6677 (N_6677,N_3654,N_5191);
or U6678 (N_6678,N_5619,N_5896);
and U6679 (N_6679,N_4275,N_5700);
nor U6680 (N_6680,N_3475,N_4819);
and U6681 (N_6681,N_5178,N_4107);
nor U6682 (N_6682,N_5984,N_4338);
nor U6683 (N_6683,N_5775,N_5074);
and U6684 (N_6684,N_3547,N_4739);
xor U6685 (N_6685,N_3728,N_3742);
and U6686 (N_6686,N_4136,N_4110);
or U6687 (N_6687,N_3512,N_3008);
nor U6688 (N_6688,N_4815,N_5063);
or U6689 (N_6689,N_3766,N_5460);
xnor U6690 (N_6690,N_5791,N_3732);
and U6691 (N_6691,N_4067,N_4931);
nor U6692 (N_6692,N_5261,N_5587);
nor U6693 (N_6693,N_5770,N_4098);
and U6694 (N_6694,N_3983,N_5681);
nor U6695 (N_6695,N_5211,N_4615);
nand U6696 (N_6696,N_4929,N_3959);
nand U6697 (N_6697,N_5407,N_5511);
and U6698 (N_6698,N_4017,N_5534);
and U6699 (N_6699,N_5081,N_5972);
xnor U6700 (N_6700,N_5334,N_5343);
nand U6701 (N_6701,N_5766,N_5726);
xnor U6702 (N_6702,N_3736,N_3175);
and U6703 (N_6703,N_3341,N_3261);
or U6704 (N_6704,N_3954,N_3687);
or U6705 (N_6705,N_3283,N_5013);
and U6706 (N_6706,N_3878,N_4917);
or U6707 (N_6707,N_5172,N_4675);
nand U6708 (N_6708,N_5012,N_4105);
xnor U6709 (N_6709,N_3855,N_4858);
or U6710 (N_6710,N_4157,N_4782);
xor U6711 (N_6711,N_5356,N_4776);
or U6712 (N_6712,N_3035,N_3592);
xnor U6713 (N_6713,N_5977,N_4781);
and U6714 (N_6714,N_3644,N_5196);
nand U6715 (N_6715,N_3912,N_5461);
nand U6716 (N_6716,N_4438,N_4194);
or U6717 (N_6717,N_3372,N_4362);
or U6718 (N_6718,N_4832,N_3936);
nand U6719 (N_6719,N_3392,N_3327);
nand U6720 (N_6720,N_3821,N_3270);
xor U6721 (N_6721,N_4853,N_5061);
or U6722 (N_6722,N_5903,N_4177);
nand U6723 (N_6723,N_4985,N_5439);
or U6724 (N_6724,N_4586,N_4896);
nand U6725 (N_6725,N_3135,N_4852);
or U6726 (N_6726,N_4439,N_4881);
or U6727 (N_6727,N_5103,N_4735);
nand U6728 (N_6728,N_3973,N_3041);
and U6729 (N_6729,N_3142,N_3624);
nor U6730 (N_6730,N_4401,N_4315);
nand U6731 (N_6731,N_5616,N_5997);
xnor U6732 (N_6732,N_5193,N_4124);
and U6733 (N_6733,N_4755,N_5271);
nand U6734 (N_6734,N_4684,N_3040);
xnor U6735 (N_6735,N_4149,N_4702);
or U6736 (N_6736,N_4416,N_3717);
nand U6737 (N_6737,N_4486,N_5705);
nand U6738 (N_6738,N_4268,N_4428);
nand U6739 (N_6739,N_4122,N_4307);
and U6740 (N_6740,N_5029,N_3173);
or U6741 (N_6741,N_5052,N_4141);
and U6742 (N_6742,N_5610,N_3153);
and U6743 (N_6743,N_4563,N_5120);
xor U6744 (N_6744,N_5959,N_3430);
nand U6745 (N_6745,N_4767,N_3819);
nand U6746 (N_6746,N_5725,N_3242);
nor U6747 (N_6747,N_4309,N_4664);
or U6748 (N_6748,N_5818,N_4592);
nor U6749 (N_6749,N_5965,N_5823);
nor U6750 (N_6750,N_4417,N_3799);
or U6751 (N_6751,N_3255,N_5599);
xnor U6752 (N_6752,N_4519,N_4691);
and U6753 (N_6753,N_5311,N_5558);
xnor U6754 (N_6754,N_4946,N_5184);
or U6755 (N_6755,N_5487,N_5317);
nand U6756 (N_6756,N_4407,N_3614);
nor U6757 (N_6757,N_5626,N_5826);
nor U6758 (N_6758,N_5739,N_5597);
nor U6759 (N_6759,N_4368,N_3741);
or U6760 (N_6760,N_4830,N_5040);
nand U6761 (N_6761,N_4153,N_4014);
and U6762 (N_6762,N_3151,N_4676);
nor U6763 (N_6763,N_4311,N_3187);
and U6764 (N_6764,N_5368,N_4988);
nand U6765 (N_6765,N_5518,N_3103);
or U6766 (N_6766,N_5224,N_5877);
or U6767 (N_6767,N_3476,N_5185);
nand U6768 (N_6768,N_3143,N_5992);
or U6769 (N_6769,N_3816,N_3320);
nand U6770 (N_6770,N_4748,N_4637);
nor U6771 (N_6771,N_3646,N_4695);
nand U6772 (N_6772,N_5594,N_3779);
xnor U6773 (N_6773,N_4329,N_4186);
xnor U6774 (N_6774,N_4549,N_4580);
or U6775 (N_6775,N_5381,N_3496);
or U6776 (N_6776,N_4224,N_4126);
nand U6777 (N_6777,N_3204,N_4838);
xor U6778 (N_6778,N_4072,N_3231);
or U6779 (N_6779,N_5281,N_5232);
and U6780 (N_6780,N_5714,N_5666);
nand U6781 (N_6781,N_4656,N_4040);
nand U6782 (N_6782,N_3830,N_5905);
xor U6783 (N_6783,N_5884,N_4146);
nand U6784 (N_6784,N_3451,N_4737);
or U6785 (N_6785,N_4693,N_4092);
nand U6786 (N_6786,N_3326,N_5933);
xor U6787 (N_6787,N_3156,N_3781);
nand U6788 (N_6788,N_5669,N_5485);
nand U6789 (N_6789,N_3786,N_3298);
xnor U6790 (N_6790,N_3857,N_3621);
nor U6791 (N_6791,N_5663,N_3948);
and U6792 (N_6792,N_3739,N_3943);
xor U6793 (N_6793,N_3113,N_3636);
nand U6794 (N_6794,N_4058,N_3253);
nor U6795 (N_6795,N_5872,N_3265);
and U6796 (N_6796,N_5047,N_3124);
nand U6797 (N_6797,N_4252,N_5973);
and U6798 (N_6798,N_3879,N_3535);
or U6799 (N_6799,N_3050,N_3996);
nor U6800 (N_6800,N_4959,N_4557);
or U6801 (N_6801,N_3474,N_4907);
nor U6802 (N_6802,N_5151,N_5022);
or U6803 (N_6803,N_3054,N_3160);
nor U6804 (N_6804,N_4181,N_5673);
nand U6805 (N_6805,N_5812,N_3498);
or U6806 (N_6806,N_5206,N_5118);
nor U6807 (N_6807,N_4784,N_3740);
nand U6808 (N_6808,N_3951,N_5874);
nand U6809 (N_6809,N_4923,N_4459);
nand U6810 (N_6810,N_4719,N_3081);
xor U6811 (N_6811,N_3292,N_5235);
nand U6812 (N_6812,N_3257,N_3281);
xnor U6813 (N_6813,N_5157,N_5067);
xor U6814 (N_6814,N_4364,N_5565);
xnor U6815 (N_6815,N_4031,N_4944);
or U6816 (N_6816,N_3925,N_3105);
and U6817 (N_6817,N_4538,N_4892);
or U6818 (N_6818,N_4183,N_5875);
nand U6819 (N_6819,N_5476,N_4044);
nor U6820 (N_6820,N_3409,N_5654);
nand U6821 (N_6821,N_4002,N_5794);
nor U6822 (N_6822,N_5806,N_5910);
or U6823 (N_6823,N_5075,N_4559);
or U6824 (N_6824,N_5069,N_5073);
or U6825 (N_6825,N_5025,N_4824);
or U6826 (N_6826,N_4677,N_3371);
nand U6827 (N_6827,N_5921,N_5825);
and U6828 (N_6828,N_4826,N_3554);
and U6829 (N_6829,N_5354,N_4629);
xor U6830 (N_6830,N_4290,N_5176);
or U6831 (N_6831,N_4097,N_5059);
or U6832 (N_6832,N_4763,N_4621);
xnor U6833 (N_6833,N_3840,N_4170);
xnor U6834 (N_6834,N_5622,N_4251);
and U6835 (N_6835,N_5632,N_4982);
and U6836 (N_6836,N_5740,N_5828);
or U6837 (N_6837,N_5639,N_5389);
nand U6838 (N_6838,N_4997,N_5956);
and U6839 (N_6839,N_3927,N_5413);
and U6840 (N_6840,N_4166,N_4831);
xnor U6841 (N_6841,N_4089,N_5885);
xor U6842 (N_6842,N_5869,N_5266);
or U6843 (N_6843,N_4582,N_5975);
and U6844 (N_6844,N_3806,N_3935);
nand U6845 (N_6845,N_3223,N_4144);
and U6846 (N_6846,N_4915,N_4085);
nor U6847 (N_6847,N_5986,N_5429);
nand U6848 (N_6848,N_3189,N_4263);
xnor U6849 (N_6849,N_5799,N_3049);
nor U6850 (N_6850,N_3428,N_4847);
or U6851 (N_6851,N_4453,N_4860);
or U6852 (N_6852,N_3562,N_4544);
nand U6853 (N_6853,N_3432,N_3955);
or U6854 (N_6854,N_4620,N_4355);
nand U6855 (N_6855,N_3798,N_5964);
nand U6856 (N_6856,N_4986,N_4957);
and U6857 (N_6857,N_5809,N_3903);
xnor U6858 (N_6858,N_5528,N_5870);
xor U6859 (N_6859,N_4589,N_4864);
and U6860 (N_6860,N_4889,N_3211);
and U6861 (N_6861,N_4269,N_5715);
nand U6862 (N_6862,N_5143,N_5377);
or U6863 (N_6863,N_4546,N_4522);
xnor U6864 (N_6864,N_3473,N_5114);
or U6865 (N_6865,N_5506,N_3699);
nor U6866 (N_6866,N_4296,N_5288);
nand U6867 (N_6867,N_3452,N_4188);
and U6868 (N_6868,N_4139,N_4000);
nand U6869 (N_6869,N_5053,N_5843);
or U6870 (N_6870,N_5643,N_5723);
xnor U6871 (N_6871,N_3166,N_5195);
nor U6872 (N_6872,N_4288,N_4809);
nor U6873 (N_6873,N_5569,N_5935);
or U6874 (N_6874,N_3583,N_4020);
nor U6875 (N_6875,N_5236,N_4569);
or U6876 (N_6876,N_4270,N_3244);
and U6877 (N_6877,N_5423,N_3611);
nor U6878 (N_6878,N_4458,N_3425);
or U6879 (N_6879,N_5249,N_3579);
or U6880 (N_6880,N_4952,N_4936);
nand U6881 (N_6881,N_5137,N_4345);
xnor U6882 (N_6882,N_3933,N_5560);
or U6883 (N_6883,N_5230,N_5495);
nor U6884 (N_6884,N_3332,N_3274);
and U6885 (N_6885,N_5418,N_4596);
nand U6886 (N_6886,N_4496,N_5748);
xor U6887 (N_6887,N_5141,N_4599);
xor U6888 (N_6888,N_3920,N_4325);
or U6889 (N_6889,N_3152,N_3601);
xnor U6890 (N_6890,N_4393,N_4780);
nand U6891 (N_6891,N_5882,N_3338);
and U6892 (N_6892,N_3026,N_3115);
nor U6893 (N_6893,N_3658,N_5513);
xor U6894 (N_6894,N_5344,N_5221);
nor U6895 (N_6895,N_5432,N_5338);
xnor U6896 (N_6896,N_3043,N_4217);
nand U6897 (N_6897,N_3383,N_4728);
and U6898 (N_6898,N_5051,N_5160);
xor U6899 (N_6899,N_3829,N_4467);
and U6900 (N_6900,N_3979,N_5123);
and U6901 (N_6901,N_3344,N_5756);
nand U6902 (N_6902,N_3357,N_5503);
and U6903 (N_6903,N_3365,N_3080);
nor U6904 (N_6904,N_5536,N_5417);
xnor U6905 (N_6905,N_4662,N_4435);
xnor U6906 (N_6906,N_4846,N_5300);
xor U6907 (N_6907,N_5267,N_4898);
nand U6908 (N_6908,N_4162,N_3184);
or U6909 (N_6909,N_4113,N_4095);
and U6910 (N_6910,N_4682,N_5735);
nand U6911 (N_6911,N_5364,N_4857);
xor U6912 (N_6912,N_5652,N_3404);
nand U6913 (N_6913,N_5148,N_5795);
xor U6914 (N_6914,N_3749,N_5391);
and U6915 (N_6915,N_5893,N_3440);
nor U6916 (N_6916,N_5062,N_5580);
or U6917 (N_6917,N_3672,N_4413);
and U6918 (N_6918,N_5322,N_4421);
and U6919 (N_6919,N_4115,N_4109);
xor U6920 (N_6920,N_4745,N_4764);
and U6921 (N_6921,N_4584,N_3092);
xnor U6922 (N_6922,N_5502,N_5046);
nor U6923 (N_6923,N_3226,N_3328);
xnor U6924 (N_6924,N_3594,N_4447);
nor U6925 (N_6925,N_3945,N_4981);
or U6926 (N_6926,N_5803,N_4969);
and U6927 (N_6927,N_4197,N_5520);
nand U6928 (N_6928,N_4164,N_5136);
nor U6929 (N_6929,N_4204,N_3019);
and U6930 (N_6930,N_5034,N_5146);
nand U6931 (N_6931,N_4743,N_3258);
nand U6932 (N_6932,N_5353,N_5326);
nand U6933 (N_6933,N_3706,N_5111);
xor U6934 (N_6934,N_5110,N_5350);
nor U6935 (N_6935,N_3940,N_4680);
and U6936 (N_6936,N_3201,N_5731);
or U6937 (N_6937,N_4996,N_5546);
xnor U6938 (N_6938,N_3881,N_5227);
nor U6939 (N_6939,N_5253,N_5009);
xor U6940 (N_6940,N_5318,N_3530);
nor U6941 (N_6941,N_3856,N_4645);
nand U6942 (N_6942,N_3006,N_5804);
or U6943 (N_6943,N_3842,N_4145);
or U6944 (N_6944,N_4213,N_3398);
and U6945 (N_6945,N_3998,N_3107);
and U6946 (N_6946,N_3631,N_5819);
and U6947 (N_6947,N_3289,N_4566);
or U6948 (N_6948,N_5909,N_4293);
nor U6949 (N_6949,N_4753,N_3557);
nor U6950 (N_6950,N_3521,N_3974);
or U6951 (N_6951,N_4463,N_5509);
nand U6952 (N_6952,N_5140,N_3023);
nand U6953 (N_6953,N_4623,N_3086);
nor U6954 (N_6954,N_5064,N_3722);
nand U6955 (N_6955,N_3273,N_3408);
nor U6956 (N_6956,N_3016,N_5405);
and U6957 (N_6957,N_4219,N_3259);
or U6958 (N_6958,N_3866,N_3319);
and U6959 (N_6959,N_3783,N_5782);
xor U6960 (N_6960,N_4602,N_5881);
nor U6961 (N_6961,N_5192,N_3975);
or U6962 (N_6962,N_3463,N_4234);
and U6963 (N_6963,N_4845,N_4633);
and U6964 (N_6964,N_3663,N_5584);
xnor U6965 (N_6965,N_3754,N_3852);
and U6966 (N_6966,N_5165,N_4861);
or U6967 (N_6967,N_3137,N_4332);
nor U6968 (N_6968,N_4312,N_4096);
or U6969 (N_6969,N_5200,N_5543);
xor U6970 (N_6970,N_4371,N_4075);
nor U6971 (N_6971,N_4610,N_5526);
or U6972 (N_6972,N_4886,N_5653);
and U6973 (N_6973,N_3757,N_5952);
and U6974 (N_6974,N_5829,N_3705);
nor U6975 (N_6975,N_4647,N_4326);
or U6976 (N_6976,N_3610,N_5091);
or U6977 (N_6977,N_4001,N_5719);
nor U6978 (N_6978,N_3033,N_5106);
xnor U6979 (N_6979,N_3593,N_4237);
xor U6980 (N_6980,N_4317,N_5522);
xor U6981 (N_6981,N_5647,N_4612);
or U6982 (N_6982,N_5631,N_5098);
nor U6983 (N_6983,N_4030,N_4179);
or U6984 (N_6984,N_3875,N_4442);
xor U6985 (N_6985,N_4601,N_3001);
or U6986 (N_6986,N_4322,N_4259);
or U6987 (N_6987,N_3890,N_4825);
xor U6988 (N_6988,N_5412,N_4366);
nor U6989 (N_6989,N_5864,N_3376);
or U6990 (N_6990,N_4130,N_4372);
nor U6991 (N_6991,N_3723,N_4073);
nand U6992 (N_6992,N_4518,N_3158);
and U6993 (N_6993,N_4267,N_3660);
nor U6994 (N_6994,N_5732,N_3659);
nor U6995 (N_6995,N_4509,N_5540);
or U6996 (N_6996,N_5555,N_4553);
and U6997 (N_6997,N_3608,N_5250);
nor U6998 (N_6998,N_4794,N_5445);
xnor U6999 (N_6999,N_3871,N_3046);
or U7000 (N_7000,N_4468,N_5207);
or U7001 (N_7001,N_5139,N_5071);
xor U7002 (N_7002,N_4357,N_5280);
nor U7003 (N_7003,N_4705,N_5861);
xnor U7004 (N_7004,N_3042,N_4331);
nor U7005 (N_7005,N_4158,N_5698);
and U7006 (N_7006,N_3481,N_5480);
and U7007 (N_7007,N_4698,N_4607);
nor U7008 (N_7008,N_3590,N_3941);
and U7009 (N_7009,N_5199,N_3400);
nand U7010 (N_7010,N_4206,N_5214);
or U7011 (N_7011,N_5810,N_5545);
xor U7012 (N_7012,N_4792,N_5088);
nand U7013 (N_7013,N_4998,N_3981);
nor U7014 (N_7014,N_4795,N_5084);
and U7015 (N_7015,N_5836,N_5216);
nand U7016 (N_7016,N_3267,N_3793);
or U7017 (N_7017,N_4101,N_5853);
or U7018 (N_7018,N_5692,N_4555);
xor U7019 (N_7019,N_5934,N_5596);
xor U7020 (N_7020,N_4906,N_5949);
or U7021 (N_7021,N_3815,N_4165);
nand U7022 (N_7022,N_4078,N_3421);
xor U7023 (N_7023,N_3264,N_5634);
nor U7024 (N_7024,N_4452,N_5256);
nand U7025 (N_7025,N_5297,N_5707);
or U7026 (N_7026,N_3366,N_4349);
nor U7027 (N_7027,N_4385,N_4539);
nand U7028 (N_7028,N_3796,N_5105);
nor U7029 (N_7029,N_3653,N_4918);
nor U7030 (N_7030,N_5168,N_4527);
nand U7031 (N_7031,N_4376,N_4065);
or U7032 (N_7032,N_5228,N_3029);
or U7033 (N_7033,N_4694,N_3566);
or U7034 (N_7034,N_5325,N_5127);
nand U7035 (N_7035,N_3370,N_4391);
nor U7036 (N_7036,N_4048,N_5920);
or U7037 (N_7037,N_3666,N_3410);
nand U7038 (N_7038,N_4869,N_3472);
xnor U7039 (N_7039,N_5548,N_3895);
xor U7040 (N_7040,N_3897,N_3438);
or U7041 (N_7041,N_5850,N_5159);
nand U7042 (N_7042,N_5449,N_3228);
nor U7043 (N_7043,N_3218,N_4958);
and U7044 (N_7044,N_4738,N_3091);
xor U7045 (N_7045,N_4697,N_5453);
or U7046 (N_7046,N_4634,N_5805);
nor U7047 (N_7047,N_4233,N_4025);
xor U7048 (N_7048,N_5842,N_4711);
nand U7049 (N_7049,N_5399,N_5888);
nor U7050 (N_7050,N_5682,N_4909);
and U7051 (N_7051,N_3093,N_3828);
nand U7052 (N_7052,N_3351,N_5954);
xor U7053 (N_7053,N_4411,N_5373);
nand U7054 (N_7054,N_4240,N_4249);
nand U7055 (N_7055,N_5142,N_3862);
nand U7056 (N_7056,N_4489,N_3823);
or U7057 (N_7057,N_3772,N_5706);
nand U7058 (N_7058,N_5886,N_4492);
and U7059 (N_7059,N_3639,N_3581);
nand U7060 (N_7060,N_3102,N_5859);
xor U7061 (N_7061,N_5936,N_5359);
nand U7062 (N_7062,N_4225,N_3597);
and U7063 (N_7063,N_3346,N_5641);
xnor U7064 (N_7064,N_3774,N_3684);
xor U7065 (N_7065,N_4318,N_3234);
nand U7066 (N_7066,N_5027,N_5058);
and U7067 (N_7067,N_3076,N_3946);
or U7068 (N_7068,N_3791,N_5395);
or U7069 (N_7069,N_5922,N_4490);
nand U7070 (N_7070,N_3467,N_4967);
and U7071 (N_7071,N_4690,N_5902);
or U7072 (N_7072,N_3126,N_3278);
and U7073 (N_7073,N_5471,N_3984);
xnor U7074 (N_7074,N_5463,N_4963);
or U7075 (N_7075,N_4880,N_3502);
or U7076 (N_7076,N_4049,N_3576);
and U7077 (N_7077,N_4477,N_3282);
or U7078 (N_7078,N_3701,N_5790);
nand U7079 (N_7079,N_5415,N_4328);
xnor U7080 (N_7080,N_5764,N_3479);
nand U7081 (N_7081,N_3060,N_3206);
xnor U7082 (N_7082,N_4540,N_5722);
or U7083 (N_7083,N_3548,N_5854);
xnor U7084 (N_7084,N_3057,N_3492);
or U7085 (N_7085,N_3004,N_3976);
or U7086 (N_7086,N_4617,N_5979);
and U7087 (N_7087,N_5720,N_3596);
nor U7088 (N_7088,N_3898,N_4510);
nand U7089 (N_7089,N_5801,N_5054);
xor U7090 (N_7090,N_5292,N_5679);
nand U7091 (N_7091,N_3000,N_4822);
nor U7092 (N_7092,N_4716,N_3038);
nand U7093 (N_7093,N_4045,N_3036);
xnor U7094 (N_7094,N_4992,N_4482);
or U7095 (N_7095,N_5687,N_3155);
nor U7096 (N_7096,N_5618,N_4631);
or U7097 (N_7097,N_5107,N_3664);
nand U7098 (N_7098,N_4948,N_5532);
nor U7099 (N_7099,N_5394,N_3737);
and U7100 (N_7100,N_4840,N_4773);
or U7101 (N_7101,N_3311,N_3509);
nand U7102 (N_7102,N_4808,N_3768);
nand U7103 (N_7103,N_3673,N_4672);
nand U7104 (N_7104,N_4175,N_5750);
xor U7105 (N_7105,N_5426,N_5131);
and U7106 (N_7106,N_5254,N_5385);
and U7107 (N_7107,N_4579,N_4382);
or U7108 (N_7108,N_3350,N_5824);
or U7109 (N_7109,N_3405,N_5183);
or U7110 (N_7110,N_5929,N_4867);
nand U7111 (N_7111,N_5574,N_4829);
nand U7112 (N_7112,N_4304,N_4961);
and U7113 (N_7113,N_5290,N_4425);
nand U7114 (N_7114,N_4056,N_3628);
xnor U7115 (N_7115,N_3164,N_5077);
or U7116 (N_7116,N_5121,N_3773);
xor U7117 (N_7117,N_5257,N_5671);
and U7118 (N_7118,N_4011,N_4729);
or U7119 (N_7119,N_5425,N_3089);
nor U7120 (N_7120,N_3843,N_3183);
xnor U7121 (N_7121,N_3181,N_4108);
nor U7122 (N_7122,N_5375,N_4034);
and U7123 (N_7123,N_4295,N_4212);
nand U7124 (N_7124,N_5684,N_5976);
or U7125 (N_7125,N_3078,N_3671);
and U7126 (N_7126,N_5466,N_3434);
nor U7127 (N_7127,N_4100,N_3977);
nand U7128 (N_7128,N_3470,N_3989);
nor U7129 (N_7129,N_4778,N_4314);
nand U7130 (N_7130,N_3641,N_4350);
nor U7131 (N_7131,N_3300,N_5932);
xor U7132 (N_7132,N_4419,N_3810);
nor U7133 (N_7133,N_5167,N_4430);
and U7134 (N_7134,N_3780,N_5862);
and U7135 (N_7135,N_3572,N_4661);
xor U7136 (N_7136,N_3097,N_3887);
nand U7137 (N_7137,N_4133,N_3230);
and U7138 (N_7138,N_3121,N_3558);
or U7139 (N_7139,N_4726,N_5299);
nor U7140 (N_7140,N_4624,N_5465);
or U7141 (N_7141,N_4887,N_3880);
and U7142 (N_7142,N_3618,N_5149);
nor U7143 (N_7143,N_5007,N_4970);
and U7144 (N_7144,N_5908,N_4710);
and U7145 (N_7145,N_3445,N_5372);
and U7146 (N_7146,N_5968,N_4377);
or U7147 (N_7147,N_5784,N_3961);
and U7148 (N_7148,N_5838,N_5568);
xor U7149 (N_7149,N_4159,N_5171);
xnor U7150 (N_7150,N_4820,N_3090);
xor U7151 (N_7151,N_4265,N_5469);
xnor U7152 (N_7152,N_4294,N_5945);
xnor U7153 (N_7153,N_4650,N_5724);
or U7154 (N_7154,N_3069,N_3811);
nor U7155 (N_7155,N_5295,N_3441);
xor U7156 (N_7156,N_4135,N_3518);
and U7157 (N_7157,N_4327,N_5122);
or U7158 (N_7158,N_3991,N_4052);
xnor U7159 (N_7159,N_5434,N_5562);
nor U7160 (N_7160,N_4491,N_4941);
nand U7161 (N_7161,N_5745,N_3744);
nor U7162 (N_7162,N_4291,N_5674);
nor U7163 (N_7163,N_3545,N_5109);
nand U7164 (N_7164,N_5363,N_3531);
nand U7165 (N_7165,N_5124,N_4446);
xnor U7166 (N_7166,N_4455,N_3127);
nor U7167 (N_7167,N_3238,N_4520);
xnor U7168 (N_7168,N_3648,N_5162);
or U7169 (N_7169,N_3224,N_3199);
xnor U7170 (N_7170,N_3716,N_4879);
nor U7171 (N_7171,N_5592,N_5298);
nor U7172 (N_7172,N_4022,N_5994);
nand U7173 (N_7173,N_5974,N_5777);
xor U7174 (N_7174,N_5717,N_5667);
xnor U7175 (N_7175,N_3188,N_5147);
nand U7176 (N_7176,N_4883,N_3848);
nand U7177 (N_7177,N_3098,N_3609);
nor U7178 (N_7178,N_5894,N_3763);
or U7179 (N_7179,N_3683,N_3575);
and U7180 (N_7180,N_4281,N_3275);
and U7181 (N_7181,N_4585,N_3670);
nor U7182 (N_7182,N_5948,N_5970);
xnor U7183 (N_7183,N_5440,N_5032);
nor U7184 (N_7184,N_4167,N_3886);
xor U7185 (N_7185,N_4594,N_5378);
or U7186 (N_7186,N_5264,N_5871);
or U7187 (N_7187,N_3939,N_5744);
nor U7188 (N_7188,N_4013,N_5797);
nand U7189 (N_7189,N_3702,N_5213);
or U7190 (N_7190,N_4047,N_3905);
xnor U7191 (N_7191,N_3051,N_3293);
nand U7192 (N_7192,N_3310,N_3299);
xor U7193 (N_7193,N_5008,N_4856);
or U7194 (N_7194,N_5772,N_5279);
and U7195 (N_7195,N_3182,N_5346);
nand U7196 (N_7196,N_3727,N_4289);
xnor U7197 (N_7197,N_4574,N_5345);
or U7198 (N_7198,N_4639,N_4004);
xnor U7199 (N_7199,N_3551,N_4786);
and U7200 (N_7200,N_3085,N_4347);
nor U7201 (N_7201,N_4556,N_4258);
nand U7202 (N_7202,N_4686,N_3106);
and U7203 (N_7203,N_3296,N_4899);
nor U7204 (N_7204,N_3643,N_4977);
or U7205 (N_7205,N_3650,N_4653);
nor U7206 (N_7206,N_5233,N_3251);
or U7207 (N_7207,N_5486,N_4508);
and U7208 (N_7208,N_3381,N_4533);
and U7209 (N_7209,N_4348,N_4125);
nor U7210 (N_7210,N_4006,N_3222);
xnor U7211 (N_7211,N_4868,N_3623);
nor U7212 (N_7212,N_3419,N_4494);
nand U7213 (N_7213,N_3526,N_3726);
xor U7214 (N_7214,N_3307,N_4524);
xnor U7215 (N_7215,N_4640,N_4788);
xor U7216 (N_7216,N_5396,N_5308);
nor U7217 (N_7217,N_5786,N_5166);
xnor U7218 (N_7218,N_5633,N_5773);
xnor U7219 (N_7219,N_4039,N_4301);
xnor U7220 (N_7220,N_3520,N_5590);
nand U7221 (N_7221,N_5928,N_5898);
xor U7222 (N_7222,N_5556,N_4418);
xnor U7223 (N_7223,N_5998,N_5332);
and U7224 (N_7224,N_3990,N_5031);
xnor U7225 (N_7225,N_5314,N_4026);
nand U7226 (N_7226,N_3669,N_3325);
xor U7227 (N_7227,N_4914,N_5488);
or U7228 (N_7228,N_4523,N_3573);
nor U7229 (N_7229,N_5458,N_4785);
nor U7230 (N_7230,N_5245,N_5208);
and U7231 (N_7231,N_3504,N_3598);
xor U7232 (N_7232,N_3168,N_3994);
or U7233 (N_7233,N_4673,N_5581);
or U7234 (N_7234,N_4399,N_3229);
or U7235 (N_7235,N_3489,N_3689);
xor U7236 (N_7236,N_3243,N_5636);
or U7237 (N_7237,N_3778,N_5704);
or U7238 (N_7238,N_3068,N_4476);
xnor U7239 (N_7239,N_4772,N_3704);
nor U7240 (N_7240,N_5301,N_5676);
nand U7241 (N_7241,N_5240,N_3095);
nor U7242 (N_7242,N_3697,N_3718);
xnor U7243 (N_7243,N_5856,N_5629);
or U7244 (N_7244,N_3117,N_4919);
and U7245 (N_7245,N_5036,N_5275);
xor U7246 (N_7246,N_3539,N_5606);
nor U7247 (N_7247,N_4754,N_3256);
or U7248 (N_7248,N_3910,N_4513);
nand U7249 (N_7249,N_3847,N_5229);
or U7250 (N_7250,N_5499,N_4551);
nor U7251 (N_7251,N_4043,N_4143);
nor U7252 (N_7252,N_3139,N_3011);
xnor U7253 (N_7253,N_3982,N_3207);
nor U7254 (N_7254,N_5579,N_5138);
or U7255 (N_7255,N_5847,N_4503);
nand U7256 (N_7256,N_3272,N_4707);
or U7257 (N_7257,N_5504,N_5263);
xor U7258 (N_7258,N_4209,N_5557);
or U7259 (N_7259,N_3599,N_4187);
xor U7260 (N_7260,N_5361,N_5989);
or U7261 (N_7261,N_4842,N_3302);
and U7262 (N_7262,N_3237,N_4926);
nor U7263 (N_7263,N_3462,N_3088);
or U7264 (N_7264,N_5282,N_5553);
nor U7265 (N_7265,N_5578,N_5958);
or U7266 (N_7266,N_3752,N_3245);
or U7267 (N_7267,N_4472,N_3603);
xor U7268 (N_7268,N_3284,N_4802);
nand U7269 (N_7269,N_4526,N_4106);
or U7270 (N_7270,N_4609,N_3014);
nor U7271 (N_7271,N_4370,N_3874);
xor U7272 (N_7272,N_3007,N_3116);
or U7273 (N_7273,N_4850,N_5155);
and U7274 (N_7274,N_3003,N_4285);
or U7275 (N_7275,N_3291,N_3568);
xor U7276 (N_7276,N_5566,N_3220);
xnor U7277 (N_7277,N_3714,N_4464);
and U7278 (N_7278,N_5369,N_4811);
or U7279 (N_7279,N_4163,N_5880);
xnor U7280 (N_7280,N_4649,N_3525);
nand U7281 (N_7281,N_3249,N_4445);
nand U7282 (N_7282,N_4516,N_3125);
and U7283 (N_7283,N_3070,N_5542);
nand U7284 (N_7284,N_4863,N_5646);
nand U7285 (N_7285,N_3316,N_5559);
nand U7286 (N_7286,N_5533,N_5879);
xor U7287 (N_7287,N_3172,N_4642);
nand U7288 (N_7288,N_4700,N_3170);
nor U7289 (N_7289,N_5529,N_4343);
nand U7290 (N_7290,N_3956,N_5713);
nor U7291 (N_7291,N_4150,N_3952);
and U7292 (N_7292,N_5398,N_3285);
nor U7293 (N_7293,N_5367,N_3620);
xor U7294 (N_7294,N_4791,N_3657);
nand U7295 (N_7295,N_4500,N_3375);
nor U7296 (N_7296,N_3308,N_4960);
or U7297 (N_7297,N_3373,N_5170);
nor U7298 (N_7298,N_3711,N_4239);
or U7299 (N_7299,N_5960,N_3625);
xnor U7300 (N_7300,N_4054,N_4473);
and U7301 (N_7301,N_3108,N_4266);
xor U7302 (N_7302,N_4423,N_3442);
xnor U7303 (N_7303,N_3784,N_5180);
nor U7304 (N_7304,N_3782,N_4408);
nor U7305 (N_7305,N_4927,N_5384);
nor U7306 (N_7306,N_3414,N_4231);
nand U7307 (N_7307,N_5672,N_5475);
or U7308 (N_7308,N_3873,N_3584);
nor U7309 (N_7309,N_3800,N_3771);
or U7310 (N_7310,N_4127,N_5270);
nand U7311 (N_7311,N_4932,N_3652);
nor U7312 (N_7312,N_5851,N_5376);
or U7313 (N_7313,N_3745,N_4203);
nand U7314 (N_7314,N_5787,N_3487);
and U7315 (N_7315,N_3179,N_3949);
xor U7316 (N_7316,N_5400,N_4950);
nor U7317 (N_7317,N_4444,N_5891);
nor U7318 (N_7318,N_4066,N_5779);
nand U7319 (N_7319,N_5262,N_5150);
and U7320 (N_7320,N_4973,N_5752);
xnor U7321 (N_7321,N_4226,N_3846);
xor U7322 (N_7322,N_4079,N_3236);
nand U7323 (N_7323,N_5655,N_5060);
nor U7324 (N_7324,N_5531,N_3587);
nand U7325 (N_7325,N_3913,N_3735);
xor U7326 (N_7326,N_5916,N_3929);
and U7327 (N_7327,N_5085,N_3411);
xor U7328 (N_7328,N_4913,N_4174);
or U7329 (N_7329,N_3382,N_5694);
and U7330 (N_7330,N_4283,N_4561);
nand U7331 (N_7331,N_3186,N_3101);
and U7332 (N_7332,N_4324,N_4504);
and U7333 (N_7333,N_5099,N_5586);
nor U7334 (N_7334,N_5442,N_5736);
or U7335 (N_7335,N_5068,N_4112);
xor U7336 (N_7336,N_5576,N_3024);
or U7337 (N_7337,N_4460,N_4572);
nor U7338 (N_7338,N_3824,N_5944);
nor U7339 (N_7339,N_4344,N_3047);
xnor U7340 (N_7340,N_3084,N_5209);
xnor U7341 (N_7341,N_5890,N_3214);
or U7342 (N_7342,N_3734,N_5635);
nor U7343 (N_7343,N_4942,N_3343);
or U7344 (N_7344,N_3606,N_4375);
xnor U7345 (N_7345,N_5490,N_3074);
nor U7346 (N_7346,N_3140,N_4063);
xnor U7347 (N_7347,N_3271,N_4248);
or U7348 (N_7348,N_5276,N_4208);
xor U7349 (N_7349,N_5860,N_5468);
nand U7350 (N_7350,N_3615,N_5337);
nor U7351 (N_7351,N_5802,N_5549);
nand U7352 (N_7352,N_4119,N_3775);
nor U7353 (N_7353,N_5591,N_5742);
nor U7354 (N_7354,N_4111,N_5443);
nor U7355 (N_7355,N_4548,N_3213);
nand U7356 (N_7356,N_5925,N_5323);
and U7357 (N_7357,N_5498,N_4659);
nand U7358 (N_7358,N_4660,N_4180);
nor U7359 (N_7359,N_4627,N_5519);
and U7360 (N_7360,N_3385,N_4176);
and U7361 (N_7361,N_3833,N_3988);
and U7362 (N_7362,N_3318,N_4873);
xnor U7363 (N_7363,N_5481,N_3053);
and U7364 (N_7364,N_3589,N_3921);
xor U7365 (N_7365,N_3622,N_5309);
nor U7366 (N_7366,N_3192,N_5855);
nand U7367 (N_7367,N_5525,N_4415);
nor U7368 (N_7368,N_5424,N_5609);
nand U7369 (N_7369,N_4059,N_4221);
nand U7370 (N_7370,N_4155,N_5265);
or U7371 (N_7371,N_3471,N_5867);
or U7372 (N_7372,N_5541,N_3210);
and U7373 (N_7373,N_4352,N_3486);
or U7374 (N_7374,N_4733,N_4297);
nor U7375 (N_7375,N_5780,N_3450);
xnor U7376 (N_7376,N_4924,N_3892);
nand U7377 (N_7377,N_3841,N_4018);
or U7378 (N_7378,N_5962,N_3527);
nor U7379 (N_7379,N_4215,N_3709);
or U7380 (N_7380,N_5913,N_5010);
xnor U7381 (N_7381,N_3693,N_4843);
nand U7382 (N_7382,N_3908,N_3339);
or U7383 (N_7383,N_3423,N_5158);
or U7384 (N_7384,N_4337,N_3159);
and U7385 (N_7385,N_5002,N_4403);
nand U7386 (N_7386,N_3396,N_4475);
and U7387 (N_7387,N_5716,N_5024);
nor U7388 (N_7388,N_3247,N_3447);
or U7389 (N_7389,N_5428,N_3415);
nand U7390 (N_7390,N_3377,N_5814);
nand U7391 (N_7391,N_3532,N_5386);
and U7392 (N_7392,N_4801,N_3219);
nor U7393 (N_7393,N_5050,N_5177);
nor U7394 (N_7394,N_4558,N_4756);
xnor U7395 (N_7395,N_3528,N_4535);
nor U7396 (N_7396,N_3052,N_3288);
or U7397 (N_7397,N_4904,N_5379);
or U7398 (N_7398,N_3161,N_3561);
or U7399 (N_7399,N_5762,N_4712);
xor U7400 (N_7400,N_5582,N_5708);
nor U7401 (N_7401,N_5161,N_3312);
or U7402 (N_7402,N_5620,N_5015);
and U7403 (N_7403,N_4849,N_4356);
xor U7404 (N_7404,N_5119,N_5630);
nand U7405 (N_7405,N_4901,N_3633);
or U7406 (N_7406,N_4373,N_3072);
and U7407 (N_7407,N_3677,N_4238);
or U7408 (N_7408,N_3100,N_4374);
or U7409 (N_7409,N_4814,N_4949);
and U7410 (N_7410,N_5755,N_5154);
nor U7411 (N_7411,N_4190,N_5037);
or U7412 (N_7412,N_5561,N_3703);
xor U7413 (N_7413,N_3048,N_5448);
nand U7414 (N_7414,N_5611,N_3455);
or U7415 (N_7415,N_5212,N_3482);
xor U7416 (N_7416,N_5621,N_3147);
xor U7417 (N_7417,N_5953,N_3872);
or U7418 (N_7418,N_4570,N_4483);
and U7419 (N_7419,N_4606,N_4121);
nand U7420 (N_7420,N_5028,N_4703);
nor U7421 (N_7421,N_3993,N_3785);
or U7422 (N_7422,N_5927,N_4717);
xnor U7423 (N_7423,N_5358,N_3132);
xnor U7424 (N_7424,N_4581,N_4273);
or U7425 (N_7425,N_4714,N_5409);
or U7426 (N_7426,N_3077,N_3969);
xor U7427 (N_7427,N_4319,N_3555);
nand U7428 (N_7428,N_4989,N_5729);
nand U7429 (N_7429,N_5637,N_3388);
and U7430 (N_7430,N_4287,N_4316);
nand U7431 (N_7431,N_4488,N_4214);
xor U7432 (N_7432,N_3607,N_5623);
or U7433 (N_7433,N_4875,N_3391);
nor U7434 (N_7434,N_5011,N_5422);
xor U7435 (N_7435,N_5446,N_4076);
xnor U7436 (N_7436,N_5333,N_3712);
xnor U7437 (N_7437,N_5402,N_4968);
or U7438 (N_7438,N_3225,N_4903);
xnor U7439 (N_7439,N_5306,N_5342);
nand U7440 (N_7440,N_5380,N_4068);
nand U7441 (N_7441,N_5751,N_4757);
and U7442 (N_7442,N_3485,N_5202);
nor U7443 (N_7443,N_5450,N_5901);
or U7444 (N_7444,N_4657,N_3212);
nor U7445 (N_7445,N_4422,N_5404);
xnor U7446 (N_7446,N_5798,N_4339);
xnor U7447 (N_7447,N_3710,N_4274);
and U7448 (N_7448,N_4454,N_5971);
and U7449 (N_7449,N_4769,N_3254);
xor U7450 (N_7450,N_3888,N_5320);
xnor U7451 (N_7451,N_5315,N_3099);
nor U7452 (N_7452,N_3536,N_3277);
xnor U7453 (N_7453,N_4552,N_4093);
xnor U7454 (N_7454,N_4972,N_5331);
or U7455 (N_7455,N_3005,N_4114);
nor U7456 (N_7456,N_5665,N_3861);
nand U7457 (N_7457,N_4041,N_3355);
nand U7458 (N_7458,N_3759,N_3336);
or U7459 (N_7459,N_4380,N_3305);
nand U7460 (N_7460,N_4622,N_5702);
or U7461 (N_7461,N_3337,N_5675);
nand U7462 (N_7462,N_5260,N_5628);
and U7463 (N_7463,N_4954,N_4865);
and U7464 (N_7464,N_4182,N_4196);
nor U7465 (N_7465,N_3553,N_3832);
xnor U7466 (N_7466,N_3205,N_3642);
or U7467 (N_7467,N_3835,N_4567);
or U7468 (N_7468,N_4161,N_4679);
or U7469 (N_7469,N_5113,N_4900);
nor U7470 (N_7470,N_5153,N_3250);
xnor U7471 (N_7471,N_4341,N_4171);
nor U7472 (N_7472,N_4771,N_4051);
nand U7473 (N_7473,N_4816,N_5961);
and U7474 (N_7474,N_4817,N_3844);
nor U7475 (N_7475,N_4202,N_5759);
xor U7476 (N_7476,N_3765,N_3200);
or U7477 (N_7477,N_4787,N_4652);
nand U7478 (N_7478,N_4429,N_4414);
nor U7479 (N_7479,N_3696,N_3513);
nand U7480 (N_7480,N_4797,N_3075);
nand U7481 (N_7481,N_5231,N_5478);
nor U7482 (N_7482,N_3280,N_3604);
nor U7483 (N_7483,N_4481,N_5996);
and U7484 (N_7484,N_3345,N_5567);
xnor U7485 (N_7485,N_5848,N_4604);
xnor U7486 (N_7486,N_5741,N_4207);
or U7487 (N_7487,N_4008,N_3197);
xor U7488 (N_7488,N_5539,N_4062);
and U7489 (N_7489,N_5021,N_4512);
or U7490 (N_7490,N_3239,N_3037);
xnor U7491 (N_7491,N_4897,N_3854);
nor U7492 (N_7492,N_3987,N_4562);
nand U7493 (N_7493,N_4704,N_4955);
xor U7494 (N_7494,N_3761,N_3510);
xnor U7495 (N_7495,N_5660,N_3235);
nand U7496 (N_7496,N_5420,N_3317);
xnor U7497 (N_7497,N_3968,N_3980);
or U7498 (N_7498,N_4894,N_4841);
and U7499 (N_7499,N_3966,N_3827);
nor U7500 (N_7500,N_5134,N_5656);
or U7501 (N_7501,N_5527,N_5043);
and U7502 (N_7502,N_5008,N_5276);
and U7503 (N_7503,N_5841,N_4149);
nand U7504 (N_7504,N_5959,N_4411);
nand U7505 (N_7505,N_5340,N_4382);
or U7506 (N_7506,N_5123,N_4747);
and U7507 (N_7507,N_4899,N_4095);
nor U7508 (N_7508,N_4716,N_3161);
xor U7509 (N_7509,N_4294,N_5697);
and U7510 (N_7510,N_4620,N_3840);
nor U7511 (N_7511,N_3928,N_3224);
nand U7512 (N_7512,N_3100,N_5433);
xor U7513 (N_7513,N_5635,N_5585);
or U7514 (N_7514,N_3834,N_4678);
nor U7515 (N_7515,N_3027,N_4358);
xor U7516 (N_7516,N_5607,N_4992);
xnor U7517 (N_7517,N_3961,N_4699);
and U7518 (N_7518,N_4103,N_5060);
xnor U7519 (N_7519,N_4119,N_5234);
and U7520 (N_7520,N_5740,N_4962);
and U7521 (N_7521,N_3035,N_5722);
xor U7522 (N_7522,N_4670,N_3780);
nor U7523 (N_7523,N_4698,N_3787);
xnor U7524 (N_7524,N_5074,N_3451);
xor U7525 (N_7525,N_3149,N_3327);
nand U7526 (N_7526,N_3369,N_3687);
nor U7527 (N_7527,N_5772,N_3802);
or U7528 (N_7528,N_3149,N_5832);
xnor U7529 (N_7529,N_3950,N_5159);
nor U7530 (N_7530,N_5163,N_3663);
nand U7531 (N_7531,N_3552,N_5627);
or U7532 (N_7532,N_5441,N_4879);
and U7533 (N_7533,N_4722,N_5038);
or U7534 (N_7534,N_3717,N_4136);
and U7535 (N_7535,N_5101,N_5359);
nor U7536 (N_7536,N_5591,N_3023);
or U7537 (N_7537,N_3387,N_3182);
and U7538 (N_7538,N_3850,N_5027);
nor U7539 (N_7539,N_4920,N_4152);
nor U7540 (N_7540,N_5023,N_5950);
nor U7541 (N_7541,N_3279,N_3517);
nor U7542 (N_7542,N_5261,N_3496);
xnor U7543 (N_7543,N_5340,N_3223);
nor U7544 (N_7544,N_5984,N_5220);
nand U7545 (N_7545,N_4750,N_3374);
or U7546 (N_7546,N_4121,N_3181);
nand U7547 (N_7547,N_4830,N_4432);
and U7548 (N_7548,N_3479,N_4845);
and U7549 (N_7549,N_4900,N_5040);
nor U7550 (N_7550,N_5054,N_4521);
nand U7551 (N_7551,N_3281,N_4996);
xor U7552 (N_7552,N_5953,N_5934);
or U7553 (N_7553,N_5479,N_4935);
xnor U7554 (N_7554,N_3454,N_3516);
nand U7555 (N_7555,N_5466,N_4809);
nor U7556 (N_7556,N_4112,N_4477);
and U7557 (N_7557,N_5003,N_3295);
or U7558 (N_7558,N_3255,N_4362);
nand U7559 (N_7559,N_3554,N_3082);
and U7560 (N_7560,N_4278,N_4848);
or U7561 (N_7561,N_3526,N_4458);
and U7562 (N_7562,N_5265,N_5341);
xnor U7563 (N_7563,N_5533,N_5320);
xnor U7564 (N_7564,N_3986,N_3944);
and U7565 (N_7565,N_4997,N_5213);
and U7566 (N_7566,N_3484,N_3962);
and U7567 (N_7567,N_3962,N_5641);
and U7568 (N_7568,N_3352,N_5582);
or U7569 (N_7569,N_5283,N_4704);
and U7570 (N_7570,N_3321,N_5969);
and U7571 (N_7571,N_4078,N_5608);
or U7572 (N_7572,N_5449,N_5540);
and U7573 (N_7573,N_5845,N_3354);
and U7574 (N_7574,N_4453,N_4810);
nand U7575 (N_7575,N_3494,N_3224);
nand U7576 (N_7576,N_3742,N_3167);
nand U7577 (N_7577,N_4036,N_3611);
nand U7578 (N_7578,N_4505,N_4384);
or U7579 (N_7579,N_5031,N_4530);
nand U7580 (N_7580,N_4844,N_3671);
xor U7581 (N_7581,N_4556,N_3416);
nand U7582 (N_7582,N_3175,N_3752);
nor U7583 (N_7583,N_4205,N_3555);
xor U7584 (N_7584,N_4938,N_4253);
xor U7585 (N_7585,N_4578,N_3687);
xor U7586 (N_7586,N_5619,N_3315);
nor U7587 (N_7587,N_3922,N_5152);
nor U7588 (N_7588,N_4536,N_4339);
or U7589 (N_7589,N_4853,N_5493);
or U7590 (N_7590,N_5663,N_5135);
and U7591 (N_7591,N_4391,N_5643);
or U7592 (N_7592,N_4707,N_3102);
and U7593 (N_7593,N_4093,N_4683);
and U7594 (N_7594,N_4287,N_3248);
nor U7595 (N_7595,N_4690,N_3776);
nand U7596 (N_7596,N_3248,N_4976);
xnor U7597 (N_7597,N_5761,N_3853);
and U7598 (N_7598,N_3259,N_4563);
and U7599 (N_7599,N_5439,N_5590);
nand U7600 (N_7600,N_3573,N_5055);
and U7601 (N_7601,N_3059,N_4029);
nor U7602 (N_7602,N_5127,N_5467);
nand U7603 (N_7603,N_3282,N_5926);
xnor U7604 (N_7604,N_4512,N_4356);
nand U7605 (N_7605,N_3182,N_5753);
or U7606 (N_7606,N_3042,N_4018);
nand U7607 (N_7607,N_4246,N_3397);
or U7608 (N_7608,N_5410,N_5536);
nand U7609 (N_7609,N_4403,N_3058);
xor U7610 (N_7610,N_3429,N_4121);
xor U7611 (N_7611,N_4494,N_3867);
and U7612 (N_7612,N_4745,N_3769);
nand U7613 (N_7613,N_3774,N_3866);
nor U7614 (N_7614,N_3612,N_5144);
or U7615 (N_7615,N_4122,N_4523);
xnor U7616 (N_7616,N_4064,N_5305);
nor U7617 (N_7617,N_4798,N_5996);
xnor U7618 (N_7618,N_5758,N_5906);
nor U7619 (N_7619,N_3847,N_4108);
xor U7620 (N_7620,N_3327,N_5988);
and U7621 (N_7621,N_3245,N_4662);
xnor U7622 (N_7622,N_5587,N_4584);
nand U7623 (N_7623,N_5245,N_5770);
xnor U7624 (N_7624,N_5251,N_5013);
and U7625 (N_7625,N_4157,N_5444);
xnor U7626 (N_7626,N_5378,N_3923);
nand U7627 (N_7627,N_3089,N_4474);
or U7628 (N_7628,N_5183,N_4705);
or U7629 (N_7629,N_3053,N_3112);
nor U7630 (N_7630,N_3296,N_4973);
or U7631 (N_7631,N_4884,N_3270);
nand U7632 (N_7632,N_3227,N_5521);
nand U7633 (N_7633,N_5766,N_3108);
nand U7634 (N_7634,N_3922,N_4644);
nand U7635 (N_7635,N_5431,N_5553);
xor U7636 (N_7636,N_3274,N_4791);
nand U7637 (N_7637,N_4675,N_3317);
nand U7638 (N_7638,N_3051,N_4095);
and U7639 (N_7639,N_5017,N_5071);
or U7640 (N_7640,N_3329,N_5122);
nand U7641 (N_7641,N_5380,N_4825);
nor U7642 (N_7642,N_4663,N_3889);
nor U7643 (N_7643,N_5909,N_4602);
nand U7644 (N_7644,N_5639,N_4233);
and U7645 (N_7645,N_4808,N_5957);
nor U7646 (N_7646,N_4348,N_5121);
and U7647 (N_7647,N_3829,N_3159);
or U7648 (N_7648,N_5674,N_4460);
nand U7649 (N_7649,N_3352,N_4980);
nand U7650 (N_7650,N_4480,N_3084);
nor U7651 (N_7651,N_5163,N_5048);
and U7652 (N_7652,N_5145,N_5123);
and U7653 (N_7653,N_3019,N_4806);
nor U7654 (N_7654,N_3236,N_4869);
nor U7655 (N_7655,N_3555,N_5395);
or U7656 (N_7656,N_4089,N_4024);
or U7657 (N_7657,N_3301,N_3703);
xor U7658 (N_7658,N_3099,N_5938);
nor U7659 (N_7659,N_3632,N_3126);
nand U7660 (N_7660,N_3682,N_3943);
and U7661 (N_7661,N_5769,N_3415);
and U7662 (N_7662,N_3005,N_4735);
and U7663 (N_7663,N_5332,N_3226);
nand U7664 (N_7664,N_5594,N_4752);
or U7665 (N_7665,N_4361,N_3861);
or U7666 (N_7666,N_5183,N_5710);
or U7667 (N_7667,N_5590,N_4064);
xor U7668 (N_7668,N_3938,N_4939);
nor U7669 (N_7669,N_4541,N_4186);
nor U7670 (N_7670,N_3609,N_5487);
and U7671 (N_7671,N_5111,N_4912);
xnor U7672 (N_7672,N_3328,N_4294);
or U7673 (N_7673,N_5964,N_4417);
nand U7674 (N_7674,N_5399,N_5439);
xor U7675 (N_7675,N_3244,N_5875);
xnor U7676 (N_7676,N_3277,N_4678);
or U7677 (N_7677,N_5502,N_4011);
and U7678 (N_7678,N_4878,N_4549);
xor U7679 (N_7679,N_5197,N_4296);
or U7680 (N_7680,N_4376,N_3743);
xnor U7681 (N_7681,N_4387,N_5070);
nand U7682 (N_7682,N_5902,N_4280);
and U7683 (N_7683,N_3013,N_5153);
nor U7684 (N_7684,N_5955,N_5247);
and U7685 (N_7685,N_3342,N_4294);
xnor U7686 (N_7686,N_4092,N_3998);
xor U7687 (N_7687,N_4750,N_3892);
nor U7688 (N_7688,N_5483,N_5149);
xor U7689 (N_7689,N_5279,N_5351);
or U7690 (N_7690,N_5948,N_3754);
or U7691 (N_7691,N_3742,N_3816);
nand U7692 (N_7692,N_5945,N_3892);
and U7693 (N_7693,N_3348,N_4918);
nor U7694 (N_7694,N_3950,N_3654);
or U7695 (N_7695,N_4651,N_5418);
nand U7696 (N_7696,N_4060,N_3139);
xnor U7697 (N_7697,N_5092,N_4800);
or U7698 (N_7698,N_5403,N_3182);
nand U7699 (N_7699,N_3775,N_5269);
nand U7700 (N_7700,N_5188,N_5698);
xor U7701 (N_7701,N_3277,N_4510);
and U7702 (N_7702,N_4432,N_3382);
nor U7703 (N_7703,N_3497,N_3830);
or U7704 (N_7704,N_4901,N_4379);
nor U7705 (N_7705,N_3434,N_3191);
nor U7706 (N_7706,N_4581,N_5787);
or U7707 (N_7707,N_4842,N_4878);
nand U7708 (N_7708,N_5875,N_4224);
or U7709 (N_7709,N_4311,N_5166);
and U7710 (N_7710,N_3427,N_4714);
nor U7711 (N_7711,N_3710,N_5517);
or U7712 (N_7712,N_3403,N_5256);
xnor U7713 (N_7713,N_5327,N_3423);
nor U7714 (N_7714,N_3450,N_3209);
or U7715 (N_7715,N_5343,N_3790);
nor U7716 (N_7716,N_4628,N_3487);
or U7717 (N_7717,N_4916,N_4887);
or U7718 (N_7718,N_4609,N_5581);
nand U7719 (N_7719,N_3836,N_3547);
nand U7720 (N_7720,N_5949,N_5529);
or U7721 (N_7721,N_5641,N_5833);
or U7722 (N_7722,N_5034,N_4404);
and U7723 (N_7723,N_5613,N_3287);
and U7724 (N_7724,N_5543,N_5961);
nand U7725 (N_7725,N_5401,N_3277);
and U7726 (N_7726,N_4868,N_4648);
nand U7727 (N_7727,N_5439,N_3565);
and U7728 (N_7728,N_5291,N_4839);
or U7729 (N_7729,N_5647,N_5462);
nand U7730 (N_7730,N_3474,N_4338);
and U7731 (N_7731,N_4651,N_3620);
and U7732 (N_7732,N_3911,N_4730);
nor U7733 (N_7733,N_4988,N_4429);
nand U7734 (N_7734,N_4704,N_5268);
nand U7735 (N_7735,N_4008,N_3553);
nor U7736 (N_7736,N_3474,N_3157);
and U7737 (N_7737,N_4464,N_3257);
or U7738 (N_7738,N_3599,N_5431);
nand U7739 (N_7739,N_3438,N_5885);
or U7740 (N_7740,N_4457,N_5630);
or U7741 (N_7741,N_3812,N_5198);
nand U7742 (N_7742,N_5912,N_3012);
and U7743 (N_7743,N_5381,N_4925);
or U7744 (N_7744,N_4381,N_3872);
or U7745 (N_7745,N_3505,N_4750);
and U7746 (N_7746,N_4731,N_4750);
and U7747 (N_7747,N_4396,N_3282);
nand U7748 (N_7748,N_3110,N_5156);
and U7749 (N_7749,N_4685,N_5285);
xor U7750 (N_7750,N_3360,N_4173);
and U7751 (N_7751,N_5298,N_4947);
and U7752 (N_7752,N_3198,N_4256);
or U7753 (N_7753,N_5958,N_5767);
and U7754 (N_7754,N_4346,N_5761);
nor U7755 (N_7755,N_4790,N_5496);
or U7756 (N_7756,N_4764,N_5776);
xnor U7757 (N_7757,N_3538,N_3729);
and U7758 (N_7758,N_5230,N_4837);
and U7759 (N_7759,N_5374,N_4398);
or U7760 (N_7760,N_5919,N_4212);
nor U7761 (N_7761,N_4107,N_4149);
and U7762 (N_7762,N_4379,N_3276);
or U7763 (N_7763,N_4212,N_3352);
nor U7764 (N_7764,N_4797,N_3597);
nor U7765 (N_7765,N_4904,N_3775);
xor U7766 (N_7766,N_3965,N_3199);
xor U7767 (N_7767,N_4521,N_5313);
nor U7768 (N_7768,N_5483,N_3699);
xnor U7769 (N_7769,N_5287,N_3376);
nor U7770 (N_7770,N_5151,N_4174);
nor U7771 (N_7771,N_3906,N_5344);
nand U7772 (N_7772,N_3207,N_3505);
or U7773 (N_7773,N_3189,N_3566);
xnor U7774 (N_7774,N_5879,N_4922);
xor U7775 (N_7775,N_4827,N_3227);
and U7776 (N_7776,N_4808,N_3990);
and U7777 (N_7777,N_5803,N_5743);
nor U7778 (N_7778,N_4660,N_5574);
or U7779 (N_7779,N_5581,N_5099);
nand U7780 (N_7780,N_5852,N_5907);
xor U7781 (N_7781,N_5461,N_5189);
nand U7782 (N_7782,N_5410,N_3711);
or U7783 (N_7783,N_3129,N_4787);
nor U7784 (N_7784,N_4071,N_3778);
and U7785 (N_7785,N_3798,N_3367);
and U7786 (N_7786,N_5776,N_3144);
or U7787 (N_7787,N_3150,N_3006);
nor U7788 (N_7788,N_3618,N_4014);
nand U7789 (N_7789,N_5331,N_3896);
xor U7790 (N_7790,N_4766,N_4487);
xor U7791 (N_7791,N_5962,N_4999);
and U7792 (N_7792,N_5228,N_5655);
and U7793 (N_7793,N_4914,N_5876);
and U7794 (N_7794,N_3132,N_3736);
and U7795 (N_7795,N_4032,N_5559);
nand U7796 (N_7796,N_4725,N_4120);
and U7797 (N_7797,N_4652,N_4934);
or U7798 (N_7798,N_3358,N_4945);
nand U7799 (N_7799,N_5187,N_4641);
nand U7800 (N_7800,N_3947,N_5142);
or U7801 (N_7801,N_3827,N_4193);
xor U7802 (N_7802,N_4261,N_4433);
xor U7803 (N_7803,N_5410,N_5681);
or U7804 (N_7804,N_3748,N_4274);
or U7805 (N_7805,N_4517,N_4996);
and U7806 (N_7806,N_5761,N_4866);
nand U7807 (N_7807,N_3234,N_4825);
nor U7808 (N_7808,N_3104,N_3483);
xnor U7809 (N_7809,N_5039,N_5825);
nand U7810 (N_7810,N_3442,N_4535);
or U7811 (N_7811,N_3765,N_4208);
nand U7812 (N_7812,N_4102,N_3922);
and U7813 (N_7813,N_5732,N_5680);
or U7814 (N_7814,N_4699,N_5656);
or U7815 (N_7815,N_5428,N_4387);
nor U7816 (N_7816,N_3758,N_4218);
or U7817 (N_7817,N_5271,N_4457);
nor U7818 (N_7818,N_3425,N_3306);
or U7819 (N_7819,N_5391,N_4157);
xnor U7820 (N_7820,N_4056,N_4671);
or U7821 (N_7821,N_4771,N_5417);
or U7822 (N_7822,N_3131,N_3156);
xnor U7823 (N_7823,N_4819,N_3700);
xor U7824 (N_7824,N_5490,N_4294);
or U7825 (N_7825,N_4572,N_4765);
or U7826 (N_7826,N_4679,N_3094);
and U7827 (N_7827,N_4244,N_4982);
nor U7828 (N_7828,N_3906,N_4614);
xnor U7829 (N_7829,N_5501,N_4715);
nand U7830 (N_7830,N_3064,N_5496);
nand U7831 (N_7831,N_5824,N_5356);
nor U7832 (N_7832,N_3909,N_3499);
xnor U7833 (N_7833,N_3456,N_3208);
nor U7834 (N_7834,N_4410,N_4902);
nor U7835 (N_7835,N_4746,N_4376);
xnor U7836 (N_7836,N_4269,N_3476);
xnor U7837 (N_7837,N_4547,N_4259);
nand U7838 (N_7838,N_5158,N_3350);
nand U7839 (N_7839,N_5987,N_3912);
and U7840 (N_7840,N_3861,N_3812);
and U7841 (N_7841,N_3465,N_4478);
and U7842 (N_7842,N_5252,N_4650);
and U7843 (N_7843,N_5554,N_3516);
nand U7844 (N_7844,N_3465,N_3712);
xor U7845 (N_7845,N_5494,N_5924);
and U7846 (N_7846,N_5314,N_3656);
and U7847 (N_7847,N_3564,N_5856);
or U7848 (N_7848,N_3862,N_5413);
nor U7849 (N_7849,N_5061,N_3026);
nand U7850 (N_7850,N_4267,N_4266);
or U7851 (N_7851,N_4132,N_4048);
and U7852 (N_7852,N_5296,N_4788);
and U7853 (N_7853,N_4489,N_4793);
nand U7854 (N_7854,N_5126,N_3435);
nor U7855 (N_7855,N_5848,N_3158);
and U7856 (N_7856,N_5276,N_5152);
nand U7857 (N_7857,N_4471,N_4542);
xnor U7858 (N_7858,N_5680,N_5647);
xnor U7859 (N_7859,N_5899,N_3671);
nor U7860 (N_7860,N_5848,N_3698);
and U7861 (N_7861,N_4394,N_5310);
xnor U7862 (N_7862,N_5252,N_4051);
xor U7863 (N_7863,N_4750,N_3700);
nor U7864 (N_7864,N_3173,N_3469);
xor U7865 (N_7865,N_4948,N_5505);
and U7866 (N_7866,N_3724,N_4087);
nor U7867 (N_7867,N_5254,N_5221);
or U7868 (N_7868,N_3168,N_3457);
and U7869 (N_7869,N_3518,N_5225);
nor U7870 (N_7870,N_3931,N_4647);
nor U7871 (N_7871,N_5262,N_4735);
xor U7872 (N_7872,N_4059,N_4623);
xnor U7873 (N_7873,N_4954,N_5985);
or U7874 (N_7874,N_5272,N_3303);
and U7875 (N_7875,N_5788,N_5207);
nor U7876 (N_7876,N_3656,N_5896);
nor U7877 (N_7877,N_5640,N_3664);
and U7878 (N_7878,N_5656,N_3578);
xor U7879 (N_7879,N_4688,N_3783);
or U7880 (N_7880,N_4222,N_3042);
or U7881 (N_7881,N_5234,N_3807);
nand U7882 (N_7882,N_5515,N_5852);
and U7883 (N_7883,N_5252,N_5761);
xor U7884 (N_7884,N_5440,N_5743);
xnor U7885 (N_7885,N_4091,N_4902);
xnor U7886 (N_7886,N_4859,N_5409);
nand U7887 (N_7887,N_5639,N_4343);
xnor U7888 (N_7888,N_4101,N_4357);
or U7889 (N_7889,N_4600,N_5189);
and U7890 (N_7890,N_3983,N_3280);
nor U7891 (N_7891,N_4933,N_5442);
nand U7892 (N_7892,N_4764,N_4250);
nor U7893 (N_7893,N_5104,N_3753);
nand U7894 (N_7894,N_5192,N_3041);
nand U7895 (N_7895,N_3228,N_4066);
nor U7896 (N_7896,N_4065,N_4994);
or U7897 (N_7897,N_5007,N_4400);
and U7898 (N_7898,N_5446,N_4168);
and U7899 (N_7899,N_3204,N_3946);
xnor U7900 (N_7900,N_4986,N_3459);
nand U7901 (N_7901,N_3289,N_4263);
or U7902 (N_7902,N_3856,N_5879);
and U7903 (N_7903,N_4822,N_4236);
nor U7904 (N_7904,N_4772,N_5827);
nor U7905 (N_7905,N_5779,N_4364);
nand U7906 (N_7906,N_4936,N_5193);
or U7907 (N_7907,N_4491,N_3207);
and U7908 (N_7908,N_3759,N_5786);
xnor U7909 (N_7909,N_4933,N_3010);
nand U7910 (N_7910,N_3792,N_3231);
nor U7911 (N_7911,N_3204,N_3346);
nor U7912 (N_7912,N_5231,N_3173);
nand U7913 (N_7913,N_4344,N_5765);
nor U7914 (N_7914,N_3642,N_3027);
xor U7915 (N_7915,N_5224,N_5086);
nand U7916 (N_7916,N_4140,N_4776);
xor U7917 (N_7917,N_3589,N_4147);
xnor U7918 (N_7918,N_5756,N_4566);
and U7919 (N_7919,N_5248,N_4658);
and U7920 (N_7920,N_5424,N_5017);
xnor U7921 (N_7921,N_3306,N_3083);
and U7922 (N_7922,N_4231,N_5615);
nand U7923 (N_7923,N_5652,N_5629);
nand U7924 (N_7924,N_3766,N_4523);
or U7925 (N_7925,N_5280,N_3640);
and U7926 (N_7926,N_3821,N_4439);
nor U7927 (N_7927,N_5511,N_5205);
or U7928 (N_7928,N_4325,N_3025);
and U7929 (N_7929,N_3609,N_5775);
or U7930 (N_7930,N_5521,N_4545);
or U7931 (N_7931,N_4964,N_5020);
or U7932 (N_7932,N_5152,N_3372);
xor U7933 (N_7933,N_5270,N_4392);
and U7934 (N_7934,N_3254,N_4946);
nand U7935 (N_7935,N_4256,N_4961);
or U7936 (N_7936,N_3090,N_3844);
nor U7937 (N_7937,N_3425,N_3057);
or U7938 (N_7938,N_3103,N_5113);
and U7939 (N_7939,N_3473,N_5321);
nor U7940 (N_7940,N_5374,N_5648);
xnor U7941 (N_7941,N_3345,N_4859);
xor U7942 (N_7942,N_3480,N_5061);
or U7943 (N_7943,N_3126,N_4945);
or U7944 (N_7944,N_3286,N_3243);
xnor U7945 (N_7945,N_3873,N_4286);
xor U7946 (N_7946,N_3673,N_3064);
xnor U7947 (N_7947,N_5976,N_5370);
and U7948 (N_7948,N_4454,N_4071);
or U7949 (N_7949,N_5067,N_4118);
and U7950 (N_7950,N_4954,N_5173);
xnor U7951 (N_7951,N_4217,N_5732);
nand U7952 (N_7952,N_3858,N_4422);
or U7953 (N_7953,N_5356,N_3753);
or U7954 (N_7954,N_3540,N_4331);
nor U7955 (N_7955,N_4617,N_4314);
xor U7956 (N_7956,N_5944,N_4449);
xnor U7957 (N_7957,N_4545,N_3296);
or U7958 (N_7958,N_5089,N_4704);
xnor U7959 (N_7959,N_3257,N_4066);
nand U7960 (N_7960,N_4134,N_4132);
nor U7961 (N_7961,N_3807,N_5784);
nor U7962 (N_7962,N_3062,N_3007);
and U7963 (N_7963,N_3678,N_4868);
and U7964 (N_7964,N_4579,N_4954);
nor U7965 (N_7965,N_3262,N_5338);
or U7966 (N_7966,N_3181,N_3368);
nand U7967 (N_7967,N_5632,N_4417);
or U7968 (N_7968,N_5849,N_4887);
and U7969 (N_7969,N_4023,N_5564);
or U7970 (N_7970,N_5572,N_4773);
xnor U7971 (N_7971,N_3021,N_4480);
and U7972 (N_7972,N_4234,N_4141);
or U7973 (N_7973,N_3869,N_5646);
xnor U7974 (N_7974,N_5169,N_3012);
xor U7975 (N_7975,N_5831,N_5414);
xor U7976 (N_7976,N_5832,N_3424);
nand U7977 (N_7977,N_3978,N_5217);
and U7978 (N_7978,N_3573,N_3196);
and U7979 (N_7979,N_5808,N_3770);
or U7980 (N_7980,N_3136,N_5356);
nor U7981 (N_7981,N_5261,N_5372);
xor U7982 (N_7982,N_3278,N_4874);
nor U7983 (N_7983,N_5232,N_3164);
and U7984 (N_7984,N_3422,N_3977);
nor U7985 (N_7985,N_3427,N_4214);
and U7986 (N_7986,N_5891,N_5147);
xor U7987 (N_7987,N_4995,N_3526);
and U7988 (N_7988,N_4113,N_5209);
xnor U7989 (N_7989,N_4853,N_3292);
nand U7990 (N_7990,N_3540,N_3794);
xor U7991 (N_7991,N_4933,N_5423);
and U7992 (N_7992,N_3684,N_5141);
and U7993 (N_7993,N_5818,N_5098);
and U7994 (N_7994,N_3606,N_3680);
or U7995 (N_7995,N_4164,N_3258);
nand U7996 (N_7996,N_4188,N_5245);
nor U7997 (N_7997,N_5514,N_3851);
nand U7998 (N_7998,N_5148,N_4640);
or U7999 (N_7999,N_5415,N_4465);
and U8000 (N_8000,N_5197,N_4171);
nor U8001 (N_8001,N_5617,N_5934);
nand U8002 (N_8002,N_4886,N_4503);
nand U8003 (N_8003,N_3472,N_5217);
or U8004 (N_8004,N_3895,N_3295);
xnor U8005 (N_8005,N_3500,N_5890);
nand U8006 (N_8006,N_4818,N_3704);
and U8007 (N_8007,N_5195,N_4506);
or U8008 (N_8008,N_4001,N_3502);
and U8009 (N_8009,N_3698,N_3934);
nor U8010 (N_8010,N_5177,N_3041);
nor U8011 (N_8011,N_5400,N_5462);
or U8012 (N_8012,N_4361,N_5697);
or U8013 (N_8013,N_4089,N_3797);
nand U8014 (N_8014,N_5296,N_5094);
or U8015 (N_8015,N_3565,N_5928);
nor U8016 (N_8016,N_4173,N_5485);
or U8017 (N_8017,N_4974,N_3078);
and U8018 (N_8018,N_5100,N_4183);
nor U8019 (N_8019,N_3783,N_5824);
and U8020 (N_8020,N_4545,N_5149);
or U8021 (N_8021,N_3521,N_4783);
xnor U8022 (N_8022,N_3557,N_3998);
xnor U8023 (N_8023,N_4365,N_3796);
xnor U8024 (N_8024,N_5331,N_3474);
nor U8025 (N_8025,N_4620,N_5557);
xor U8026 (N_8026,N_5836,N_5924);
xnor U8027 (N_8027,N_4044,N_5136);
and U8028 (N_8028,N_5965,N_5329);
and U8029 (N_8029,N_5963,N_3810);
nor U8030 (N_8030,N_5454,N_5155);
or U8031 (N_8031,N_3517,N_5471);
and U8032 (N_8032,N_3540,N_3272);
or U8033 (N_8033,N_3769,N_4540);
or U8034 (N_8034,N_4734,N_3658);
xnor U8035 (N_8035,N_3227,N_5276);
xnor U8036 (N_8036,N_3472,N_4921);
nor U8037 (N_8037,N_3585,N_3095);
nor U8038 (N_8038,N_4071,N_3880);
xor U8039 (N_8039,N_5775,N_4137);
and U8040 (N_8040,N_4558,N_3022);
nor U8041 (N_8041,N_4202,N_4457);
nand U8042 (N_8042,N_5206,N_4956);
xnor U8043 (N_8043,N_5033,N_4325);
xnor U8044 (N_8044,N_3625,N_5457);
xor U8045 (N_8045,N_3958,N_4901);
or U8046 (N_8046,N_4002,N_5118);
nand U8047 (N_8047,N_5000,N_3087);
and U8048 (N_8048,N_4654,N_5371);
or U8049 (N_8049,N_5260,N_4167);
nor U8050 (N_8050,N_4366,N_3355);
and U8051 (N_8051,N_3431,N_3642);
and U8052 (N_8052,N_5721,N_4288);
nand U8053 (N_8053,N_4018,N_5948);
or U8054 (N_8054,N_4315,N_4033);
nor U8055 (N_8055,N_5322,N_3673);
nor U8056 (N_8056,N_5512,N_5830);
and U8057 (N_8057,N_3090,N_3797);
nand U8058 (N_8058,N_5076,N_3864);
nand U8059 (N_8059,N_4557,N_3351);
xnor U8060 (N_8060,N_3802,N_3740);
or U8061 (N_8061,N_5699,N_5370);
and U8062 (N_8062,N_3454,N_3687);
nand U8063 (N_8063,N_4780,N_3322);
nand U8064 (N_8064,N_3964,N_5509);
or U8065 (N_8065,N_3121,N_4797);
nand U8066 (N_8066,N_3911,N_5814);
or U8067 (N_8067,N_3655,N_5648);
xnor U8068 (N_8068,N_3875,N_4460);
nand U8069 (N_8069,N_5090,N_5474);
nor U8070 (N_8070,N_5536,N_4438);
or U8071 (N_8071,N_3647,N_3217);
nand U8072 (N_8072,N_3042,N_3830);
xnor U8073 (N_8073,N_3542,N_3786);
nand U8074 (N_8074,N_3517,N_3199);
nor U8075 (N_8075,N_3602,N_5449);
and U8076 (N_8076,N_5016,N_3990);
or U8077 (N_8077,N_4427,N_5375);
and U8078 (N_8078,N_4083,N_4967);
or U8079 (N_8079,N_4329,N_5851);
or U8080 (N_8080,N_5280,N_3379);
or U8081 (N_8081,N_3211,N_4796);
and U8082 (N_8082,N_4614,N_4684);
nand U8083 (N_8083,N_5577,N_3704);
or U8084 (N_8084,N_4171,N_5928);
or U8085 (N_8085,N_3303,N_3343);
xnor U8086 (N_8086,N_4671,N_5372);
and U8087 (N_8087,N_5809,N_5380);
and U8088 (N_8088,N_4134,N_3549);
nor U8089 (N_8089,N_3107,N_4945);
xor U8090 (N_8090,N_4590,N_3695);
xnor U8091 (N_8091,N_3759,N_3259);
xor U8092 (N_8092,N_3087,N_3170);
nand U8093 (N_8093,N_4611,N_3015);
xor U8094 (N_8094,N_5514,N_4396);
nor U8095 (N_8095,N_4397,N_4272);
xnor U8096 (N_8096,N_4714,N_5687);
or U8097 (N_8097,N_3926,N_3686);
and U8098 (N_8098,N_3309,N_4401);
xor U8099 (N_8099,N_5609,N_5246);
and U8100 (N_8100,N_3193,N_5056);
nand U8101 (N_8101,N_4291,N_3192);
xor U8102 (N_8102,N_4127,N_3626);
nand U8103 (N_8103,N_5462,N_3184);
nand U8104 (N_8104,N_4023,N_4936);
or U8105 (N_8105,N_4219,N_5569);
and U8106 (N_8106,N_4884,N_3980);
nor U8107 (N_8107,N_4698,N_5851);
nand U8108 (N_8108,N_3682,N_4884);
or U8109 (N_8109,N_4661,N_4732);
nor U8110 (N_8110,N_5299,N_5726);
nor U8111 (N_8111,N_4189,N_3286);
nor U8112 (N_8112,N_3621,N_4830);
nand U8113 (N_8113,N_4595,N_3054);
nor U8114 (N_8114,N_3562,N_3073);
xor U8115 (N_8115,N_5617,N_5086);
xnor U8116 (N_8116,N_3564,N_4784);
nor U8117 (N_8117,N_5474,N_4281);
nor U8118 (N_8118,N_3460,N_5224);
or U8119 (N_8119,N_3628,N_3525);
xor U8120 (N_8120,N_4682,N_4523);
or U8121 (N_8121,N_4807,N_4553);
or U8122 (N_8122,N_4172,N_5751);
and U8123 (N_8123,N_4810,N_5132);
or U8124 (N_8124,N_5284,N_3890);
nand U8125 (N_8125,N_5835,N_5054);
or U8126 (N_8126,N_5569,N_4610);
nand U8127 (N_8127,N_5025,N_3214);
and U8128 (N_8128,N_4492,N_5981);
nor U8129 (N_8129,N_5790,N_4130);
xor U8130 (N_8130,N_5191,N_5373);
xor U8131 (N_8131,N_5606,N_4939);
nor U8132 (N_8132,N_3292,N_4686);
xor U8133 (N_8133,N_4440,N_3119);
xnor U8134 (N_8134,N_5666,N_4943);
and U8135 (N_8135,N_3465,N_5551);
or U8136 (N_8136,N_4318,N_4728);
xnor U8137 (N_8137,N_4670,N_3581);
nor U8138 (N_8138,N_5444,N_4465);
nand U8139 (N_8139,N_3843,N_5676);
xnor U8140 (N_8140,N_4705,N_5700);
xnor U8141 (N_8141,N_5849,N_3401);
and U8142 (N_8142,N_4708,N_3805);
and U8143 (N_8143,N_4708,N_4067);
and U8144 (N_8144,N_3953,N_5761);
nor U8145 (N_8145,N_3198,N_5785);
xor U8146 (N_8146,N_3139,N_5397);
xnor U8147 (N_8147,N_4082,N_4530);
nor U8148 (N_8148,N_4150,N_5657);
and U8149 (N_8149,N_3945,N_3668);
and U8150 (N_8150,N_3650,N_4523);
or U8151 (N_8151,N_3084,N_5322);
nand U8152 (N_8152,N_5800,N_3841);
nor U8153 (N_8153,N_3374,N_5010);
xor U8154 (N_8154,N_5758,N_3725);
nand U8155 (N_8155,N_3713,N_3066);
nor U8156 (N_8156,N_3807,N_5470);
and U8157 (N_8157,N_4723,N_5345);
and U8158 (N_8158,N_5691,N_5076);
xor U8159 (N_8159,N_5113,N_4462);
xor U8160 (N_8160,N_3128,N_4910);
or U8161 (N_8161,N_4237,N_3575);
nor U8162 (N_8162,N_3674,N_4588);
nand U8163 (N_8163,N_5250,N_5409);
nand U8164 (N_8164,N_3362,N_4586);
nand U8165 (N_8165,N_5404,N_5414);
nand U8166 (N_8166,N_4493,N_5274);
xor U8167 (N_8167,N_5597,N_5875);
nand U8168 (N_8168,N_4335,N_4296);
xnor U8169 (N_8169,N_3668,N_3564);
nor U8170 (N_8170,N_4854,N_4037);
and U8171 (N_8171,N_5550,N_3276);
nand U8172 (N_8172,N_3150,N_3648);
and U8173 (N_8173,N_4670,N_4912);
nand U8174 (N_8174,N_4448,N_5252);
nand U8175 (N_8175,N_3655,N_3375);
nand U8176 (N_8176,N_3090,N_4150);
xnor U8177 (N_8177,N_3793,N_4272);
and U8178 (N_8178,N_4606,N_4123);
xor U8179 (N_8179,N_5490,N_3695);
nand U8180 (N_8180,N_4217,N_4357);
xor U8181 (N_8181,N_4022,N_4850);
nand U8182 (N_8182,N_4073,N_5571);
nand U8183 (N_8183,N_4579,N_5309);
or U8184 (N_8184,N_3880,N_5577);
or U8185 (N_8185,N_3723,N_3284);
and U8186 (N_8186,N_3522,N_3837);
nand U8187 (N_8187,N_4617,N_3280);
xnor U8188 (N_8188,N_3231,N_5713);
and U8189 (N_8189,N_4293,N_4208);
nand U8190 (N_8190,N_5759,N_5569);
xor U8191 (N_8191,N_3141,N_3785);
and U8192 (N_8192,N_4392,N_4170);
and U8193 (N_8193,N_5811,N_3002);
xnor U8194 (N_8194,N_5889,N_5369);
xnor U8195 (N_8195,N_5387,N_4751);
xnor U8196 (N_8196,N_3888,N_4097);
xnor U8197 (N_8197,N_4040,N_4079);
and U8198 (N_8198,N_4365,N_3010);
xnor U8199 (N_8199,N_4232,N_4016);
nand U8200 (N_8200,N_3013,N_3114);
nor U8201 (N_8201,N_5626,N_4914);
xnor U8202 (N_8202,N_3311,N_4626);
nand U8203 (N_8203,N_3712,N_3806);
nand U8204 (N_8204,N_4566,N_3978);
or U8205 (N_8205,N_3615,N_4754);
xnor U8206 (N_8206,N_5894,N_5429);
xor U8207 (N_8207,N_5444,N_5120);
xnor U8208 (N_8208,N_3067,N_5117);
or U8209 (N_8209,N_5604,N_5050);
nand U8210 (N_8210,N_5166,N_4577);
nor U8211 (N_8211,N_3021,N_5491);
or U8212 (N_8212,N_3155,N_4764);
nand U8213 (N_8213,N_3652,N_5487);
or U8214 (N_8214,N_3091,N_3954);
or U8215 (N_8215,N_4930,N_3788);
xor U8216 (N_8216,N_3763,N_5313);
nor U8217 (N_8217,N_5761,N_3113);
nor U8218 (N_8218,N_5478,N_4284);
nand U8219 (N_8219,N_4463,N_3804);
and U8220 (N_8220,N_3435,N_5553);
or U8221 (N_8221,N_5584,N_3376);
xor U8222 (N_8222,N_3116,N_5814);
and U8223 (N_8223,N_4693,N_4877);
and U8224 (N_8224,N_5226,N_3381);
nor U8225 (N_8225,N_4694,N_5307);
nor U8226 (N_8226,N_5618,N_3905);
nand U8227 (N_8227,N_3611,N_3930);
xor U8228 (N_8228,N_3039,N_5214);
xor U8229 (N_8229,N_3891,N_3216);
nand U8230 (N_8230,N_3975,N_3891);
nand U8231 (N_8231,N_3178,N_5995);
xnor U8232 (N_8232,N_3693,N_3841);
nand U8233 (N_8233,N_4415,N_5371);
or U8234 (N_8234,N_4168,N_3425);
and U8235 (N_8235,N_3538,N_3324);
xor U8236 (N_8236,N_5308,N_5845);
nand U8237 (N_8237,N_5969,N_5310);
xor U8238 (N_8238,N_5251,N_5712);
xnor U8239 (N_8239,N_5767,N_4525);
nor U8240 (N_8240,N_5889,N_5833);
xnor U8241 (N_8241,N_4455,N_4785);
nor U8242 (N_8242,N_5291,N_5446);
nand U8243 (N_8243,N_5483,N_4241);
and U8244 (N_8244,N_5587,N_5858);
or U8245 (N_8245,N_4136,N_3453);
xnor U8246 (N_8246,N_3287,N_4654);
and U8247 (N_8247,N_4321,N_4846);
or U8248 (N_8248,N_5557,N_5568);
xor U8249 (N_8249,N_5302,N_5938);
xnor U8250 (N_8250,N_4331,N_4394);
or U8251 (N_8251,N_5572,N_3531);
xor U8252 (N_8252,N_5842,N_5009);
nand U8253 (N_8253,N_5870,N_4916);
nand U8254 (N_8254,N_5304,N_4888);
nor U8255 (N_8255,N_3396,N_3632);
or U8256 (N_8256,N_5748,N_3062);
xnor U8257 (N_8257,N_3737,N_3591);
or U8258 (N_8258,N_5638,N_4161);
and U8259 (N_8259,N_5604,N_5160);
or U8260 (N_8260,N_5344,N_5802);
and U8261 (N_8261,N_4449,N_4320);
nor U8262 (N_8262,N_4986,N_5164);
nand U8263 (N_8263,N_4446,N_4083);
and U8264 (N_8264,N_3298,N_5788);
and U8265 (N_8265,N_3910,N_4773);
and U8266 (N_8266,N_4147,N_3896);
xor U8267 (N_8267,N_5725,N_4675);
and U8268 (N_8268,N_4898,N_3569);
and U8269 (N_8269,N_3677,N_3558);
and U8270 (N_8270,N_5671,N_3065);
and U8271 (N_8271,N_3045,N_3758);
or U8272 (N_8272,N_3795,N_3735);
nor U8273 (N_8273,N_3218,N_5655);
nor U8274 (N_8274,N_3551,N_4284);
xnor U8275 (N_8275,N_3225,N_3622);
xnor U8276 (N_8276,N_3141,N_5261);
or U8277 (N_8277,N_5756,N_5743);
nand U8278 (N_8278,N_4574,N_3357);
or U8279 (N_8279,N_3121,N_3182);
and U8280 (N_8280,N_5469,N_5875);
or U8281 (N_8281,N_4828,N_3914);
and U8282 (N_8282,N_5515,N_5098);
or U8283 (N_8283,N_3133,N_4454);
nand U8284 (N_8284,N_3344,N_3714);
and U8285 (N_8285,N_5548,N_4937);
nand U8286 (N_8286,N_4429,N_3689);
or U8287 (N_8287,N_5614,N_3282);
and U8288 (N_8288,N_5970,N_5429);
and U8289 (N_8289,N_4838,N_3981);
nand U8290 (N_8290,N_4006,N_3479);
and U8291 (N_8291,N_4499,N_5305);
or U8292 (N_8292,N_3944,N_4494);
and U8293 (N_8293,N_4550,N_5013);
and U8294 (N_8294,N_5312,N_4064);
nor U8295 (N_8295,N_5428,N_4066);
nand U8296 (N_8296,N_4674,N_3955);
nor U8297 (N_8297,N_4526,N_3242);
or U8298 (N_8298,N_4008,N_5279);
nand U8299 (N_8299,N_3230,N_5286);
and U8300 (N_8300,N_3207,N_5706);
and U8301 (N_8301,N_3148,N_3105);
xor U8302 (N_8302,N_4141,N_4941);
nand U8303 (N_8303,N_4898,N_4074);
nor U8304 (N_8304,N_5200,N_3083);
and U8305 (N_8305,N_4590,N_3107);
and U8306 (N_8306,N_3833,N_3201);
nand U8307 (N_8307,N_3899,N_4219);
and U8308 (N_8308,N_4838,N_3959);
xnor U8309 (N_8309,N_3701,N_5719);
nand U8310 (N_8310,N_4060,N_3435);
xnor U8311 (N_8311,N_3489,N_4785);
and U8312 (N_8312,N_4434,N_4298);
nor U8313 (N_8313,N_5786,N_4270);
or U8314 (N_8314,N_4248,N_5293);
xnor U8315 (N_8315,N_5751,N_5793);
nand U8316 (N_8316,N_5718,N_3294);
xnor U8317 (N_8317,N_5004,N_5568);
nor U8318 (N_8318,N_4549,N_4930);
and U8319 (N_8319,N_3048,N_4263);
xor U8320 (N_8320,N_4034,N_4500);
nor U8321 (N_8321,N_3566,N_3470);
and U8322 (N_8322,N_4315,N_3662);
and U8323 (N_8323,N_4936,N_3116);
xnor U8324 (N_8324,N_4672,N_5441);
nor U8325 (N_8325,N_4618,N_4368);
or U8326 (N_8326,N_3728,N_3093);
xor U8327 (N_8327,N_5754,N_4453);
nand U8328 (N_8328,N_5976,N_5095);
or U8329 (N_8329,N_4647,N_4954);
nor U8330 (N_8330,N_5504,N_3277);
nor U8331 (N_8331,N_5292,N_5817);
xor U8332 (N_8332,N_5662,N_4297);
nor U8333 (N_8333,N_3102,N_3715);
or U8334 (N_8334,N_3193,N_5811);
nor U8335 (N_8335,N_3467,N_3755);
and U8336 (N_8336,N_5078,N_4824);
xor U8337 (N_8337,N_4000,N_4981);
and U8338 (N_8338,N_4129,N_5109);
nor U8339 (N_8339,N_3212,N_5279);
xnor U8340 (N_8340,N_4136,N_5349);
and U8341 (N_8341,N_3640,N_4587);
xor U8342 (N_8342,N_3125,N_4162);
xnor U8343 (N_8343,N_5517,N_4923);
nand U8344 (N_8344,N_3540,N_3562);
or U8345 (N_8345,N_4058,N_4682);
or U8346 (N_8346,N_3238,N_5410);
or U8347 (N_8347,N_5096,N_3166);
nor U8348 (N_8348,N_3219,N_4906);
or U8349 (N_8349,N_5714,N_5731);
nand U8350 (N_8350,N_5981,N_4922);
nand U8351 (N_8351,N_3649,N_4676);
or U8352 (N_8352,N_3198,N_3583);
xor U8353 (N_8353,N_3303,N_3100);
xnor U8354 (N_8354,N_3211,N_3309);
nor U8355 (N_8355,N_5364,N_3830);
and U8356 (N_8356,N_3244,N_3561);
xor U8357 (N_8357,N_5599,N_3877);
and U8358 (N_8358,N_5061,N_3761);
and U8359 (N_8359,N_4525,N_4181);
nor U8360 (N_8360,N_5675,N_3793);
or U8361 (N_8361,N_4122,N_5486);
nor U8362 (N_8362,N_3293,N_3673);
nor U8363 (N_8363,N_4725,N_4299);
xor U8364 (N_8364,N_4113,N_3871);
or U8365 (N_8365,N_4236,N_5295);
or U8366 (N_8366,N_4165,N_3265);
nor U8367 (N_8367,N_4886,N_3282);
and U8368 (N_8368,N_5612,N_4024);
and U8369 (N_8369,N_3192,N_4755);
or U8370 (N_8370,N_4950,N_4925);
xnor U8371 (N_8371,N_4855,N_5445);
or U8372 (N_8372,N_5623,N_3489);
nand U8373 (N_8373,N_5807,N_3875);
and U8374 (N_8374,N_4260,N_4304);
xor U8375 (N_8375,N_4511,N_4302);
nor U8376 (N_8376,N_3485,N_5233);
and U8377 (N_8377,N_4861,N_3235);
xor U8378 (N_8378,N_5906,N_5013);
nand U8379 (N_8379,N_4840,N_3122);
nand U8380 (N_8380,N_5858,N_3767);
or U8381 (N_8381,N_3591,N_3197);
and U8382 (N_8382,N_4685,N_5523);
or U8383 (N_8383,N_5106,N_5132);
and U8384 (N_8384,N_4675,N_5069);
or U8385 (N_8385,N_5933,N_3780);
and U8386 (N_8386,N_5706,N_5893);
and U8387 (N_8387,N_5197,N_5622);
nand U8388 (N_8388,N_3516,N_4777);
nand U8389 (N_8389,N_4611,N_4662);
nor U8390 (N_8390,N_4140,N_4904);
or U8391 (N_8391,N_5114,N_4851);
nor U8392 (N_8392,N_3704,N_5333);
or U8393 (N_8393,N_5279,N_3084);
and U8394 (N_8394,N_5502,N_4299);
nor U8395 (N_8395,N_3032,N_5165);
nor U8396 (N_8396,N_3347,N_4162);
and U8397 (N_8397,N_5652,N_4313);
xnor U8398 (N_8398,N_5278,N_5491);
xnor U8399 (N_8399,N_3933,N_4242);
xor U8400 (N_8400,N_5904,N_3909);
xor U8401 (N_8401,N_5119,N_4046);
nor U8402 (N_8402,N_4146,N_4833);
nor U8403 (N_8403,N_3212,N_4304);
nor U8404 (N_8404,N_3941,N_4455);
or U8405 (N_8405,N_5449,N_3216);
nor U8406 (N_8406,N_3574,N_4088);
nand U8407 (N_8407,N_3324,N_5600);
nor U8408 (N_8408,N_4834,N_4215);
and U8409 (N_8409,N_4761,N_4554);
nor U8410 (N_8410,N_3198,N_5789);
or U8411 (N_8411,N_3050,N_5484);
nor U8412 (N_8412,N_3001,N_3221);
and U8413 (N_8413,N_5062,N_5908);
nor U8414 (N_8414,N_3461,N_5087);
or U8415 (N_8415,N_4488,N_5333);
and U8416 (N_8416,N_3789,N_3736);
and U8417 (N_8417,N_5278,N_4307);
xor U8418 (N_8418,N_5650,N_3973);
xnor U8419 (N_8419,N_4524,N_3161);
nand U8420 (N_8420,N_4350,N_3005);
nor U8421 (N_8421,N_3642,N_4032);
and U8422 (N_8422,N_4204,N_3469);
and U8423 (N_8423,N_5733,N_5491);
xor U8424 (N_8424,N_5323,N_5730);
and U8425 (N_8425,N_3755,N_3418);
nand U8426 (N_8426,N_5528,N_5172);
nand U8427 (N_8427,N_3096,N_4274);
nand U8428 (N_8428,N_5073,N_4359);
nor U8429 (N_8429,N_3862,N_4886);
and U8430 (N_8430,N_5729,N_3872);
xor U8431 (N_8431,N_5124,N_3696);
xor U8432 (N_8432,N_4797,N_5740);
or U8433 (N_8433,N_5567,N_5651);
nor U8434 (N_8434,N_5901,N_4566);
nand U8435 (N_8435,N_3711,N_3789);
and U8436 (N_8436,N_3605,N_4581);
nor U8437 (N_8437,N_4356,N_4799);
nand U8438 (N_8438,N_3337,N_3822);
and U8439 (N_8439,N_3674,N_4187);
nor U8440 (N_8440,N_4839,N_4316);
or U8441 (N_8441,N_3835,N_3648);
or U8442 (N_8442,N_3749,N_5781);
and U8443 (N_8443,N_4594,N_5131);
xor U8444 (N_8444,N_3270,N_4138);
xnor U8445 (N_8445,N_4146,N_5133);
nand U8446 (N_8446,N_5709,N_5218);
or U8447 (N_8447,N_5154,N_5180);
nand U8448 (N_8448,N_3026,N_5949);
nand U8449 (N_8449,N_5300,N_4834);
and U8450 (N_8450,N_5754,N_4049);
nor U8451 (N_8451,N_4917,N_5514);
nand U8452 (N_8452,N_5894,N_4443);
and U8453 (N_8453,N_5953,N_5305);
xnor U8454 (N_8454,N_5436,N_3083);
nor U8455 (N_8455,N_5494,N_5768);
nand U8456 (N_8456,N_3677,N_5407);
nand U8457 (N_8457,N_5912,N_4319);
nor U8458 (N_8458,N_3733,N_5770);
nand U8459 (N_8459,N_4890,N_4250);
nor U8460 (N_8460,N_5255,N_3031);
nor U8461 (N_8461,N_5552,N_3293);
nand U8462 (N_8462,N_5559,N_4659);
and U8463 (N_8463,N_4927,N_4548);
nand U8464 (N_8464,N_4194,N_3957);
nand U8465 (N_8465,N_3086,N_4393);
and U8466 (N_8466,N_3171,N_3840);
nand U8467 (N_8467,N_3481,N_3009);
xnor U8468 (N_8468,N_5400,N_4297);
and U8469 (N_8469,N_3804,N_3469);
and U8470 (N_8470,N_3157,N_5486);
and U8471 (N_8471,N_5962,N_4144);
xnor U8472 (N_8472,N_3859,N_4585);
nand U8473 (N_8473,N_3173,N_3632);
and U8474 (N_8474,N_3060,N_5190);
nand U8475 (N_8475,N_3600,N_4786);
and U8476 (N_8476,N_3718,N_5125);
xor U8477 (N_8477,N_3721,N_4436);
xor U8478 (N_8478,N_5088,N_5554);
or U8479 (N_8479,N_5202,N_4431);
xnor U8480 (N_8480,N_5240,N_5540);
or U8481 (N_8481,N_5565,N_3591);
nor U8482 (N_8482,N_4710,N_5431);
nor U8483 (N_8483,N_3486,N_5816);
or U8484 (N_8484,N_5533,N_3313);
or U8485 (N_8485,N_4730,N_4239);
nor U8486 (N_8486,N_5843,N_5021);
nand U8487 (N_8487,N_3574,N_5686);
xnor U8488 (N_8488,N_5992,N_5228);
nand U8489 (N_8489,N_4291,N_4302);
nand U8490 (N_8490,N_3293,N_4982);
xnor U8491 (N_8491,N_5717,N_3203);
nor U8492 (N_8492,N_3506,N_4995);
xor U8493 (N_8493,N_3615,N_5217);
nor U8494 (N_8494,N_3545,N_4992);
and U8495 (N_8495,N_5747,N_5143);
or U8496 (N_8496,N_3842,N_4878);
xnor U8497 (N_8497,N_4821,N_3175);
nand U8498 (N_8498,N_5030,N_4491);
and U8499 (N_8499,N_5372,N_4669);
and U8500 (N_8500,N_3723,N_4333);
nor U8501 (N_8501,N_3291,N_3465);
nor U8502 (N_8502,N_3015,N_5548);
xor U8503 (N_8503,N_3623,N_5137);
nor U8504 (N_8504,N_4753,N_3377);
and U8505 (N_8505,N_4589,N_5026);
or U8506 (N_8506,N_5478,N_3925);
nor U8507 (N_8507,N_3726,N_3457);
and U8508 (N_8508,N_3595,N_3308);
and U8509 (N_8509,N_3603,N_3410);
xnor U8510 (N_8510,N_3493,N_4100);
and U8511 (N_8511,N_4249,N_3942);
xnor U8512 (N_8512,N_3516,N_4834);
nor U8513 (N_8513,N_5792,N_4322);
and U8514 (N_8514,N_4882,N_4085);
or U8515 (N_8515,N_5346,N_5010);
and U8516 (N_8516,N_5169,N_3330);
and U8517 (N_8517,N_4947,N_4230);
xnor U8518 (N_8518,N_5336,N_3974);
nand U8519 (N_8519,N_4336,N_4612);
nor U8520 (N_8520,N_3445,N_4060);
nor U8521 (N_8521,N_3381,N_3519);
nor U8522 (N_8522,N_4825,N_5746);
xor U8523 (N_8523,N_5060,N_5132);
xnor U8524 (N_8524,N_4280,N_4568);
nand U8525 (N_8525,N_4202,N_5335);
xor U8526 (N_8526,N_3634,N_5375);
xor U8527 (N_8527,N_5397,N_3114);
nor U8528 (N_8528,N_5029,N_5738);
and U8529 (N_8529,N_4280,N_5282);
nor U8530 (N_8530,N_5924,N_4250);
xnor U8531 (N_8531,N_3002,N_5769);
nor U8532 (N_8532,N_3734,N_4182);
xor U8533 (N_8533,N_5837,N_4104);
nor U8534 (N_8534,N_3843,N_4565);
or U8535 (N_8535,N_4383,N_4980);
nand U8536 (N_8536,N_3436,N_5955);
or U8537 (N_8537,N_5590,N_3024);
xnor U8538 (N_8538,N_4755,N_3698);
and U8539 (N_8539,N_5907,N_3956);
and U8540 (N_8540,N_5909,N_3514);
or U8541 (N_8541,N_3078,N_4970);
or U8542 (N_8542,N_5215,N_3899);
xnor U8543 (N_8543,N_5495,N_3868);
xnor U8544 (N_8544,N_5357,N_4206);
xnor U8545 (N_8545,N_5200,N_4514);
xnor U8546 (N_8546,N_3770,N_3031);
nand U8547 (N_8547,N_4709,N_5584);
nor U8548 (N_8548,N_4099,N_4234);
xor U8549 (N_8549,N_3356,N_3090);
or U8550 (N_8550,N_5137,N_3462);
nand U8551 (N_8551,N_4372,N_5130);
nor U8552 (N_8552,N_5807,N_3748);
nand U8553 (N_8553,N_4469,N_5683);
nor U8554 (N_8554,N_4000,N_4262);
nor U8555 (N_8555,N_5338,N_5403);
and U8556 (N_8556,N_3846,N_4100);
and U8557 (N_8557,N_3458,N_3680);
nor U8558 (N_8558,N_4595,N_3700);
nand U8559 (N_8559,N_5591,N_5607);
or U8560 (N_8560,N_5585,N_4798);
and U8561 (N_8561,N_5805,N_5134);
and U8562 (N_8562,N_3295,N_5291);
xor U8563 (N_8563,N_3953,N_3368);
nand U8564 (N_8564,N_5319,N_5910);
nand U8565 (N_8565,N_4387,N_3832);
nor U8566 (N_8566,N_3227,N_3940);
and U8567 (N_8567,N_5378,N_4242);
nor U8568 (N_8568,N_4379,N_3247);
and U8569 (N_8569,N_4937,N_5727);
nand U8570 (N_8570,N_5376,N_3590);
nand U8571 (N_8571,N_3497,N_5262);
nand U8572 (N_8572,N_5603,N_4954);
nand U8573 (N_8573,N_4714,N_4871);
and U8574 (N_8574,N_5091,N_5900);
or U8575 (N_8575,N_3292,N_4001);
nor U8576 (N_8576,N_3986,N_5446);
or U8577 (N_8577,N_4693,N_4997);
or U8578 (N_8578,N_4656,N_3926);
nand U8579 (N_8579,N_3857,N_4064);
xnor U8580 (N_8580,N_5813,N_4507);
and U8581 (N_8581,N_3843,N_3659);
xnor U8582 (N_8582,N_4673,N_5023);
xor U8583 (N_8583,N_3728,N_4987);
nor U8584 (N_8584,N_3144,N_3774);
nor U8585 (N_8585,N_4304,N_5809);
nor U8586 (N_8586,N_5961,N_4781);
and U8587 (N_8587,N_5333,N_3123);
xnor U8588 (N_8588,N_3163,N_3981);
or U8589 (N_8589,N_3525,N_3137);
nor U8590 (N_8590,N_3705,N_3610);
nor U8591 (N_8591,N_3613,N_5321);
or U8592 (N_8592,N_3732,N_4489);
or U8593 (N_8593,N_5698,N_5098);
and U8594 (N_8594,N_5008,N_3223);
xnor U8595 (N_8595,N_5308,N_5931);
and U8596 (N_8596,N_4235,N_3536);
or U8597 (N_8597,N_4645,N_4421);
nor U8598 (N_8598,N_5451,N_5423);
nor U8599 (N_8599,N_4586,N_4575);
nand U8600 (N_8600,N_5296,N_4526);
or U8601 (N_8601,N_3842,N_3346);
and U8602 (N_8602,N_4673,N_3067);
xor U8603 (N_8603,N_4816,N_3875);
xor U8604 (N_8604,N_4683,N_4223);
nand U8605 (N_8605,N_4689,N_3795);
or U8606 (N_8606,N_4623,N_5034);
nor U8607 (N_8607,N_4597,N_5457);
and U8608 (N_8608,N_5182,N_3422);
nor U8609 (N_8609,N_4925,N_3367);
nand U8610 (N_8610,N_4855,N_3514);
nor U8611 (N_8611,N_3117,N_3037);
and U8612 (N_8612,N_5669,N_4038);
nand U8613 (N_8613,N_5229,N_4848);
or U8614 (N_8614,N_3015,N_3839);
nor U8615 (N_8615,N_3656,N_3789);
xnor U8616 (N_8616,N_5915,N_5216);
nor U8617 (N_8617,N_4904,N_4188);
or U8618 (N_8618,N_5416,N_3337);
and U8619 (N_8619,N_4231,N_5136);
or U8620 (N_8620,N_3069,N_5329);
xnor U8621 (N_8621,N_4348,N_4487);
or U8622 (N_8622,N_3285,N_5617);
or U8623 (N_8623,N_3777,N_3813);
nand U8624 (N_8624,N_3623,N_4923);
xor U8625 (N_8625,N_4782,N_5831);
and U8626 (N_8626,N_3873,N_5550);
and U8627 (N_8627,N_5917,N_5674);
nor U8628 (N_8628,N_4810,N_3274);
xnor U8629 (N_8629,N_3407,N_5844);
and U8630 (N_8630,N_3965,N_5437);
nand U8631 (N_8631,N_3938,N_4312);
nand U8632 (N_8632,N_5133,N_3694);
xnor U8633 (N_8633,N_4797,N_3488);
or U8634 (N_8634,N_5510,N_5406);
nand U8635 (N_8635,N_5168,N_3339);
and U8636 (N_8636,N_3019,N_5040);
nor U8637 (N_8637,N_5158,N_5291);
xor U8638 (N_8638,N_3431,N_4411);
and U8639 (N_8639,N_5434,N_5365);
xor U8640 (N_8640,N_3393,N_4712);
or U8641 (N_8641,N_5914,N_3664);
and U8642 (N_8642,N_5506,N_4418);
or U8643 (N_8643,N_4274,N_4123);
xnor U8644 (N_8644,N_4216,N_3968);
xor U8645 (N_8645,N_5373,N_3558);
nand U8646 (N_8646,N_3725,N_3746);
and U8647 (N_8647,N_4782,N_3496);
nor U8648 (N_8648,N_4499,N_4162);
nand U8649 (N_8649,N_4331,N_4744);
and U8650 (N_8650,N_3937,N_4172);
or U8651 (N_8651,N_5138,N_5440);
nor U8652 (N_8652,N_3494,N_3746);
nand U8653 (N_8653,N_4914,N_5614);
nand U8654 (N_8654,N_5712,N_5325);
or U8655 (N_8655,N_5542,N_3116);
or U8656 (N_8656,N_3652,N_5737);
or U8657 (N_8657,N_3328,N_3578);
or U8658 (N_8658,N_4560,N_5928);
nand U8659 (N_8659,N_5785,N_4362);
xor U8660 (N_8660,N_4104,N_3902);
xor U8661 (N_8661,N_5601,N_4507);
and U8662 (N_8662,N_5625,N_3589);
xnor U8663 (N_8663,N_5099,N_4383);
nand U8664 (N_8664,N_5403,N_4700);
xnor U8665 (N_8665,N_4273,N_4430);
nor U8666 (N_8666,N_4556,N_4736);
xor U8667 (N_8667,N_3672,N_5986);
nand U8668 (N_8668,N_4684,N_4732);
nand U8669 (N_8669,N_3956,N_3172);
and U8670 (N_8670,N_3534,N_5068);
nand U8671 (N_8671,N_4675,N_3659);
and U8672 (N_8672,N_4696,N_4439);
nand U8673 (N_8673,N_4570,N_3952);
nand U8674 (N_8674,N_4111,N_5180);
nand U8675 (N_8675,N_3508,N_3311);
xor U8676 (N_8676,N_4461,N_3253);
nand U8677 (N_8677,N_4378,N_3607);
and U8678 (N_8678,N_4999,N_4776);
and U8679 (N_8679,N_3219,N_5949);
nor U8680 (N_8680,N_3636,N_3909);
xnor U8681 (N_8681,N_5230,N_4778);
and U8682 (N_8682,N_5713,N_3428);
or U8683 (N_8683,N_5336,N_5547);
nand U8684 (N_8684,N_3410,N_4563);
and U8685 (N_8685,N_4282,N_4583);
xor U8686 (N_8686,N_3570,N_5821);
xor U8687 (N_8687,N_3671,N_3899);
or U8688 (N_8688,N_3201,N_5257);
or U8689 (N_8689,N_4168,N_5053);
nor U8690 (N_8690,N_5861,N_3880);
or U8691 (N_8691,N_5650,N_3673);
xor U8692 (N_8692,N_5423,N_3639);
or U8693 (N_8693,N_5522,N_3151);
xor U8694 (N_8694,N_4776,N_3644);
and U8695 (N_8695,N_4187,N_5783);
xnor U8696 (N_8696,N_4006,N_3185);
or U8697 (N_8697,N_3701,N_3311);
or U8698 (N_8698,N_3154,N_3211);
or U8699 (N_8699,N_3590,N_4733);
nor U8700 (N_8700,N_4112,N_5906);
nor U8701 (N_8701,N_4390,N_3031);
xor U8702 (N_8702,N_4031,N_4991);
xor U8703 (N_8703,N_3282,N_3238);
nor U8704 (N_8704,N_5345,N_3154);
xor U8705 (N_8705,N_4321,N_4780);
and U8706 (N_8706,N_3908,N_3686);
xor U8707 (N_8707,N_3801,N_3432);
and U8708 (N_8708,N_5193,N_3372);
nor U8709 (N_8709,N_3235,N_4726);
xnor U8710 (N_8710,N_5271,N_5251);
nor U8711 (N_8711,N_4549,N_5468);
nor U8712 (N_8712,N_4789,N_5231);
xnor U8713 (N_8713,N_4286,N_3318);
nand U8714 (N_8714,N_5516,N_3525);
nand U8715 (N_8715,N_4710,N_3978);
nand U8716 (N_8716,N_4669,N_5114);
nor U8717 (N_8717,N_3254,N_4695);
nor U8718 (N_8718,N_3826,N_3767);
xor U8719 (N_8719,N_5313,N_3403);
and U8720 (N_8720,N_3804,N_3828);
nand U8721 (N_8721,N_4117,N_5766);
nand U8722 (N_8722,N_3621,N_4522);
nor U8723 (N_8723,N_5711,N_3924);
nand U8724 (N_8724,N_4656,N_3602);
nand U8725 (N_8725,N_4531,N_4299);
and U8726 (N_8726,N_5316,N_4624);
or U8727 (N_8727,N_5759,N_3069);
or U8728 (N_8728,N_5945,N_3296);
or U8729 (N_8729,N_5537,N_5486);
nor U8730 (N_8730,N_5409,N_3777);
xor U8731 (N_8731,N_3737,N_4005);
or U8732 (N_8732,N_4792,N_3355);
and U8733 (N_8733,N_5759,N_5872);
nand U8734 (N_8734,N_4656,N_4971);
and U8735 (N_8735,N_5196,N_4714);
nand U8736 (N_8736,N_3194,N_4710);
and U8737 (N_8737,N_4463,N_3234);
nand U8738 (N_8738,N_4258,N_4595);
nor U8739 (N_8739,N_5096,N_5687);
nand U8740 (N_8740,N_5397,N_5853);
nor U8741 (N_8741,N_4148,N_3791);
or U8742 (N_8742,N_4239,N_5725);
or U8743 (N_8743,N_3225,N_3249);
xor U8744 (N_8744,N_3421,N_4806);
nor U8745 (N_8745,N_4210,N_5198);
and U8746 (N_8746,N_5527,N_4342);
or U8747 (N_8747,N_4530,N_4631);
or U8748 (N_8748,N_3481,N_3840);
nand U8749 (N_8749,N_4447,N_3246);
and U8750 (N_8750,N_5334,N_4511);
xor U8751 (N_8751,N_5021,N_3882);
and U8752 (N_8752,N_5616,N_3909);
and U8753 (N_8753,N_4391,N_3459);
nor U8754 (N_8754,N_4991,N_4693);
nor U8755 (N_8755,N_3319,N_3128);
xor U8756 (N_8756,N_5518,N_3956);
or U8757 (N_8757,N_5413,N_5160);
nand U8758 (N_8758,N_4823,N_4258);
nand U8759 (N_8759,N_3012,N_3362);
xnor U8760 (N_8760,N_5326,N_5746);
or U8761 (N_8761,N_5964,N_3114);
or U8762 (N_8762,N_4406,N_3932);
or U8763 (N_8763,N_3384,N_3444);
or U8764 (N_8764,N_4006,N_5899);
nor U8765 (N_8765,N_4574,N_5059);
and U8766 (N_8766,N_5084,N_4923);
nand U8767 (N_8767,N_3167,N_4598);
nand U8768 (N_8768,N_5510,N_5986);
nand U8769 (N_8769,N_3167,N_5531);
xor U8770 (N_8770,N_4240,N_5432);
xor U8771 (N_8771,N_5511,N_5765);
or U8772 (N_8772,N_5560,N_3126);
nand U8773 (N_8773,N_5921,N_3468);
nor U8774 (N_8774,N_4047,N_5943);
or U8775 (N_8775,N_4064,N_4953);
xnor U8776 (N_8776,N_5046,N_4182);
nand U8777 (N_8777,N_5741,N_4745);
xor U8778 (N_8778,N_3263,N_5054);
xnor U8779 (N_8779,N_3417,N_3062);
nand U8780 (N_8780,N_5260,N_5875);
xnor U8781 (N_8781,N_3619,N_4613);
and U8782 (N_8782,N_3765,N_5895);
or U8783 (N_8783,N_3219,N_5044);
nand U8784 (N_8784,N_3110,N_5833);
nor U8785 (N_8785,N_5683,N_3270);
or U8786 (N_8786,N_4483,N_5873);
xnor U8787 (N_8787,N_3120,N_5814);
nor U8788 (N_8788,N_3918,N_3755);
nand U8789 (N_8789,N_3854,N_3107);
xor U8790 (N_8790,N_3323,N_5649);
and U8791 (N_8791,N_3900,N_4003);
and U8792 (N_8792,N_5147,N_4740);
xnor U8793 (N_8793,N_5179,N_3751);
or U8794 (N_8794,N_5703,N_4859);
nand U8795 (N_8795,N_4386,N_5838);
nand U8796 (N_8796,N_3408,N_5932);
nor U8797 (N_8797,N_4569,N_3698);
xnor U8798 (N_8798,N_3666,N_5041);
nand U8799 (N_8799,N_4643,N_5973);
xor U8800 (N_8800,N_4028,N_3779);
xnor U8801 (N_8801,N_5703,N_3836);
nand U8802 (N_8802,N_5745,N_4530);
and U8803 (N_8803,N_5301,N_3630);
xnor U8804 (N_8804,N_5467,N_5920);
or U8805 (N_8805,N_3090,N_3707);
nand U8806 (N_8806,N_4875,N_3487);
nor U8807 (N_8807,N_3404,N_3774);
nor U8808 (N_8808,N_4967,N_5366);
or U8809 (N_8809,N_4049,N_4918);
xor U8810 (N_8810,N_3315,N_3542);
nor U8811 (N_8811,N_5873,N_3323);
xor U8812 (N_8812,N_5156,N_4504);
xor U8813 (N_8813,N_5849,N_4087);
or U8814 (N_8814,N_3428,N_4360);
nor U8815 (N_8815,N_3918,N_3127);
or U8816 (N_8816,N_3029,N_4913);
or U8817 (N_8817,N_5688,N_3465);
or U8818 (N_8818,N_5983,N_5831);
nand U8819 (N_8819,N_5655,N_4659);
or U8820 (N_8820,N_5410,N_5137);
or U8821 (N_8821,N_4475,N_5914);
or U8822 (N_8822,N_4170,N_4663);
xor U8823 (N_8823,N_4966,N_4718);
and U8824 (N_8824,N_4851,N_4417);
nor U8825 (N_8825,N_3513,N_3408);
nor U8826 (N_8826,N_3491,N_4411);
or U8827 (N_8827,N_4764,N_5430);
xor U8828 (N_8828,N_3823,N_4988);
xor U8829 (N_8829,N_5584,N_5041);
nor U8830 (N_8830,N_3609,N_4255);
nand U8831 (N_8831,N_3934,N_4534);
nor U8832 (N_8832,N_4242,N_3206);
or U8833 (N_8833,N_5652,N_5536);
xor U8834 (N_8834,N_5684,N_4898);
and U8835 (N_8835,N_5997,N_3401);
or U8836 (N_8836,N_3685,N_3680);
xor U8837 (N_8837,N_5988,N_3850);
or U8838 (N_8838,N_3407,N_4140);
xnor U8839 (N_8839,N_4626,N_3073);
nor U8840 (N_8840,N_4982,N_4229);
and U8841 (N_8841,N_3226,N_4643);
and U8842 (N_8842,N_4415,N_5408);
nor U8843 (N_8843,N_4302,N_5295);
or U8844 (N_8844,N_3141,N_3726);
or U8845 (N_8845,N_4215,N_4528);
nor U8846 (N_8846,N_4271,N_4876);
or U8847 (N_8847,N_4198,N_3425);
nand U8848 (N_8848,N_4295,N_3963);
xor U8849 (N_8849,N_4852,N_3418);
nor U8850 (N_8850,N_4993,N_4074);
nor U8851 (N_8851,N_5123,N_4952);
nor U8852 (N_8852,N_4296,N_4547);
and U8853 (N_8853,N_5784,N_3652);
nand U8854 (N_8854,N_4958,N_3731);
and U8855 (N_8855,N_3826,N_3765);
or U8856 (N_8856,N_4171,N_4814);
xnor U8857 (N_8857,N_4805,N_4826);
or U8858 (N_8858,N_4407,N_5071);
and U8859 (N_8859,N_5032,N_3121);
xor U8860 (N_8860,N_5316,N_3713);
nand U8861 (N_8861,N_3921,N_3235);
nor U8862 (N_8862,N_3743,N_4865);
and U8863 (N_8863,N_3537,N_5913);
or U8864 (N_8864,N_4527,N_4228);
xor U8865 (N_8865,N_5306,N_3692);
xnor U8866 (N_8866,N_4944,N_5994);
nand U8867 (N_8867,N_5755,N_4252);
nand U8868 (N_8868,N_3960,N_5958);
and U8869 (N_8869,N_3913,N_3356);
nand U8870 (N_8870,N_5856,N_5847);
nand U8871 (N_8871,N_4612,N_4650);
xnor U8872 (N_8872,N_4960,N_5758);
or U8873 (N_8873,N_5307,N_3816);
xor U8874 (N_8874,N_3031,N_3768);
or U8875 (N_8875,N_4777,N_3143);
or U8876 (N_8876,N_4363,N_4218);
and U8877 (N_8877,N_5306,N_4925);
nand U8878 (N_8878,N_3542,N_5720);
nor U8879 (N_8879,N_4830,N_4018);
or U8880 (N_8880,N_3643,N_5146);
nor U8881 (N_8881,N_3134,N_5612);
nor U8882 (N_8882,N_5230,N_3767);
or U8883 (N_8883,N_3988,N_3805);
xor U8884 (N_8884,N_4156,N_5536);
or U8885 (N_8885,N_5697,N_4752);
and U8886 (N_8886,N_4779,N_4851);
and U8887 (N_8887,N_5137,N_3867);
or U8888 (N_8888,N_3844,N_3603);
or U8889 (N_8889,N_5954,N_3000);
xnor U8890 (N_8890,N_3310,N_3490);
nor U8891 (N_8891,N_4321,N_5884);
nor U8892 (N_8892,N_4901,N_3871);
xnor U8893 (N_8893,N_5050,N_4745);
or U8894 (N_8894,N_4698,N_5760);
xnor U8895 (N_8895,N_3076,N_5222);
nand U8896 (N_8896,N_5565,N_3147);
xnor U8897 (N_8897,N_4082,N_3013);
nand U8898 (N_8898,N_4753,N_4986);
nand U8899 (N_8899,N_4353,N_3759);
nor U8900 (N_8900,N_5912,N_5766);
xor U8901 (N_8901,N_4545,N_5730);
nor U8902 (N_8902,N_4348,N_4734);
nand U8903 (N_8903,N_4345,N_4131);
or U8904 (N_8904,N_3224,N_4999);
and U8905 (N_8905,N_3342,N_4759);
or U8906 (N_8906,N_5342,N_5919);
nor U8907 (N_8907,N_5705,N_5248);
and U8908 (N_8908,N_5292,N_3854);
nor U8909 (N_8909,N_5111,N_4503);
nor U8910 (N_8910,N_5644,N_4337);
xor U8911 (N_8911,N_3170,N_4432);
and U8912 (N_8912,N_4995,N_4803);
xor U8913 (N_8913,N_5265,N_4750);
and U8914 (N_8914,N_3722,N_3874);
nor U8915 (N_8915,N_5150,N_3864);
xnor U8916 (N_8916,N_4363,N_4274);
xor U8917 (N_8917,N_4788,N_4239);
nor U8918 (N_8918,N_3048,N_5419);
nor U8919 (N_8919,N_5176,N_5092);
nand U8920 (N_8920,N_5907,N_3466);
or U8921 (N_8921,N_3752,N_5986);
and U8922 (N_8922,N_3111,N_5017);
nand U8923 (N_8923,N_4372,N_5502);
and U8924 (N_8924,N_3040,N_4148);
xnor U8925 (N_8925,N_4110,N_3254);
and U8926 (N_8926,N_5896,N_5311);
nor U8927 (N_8927,N_5124,N_5297);
nand U8928 (N_8928,N_5167,N_5119);
or U8929 (N_8929,N_3773,N_4409);
nand U8930 (N_8930,N_3578,N_5506);
nor U8931 (N_8931,N_5247,N_4881);
xnor U8932 (N_8932,N_4359,N_3119);
nand U8933 (N_8933,N_3332,N_5427);
xnor U8934 (N_8934,N_4795,N_5035);
and U8935 (N_8935,N_5204,N_5312);
nor U8936 (N_8936,N_3629,N_3573);
xor U8937 (N_8937,N_3651,N_3501);
xor U8938 (N_8938,N_5220,N_5067);
or U8939 (N_8939,N_4830,N_4819);
nand U8940 (N_8940,N_4997,N_5636);
xnor U8941 (N_8941,N_3615,N_3943);
nand U8942 (N_8942,N_4161,N_3499);
nor U8943 (N_8943,N_3815,N_5935);
or U8944 (N_8944,N_3632,N_5465);
xor U8945 (N_8945,N_5622,N_3131);
nor U8946 (N_8946,N_3137,N_3161);
and U8947 (N_8947,N_3179,N_5623);
nor U8948 (N_8948,N_4828,N_4061);
nand U8949 (N_8949,N_5825,N_3202);
nor U8950 (N_8950,N_5577,N_4419);
and U8951 (N_8951,N_4237,N_3179);
or U8952 (N_8952,N_3521,N_4511);
nor U8953 (N_8953,N_4147,N_4638);
and U8954 (N_8954,N_4295,N_5878);
nor U8955 (N_8955,N_5115,N_5316);
or U8956 (N_8956,N_5398,N_4537);
or U8957 (N_8957,N_4098,N_5703);
nand U8958 (N_8958,N_3514,N_5366);
or U8959 (N_8959,N_4927,N_4192);
xor U8960 (N_8960,N_4860,N_3015);
xor U8961 (N_8961,N_3665,N_5921);
or U8962 (N_8962,N_4989,N_5219);
xor U8963 (N_8963,N_3174,N_4285);
or U8964 (N_8964,N_5920,N_4698);
xor U8965 (N_8965,N_4391,N_4167);
or U8966 (N_8966,N_4683,N_3296);
or U8967 (N_8967,N_5920,N_3006);
or U8968 (N_8968,N_3414,N_3029);
xnor U8969 (N_8969,N_3971,N_5333);
nand U8970 (N_8970,N_5981,N_5404);
nand U8971 (N_8971,N_5546,N_4266);
xor U8972 (N_8972,N_4199,N_5192);
xor U8973 (N_8973,N_3319,N_5106);
or U8974 (N_8974,N_3674,N_5923);
or U8975 (N_8975,N_5565,N_3358);
nand U8976 (N_8976,N_4373,N_5215);
and U8977 (N_8977,N_5224,N_4324);
nor U8978 (N_8978,N_4860,N_4213);
or U8979 (N_8979,N_4282,N_3410);
or U8980 (N_8980,N_4103,N_3542);
or U8981 (N_8981,N_4020,N_3156);
nand U8982 (N_8982,N_3682,N_5635);
nand U8983 (N_8983,N_3014,N_5589);
nand U8984 (N_8984,N_5619,N_3295);
nand U8985 (N_8985,N_3981,N_5745);
or U8986 (N_8986,N_4848,N_4053);
xor U8987 (N_8987,N_3915,N_3249);
or U8988 (N_8988,N_5643,N_5012);
xor U8989 (N_8989,N_4650,N_5031);
xnor U8990 (N_8990,N_5663,N_3260);
or U8991 (N_8991,N_3594,N_5359);
xnor U8992 (N_8992,N_5953,N_5078);
and U8993 (N_8993,N_3463,N_3809);
nand U8994 (N_8994,N_3713,N_4567);
or U8995 (N_8995,N_4419,N_5684);
nand U8996 (N_8996,N_4323,N_5884);
or U8997 (N_8997,N_5864,N_3354);
nand U8998 (N_8998,N_5843,N_5265);
and U8999 (N_8999,N_4983,N_4822);
nor U9000 (N_9000,N_8923,N_7763);
xnor U9001 (N_9001,N_7836,N_6601);
or U9002 (N_9002,N_6057,N_8686);
xnor U9003 (N_9003,N_6400,N_7645);
or U9004 (N_9004,N_8734,N_7270);
xor U9005 (N_9005,N_6841,N_8294);
xnor U9006 (N_9006,N_8284,N_7443);
or U9007 (N_9007,N_8693,N_8224);
or U9008 (N_9008,N_6399,N_6779);
nor U9009 (N_9009,N_7362,N_7091);
nand U9010 (N_9010,N_6247,N_6036);
nor U9011 (N_9011,N_7812,N_6404);
xor U9012 (N_9012,N_6969,N_8092);
or U9013 (N_9013,N_8278,N_7429);
nor U9014 (N_9014,N_6480,N_7550);
xnor U9015 (N_9015,N_7993,N_6052);
xnor U9016 (N_9016,N_6739,N_8003);
and U9017 (N_9017,N_8879,N_8221);
nor U9018 (N_9018,N_6003,N_8559);
nand U9019 (N_9019,N_7949,N_6960);
and U9020 (N_9020,N_7038,N_6668);
xnor U9021 (N_9021,N_8317,N_6890);
xnor U9022 (N_9022,N_7857,N_6616);
or U9023 (N_9023,N_8679,N_8688);
and U9024 (N_9024,N_7026,N_7722);
or U9025 (N_9025,N_7405,N_8189);
nor U9026 (N_9026,N_7962,N_6314);
or U9027 (N_9027,N_7285,N_8235);
nor U9028 (N_9028,N_6059,N_8549);
nand U9029 (N_9029,N_8727,N_7428);
xnor U9030 (N_9030,N_7290,N_6958);
and U9031 (N_9031,N_7663,N_8053);
or U9032 (N_9032,N_6849,N_8920);
nand U9033 (N_9033,N_6845,N_8709);
and U9034 (N_9034,N_6575,N_6089);
or U9035 (N_9035,N_7977,N_8758);
or U9036 (N_9036,N_8756,N_6352);
and U9037 (N_9037,N_8625,N_8861);
or U9038 (N_9038,N_8641,N_6632);
and U9039 (N_9039,N_8367,N_6118);
or U9040 (N_9040,N_6361,N_8319);
and U9041 (N_9041,N_8000,N_6800);
xor U9042 (N_9042,N_6097,N_7462);
nand U9043 (N_9043,N_7538,N_6513);
and U9044 (N_9044,N_8328,N_7546);
xnor U9045 (N_9045,N_8543,N_8241);
xor U9046 (N_9046,N_8884,N_8710);
or U9047 (N_9047,N_6514,N_7395);
xor U9048 (N_9048,N_8155,N_7080);
or U9049 (N_9049,N_8350,N_7626);
nand U9050 (N_9050,N_7312,N_6984);
nor U9051 (N_9051,N_7005,N_8311);
or U9052 (N_9052,N_7394,N_7619);
or U9053 (N_9053,N_8237,N_6682);
nand U9054 (N_9054,N_8843,N_6666);
and U9055 (N_9055,N_7522,N_8115);
xor U9056 (N_9056,N_6588,N_6294);
xnor U9057 (N_9057,N_7343,N_8131);
nor U9058 (N_9058,N_8841,N_8208);
and U9059 (N_9059,N_8724,N_7628);
xor U9060 (N_9060,N_8029,N_6270);
nand U9061 (N_9061,N_7473,N_6167);
nor U9062 (N_9062,N_7720,N_7564);
and U9063 (N_9063,N_7688,N_8965);
nor U9064 (N_9064,N_6913,N_7810);
nand U9065 (N_9065,N_7039,N_6406);
nand U9066 (N_9066,N_6563,N_7381);
nor U9067 (N_9067,N_7704,N_6181);
and U9068 (N_9068,N_8112,N_6851);
nor U9069 (N_9069,N_6536,N_6690);
or U9070 (N_9070,N_6872,N_6233);
xnor U9071 (N_9071,N_6834,N_8658);
or U9072 (N_9072,N_6810,N_7639);
nand U9073 (N_9073,N_8216,N_7274);
xnor U9074 (N_9074,N_7438,N_6466);
and U9075 (N_9075,N_8874,N_8139);
xnor U9076 (N_9076,N_8306,N_8191);
xor U9077 (N_9077,N_6805,N_7811);
xnor U9078 (N_9078,N_8668,N_6732);
nor U9079 (N_9079,N_7107,N_7533);
or U9080 (N_9080,N_6844,N_8816);
nand U9081 (N_9081,N_8747,N_7690);
nor U9082 (N_9082,N_8618,N_6101);
nor U9083 (N_9083,N_6398,N_8215);
nor U9084 (N_9084,N_7154,N_6564);
nor U9085 (N_9085,N_6343,N_8667);
nor U9086 (N_9086,N_8070,N_8116);
nor U9087 (N_9087,N_7576,N_6462);
nand U9088 (N_9088,N_6121,N_8381);
xnor U9089 (N_9089,N_6006,N_6134);
nor U9090 (N_9090,N_8907,N_6238);
and U9091 (N_9091,N_8852,N_7847);
and U9092 (N_9092,N_6223,N_8413);
nand U9093 (N_9093,N_8819,N_7435);
xor U9094 (N_9094,N_8334,N_7583);
nor U9095 (N_9095,N_8578,N_8105);
xor U9096 (N_9096,N_6370,N_8595);
and U9097 (N_9097,N_7127,N_7033);
and U9098 (N_9098,N_6735,N_7013);
nor U9099 (N_9099,N_8056,N_6344);
and U9100 (N_9100,N_8863,N_7212);
or U9101 (N_9101,N_8422,N_7465);
nand U9102 (N_9102,N_7578,N_8295);
nand U9103 (N_9103,N_7779,N_7043);
nor U9104 (N_9104,N_6329,N_6137);
nand U9105 (N_9105,N_8229,N_6792);
and U9106 (N_9106,N_7792,N_6371);
and U9107 (N_9107,N_8254,N_6642);
or U9108 (N_9108,N_6850,N_6523);
xor U9109 (N_9109,N_8050,N_7877);
and U9110 (N_9110,N_6700,N_7934);
or U9111 (N_9111,N_6661,N_6525);
nand U9112 (N_9112,N_7728,N_8486);
nor U9113 (N_9113,N_7407,N_6420);
xnor U9114 (N_9114,N_7320,N_8099);
nor U9115 (N_9115,N_6931,N_8028);
nor U9116 (N_9116,N_7958,N_7046);
nor U9117 (N_9117,N_8992,N_7304);
nand U9118 (N_9118,N_6983,N_8958);
nand U9119 (N_9119,N_8629,N_7859);
and U9120 (N_9120,N_6957,N_7928);
and U9121 (N_9121,N_8645,N_8019);
nor U9122 (N_9122,N_8172,N_7944);
and U9123 (N_9123,N_6771,N_8013);
or U9124 (N_9124,N_7382,N_8656);
xnor U9125 (N_9125,N_7062,N_8488);
and U9126 (N_9126,N_6533,N_8057);
nor U9127 (N_9127,N_6893,N_7879);
nand U9128 (N_9128,N_7537,N_6482);
nor U9129 (N_9129,N_6947,N_7098);
and U9130 (N_9130,N_8401,N_7016);
nor U9131 (N_9131,N_8630,N_8525);
xor U9132 (N_9132,N_7111,N_8010);
nand U9133 (N_9133,N_6070,N_6785);
and U9134 (N_9134,N_6626,N_7484);
and U9135 (N_9135,N_7729,N_6244);
xnor U9136 (N_9136,N_7229,N_6350);
nand U9137 (N_9137,N_6419,N_8123);
or U9138 (N_9138,N_6449,N_8394);
nor U9139 (N_9139,N_7331,N_6441);
or U9140 (N_9140,N_7641,N_7317);
xor U9141 (N_9141,N_8272,N_8043);
xnor U9142 (N_9142,N_6349,N_7615);
and U9143 (N_9143,N_6472,N_7687);
or U9144 (N_9144,N_6448,N_7444);
xor U9145 (N_9145,N_6226,N_7116);
nand U9146 (N_9146,N_6009,N_8507);
nand U9147 (N_9147,N_6055,N_6046);
and U9148 (N_9148,N_6173,N_8713);
nand U9149 (N_9149,N_6819,N_6393);
nand U9150 (N_9150,N_7432,N_8151);
nand U9151 (N_9151,N_6022,N_7825);
or U9152 (N_9152,N_8142,N_7195);
nand U9153 (N_9153,N_8416,N_7667);
or U9154 (N_9154,N_6993,N_8436);
xnor U9155 (N_9155,N_7560,N_8526);
and U9156 (N_9156,N_6122,N_6622);
and U9157 (N_9157,N_7893,N_7748);
xor U9158 (N_9158,N_8518,N_7913);
nand U9159 (N_9159,N_7677,N_8893);
nor U9160 (N_9160,N_7453,N_8736);
nor U9161 (N_9161,N_6534,N_6655);
or U9162 (N_9162,N_6997,N_7246);
nor U9163 (N_9163,N_7308,N_6681);
or U9164 (N_9164,N_6861,N_6551);
nand U9165 (N_9165,N_6503,N_7617);
and U9166 (N_9166,N_7069,N_6675);
nand U9167 (N_9167,N_7972,N_7796);
nor U9168 (N_9168,N_6092,N_8665);
nor U9169 (N_9169,N_6296,N_6593);
or U9170 (N_9170,N_7955,N_8828);
and U9171 (N_9171,N_7735,N_7581);
and U9172 (N_9172,N_6612,N_8210);
xnor U9173 (N_9173,N_8801,N_7151);
nand U9174 (N_9174,N_7666,N_6346);
xor U9175 (N_9175,N_7721,N_7723);
nor U9176 (N_9176,N_7064,N_7767);
nor U9177 (N_9177,N_8402,N_8777);
nor U9178 (N_9178,N_6124,N_6120);
or U9179 (N_9179,N_8046,N_6102);
xor U9180 (N_9180,N_7622,N_8261);
and U9181 (N_9181,N_7740,N_7500);
nor U9182 (N_9182,N_7613,N_6227);
and U9183 (N_9183,N_8240,N_8101);
nand U9184 (N_9184,N_6895,N_7421);
xor U9185 (N_9185,N_6859,N_6965);
xnor U9186 (N_9186,N_8790,N_8813);
nor U9187 (N_9187,N_6737,N_6899);
nand U9188 (N_9188,N_8459,N_6948);
nand U9189 (N_9189,N_6925,N_6922);
or U9190 (N_9190,N_7076,N_8177);
and U9191 (N_9191,N_6529,N_6248);
nand U9192 (N_9192,N_8792,N_6279);
nand U9193 (N_9193,N_6029,N_6475);
xnor U9194 (N_9194,N_8853,N_8798);
or U9195 (N_9195,N_7020,N_7670);
or U9196 (N_9196,N_6407,N_6772);
or U9197 (N_9197,N_6255,N_7717);
or U9198 (N_9198,N_7319,N_6709);
nor U9199 (N_9199,N_7142,N_7017);
nand U9200 (N_9200,N_6724,N_7650);
and U9201 (N_9201,N_7349,N_7359);
nor U9202 (N_9202,N_7420,N_7774);
and U9203 (N_9203,N_6162,N_6253);
nand U9204 (N_9204,N_8163,N_7618);
or U9205 (N_9205,N_6887,N_7526);
and U9206 (N_9206,N_6087,N_8995);
nor U9207 (N_9207,N_8829,N_6574);
or U9208 (N_9208,N_7542,N_6447);
or U9209 (N_9209,N_7237,N_6094);
or U9210 (N_9210,N_8972,N_6379);
nor U9211 (N_9211,N_6033,N_7745);
xor U9212 (N_9212,N_8872,N_6417);
xor U9213 (N_9213,N_8415,N_6275);
or U9214 (N_9214,N_7267,N_8657);
nand U9215 (N_9215,N_7345,N_8672);
xnor U9216 (N_9216,N_7881,N_7858);
nor U9217 (N_9217,N_8063,N_7335);
nor U9218 (N_9218,N_8204,N_7959);
and U9219 (N_9219,N_8122,N_7252);
xor U9220 (N_9220,N_8468,N_6694);
or U9221 (N_9221,N_8207,N_7263);
or U9222 (N_9222,N_8467,N_7146);
nand U9223 (N_9223,N_6271,N_7731);
nor U9224 (N_9224,N_7978,N_6334);
xnor U9225 (N_9225,N_7556,N_7070);
and U9226 (N_9226,N_8069,N_8379);
or U9227 (N_9227,N_8450,N_8639);
nor U9228 (N_9228,N_8303,N_6424);
or U9229 (N_9229,N_6035,N_7756);
nand U9230 (N_9230,N_7414,N_7044);
xnor U9231 (N_9231,N_6459,N_7848);
or U9232 (N_9232,N_8870,N_7943);
and U9233 (N_9233,N_7314,N_6421);
and U9234 (N_9234,N_6826,N_7430);
and U9235 (N_9235,N_6813,N_8466);
xnor U9236 (N_9236,N_6285,N_7684);
xor U9237 (N_9237,N_7783,N_6921);
nor U9238 (N_9238,N_8939,N_7964);
nor U9239 (N_9239,N_7924,N_6451);
nand U9240 (N_9240,N_6883,N_8458);
nand U9241 (N_9241,N_8347,N_8062);
nor U9242 (N_9242,N_6490,N_8624);
xor U9243 (N_9243,N_8596,N_7367);
nand U9244 (N_9244,N_7037,N_8969);
nor U9245 (N_9245,N_7544,N_8517);
or U9246 (N_9246,N_8814,N_8921);
and U9247 (N_9247,N_8882,N_7168);
xor U9248 (N_9248,N_7268,N_8095);
nor U9249 (N_9249,N_7074,N_8840);
nand U9250 (N_9250,N_8600,N_8901);
xor U9251 (N_9251,N_6532,N_7839);
or U9252 (N_9252,N_6967,N_7660);
xor U9253 (N_9253,N_8358,N_7036);
and U9254 (N_9254,N_6602,N_8546);
nor U9255 (N_9255,N_6540,N_8147);
or U9256 (N_9256,N_6438,N_7915);
nor U9257 (N_9257,N_8481,N_8904);
nor U9258 (N_9258,N_6064,N_7061);
nor U9259 (N_9259,N_8186,N_7797);
xnor U9260 (N_9260,N_6187,N_8502);
nand U9261 (N_9261,N_6415,N_7185);
xor U9262 (N_9262,N_6198,N_7876);
or U9263 (N_9263,N_8552,N_6988);
or U9264 (N_9264,N_7235,N_8523);
nand U9265 (N_9265,N_6986,N_7374);
nand U9266 (N_9266,N_7342,N_8375);
xor U9267 (N_9267,N_7310,N_7370);
nand U9268 (N_9268,N_6467,N_8434);
and U9269 (N_9269,N_6911,N_8174);
nand U9270 (N_9270,N_7002,N_7662);
xor U9271 (N_9271,N_6453,N_7422);
nor U9272 (N_9272,N_6470,N_8547);
and U9273 (N_9273,N_6541,N_8701);
and U9274 (N_9274,N_7824,N_8324);
nand U9275 (N_9275,N_8584,N_7883);
nor U9276 (N_9276,N_7244,N_6425);
xnor U9277 (N_9277,N_7031,N_6949);
xnor U9278 (N_9278,N_8789,N_8232);
nor U9279 (N_9279,N_7115,N_8566);
and U9280 (N_9280,N_7378,N_8049);
xor U9281 (N_9281,N_7179,N_6131);
nand U9282 (N_9282,N_6069,N_8737);
and U9283 (N_9283,N_8463,N_7592);
xnor U9284 (N_9284,N_6317,N_8193);
or U9285 (N_9285,N_8022,N_7770);
and U9286 (N_9286,N_8587,N_8397);
and U9287 (N_9287,N_7808,N_8760);
xnor U9288 (N_9288,N_6224,N_7322);
or U9289 (N_9289,N_7124,N_7806);
nor U9290 (N_9290,N_6816,N_8108);
xnor U9291 (N_9291,N_6138,N_6446);
xor U9292 (N_9292,N_8471,N_7776);
xor U9293 (N_9293,N_8589,N_6686);
and U9294 (N_9294,N_7846,N_8746);
nand U9295 (N_9295,N_7141,N_7777);
and U9296 (N_9296,N_8461,N_8900);
xnor U9297 (N_9297,N_6589,N_7574);
and U9298 (N_9298,N_6491,N_7898);
nor U9299 (N_9299,N_8372,N_6985);
nor U9300 (N_9300,N_7008,N_6896);
nor U9301 (N_9301,N_7910,N_7132);
nor U9302 (N_9302,N_7878,N_8527);
xnor U9303 (N_9303,N_8702,N_6943);
xor U9304 (N_9304,N_8411,N_7027);
nor U9305 (N_9305,N_8579,N_8539);
xnor U9306 (N_9306,N_7390,N_6873);
or U9307 (N_9307,N_7216,N_7372);
nor U9308 (N_9308,N_6879,N_7644);
and U9309 (N_9309,N_7239,N_7273);
nand U9310 (N_9310,N_8133,N_6869);
and U9311 (N_9311,N_8329,N_7392);
xnor U9312 (N_9312,N_8574,N_6099);
xor U9313 (N_9313,N_6782,N_7052);
or U9314 (N_9314,N_6904,N_6026);
nor U9315 (N_9315,N_8102,N_6875);
or U9316 (N_9316,N_6697,N_6038);
and U9317 (N_9317,N_8860,N_6884);
and U9318 (N_9318,N_8866,N_8898);
nor U9319 (N_9319,N_6372,N_6061);
nor U9320 (N_9320,N_6596,N_8794);
nand U9321 (N_9321,N_8945,N_6531);
nor U9322 (N_9322,N_8234,N_6355);
nand U9323 (N_9323,N_8824,N_8895);
xor U9324 (N_9324,N_8537,N_7819);
or U9325 (N_9325,N_8170,N_8779);
nor U9326 (N_9326,N_6753,N_6801);
and U9327 (N_9327,N_7575,N_7330);
and U9328 (N_9328,N_6456,N_8275);
nand U9329 (N_9329,N_7814,N_7693);
nand U9330 (N_9330,N_7327,N_7681);
or U9331 (N_9331,N_7144,N_7326);
nor U9332 (N_9332,N_7694,N_7358);
and U9333 (N_9333,N_7103,N_8808);
nor U9334 (N_9334,N_8017,N_7408);
nor U9335 (N_9335,N_7371,N_7366);
xor U9336 (N_9336,N_7925,N_8722);
nand U9337 (N_9337,N_8041,N_8273);
nand U9338 (N_9338,N_8716,N_7206);
and U9339 (N_9339,N_7266,N_7999);
or U9340 (N_9340,N_7213,N_6611);
and U9341 (N_9341,N_8058,N_6183);
nand U9342 (N_9342,N_6714,N_6920);
nor U9343 (N_9343,N_7968,N_8075);
nor U9344 (N_9344,N_7092,N_7869);
and U9345 (N_9345,N_7961,N_6923);
and U9346 (N_9346,N_6461,N_6288);
or U9347 (N_9347,N_7114,N_6790);
nor U9348 (N_9348,N_6292,N_8906);
and U9349 (N_9349,N_6074,N_8892);
or U9350 (N_9350,N_7799,N_6867);
nand U9351 (N_9351,N_6506,N_8280);
and U9352 (N_9352,N_7090,N_8339);
and U9353 (N_9353,N_6423,N_6062);
nor U9354 (N_9354,N_7710,N_7035);
nor U9355 (N_9355,N_6505,N_7531);
xnor U9356 (N_9356,N_8555,N_8869);
nor U9357 (N_9357,N_8944,N_8940);
or U9358 (N_9358,N_6312,N_8754);
nor U9359 (N_9359,N_6888,N_8961);
xnor U9360 (N_9360,N_7634,N_6569);
nand U9361 (N_9361,N_7354,N_6909);
nand U9362 (N_9362,N_8289,N_7757);
nand U9363 (N_9363,N_6336,N_7954);
nand U9364 (N_9364,N_6469,N_7389);
and U9365 (N_9365,N_7772,N_7614);
xnor U9366 (N_9366,N_6373,N_6658);
nand U9367 (N_9367,N_6796,N_8744);
or U9368 (N_9368,N_6818,N_6037);
and U9369 (N_9369,N_6460,N_7970);
nand U9370 (N_9370,N_7568,N_6761);
and U9371 (N_9371,N_8315,N_8187);
xnor U9372 (N_9372,N_8815,N_7336);
nand U9373 (N_9373,N_7908,N_7073);
and U9374 (N_9374,N_6866,N_6231);
and U9375 (N_9375,N_6891,N_6580);
nand U9376 (N_9376,N_8694,N_8855);
nor U9377 (N_9377,N_6959,N_8001);
or U9378 (N_9378,N_8363,N_6304);
or U9379 (N_9379,N_8117,N_7988);
nand U9380 (N_9380,N_8928,N_8960);
or U9381 (N_9381,N_7922,N_8627);
nor U9382 (N_9382,N_8955,N_8909);
xor U9383 (N_9383,N_8024,N_8532);
and U9384 (N_9384,N_7623,N_6797);
xor U9385 (N_9385,N_7328,N_7761);
nor U9386 (N_9386,N_7605,N_7313);
or U9387 (N_9387,N_6865,N_7265);
nor U9388 (N_9388,N_7837,N_8602);
nand U9389 (N_9389,N_8757,N_7021);
xor U9390 (N_9390,N_8642,N_7165);
or U9391 (N_9391,N_8188,N_6075);
or U9392 (N_9392,N_7384,N_7896);
nor U9393 (N_9393,N_8809,N_6090);
nand U9394 (N_9394,N_8355,N_8078);
xor U9395 (N_9395,N_6148,N_6045);
and U9396 (N_9396,N_8690,N_8932);
xnor U9397 (N_9397,N_6486,N_6669);
nor U9398 (N_9398,N_8292,N_8180);
xor U9399 (N_9399,N_6319,N_7991);
or U9400 (N_9400,N_8084,N_8290);
nand U9401 (N_9401,N_6678,N_8321);
nor U9402 (N_9402,N_8025,N_8055);
xor U9403 (N_9403,N_6998,N_6008);
nor U9404 (N_9404,N_6305,N_8395);
xor U9405 (N_9405,N_7034,N_7459);
and U9406 (N_9406,N_8141,N_7791);
or U9407 (N_9407,N_7351,N_7668);
and U9408 (N_9408,N_7937,N_6409);
nor U9409 (N_9409,N_6284,N_7191);
xor U9410 (N_9410,N_6807,N_6956);
xor U9411 (N_9411,N_6110,N_7109);
nand U9412 (N_9412,N_8603,N_7516);
and U9413 (N_9413,N_6591,N_8330);
nand U9414 (N_9414,N_8873,N_7441);
or U9415 (N_9415,N_6507,N_6430);
or U9416 (N_9416,N_7306,N_8501);
or U9417 (N_9417,N_6768,N_6144);
nor U9418 (N_9418,N_8717,N_7673);
nor U9419 (N_9419,N_6154,N_6366);
nand U9420 (N_9420,N_8382,N_6071);
or U9421 (N_9421,N_7227,N_6687);
xor U9422 (N_9422,N_7169,N_7249);
nor U9423 (N_9423,N_7851,N_8277);
xnor U9424 (N_9424,N_8785,N_6488);
xor U9425 (N_9425,N_7502,N_6358);
xor U9426 (N_9426,N_8137,N_6951);
and U9427 (N_9427,N_6060,N_7903);
nor U9428 (N_9428,N_6500,N_7852);
nand U9429 (N_9429,N_6915,N_8606);
nand U9430 (N_9430,N_6740,N_7000);
nor U9431 (N_9431,N_8726,N_7921);
or U9432 (N_9432,N_7765,N_6539);
or U9433 (N_9433,N_8862,N_8265);
and U9434 (N_9434,N_8033,N_8836);
nand U9435 (N_9435,N_7637,N_8570);
xor U9436 (N_9436,N_8268,N_7601);
xnor U9437 (N_9437,N_6163,N_6741);
nor U9438 (N_9438,N_6520,N_8362);
xnor U9439 (N_9439,N_6696,N_7809);
nand U9440 (N_9440,N_8993,N_7198);
and U9441 (N_9441,N_8765,N_6995);
and U9442 (N_9442,N_6197,N_6780);
nand U9443 (N_9443,N_7579,N_7099);
nand U9444 (N_9444,N_8957,N_7084);
xnor U9445 (N_9445,N_7167,N_7815);
and U9446 (N_9446,N_7888,N_8633);
nand U9447 (N_9447,N_8768,N_8035);
nor U9448 (N_9448,N_7256,N_8729);
xnor U9449 (N_9449,N_8244,N_8966);
xor U9450 (N_9450,N_6458,N_7194);
xnor U9451 (N_9451,N_8905,N_6202);
nand U9452 (N_9452,N_7163,N_6261);
nand U9453 (N_9453,N_6839,N_7510);
xnor U9454 (N_9454,N_7255,N_7205);
nor U9455 (N_9455,N_7834,N_6360);
xnor U9456 (N_9456,N_7166,N_6135);
nand U9457 (N_9457,N_8061,N_8634);
or U9458 (N_9458,N_6628,N_6191);
nor U9459 (N_9459,N_7451,N_7171);
nand U9460 (N_9460,N_6734,N_8264);
nor U9461 (N_9461,N_8257,N_7741);
xor U9462 (N_9462,N_7023,N_6684);
nand U9463 (N_9463,N_7347,N_8669);
and U9464 (N_9464,N_8671,N_8886);
nand U9465 (N_9465,N_6030,N_7009);
nor U9466 (N_9466,N_6338,N_7143);
nor U9467 (N_9467,N_6463,N_8298);
nand U9468 (N_9468,N_8619,N_7826);
nor U9469 (N_9469,N_8697,N_8357);
and U9470 (N_9470,N_6212,N_6321);
or U9471 (N_9471,N_6830,N_6141);
nand U9472 (N_9472,N_8090,N_7129);
nor U9473 (N_9473,N_6186,N_6710);
nand U9474 (N_9474,N_8585,N_8930);
nor U9475 (N_9475,N_7041,N_8512);
nor U9476 (N_9476,N_7685,N_6422);
nand U9477 (N_9477,N_6001,N_6776);
and U9478 (N_9478,N_7584,N_6232);
nor U9479 (N_9479,N_6243,N_8677);
or U9480 (N_9480,N_6190,N_7679);
nand U9481 (N_9481,N_7203,N_6679);
and U9482 (N_9482,N_6041,N_8296);
nor U9483 (N_9483,N_8089,N_7174);
and U9484 (N_9484,N_6582,N_8408);
or U9485 (N_9485,N_6556,N_6145);
nand U9486 (N_9486,N_7802,N_7751);
and U9487 (N_9487,N_7104,N_8446);
xnor U9488 (N_9488,N_7933,N_6147);
nand U9489 (N_9489,N_6157,N_6149);
or U9490 (N_9490,N_7400,N_8857);
and U9491 (N_9491,N_6201,N_7736);
nor U9492 (N_9492,N_8494,N_8389);
or U9493 (N_9493,N_7277,N_6013);
xnor U9494 (N_9494,N_7178,N_6499);
and U9495 (N_9495,N_6667,N_6395);
or U9496 (N_9496,N_6603,N_7133);
and U9497 (N_9497,N_6019,N_6620);
or U9498 (N_9498,N_7475,N_8127);
nor U9499 (N_9499,N_6953,N_7953);
and U9500 (N_9500,N_7085,N_6765);
and U9501 (N_9501,N_6111,N_8655);
xnor U9502 (N_9502,N_8676,N_7515);
and U9503 (N_9503,N_6560,N_8077);
nor U9504 (N_9504,N_8691,N_8822);
and U9505 (N_9505,N_7676,N_6128);
or U9506 (N_9506,N_8313,N_6945);
or U9507 (N_9507,N_6236,N_6471);
nand U9508 (N_9508,N_6929,N_6527);
xnor U9509 (N_9509,N_6464,N_8751);
nand U9510 (N_9510,N_7674,N_7134);
nand U9511 (N_9511,N_8225,N_7495);
nand U9512 (N_9512,N_7786,N_8659);
xor U9513 (N_9513,N_7539,N_8154);
and U9514 (N_9514,N_7973,N_6924);
xor U9515 (N_9515,N_8250,N_6397);
or U9516 (N_9516,N_8333,N_7631);
nor U9517 (N_9517,N_6707,N_8536);
xor U9518 (N_9518,N_8610,N_8803);
xor U9519 (N_9519,N_6117,N_7996);
nor U9520 (N_9520,N_6543,N_7042);
nor U9521 (N_9521,N_8977,N_7590);
nor U9522 (N_9522,N_6384,N_8636);
and U9523 (N_9523,N_8800,N_8811);
nor U9524 (N_9524,N_7892,N_6939);
nor U9525 (N_9525,N_8414,N_7785);
xor U9526 (N_9526,N_8678,N_7920);
nor U9527 (N_9527,N_6809,N_6129);
and U9528 (N_9528,N_7175,N_6368);
nand U9529 (N_9529,N_6367,N_6802);
and U9530 (N_9530,N_6085,N_7425);
or U9531 (N_9531,N_8767,N_8598);
and U9532 (N_9532,N_8877,N_8554);
xnor U9533 (N_9533,N_6583,N_7573);
nor U9534 (N_9534,N_6854,N_6014);
xor U9535 (N_9535,N_7596,N_7822);
or U9536 (N_9536,N_7749,N_6429);
nand U9537 (N_9537,N_6562,N_8297);
nand U9538 (N_9538,N_6511,N_6629);
nor U9539 (N_9539,N_8764,N_7353);
or U9540 (N_9540,N_7672,N_7396);
nand U9541 (N_9541,N_6114,N_8192);
xor U9542 (N_9542,N_8424,N_8071);
and U9543 (N_9543,N_7849,N_6932);
nor U9544 (N_9544,N_7015,N_6440);
and U9545 (N_9545,N_7329,N_6299);
xor U9546 (N_9546,N_6205,N_6342);
nand U9547 (N_9547,N_6389,N_8370);
nor U9548 (N_9548,N_8715,N_6549);
or U9549 (N_9549,N_7466,N_7967);
nand U9550 (N_9550,N_8844,N_8996);
and U9551 (N_9551,N_7007,N_7057);
nand U9552 (N_9552,N_6260,N_8111);
or U9553 (N_9553,N_6068,N_8439);
nand U9554 (N_9554,N_8426,N_8138);
or U9555 (N_9555,N_7240,N_8612);
or U9556 (N_9556,N_7818,N_8432);
xnor U9557 (N_9557,N_6699,N_8699);
xor U9558 (N_9558,N_7804,N_6952);
or U9559 (N_9559,N_6307,N_6095);
nor U9560 (N_9560,N_6657,N_6894);
nand U9561 (N_9561,N_8851,N_8005);
nor U9562 (N_9562,N_8968,N_6538);
nand U9563 (N_9563,N_7840,N_6199);
nor U9564 (N_9564,N_6643,N_7498);
nor U9565 (N_9565,N_7629,N_7207);
and U9566 (N_9566,N_7437,N_7984);
xor U9567 (N_9567,N_8008,N_6572);
xnor U9568 (N_9568,N_8302,N_6347);
or U9569 (N_9569,N_8827,N_8805);
xnor U9570 (N_9570,N_8399,N_7279);
xor U9571 (N_9571,N_7552,N_7162);
nand U9572 (N_9572,N_7588,N_8664);
and U9573 (N_9573,N_7535,N_6954);
and U9574 (N_9574,N_8875,N_7932);
xor U9575 (N_9575,N_7901,N_6719);
xor U9576 (N_9576,N_7415,N_6457);
or U9577 (N_9577,N_8126,N_7222);
or U9578 (N_9578,N_6573,N_6266);
xor U9579 (N_9579,N_6254,N_8941);
xnor U9580 (N_9580,N_8839,N_7398);
xnor U9581 (N_9581,N_6341,N_7974);
nand U9582 (N_9582,N_8750,N_8136);
or U9583 (N_9583,N_7211,N_8073);
xnor U9584 (N_9584,N_7594,N_7145);
and U9585 (N_9585,N_7947,N_6720);
nand U9586 (N_9586,N_7833,N_8037);
nor U9587 (N_9587,N_7773,N_8183);
or U9588 (N_9588,N_8868,N_8107);
and U9589 (N_9589,N_8020,N_6208);
nand U9590 (N_9590,N_8454,N_6310);
or U9591 (N_9591,N_8119,N_7449);
xnor U9592 (N_9592,N_6885,N_8648);
nor U9593 (N_9593,N_7737,N_7902);
and U9594 (N_9594,N_6633,N_7176);
nand U9595 (N_9595,N_8453,N_6824);
nand U9596 (N_9596,N_7880,N_7714);
nor U9597 (N_9597,N_6717,N_8711);
nand U9598 (N_9598,N_7764,N_6857);
or U9599 (N_9599,N_6320,N_6808);
or U9600 (N_9600,N_8451,N_6789);
xnor U9601 (N_9601,N_6412,N_8376);
or U9602 (N_9602,N_8462,N_7391);
or U9603 (N_9603,N_8769,N_6192);
nor U9604 (N_9604,N_8165,N_6093);
xor U9605 (N_9605,N_7344,N_8963);
xnor U9606 (N_9606,N_7950,N_6903);
xnor U9607 (N_9607,N_6091,N_7957);
nand U9608 (N_9608,N_7760,N_8258);
nand U9609 (N_9609,N_6812,N_7558);
or U9610 (N_9610,N_7884,N_8807);
nand U9611 (N_9611,N_6084,N_7204);
xor U9612 (N_9612,N_8674,N_6002);
and U9613 (N_9613,N_6829,N_7669);
xnor U9614 (N_9614,N_6553,N_6123);
or U9615 (N_9615,N_8040,N_6301);
and U9616 (N_9616,N_8293,N_6786);
and U9617 (N_9617,N_6970,N_7938);
and U9618 (N_9618,N_7768,N_8034);
nor U9619 (N_9619,N_6476,N_6578);
nand U9620 (N_9620,N_8983,N_6215);
nand U9621 (N_9621,N_8149,N_7985);
xor U9622 (N_9622,N_6179,N_7380);
and U9623 (N_9623,N_6241,N_7828);
and U9624 (N_9624,N_8572,N_7769);
or U9625 (N_9625,N_7753,N_7295);
or U9626 (N_9626,N_6585,N_8247);
or U9627 (N_9627,N_6736,N_6918);
or U9628 (N_9628,N_7457,N_7247);
xor U9629 (N_9629,N_7424,N_8222);
xor U9630 (N_9630,N_6762,N_6676);
nor U9631 (N_9631,N_7060,N_8903);
nand U9632 (N_9632,N_8644,N_8964);
nand U9633 (N_9633,N_7989,N_7572);
nand U9634 (N_9634,N_8212,N_8514);
nand U9635 (N_9635,N_8430,N_6252);
nor U9636 (N_9636,N_6160,N_8283);
or U9637 (N_9637,N_8745,N_6671);
nor U9638 (N_9638,N_6518,N_8156);
and U9639 (N_9639,N_6176,N_6004);
or U9640 (N_9640,N_6437,N_8014);
xnor U9641 (N_9641,N_7598,N_7707);
xor U9642 (N_9642,N_6515,N_8135);
nor U9643 (N_9643,N_7136,N_8684);
nand U9644 (N_9644,N_6431,N_8325);
xor U9645 (N_9645,N_6664,N_8490);
and U9646 (N_9646,N_7232,N_6049);
nor U9647 (N_9647,N_7416,N_6597);
nand U9648 (N_9648,N_7245,N_8447);
xor U9649 (N_9649,N_7128,N_7460);
or U9650 (N_9650,N_6015,N_8615);
or U9651 (N_9651,N_8643,N_6392);
nand U9652 (N_9652,N_6230,N_7160);
and U9653 (N_9653,N_6638,N_8652);
and U9654 (N_9654,N_6610,N_8831);
xor U9655 (N_9655,N_7325,N_7942);
nor U9656 (N_9656,N_6249,N_8125);
and U9657 (N_9657,N_6258,N_6337);
xnor U9658 (N_9658,N_7602,N_8505);
and U9659 (N_9659,N_6853,N_6917);
xnor U9660 (N_9660,N_7047,N_8609);
or U9661 (N_9661,N_7716,N_8740);
nand U9662 (N_9662,N_6222,N_6674);
or U9663 (N_9663,N_7611,N_6308);
nand U9664 (N_9664,N_6938,N_7916);
and U9665 (N_9665,N_8167,N_6414);
or U9666 (N_9666,N_8196,N_6537);
nor U9667 (N_9667,N_6428,N_7965);
xor U9668 (N_9668,N_7816,N_8924);
or U9669 (N_9669,N_7789,N_6277);
nand U9670 (N_9670,N_8804,N_7093);
xnor U9671 (N_9671,N_7140,N_8530);
nand U9672 (N_9672,N_8558,N_6754);
xor U9673 (N_9673,N_6439,N_6332);
xor U9674 (N_9674,N_6862,N_8739);
and U9675 (N_9675,N_8067,N_8281);
and U9676 (N_9676,N_6433,N_8442);
xnor U9677 (N_9677,N_6498,N_8495);
nand U9678 (N_9678,N_6587,N_6774);
nand U9679 (N_9679,N_7724,N_8120);
nor U9680 (N_9680,N_8299,N_7895);
xor U9681 (N_9681,N_7711,N_8012);
and U9682 (N_9682,N_6526,N_6650);
nor U9683 (N_9683,N_7800,N_7001);
nand U9684 (N_9684,N_8556,N_6053);
nor U9685 (N_9685,N_8477,N_6760);
nor U9686 (N_9686,N_6185,N_6410);
nor U9687 (N_9687,N_8304,N_6711);
nor U9688 (N_9688,N_8557,N_7272);
nand U9689 (N_9689,N_6979,N_7096);
nand U9690 (N_9690,N_8007,N_6528);
xnor U9691 (N_9691,N_8931,N_8799);
or U9692 (N_9692,N_8400,N_7242);
or U9693 (N_9693,N_7488,N_7433);
nand U9694 (N_9694,N_7383,N_7653);
nor U9695 (N_9695,N_8047,N_8974);
or U9696 (N_9696,N_8475,N_7439);
and U9697 (N_9697,N_8988,N_6113);
and U9698 (N_9698,N_7333,N_6827);
and U9699 (N_9699,N_6391,N_6554);
xnor U9700 (N_9700,N_8223,N_6325);
nor U9701 (N_9701,N_8646,N_7838);
nand U9702 (N_9702,N_6713,N_6758);
nor U9703 (N_9703,N_8337,N_7744);
xnor U9704 (N_9704,N_8979,N_7940);
nor U9705 (N_9705,N_6592,N_7927);
or U9706 (N_9706,N_8953,N_6881);
nor U9707 (N_9707,N_6725,N_7734);
or U9708 (N_9708,N_7431,N_7478);
nand U9709 (N_9709,N_6784,N_8184);
nor U9710 (N_9710,N_6432,N_7939);
xor U9711 (N_9711,N_8348,N_6571);
xor U9712 (N_9712,N_7226,N_6262);
and U9713 (N_9713,N_6550,N_8231);
nor U9714 (N_9714,N_8696,N_6302);
and U9715 (N_9715,N_8548,N_6474);
or U9716 (N_9716,N_6973,N_8285);
nor U9717 (N_9717,N_7998,N_6027);
nand U9718 (N_9718,N_8894,N_6644);
and U9719 (N_9719,N_7496,N_8509);
nor U9720 (N_9720,N_7455,N_8956);
nand U9721 (N_9721,N_6450,N_6383);
nor U9722 (N_9722,N_8718,N_8692);
xor U9723 (N_9723,N_8535,N_6443);
nor U9724 (N_9724,N_6625,N_6673);
and U9725 (N_9725,N_7562,N_8899);
nand U9726 (N_9726,N_7610,N_8749);
xnor U9727 (N_9727,N_6656,N_7040);
nor U9728 (N_9728,N_8480,N_6799);
or U9729 (N_9729,N_6509,N_8551);
xnor U9730 (N_9730,N_7149,N_6989);
xor U9731 (N_9731,N_7332,N_7885);
nor U9732 (N_9732,N_7491,N_6142);
nor U9733 (N_9733,N_8386,N_6811);
xor U9734 (N_9734,N_6568,N_7208);
xor U9735 (N_9735,N_8622,N_7807);
and U9736 (N_9736,N_8307,N_6729);
nand U9737 (N_9737,N_7117,N_7508);
xor U9738 (N_9738,N_8858,N_6005);
nand U9739 (N_9739,N_8211,N_7147);
xnor U9740 (N_9740,N_6274,N_8218);
or U9741 (N_9741,N_7250,N_6240);
xnor U9742 (N_9742,N_6382,N_6100);
nand U9743 (N_9743,N_7682,N_8663);
or U9744 (N_9744,N_7919,N_8914);
nor U9745 (N_9745,N_6139,N_6411);
or U9746 (N_9746,N_8593,N_6695);
nor U9747 (N_9747,N_7640,N_6290);
nand U9748 (N_9748,N_8775,N_8885);
nor U9749 (N_9749,N_6501,N_7671);
nor U9750 (N_9750,N_6598,N_8360);
xnor U9751 (N_9751,N_6207,N_8795);
xor U9752 (N_9752,N_6031,N_8344);
nand U9753 (N_9753,N_7570,N_8732);
or U9754 (N_9754,N_8152,N_6976);
or U9755 (N_9755,N_6722,N_6946);
nor U9756 (N_9756,N_6645,N_7340);
or U9757 (N_9757,N_7385,N_8999);
nand U9758 (N_9758,N_7221,N_8823);
or U9759 (N_9759,N_8708,N_6825);
nand U9760 (N_9760,N_6318,N_8985);
nand U9761 (N_9761,N_6613,N_7647);
and U9762 (N_9762,N_7830,N_7705);
nand U9763 (N_9763,N_6619,N_8452);
nor U9764 (N_9764,N_6390,N_8651);
nor U9765 (N_9765,N_7643,N_8849);
and U9766 (N_9766,N_6376,N_7440);
xnor U9767 (N_9767,N_8087,N_8243);
xnor U9768 (N_9768,N_8607,N_8908);
or U9769 (N_9769,N_6933,N_8410);
nand U9770 (N_9770,N_6795,N_7680);
xnor U9771 (N_9771,N_8145,N_6287);
xor U9772 (N_9772,N_8169,N_7102);
xor U9773 (N_9773,N_6333,N_6775);
xor U9774 (N_9774,N_7831,N_7130);
or U9775 (N_9775,N_7291,N_6685);
nand U9776 (N_9776,N_7202,N_8378);
nand U9777 (N_9777,N_6189,N_8383);
and U9778 (N_9778,N_6750,N_8393);
nand U9779 (N_9779,N_8233,N_6659);
nand U9780 (N_9780,N_6755,N_6401);
and U9781 (N_9781,N_8103,N_6096);
xnor U9782 (N_9782,N_6018,N_6738);
or U9783 (N_9783,N_7604,N_6703);
or U9784 (N_9784,N_6213,N_7311);
or U9785 (N_9785,N_8065,N_6555);
or U9786 (N_9786,N_8279,N_8009);
xor U9787 (N_9787,N_8605,N_7719);
xor U9788 (N_9788,N_6257,N_6126);
or U9789 (N_9789,N_7845,N_7254);
and U9790 (N_9790,N_7150,N_7118);
xnor U9791 (N_9791,N_6007,N_7119);
nor U9792 (N_9792,N_6856,N_7339);
nor U9793 (N_9793,N_8922,N_8553);
nor U9794 (N_9794,N_7190,N_7832);
xnor U9795 (N_9795,N_7675,N_6219);
nor U9796 (N_9796,N_8085,N_7821);
and U9797 (N_9797,N_6751,N_6848);
or U9798 (N_9798,N_7784,N_6815);
nand U9799 (N_9799,N_8842,N_7402);
xnor U9800 (N_9800,N_7071,N_6637);
and U9801 (N_9801,N_8687,N_6649);
and U9802 (N_9802,N_7159,N_8361);
and U9803 (N_9803,N_8632,N_7914);
and U9804 (N_9804,N_7813,N_6728);
or U9805 (N_9805,N_6492,N_8946);
and U9806 (N_9806,N_6054,N_8194);
nand U9807 (N_9807,N_8044,N_6930);
or U9808 (N_9808,N_6987,N_7951);
or U9809 (N_9809,N_6178,N_8542);
or U9810 (N_9810,N_6088,N_7561);
nor U9811 (N_9811,N_6590,N_6328);
nand U9812 (N_9812,N_6174,N_6636);
nor U9813 (N_9813,N_7513,N_6759);
nor U9814 (N_9814,N_8948,N_8052);
nor U9815 (N_9815,N_6340,N_8762);
xor U9816 (N_9816,N_6436,N_7890);
xor U9817 (N_9817,N_8797,N_7199);
and U9818 (N_9818,N_8976,N_6493);
and U9819 (N_9819,N_6056,N_8385);
and U9820 (N_9820,N_7587,N_7599);
nand U9821 (N_9821,N_8185,N_6991);
and U9822 (N_9822,N_8576,N_8878);
or U9823 (N_9823,N_8002,N_7122);
nor U9824 (N_9824,N_8031,N_7862);
nor U9825 (N_9825,N_8146,N_6586);
nor U9826 (N_9826,N_8251,N_8286);
nor U9827 (N_9827,N_7689,N_8096);
nor U9828 (N_9828,N_8081,N_6028);
or U9829 (N_9829,N_8631,N_8997);
or U9830 (N_9830,N_8440,N_6311);
or U9831 (N_9831,N_7417,N_7823);
or U9832 (N_9832,N_8457,N_6452);
nor U9833 (N_9833,N_8195,N_8124);
nor U9834 (N_9834,N_8580,N_7929);
nor U9835 (N_9835,N_6086,N_8253);
nor U9836 (N_9836,N_6184,N_7926);
or U9837 (N_9837,N_8919,N_7193);
nor U9838 (N_9838,N_8500,N_6251);
nand U9839 (N_9839,N_6820,N_8106);
and U9840 (N_9840,N_7448,N_8533);
or U9841 (N_9841,N_8916,N_6221);
or U9842 (N_9842,N_6621,N_6599);
nor U9843 (N_9843,N_6177,N_7324);
or U9844 (N_9844,N_7423,N_8524);
and U9845 (N_9845,N_6651,N_6897);
and U9846 (N_9846,N_8577,N_8788);
nor U9847 (N_9847,N_8733,N_8912);
xnor U9848 (N_9848,N_8342,N_7960);
nor U9849 (N_9849,N_7886,N_7905);
nand U9850 (N_9850,N_6021,N_7871);
nor U9851 (N_9851,N_6652,N_7079);
nand U9852 (N_9852,N_6581,N_6444);
xor U9853 (N_9853,N_6521,N_6115);
nor U9854 (N_9854,N_8217,N_7600);
or U9855 (N_9855,N_7126,N_7766);
and U9856 (N_9856,N_7727,N_7012);
nand U9857 (N_9857,N_6152,N_8917);
nor U9858 (N_9858,N_8158,N_8973);
xnor U9859 (N_9859,N_6963,N_8926);
xnor U9860 (N_9860,N_8226,N_8781);
and U9861 (N_9861,N_8685,N_8538);
and U9862 (N_9862,N_6704,N_6216);
nor U9863 (N_9863,N_7183,N_7373);
nand U9864 (N_9864,N_7472,N_8168);
nand U9865 (N_9865,N_6264,N_6039);
xnor U9866 (N_9866,N_8343,N_7307);
nand U9867 (N_9867,N_8366,N_7712);
xnor U9868 (N_9868,N_7220,N_6306);
or U9869 (N_9869,N_6748,N_8594);
or U9870 (N_9870,N_8975,N_6919);
and U9871 (N_9871,N_7616,N_6777);
nor U9872 (N_9872,N_7780,N_7271);
or U9873 (N_9873,N_8755,N_6364);
or U9874 (N_9874,N_7482,N_6335);
nor U9875 (N_9875,N_8620,N_6180);
xor U9876 (N_9876,N_7621,N_6326);
nor U9877 (N_9877,N_8316,N_7309);
and U9878 (N_9878,N_8282,N_8396);
xor U9879 (N_9879,N_6295,N_8817);
and U9880 (N_9880,N_7413,N_7555);
nand U9881 (N_9881,N_7844,N_7248);
and U9882 (N_9882,N_8472,N_7755);
or U9883 (N_9883,N_8407,N_8082);
nor U9884 (N_9884,N_7580,N_8771);
nor U9885 (N_9885,N_8510,N_8971);
nor U9886 (N_9886,N_6182,N_8435);
and U9887 (N_9887,N_6273,N_8088);
nor U9888 (N_9888,N_8649,N_7125);
or U9889 (N_9889,N_7658,N_6298);
xnor U9890 (N_9890,N_8433,N_7157);
nand U9891 (N_9891,N_8214,N_8438);
or U9892 (N_9892,N_8478,N_7262);
xor U9893 (N_9893,N_6898,N_6980);
and U9894 (N_9894,N_7006,N_8647);
or U9895 (N_9895,N_8938,N_7497);
and U9896 (N_9896,N_6516,N_8201);
and U9897 (N_9897,N_6975,N_8130);
xor U9898 (N_9898,N_8465,N_8032);
or U9899 (N_9899,N_8338,N_7519);
nor U9900 (N_9900,N_8114,N_7665);
xor U9901 (N_9901,N_6104,N_6557);
and U9902 (N_9902,N_6125,N_8064);
nand U9903 (N_9903,N_8140,N_8178);
nor U9904 (N_9904,N_7608,N_7725);
nor U9905 (N_9905,N_8617,N_7747);
and U9906 (N_9906,N_8545,N_7100);
nand U9907 (N_9907,N_8181,N_7781);
and U9908 (N_9908,N_6691,N_8770);
nor U9909 (N_9909,N_7872,N_6237);
nand U9910 (N_9910,N_6688,N_8190);
or U9911 (N_9911,N_6937,N_6706);
xnor U9912 (N_9912,N_8270,N_6345);
or U9913 (N_9913,N_7030,N_7251);
nand U9914 (N_9914,N_8913,N_6377);
and U9915 (N_9915,N_7072,N_7853);
nand U9916 (N_9916,N_6434,N_6646);
nor U9917 (N_9917,N_6502,N_7158);
or U9918 (N_9918,N_6473,N_8949);
and U9919 (N_9919,N_7699,N_8118);
nor U9920 (N_9920,N_8575,N_8015);
and U9921 (N_9921,N_6303,N_7131);
or U9922 (N_9922,N_6194,N_6746);
and U9923 (N_9923,N_6378,N_8859);
or U9924 (N_9924,N_6106,N_7388);
xnor U9925 (N_9925,N_6992,N_8623);
or U9926 (N_9926,N_8318,N_8262);
nor U9927 (N_9927,N_7697,N_8680);
nand U9928 (N_9928,N_7540,N_7794);
nand U9929 (N_9929,N_6217,N_8735);
nor U9930 (N_9930,N_6577,N_8883);
and U9931 (N_9931,N_6981,N_8511);
xor U9932 (N_9932,N_7258,N_7509);
nor U9933 (N_9933,N_6874,N_7790);
xnor U9934 (N_9934,N_7917,N_6322);
nor U9935 (N_9935,N_8568,N_6608);
nand U9936 (N_9936,N_7170,N_8871);
nor U9937 (N_9937,N_6723,N_8821);
xnor U9938 (N_9938,N_7586,N_7805);
nor U9939 (N_9939,N_8406,N_8419);
nor U9940 (N_9940,N_8856,N_6968);
and U9941 (N_9941,N_6485,N_8148);
xnor U9942 (N_9942,N_6098,N_7156);
and U9943 (N_9943,N_8978,N_7743);
and U9944 (N_9944,N_7173,N_8832);
nand U9945 (N_9945,N_6773,N_8030);
xor U9946 (N_9946,N_6465,N_7952);
xor U9947 (N_9947,N_6552,N_7419);
and U9948 (N_9948,N_8470,N_6977);
xnor U9949 (N_9949,N_7762,N_7357);
nand U9950 (N_9950,N_6132,N_8522);
nor U9951 (N_9951,N_7992,N_8714);
nand U9952 (N_9952,N_8404,N_8418);
nand U9953 (N_9953,N_8209,N_6204);
or U9954 (N_9954,N_8650,N_6362);
nand U9955 (N_9955,N_6127,N_6654);
or U9956 (N_9956,N_7518,N_8080);
or U9957 (N_9957,N_7935,N_6220);
nor U9958 (N_9958,N_7715,N_7941);
or U9959 (N_9959,N_7788,N_6727);
xnor U9960 (N_9960,N_6331,N_8100);
and U9961 (N_9961,N_7418,N_6150);
xnor U9962 (N_9962,N_8309,N_7855);
nor U9963 (N_9963,N_8485,N_6966);
and U9964 (N_9964,N_7075,N_6403);
nand U9965 (N_9965,N_6770,N_7106);
xnor U9966 (N_9966,N_6900,N_8591);
or U9967 (N_9967,N_7218,N_7316);
or U9968 (N_9968,N_8016,N_8323);
nor U9969 (N_9969,N_7738,N_8301);
nor U9970 (N_9970,N_8074,N_7843);
nand U9971 (N_9971,N_8989,N_8489);
or U9972 (N_9972,N_8786,N_8780);
and U9973 (N_9973,N_7172,N_6496);
or U9974 (N_9974,N_7529,N_7210);
nor U9975 (N_9975,N_8588,N_8132);
and U9976 (N_9976,N_7137,N_7476);
xnor U9977 (N_9977,N_6764,N_6522);
and U9978 (N_9978,N_8403,N_8962);
xor U9979 (N_9979,N_7904,N_7483);
or U9980 (N_9980,N_8608,N_8220);
nor U9981 (N_9981,N_7302,N_8635);
nand U9982 (N_9982,N_7863,N_8420);
and U9983 (N_9983,N_6999,N_7470);
or U9984 (N_9984,N_7375,N_8929);
nand U9985 (N_9985,N_8038,N_6718);
nand U9986 (N_9986,N_6745,N_6683);
nor U9987 (N_9987,N_8683,N_8072);
nor U9988 (N_9988,N_7551,N_8936);
nor U9989 (N_9989,N_8364,N_8890);
or U9990 (N_9990,N_7505,N_6955);
or U9991 (N_9991,N_8091,N_6316);
nor U9992 (N_9992,N_6788,N_8287);
or U9993 (N_9993,N_6455,N_6901);
nor U9994 (N_9994,N_7305,N_6229);
or U9995 (N_9995,N_6363,N_7517);
or U9996 (N_9996,N_7294,N_7520);
or U9997 (N_9997,N_7189,N_7404);
nand U9998 (N_9998,N_6701,N_7648);
nor U9999 (N_9999,N_6828,N_7303);
and U10000 (N_10000,N_8583,N_7625);
xor U10001 (N_10001,N_8743,N_7678);
nor U10002 (N_10002,N_7534,N_6689);
xnor U10003 (N_10003,N_6806,N_6648);
xor U10004 (N_10004,N_7566,N_6961);
nor U10005 (N_10005,N_6080,N_6369);
xnor U10006 (N_10006,N_8611,N_7014);
nor U10007 (N_10007,N_8621,N_6545);
nor U10008 (N_10008,N_6354,N_8791);
nor U10009 (N_10009,N_6640,N_8567);
xor U10010 (N_10010,N_7657,N_6868);
nand U10011 (N_10011,N_7530,N_7238);
or U10012 (N_10012,N_7361,N_6140);
nor U10013 (N_10013,N_8590,N_8934);
nor U10014 (N_10014,N_8161,N_6188);
or U10015 (N_10015,N_8582,N_7945);
xor U10016 (N_10016,N_8487,N_7525);
nor U10017 (N_10017,N_7536,N_6386);
and U10018 (N_10018,N_7686,N_6747);
nand U10019 (N_10019,N_8848,N_7048);
nand U10020 (N_10020,N_8351,N_6050);
or U10021 (N_10021,N_6677,N_6143);
nand U10022 (N_10022,N_8369,N_6210);
nand U10023 (N_10023,N_7490,N_8573);
and U10024 (N_10024,N_8867,N_6605);
xor U10025 (N_10025,N_8482,N_7624);
nand U10026 (N_10026,N_6291,N_8806);
nor U10027 (N_10027,N_6902,N_8845);
and U10028 (N_10028,N_8352,N_7095);
nand U10029 (N_10029,N_8544,N_6889);
xor U10030 (N_10030,N_6594,N_6000);
nor U10031 (N_10031,N_8171,N_6858);
or U10032 (N_10032,N_7504,N_6375);
nor U10033 (N_10033,N_7801,N_8660);
or U10034 (N_10034,N_7899,N_7411);
nor U10035 (N_10035,N_6175,N_6823);
nand U10036 (N_10036,N_7296,N_8731);
or U10037 (N_10037,N_6641,N_6907);
xor U10038 (N_10038,N_7300,N_6484);
and U10039 (N_10039,N_6936,N_7088);
nand U10040 (N_10040,N_7298,N_7918);
and U10041 (N_10041,N_7108,N_6077);
or U10042 (N_10042,N_6339,N_8004);
nand U10043 (N_10043,N_8508,N_8464);
nand U10044 (N_10044,N_8349,N_8202);
and U10045 (N_10045,N_6478,N_6435);
or U10046 (N_10046,N_8561,N_6477);
xor U10047 (N_10047,N_6196,N_8443);
and U10048 (N_10048,N_6297,N_6971);
nor U10049 (N_10049,N_6814,N_7582);
nor U10050 (N_10050,N_8354,N_7636);
nor U10051 (N_10051,N_6595,N_8230);
nand U10052 (N_10052,N_7087,N_8818);
nor U10053 (N_10053,N_7507,N_6756);
nor U10054 (N_10054,N_8143,N_8721);
xnor U10055 (N_10055,N_6798,N_8437);
and U10056 (N_10056,N_6766,N_6692);
and U10057 (N_10057,N_7541,N_7257);
or U10058 (N_10058,N_6864,N_8889);
and U10059 (N_10059,N_7177,N_7702);
xor U10060 (N_10060,N_6130,N_6855);
xnor U10061 (N_10061,N_7468,N_7865);
nor U10062 (N_10062,N_6203,N_6010);
and U10063 (N_10063,N_6313,N_7887);
or U10064 (N_10064,N_8242,N_6330);
and U10065 (N_10065,N_8259,N_7463);
xor U10066 (N_10066,N_6206,N_7553);
nand U10067 (N_10067,N_6195,N_8761);
nand U10068 (N_10068,N_8707,N_7436);
and U10069 (N_10069,N_7512,N_7549);
xnor U10070 (N_10070,N_8796,N_6994);
or U10071 (N_10071,N_8748,N_8704);
nand U10072 (N_10072,N_7718,N_6905);
xor U10073 (N_10073,N_6852,N_6268);
or U10074 (N_10074,N_8521,N_7334);
or U10075 (N_10075,N_6744,N_7182);
or U10076 (N_10076,N_7363,N_6721);
and U10077 (N_10077,N_7427,N_7018);
nor U10078 (N_10078,N_8864,N_6906);
nand U10079 (N_10079,N_8445,N_7261);
nor U10080 (N_10080,N_8045,N_6159);
xnor U10081 (N_10081,N_6267,N_7399);
and U10082 (N_10082,N_8384,N_6512);
nand U10083 (N_10083,N_6803,N_7297);
nand U10084 (N_10084,N_6228,N_8335);
and U10085 (N_10085,N_6670,N_7545);
xor U10086 (N_10086,N_7692,N_6246);
or U10087 (N_10087,N_8835,N_6607);
nor U10088 (N_10088,N_7696,N_7078);
or U10089 (N_10089,N_6833,N_8787);
or U10090 (N_10090,N_7906,N_6510);
or U10091 (N_10091,N_7835,N_6278);
and U10092 (N_10092,N_8493,N_6680);
nor U10093 (N_10093,N_8880,N_7138);
nor U10094 (N_10094,N_8391,N_6631);
xor U10095 (N_10095,N_7969,N_7850);
nor U10096 (N_10096,N_8902,N_8592);
nand U10097 (N_10097,N_6886,N_8626);
or U10098 (N_10098,N_7081,N_7186);
xnor U10099 (N_10099,N_6081,N_8455);
or U10100 (N_10100,N_8039,N_7181);
and U10101 (N_10101,N_8483,N_6324);
xnor U10102 (N_10102,N_6519,N_8987);
or U10103 (N_10103,N_7323,N_7638);
xnor U10104 (N_10104,N_8637,N_8079);
xnor U10105 (N_10105,N_7259,N_8504);
nand U10106 (N_10106,N_7386,N_8950);
and U10107 (N_10107,N_6300,N_7649);
nand U10108 (N_10108,N_8051,N_7164);
nand U10109 (N_10109,N_6109,N_6405);
xnor U10110 (N_10110,N_7217,N_8563);
and U10111 (N_10111,N_7234,N_8431);
nand U10112 (N_10112,N_6082,N_7456);
or U10113 (N_10113,N_8712,N_6663);
and U10114 (N_10114,N_7010,N_6170);
and U10115 (N_10115,N_7293,N_8166);
nand U10116 (N_10116,N_6942,N_8519);
nand U10117 (N_10117,N_8766,N_7981);
and U10118 (N_10118,N_7086,N_6315);
nor U10119 (N_10119,N_6225,N_7376);
or U10120 (N_10120,N_6281,N_8725);
nand U10121 (N_10121,N_7401,N_6169);
xor U10122 (N_10122,N_7759,N_8571);
and U10123 (N_10123,N_6164,N_8837);
nor U10124 (N_10124,N_7936,N_7543);
nand U10125 (N_10125,N_8173,N_8833);
xor U10126 (N_10126,N_8752,N_6276);
nand U10127 (N_10127,N_8249,N_7022);
or U10128 (N_10128,N_7360,N_8981);
and U10129 (N_10129,N_7911,N_8083);
xnor U10130 (N_10130,N_6073,N_8006);
xnor U10131 (N_10131,N_8742,N_8763);
or U10132 (N_10132,N_8782,N_8947);
xor U10133 (N_10133,N_7321,N_7121);
nand U10134 (N_10134,N_7355,N_6882);
xnor U10135 (N_10135,N_7492,N_7524);
or U10136 (N_10136,N_8497,N_8104);
or U10137 (N_10137,N_6927,N_6914);
xor U10138 (N_10138,N_7110,N_6832);
or U10139 (N_10139,N_7066,N_8910);
nor U10140 (N_10140,N_7113,N_6752);
nor U10141 (N_10141,N_6153,N_7474);
nand U10142 (N_10142,N_7817,N_6836);
nand U10143 (N_10143,N_6239,N_8312);
or U10144 (N_10144,N_7554,N_7387);
or U10145 (N_10145,N_8398,N_6327);
or U10146 (N_10146,N_8110,N_7571);
nor U10147 (N_10147,N_6878,N_8887);
nand U10148 (N_10148,N_7514,N_8098);
nand U10149 (N_10149,N_8614,N_6964);
or U10150 (N_10150,N_8353,N_6653);
nor U10151 (N_10151,N_8531,N_6048);
nand U10152 (N_10152,N_8059,N_8970);
and U10153 (N_10153,N_8498,N_6517);
and U10154 (N_10154,N_8730,N_6712);
or U10155 (N_10155,N_6165,N_6548);
nor U10156 (N_10156,N_7260,N_7889);
and U10157 (N_10157,N_7054,N_7051);
or U10158 (N_10158,N_8891,N_8162);
xnor U10159 (N_10159,N_7795,N_6730);
nor U10160 (N_10160,N_6566,N_6116);
nand U10161 (N_10161,N_7864,N_8164);
nand U10162 (N_10162,N_6133,N_7135);
nor U10163 (N_10163,N_7793,N_7565);
and U10164 (N_10164,N_7948,N_6835);
or U10165 (N_10165,N_6600,N_7695);
nor U10166 (N_10166,N_6044,N_6693);
nor U10167 (N_10167,N_6831,N_8846);
nand U10168 (N_10168,N_6047,N_7975);
and U10169 (N_10169,N_7511,N_6034);
xnor U10170 (N_10170,N_8236,N_6402);
or U10171 (N_10171,N_7442,N_6639);
or U10172 (N_10172,N_7341,N_8534);
or U10173 (N_10173,N_8340,N_7655);
and U10174 (N_10174,N_7652,N_6483);
or U10175 (N_10175,N_6283,N_7569);
and U10176 (N_10176,N_8793,N_6454);
nand U10177 (N_10177,N_8036,N_7597);
nand U10178 (N_10178,N_7983,N_8541);
and U10179 (N_10179,N_7481,N_7532);
and U10180 (N_10180,N_7607,N_8448);
nand U10181 (N_10181,N_7469,N_8271);
or U10182 (N_10182,N_8336,N_6348);
nand U10183 (N_10183,N_7868,N_8773);
or U10184 (N_10184,N_8951,N_6698);
nand U10185 (N_10185,N_8990,N_7011);
or U10186 (N_10186,N_7820,N_6272);
or U10187 (N_10187,N_7620,N_6547);
or U10188 (N_10188,N_8456,N_7577);
xor U10189 (N_10189,N_8954,N_8429);
and U10190 (N_10190,N_8915,N_8054);
and U10191 (N_10191,N_6742,N_7995);
nor U10192 (N_10192,N_6544,N_8925);
nor U10193 (N_10193,N_7101,N_7477);
nor U10194 (N_10194,N_7963,N_8373);
nor U10195 (N_10195,N_8449,N_7841);
nand U10196 (N_10196,N_8341,N_7499);
nand U10197 (N_10197,N_8943,N_6235);
nor U10198 (N_10198,N_6020,N_6388);
nand U10199 (N_10199,N_8515,N_7506);
nand U10200 (N_10200,N_7068,N_8248);
and U10201 (N_10201,N_7028,N_8759);
xor U10202 (N_10202,N_6489,N_6837);
nor U10203 (N_10203,N_8562,N_8276);
and U10204 (N_10204,N_8359,N_6617);
nand U10205 (N_10205,N_8653,N_6413);
nor U10206 (N_10206,N_6487,N_6567);
nor U10207 (N_10207,N_6940,N_6076);
nor U10208 (N_10208,N_7733,N_7236);
or U10209 (N_10209,N_8068,N_6263);
nor U10210 (N_10210,N_7446,N_6200);
or U10211 (N_10211,N_8927,N_6624);
and U10212 (N_10212,N_8826,N_7192);
nor U10213 (N_10213,N_7049,N_6892);
and U10214 (N_10214,N_7787,N_8854);
xnor U10215 (N_10215,N_8128,N_8783);
xor U10216 (N_10216,N_8473,N_8094);
and U10217 (N_10217,N_6119,N_7606);
nand U10218 (N_10218,N_7557,N_6847);
nor U10219 (N_10219,N_7654,N_8778);
nand U10220 (N_10220,N_7025,N_7276);
or U10221 (N_10221,N_7379,N_7730);
nor U10222 (N_10222,N_6559,N_7503);
nand U10223 (N_10223,N_8738,N_6990);
and U10224 (N_10224,N_8365,N_7713);
or U10225 (N_10225,N_8274,N_8441);
or U10226 (N_10226,N_8256,N_8310);
nand U10227 (N_10227,N_7077,N_8356);
nand U10228 (N_10228,N_7188,N_7346);
nand U10229 (N_10229,N_8774,N_6793);
and U10230 (N_10230,N_7523,N_7708);
or U10231 (N_10231,N_7338,N_6530);
or U10232 (N_10232,N_6504,N_6381);
and U10233 (N_10233,N_7426,N_8720);
and U10234 (N_10234,N_8681,N_8159);
nand U10235 (N_10235,N_7897,N_6256);
xnor U10236 (N_10236,N_6647,N_7976);
xnor U10237 (N_10237,N_7225,N_6870);
nor U10238 (N_10238,N_8066,N_6561);
nor U10239 (N_10239,N_6565,N_8540);
nand U10240 (N_10240,N_6623,N_8327);
xnor U10241 (N_10241,N_8252,N_6908);
nor U10242 (N_10242,N_7348,N_7283);
or U10243 (N_10243,N_8332,N_6155);
xnor U10244 (N_10244,N_8200,N_8876);
xor U10245 (N_10245,N_6112,N_7083);
nand U10246 (N_10246,N_7480,N_7461);
or U10247 (N_10247,N_6778,N_6209);
nor U10248 (N_10248,N_7726,N_6584);
nand U10249 (N_10249,N_7447,N_7299);
nand U10250 (N_10250,N_6359,N_6063);
nor U10251 (N_10251,N_7612,N_7045);
nand U10252 (N_10252,N_8673,N_6749);
nand U10253 (N_10253,N_7882,N_6394);
xnor U10254 (N_10254,N_6146,N_6916);
or U10255 (N_10255,N_7891,N_7288);
or U10256 (N_10256,N_8390,N_7120);
and U10257 (N_10257,N_7282,N_8741);
xor U10258 (N_10258,N_7241,N_6418);
xor U10259 (N_10259,N_8263,N_8496);
nor U10260 (N_10260,N_7219,N_8967);
nand U10261 (N_10261,N_8346,N_7286);
xnor U10262 (N_10262,N_7063,N_7368);
and U10263 (N_10263,N_7161,N_8492);
or U10264 (N_10264,N_7860,N_7664);
nor U10265 (N_10265,N_8121,N_8093);
or U10266 (N_10266,N_6604,N_7187);
and U10267 (N_10267,N_6757,N_6151);
nand U10268 (N_10268,N_6817,N_6576);
xor U10269 (N_10269,N_6609,N_7867);
or U10270 (N_10270,N_7253,N_6445);
or U10271 (N_10271,N_6618,N_6479);
xnor U10272 (N_10272,N_6926,N_7701);
nor U10273 (N_10273,N_6627,N_6863);
or U10274 (N_10274,N_7393,N_7369);
xnor U10275 (N_10275,N_6353,N_6662);
xor U10276 (N_10276,N_8027,N_8011);
nor U10277 (N_10277,N_8654,N_7112);
or U10278 (N_10278,N_8689,N_8896);
and U10279 (N_10279,N_6396,N_6079);
nand U10280 (N_10280,N_8675,N_7089);
and U10281 (N_10281,N_7280,N_7706);
or U10282 (N_10282,N_8601,N_6078);
xnor U10283 (N_10283,N_8703,N_6105);
or U10284 (N_10284,N_8157,N_7642);
and U10285 (N_10285,N_8810,N_8392);
nor U10286 (N_10286,N_8377,N_8911);
or U10287 (N_10287,N_7997,N_8371);
nand U10288 (N_10288,N_7798,N_6767);
xnor U10289 (N_10289,N_6156,N_6168);
and U10290 (N_10290,N_6769,N_7224);
or U10291 (N_10291,N_6781,N_6282);
nand U10292 (N_10292,N_6214,N_6570);
nand U10293 (N_10293,N_8550,N_7912);
nand U10294 (N_10294,N_8937,N_6374);
and U10295 (N_10295,N_6606,N_8428);
nor U10296 (N_10296,N_6365,N_6910);
nand U10297 (N_10297,N_6783,N_8266);
nor U10298 (N_10298,N_6380,N_7842);
nor U10299 (N_10299,N_6672,N_7467);
nor U10300 (N_10300,N_7527,N_6716);
or U10301 (N_10301,N_7410,N_7148);
and U10302 (N_10302,N_8474,N_7651);
nor U10303 (N_10303,N_6058,N_6542);
and U10304 (N_10304,N_8387,N_7966);
nor U10305 (N_10305,N_6705,N_7609);
nor U10306 (N_10306,N_8628,N_6614);
or U10307 (N_10307,N_8314,N_8476);
nand U10308 (N_10308,N_8246,N_7746);
xnor U10309 (N_10309,N_6172,N_8150);
nand U10310 (N_10310,N_8203,N_8269);
nand U10311 (N_10311,N_6524,N_8850);
xnor U10312 (N_10312,N_7315,N_8326);
or U10313 (N_10313,N_6408,N_6558);
and U10314 (N_10314,N_7979,N_7547);
nand U10315 (N_10315,N_8042,N_8991);
nand U10316 (N_10316,N_7287,N_7589);
xnor U10317 (N_10317,N_8484,N_8380);
nor U10318 (N_10318,N_7866,N_7595);
nand U10319 (N_10319,N_8291,N_7771);
or U10320 (N_10320,N_6630,N_7563);
nor U10321 (N_10321,N_7659,N_8021);
and U10322 (N_10322,N_6259,N_8086);
or U10323 (N_10323,N_6158,N_8479);
xor U10324 (N_10324,N_8460,N_7487);
nor U10325 (N_10325,N_8499,N_8109);
or U10326 (N_10326,N_8935,N_8784);
xor U10327 (N_10327,N_6733,N_7458);
nor U10328 (N_10328,N_8374,N_7656);
and U10329 (N_10329,N_8076,N_8239);
and U10330 (N_10330,N_8144,N_6546);
nor U10331 (N_10331,N_6171,N_6040);
nand U10332 (N_10332,N_8026,N_7732);
nand U10333 (N_10333,N_6108,N_8918);
nor U10334 (N_10334,N_8897,N_7214);
or U10335 (N_10335,N_6323,N_8469);
nand U10336 (N_10336,N_8308,N_6791);
or U10337 (N_10337,N_8300,N_7683);
nor U10338 (N_10338,N_8176,N_6877);
and U10339 (N_10339,N_7318,N_8097);
or U10340 (N_10340,N_8812,N_8425);
nor U10341 (N_10341,N_6660,N_8503);
nor U10342 (N_10342,N_7856,N_7971);
and U10343 (N_10343,N_6962,N_6066);
xnor U10344 (N_10344,N_8772,N_8666);
nor U10345 (N_10345,N_7123,N_6702);
nand U10346 (N_10346,N_8153,N_8723);
or U10347 (N_10347,N_6880,N_6286);
nor U10348 (N_10348,N_8661,N_6804);
nor U10349 (N_10349,N_6497,N_6468);
or U10350 (N_10350,N_6934,N_8113);
xor U10351 (N_10351,N_8682,N_7450);
or U10352 (N_10352,N_6023,N_8175);
or U10353 (N_10353,N_6635,N_6017);
xor U10354 (N_10354,N_8227,N_8405);
and U10355 (N_10355,N_7223,N_7152);
nor U10356 (N_10356,N_7412,N_8516);
and U10357 (N_10357,N_7032,N_8427);
or U10358 (N_10358,N_7754,N_8700);
nor U10359 (N_10359,N_7184,N_6495);
nand U10360 (N_10360,N_6708,N_6042);
xor U10361 (N_10361,N_6043,N_8564);
and U10362 (N_10362,N_8288,N_8134);
nand U10363 (N_10363,N_8565,N_7709);
nor U10364 (N_10364,N_8182,N_7627);
nor U10365 (N_10365,N_7923,N_7567);
xnor U10366 (N_10366,N_6065,N_8228);
nand U10367 (N_10367,N_7434,N_7994);
or U10368 (N_10368,N_7854,N_8506);
xnor U10369 (N_10369,N_7356,N_8023);
and U10370 (N_10370,N_6166,N_6011);
nand U10371 (N_10371,N_7452,N_8417);
xnor U10372 (N_10372,N_8802,N_7269);
xnor U10373 (N_10373,N_8952,N_7201);
nor U10374 (N_10374,N_7055,N_6928);
nand U10375 (N_10375,N_6950,N_6508);
and U10376 (N_10376,N_6871,N_6067);
and U10377 (N_10377,N_6161,N_6442);
and U10378 (N_10378,N_7494,N_8986);
and U10379 (N_10379,N_7493,N_6787);
nor U10380 (N_10380,N_6665,N_7646);
xnor U10381 (N_10381,N_6843,N_7900);
and U10382 (N_10382,N_8219,N_7056);
or U10383 (N_10383,N_7284,N_6309);
nand U10384 (N_10384,N_8412,N_6289);
or U10385 (N_10385,N_7775,N_7635);
nand U10386 (N_10386,N_7698,N_7228);
or U10387 (N_10387,N_8830,N_7986);
xor U10388 (N_10388,N_7931,N_7243);
nor U10389 (N_10389,N_7987,N_7521);
nand U10390 (N_10390,N_8529,N_6016);
nor U10391 (N_10391,N_7585,N_7365);
or U10392 (N_10392,N_8388,N_8368);
nor U10393 (N_10393,N_7024,N_7591);
and U10394 (N_10394,N_8320,N_6265);
and U10395 (N_10395,N_7289,N_8980);
nand U10396 (N_10396,N_7454,N_8994);
nand U10397 (N_10397,N_8060,N_7364);
nand U10398 (N_10398,N_6385,N_7548);
xnor U10399 (N_10399,N_6351,N_7215);
xnor U10400 (N_10400,N_8423,N_8421);
nor U10401 (N_10401,N_7053,N_6357);
or U10402 (N_10402,N_7501,N_6996);
or U10403 (N_10403,N_8048,N_6731);
xnor U10404 (N_10404,N_6426,N_7603);
nand U10405 (N_10405,N_8255,N_6634);
or U10406 (N_10406,N_8776,N_8581);
or U10407 (N_10407,N_7946,N_8753);
nor U10408 (N_10408,N_8982,N_7471);
or U10409 (N_10409,N_8528,N_6387);
and U10410 (N_10410,N_6860,N_8179);
and U10411 (N_10411,N_7097,N_7067);
or U10412 (N_10412,N_7301,N_6269);
xor U10413 (N_10413,N_6356,N_6715);
and U10414 (N_10414,N_7528,N_8888);
nand U10415 (N_10415,N_7409,N_7873);
nand U10416 (N_10416,N_8197,N_7875);
nand U10417 (N_10417,N_7633,N_7377);
nand U10418 (N_10418,N_7980,N_8838);
nor U10419 (N_10419,N_8638,N_7691);
nor U10420 (N_10420,N_7352,N_6250);
nor U10421 (N_10421,N_7782,N_7752);
xor U10422 (N_10422,N_6821,N_8662);
or U10423 (N_10423,N_8695,N_7485);
nand U10424 (N_10424,N_7909,N_7153);
and U10425 (N_10425,N_6941,N_6242);
and U10426 (N_10426,N_7209,N_7778);
xnor U10427 (N_10427,N_7180,N_7350);
or U10428 (N_10428,N_8706,N_8213);
xnor U10429 (N_10429,N_8942,N_7829);
nor U10430 (N_10430,N_7233,N_7956);
nand U10431 (N_10431,N_7739,N_6822);
xor U10432 (N_10432,N_8331,N_8984);
or U10433 (N_10433,N_8604,N_7990);
or U10434 (N_10434,N_6876,N_6012);
nor U10435 (N_10435,N_8825,N_8322);
and U10436 (N_10436,N_7742,N_8847);
and U10437 (N_10437,N_8670,N_7281);
nor U10438 (N_10438,N_6935,N_6193);
nor U10439 (N_10439,N_8998,N_6743);
xor U10440 (N_10440,N_6481,N_7337);
nor U10441 (N_10441,N_6025,N_7403);
nor U10442 (N_10442,N_7050,N_6245);
and U10443 (N_10443,N_8018,N_6032);
nand U10444 (N_10444,N_7275,N_6051);
nor U10445 (N_10445,N_6083,N_6944);
and U10446 (N_10446,N_6726,N_8599);
or U10447 (N_10447,N_7094,N_8698);
and U10448 (N_10448,N_7200,N_6838);
or U10449 (N_10449,N_6912,N_6763);
xnor U10450 (N_10450,N_6846,N_8345);
nand U10451 (N_10451,N_8640,N_8616);
and U10452 (N_10452,N_7278,N_6218);
and U10453 (N_10453,N_7464,N_8881);
or U10454 (N_10454,N_7230,N_8199);
xor U10455 (N_10455,N_6974,N_7004);
and U10456 (N_10456,N_7058,N_7930);
nor U10457 (N_10457,N_6840,N_8820);
xnor U10458 (N_10458,N_8260,N_8245);
nor U10459 (N_10459,N_6072,N_7486);
or U10460 (N_10460,N_6982,N_7406);
nor U10461 (N_10461,N_7593,N_8719);
xor U10462 (N_10462,N_8865,N_6842);
xor U10463 (N_10463,N_7082,N_6211);
and U10464 (N_10464,N_6972,N_7827);
xor U10465 (N_10465,N_6293,N_8520);
nand U10466 (N_10466,N_7445,N_8205);
nand U10467 (N_10467,N_6427,N_8728);
and U10468 (N_10468,N_8933,N_8409);
and U10469 (N_10469,N_8597,N_6136);
and U10470 (N_10470,N_7750,N_7630);
nor U10471 (N_10471,N_6494,N_7632);
and U10472 (N_10472,N_6234,N_8160);
nor U10473 (N_10473,N_8586,N_7700);
xnor U10474 (N_10474,N_8560,N_7105);
nor U10475 (N_10475,N_6978,N_7907);
nor U10476 (N_10476,N_8705,N_7703);
or U10477 (N_10477,N_7874,N_6535);
nor U10478 (N_10478,N_8834,N_7803);
and U10479 (N_10479,N_8569,N_7264);
nor U10480 (N_10480,N_7292,N_8513);
xnor U10481 (N_10481,N_8613,N_7231);
xor U10482 (N_10482,N_7661,N_8959);
nor U10483 (N_10483,N_8444,N_7029);
nor U10484 (N_10484,N_8238,N_8206);
nand U10485 (N_10485,N_8129,N_8491);
xor U10486 (N_10486,N_7019,N_6024);
and U10487 (N_10487,N_6416,N_7155);
xor U10488 (N_10488,N_7196,N_6794);
or U10489 (N_10489,N_6615,N_8198);
xor U10490 (N_10490,N_7397,N_7003);
nor U10491 (N_10491,N_7758,N_7059);
nor U10492 (N_10492,N_7559,N_6107);
or U10493 (N_10493,N_7489,N_7479);
and U10494 (N_10494,N_6103,N_6579);
nand U10495 (N_10495,N_7861,N_7065);
xnor U10496 (N_10496,N_7982,N_7894);
nor U10497 (N_10497,N_8305,N_8267);
or U10498 (N_10498,N_7197,N_7139);
nor U10499 (N_10499,N_7870,N_6280);
and U10500 (N_10500,N_7805,N_6285);
nor U10501 (N_10501,N_7075,N_7751);
nor U10502 (N_10502,N_7896,N_7952);
nor U10503 (N_10503,N_6261,N_7552);
nand U10504 (N_10504,N_7548,N_7549);
nor U10505 (N_10505,N_7930,N_6743);
xor U10506 (N_10506,N_7528,N_8777);
nor U10507 (N_10507,N_6278,N_7093);
and U10508 (N_10508,N_6376,N_6176);
or U10509 (N_10509,N_6495,N_6498);
or U10510 (N_10510,N_6865,N_8464);
xnor U10511 (N_10511,N_8493,N_8602);
nor U10512 (N_10512,N_7443,N_8562);
nor U10513 (N_10513,N_6723,N_6200);
or U10514 (N_10514,N_6093,N_6237);
xnor U10515 (N_10515,N_7968,N_7908);
and U10516 (N_10516,N_7826,N_6912);
and U10517 (N_10517,N_6375,N_6023);
and U10518 (N_10518,N_6959,N_8976);
xor U10519 (N_10519,N_6291,N_7422);
nand U10520 (N_10520,N_6822,N_7059);
xnor U10521 (N_10521,N_7740,N_7793);
or U10522 (N_10522,N_6122,N_6620);
nand U10523 (N_10523,N_6771,N_7977);
nand U10524 (N_10524,N_7295,N_8673);
nor U10525 (N_10525,N_8692,N_8788);
nand U10526 (N_10526,N_6953,N_7488);
xnor U10527 (N_10527,N_8147,N_8546);
and U10528 (N_10528,N_7942,N_6616);
nand U10529 (N_10529,N_8416,N_8069);
or U10530 (N_10530,N_6332,N_6683);
and U10531 (N_10531,N_6304,N_8660);
xor U10532 (N_10532,N_6725,N_6921);
nor U10533 (N_10533,N_6980,N_6242);
and U10534 (N_10534,N_8031,N_8859);
nand U10535 (N_10535,N_7269,N_6169);
or U10536 (N_10536,N_8681,N_6954);
or U10537 (N_10537,N_8829,N_8741);
or U10538 (N_10538,N_7894,N_7530);
and U10539 (N_10539,N_6852,N_7454);
nor U10540 (N_10540,N_8041,N_6387);
nor U10541 (N_10541,N_7930,N_8550);
and U10542 (N_10542,N_6771,N_6680);
nand U10543 (N_10543,N_8057,N_8118);
nand U10544 (N_10544,N_8567,N_8174);
and U10545 (N_10545,N_6026,N_8717);
nand U10546 (N_10546,N_6909,N_7721);
and U10547 (N_10547,N_8277,N_8457);
nor U10548 (N_10548,N_7201,N_8117);
nor U10549 (N_10549,N_6307,N_6002);
xnor U10550 (N_10550,N_6776,N_8847);
or U10551 (N_10551,N_8459,N_8194);
xor U10552 (N_10552,N_7268,N_8660);
nor U10553 (N_10553,N_8487,N_8355);
or U10554 (N_10554,N_6778,N_8375);
xnor U10555 (N_10555,N_7751,N_6588);
nor U10556 (N_10556,N_8416,N_6643);
or U10557 (N_10557,N_7485,N_7995);
xnor U10558 (N_10558,N_7453,N_8336);
or U10559 (N_10559,N_7474,N_7893);
nand U10560 (N_10560,N_8395,N_8390);
nand U10561 (N_10561,N_7658,N_8899);
nand U10562 (N_10562,N_8716,N_6242);
nor U10563 (N_10563,N_6522,N_8132);
and U10564 (N_10564,N_6282,N_6053);
nand U10565 (N_10565,N_7002,N_7401);
nor U10566 (N_10566,N_6320,N_7530);
or U10567 (N_10567,N_6936,N_6226);
or U10568 (N_10568,N_8388,N_6877);
xnor U10569 (N_10569,N_6374,N_7977);
nor U10570 (N_10570,N_8442,N_8155);
or U10571 (N_10571,N_6259,N_7047);
nor U10572 (N_10572,N_7428,N_8721);
and U10573 (N_10573,N_8666,N_8618);
and U10574 (N_10574,N_6717,N_7447);
or U10575 (N_10575,N_7785,N_8504);
nor U10576 (N_10576,N_6406,N_8274);
or U10577 (N_10577,N_6161,N_6883);
nor U10578 (N_10578,N_7593,N_7047);
nor U10579 (N_10579,N_8585,N_7829);
xor U10580 (N_10580,N_6859,N_8133);
and U10581 (N_10581,N_8153,N_7906);
nand U10582 (N_10582,N_7853,N_7969);
or U10583 (N_10583,N_6624,N_6460);
and U10584 (N_10584,N_8431,N_8333);
xnor U10585 (N_10585,N_8243,N_7589);
or U10586 (N_10586,N_8770,N_7344);
and U10587 (N_10587,N_6999,N_8862);
nand U10588 (N_10588,N_8937,N_7670);
and U10589 (N_10589,N_7024,N_7302);
and U10590 (N_10590,N_6472,N_8832);
xor U10591 (N_10591,N_7684,N_6170);
and U10592 (N_10592,N_6108,N_7768);
and U10593 (N_10593,N_7273,N_8847);
nand U10594 (N_10594,N_8724,N_7865);
and U10595 (N_10595,N_7630,N_7151);
xor U10596 (N_10596,N_6055,N_8484);
nand U10597 (N_10597,N_6455,N_7984);
or U10598 (N_10598,N_6281,N_7281);
or U10599 (N_10599,N_7312,N_8449);
xnor U10600 (N_10600,N_8602,N_6354);
or U10601 (N_10601,N_7296,N_8822);
and U10602 (N_10602,N_8069,N_8099);
xor U10603 (N_10603,N_6794,N_8521);
and U10604 (N_10604,N_8170,N_7290);
or U10605 (N_10605,N_6786,N_6266);
and U10606 (N_10606,N_8138,N_7381);
xnor U10607 (N_10607,N_6886,N_7611);
nor U10608 (N_10608,N_7799,N_8268);
nand U10609 (N_10609,N_6566,N_7186);
xor U10610 (N_10610,N_7163,N_8813);
nand U10611 (N_10611,N_6498,N_8976);
or U10612 (N_10612,N_7731,N_8886);
nand U10613 (N_10613,N_6825,N_7475);
or U10614 (N_10614,N_6174,N_8992);
or U10615 (N_10615,N_8151,N_8080);
xnor U10616 (N_10616,N_8641,N_7555);
nand U10617 (N_10617,N_6912,N_6645);
nor U10618 (N_10618,N_8726,N_7402);
xnor U10619 (N_10619,N_7275,N_8469);
nand U10620 (N_10620,N_8886,N_7851);
xnor U10621 (N_10621,N_6948,N_7577);
nand U10622 (N_10622,N_6281,N_7062);
and U10623 (N_10623,N_6818,N_6155);
xor U10624 (N_10624,N_8846,N_8913);
nor U10625 (N_10625,N_8687,N_7743);
nand U10626 (N_10626,N_7910,N_7257);
and U10627 (N_10627,N_7081,N_8974);
xor U10628 (N_10628,N_7584,N_7316);
xor U10629 (N_10629,N_8458,N_7462);
or U10630 (N_10630,N_7872,N_7330);
xnor U10631 (N_10631,N_8730,N_7381);
xnor U10632 (N_10632,N_7199,N_8281);
xor U10633 (N_10633,N_7520,N_8769);
or U10634 (N_10634,N_8565,N_7814);
xnor U10635 (N_10635,N_8794,N_6505);
xor U10636 (N_10636,N_7531,N_6055);
nor U10637 (N_10637,N_7493,N_8342);
xnor U10638 (N_10638,N_8490,N_7017);
or U10639 (N_10639,N_8249,N_8171);
and U10640 (N_10640,N_7226,N_6730);
or U10641 (N_10641,N_6486,N_6209);
nand U10642 (N_10642,N_6286,N_7156);
or U10643 (N_10643,N_7816,N_7760);
and U10644 (N_10644,N_7933,N_7663);
or U10645 (N_10645,N_8829,N_8695);
nand U10646 (N_10646,N_7643,N_8616);
nor U10647 (N_10647,N_6147,N_7040);
or U10648 (N_10648,N_6425,N_8955);
and U10649 (N_10649,N_6357,N_8219);
and U10650 (N_10650,N_6044,N_7688);
and U10651 (N_10651,N_8350,N_6076);
or U10652 (N_10652,N_6781,N_6530);
and U10653 (N_10653,N_8644,N_8391);
nand U10654 (N_10654,N_8979,N_8940);
xnor U10655 (N_10655,N_7339,N_6185);
xnor U10656 (N_10656,N_8599,N_6232);
nand U10657 (N_10657,N_7082,N_7877);
or U10658 (N_10658,N_6397,N_8152);
nand U10659 (N_10659,N_6220,N_8205);
or U10660 (N_10660,N_7922,N_7321);
xnor U10661 (N_10661,N_7297,N_8833);
and U10662 (N_10662,N_7961,N_7889);
or U10663 (N_10663,N_8264,N_8717);
nor U10664 (N_10664,N_7163,N_6886);
nand U10665 (N_10665,N_7501,N_8112);
xnor U10666 (N_10666,N_7326,N_8561);
nand U10667 (N_10667,N_7870,N_8824);
xor U10668 (N_10668,N_7649,N_8179);
or U10669 (N_10669,N_7426,N_7862);
nand U10670 (N_10670,N_8411,N_8469);
nor U10671 (N_10671,N_6980,N_6642);
xnor U10672 (N_10672,N_8839,N_7373);
nand U10673 (N_10673,N_6903,N_8785);
or U10674 (N_10674,N_6935,N_8393);
and U10675 (N_10675,N_8828,N_6441);
or U10676 (N_10676,N_6560,N_7202);
xor U10677 (N_10677,N_8783,N_8403);
nand U10678 (N_10678,N_6753,N_7909);
nand U10679 (N_10679,N_7333,N_8698);
xor U10680 (N_10680,N_8197,N_6025);
nor U10681 (N_10681,N_6695,N_8608);
nor U10682 (N_10682,N_8625,N_6018);
and U10683 (N_10683,N_7961,N_6360);
and U10684 (N_10684,N_7370,N_8372);
or U10685 (N_10685,N_8449,N_7843);
or U10686 (N_10686,N_6621,N_8195);
xnor U10687 (N_10687,N_8602,N_6535);
xor U10688 (N_10688,N_7975,N_6393);
nand U10689 (N_10689,N_6765,N_8855);
nand U10690 (N_10690,N_7143,N_7598);
nand U10691 (N_10691,N_6777,N_7436);
nand U10692 (N_10692,N_8316,N_8984);
nand U10693 (N_10693,N_6248,N_7100);
and U10694 (N_10694,N_8775,N_6789);
nand U10695 (N_10695,N_6721,N_8298);
and U10696 (N_10696,N_8935,N_6495);
or U10697 (N_10697,N_6612,N_7690);
nor U10698 (N_10698,N_7002,N_6124);
and U10699 (N_10699,N_7093,N_6480);
nand U10700 (N_10700,N_8360,N_6676);
nor U10701 (N_10701,N_6954,N_6117);
and U10702 (N_10702,N_8444,N_8785);
nor U10703 (N_10703,N_8257,N_7950);
nor U10704 (N_10704,N_6136,N_6297);
nand U10705 (N_10705,N_7935,N_6147);
nor U10706 (N_10706,N_8118,N_7705);
and U10707 (N_10707,N_8752,N_7725);
nand U10708 (N_10708,N_8867,N_8876);
nor U10709 (N_10709,N_8881,N_8457);
xnor U10710 (N_10710,N_7474,N_8679);
nor U10711 (N_10711,N_8803,N_8035);
or U10712 (N_10712,N_8907,N_8722);
nor U10713 (N_10713,N_8357,N_7051);
xnor U10714 (N_10714,N_6390,N_7494);
and U10715 (N_10715,N_8914,N_6002);
or U10716 (N_10716,N_7401,N_6931);
xnor U10717 (N_10717,N_6923,N_6548);
nor U10718 (N_10718,N_8673,N_7250);
xnor U10719 (N_10719,N_8894,N_7025);
nor U10720 (N_10720,N_8899,N_8257);
and U10721 (N_10721,N_8059,N_7422);
or U10722 (N_10722,N_7131,N_6667);
or U10723 (N_10723,N_6192,N_8587);
nor U10724 (N_10724,N_8296,N_7067);
xor U10725 (N_10725,N_6105,N_6402);
nand U10726 (N_10726,N_6911,N_6297);
and U10727 (N_10727,N_6970,N_8544);
or U10728 (N_10728,N_8021,N_6269);
xor U10729 (N_10729,N_6363,N_6674);
xnor U10730 (N_10730,N_8183,N_6634);
xnor U10731 (N_10731,N_6741,N_6194);
xnor U10732 (N_10732,N_6969,N_7543);
or U10733 (N_10733,N_6410,N_8799);
and U10734 (N_10734,N_7296,N_8052);
nand U10735 (N_10735,N_8761,N_6353);
xnor U10736 (N_10736,N_7867,N_8888);
nor U10737 (N_10737,N_6084,N_7486);
and U10738 (N_10738,N_6011,N_6359);
nand U10739 (N_10739,N_7718,N_8014);
and U10740 (N_10740,N_8328,N_7679);
and U10741 (N_10741,N_8646,N_7808);
nor U10742 (N_10742,N_7962,N_6626);
nand U10743 (N_10743,N_7750,N_8731);
or U10744 (N_10744,N_7526,N_6098);
or U10745 (N_10745,N_7533,N_7127);
and U10746 (N_10746,N_7626,N_8557);
or U10747 (N_10747,N_7730,N_7995);
xor U10748 (N_10748,N_8745,N_6684);
xnor U10749 (N_10749,N_6955,N_8910);
or U10750 (N_10750,N_6388,N_6313);
or U10751 (N_10751,N_7979,N_8073);
xnor U10752 (N_10752,N_6508,N_8514);
and U10753 (N_10753,N_6774,N_6145);
xnor U10754 (N_10754,N_7792,N_6909);
nand U10755 (N_10755,N_7644,N_7343);
xor U10756 (N_10756,N_8085,N_8081);
xnor U10757 (N_10757,N_8765,N_6312);
and U10758 (N_10758,N_8600,N_7840);
or U10759 (N_10759,N_8378,N_6364);
xor U10760 (N_10760,N_7123,N_7959);
xor U10761 (N_10761,N_8271,N_8884);
xor U10762 (N_10762,N_8645,N_7505);
or U10763 (N_10763,N_7155,N_7236);
nor U10764 (N_10764,N_7932,N_7187);
and U10765 (N_10765,N_7755,N_7553);
nand U10766 (N_10766,N_7833,N_7409);
nor U10767 (N_10767,N_6195,N_7047);
nand U10768 (N_10768,N_7128,N_7864);
or U10769 (N_10769,N_7305,N_7002);
nand U10770 (N_10770,N_8944,N_7670);
xor U10771 (N_10771,N_7069,N_8704);
or U10772 (N_10772,N_7030,N_8833);
nor U10773 (N_10773,N_6328,N_8597);
nand U10774 (N_10774,N_7122,N_8013);
or U10775 (N_10775,N_7476,N_8260);
nand U10776 (N_10776,N_7688,N_7673);
xnor U10777 (N_10777,N_6372,N_8344);
and U10778 (N_10778,N_6528,N_8767);
xnor U10779 (N_10779,N_6432,N_7067);
nor U10780 (N_10780,N_8473,N_8716);
nor U10781 (N_10781,N_8682,N_8551);
nor U10782 (N_10782,N_6371,N_7664);
nor U10783 (N_10783,N_6492,N_6384);
nor U10784 (N_10784,N_8450,N_8764);
and U10785 (N_10785,N_7426,N_7173);
nor U10786 (N_10786,N_7073,N_7848);
nor U10787 (N_10787,N_8535,N_7422);
nand U10788 (N_10788,N_7668,N_8134);
nand U10789 (N_10789,N_8184,N_7548);
or U10790 (N_10790,N_8139,N_8620);
and U10791 (N_10791,N_8623,N_6349);
nor U10792 (N_10792,N_8947,N_7076);
and U10793 (N_10793,N_7247,N_6005);
nand U10794 (N_10794,N_6803,N_8207);
xnor U10795 (N_10795,N_6325,N_7540);
nor U10796 (N_10796,N_7870,N_6279);
nand U10797 (N_10797,N_8405,N_6525);
xnor U10798 (N_10798,N_6043,N_7231);
or U10799 (N_10799,N_6853,N_7372);
nor U10800 (N_10800,N_7949,N_7538);
and U10801 (N_10801,N_8079,N_6280);
nand U10802 (N_10802,N_7196,N_7001);
or U10803 (N_10803,N_7638,N_8343);
xnor U10804 (N_10804,N_6010,N_6357);
xor U10805 (N_10805,N_7440,N_6924);
nand U10806 (N_10806,N_7794,N_6962);
nor U10807 (N_10807,N_6979,N_8494);
nand U10808 (N_10808,N_7075,N_6108);
nor U10809 (N_10809,N_7001,N_6201);
or U10810 (N_10810,N_7247,N_8210);
and U10811 (N_10811,N_8996,N_8316);
or U10812 (N_10812,N_8881,N_7273);
nand U10813 (N_10813,N_6230,N_7043);
nand U10814 (N_10814,N_8142,N_6751);
xnor U10815 (N_10815,N_7891,N_7623);
nand U10816 (N_10816,N_6702,N_8741);
nand U10817 (N_10817,N_8521,N_6892);
or U10818 (N_10818,N_6461,N_8261);
or U10819 (N_10819,N_6743,N_8840);
nor U10820 (N_10820,N_7876,N_8147);
and U10821 (N_10821,N_6325,N_8252);
nand U10822 (N_10822,N_7167,N_8656);
and U10823 (N_10823,N_8139,N_6172);
or U10824 (N_10824,N_7498,N_7438);
or U10825 (N_10825,N_6447,N_8863);
or U10826 (N_10826,N_8187,N_6315);
nor U10827 (N_10827,N_6441,N_6413);
nand U10828 (N_10828,N_6930,N_6204);
or U10829 (N_10829,N_6010,N_6242);
xor U10830 (N_10830,N_8502,N_8011);
xnor U10831 (N_10831,N_8838,N_7275);
nor U10832 (N_10832,N_6885,N_7465);
nand U10833 (N_10833,N_6199,N_6017);
and U10834 (N_10834,N_7755,N_6466);
and U10835 (N_10835,N_8956,N_7457);
and U10836 (N_10836,N_8482,N_6476);
or U10837 (N_10837,N_6740,N_8257);
nand U10838 (N_10838,N_6905,N_8519);
or U10839 (N_10839,N_7556,N_8561);
nand U10840 (N_10840,N_8451,N_8126);
and U10841 (N_10841,N_8258,N_7782);
or U10842 (N_10842,N_7132,N_8560);
nor U10843 (N_10843,N_7092,N_6815);
xor U10844 (N_10844,N_7057,N_8963);
or U10845 (N_10845,N_7432,N_6888);
nand U10846 (N_10846,N_6151,N_7780);
xnor U10847 (N_10847,N_6293,N_8954);
or U10848 (N_10848,N_7440,N_8231);
nor U10849 (N_10849,N_6325,N_7245);
and U10850 (N_10850,N_7639,N_8903);
and U10851 (N_10851,N_6298,N_7652);
or U10852 (N_10852,N_6139,N_8033);
nor U10853 (N_10853,N_8401,N_6799);
or U10854 (N_10854,N_6531,N_6278);
nor U10855 (N_10855,N_6412,N_6851);
xor U10856 (N_10856,N_8785,N_6067);
and U10857 (N_10857,N_8667,N_6592);
xnor U10858 (N_10858,N_7611,N_7812);
nand U10859 (N_10859,N_7314,N_7831);
nor U10860 (N_10860,N_7190,N_6669);
and U10861 (N_10861,N_8642,N_7082);
and U10862 (N_10862,N_8439,N_6046);
nor U10863 (N_10863,N_6609,N_7684);
nor U10864 (N_10864,N_8689,N_8085);
or U10865 (N_10865,N_7635,N_7539);
nor U10866 (N_10866,N_8151,N_6054);
nand U10867 (N_10867,N_7648,N_7230);
nand U10868 (N_10868,N_8603,N_6494);
or U10869 (N_10869,N_8799,N_8175);
xor U10870 (N_10870,N_6567,N_7985);
and U10871 (N_10871,N_7287,N_7227);
nand U10872 (N_10872,N_7978,N_7551);
or U10873 (N_10873,N_6440,N_7359);
xor U10874 (N_10874,N_8011,N_7987);
or U10875 (N_10875,N_8581,N_6636);
or U10876 (N_10876,N_6227,N_7735);
or U10877 (N_10877,N_7424,N_7131);
and U10878 (N_10878,N_8185,N_7691);
xor U10879 (N_10879,N_7452,N_6705);
nand U10880 (N_10880,N_8716,N_8585);
and U10881 (N_10881,N_8692,N_7204);
nand U10882 (N_10882,N_7764,N_8086);
or U10883 (N_10883,N_6137,N_6893);
and U10884 (N_10884,N_8320,N_6000);
nor U10885 (N_10885,N_7605,N_6485);
xnor U10886 (N_10886,N_8970,N_6181);
xnor U10887 (N_10887,N_7536,N_8663);
or U10888 (N_10888,N_7507,N_8428);
or U10889 (N_10889,N_7675,N_8916);
xnor U10890 (N_10890,N_6361,N_6970);
nor U10891 (N_10891,N_7263,N_6922);
nand U10892 (N_10892,N_7211,N_8120);
nor U10893 (N_10893,N_7155,N_7779);
or U10894 (N_10894,N_7025,N_7482);
or U10895 (N_10895,N_8524,N_7535);
nor U10896 (N_10896,N_7590,N_6550);
and U10897 (N_10897,N_8950,N_8207);
nor U10898 (N_10898,N_7526,N_6499);
nand U10899 (N_10899,N_7167,N_7931);
xnor U10900 (N_10900,N_8318,N_8723);
and U10901 (N_10901,N_6295,N_6612);
nand U10902 (N_10902,N_6335,N_6956);
or U10903 (N_10903,N_8584,N_7838);
or U10904 (N_10904,N_6946,N_6902);
and U10905 (N_10905,N_6766,N_6217);
or U10906 (N_10906,N_7852,N_8372);
and U10907 (N_10907,N_6033,N_7162);
nor U10908 (N_10908,N_6821,N_8251);
and U10909 (N_10909,N_8601,N_6573);
nor U10910 (N_10910,N_6118,N_7720);
xor U10911 (N_10911,N_6662,N_6363);
nor U10912 (N_10912,N_8927,N_6502);
or U10913 (N_10913,N_6404,N_6919);
nor U10914 (N_10914,N_8857,N_7514);
nand U10915 (N_10915,N_8564,N_6025);
nand U10916 (N_10916,N_6375,N_8346);
and U10917 (N_10917,N_8574,N_8585);
and U10918 (N_10918,N_6244,N_8919);
xnor U10919 (N_10919,N_7839,N_6462);
nand U10920 (N_10920,N_7114,N_7100);
xnor U10921 (N_10921,N_6513,N_7744);
nand U10922 (N_10922,N_7723,N_7616);
and U10923 (N_10923,N_6859,N_8508);
nand U10924 (N_10924,N_6229,N_7249);
or U10925 (N_10925,N_7287,N_6517);
nand U10926 (N_10926,N_8150,N_8280);
and U10927 (N_10927,N_7738,N_7749);
and U10928 (N_10928,N_7232,N_8104);
xor U10929 (N_10929,N_8546,N_6963);
nand U10930 (N_10930,N_7687,N_7202);
nor U10931 (N_10931,N_6186,N_8137);
nand U10932 (N_10932,N_6800,N_7689);
xnor U10933 (N_10933,N_7266,N_8495);
nand U10934 (N_10934,N_8685,N_7445);
xor U10935 (N_10935,N_8976,N_8677);
or U10936 (N_10936,N_7444,N_7410);
or U10937 (N_10937,N_8897,N_6582);
xnor U10938 (N_10938,N_6614,N_6826);
nand U10939 (N_10939,N_7225,N_6983);
and U10940 (N_10940,N_8439,N_6342);
nand U10941 (N_10941,N_8415,N_6675);
nor U10942 (N_10942,N_7539,N_8144);
nand U10943 (N_10943,N_8080,N_8035);
nand U10944 (N_10944,N_7545,N_8156);
nand U10945 (N_10945,N_7199,N_8308);
or U10946 (N_10946,N_7385,N_7335);
and U10947 (N_10947,N_7338,N_8317);
and U10948 (N_10948,N_7069,N_7281);
xnor U10949 (N_10949,N_6975,N_7148);
nand U10950 (N_10950,N_6445,N_8082);
or U10951 (N_10951,N_6866,N_7176);
or U10952 (N_10952,N_7205,N_7519);
nor U10953 (N_10953,N_6581,N_6911);
or U10954 (N_10954,N_6508,N_7896);
nor U10955 (N_10955,N_7937,N_7781);
nor U10956 (N_10956,N_8065,N_8810);
and U10957 (N_10957,N_8465,N_7324);
or U10958 (N_10958,N_8030,N_8434);
or U10959 (N_10959,N_6860,N_7658);
nand U10960 (N_10960,N_6407,N_7616);
or U10961 (N_10961,N_8051,N_6294);
or U10962 (N_10962,N_6484,N_6201);
or U10963 (N_10963,N_6210,N_7603);
nor U10964 (N_10964,N_7202,N_7233);
or U10965 (N_10965,N_6692,N_8669);
xor U10966 (N_10966,N_6157,N_7138);
xor U10967 (N_10967,N_8863,N_7987);
xnor U10968 (N_10968,N_7278,N_7474);
or U10969 (N_10969,N_6298,N_8441);
nor U10970 (N_10970,N_7651,N_8367);
and U10971 (N_10971,N_7500,N_8102);
xnor U10972 (N_10972,N_8012,N_8911);
nand U10973 (N_10973,N_8072,N_6145);
xnor U10974 (N_10974,N_6203,N_7932);
xnor U10975 (N_10975,N_8023,N_7908);
nand U10976 (N_10976,N_6687,N_6500);
and U10977 (N_10977,N_6378,N_8750);
or U10978 (N_10978,N_7862,N_8978);
or U10979 (N_10979,N_7298,N_6528);
or U10980 (N_10980,N_8982,N_6459);
nand U10981 (N_10981,N_7651,N_6950);
or U10982 (N_10982,N_7139,N_7876);
xnor U10983 (N_10983,N_8255,N_7399);
or U10984 (N_10984,N_7420,N_7640);
nor U10985 (N_10985,N_6702,N_7836);
and U10986 (N_10986,N_8201,N_6183);
or U10987 (N_10987,N_8370,N_7708);
xnor U10988 (N_10988,N_6319,N_8756);
nor U10989 (N_10989,N_8231,N_6117);
nor U10990 (N_10990,N_8856,N_7725);
nand U10991 (N_10991,N_8484,N_7546);
or U10992 (N_10992,N_8314,N_7289);
and U10993 (N_10993,N_8449,N_6284);
nand U10994 (N_10994,N_6086,N_7851);
and U10995 (N_10995,N_6548,N_8322);
nand U10996 (N_10996,N_6762,N_7910);
or U10997 (N_10997,N_8003,N_6646);
or U10998 (N_10998,N_8795,N_8180);
xnor U10999 (N_10999,N_7095,N_8246);
nor U11000 (N_11000,N_8026,N_6301);
nand U11001 (N_11001,N_7508,N_6690);
or U11002 (N_11002,N_8959,N_7940);
xor U11003 (N_11003,N_8132,N_6302);
or U11004 (N_11004,N_8523,N_6764);
nand U11005 (N_11005,N_8007,N_6970);
xnor U11006 (N_11006,N_7614,N_7142);
xnor U11007 (N_11007,N_7103,N_8378);
and U11008 (N_11008,N_8791,N_7265);
nor U11009 (N_11009,N_8169,N_7813);
or U11010 (N_11010,N_6193,N_6082);
nand U11011 (N_11011,N_6991,N_7855);
nor U11012 (N_11012,N_8985,N_8476);
nor U11013 (N_11013,N_8503,N_7202);
xnor U11014 (N_11014,N_7432,N_6064);
nand U11015 (N_11015,N_8069,N_7229);
or U11016 (N_11016,N_8058,N_8139);
nor U11017 (N_11017,N_7358,N_7114);
xor U11018 (N_11018,N_8224,N_6057);
and U11019 (N_11019,N_6175,N_8097);
nor U11020 (N_11020,N_7781,N_6333);
and U11021 (N_11021,N_6403,N_8024);
xnor U11022 (N_11022,N_6940,N_7020);
or U11023 (N_11023,N_7214,N_8702);
nor U11024 (N_11024,N_7242,N_8556);
xor U11025 (N_11025,N_7403,N_6236);
nand U11026 (N_11026,N_7976,N_6886);
nor U11027 (N_11027,N_7867,N_6711);
nand U11028 (N_11028,N_7446,N_7757);
xor U11029 (N_11029,N_6507,N_6069);
nand U11030 (N_11030,N_8543,N_8763);
and U11031 (N_11031,N_7085,N_6255);
and U11032 (N_11032,N_8576,N_7128);
or U11033 (N_11033,N_7302,N_7878);
or U11034 (N_11034,N_8651,N_7512);
and U11035 (N_11035,N_8972,N_7852);
xor U11036 (N_11036,N_6808,N_8784);
and U11037 (N_11037,N_6958,N_8095);
xnor U11038 (N_11038,N_8569,N_7236);
nand U11039 (N_11039,N_8240,N_8756);
nand U11040 (N_11040,N_7657,N_6921);
and U11041 (N_11041,N_8880,N_6571);
xnor U11042 (N_11042,N_7217,N_8836);
nor U11043 (N_11043,N_8402,N_8589);
xnor U11044 (N_11044,N_7747,N_8321);
or U11045 (N_11045,N_6505,N_6573);
nand U11046 (N_11046,N_8407,N_6000);
or U11047 (N_11047,N_8351,N_6063);
nor U11048 (N_11048,N_6998,N_6192);
and U11049 (N_11049,N_6184,N_8682);
or U11050 (N_11050,N_8406,N_6481);
xnor U11051 (N_11051,N_7948,N_6895);
nor U11052 (N_11052,N_6261,N_6827);
nor U11053 (N_11053,N_8996,N_7788);
xnor U11054 (N_11054,N_8216,N_7666);
and U11055 (N_11055,N_7776,N_6122);
or U11056 (N_11056,N_6695,N_6964);
nand U11057 (N_11057,N_7063,N_7541);
or U11058 (N_11058,N_8597,N_8149);
nand U11059 (N_11059,N_6688,N_6677);
nor U11060 (N_11060,N_7753,N_6425);
nor U11061 (N_11061,N_8585,N_8057);
or U11062 (N_11062,N_6960,N_8305);
nor U11063 (N_11063,N_7489,N_6786);
or U11064 (N_11064,N_7001,N_8633);
and U11065 (N_11065,N_6010,N_7566);
and U11066 (N_11066,N_8837,N_8809);
and U11067 (N_11067,N_8062,N_7352);
nand U11068 (N_11068,N_8648,N_8416);
or U11069 (N_11069,N_7711,N_6735);
or U11070 (N_11070,N_6104,N_6541);
xor U11071 (N_11071,N_7191,N_7571);
nand U11072 (N_11072,N_8971,N_7846);
xor U11073 (N_11073,N_7314,N_8405);
xor U11074 (N_11074,N_6671,N_8062);
nand U11075 (N_11075,N_6817,N_7348);
xnor U11076 (N_11076,N_6697,N_8712);
or U11077 (N_11077,N_7581,N_6525);
nand U11078 (N_11078,N_6230,N_8636);
xnor U11079 (N_11079,N_6490,N_6770);
and U11080 (N_11080,N_6492,N_7721);
nor U11081 (N_11081,N_8022,N_8463);
and U11082 (N_11082,N_8504,N_7361);
and U11083 (N_11083,N_8033,N_6539);
or U11084 (N_11084,N_8735,N_7826);
or U11085 (N_11085,N_8265,N_7461);
xor U11086 (N_11086,N_6255,N_6139);
nor U11087 (N_11087,N_6686,N_8023);
nand U11088 (N_11088,N_6216,N_6351);
xnor U11089 (N_11089,N_8489,N_8683);
or U11090 (N_11090,N_6086,N_8494);
xor U11091 (N_11091,N_6573,N_6222);
and U11092 (N_11092,N_8956,N_8045);
nand U11093 (N_11093,N_7339,N_7415);
nor U11094 (N_11094,N_8966,N_6439);
nand U11095 (N_11095,N_7228,N_6166);
or U11096 (N_11096,N_8353,N_6909);
nor U11097 (N_11097,N_8798,N_8449);
nand U11098 (N_11098,N_8391,N_6824);
or U11099 (N_11099,N_6225,N_8158);
nor U11100 (N_11100,N_6487,N_7441);
nand U11101 (N_11101,N_7782,N_7502);
nand U11102 (N_11102,N_8571,N_7667);
and U11103 (N_11103,N_6694,N_8844);
or U11104 (N_11104,N_6703,N_6445);
nand U11105 (N_11105,N_6653,N_6164);
nor U11106 (N_11106,N_6771,N_8912);
nand U11107 (N_11107,N_6682,N_7526);
xor U11108 (N_11108,N_7479,N_6703);
or U11109 (N_11109,N_6867,N_7113);
xor U11110 (N_11110,N_6438,N_7475);
and U11111 (N_11111,N_6558,N_8302);
and U11112 (N_11112,N_7427,N_6518);
and U11113 (N_11113,N_8967,N_6325);
or U11114 (N_11114,N_8225,N_6580);
or U11115 (N_11115,N_7620,N_6270);
xnor U11116 (N_11116,N_6491,N_6345);
or U11117 (N_11117,N_8402,N_7229);
or U11118 (N_11118,N_7803,N_8556);
nor U11119 (N_11119,N_7864,N_6987);
or U11120 (N_11120,N_8434,N_7763);
nand U11121 (N_11121,N_8622,N_8263);
xnor U11122 (N_11122,N_8367,N_6539);
and U11123 (N_11123,N_8561,N_6427);
xor U11124 (N_11124,N_8071,N_8481);
and U11125 (N_11125,N_6279,N_8445);
nand U11126 (N_11126,N_7524,N_7913);
nand U11127 (N_11127,N_8754,N_7197);
or U11128 (N_11128,N_7379,N_7271);
nand U11129 (N_11129,N_7648,N_7720);
xnor U11130 (N_11130,N_7810,N_8969);
xnor U11131 (N_11131,N_7384,N_6226);
or U11132 (N_11132,N_6824,N_6627);
or U11133 (N_11133,N_8039,N_7366);
nand U11134 (N_11134,N_7275,N_6094);
xnor U11135 (N_11135,N_7188,N_8198);
nor U11136 (N_11136,N_6784,N_6760);
nor U11137 (N_11137,N_6698,N_7656);
or U11138 (N_11138,N_8338,N_8564);
or U11139 (N_11139,N_6730,N_6915);
xor U11140 (N_11140,N_7804,N_6123);
or U11141 (N_11141,N_7628,N_7564);
and U11142 (N_11142,N_8688,N_6209);
nand U11143 (N_11143,N_6716,N_8430);
nor U11144 (N_11144,N_6112,N_6799);
nor U11145 (N_11145,N_8692,N_8614);
xnor U11146 (N_11146,N_8078,N_6216);
and U11147 (N_11147,N_6738,N_6381);
or U11148 (N_11148,N_8733,N_6188);
nor U11149 (N_11149,N_6866,N_6803);
xnor U11150 (N_11150,N_6039,N_8041);
or U11151 (N_11151,N_6695,N_7331);
and U11152 (N_11152,N_6612,N_8310);
nand U11153 (N_11153,N_8404,N_8080);
or U11154 (N_11154,N_6000,N_6099);
and U11155 (N_11155,N_8368,N_8065);
nand U11156 (N_11156,N_8116,N_8273);
nor U11157 (N_11157,N_7664,N_8646);
xnor U11158 (N_11158,N_6766,N_7043);
xnor U11159 (N_11159,N_7996,N_7729);
nand U11160 (N_11160,N_8853,N_7934);
nor U11161 (N_11161,N_8486,N_7597);
or U11162 (N_11162,N_6345,N_6278);
nand U11163 (N_11163,N_8964,N_8764);
nand U11164 (N_11164,N_7200,N_8699);
and U11165 (N_11165,N_7877,N_8420);
xnor U11166 (N_11166,N_8896,N_6740);
nand U11167 (N_11167,N_8775,N_6675);
and U11168 (N_11168,N_8977,N_7773);
nor U11169 (N_11169,N_8217,N_6073);
or U11170 (N_11170,N_7967,N_7667);
nor U11171 (N_11171,N_7009,N_6665);
and U11172 (N_11172,N_8640,N_8770);
and U11173 (N_11173,N_8689,N_6820);
and U11174 (N_11174,N_8793,N_6679);
or U11175 (N_11175,N_8280,N_6675);
or U11176 (N_11176,N_6955,N_6183);
nand U11177 (N_11177,N_7757,N_7510);
nor U11178 (N_11178,N_7400,N_8357);
xor U11179 (N_11179,N_6079,N_8256);
xnor U11180 (N_11180,N_6383,N_6758);
nand U11181 (N_11181,N_8923,N_7849);
nor U11182 (N_11182,N_7721,N_6342);
nand U11183 (N_11183,N_7600,N_7767);
or U11184 (N_11184,N_6137,N_7848);
nor U11185 (N_11185,N_6849,N_7481);
and U11186 (N_11186,N_6056,N_6998);
and U11187 (N_11187,N_6484,N_7770);
or U11188 (N_11188,N_6664,N_8178);
or U11189 (N_11189,N_7466,N_7988);
nand U11190 (N_11190,N_8910,N_7328);
xnor U11191 (N_11191,N_7531,N_7773);
nor U11192 (N_11192,N_7659,N_6445);
nand U11193 (N_11193,N_6459,N_6389);
nand U11194 (N_11194,N_8083,N_8832);
nor U11195 (N_11195,N_7102,N_7961);
nand U11196 (N_11196,N_7789,N_8004);
nor U11197 (N_11197,N_8570,N_6355);
nor U11198 (N_11198,N_8768,N_6546);
nor U11199 (N_11199,N_7964,N_7267);
and U11200 (N_11200,N_7147,N_8670);
nand U11201 (N_11201,N_6735,N_8928);
or U11202 (N_11202,N_8161,N_7519);
or U11203 (N_11203,N_7984,N_8745);
xor U11204 (N_11204,N_7470,N_6749);
nor U11205 (N_11205,N_7396,N_8712);
nand U11206 (N_11206,N_8382,N_7674);
or U11207 (N_11207,N_6240,N_6899);
and U11208 (N_11208,N_6156,N_7208);
nor U11209 (N_11209,N_8201,N_8133);
nand U11210 (N_11210,N_8128,N_8672);
nand U11211 (N_11211,N_8247,N_7443);
and U11212 (N_11212,N_8320,N_6386);
or U11213 (N_11213,N_8377,N_7175);
or U11214 (N_11214,N_8480,N_7433);
nor U11215 (N_11215,N_6783,N_7837);
and U11216 (N_11216,N_7057,N_6321);
nor U11217 (N_11217,N_8810,N_6313);
xor U11218 (N_11218,N_7064,N_6313);
xor U11219 (N_11219,N_8490,N_7893);
nor U11220 (N_11220,N_6683,N_6131);
and U11221 (N_11221,N_8335,N_6389);
xor U11222 (N_11222,N_7090,N_8290);
nand U11223 (N_11223,N_7064,N_7880);
nor U11224 (N_11224,N_7327,N_6299);
or U11225 (N_11225,N_8655,N_7632);
xnor U11226 (N_11226,N_6469,N_6962);
nor U11227 (N_11227,N_6760,N_8294);
xnor U11228 (N_11228,N_7185,N_7812);
or U11229 (N_11229,N_8589,N_7091);
nand U11230 (N_11230,N_7096,N_7281);
xnor U11231 (N_11231,N_8550,N_8791);
nand U11232 (N_11232,N_8585,N_8098);
xnor U11233 (N_11233,N_7213,N_7689);
nand U11234 (N_11234,N_6954,N_6176);
or U11235 (N_11235,N_7733,N_8939);
or U11236 (N_11236,N_6162,N_7037);
and U11237 (N_11237,N_7293,N_8155);
nor U11238 (N_11238,N_8672,N_7573);
nor U11239 (N_11239,N_8899,N_8351);
and U11240 (N_11240,N_8743,N_6656);
and U11241 (N_11241,N_6875,N_8553);
or U11242 (N_11242,N_7126,N_8934);
and U11243 (N_11243,N_6192,N_7342);
xnor U11244 (N_11244,N_6069,N_6640);
or U11245 (N_11245,N_6652,N_8391);
nor U11246 (N_11246,N_7764,N_6394);
and U11247 (N_11247,N_8911,N_8381);
or U11248 (N_11248,N_6139,N_6895);
and U11249 (N_11249,N_6812,N_8764);
and U11250 (N_11250,N_7129,N_8531);
or U11251 (N_11251,N_6678,N_6345);
xnor U11252 (N_11252,N_8705,N_8390);
nand U11253 (N_11253,N_7669,N_7886);
and U11254 (N_11254,N_8349,N_8166);
xnor U11255 (N_11255,N_7651,N_7322);
or U11256 (N_11256,N_7344,N_6930);
nand U11257 (N_11257,N_6630,N_6280);
nand U11258 (N_11258,N_8348,N_6694);
and U11259 (N_11259,N_6001,N_6747);
nor U11260 (N_11260,N_7528,N_6252);
nand U11261 (N_11261,N_8216,N_7047);
xnor U11262 (N_11262,N_7280,N_7301);
and U11263 (N_11263,N_8308,N_8923);
nand U11264 (N_11264,N_8260,N_7675);
and U11265 (N_11265,N_6499,N_6311);
nand U11266 (N_11266,N_7890,N_8564);
nand U11267 (N_11267,N_7882,N_6950);
nor U11268 (N_11268,N_7406,N_8845);
and U11269 (N_11269,N_6779,N_7868);
nand U11270 (N_11270,N_7161,N_8061);
nor U11271 (N_11271,N_8541,N_6174);
and U11272 (N_11272,N_7131,N_6852);
xor U11273 (N_11273,N_8780,N_6426);
nand U11274 (N_11274,N_8429,N_7129);
and U11275 (N_11275,N_6683,N_7341);
and U11276 (N_11276,N_8988,N_6723);
or U11277 (N_11277,N_8981,N_8418);
nor U11278 (N_11278,N_6801,N_6260);
nand U11279 (N_11279,N_6729,N_8384);
nand U11280 (N_11280,N_7422,N_8213);
and U11281 (N_11281,N_8724,N_7454);
nor U11282 (N_11282,N_6945,N_8521);
xnor U11283 (N_11283,N_7723,N_8564);
and U11284 (N_11284,N_6785,N_6432);
or U11285 (N_11285,N_6736,N_8752);
nor U11286 (N_11286,N_6096,N_7664);
or U11287 (N_11287,N_7430,N_6947);
xnor U11288 (N_11288,N_6796,N_8092);
nor U11289 (N_11289,N_7162,N_6736);
nor U11290 (N_11290,N_6009,N_7503);
nor U11291 (N_11291,N_6504,N_8816);
and U11292 (N_11292,N_7426,N_6408);
nand U11293 (N_11293,N_7886,N_7594);
or U11294 (N_11294,N_8592,N_7331);
and U11295 (N_11295,N_8336,N_7965);
nor U11296 (N_11296,N_6406,N_6313);
nand U11297 (N_11297,N_6234,N_8246);
nand U11298 (N_11298,N_8645,N_8218);
xnor U11299 (N_11299,N_8953,N_7983);
nand U11300 (N_11300,N_7954,N_6400);
nor U11301 (N_11301,N_7146,N_8535);
nor U11302 (N_11302,N_8563,N_7698);
xor U11303 (N_11303,N_7900,N_8980);
nand U11304 (N_11304,N_6771,N_6316);
nor U11305 (N_11305,N_7248,N_7508);
xnor U11306 (N_11306,N_8082,N_8047);
nor U11307 (N_11307,N_7654,N_6957);
nand U11308 (N_11308,N_6586,N_7087);
and U11309 (N_11309,N_6545,N_8108);
and U11310 (N_11310,N_7690,N_6549);
and U11311 (N_11311,N_7894,N_8628);
nor U11312 (N_11312,N_6710,N_6378);
nand U11313 (N_11313,N_6594,N_8309);
or U11314 (N_11314,N_7517,N_7552);
nor U11315 (N_11315,N_8782,N_6116);
xor U11316 (N_11316,N_6306,N_6677);
nand U11317 (N_11317,N_8393,N_6420);
nor U11318 (N_11318,N_7823,N_6182);
and U11319 (N_11319,N_6272,N_8184);
and U11320 (N_11320,N_8292,N_7525);
nor U11321 (N_11321,N_8327,N_8886);
xnor U11322 (N_11322,N_7308,N_8313);
xnor U11323 (N_11323,N_6938,N_7056);
or U11324 (N_11324,N_7014,N_6873);
nor U11325 (N_11325,N_6042,N_7954);
nor U11326 (N_11326,N_6483,N_8398);
xor U11327 (N_11327,N_7216,N_8722);
or U11328 (N_11328,N_8853,N_8448);
xor U11329 (N_11329,N_8574,N_8963);
nand U11330 (N_11330,N_6669,N_7771);
xnor U11331 (N_11331,N_7978,N_6469);
nor U11332 (N_11332,N_6834,N_8673);
nor U11333 (N_11333,N_7752,N_8222);
nor U11334 (N_11334,N_8962,N_8250);
nand U11335 (N_11335,N_7647,N_8821);
or U11336 (N_11336,N_8453,N_8207);
or U11337 (N_11337,N_6927,N_8862);
nor U11338 (N_11338,N_7068,N_7073);
and U11339 (N_11339,N_8587,N_7089);
xnor U11340 (N_11340,N_8463,N_8260);
and U11341 (N_11341,N_6841,N_6382);
nand U11342 (N_11342,N_8902,N_6935);
xnor U11343 (N_11343,N_7545,N_6554);
nor U11344 (N_11344,N_8276,N_8145);
xnor U11345 (N_11345,N_8112,N_7791);
and U11346 (N_11346,N_8696,N_6065);
xor U11347 (N_11347,N_8761,N_7221);
and U11348 (N_11348,N_8557,N_6333);
or U11349 (N_11349,N_7272,N_8969);
nor U11350 (N_11350,N_7910,N_7790);
or U11351 (N_11351,N_7750,N_7242);
and U11352 (N_11352,N_8272,N_6096);
nor U11353 (N_11353,N_7566,N_7786);
nor U11354 (N_11354,N_8997,N_8176);
or U11355 (N_11355,N_7029,N_8037);
nor U11356 (N_11356,N_6794,N_8095);
and U11357 (N_11357,N_7317,N_7737);
and U11358 (N_11358,N_8975,N_8695);
xor U11359 (N_11359,N_8692,N_8789);
xor U11360 (N_11360,N_8249,N_7170);
or U11361 (N_11361,N_6246,N_7652);
xnor U11362 (N_11362,N_8237,N_7428);
and U11363 (N_11363,N_6792,N_8329);
xnor U11364 (N_11364,N_7445,N_6799);
nor U11365 (N_11365,N_8973,N_8463);
nand U11366 (N_11366,N_7437,N_8291);
or U11367 (N_11367,N_7580,N_7650);
nor U11368 (N_11368,N_7390,N_7970);
and U11369 (N_11369,N_7015,N_6836);
and U11370 (N_11370,N_6604,N_6295);
xnor U11371 (N_11371,N_7073,N_6776);
xor U11372 (N_11372,N_6814,N_7482);
xor U11373 (N_11373,N_8946,N_8600);
xnor U11374 (N_11374,N_8956,N_7904);
and U11375 (N_11375,N_6618,N_6401);
xor U11376 (N_11376,N_8901,N_6477);
and U11377 (N_11377,N_7984,N_6854);
and U11378 (N_11378,N_7730,N_6170);
nand U11379 (N_11379,N_8446,N_8149);
and U11380 (N_11380,N_8849,N_8458);
or U11381 (N_11381,N_7635,N_7987);
nand U11382 (N_11382,N_7388,N_7357);
nor U11383 (N_11383,N_6104,N_7606);
and U11384 (N_11384,N_7588,N_8179);
or U11385 (N_11385,N_7016,N_8732);
nand U11386 (N_11386,N_7852,N_8989);
nand U11387 (N_11387,N_7985,N_8005);
nor U11388 (N_11388,N_6953,N_8150);
and U11389 (N_11389,N_8123,N_6798);
nor U11390 (N_11390,N_6833,N_8818);
xnor U11391 (N_11391,N_8253,N_6446);
or U11392 (N_11392,N_7096,N_6406);
and U11393 (N_11393,N_8952,N_6523);
or U11394 (N_11394,N_7295,N_7923);
or U11395 (N_11395,N_8227,N_7019);
nand U11396 (N_11396,N_7479,N_8501);
or U11397 (N_11397,N_8790,N_6793);
xor U11398 (N_11398,N_8429,N_7098);
and U11399 (N_11399,N_6924,N_6239);
nor U11400 (N_11400,N_7768,N_7514);
or U11401 (N_11401,N_7902,N_6866);
nor U11402 (N_11402,N_6015,N_7263);
nand U11403 (N_11403,N_8831,N_6539);
or U11404 (N_11404,N_6874,N_8217);
nor U11405 (N_11405,N_6530,N_8936);
nor U11406 (N_11406,N_7242,N_8440);
nor U11407 (N_11407,N_7119,N_8395);
and U11408 (N_11408,N_8496,N_7615);
and U11409 (N_11409,N_7931,N_8640);
nand U11410 (N_11410,N_8492,N_6630);
xnor U11411 (N_11411,N_8969,N_6855);
or U11412 (N_11412,N_6841,N_8398);
or U11413 (N_11413,N_6233,N_6361);
xnor U11414 (N_11414,N_8216,N_6217);
xor U11415 (N_11415,N_7430,N_6398);
xnor U11416 (N_11416,N_6667,N_8784);
nor U11417 (N_11417,N_7307,N_8000);
xnor U11418 (N_11418,N_8178,N_6663);
nor U11419 (N_11419,N_8693,N_7445);
nand U11420 (N_11420,N_6617,N_6397);
or U11421 (N_11421,N_8002,N_6340);
nor U11422 (N_11422,N_6327,N_6028);
xnor U11423 (N_11423,N_6932,N_6471);
and U11424 (N_11424,N_6140,N_6509);
nor U11425 (N_11425,N_8155,N_6932);
nand U11426 (N_11426,N_8013,N_7344);
nor U11427 (N_11427,N_6839,N_7768);
nand U11428 (N_11428,N_8390,N_8506);
and U11429 (N_11429,N_7062,N_8140);
nor U11430 (N_11430,N_8299,N_8122);
nor U11431 (N_11431,N_6833,N_6810);
nand U11432 (N_11432,N_7193,N_8467);
or U11433 (N_11433,N_8599,N_6121);
nand U11434 (N_11434,N_7219,N_8385);
or U11435 (N_11435,N_8185,N_6462);
and U11436 (N_11436,N_7584,N_6829);
or U11437 (N_11437,N_7731,N_8112);
nor U11438 (N_11438,N_7832,N_7644);
nand U11439 (N_11439,N_8662,N_6923);
and U11440 (N_11440,N_8737,N_6632);
nor U11441 (N_11441,N_8014,N_6946);
xnor U11442 (N_11442,N_8677,N_8231);
nor U11443 (N_11443,N_7536,N_7739);
and U11444 (N_11444,N_8151,N_8406);
or U11445 (N_11445,N_8175,N_7189);
and U11446 (N_11446,N_8852,N_8439);
nor U11447 (N_11447,N_8678,N_6525);
or U11448 (N_11448,N_6828,N_8442);
xor U11449 (N_11449,N_6227,N_8981);
nand U11450 (N_11450,N_6737,N_6566);
or U11451 (N_11451,N_6919,N_8413);
and U11452 (N_11452,N_7457,N_7196);
nand U11453 (N_11453,N_6411,N_7624);
nor U11454 (N_11454,N_6669,N_7648);
nor U11455 (N_11455,N_7759,N_8924);
xnor U11456 (N_11456,N_7891,N_6927);
xnor U11457 (N_11457,N_7524,N_7702);
nor U11458 (N_11458,N_8057,N_8417);
nor U11459 (N_11459,N_6808,N_7595);
and U11460 (N_11460,N_6627,N_8685);
and U11461 (N_11461,N_6387,N_6348);
or U11462 (N_11462,N_8441,N_7144);
nor U11463 (N_11463,N_6559,N_7325);
xor U11464 (N_11464,N_8832,N_6890);
or U11465 (N_11465,N_7121,N_6726);
or U11466 (N_11466,N_8860,N_8558);
nor U11467 (N_11467,N_8803,N_6019);
xor U11468 (N_11468,N_7230,N_7337);
or U11469 (N_11469,N_7017,N_6543);
or U11470 (N_11470,N_6744,N_8568);
xnor U11471 (N_11471,N_7973,N_8007);
nand U11472 (N_11472,N_8028,N_6723);
and U11473 (N_11473,N_6811,N_6573);
xnor U11474 (N_11474,N_6839,N_8203);
and U11475 (N_11475,N_8929,N_8446);
xor U11476 (N_11476,N_8907,N_7993);
or U11477 (N_11477,N_6561,N_7493);
and U11478 (N_11478,N_6777,N_7781);
or U11479 (N_11479,N_8954,N_6066);
or U11480 (N_11480,N_7171,N_6543);
and U11481 (N_11481,N_7756,N_8511);
nand U11482 (N_11482,N_6486,N_7197);
or U11483 (N_11483,N_7991,N_6910);
nor U11484 (N_11484,N_8955,N_7460);
nand U11485 (N_11485,N_8532,N_7659);
xor U11486 (N_11486,N_6564,N_8267);
and U11487 (N_11487,N_8371,N_6822);
and U11488 (N_11488,N_7828,N_6312);
nor U11489 (N_11489,N_8399,N_8590);
xor U11490 (N_11490,N_6339,N_8737);
nor U11491 (N_11491,N_7809,N_7482);
xor U11492 (N_11492,N_7908,N_8732);
and U11493 (N_11493,N_8130,N_6096);
and U11494 (N_11494,N_6419,N_6609);
nand U11495 (N_11495,N_7006,N_6027);
nand U11496 (N_11496,N_7917,N_8939);
and U11497 (N_11497,N_8581,N_8088);
xnor U11498 (N_11498,N_6884,N_6701);
nand U11499 (N_11499,N_6187,N_6735);
xnor U11500 (N_11500,N_8773,N_7348);
nand U11501 (N_11501,N_8660,N_8532);
and U11502 (N_11502,N_6047,N_6605);
nor U11503 (N_11503,N_7284,N_8913);
and U11504 (N_11504,N_8271,N_8338);
xnor U11505 (N_11505,N_8377,N_7354);
nor U11506 (N_11506,N_7504,N_7643);
nand U11507 (N_11507,N_6192,N_8877);
and U11508 (N_11508,N_6397,N_7292);
or U11509 (N_11509,N_8063,N_7913);
xnor U11510 (N_11510,N_8700,N_6892);
xnor U11511 (N_11511,N_6516,N_8006);
or U11512 (N_11512,N_7481,N_8375);
xor U11513 (N_11513,N_6657,N_6014);
nor U11514 (N_11514,N_8876,N_7085);
nor U11515 (N_11515,N_8729,N_8423);
and U11516 (N_11516,N_6867,N_8690);
nand U11517 (N_11517,N_6524,N_8582);
nor U11518 (N_11518,N_8691,N_6674);
or U11519 (N_11519,N_6137,N_6828);
nor U11520 (N_11520,N_6714,N_6374);
nand U11521 (N_11521,N_8881,N_7543);
xor U11522 (N_11522,N_8181,N_7416);
nand U11523 (N_11523,N_6715,N_8436);
xor U11524 (N_11524,N_6046,N_8624);
xor U11525 (N_11525,N_8962,N_7528);
or U11526 (N_11526,N_8019,N_8308);
nand U11527 (N_11527,N_8657,N_7722);
nor U11528 (N_11528,N_6580,N_8157);
nand U11529 (N_11529,N_8668,N_6376);
nand U11530 (N_11530,N_7903,N_7665);
nand U11531 (N_11531,N_6401,N_7829);
xnor U11532 (N_11532,N_8007,N_7658);
nor U11533 (N_11533,N_7992,N_8257);
nor U11534 (N_11534,N_7850,N_8440);
and U11535 (N_11535,N_6897,N_6252);
nand U11536 (N_11536,N_6995,N_7175);
nand U11537 (N_11537,N_8175,N_8230);
xor U11538 (N_11538,N_7760,N_7356);
xor U11539 (N_11539,N_8857,N_7920);
nor U11540 (N_11540,N_8175,N_7571);
nand U11541 (N_11541,N_6231,N_6542);
and U11542 (N_11542,N_6438,N_8300);
and U11543 (N_11543,N_8272,N_8193);
xor U11544 (N_11544,N_8655,N_6118);
nand U11545 (N_11545,N_8329,N_6715);
or U11546 (N_11546,N_8171,N_8349);
or U11547 (N_11547,N_8499,N_7129);
or U11548 (N_11548,N_6446,N_7548);
nor U11549 (N_11549,N_8022,N_8537);
nor U11550 (N_11550,N_7285,N_8118);
nand U11551 (N_11551,N_8421,N_7811);
and U11552 (N_11552,N_6836,N_8190);
nand U11553 (N_11553,N_8462,N_8731);
and U11554 (N_11554,N_8586,N_8410);
or U11555 (N_11555,N_7966,N_7113);
nand U11556 (N_11556,N_8125,N_7939);
nand U11557 (N_11557,N_6231,N_7425);
xnor U11558 (N_11558,N_6388,N_6638);
nor U11559 (N_11559,N_7435,N_6370);
nand U11560 (N_11560,N_8702,N_6516);
xor U11561 (N_11561,N_7342,N_6565);
nor U11562 (N_11562,N_7385,N_8096);
nand U11563 (N_11563,N_6960,N_6996);
nand U11564 (N_11564,N_8435,N_7975);
and U11565 (N_11565,N_6165,N_7268);
or U11566 (N_11566,N_6879,N_7866);
or U11567 (N_11567,N_6919,N_6305);
xnor U11568 (N_11568,N_8529,N_8931);
xor U11569 (N_11569,N_7846,N_7180);
or U11570 (N_11570,N_8244,N_6790);
and U11571 (N_11571,N_8526,N_8884);
or U11572 (N_11572,N_8407,N_8681);
nor U11573 (N_11573,N_7537,N_7458);
or U11574 (N_11574,N_7335,N_7042);
or U11575 (N_11575,N_7374,N_6035);
xor U11576 (N_11576,N_8218,N_6055);
nor U11577 (N_11577,N_8964,N_6982);
nor U11578 (N_11578,N_8240,N_7043);
nand U11579 (N_11579,N_6099,N_8877);
or U11580 (N_11580,N_8360,N_6914);
xor U11581 (N_11581,N_8255,N_6995);
nand U11582 (N_11582,N_8515,N_6361);
nor U11583 (N_11583,N_7340,N_8205);
nor U11584 (N_11584,N_7673,N_6745);
and U11585 (N_11585,N_6027,N_6215);
nor U11586 (N_11586,N_7007,N_8527);
nor U11587 (N_11587,N_6875,N_8905);
or U11588 (N_11588,N_8871,N_6978);
and U11589 (N_11589,N_8073,N_7358);
nor U11590 (N_11590,N_8615,N_6853);
nor U11591 (N_11591,N_7749,N_8340);
and U11592 (N_11592,N_7144,N_7648);
nand U11593 (N_11593,N_6186,N_6151);
xor U11594 (N_11594,N_6501,N_8162);
and U11595 (N_11595,N_6570,N_7957);
xnor U11596 (N_11596,N_6689,N_8759);
nor U11597 (N_11597,N_7572,N_7930);
nand U11598 (N_11598,N_6074,N_8586);
nand U11599 (N_11599,N_8561,N_6532);
or U11600 (N_11600,N_6166,N_6681);
nand U11601 (N_11601,N_8984,N_8734);
xnor U11602 (N_11602,N_7359,N_8681);
xor U11603 (N_11603,N_7431,N_7784);
xnor U11604 (N_11604,N_6939,N_7239);
nand U11605 (N_11605,N_6417,N_8770);
nand U11606 (N_11606,N_8610,N_7482);
or U11607 (N_11607,N_6348,N_6951);
xor U11608 (N_11608,N_7087,N_6620);
nor U11609 (N_11609,N_6661,N_8761);
nand U11610 (N_11610,N_6847,N_6431);
nand U11611 (N_11611,N_6209,N_8516);
nor U11612 (N_11612,N_8564,N_6575);
or U11613 (N_11613,N_6129,N_6284);
or U11614 (N_11614,N_7562,N_6937);
or U11615 (N_11615,N_6312,N_7580);
or U11616 (N_11616,N_6632,N_7658);
or U11617 (N_11617,N_7050,N_8676);
or U11618 (N_11618,N_7635,N_6175);
xnor U11619 (N_11619,N_7788,N_8037);
nand U11620 (N_11620,N_6708,N_8745);
nor U11621 (N_11621,N_6011,N_8663);
nand U11622 (N_11622,N_7756,N_6813);
xor U11623 (N_11623,N_6328,N_6390);
or U11624 (N_11624,N_7419,N_8671);
nor U11625 (N_11625,N_6926,N_8281);
or U11626 (N_11626,N_7448,N_7506);
xnor U11627 (N_11627,N_8487,N_6604);
xnor U11628 (N_11628,N_8913,N_8709);
nand U11629 (N_11629,N_6591,N_6040);
nor U11630 (N_11630,N_6162,N_7155);
or U11631 (N_11631,N_7112,N_6280);
xor U11632 (N_11632,N_8137,N_6920);
or U11633 (N_11633,N_8722,N_6830);
xor U11634 (N_11634,N_8098,N_7483);
or U11635 (N_11635,N_7575,N_6848);
and U11636 (N_11636,N_8173,N_8783);
xnor U11637 (N_11637,N_7828,N_6071);
or U11638 (N_11638,N_8558,N_7859);
nor U11639 (N_11639,N_8935,N_6058);
nand U11640 (N_11640,N_6272,N_7044);
and U11641 (N_11641,N_6601,N_6232);
xor U11642 (N_11642,N_7969,N_8532);
nor U11643 (N_11643,N_6198,N_6172);
and U11644 (N_11644,N_8314,N_6912);
nand U11645 (N_11645,N_8858,N_6764);
nor U11646 (N_11646,N_8152,N_7374);
and U11647 (N_11647,N_6492,N_8954);
or U11648 (N_11648,N_7209,N_6949);
and U11649 (N_11649,N_6047,N_7899);
nand U11650 (N_11650,N_8643,N_7315);
nand U11651 (N_11651,N_8513,N_6968);
nand U11652 (N_11652,N_8715,N_7783);
nor U11653 (N_11653,N_6157,N_7758);
or U11654 (N_11654,N_8052,N_8420);
nor U11655 (N_11655,N_7191,N_7280);
and U11656 (N_11656,N_6938,N_7481);
nor U11657 (N_11657,N_7165,N_6826);
xor U11658 (N_11658,N_8053,N_6229);
and U11659 (N_11659,N_8719,N_6257);
xnor U11660 (N_11660,N_8229,N_6377);
and U11661 (N_11661,N_8430,N_6082);
xor U11662 (N_11662,N_8684,N_8266);
or U11663 (N_11663,N_7461,N_8883);
nand U11664 (N_11664,N_6005,N_7574);
xnor U11665 (N_11665,N_6729,N_8505);
nand U11666 (N_11666,N_6930,N_7482);
nor U11667 (N_11667,N_8536,N_8806);
xnor U11668 (N_11668,N_7417,N_7827);
xor U11669 (N_11669,N_8292,N_6373);
nor U11670 (N_11670,N_8498,N_7660);
nand U11671 (N_11671,N_7724,N_6253);
nor U11672 (N_11672,N_7921,N_7059);
nand U11673 (N_11673,N_6215,N_8418);
xnor U11674 (N_11674,N_6005,N_8859);
xor U11675 (N_11675,N_7488,N_6530);
or U11676 (N_11676,N_6901,N_8704);
nand U11677 (N_11677,N_6843,N_7270);
xor U11678 (N_11678,N_6874,N_7938);
or U11679 (N_11679,N_6398,N_6142);
nor U11680 (N_11680,N_7606,N_7711);
nand U11681 (N_11681,N_6798,N_8072);
xnor U11682 (N_11682,N_8545,N_6089);
nand U11683 (N_11683,N_8827,N_6640);
nand U11684 (N_11684,N_7509,N_7457);
or U11685 (N_11685,N_6074,N_6763);
nand U11686 (N_11686,N_7367,N_8432);
or U11687 (N_11687,N_7319,N_7596);
nor U11688 (N_11688,N_6616,N_8227);
nand U11689 (N_11689,N_7742,N_8905);
xnor U11690 (N_11690,N_7864,N_8996);
nand U11691 (N_11691,N_7897,N_7438);
nor U11692 (N_11692,N_6456,N_7013);
or U11693 (N_11693,N_7410,N_6375);
xnor U11694 (N_11694,N_6640,N_7735);
or U11695 (N_11695,N_8428,N_8691);
or U11696 (N_11696,N_6115,N_6562);
and U11697 (N_11697,N_8792,N_8967);
xnor U11698 (N_11698,N_7033,N_6029);
or U11699 (N_11699,N_8860,N_7743);
and U11700 (N_11700,N_6043,N_8962);
nor U11701 (N_11701,N_7677,N_8535);
nor U11702 (N_11702,N_7108,N_6562);
or U11703 (N_11703,N_7893,N_6653);
or U11704 (N_11704,N_8967,N_6717);
nor U11705 (N_11705,N_8470,N_6026);
nor U11706 (N_11706,N_6185,N_8911);
and U11707 (N_11707,N_7560,N_7734);
xnor U11708 (N_11708,N_6829,N_7415);
nand U11709 (N_11709,N_6673,N_8151);
or U11710 (N_11710,N_6202,N_8819);
xnor U11711 (N_11711,N_6204,N_8676);
and U11712 (N_11712,N_6632,N_8761);
nor U11713 (N_11713,N_6562,N_8900);
and U11714 (N_11714,N_7658,N_6079);
and U11715 (N_11715,N_8917,N_6060);
nor U11716 (N_11716,N_7617,N_7305);
or U11717 (N_11717,N_8887,N_7236);
nor U11718 (N_11718,N_7882,N_8591);
xor U11719 (N_11719,N_8850,N_6208);
or U11720 (N_11720,N_8339,N_6893);
or U11721 (N_11721,N_7341,N_7558);
nand U11722 (N_11722,N_8979,N_8488);
or U11723 (N_11723,N_7957,N_7633);
or U11724 (N_11724,N_8477,N_6332);
nor U11725 (N_11725,N_8337,N_7858);
and U11726 (N_11726,N_8928,N_8942);
nand U11727 (N_11727,N_8551,N_8210);
nand U11728 (N_11728,N_7951,N_6094);
nor U11729 (N_11729,N_8616,N_7649);
nor U11730 (N_11730,N_6351,N_6377);
nor U11731 (N_11731,N_7190,N_8480);
xor U11732 (N_11732,N_8521,N_7112);
and U11733 (N_11733,N_6518,N_6198);
xor U11734 (N_11734,N_6043,N_8047);
xnor U11735 (N_11735,N_7656,N_6076);
and U11736 (N_11736,N_8510,N_7369);
nand U11737 (N_11737,N_6383,N_6660);
nand U11738 (N_11738,N_8977,N_7473);
nand U11739 (N_11739,N_6630,N_8923);
nor U11740 (N_11740,N_8099,N_7463);
nor U11741 (N_11741,N_6673,N_8370);
xor U11742 (N_11742,N_7089,N_8411);
nor U11743 (N_11743,N_8929,N_8711);
and U11744 (N_11744,N_6257,N_7231);
or U11745 (N_11745,N_8379,N_7650);
nand U11746 (N_11746,N_7623,N_6645);
nand U11747 (N_11747,N_6371,N_6195);
nor U11748 (N_11748,N_7213,N_7444);
nor U11749 (N_11749,N_7458,N_8110);
nor U11750 (N_11750,N_7233,N_7926);
nand U11751 (N_11751,N_6571,N_8250);
or U11752 (N_11752,N_6640,N_8023);
nor U11753 (N_11753,N_6321,N_6283);
and U11754 (N_11754,N_6124,N_7199);
nor U11755 (N_11755,N_8024,N_6504);
xnor U11756 (N_11756,N_7925,N_7743);
xor U11757 (N_11757,N_8850,N_6568);
or U11758 (N_11758,N_8024,N_6114);
or U11759 (N_11759,N_6265,N_7198);
or U11760 (N_11760,N_6175,N_8498);
nand U11761 (N_11761,N_7112,N_8997);
xor U11762 (N_11762,N_7762,N_7498);
and U11763 (N_11763,N_6053,N_8630);
and U11764 (N_11764,N_7977,N_8220);
nor U11765 (N_11765,N_7498,N_7705);
nand U11766 (N_11766,N_8987,N_7815);
and U11767 (N_11767,N_7876,N_8991);
or U11768 (N_11768,N_6597,N_6981);
xor U11769 (N_11769,N_6857,N_7457);
nand U11770 (N_11770,N_7206,N_6340);
or U11771 (N_11771,N_8002,N_7701);
and U11772 (N_11772,N_8660,N_7488);
xor U11773 (N_11773,N_7630,N_6059);
nand U11774 (N_11774,N_6935,N_7308);
nand U11775 (N_11775,N_7345,N_6438);
nor U11776 (N_11776,N_7228,N_7073);
nor U11777 (N_11777,N_6098,N_7404);
xnor U11778 (N_11778,N_6490,N_7202);
nand U11779 (N_11779,N_6344,N_7227);
nor U11780 (N_11780,N_6941,N_7339);
and U11781 (N_11781,N_8764,N_8954);
nand U11782 (N_11782,N_6692,N_8399);
and U11783 (N_11783,N_6085,N_8701);
xnor U11784 (N_11784,N_7003,N_6934);
nor U11785 (N_11785,N_8983,N_7183);
and U11786 (N_11786,N_6112,N_7853);
nand U11787 (N_11787,N_7659,N_8267);
nand U11788 (N_11788,N_6281,N_6907);
nor U11789 (N_11789,N_7979,N_8969);
and U11790 (N_11790,N_7962,N_7693);
or U11791 (N_11791,N_6213,N_8927);
xnor U11792 (N_11792,N_6407,N_8479);
xor U11793 (N_11793,N_8023,N_7759);
xor U11794 (N_11794,N_8749,N_8630);
nand U11795 (N_11795,N_7198,N_8518);
nand U11796 (N_11796,N_8501,N_6833);
or U11797 (N_11797,N_6089,N_6821);
xnor U11798 (N_11798,N_8387,N_7488);
xnor U11799 (N_11799,N_7182,N_8777);
xnor U11800 (N_11800,N_7061,N_8722);
and U11801 (N_11801,N_8277,N_8072);
or U11802 (N_11802,N_7839,N_6540);
xnor U11803 (N_11803,N_8061,N_6951);
nor U11804 (N_11804,N_6672,N_6432);
and U11805 (N_11805,N_7007,N_8013);
nand U11806 (N_11806,N_8831,N_6241);
xnor U11807 (N_11807,N_7194,N_8106);
or U11808 (N_11808,N_7134,N_7973);
nand U11809 (N_11809,N_7712,N_7639);
nor U11810 (N_11810,N_7379,N_6973);
nor U11811 (N_11811,N_8400,N_6860);
xor U11812 (N_11812,N_7856,N_7258);
xor U11813 (N_11813,N_7419,N_7482);
nand U11814 (N_11814,N_6545,N_6095);
and U11815 (N_11815,N_6393,N_8848);
or U11816 (N_11816,N_6760,N_6857);
and U11817 (N_11817,N_8111,N_8922);
and U11818 (N_11818,N_7424,N_6559);
or U11819 (N_11819,N_6733,N_8887);
nor U11820 (N_11820,N_7847,N_7674);
nand U11821 (N_11821,N_6497,N_8929);
and U11822 (N_11822,N_6827,N_6841);
xor U11823 (N_11823,N_8221,N_7604);
or U11824 (N_11824,N_7021,N_6520);
or U11825 (N_11825,N_8781,N_7911);
nand U11826 (N_11826,N_7202,N_7260);
and U11827 (N_11827,N_8338,N_8804);
and U11828 (N_11828,N_7633,N_6337);
xor U11829 (N_11829,N_6130,N_7479);
nand U11830 (N_11830,N_8043,N_6650);
nand U11831 (N_11831,N_8984,N_8147);
nand U11832 (N_11832,N_7956,N_6707);
nor U11833 (N_11833,N_8444,N_7549);
nor U11834 (N_11834,N_8157,N_6514);
or U11835 (N_11835,N_8545,N_8569);
and U11836 (N_11836,N_8809,N_7205);
nand U11837 (N_11837,N_6750,N_6356);
nor U11838 (N_11838,N_8923,N_8686);
nor U11839 (N_11839,N_8712,N_7846);
nand U11840 (N_11840,N_6325,N_8745);
or U11841 (N_11841,N_6838,N_7466);
xor U11842 (N_11842,N_6225,N_8897);
nor U11843 (N_11843,N_8210,N_6731);
nor U11844 (N_11844,N_6123,N_8413);
nand U11845 (N_11845,N_6672,N_7474);
or U11846 (N_11846,N_6795,N_6957);
nand U11847 (N_11847,N_7990,N_8637);
nand U11848 (N_11848,N_7092,N_6616);
nor U11849 (N_11849,N_6435,N_6458);
or U11850 (N_11850,N_8946,N_6056);
and U11851 (N_11851,N_6749,N_6546);
and U11852 (N_11852,N_7403,N_7202);
nand U11853 (N_11853,N_8389,N_7698);
nor U11854 (N_11854,N_7020,N_7503);
nor U11855 (N_11855,N_7998,N_7439);
xor U11856 (N_11856,N_6985,N_6324);
xor U11857 (N_11857,N_6588,N_7867);
nand U11858 (N_11858,N_8758,N_6900);
and U11859 (N_11859,N_6199,N_6178);
xnor U11860 (N_11860,N_6356,N_7736);
and U11861 (N_11861,N_8352,N_7841);
xnor U11862 (N_11862,N_7525,N_7092);
nand U11863 (N_11863,N_7293,N_7039);
or U11864 (N_11864,N_7080,N_7361);
and U11865 (N_11865,N_6673,N_7753);
or U11866 (N_11866,N_7810,N_7336);
nor U11867 (N_11867,N_8080,N_6205);
or U11868 (N_11868,N_7103,N_6240);
and U11869 (N_11869,N_8864,N_6990);
or U11870 (N_11870,N_7425,N_7811);
nor U11871 (N_11871,N_6262,N_8000);
and U11872 (N_11872,N_8946,N_7117);
and U11873 (N_11873,N_7960,N_8216);
nor U11874 (N_11874,N_6575,N_8188);
xor U11875 (N_11875,N_7642,N_6714);
xor U11876 (N_11876,N_6194,N_6143);
nand U11877 (N_11877,N_8848,N_7086);
nand U11878 (N_11878,N_7613,N_8650);
or U11879 (N_11879,N_8045,N_8675);
nor U11880 (N_11880,N_8597,N_7369);
xnor U11881 (N_11881,N_6620,N_8857);
and U11882 (N_11882,N_6508,N_7915);
xor U11883 (N_11883,N_6244,N_6556);
and U11884 (N_11884,N_7494,N_6073);
and U11885 (N_11885,N_8929,N_8642);
nand U11886 (N_11886,N_8976,N_6842);
xor U11887 (N_11887,N_7701,N_8427);
nor U11888 (N_11888,N_6006,N_7378);
or U11889 (N_11889,N_7498,N_8613);
or U11890 (N_11890,N_8871,N_8486);
and U11891 (N_11891,N_6268,N_8242);
nand U11892 (N_11892,N_8553,N_7365);
nor U11893 (N_11893,N_8981,N_6256);
and U11894 (N_11894,N_6699,N_8929);
and U11895 (N_11895,N_6017,N_6891);
and U11896 (N_11896,N_6129,N_6114);
xnor U11897 (N_11897,N_8404,N_8760);
or U11898 (N_11898,N_8415,N_7285);
nor U11899 (N_11899,N_6156,N_8056);
and U11900 (N_11900,N_8972,N_6034);
xnor U11901 (N_11901,N_8286,N_6629);
nand U11902 (N_11902,N_6197,N_6077);
xor U11903 (N_11903,N_7754,N_7696);
xnor U11904 (N_11904,N_8322,N_7809);
or U11905 (N_11905,N_8898,N_7102);
or U11906 (N_11906,N_8492,N_7054);
nor U11907 (N_11907,N_6099,N_8185);
nand U11908 (N_11908,N_7417,N_6046);
or U11909 (N_11909,N_6470,N_7978);
or U11910 (N_11910,N_8374,N_6284);
and U11911 (N_11911,N_6966,N_6038);
xnor U11912 (N_11912,N_6955,N_7273);
or U11913 (N_11913,N_6020,N_8149);
nand U11914 (N_11914,N_6157,N_7772);
nand U11915 (N_11915,N_7157,N_6386);
or U11916 (N_11916,N_8679,N_7704);
nor U11917 (N_11917,N_6865,N_6235);
nand U11918 (N_11918,N_8321,N_6693);
xnor U11919 (N_11919,N_6271,N_7870);
and U11920 (N_11920,N_8843,N_7895);
and U11921 (N_11921,N_7675,N_8782);
or U11922 (N_11922,N_7107,N_6068);
and U11923 (N_11923,N_8398,N_8007);
and U11924 (N_11924,N_6339,N_8113);
nand U11925 (N_11925,N_7448,N_6489);
nand U11926 (N_11926,N_6588,N_8517);
xor U11927 (N_11927,N_7853,N_7289);
or U11928 (N_11928,N_7681,N_7929);
xnor U11929 (N_11929,N_7861,N_8039);
and U11930 (N_11930,N_6390,N_7527);
nand U11931 (N_11931,N_7654,N_8479);
nand U11932 (N_11932,N_7125,N_7298);
xor U11933 (N_11933,N_8435,N_7777);
nor U11934 (N_11934,N_6812,N_6786);
xnor U11935 (N_11935,N_8654,N_7707);
nand U11936 (N_11936,N_7178,N_6683);
nand U11937 (N_11937,N_6033,N_7285);
nor U11938 (N_11938,N_6388,N_7658);
xor U11939 (N_11939,N_6965,N_7589);
xnor U11940 (N_11940,N_7838,N_6126);
xor U11941 (N_11941,N_8932,N_6586);
and U11942 (N_11942,N_8022,N_8850);
nand U11943 (N_11943,N_8636,N_6038);
xor U11944 (N_11944,N_6156,N_8695);
or U11945 (N_11945,N_7828,N_8917);
and U11946 (N_11946,N_7233,N_8577);
nor U11947 (N_11947,N_6792,N_7675);
and U11948 (N_11948,N_8716,N_8447);
xnor U11949 (N_11949,N_8308,N_6697);
xnor U11950 (N_11950,N_8039,N_6192);
or U11951 (N_11951,N_7425,N_8150);
nor U11952 (N_11952,N_8361,N_6252);
or U11953 (N_11953,N_6951,N_6636);
nand U11954 (N_11954,N_7413,N_6840);
nor U11955 (N_11955,N_6326,N_6294);
xnor U11956 (N_11956,N_7616,N_6792);
xor U11957 (N_11957,N_8824,N_8678);
nand U11958 (N_11958,N_6294,N_8589);
nand U11959 (N_11959,N_6269,N_7878);
or U11960 (N_11960,N_6416,N_7746);
nand U11961 (N_11961,N_6035,N_6960);
nand U11962 (N_11962,N_8062,N_8842);
or U11963 (N_11963,N_7738,N_7286);
and U11964 (N_11964,N_7064,N_7884);
and U11965 (N_11965,N_6737,N_6081);
nor U11966 (N_11966,N_8544,N_6720);
and U11967 (N_11967,N_7270,N_7110);
or U11968 (N_11968,N_6485,N_7432);
xor U11969 (N_11969,N_8481,N_6091);
and U11970 (N_11970,N_6512,N_7597);
or U11971 (N_11971,N_6059,N_8544);
nand U11972 (N_11972,N_8309,N_6149);
xor U11973 (N_11973,N_7185,N_8237);
nand U11974 (N_11974,N_8923,N_8576);
nor U11975 (N_11975,N_6638,N_6512);
or U11976 (N_11976,N_6033,N_8572);
or U11977 (N_11977,N_6142,N_6377);
or U11978 (N_11978,N_8546,N_6909);
nand U11979 (N_11979,N_7304,N_6188);
nor U11980 (N_11980,N_7774,N_7607);
nor U11981 (N_11981,N_8102,N_7617);
nor U11982 (N_11982,N_8032,N_6589);
xor U11983 (N_11983,N_7234,N_7444);
nand U11984 (N_11984,N_8525,N_7835);
xnor U11985 (N_11985,N_7834,N_7024);
nand U11986 (N_11986,N_7663,N_7051);
or U11987 (N_11987,N_7753,N_6538);
xor U11988 (N_11988,N_7085,N_7448);
and U11989 (N_11989,N_6082,N_8577);
nor U11990 (N_11990,N_7790,N_8952);
or U11991 (N_11991,N_7407,N_8264);
nand U11992 (N_11992,N_7695,N_6720);
nor U11993 (N_11993,N_8908,N_6742);
nor U11994 (N_11994,N_7594,N_8516);
and U11995 (N_11995,N_7628,N_6013);
xnor U11996 (N_11996,N_6145,N_6601);
xor U11997 (N_11997,N_6497,N_8093);
nor U11998 (N_11998,N_8169,N_6324);
and U11999 (N_11999,N_7421,N_7253);
or U12000 (N_12000,N_11826,N_11659);
nand U12001 (N_12001,N_10630,N_10152);
or U12002 (N_12002,N_10284,N_9676);
or U12003 (N_12003,N_10210,N_10260);
nand U12004 (N_12004,N_10746,N_10449);
nand U12005 (N_12005,N_10215,N_9493);
nor U12006 (N_12006,N_11249,N_11097);
and U12007 (N_12007,N_11535,N_10920);
and U12008 (N_12008,N_9634,N_9480);
nor U12009 (N_12009,N_9958,N_9193);
nand U12010 (N_12010,N_10151,N_9766);
and U12011 (N_12011,N_11503,N_9035);
xor U12012 (N_12012,N_9448,N_10939);
xnor U12013 (N_12013,N_10039,N_9464);
xnor U12014 (N_12014,N_9862,N_9875);
nor U12015 (N_12015,N_10744,N_10809);
nand U12016 (N_12016,N_10280,N_11466);
and U12017 (N_12017,N_11305,N_10701);
and U12018 (N_12018,N_9787,N_9533);
nand U12019 (N_12019,N_9824,N_11151);
xnor U12020 (N_12020,N_11206,N_9739);
nor U12021 (N_12021,N_11464,N_11759);
nand U12022 (N_12022,N_9281,N_11079);
or U12023 (N_12023,N_10930,N_11121);
xnor U12024 (N_12024,N_9165,N_11420);
or U12025 (N_12025,N_10826,N_10241);
and U12026 (N_12026,N_10243,N_10803);
nand U12027 (N_12027,N_10897,N_9659);
xor U12028 (N_12028,N_10177,N_9941);
nor U12029 (N_12029,N_9428,N_9772);
nand U12030 (N_12030,N_10383,N_9934);
or U12031 (N_12031,N_9065,N_10410);
nor U12032 (N_12032,N_10504,N_10348);
nor U12033 (N_12033,N_9970,N_11601);
nand U12034 (N_12034,N_10121,N_11877);
or U12035 (N_12035,N_9172,N_10714);
nor U12036 (N_12036,N_9138,N_9842);
and U12037 (N_12037,N_9455,N_11895);
or U12038 (N_12038,N_11513,N_9123);
nand U12039 (N_12039,N_10153,N_10176);
xnor U12040 (N_12040,N_11239,N_11606);
xor U12041 (N_12041,N_11525,N_9411);
xor U12042 (N_12042,N_9174,N_11125);
and U12043 (N_12043,N_9328,N_10211);
or U12044 (N_12044,N_10567,N_10428);
and U12045 (N_12045,N_10984,N_9154);
nor U12046 (N_12046,N_9628,N_10108);
or U12047 (N_12047,N_9277,N_9614);
and U12048 (N_12048,N_9967,N_9056);
nand U12049 (N_12049,N_11011,N_9732);
nand U12050 (N_12050,N_11709,N_10943);
and U12051 (N_12051,N_11959,N_11120);
xor U12052 (N_12052,N_11123,N_11428);
and U12053 (N_12053,N_9489,N_11894);
nor U12054 (N_12054,N_9609,N_11431);
and U12055 (N_12055,N_11155,N_10040);
and U12056 (N_12056,N_11360,N_10795);
and U12057 (N_12057,N_11716,N_11068);
xnor U12058 (N_12058,N_10435,N_9948);
xor U12059 (N_12059,N_9519,N_9048);
nand U12060 (N_12060,N_11507,N_10288);
nand U12061 (N_12061,N_9517,N_9271);
nor U12062 (N_12062,N_10534,N_11396);
or U12063 (N_12063,N_11113,N_9479);
and U12064 (N_12064,N_10818,N_9134);
xnor U12065 (N_12065,N_10952,N_9699);
and U12066 (N_12066,N_11622,N_9837);
nor U12067 (N_12067,N_10379,N_10069);
nor U12068 (N_12068,N_10485,N_11742);
or U12069 (N_12069,N_11336,N_9522);
xnor U12070 (N_12070,N_9831,N_10450);
or U12071 (N_12071,N_11806,N_10443);
nand U12072 (N_12072,N_11133,N_11695);
or U12073 (N_12073,N_9832,N_10753);
xnor U12074 (N_12074,N_10910,N_10513);
and U12075 (N_12075,N_10345,N_9598);
nor U12076 (N_12076,N_10518,N_10692);
and U12077 (N_12077,N_9949,N_10834);
xor U12078 (N_12078,N_9327,N_10408);
and U12079 (N_12079,N_9213,N_10465);
nor U12080 (N_12080,N_9765,N_11276);
and U12081 (N_12081,N_9496,N_10591);
nor U12082 (N_12082,N_10977,N_10095);
nand U12083 (N_12083,N_11588,N_10166);
xnor U12084 (N_12084,N_11673,N_10104);
nor U12085 (N_12085,N_11519,N_10311);
nor U12086 (N_12086,N_11354,N_11453);
or U12087 (N_12087,N_11975,N_11812);
xor U12088 (N_12088,N_9243,N_9266);
and U12089 (N_12089,N_10271,N_10578);
and U12090 (N_12090,N_9656,N_10643);
and U12091 (N_12091,N_10261,N_10906);
nor U12092 (N_12092,N_9442,N_10232);
and U12093 (N_12093,N_11551,N_9801);
nand U12094 (N_12094,N_9137,N_10283);
nand U12095 (N_12095,N_11747,N_11544);
or U12096 (N_12096,N_10392,N_11470);
xnor U12097 (N_12097,N_9023,N_10937);
nor U12098 (N_12098,N_11033,N_9576);
xor U12099 (N_12099,N_11433,N_9346);
or U12100 (N_12100,N_11928,N_9921);
and U12101 (N_12101,N_11815,N_9369);
and U12102 (N_12102,N_10594,N_11979);
or U12103 (N_12103,N_10031,N_10880);
nor U12104 (N_12104,N_9190,N_10606);
nor U12105 (N_12105,N_9977,N_9552);
xnor U12106 (N_12106,N_11728,N_10479);
or U12107 (N_12107,N_10003,N_9555);
and U12108 (N_12108,N_9582,N_9405);
and U12109 (N_12109,N_11614,N_11108);
nor U12110 (N_12110,N_10086,N_10498);
xor U12111 (N_12111,N_9904,N_11858);
nand U12112 (N_12112,N_9413,N_11740);
or U12113 (N_12113,N_11139,N_10777);
nand U12114 (N_12114,N_11722,N_9878);
and U12115 (N_12115,N_10884,N_10586);
nand U12116 (N_12116,N_11825,N_9159);
nand U12117 (N_12117,N_10360,N_9458);
or U12118 (N_12118,N_9141,N_9201);
and U12119 (N_12119,N_9913,N_11445);
or U12120 (N_12120,N_10363,N_10709);
nor U12121 (N_12121,N_11110,N_10853);
and U12122 (N_12122,N_9839,N_9096);
xor U12123 (N_12123,N_10509,N_10660);
nor U12124 (N_12124,N_11390,N_9286);
xor U12125 (N_12125,N_9537,N_10782);
xor U12126 (N_12126,N_10446,N_11328);
nor U12127 (N_12127,N_9619,N_9241);
or U12128 (N_12128,N_11945,N_11363);
nand U12129 (N_12129,N_11048,N_9392);
or U12130 (N_12130,N_11751,N_9214);
nand U12131 (N_12131,N_11577,N_11212);
nor U12132 (N_12132,N_11765,N_10342);
and U12133 (N_12133,N_11261,N_10366);
and U12134 (N_12134,N_9362,N_11972);
and U12135 (N_12135,N_11412,N_10116);
or U12136 (N_12136,N_11392,N_9916);
nor U12137 (N_12137,N_9347,N_10061);
nor U12138 (N_12138,N_9974,N_11042);
and U12139 (N_12139,N_10830,N_10090);
xor U12140 (N_12140,N_9162,N_10564);
xnor U12141 (N_12141,N_11809,N_9407);
or U12142 (N_12142,N_11312,N_10332);
and U12143 (N_12143,N_9014,N_9982);
or U12144 (N_12144,N_11834,N_10973);
and U12145 (N_12145,N_9210,N_11738);
or U12146 (N_12146,N_10060,N_10367);
xnor U12147 (N_12147,N_10337,N_11065);
nand U12148 (N_12148,N_10820,N_9639);
or U12149 (N_12149,N_11521,N_10255);
nor U12150 (N_12150,N_11849,N_10601);
and U12151 (N_12151,N_9888,N_9964);
nor U12152 (N_12152,N_11088,N_9804);
nor U12153 (N_12153,N_9185,N_11313);
and U12154 (N_12154,N_10636,N_11938);
xor U12155 (N_12155,N_11447,N_9840);
nand U12156 (N_12156,N_10511,N_10480);
nor U12157 (N_12157,N_10323,N_10272);
or U12158 (N_12158,N_9384,N_9494);
xnor U12159 (N_12159,N_11002,N_10196);
xor U12160 (N_12160,N_11656,N_11511);
and U12161 (N_12161,N_9693,N_9754);
or U12162 (N_12162,N_11529,N_9044);
xor U12163 (N_12163,N_10793,N_9993);
or U12164 (N_12164,N_11753,N_10142);
nand U12165 (N_12165,N_11892,N_10565);
and U12166 (N_12166,N_11773,N_11457);
xor U12167 (N_12167,N_11666,N_10021);
or U12168 (N_12168,N_9939,N_9655);
xor U12169 (N_12169,N_9567,N_10277);
xor U12170 (N_12170,N_10224,N_11427);
nor U12171 (N_12171,N_9503,N_10481);
or U12172 (N_12172,N_9780,N_9730);
xor U12173 (N_12173,N_11735,N_10571);
nand U12174 (N_12174,N_9223,N_9991);
and U12175 (N_12175,N_10494,N_9870);
nor U12176 (N_12176,N_9534,N_9924);
xor U12177 (N_12177,N_11395,N_9254);
or U12178 (N_12178,N_9120,N_11402);
nor U12179 (N_12179,N_10862,N_9922);
or U12180 (N_12180,N_9771,N_10599);
xor U12181 (N_12181,N_9351,N_11718);
nand U12182 (N_12182,N_11438,N_11271);
nor U12183 (N_12183,N_9729,N_10524);
nand U12184 (N_12184,N_11164,N_10497);
nor U12185 (N_12185,N_9128,N_9985);
nor U12186 (N_12186,N_11282,N_9475);
and U12187 (N_12187,N_9572,N_11407);
nand U12188 (N_12188,N_9690,N_10429);
nor U12189 (N_12189,N_11855,N_10874);
nor U12190 (N_12190,N_9219,N_9244);
or U12191 (N_12191,N_9393,N_9653);
nor U12192 (N_12192,N_9389,N_11217);
xnor U12193 (N_12193,N_11626,N_9390);
nand U12194 (N_12194,N_10851,N_10091);
and U12195 (N_12195,N_10233,N_9456);
xnor U12196 (N_12196,N_10197,N_11550);
xor U12197 (N_12197,N_10759,N_9333);
or U12198 (N_12198,N_9177,N_10893);
and U12199 (N_12199,N_9672,N_10161);
nor U12200 (N_12200,N_11910,N_10626);
or U12201 (N_12201,N_11440,N_9060);
xnor U12202 (N_12202,N_11421,N_9476);
and U12203 (N_12203,N_10106,N_9615);
nor U12204 (N_12204,N_10129,N_11852);
xnor U12205 (N_12205,N_9097,N_10434);
nand U12206 (N_12206,N_10831,N_9148);
or U12207 (N_12207,N_10922,N_11838);
nor U12208 (N_12208,N_9115,N_10929);
nand U12209 (N_12209,N_11029,N_11311);
nand U12210 (N_12210,N_11671,N_9980);
or U12211 (N_12211,N_11708,N_9136);
xnor U12212 (N_12212,N_11099,N_10604);
nor U12213 (N_12213,N_10837,N_11701);
xnor U12214 (N_12214,N_11302,N_9835);
or U12215 (N_12215,N_9554,N_10926);
nor U12216 (N_12216,N_9258,N_10122);
nor U12217 (N_12217,N_10781,N_9834);
xor U12218 (N_12218,N_10967,N_11231);
or U12219 (N_12219,N_10775,N_9003);
and U12220 (N_12220,N_9529,N_10209);
nor U12221 (N_12221,N_10466,N_9481);
nor U12222 (N_12222,N_10841,N_9121);
nor U12223 (N_12223,N_10708,N_9047);
xor U12224 (N_12224,N_10011,N_9221);
xor U12225 (N_12225,N_9220,N_11814);
xnor U12226 (N_12226,N_9045,N_9767);
and U12227 (N_12227,N_9830,N_9228);
nand U12228 (N_12228,N_9813,N_9415);
and U12229 (N_12229,N_9043,N_9378);
xor U12230 (N_12230,N_9100,N_11300);
xnor U12231 (N_12231,N_11679,N_11787);
xnor U12232 (N_12232,N_9911,N_9098);
nor U12233 (N_12233,N_11208,N_10621);
nor U12234 (N_12234,N_9033,N_10115);
xor U12235 (N_12235,N_11982,N_11129);
nand U12236 (N_12236,N_9288,N_11946);
xnor U12237 (N_12237,N_10340,N_10027);
nand U12238 (N_12238,N_10216,N_9426);
and U12239 (N_12239,N_11497,N_9709);
nand U12240 (N_12240,N_11411,N_10240);
nor U12241 (N_12241,N_10319,N_11677);
or U12242 (N_12242,N_9790,N_10117);
nor U12243 (N_12243,N_9737,N_9617);
nor U12244 (N_12244,N_9250,N_9486);
nand U12245 (N_12245,N_9714,N_11038);
nand U12246 (N_12246,N_10290,N_10310);
xnor U12247 (N_12247,N_11788,N_10084);
nor U12248 (N_12248,N_10928,N_10105);
or U12249 (N_12249,N_11181,N_10038);
xnor U12250 (N_12250,N_11926,N_9026);
and U12251 (N_12251,N_10451,N_9838);
or U12252 (N_12252,N_11031,N_9589);
nand U12253 (N_12253,N_11253,N_10155);
xnor U12254 (N_12254,N_10935,N_9302);
nor U12255 (N_12255,N_11278,N_10220);
nor U12256 (N_12256,N_11114,N_9158);
xor U12257 (N_12257,N_9414,N_9160);
or U12258 (N_12258,N_9526,N_10032);
nor U12259 (N_12259,N_9110,N_10526);
nand U12260 (N_12260,N_11797,N_10532);
and U12261 (N_12261,N_11487,N_10322);
nand U12262 (N_12262,N_11488,N_10373);
or U12263 (N_12263,N_11291,N_9133);
or U12264 (N_12264,N_10458,N_10048);
and U12265 (N_12265,N_11280,N_11929);
nor U12266 (N_12266,N_11066,N_10415);
or U12267 (N_12267,N_9925,N_10710);
and U12268 (N_12268,N_9039,N_11010);
nand U12269 (N_12269,N_10720,N_10202);
xnor U12270 (N_12270,N_11732,N_11856);
xnor U12271 (N_12271,N_11973,N_9126);
or U12272 (N_12272,N_10163,N_9200);
and U12273 (N_12273,N_11260,N_11839);
xor U12274 (N_12274,N_10572,N_9037);
and U12275 (N_12275,N_11911,N_11352);
nand U12276 (N_12276,N_9109,N_9350);
nand U12277 (N_12277,N_11351,N_11172);
or U12278 (N_12278,N_11180,N_10448);
nand U12279 (N_12279,N_10993,N_10418);
or U12280 (N_12280,N_11760,N_9553);
nand U12281 (N_12281,N_10258,N_9451);
and U12282 (N_12282,N_11772,N_9587);
xnor U12283 (N_12283,N_11854,N_10832);
or U12284 (N_12284,N_10522,N_9020);
and U12285 (N_12285,N_10971,N_9966);
nor U12286 (N_12286,N_10279,N_10386);
nor U12287 (N_12287,N_11451,N_10649);
or U12288 (N_12288,N_11049,N_10346);
and U12289 (N_12289,N_11865,N_10833);
nand U12290 (N_12290,N_11537,N_11991);
nand U12291 (N_12291,N_9650,N_9192);
nor U12292 (N_12292,N_10352,N_11640);
xor U12293 (N_12293,N_11192,N_11866);
nand U12294 (N_12294,N_10245,N_10905);
and U12295 (N_12295,N_10476,N_9682);
or U12296 (N_12296,N_10114,N_9802);
nand U12297 (N_12297,N_9793,N_9929);
or U12298 (N_12298,N_10724,N_9152);
or U12299 (N_12299,N_11861,N_10460);
or U12300 (N_12300,N_9275,N_9425);
nor U12301 (N_12301,N_11661,N_11920);
nor U12302 (N_12302,N_9111,N_11102);
or U12303 (N_12303,N_11623,N_9444);
xor U12304 (N_12304,N_11279,N_9488);
and U12305 (N_12305,N_11736,N_9140);
xnor U12306 (N_12306,N_11974,N_9570);
nand U12307 (N_12307,N_11694,N_11900);
or U12308 (N_12308,N_11409,N_9910);
nand U12309 (N_12309,N_9508,N_9686);
or U12310 (N_12310,N_9588,N_11915);
or U12311 (N_12311,N_10972,N_11962);
and U12312 (N_12312,N_11729,N_9968);
or U12313 (N_12313,N_10653,N_11800);
nand U12314 (N_12314,N_10043,N_10925);
nor U12315 (N_12315,N_10535,N_10149);
nand U12316 (N_12316,N_10719,N_10400);
and U12317 (N_12317,N_11194,N_10944);
nand U12318 (N_12318,N_9715,N_10885);
or U12319 (N_12319,N_11064,N_11932);
or U12320 (N_12320,N_11107,N_9976);
nand U12321 (N_12321,N_10530,N_11980);
xnor U12322 (N_12322,N_11881,N_9706);
nand U12323 (N_12323,N_11597,N_9417);
nand U12324 (N_12324,N_11315,N_9914);
xnor U12325 (N_12325,N_9147,N_9516);
xor U12326 (N_12326,N_9996,N_11145);
or U12327 (N_12327,N_11128,N_9107);
nand U12328 (N_12328,N_9592,N_10894);
and U12329 (N_12329,N_10983,N_9283);
or U12330 (N_12330,N_10250,N_10338);
nand U12331 (N_12331,N_11157,N_11171);
or U12332 (N_12332,N_9256,N_9196);
nor U12333 (N_12333,N_9376,N_9375);
xnor U12334 (N_12334,N_10026,N_9669);
or U12335 (N_12335,N_10406,N_10327);
nor U12336 (N_12336,N_10193,N_10585);
nand U12337 (N_12337,N_9294,N_9989);
or U12338 (N_12338,N_11184,N_10609);
nor U12339 (N_12339,N_10637,N_10743);
nand U12340 (N_12340,N_10171,N_10769);
nor U12341 (N_12341,N_10459,N_9101);
xnor U12342 (N_12342,N_11222,N_9209);
nand U12343 (N_12343,N_11922,N_11940);
or U12344 (N_12344,N_9525,N_11480);
and U12345 (N_12345,N_11976,N_9226);
nand U12346 (N_12346,N_11482,N_10145);
xor U12347 (N_12347,N_9090,N_9885);
nand U12348 (N_12348,N_10073,N_11745);
or U12349 (N_12349,N_11889,N_10797);
xnor U12350 (N_12350,N_9527,N_10558);
nand U12351 (N_12351,N_10707,N_10413);
nand U12352 (N_12352,N_10072,N_10221);
nor U12353 (N_12353,N_11501,N_9088);
xor U12354 (N_12354,N_11292,N_11681);
or U12355 (N_12355,N_11560,N_10788);
and U12356 (N_12356,N_10750,N_9153);
nor U12357 (N_12357,N_9861,N_9603);
xnor U12358 (N_12358,N_10128,N_10907);
and U12359 (N_12359,N_11754,N_9716);
or U12360 (N_12360,N_11628,N_11785);
or U12361 (N_12361,N_9318,N_10886);
nand U12362 (N_12362,N_9829,N_11868);
and U12363 (N_12363,N_11131,N_9726);
nand U12364 (N_12364,N_9300,N_9398);
or U12365 (N_12365,N_11909,N_11741);
or U12366 (N_12366,N_9282,N_9343);
or U12367 (N_12367,N_9947,N_10563);
and U12368 (N_12368,N_11397,N_11688);
and U12369 (N_12369,N_10824,N_11624);
or U12370 (N_12370,N_9595,N_10985);
nand U12371 (N_12371,N_9719,N_9573);
or U12372 (N_12372,N_11651,N_9658);
nor U12373 (N_12373,N_9314,N_10351);
and U12374 (N_12374,N_9819,N_11720);
or U12375 (N_12375,N_10628,N_11565);
and U12376 (N_12376,N_9748,N_11933);
nor U12377 (N_12377,N_10908,N_10454);
xnor U12378 (N_12378,N_9180,N_10561);
or U12379 (N_12379,N_10890,N_10773);
xnor U12380 (N_12380,N_9704,N_9942);
and U12381 (N_12381,N_9216,N_10792);
nor U12382 (N_12382,N_11805,N_11674);
xnor U12383 (N_12383,N_9701,N_10470);
xor U12384 (N_12384,N_11256,N_11885);
nand U12385 (N_12385,N_11968,N_11845);
xor U12386 (N_12386,N_11725,N_10732);
nor U12387 (N_12387,N_9296,N_10722);
or U12388 (N_12388,N_9954,N_9249);
xor U12389 (N_12389,N_11642,N_10186);
nor U12390 (N_12390,N_9015,N_9053);
xor U12391 (N_12391,N_11268,N_11224);
nor U12392 (N_12392,N_11032,N_9577);
and U12393 (N_12393,N_11000,N_10647);
or U12394 (N_12394,N_10307,N_10262);
or U12395 (N_12395,N_10817,N_10184);
nor U12396 (N_12396,N_11724,N_9436);
nor U12397 (N_12397,N_11755,N_11020);
nand U12398 (N_12398,N_10941,N_9259);
nor U12399 (N_12399,N_11243,N_10137);
nand U12400 (N_12400,N_9773,N_10768);
xnor U12401 (N_12401,N_9886,N_10417);
and U12402 (N_12402,N_11017,N_10127);
and U12403 (N_12403,N_10344,N_10306);
or U12404 (N_12404,N_9688,N_11116);
or U12405 (N_12405,N_10350,N_11890);
xor U12406 (N_12406,N_11027,N_11886);
xnor U12407 (N_12407,N_9364,N_10546);
xnor U12408 (N_12408,N_11204,N_11442);
and U12409 (N_12409,N_9342,N_9708);
nor U12410 (N_12410,N_10491,N_11448);
nand U12411 (N_12411,N_10595,N_9791);
nand U12412 (N_12412,N_9085,N_11439);
nand U12413 (N_12413,N_11454,N_10389);
or U12414 (N_12414,N_11326,N_10318);
nand U12415 (N_12415,N_11556,N_9074);
xor U12416 (N_12416,N_9437,N_9331);
nand U12417 (N_12417,N_10754,N_10704);
and U12418 (N_12418,N_9736,N_11616);
or U12419 (N_12419,N_11430,N_9827);
or U12420 (N_12420,N_9454,N_9010);
nand U12421 (N_12421,N_11167,N_10807);
and U12422 (N_12422,N_11713,N_11201);
nand U12423 (N_12423,N_9545,N_11615);
xor U12424 (N_12424,N_11879,N_10191);
and U12425 (N_12425,N_9877,N_9575);
nor U12426 (N_12426,N_10829,N_11388);
xnor U12427 (N_12427,N_11853,N_10499);
nor U12428 (N_12428,N_10543,N_10783);
nand U12429 (N_12429,N_11563,N_9368);
xnor U12430 (N_12430,N_9002,N_10471);
nor U12431 (N_12431,N_10355,N_11211);
xnor U12432 (N_12432,N_11075,N_10314);
xor U12433 (N_12433,N_11764,N_9155);
nor U12434 (N_12434,N_9051,N_10811);
nor U12435 (N_12435,N_11637,N_10251);
xor U12436 (N_12436,N_10836,N_9181);
nor U12437 (N_12437,N_10638,N_11477);
and U12438 (N_12438,N_9361,N_11953);
and U12439 (N_12439,N_9170,N_9021);
or U12440 (N_12440,N_9551,N_11189);
nand U12441 (N_12441,N_9975,N_11534);
nand U12442 (N_12442,N_11119,N_9093);
and U12443 (N_12443,N_11964,N_10916);
and U12444 (N_12444,N_9559,N_11061);
xor U12445 (N_12445,N_9779,N_10388);
and U12446 (N_12446,N_10876,N_10253);
and U12447 (N_12447,N_9943,N_9741);
or U12448 (N_12448,N_11818,N_9262);
nor U12449 (N_12449,N_11548,N_11594);
nand U12450 (N_12450,N_10645,N_9463);
nor U12451 (N_12451,N_9652,N_10422);
and U12452 (N_12452,N_11983,N_9700);
xor U12453 (N_12453,N_10822,N_11491);
nor U12454 (N_12454,N_10650,N_10778);
nand U12455 (N_12455,N_10713,N_10292);
nand U12456 (N_12456,N_11489,N_10933);
nor U12457 (N_12457,N_10957,N_9285);
nor U12458 (N_12458,N_11101,N_9776);
or U12459 (N_12459,N_10335,N_9124);
nor U12460 (N_12460,N_9016,N_10663);
or U12461 (N_12461,N_10597,N_10964);
xor U12462 (N_12462,N_11531,N_10462);
and U12463 (N_12463,N_9354,N_11739);
nand U12464 (N_12464,N_10089,N_11481);
and U12465 (N_12465,N_10521,N_9338);
or U12466 (N_12466,N_11219,N_11875);
nor U12467 (N_12467,N_10452,N_11842);
xor U12468 (N_12468,N_9915,N_9011);
nand U12469 (N_12469,N_10045,N_10705);
and U12470 (N_12470,N_11903,N_11483);
nor U12471 (N_12471,N_11987,N_11723);
nand U12472 (N_12472,N_11419,N_10730);
and U12473 (N_12473,N_10206,N_10050);
nor U12474 (N_12474,N_9636,N_11174);
or U12475 (N_12475,N_10402,N_9206);
or U12476 (N_12476,N_10256,N_9335);
nor U12477 (N_12477,N_11930,N_9290);
xor U12478 (N_12478,N_11160,N_9562);
nand U12479 (N_12479,N_10900,N_9883);
or U12480 (N_12480,N_11314,N_10304);
nand U12481 (N_12481,N_10102,N_10533);
nand U12482 (N_12482,N_9853,N_10828);
and U12483 (N_12483,N_10602,N_11404);
nor U12484 (N_12484,N_10079,N_9590);
and U12485 (N_12485,N_10016,N_9815);
or U12486 (N_12486,N_10537,N_11069);
and U12487 (N_12487,N_10784,N_11578);
nand U12488 (N_12488,N_10486,N_11761);
nor U12489 (N_12489,N_11286,N_11752);
nor U12490 (N_12490,N_11105,N_10684);
nand U12491 (N_12491,N_9151,N_10583);
nand U12492 (N_12492,N_11091,N_10124);
and U12493 (N_12493,N_11337,N_10286);
or U12494 (N_12494,N_11465,N_9222);
xor U12495 (N_12495,N_10912,N_11690);
nand U12496 (N_12496,N_11316,N_11634);
and U12497 (N_12497,N_11093,N_9070);
nor U12498 (N_12498,N_10000,N_11562);
nor U12499 (N_12499,N_9960,N_11663);
nor U12500 (N_12500,N_11244,N_11939);
nor U12501 (N_12501,N_10655,N_11523);
and U12502 (N_12502,N_10349,N_9322);
nor U12503 (N_12503,N_11324,N_9786);
nand U12504 (N_12504,N_10331,N_10468);
nand U12505 (N_12505,N_9440,N_10679);
and U12506 (N_12506,N_9449,N_11142);
and U12507 (N_12507,N_10855,N_11100);
nand U12508 (N_12508,N_10844,N_11413);
nor U12509 (N_12509,N_11520,N_10150);
or U12510 (N_12510,N_10440,N_10461);
xor U12511 (N_12511,N_11115,N_10640);
or U12512 (N_12512,N_9040,N_9891);
nand U12513 (N_12513,N_11587,N_10892);
xor U12514 (N_12514,N_10845,N_10875);
nand U12515 (N_12515,N_9784,N_11334);
nand U12516 (N_12516,N_9498,N_9145);
and U12517 (N_12517,N_9624,N_11387);
nand U12518 (N_12518,N_11287,N_10794);
or U12519 (N_12519,N_11643,N_9703);
nand U12520 (N_12520,N_10582,N_10819);
and U12521 (N_12521,N_10453,N_10510);
and U12522 (N_12522,N_10017,N_10394);
and U12523 (N_12523,N_11141,N_9410);
nand U12524 (N_12524,N_9324,N_9325);
xnor U12525 (N_12525,N_11092,N_9337);
and U12526 (N_12526,N_11467,N_10023);
nand U12527 (N_12527,N_10181,N_10806);
nand U12528 (N_12528,N_10222,N_10478);
and U12529 (N_12529,N_9232,N_9848);
nand U12530 (N_12530,N_10961,N_9462);
nor U12531 (N_12531,N_11799,N_11007);
xor U12532 (N_12532,N_10988,N_9971);
xor U12533 (N_12533,N_9998,N_9025);
xor U12534 (N_12534,N_10545,N_11175);
xnor U12535 (N_12535,N_10588,N_10175);
and U12536 (N_12536,N_10096,N_11087);
and U12537 (N_12537,N_9594,N_11508);
and U12538 (N_12538,N_11382,N_11076);
and U12539 (N_12539,N_11476,N_10172);
or U12540 (N_12540,N_9675,N_11796);
nand U12541 (N_12541,N_9550,N_9050);
or U12542 (N_12542,N_11285,N_9186);
xor U12543 (N_12543,N_11509,N_10396);
nand U12544 (N_12544,N_11486,N_11494);
and U12545 (N_12545,N_9168,N_10173);
or U12546 (N_12546,N_11455,N_10702);
nand U12547 (N_12547,N_11824,N_10044);
and U12548 (N_12548,N_10416,N_10752);
nand U12549 (N_12549,N_10259,N_9321);
xor U12550 (N_12550,N_11934,N_11044);
xnor U12551 (N_12551,N_9549,N_10347);
nand U12552 (N_12552,N_11984,N_10870);
and U12553 (N_12553,N_9358,N_9586);
nand U12554 (N_12554,N_10358,N_10542);
and U12555 (N_12555,N_9388,N_11234);
or U12556 (N_12556,N_11542,N_11051);
xor U12557 (N_12557,N_11422,N_9933);
nor U12558 (N_12558,N_11275,N_9189);
or U12559 (N_12559,N_9890,N_9651);
or U12560 (N_12560,N_9316,N_9308);
xnor U12561 (N_12561,N_10412,N_11530);
and U12562 (N_12562,N_11492,N_9505);
or U12563 (N_12563,N_11380,N_10536);
nand U12564 (N_12564,N_9692,N_9593);
and U12565 (N_12565,N_11216,N_9291);
nor U12566 (N_12566,N_11257,N_11775);
and U12567 (N_12567,N_10118,N_10200);
and U12568 (N_12568,N_10728,N_11490);
or U12569 (N_12569,N_9674,N_9064);
xnor U12570 (N_12570,N_9513,N_10924);
and U12571 (N_12571,N_11857,N_11552);
or U12572 (N_12572,N_11955,N_11122);
and U12573 (N_12573,N_9520,N_10147);
nand U12574 (N_12574,N_9645,N_11908);
or U12575 (N_12575,N_11098,N_10278);
nor U12576 (N_12576,N_11398,N_10382);
xor U12577 (N_12577,N_11235,N_11887);
nand U12578 (N_12578,N_11379,N_9252);
nand U12579 (N_12579,N_11630,N_9265);
or U12580 (N_12580,N_11913,N_10742);
xnor U12581 (N_12581,N_10860,N_10691);
nand U12582 (N_12582,N_11472,N_11232);
or U12583 (N_12583,N_10927,N_11377);
and U12584 (N_12584,N_11689,N_11176);
nor U12585 (N_12585,N_11954,N_11109);
or U12586 (N_12586,N_10958,N_10827);
nor U12587 (N_12587,N_10188,N_11124);
nor U12588 (N_12588,N_10821,N_10953);
nand U12589 (N_12589,N_11266,N_9560);
and U12590 (N_12590,N_9860,N_11117);
xor U12591 (N_12591,N_9268,N_11776);
and U12592 (N_12592,N_9538,N_9150);
nor U12593 (N_12593,N_9778,N_9667);
xnor U12594 (N_12594,N_9666,N_11389);
or U12595 (N_12595,N_10087,N_9034);
or U12596 (N_12596,N_9429,N_9202);
nor U12597 (N_12597,N_9905,N_10441);
nand U12598 (N_12598,N_9122,N_10223);
and U12599 (N_12599,N_10432,N_11816);
nand U12600 (N_12600,N_10328,N_11575);
and U12601 (N_12601,N_10192,N_10505);
and U12602 (N_12602,N_11299,N_10519);
xnor U12603 (N_12603,N_10403,N_9713);
or U12604 (N_12604,N_11071,N_10881);
nand U12605 (N_12605,N_9903,N_9307);
nand U12606 (N_12606,N_11668,N_10948);
and U12607 (N_12607,N_11441,N_10528);
nand U12608 (N_12608,N_10407,N_11848);
or U12609 (N_12609,N_9530,N_9907);
nor U12610 (N_12610,N_10054,N_10774);
xor U12611 (N_12611,N_10131,N_9647);
nand U12612 (N_12612,N_10666,N_9404);
and U12613 (N_12613,N_9317,N_11158);
and U12614 (N_12614,N_11050,N_9642);
and U12615 (N_12615,N_10711,N_11780);
and U12616 (N_12616,N_10654,N_11641);
and U12617 (N_12617,N_10353,N_10887);
nor U12618 (N_12618,N_11949,N_11867);
nand U12619 (N_12619,N_10354,N_9919);
xnor U12620 (N_12620,N_10931,N_10789);
nor U12621 (N_12621,N_11744,N_9932);
and U12622 (N_12622,N_9760,N_11094);
nor U12623 (N_12623,N_10294,N_9365);
nand U12624 (N_12624,N_11469,N_11456);
or U12625 (N_12625,N_10718,N_9743);
or U12626 (N_12626,N_11468,N_9979);
or U12627 (N_12627,N_11250,N_10677);
and U12628 (N_12628,N_9755,N_10997);
xnor U12629 (N_12629,N_11332,N_10786);
xnor U12630 (N_12630,N_9662,N_9401);
nand U12631 (N_12631,N_9618,N_9930);
and U12632 (N_12632,N_10757,N_10664);
or U12633 (N_12633,N_11627,N_10648);
xor U12634 (N_12634,N_10978,N_9502);
xor U12635 (N_12635,N_9453,N_10285);
nand U12636 (N_12636,N_9341,N_9826);
nor U12637 (N_12637,N_11837,N_10488);
nand U12638 (N_12638,N_10093,N_9944);
nor U12639 (N_12639,N_11084,N_10838);
or U12640 (N_12640,N_11414,N_10492);
or U12641 (N_12641,N_10405,N_11341);
xnor U12642 (N_12642,N_10399,N_9972);
and U12643 (N_12643,N_10226,N_10436);
nor U12644 (N_12644,N_9142,N_10909);
nand U12645 (N_12645,N_11957,N_9299);
or U12646 (N_12646,N_9229,N_9038);
nor U12647 (N_12647,N_11645,N_10552);
nor U12648 (N_12648,N_10861,N_9443);
nor U12649 (N_12649,N_10143,N_11346);
and U12650 (N_12650,N_10735,N_10766);
nor U12651 (N_12651,N_11273,N_11524);
or U12652 (N_12652,N_9898,N_10848);
nor U12653 (N_12653,N_9777,N_11596);
nand U12654 (N_12654,N_10555,N_10556);
or U12655 (N_12655,N_11296,N_10484);
nand U12656 (N_12656,N_10266,N_11283);
xor U12657 (N_12657,N_11459,N_9908);
or U12658 (N_12658,N_10496,N_10316);
and U12659 (N_12659,N_11040,N_11304);
and U12660 (N_12660,N_11547,N_11177);
nand U12661 (N_12661,N_10991,N_10903);
xnor U12662 (N_12662,N_11710,N_10825);
or U12663 (N_12663,N_10740,N_10100);
nand U12664 (N_12664,N_10098,N_11026);
or U12665 (N_12665,N_10620,N_10165);
or U12666 (N_12666,N_10762,N_10125);
nand U12667 (N_12667,N_10404,N_11165);
xnor U12668 (N_12668,N_9018,N_9310);
xor U12669 (N_12669,N_9528,N_10992);
and U12670 (N_12670,N_11386,N_11185);
and U12671 (N_12671,N_11829,N_10658);
and U12672 (N_12672,N_9370,N_11698);
and U12673 (N_12673,N_9808,N_11168);
and U12674 (N_12674,N_9359,N_9195);
or U12675 (N_12675,N_11053,N_9889);
nand U12676 (N_12676,N_9108,N_10483);
and U12677 (N_12677,N_10639,N_9665);
nor U12678 (N_12678,N_9876,N_11549);
xor U12679 (N_12679,N_9211,N_10296);
and U12680 (N_12680,N_9873,N_11580);
nand U12681 (N_12681,N_9531,N_10423);
xor U12682 (N_12682,N_11872,N_11156);
or U12683 (N_12683,N_9167,N_11917);
nor U12684 (N_12684,N_10756,N_9470);
nor U12685 (N_12685,N_11602,N_10430);
xor U12686 (N_12686,N_10986,N_11541);
or U12687 (N_12687,N_10878,N_9649);
xnor U12688 (N_12688,N_10659,N_9366);
and U12689 (N_12689,N_11394,N_10447);
and U12690 (N_12690,N_11700,N_9733);
nand U12691 (N_12691,N_11325,N_11408);
and U12692 (N_12692,N_11417,N_10675);
and U12693 (N_12693,N_9984,N_11138);
and U12694 (N_12694,N_10678,N_11226);
or U12695 (N_12695,N_9233,N_11603);
or U12696 (N_12696,N_10864,N_9046);
nand U12697 (N_12697,N_11229,N_11670);
and U12698 (N_12698,N_11406,N_9856);
and U12699 (N_12699,N_10872,N_9248);
nor U12700 (N_12700,N_10433,N_9825);
nand U12701 (N_12701,N_9806,N_9371);
xnor U12702 (N_12702,N_9363,N_10025);
nor U12703 (N_12703,N_11358,N_10409);
nor U12704 (N_12704,N_10763,N_10761);
xor U12705 (N_12705,N_11654,N_9036);
nor U12706 (N_12706,N_11307,N_9812);
nor U12707 (N_12707,N_11308,N_10356);
nor U12708 (N_12708,N_9487,N_11986);
and U12709 (N_12709,N_9660,N_11415);
or U12710 (N_12710,N_11635,N_10071);
xnor U12711 (N_12711,N_9717,N_10162);
or U12712 (N_12712,N_10942,N_10624);
or U12713 (N_12713,N_9858,N_9601);
and U12714 (N_12714,N_10956,N_11111);
nor U12715 (N_12715,N_10041,N_10502);
xnor U12716 (N_12716,N_10075,N_11743);
xor U12717 (N_12717,N_11958,N_9605);
and U12718 (N_12718,N_11687,N_9083);
or U12719 (N_12719,N_11749,N_11070);
nand U12720 (N_12720,N_10889,N_9467);
and U12721 (N_12721,N_9257,N_9521);
nor U12722 (N_12722,N_10974,N_10281);
nor U12723 (N_12723,N_9408,N_11237);
nand U12724 (N_12724,N_9608,N_11018);
and U12725 (N_12725,N_9353,N_10566);
or U12726 (N_12726,N_10092,N_10954);
or U12727 (N_12727,N_11182,N_9260);
xor U12728 (N_12728,N_10932,N_11786);
nand U12729 (N_12729,N_10074,N_10013);
xnor U12730 (N_12730,N_11766,N_10110);
nand U12731 (N_12731,N_9632,N_11485);
nor U12732 (N_12732,N_10330,N_11272);
and U12733 (N_12733,N_9828,N_10703);
xnor U12734 (N_12734,N_9146,N_10879);
or U12735 (N_12735,N_9817,N_11149);
nor U12736 (N_12736,N_10036,N_11610);
or U12737 (N_12737,N_9852,N_11188);
xnor U12738 (N_12738,N_10275,N_9198);
nand U12739 (N_12739,N_11543,N_11789);
or U12740 (N_12740,N_9240,N_9057);
nor U12741 (N_12741,N_9783,N_11532);
nand U12742 (N_12742,N_11166,N_9591);
xor U12743 (N_12743,N_9239,N_10273);
nand U12744 (N_12744,N_11331,N_10099);
or U12745 (N_12745,N_11479,N_9373);
nor U12746 (N_12746,N_10427,N_9616);
xnor U12747 (N_12747,N_11238,N_11609);
nor U12748 (N_12748,N_10252,N_11540);
and U12749 (N_12749,N_10706,N_9293);
or U12750 (N_12750,N_9657,N_9377);
xor U12751 (N_12751,N_10847,N_10264);
or U12752 (N_12752,N_10951,N_10815);
nand U12753 (N_12753,N_11003,N_11289);
xor U12754 (N_12754,N_9006,N_9497);
or U12755 (N_12755,N_10805,N_11103);
or U12756 (N_12756,N_10088,N_11576);
nor U12757 (N_12757,N_10899,N_11618);
nor U12758 (N_12758,N_9215,N_10608);
and U12759 (N_12759,N_11638,N_11134);
xor U12760 (N_12760,N_10945,N_10593);
or U12761 (N_12761,N_11383,N_9431);
nor U12762 (N_12762,N_9807,N_11221);
nand U12763 (N_12763,N_9116,N_9999);
xor U12764 (N_12764,N_11662,N_11223);
or U12765 (N_12765,N_11436,N_10798);
xnor U12766 (N_12766,N_11777,N_11330);
or U12767 (N_12767,N_9871,N_10646);
xnor U12768 (N_12768,N_9851,N_9751);
nor U12769 (N_12769,N_9009,N_11696);
nor U12770 (N_12770,N_10141,N_10005);
xnor U12771 (N_12771,N_10551,N_11712);
or U12772 (N_12772,N_9380,N_9013);
or U12773 (N_12773,N_11161,N_11948);
or U12774 (N_12774,N_11592,N_10070);
nor U12775 (N_12775,N_10577,N_9585);
nor U12776 (N_12776,N_9329,N_11526);
or U12777 (N_12777,N_10693,N_10493);
and U12778 (N_12778,N_11863,N_10934);
nor U12779 (N_12779,N_10438,N_10859);
nor U12780 (N_12780,N_11778,N_10377);
nand U12781 (N_12781,N_10607,N_11263);
or U12782 (N_12782,N_9086,N_11801);
nand U12783 (N_12783,N_9372,N_9792);
and U12784 (N_12784,N_9263,N_10842);
nor U12785 (N_12785,N_11950,N_9374);
nand U12786 (N_12786,N_11613,N_9445);
nor U12787 (N_12787,N_11034,N_10384);
nand U12788 (N_12788,N_9722,N_10187);
nand U12789 (N_12789,N_10758,N_11769);
and U12790 (N_12790,N_11931,N_9846);
or U12791 (N_12791,N_9119,N_9396);
nand U12792 (N_12792,N_9344,N_11078);
or U12793 (N_12793,N_10975,N_11370);
nand U12794 (N_12794,N_11147,N_10616);
and U12795 (N_12795,N_9187,N_9491);
nor U12796 (N_12796,N_11024,N_9078);
nand U12797 (N_12797,N_9809,N_10341);
xnor U12798 (N_12798,N_9602,N_11733);
or U12799 (N_12799,N_9957,N_9625);
nand U12800 (N_12800,N_10839,N_10295);
xor U12801 (N_12801,N_9450,N_9469);
or U12802 (N_12802,N_11269,N_10107);
xnor U12803 (N_12803,N_11301,N_10315);
xor U12804 (N_12804,N_10463,N_9612);
nor U12805 (N_12805,N_10083,N_10179);
xnor U12806 (N_12806,N_10712,N_9607);
nor U12807 (N_12807,N_10816,N_9543);
xnor U12808 (N_12808,N_10605,N_11495);
and U12809 (N_12809,N_9561,N_10507);
xor U12810 (N_12810,N_11350,N_11978);
xnor U12811 (N_12811,N_10868,N_11936);
and U12812 (N_12812,N_11607,N_11197);
or U12813 (N_12813,N_9477,N_9175);
nor U12814 (N_12814,N_9622,N_9633);
and U12815 (N_12815,N_9432,N_10301);
and U12816 (N_12816,N_11762,N_10725);
xor U12817 (N_12817,N_9897,N_9721);
nand U12818 (N_12818,N_11322,N_9067);
nand U12819 (N_12819,N_11475,N_11339);
and U12820 (N_12820,N_10164,N_11340);
nand U12821 (N_12821,N_9928,N_9556);
nor U12822 (N_12822,N_11774,N_11808);
and U12823 (N_12823,N_11233,N_10557);
nand U12824 (N_12824,N_11199,N_9412);
and U12825 (N_12825,N_11617,N_10671);
xnor U12826 (N_12826,N_9689,N_9680);
and U12827 (N_12827,N_10600,N_10568);
or U12828 (N_12828,N_9005,N_11822);
nand U12829 (N_12829,N_11236,N_10317);
nand U12830 (N_12830,N_11937,N_10030);
nor U12831 (N_12831,N_11012,N_11791);
or U12832 (N_12832,N_9072,N_10274);
nand U12833 (N_12833,N_10391,N_10042);
and U12834 (N_12834,N_9646,N_9000);
nor U12835 (N_12835,N_10802,N_10018);
nand U12836 (N_12836,N_10237,N_9125);
and U12837 (N_12837,N_11127,N_9424);
nand U12838 (N_12838,N_11393,N_9724);
or U12839 (N_12839,N_11359,N_10950);
nor U12840 (N_12840,N_11136,N_9422);
nand U12841 (N_12841,N_9161,N_11385);
xor U12842 (N_12842,N_9129,N_9874);
and U12843 (N_12843,N_10144,N_11990);
and U12844 (N_12844,N_11418,N_10661);
or U12845 (N_12845,N_10123,N_11633);
nand U12846 (N_12846,N_10850,N_11721);
nand U12847 (N_12847,N_11126,N_9557);
nand U12848 (N_12848,N_10508,N_9081);
xnor U12849 (N_12849,N_11081,N_9482);
or U12850 (N_12850,N_10590,N_11927);
or U12851 (N_12851,N_11361,N_11620);
nand U12852 (N_12852,N_10287,N_9075);
xnor U12853 (N_12853,N_11510,N_10631);
nand U12854 (N_12854,N_9001,N_10146);
nor U12855 (N_12855,N_10739,N_9637);
or U12856 (N_12856,N_10547,N_11281);
xnor U12857 (N_12857,N_9864,N_10982);
nand U12858 (N_12858,N_11502,N_10525);
nand U12859 (N_12859,N_10538,N_11112);
nand U12860 (N_12860,N_9238,N_11553);
nor U12861 (N_12861,N_9880,N_9761);
xor U12862 (N_12862,N_10883,N_10370);
xor U12863 (N_12863,N_9278,N_9113);
xor U12864 (N_12864,N_9710,N_9940);
or U12865 (N_12865,N_11657,N_9725);
nand U12866 (N_12866,N_9334,N_9963);
nor U12867 (N_12867,N_9077,N_11366);
or U12868 (N_12868,N_9952,N_9423);
nor U12869 (N_12869,N_9438,N_11255);
xnor U12870 (N_12870,N_9315,N_9759);
nor U12871 (N_12871,N_11461,N_11970);
or U12872 (N_12872,N_11163,N_11925);
xor U12873 (N_12873,N_11173,N_10615);
nand U12874 (N_12874,N_10130,N_9994);
or U12875 (N_12875,N_10873,N_10669);
or U12876 (N_12876,N_10665,N_10801);
or U12877 (N_12877,N_11897,N_9447);
nor U12878 (N_12878,N_9164,N_10549);
or U12879 (N_12879,N_9893,N_11568);
nor U12880 (N_12880,N_9049,N_10160);
and U12881 (N_12881,N_10056,N_10058);
and U12882 (N_12882,N_11218,N_11083);
nand U12883 (N_12883,N_10455,N_11985);
or U12884 (N_12884,N_11259,N_11817);
nor U12885 (N_12885,N_11783,N_9068);
or U12886 (N_12886,N_10562,N_11771);
nor U12887 (N_12887,N_11030,N_11499);
and U12888 (N_12888,N_11036,N_9309);
nand U12889 (N_12889,N_11921,N_9280);
nor U12890 (N_12890,N_11685,N_11557);
xnor U12891 (N_12891,N_9382,N_9623);
nor U12892 (N_12892,N_10047,N_10212);
xor U12893 (N_12893,N_11434,N_11023);
nand U12894 (N_12894,N_9188,N_11294);
xnor U12895 (N_12895,N_9978,N_9843);
nor U12896 (N_12896,N_11319,N_10913);
or U12897 (N_12897,N_11583,N_10183);
and U12898 (N_12898,N_11798,N_10246);
nor U12899 (N_12899,N_9894,N_11446);
or U12900 (N_12900,N_11170,N_11169);
or U12901 (N_12901,N_10305,N_11639);
nand U12902 (N_12902,N_11264,N_11016);
nand U12903 (N_12903,N_9409,N_9723);
nor U12904 (N_12904,N_10963,N_11367);
or U12905 (N_12905,N_9173,N_11584);
xnor U12906 (N_12906,N_11310,N_10263);
nor U12907 (N_12907,N_11647,N_9859);
or U12908 (N_12908,N_10915,N_9234);
xnor U12909 (N_12909,N_11591,N_10242);
nor U12910 (N_12910,N_10401,N_10244);
xnor U12911 (N_12911,N_11757,N_10359);
nor U12912 (N_12912,N_10472,N_10134);
nor U12913 (N_12913,N_9402,N_10230);
or U12914 (N_12914,N_11047,N_9292);
xnor U12915 (N_12915,N_10603,N_11850);
or U12916 (N_12916,N_10854,N_11137);
nor U12917 (N_12917,N_10840,N_9746);
nor U12918 (N_12918,N_10421,N_11058);
nand U12919 (N_12919,N_10297,N_9117);
nor U12920 (N_12920,N_11460,N_9684);
and U12921 (N_12921,N_9058,N_10729);
xor U12922 (N_12922,N_10437,N_11333);
xnor U12923 (N_12923,N_11833,N_9332);
nor U12924 (N_12924,N_11692,N_10190);
xor U12925 (N_12925,N_10898,N_10721);
nand U12926 (N_12926,N_10326,N_9785);
nand U12927 (N_12927,N_10747,N_9707);
nand U12928 (N_12928,N_11437,N_9069);
nand U12929 (N_12929,N_9313,N_11329);
or U12930 (N_12930,N_11284,N_9012);
nor U12931 (N_12931,N_9822,N_9135);
nor U12932 (N_12932,N_10309,N_10303);
xor U12933 (N_12933,N_9212,N_9892);
nor U12934 (N_12934,N_10634,N_10205);
xnor U12935 (N_12935,N_9157,N_9844);
nor U12936 (N_12936,N_10365,N_9242);
or U12937 (N_12937,N_11715,N_9604);
nand U12938 (N_12938,N_11348,N_10641);
nand U12939 (N_12939,N_10194,N_11598);
and U12940 (N_12940,N_10267,N_9330);
nor U12941 (N_12941,N_11251,N_10414);
or U12942 (N_12942,N_11924,N_11821);
xnor U12943 (N_12943,N_10687,N_11655);
or U12944 (N_12944,N_10014,N_10495);
nand U12945 (N_12945,N_10132,N_9774);
or U12946 (N_12946,N_10699,N_10550);
nor U12947 (N_12947,N_11621,N_9920);
nor U12948 (N_12948,N_9484,N_10895);
and U12949 (N_12949,N_9987,N_9246);
or U12950 (N_12950,N_11056,N_11009);
nand U12951 (N_12951,N_9360,N_9687);
xor U12952 (N_12952,N_10052,N_9568);
nor U12953 (N_12953,N_11449,N_11632);
and U12954 (N_12954,N_11146,N_10685);
nand U12955 (N_12955,N_10361,N_11942);
and U12956 (N_12956,N_9106,N_9019);
or U12957 (N_12957,N_10657,N_11574);
nand U12958 (N_12958,N_11343,N_11750);
and U12959 (N_12959,N_10651,N_9194);
or U12960 (N_12960,N_10683,N_11746);
nor U12961 (N_12961,N_10865,N_11148);
nand U12962 (N_12962,N_11375,N_11355);
nor U12963 (N_12963,N_11660,N_11870);
or U12964 (N_12964,N_11213,N_11579);
nor U12965 (N_12965,N_9251,N_10813);
nand U12966 (N_12966,N_11452,N_9718);
xor U12967 (N_12967,N_11365,N_10227);
nand U12968 (N_12968,N_11424,N_10808);
nor U12969 (N_12969,N_10320,N_10207);
nor U12970 (N_12970,N_10741,N_10779);
and U12971 (N_12971,N_11179,N_9394);
and U12972 (N_12972,N_10148,N_10919);
nand U12973 (N_12973,N_10994,N_11135);
nand U12974 (N_12974,N_10214,N_9055);
xnor U12975 (N_12975,N_10431,N_9564);
nand U12976 (N_12976,N_11429,N_10541);
nor U12977 (N_12977,N_11095,N_11132);
xor U12978 (N_12978,N_9901,N_9663);
nor U12979 (N_12979,N_9887,N_9797);
nor U12980 (N_12980,N_9823,N_11152);
nor U12981 (N_12981,N_10035,N_9740);
and U12982 (N_12982,N_9506,N_10823);
xor U12983 (N_12983,N_9127,N_9762);
nor U12984 (N_12984,N_10745,N_11242);
or U12985 (N_12985,N_11994,N_11399);
nor U12986 (N_12986,N_10888,N_9868);
nand U12987 (N_12987,N_9981,N_10420);
nor U12988 (N_12988,N_10667,N_10293);
and U12989 (N_12989,N_11193,N_11884);
and U12990 (N_12990,N_9540,N_10037);
nand U12991 (N_12991,N_11403,N_11060);
xor U12992 (N_12992,N_10034,N_9867);
nor U12993 (N_12993,N_10234,N_10723);
or U12994 (N_12994,N_9992,N_9547);
xnor U12995 (N_12995,N_9983,N_10612);
and U12996 (N_12996,N_10419,N_9406);
xor U12997 (N_12997,N_9004,N_10695);
xor U12998 (N_12998,N_10866,N_11888);
or U12999 (N_12999,N_10393,N_10467);
nand U13000 (N_13000,N_11041,N_10291);
or U13001 (N_13001,N_9176,N_9367);
or U13002 (N_13002,N_9945,N_9728);
or U13003 (N_13003,N_11344,N_10126);
or U13004 (N_13004,N_10208,N_10378);
or U13005 (N_13005,N_9092,N_10411);
nand U13006 (N_13006,N_9465,N_9918);
and U13007 (N_13007,N_11391,N_10066);
nand U13008 (N_13008,N_11074,N_9461);
and U13009 (N_13009,N_10727,N_9796);
xnor U13010 (N_13010,N_11650,N_10385);
nand U13011 (N_13011,N_9671,N_11515);
and U13012 (N_13012,N_9712,N_11790);
nand U13013 (N_13013,N_10046,N_11691);
and U13014 (N_13014,N_9143,N_10199);
nor U13015 (N_13015,N_9320,N_11611);
xnor U13016 (N_13016,N_11943,N_11090);
nor U13017 (N_13017,N_9895,N_9349);
and U13018 (N_13018,N_11306,N_9626);
nand U13019 (N_13019,N_11130,N_9356);
or U13020 (N_13020,N_11846,N_11793);
xor U13021 (N_13021,N_10268,N_11779);
nand U13022 (N_13022,N_9071,N_10053);
or U13023 (N_13023,N_11522,N_11426);
xor U13024 (N_13024,N_10529,N_10270);
nor U13025 (N_13025,N_11473,N_11435);
xnor U13026 (N_13026,N_11059,N_9799);
nor U13027 (N_13027,N_9841,N_11811);
nor U13028 (N_13028,N_10113,N_11768);
and U13029 (N_13029,N_9224,N_10457);
xnor U13030 (N_13030,N_9524,N_11089);
and U13031 (N_13031,N_9352,N_9566);
and U13032 (N_13032,N_11484,N_9457);
nor U13033 (N_13033,N_11295,N_9747);
nand U13034 (N_13034,N_10877,N_10501);
or U13035 (N_13035,N_9041,N_10500);
and U13036 (N_13036,N_9578,N_11252);
nand U13037 (N_13037,N_10357,N_9571);
or U13038 (N_13038,N_11203,N_9095);
xnor U13039 (N_13039,N_9357,N_11539);
xnor U13040 (N_13040,N_11841,N_9863);
nor U13041 (N_13041,N_9758,N_11086);
and U13042 (N_13042,N_10324,N_9511);
xor U13043 (N_13043,N_9512,N_10625);
xnor U13044 (N_13044,N_10236,N_11726);
xnor U13045 (N_13045,N_9912,N_9430);
and U13046 (N_13046,N_9416,N_9951);
nand U13047 (N_13047,N_10077,N_10313);
xnor U13048 (N_13048,N_11195,N_10229);
nor U13049 (N_13049,N_11080,N_9420);
xnor U13050 (N_13050,N_9836,N_11554);
nand U13051 (N_13051,N_9103,N_11559);
and U13052 (N_13052,N_10249,N_11669);
xor U13053 (N_13053,N_11254,N_11323);
or U13054 (N_13054,N_10523,N_11006);
and U13055 (N_13055,N_11923,N_10057);
or U13056 (N_13056,N_11734,N_10642);
nor U13057 (N_13057,N_10329,N_11590);
nor U13058 (N_13058,N_9931,N_10584);
and U13059 (N_13059,N_11571,N_9276);
or U13060 (N_13060,N_9460,N_11705);
nor U13061 (N_13061,N_10225,N_9483);
nand U13062 (N_13062,N_11907,N_11586);
and U13063 (N_13063,N_11246,N_10717);
nand U13064 (N_13064,N_10949,N_10955);
nor U13065 (N_13065,N_11005,N_11702);
xnor U13066 (N_13066,N_9811,N_10254);
nor U13067 (N_13067,N_9803,N_10863);
nor U13068 (N_13068,N_11104,N_9509);
nand U13069 (N_13069,N_10835,N_10103);
and U13070 (N_13070,N_11569,N_11247);
xor U13071 (N_13071,N_10914,N_9613);
nor U13072 (N_13072,N_9805,N_11327);
xor U13073 (N_13073,N_9621,N_11684);
or U13074 (N_13074,N_11293,N_11118);
nor U13075 (N_13075,N_9144,N_11697);
or U13076 (N_13076,N_9794,N_11187);
and U13077 (N_13077,N_9235,N_9678);
nand U13078 (N_13078,N_11450,N_9472);
and U13079 (N_13079,N_9548,N_11693);
nor U13080 (N_13080,N_11055,N_10213);
or U13081 (N_13081,N_11077,N_10474);
and U13082 (N_13082,N_11496,N_9400);
or U13083 (N_13083,N_10203,N_10780);
and U13084 (N_13084,N_9052,N_10397);
nor U13085 (N_13085,N_9355,N_10325);
xor U13086 (N_13086,N_11707,N_10901);
or U13087 (N_13087,N_10981,N_11996);
nand U13088 (N_13088,N_9927,N_11807);
and U13089 (N_13089,N_10078,N_10946);
nand U13090 (N_13090,N_11570,N_11008);
nor U13091 (N_13091,N_10015,N_10517);
or U13092 (N_13092,N_11400,N_9697);
nand U13093 (N_13093,N_9466,N_10623);
or U13094 (N_13094,N_10569,N_11912);
and U13095 (N_13095,N_9383,N_10334);
nor U13096 (N_13096,N_11999,N_9938);
xor U13097 (N_13097,N_11106,N_10867);
and U13098 (N_13098,N_9336,N_10520);
nand U13099 (N_13099,N_9814,N_10596);
nor U13100 (N_13100,N_9272,N_11859);
nand U13101 (N_13101,N_9536,N_9225);
xnor U13102 (N_13102,N_11368,N_10503);
nand U13103 (N_13103,N_9326,N_11150);
nand U13104 (N_13104,N_9742,N_9988);
or U13105 (N_13105,N_9900,N_9597);
nor U13106 (N_13106,N_11988,N_9702);
nand U13107 (N_13107,N_9565,N_10174);
or U13108 (N_13108,N_11599,N_10198);
nand U13109 (N_13109,N_10362,N_11941);
or U13110 (N_13110,N_11374,N_9184);
nand U13111 (N_13111,N_9935,N_10228);
and U13112 (N_13112,N_10751,N_9446);
and U13113 (N_13113,N_10081,N_9439);
or U13114 (N_13114,N_9094,N_10785);
nand U13115 (N_13115,N_11364,N_9541);
nor U13116 (N_13116,N_10911,N_10375);
nor U13117 (N_13117,N_9764,N_10598);
nand U13118 (N_13118,N_10475,N_11830);
nand U13119 (N_13119,N_9800,N_11462);
xnor U13120 (N_13120,N_11014,N_9599);
or U13121 (N_13121,N_9627,N_10575);
or U13122 (N_13122,N_10976,N_9950);
and U13123 (N_13123,N_10736,N_9105);
nand U13124 (N_13124,N_9166,N_9731);
or U13125 (N_13125,N_9923,N_11498);
or U13126 (N_13126,N_11564,N_11706);
nand U13127 (N_13127,N_11947,N_11956);
xor U13128 (N_13128,N_11369,N_9953);
xor U13129 (N_13129,N_10553,N_9149);
or U13130 (N_13130,N_10490,N_9029);
nand U13131 (N_13131,N_9218,N_11558);
nor U13132 (N_13132,N_11960,N_10726);
and U13133 (N_13133,N_10959,N_9112);
xor U13134 (N_13134,N_11085,N_9635);
or U13135 (N_13135,N_11274,N_9485);
nand U13136 (N_13136,N_9253,N_9763);
nand U13137 (N_13137,N_9066,N_11057);
xor U13138 (N_13138,N_11444,N_10843);
or U13139 (N_13139,N_10055,N_10204);
or U13140 (N_13140,N_9770,N_9881);
nand U13141 (N_13141,N_11664,N_9535);
nand U13142 (N_13142,N_11918,N_9705);
nand U13143 (N_13143,N_10686,N_10109);
nand U13144 (N_13144,N_10185,N_9087);
and U13145 (N_13145,N_11373,N_11648);
nand U13146 (N_13146,N_11649,N_9641);
or U13147 (N_13147,N_11416,N_11672);
or U13148 (N_13148,N_9217,N_9510);
nand U13149 (N_13149,N_9245,N_9171);
xor U13150 (N_13150,N_11504,N_10962);
or U13151 (N_13151,N_11880,N_10570);
xnor U13152 (N_13152,N_11993,N_10059);
and U13153 (N_13153,N_10219,N_9629);
nand U13154 (N_13154,N_9789,N_11214);
and U13155 (N_13155,N_9781,N_9273);
nand U13156 (N_13156,N_11054,N_9833);
and U13157 (N_13157,N_11321,N_11518);
nor U13158 (N_13158,N_11303,N_9490);
or U13159 (N_13159,N_11478,N_9644);
or U13160 (N_13160,N_10970,N_9865);
xnor U13161 (N_13161,N_11906,N_9884);
or U13162 (N_13162,N_9664,N_10157);
and U13163 (N_13163,N_11767,N_10716);
or U13164 (N_13164,N_10473,N_11025);
nor U13165 (N_13165,N_10938,N_11625);
nor U13166 (N_13166,N_11067,N_9323);
nor U13167 (N_13167,N_10339,N_10158);
or U13168 (N_13168,N_11714,N_10554);
or U13169 (N_13169,N_11871,N_11573);
nand U13170 (N_13170,N_9132,N_11512);
or U13171 (N_13171,N_11561,N_11899);
nand U13172 (N_13172,N_9391,N_10791);
nand U13173 (N_13173,N_11792,N_9727);
xnor U13174 (N_13174,N_10024,N_11992);
xor U13175 (N_13175,N_11898,N_10135);
or U13176 (N_13176,N_9270,N_10217);
and U13177 (N_13177,N_11683,N_9683);
and U13178 (N_13178,N_11514,N_9584);
nand U13179 (N_13179,N_9348,N_11043);
xor U13180 (N_13180,N_9435,N_9028);
or U13181 (N_13181,N_11904,N_10688);
and U13182 (N_13182,N_10111,N_9691);
and U13183 (N_13183,N_11971,N_9022);
and U13184 (N_13184,N_10622,N_10051);
nor U13185 (N_13185,N_9795,N_10008);
or U13186 (N_13186,N_11317,N_9670);
xnor U13187 (N_13187,N_11612,N_9468);
nor U13188 (N_13188,N_11631,N_9418);
and U13189 (N_13189,N_11680,N_9995);
nand U13190 (N_13190,N_11703,N_11022);
xnor U13191 (N_13191,N_10239,N_9610);
nand U13192 (N_13192,N_10700,N_9395);
or U13193 (N_13193,N_10372,N_9539);
nand U13194 (N_13194,N_9532,N_10846);
nand U13195 (N_13195,N_11202,N_9261);
or U13196 (N_13196,N_11589,N_9581);
nor U13197 (N_13197,N_9869,N_9080);
xnor U13198 (N_13198,N_10814,N_11516);
nor U13199 (N_13199,N_9775,N_9685);
and U13200 (N_13200,N_11245,N_10364);
xnor U13201 (N_13201,N_10800,N_10138);
and U13202 (N_13202,N_11981,N_10662);
nand U13203 (N_13203,N_10748,N_11241);
xnor U13204 (N_13204,N_10112,N_9399);
or U13205 (N_13205,N_10001,N_10276);
nor U13206 (N_13206,N_11646,N_10673);
nor U13207 (N_13207,N_11831,N_9061);
nand U13208 (N_13208,N_11200,N_10333);
nor U13209 (N_13209,N_10514,N_10921);
xnor U13210 (N_13210,N_11794,N_11758);
xor U13211 (N_13211,N_10308,N_11342);
and U13212 (N_13212,N_9499,N_9182);
and U13213 (N_13213,N_11240,N_10715);
nand U13214 (N_13214,N_10969,N_11037);
nor U13215 (N_13215,N_10282,N_10548);
and U13216 (N_13216,N_10618,N_11719);
and U13217 (N_13217,N_10540,N_9600);
nand U13218 (N_13218,N_10696,N_11035);
and U13219 (N_13219,N_9753,N_10904);
xor U13220 (N_13220,N_9654,N_10681);
and U13221 (N_13221,N_9452,N_9855);
xor U13222 (N_13222,N_10444,N_11803);
nand U13223 (N_13223,N_9304,N_9227);
nor U13224 (N_13224,N_11062,N_11882);
nor U13225 (N_13225,N_9459,N_9381);
xor U13226 (N_13226,N_9076,N_9745);
nand U13227 (N_13227,N_9514,N_9295);
xnor U13228 (N_13228,N_11781,N_10010);
nand U13229 (N_13229,N_9284,N_11046);
nand U13230 (N_13230,N_11967,N_11977);
nand U13231 (N_13231,N_9500,N_11401);
nor U13232 (N_13232,N_9959,N_11533);
xor U13233 (N_13233,N_9515,N_9937);
nand U13234 (N_13234,N_9973,N_10343);
or U13235 (N_13235,N_11376,N_11595);
xor U13236 (N_13236,N_10425,N_11619);
nand U13237 (N_13237,N_10136,N_10940);
nand U13238 (N_13238,N_10067,N_9620);
or U13239 (N_13239,N_9434,N_10857);
and U13240 (N_13240,N_10613,N_11658);
xor U13241 (N_13241,N_11039,N_9698);
or U13242 (N_13242,N_9303,N_10787);
or U13243 (N_13243,N_11582,N_10810);
nor U13244 (N_13244,N_11704,N_9492);
xnor U13245 (N_13245,N_10996,N_10439);
nand U13246 (N_13246,N_10852,N_10882);
xor U13247 (N_13247,N_9695,N_11183);
nand U13248 (N_13248,N_9156,N_9191);
nor U13249 (N_13249,N_9319,N_11371);
or U13250 (N_13250,N_10376,N_9042);
xnor U13251 (N_13251,N_10980,N_10371);
xnor U13252 (N_13252,N_11186,N_11474);
and U13253 (N_13253,N_9997,N_11215);
and U13254 (N_13254,N_10576,N_11667);
nand U13255 (N_13255,N_11178,N_9544);
nand U13256 (N_13256,N_9523,N_9297);
xnor U13257 (N_13257,N_9518,N_9007);
and U13258 (N_13258,N_9866,N_9917);
nand U13259 (N_13259,N_10871,N_9872);
and U13260 (N_13260,N_11159,N_10670);
nor U13261 (N_13261,N_10999,N_9471);
xnor U13262 (N_13262,N_9507,N_11969);
or U13263 (N_13263,N_11737,N_9788);
nor U13264 (N_13264,N_9681,N_11566);
nand U13265 (N_13265,N_10387,N_9030);
xnor U13266 (N_13266,N_10168,N_11963);
nor U13267 (N_13267,N_11265,N_11572);
and U13268 (N_13268,N_9569,N_10445);
nand U13269 (N_13269,N_10668,N_10269);
nor U13270 (N_13270,N_10617,N_10068);
nand U13271 (N_13271,N_11784,N_9099);
nor U13272 (N_13272,N_10248,N_10302);
xor U13273 (N_13273,N_9104,N_9638);
nand U13274 (N_13274,N_10960,N_9896);
nand U13275 (N_13275,N_9640,N_10265);
nor U13276 (N_13276,N_10987,N_10426);
xnor U13277 (N_13277,N_9936,N_11804);
and U13278 (N_13278,N_11162,N_11860);
and U13279 (N_13279,N_10442,N_10587);
xnor U13280 (N_13280,N_10936,N_10573);
or U13281 (N_13281,N_10082,N_10456);
nand U13282 (N_13282,N_9403,N_11965);
nand U13283 (N_13283,N_11862,N_11372);
and U13284 (N_13284,N_9345,N_11228);
and U13285 (N_13285,N_10515,N_9986);
and U13286 (N_13286,N_10062,N_10627);
or U13287 (N_13287,N_11013,N_10065);
or U13288 (N_13288,N_11717,N_9738);
nor U13289 (N_13289,N_10469,N_11143);
xor U13290 (N_13290,N_10398,N_10140);
nand U13291 (N_13291,N_9274,N_10544);
and U13292 (N_13292,N_10369,N_10336);
nor U13293 (N_13293,N_11500,N_9279);
nor U13294 (N_13294,N_10923,N_9926);
xor U13295 (N_13295,N_10028,N_10574);
or U13296 (N_13296,N_10698,N_9397);
or U13297 (N_13297,N_10049,N_9965);
nand U13298 (N_13298,N_10156,N_10676);
xnor U13299 (N_13299,N_9648,N_11288);
nand U13300 (N_13300,N_9379,N_10765);
xor U13301 (N_13301,N_9711,N_9301);
nand U13302 (N_13302,N_9387,N_10238);
nand U13303 (N_13303,N_10995,N_10139);
or U13304 (N_13304,N_11536,N_10298);
nor U13305 (N_13305,N_10020,N_9899);
xor U13306 (N_13306,N_10680,N_11727);
nand U13307 (N_13307,N_9946,N_11378);
nand U13308 (N_13308,N_9031,N_11699);
xor U13309 (N_13309,N_10694,N_11432);
and U13310 (N_13310,N_11297,N_9606);
or U13311 (N_13311,N_9631,N_11019);
and U13312 (N_13312,N_11277,N_10812);
xnor U13313 (N_13313,N_9063,N_11795);
nor U13314 (N_13314,N_11220,N_10767);
xor U13315 (N_13315,N_9118,N_10858);
nand U13316 (N_13316,N_9668,N_9630);
nand U13317 (N_13317,N_9419,N_11840);
xnor U13318 (N_13318,N_9818,N_11585);
or U13319 (N_13319,N_10169,N_9820);
and U13320 (N_13320,N_10697,N_11410);
nand U13321 (N_13321,N_9563,N_9734);
and U13322 (N_13322,N_11270,N_10869);
nor U13323 (N_13323,N_9909,N_10424);
nand U13324 (N_13324,N_11916,N_11353);
and U13325 (N_13325,N_11555,N_9955);
or U13326 (N_13326,N_10506,N_9441);
nand U13327 (N_13327,N_10368,N_10374);
nand U13328 (N_13328,N_10063,N_11905);
and U13329 (N_13329,N_11335,N_9130);
xnor U13330 (N_13330,N_11600,N_11309);
xor U13331 (N_13331,N_9969,N_9749);
nor U13332 (N_13332,N_10989,N_11356);
nor U13333 (N_13333,N_11844,N_11951);
nand U13334 (N_13334,N_10182,N_10312);
or U13335 (N_13335,N_11154,N_10589);
or U13336 (N_13336,N_10231,N_11995);
nor U13337 (N_13337,N_11362,N_11230);
and U13338 (N_13338,N_9062,N_9990);
nor U13339 (N_13339,N_9207,N_11608);
and U13340 (N_13340,N_9735,N_11021);
or U13341 (N_13341,N_10477,N_11073);
xnor U13342 (N_13342,N_9205,N_11493);
and U13343 (N_13343,N_11190,N_11644);
and U13344 (N_13344,N_9845,N_11196);
xor U13345 (N_13345,N_10380,N_10633);
or U13346 (N_13346,N_9230,N_11827);
or U13347 (N_13347,N_10635,N_9131);
nand U13348 (N_13348,N_9769,N_9433);
or U13349 (N_13349,N_10690,N_10804);
nand U13350 (N_13350,N_10516,N_10733);
nor U13351 (N_13351,N_11873,N_9082);
nand U13352 (N_13352,N_10579,N_10004);
nand U13353 (N_13353,N_10289,N_10902);
or U13354 (N_13354,N_11997,N_9421);
nand U13355 (N_13355,N_11593,N_11262);
xor U13356 (N_13356,N_11847,N_9091);
and U13357 (N_13357,N_10180,N_11629);
or U13358 (N_13358,N_11782,N_9961);
or U13359 (N_13359,N_10076,N_9339);
and U13360 (N_13360,N_9306,N_9474);
xor U13361 (N_13361,N_9798,N_11028);
nor U13362 (N_13362,N_11258,N_10064);
or U13363 (N_13363,N_9255,N_11527);
or U13364 (N_13364,N_9821,N_11843);
and U13365 (N_13365,N_11653,N_9810);
or U13366 (N_13366,N_10007,N_10581);
or U13367 (N_13367,N_11405,N_11902);
and U13368 (N_13368,N_9311,N_10592);
or U13369 (N_13369,N_10101,N_9247);
or U13370 (N_13370,N_9237,N_10133);
nand U13371 (N_13371,N_10737,N_11153);
and U13372 (N_13372,N_11851,N_9962);
and U13373 (N_13373,N_11458,N_10512);
nand U13374 (N_13374,N_10790,N_11144);
or U13375 (N_13375,N_10167,N_9386);
and U13376 (N_13376,N_11966,N_11756);
nor U13377 (N_13377,N_10321,N_9179);
or U13378 (N_13378,N_9473,N_9312);
or U13379 (N_13379,N_10195,N_9956);
and U13380 (N_13380,N_11813,N_10006);
or U13381 (N_13381,N_11318,N_9478);
or U13382 (N_13382,N_11471,N_9269);
and U13383 (N_13383,N_9267,N_11205);
or U13384 (N_13384,N_11730,N_9611);
and U13385 (N_13385,N_11748,N_11820);
or U13386 (N_13386,N_9583,N_10154);
nand U13387 (N_13387,N_9558,N_9596);
and U13388 (N_13388,N_9816,N_10390);
nor U13389 (N_13389,N_10489,N_9199);
and U13390 (N_13390,N_10734,N_10998);
nand U13391 (N_13391,N_9231,N_11686);
nor U13392 (N_13392,N_11538,N_10764);
nor U13393 (N_13393,N_9178,N_10395);
nand U13394 (N_13394,N_11052,N_11676);
and U13395 (N_13395,N_10009,N_10629);
nor U13396 (N_13396,N_10770,N_9756);
xnor U13397 (N_13397,N_10085,N_11874);
and U13398 (N_13398,N_10464,N_10120);
nand U13399 (N_13399,N_11528,N_10966);
xnor U13400 (N_13400,N_11298,N_11891);
xor U13401 (N_13401,N_10682,N_9768);
or U13402 (N_13402,N_10611,N_11711);
nand U13403 (N_13403,N_10731,N_9264);
xnor U13404 (N_13404,N_9054,N_10776);
nand U13405 (N_13405,N_9059,N_10610);
nor U13406 (N_13406,N_9032,N_9163);
and U13407 (N_13407,N_10531,N_11802);
nand U13408 (N_13408,N_11357,N_9679);
xor U13409 (N_13409,N_10796,N_10738);
or U13410 (N_13410,N_9850,N_10619);
xnor U13411 (N_13411,N_10580,N_11770);
or U13412 (N_13412,N_9501,N_10672);
and U13413 (N_13413,N_9902,N_11546);
nand U13414 (N_13414,N_10201,N_11210);
xnor U13415 (N_13415,N_10760,N_9882);
and U13416 (N_13416,N_9298,N_10799);
nand U13417 (N_13417,N_9017,N_11347);
and U13418 (N_13418,N_10381,N_10080);
xnor U13419 (N_13419,N_9197,N_10299);
xnor U13420 (N_13420,N_9757,N_11384);
or U13421 (N_13421,N_10771,N_11961);
nand U13422 (N_13422,N_10247,N_10652);
nor U13423 (N_13423,N_9084,N_10560);
and U13424 (N_13424,N_11763,N_10170);
or U13425 (N_13425,N_9752,N_11338);
nor U13426 (N_13426,N_9694,N_11893);
and U13427 (N_13427,N_10159,N_10891);
nand U13428 (N_13428,N_10632,N_11345);
and U13429 (N_13429,N_9504,N_11896);
or U13430 (N_13430,N_11878,N_11320);
nand U13431 (N_13431,N_11425,N_9102);
and U13432 (N_13432,N_10917,N_9024);
and U13433 (N_13433,N_9696,N_11989);
nand U13434 (N_13434,N_10614,N_10097);
or U13435 (N_13435,N_9879,N_9673);
xor U13436 (N_13436,N_10019,N_9204);
nand U13437 (N_13437,N_10689,N_10257);
xor U13438 (N_13438,N_11209,N_10539);
nor U13439 (N_13439,N_10656,N_9720);
xnor U13440 (N_13440,N_9782,N_10029);
or U13441 (N_13441,N_11604,N_10755);
or U13442 (N_13442,N_10947,N_10644);
nand U13443 (N_13443,N_9427,N_10849);
nand U13444 (N_13444,N_10189,N_10527);
nand U13445 (N_13445,N_11082,N_10990);
xor U13446 (N_13446,N_9643,N_11678);
and U13447 (N_13447,N_10979,N_10178);
nor U13448 (N_13448,N_10772,N_9385);
and U13449 (N_13449,N_9073,N_11063);
xor U13450 (N_13450,N_9114,N_9495);
xnor U13451 (N_13451,N_10482,N_11605);
or U13452 (N_13452,N_11675,N_10119);
nor U13453 (N_13453,N_11914,N_10300);
nand U13454 (N_13454,N_11072,N_11935);
nand U13455 (N_13455,N_11836,N_11883);
nand U13456 (N_13456,N_10674,N_10856);
and U13457 (N_13457,N_11381,N_11423);
nor U13458 (N_13458,N_9580,N_11001);
nand U13459 (N_13459,N_10918,N_11267);
nand U13460 (N_13460,N_11952,N_9847);
nor U13461 (N_13461,N_9574,N_11998);
nand U13462 (N_13462,N_9542,N_9139);
nand U13463 (N_13463,N_10094,N_10002);
and U13464 (N_13464,N_11901,N_9744);
nor U13465 (N_13465,N_10559,N_11045);
and U13466 (N_13466,N_11869,N_10968);
or U13467 (N_13467,N_9089,N_11443);
xnor U13468 (N_13468,N_11225,N_11567);
nand U13469 (N_13469,N_9854,N_11191);
nand U13470 (N_13470,N_11652,N_9849);
nand U13471 (N_13471,N_9208,N_9661);
or U13472 (N_13472,N_11207,N_10749);
and U13473 (N_13473,N_9857,N_9289);
or U13474 (N_13474,N_10896,N_11819);
xnor U13475 (N_13475,N_10012,N_10033);
nor U13476 (N_13476,N_11248,N_9579);
xnor U13477 (N_13477,N_10022,N_11876);
or U13478 (N_13478,N_11810,N_9008);
and U13479 (N_13479,N_11015,N_11823);
and U13480 (N_13480,N_9677,N_11828);
nand U13481 (N_13481,N_9340,N_11290);
nor U13482 (N_13482,N_11832,N_11505);
xor U13483 (N_13483,N_9287,N_11665);
and U13484 (N_13484,N_11835,N_11198);
and U13485 (N_13485,N_11096,N_11636);
nand U13486 (N_13486,N_9236,N_11506);
and U13487 (N_13487,N_11919,N_11227);
nand U13488 (N_13488,N_9203,N_10218);
nor U13489 (N_13489,N_11463,N_11349);
or U13490 (N_13490,N_11140,N_9027);
nor U13491 (N_13491,N_9750,N_11682);
nand U13492 (N_13492,N_11004,N_11864);
xor U13493 (N_13493,N_9906,N_11581);
and U13494 (N_13494,N_11944,N_11517);
nor U13495 (N_13495,N_10965,N_10487);
nor U13496 (N_13496,N_10235,N_9169);
or U13497 (N_13497,N_9546,N_9183);
or U13498 (N_13498,N_11731,N_11545);
xor U13499 (N_13499,N_9079,N_9305);
nor U13500 (N_13500,N_10569,N_9086);
or U13501 (N_13501,N_9937,N_10226);
nand U13502 (N_13502,N_11066,N_9470);
nor U13503 (N_13503,N_10098,N_11832);
or U13504 (N_13504,N_11810,N_10110);
xnor U13505 (N_13505,N_10190,N_9304);
xor U13506 (N_13506,N_11733,N_9496);
and U13507 (N_13507,N_11037,N_11176);
nand U13508 (N_13508,N_11731,N_9799);
or U13509 (N_13509,N_10663,N_9069);
nor U13510 (N_13510,N_11818,N_11674);
nor U13511 (N_13511,N_11630,N_11754);
and U13512 (N_13512,N_10126,N_11935);
nor U13513 (N_13513,N_10164,N_11232);
xor U13514 (N_13514,N_10397,N_10950);
xor U13515 (N_13515,N_9617,N_11309);
nand U13516 (N_13516,N_9979,N_9349);
and U13517 (N_13517,N_9852,N_9869);
nor U13518 (N_13518,N_9998,N_10024);
nand U13519 (N_13519,N_10797,N_10390);
xnor U13520 (N_13520,N_11810,N_10210);
nor U13521 (N_13521,N_9088,N_11766);
or U13522 (N_13522,N_9290,N_9503);
xnor U13523 (N_13523,N_11540,N_10081);
and U13524 (N_13524,N_10392,N_9442);
nor U13525 (N_13525,N_10176,N_9400);
xnor U13526 (N_13526,N_9574,N_10908);
nand U13527 (N_13527,N_11363,N_11276);
and U13528 (N_13528,N_9064,N_10765);
and U13529 (N_13529,N_11185,N_11145);
or U13530 (N_13530,N_11952,N_11458);
nand U13531 (N_13531,N_9145,N_11017);
and U13532 (N_13532,N_9048,N_9968);
and U13533 (N_13533,N_11469,N_10415);
and U13534 (N_13534,N_10596,N_11865);
or U13535 (N_13535,N_9451,N_11523);
xnor U13536 (N_13536,N_11143,N_10491);
nand U13537 (N_13537,N_10494,N_9725);
and U13538 (N_13538,N_10973,N_9756);
and U13539 (N_13539,N_10963,N_10919);
nand U13540 (N_13540,N_10763,N_10167);
nor U13541 (N_13541,N_9713,N_9978);
nor U13542 (N_13542,N_9791,N_10009);
nor U13543 (N_13543,N_11618,N_9204);
nand U13544 (N_13544,N_10955,N_9178);
xnor U13545 (N_13545,N_10009,N_9858);
and U13546 (N_13546,N_11388,N_11339);
and U13547 (N_13547,N_9124,N_9544);
nand U13548 (N_13548,N_10554,N_11745);
nand U13549 (N_13549,N_9932,N_9561);
nor U13550 (N_13550,N_10982,N_10244);
and U13551 (N_13551,N_9115,N_10372);
nand U13552 (N_13552,N_9609,N_9613);
nor U13553 (N_13553,N_11221,N_9281);
nand U13554 (N_13554,N_9258,N_11053);
xor U13555 (N_13555,N_10243,N_11412);
xor U13556 (N_13556,N_10149,N_10641);
nand U13557 (N_13557,N_10918,N_11256);
nand U13558 (N_13558,N_11908,N_10766);
or U13559 (N_13559,N_10778,N_9409);
xor U13560 (N_13560,N_10848,N_11921);
nand U13561 (N_13561,N_10631,N_9716);
xnor U13562 (N_13562,N_9336,N_11268);
nand U13563 (N_13563,N_10756,N_9274);
nand U13564 (N_13564,N_9496,N_9322);
nor U13565 (N_13565,N_9057,N_10701);
and U13566 (N_13566,N_11884,N_11604);
or U13567 (N_13567,N_11200,N_10130);
nor U13568 (N_13568,N_10694,N_11219);
and U13569 (N_13569,N_10769,N_11372);
nor U13570 (N_13570,N_10540,N_10175);
or U13571 (N_13571,N_11247,N_11151);
nand U13572 (N_13572,N_9325,N_9632);
nor U13573 (N_13573,N_10178,N_11056);
nor U13574 (N_13574,N_10548,N_9196);
and U13575 (N_13575,N_9719,N_10889);
or U13576 (N_13576,N_11303,N_9742);
and U13577 (N_13577,N_10541,N_10860);
or U13578 (N_13578,N_10689,N_10832);
nand U13579 (N_13579,N_9461,N_11013);
or U13580 (N_13580,N_11591,N_9413);
xnor U13581 (N_13581,N_10140,N_11346);
xnor U13582 (N_13582,N_10917,N_10156);
xor U13583 (N_13583,N_10300,N_10160);
and U13584 (N_13584,N_11477,N_9820);
xnor U13585 (N_13585,N_10501,N_9832);
xnor U13586 (N_13586,N_11317,N_9917);
and U13587 (N_13587,N_10749,N_10403);
xnor U13588 (N_13588,N_9004,N_9391);
or U13589 (N_13589,N_11147,N_10772);
xor U13590 (N_13590,N_10999,N_10987);
xnor U13591 (N_13591,N_9154,N_11455);
and U13592 (N_13592,N_11574,N_11470);
or U13593 (N_13593,N_9645,N_10981);
nor U13594 (N_13594,N_10147,N_9604);
xor U13595 (N_13595,N_9652,N_9459);
and U13596 (N_13596,N_11492,N_10711);
nand U13597 (N_13597,N_10306,N_9829);
or U13598 (N_13598,N_9584,N_9570);
nor U13599 (N_13599,N_10623,N_10708);
or U13600 (N_13600,N_9537,N_11938);
and U13601 (N_13601,N_11683,N_11146);
and U13602 (N_13602,N_10509,N_11499);
xnor U13603 (N_13603,N_9301,N_10379);
nor U13604 (N_13604,N_10456,N_10199);
nand U13605 (N_13605,N_9917,N_10599);
xor U13606 (N_13606,N_10073,N_11392);
or U13607 (N_13607,N_11169,N_9328);
xor U13608 (N_13608,N_9375,N_9390);
xnor U13609 (N_13609,N_9447,N_10574);
or U13610 (N_13610,N_9391,N_9010);
or U13611 (N_13611,N_11040,N_10621);
xnor U13612 (N_13612,N_10590,N_10431);
and U13613 (N_13613,N_11721,N_10974);
and U13614 (N_13614,N_9249,N_10426);
nand U13615 (N_13615,N_11916,N_10664);
or U13616 (N_13616,N_11569,N_10531);
or U13617 (N_13617,N_10331,N_10959);
xnor U13618 (N_13618,N_10395,N_10446);
or U13619 (N_13619,N_10126,N_9748);
or U13620 (N_13620,N_11594,N_9151);
nand U13621 (N_13621,N_11939,N_10460);
xor U13622 (N_13622,N_11597,N_9845);
nor U13623 (N_13623,N_10768,N_10825);
and U13624 (N_13624,N_10747,N_10282);
or U13625 (N_13625,N_11211,N_9938);
and U13626 (N_13626,N_9102,N_11223);
or U13627 (N_13627,N_11234,N_10867);
nor U13628 (N_13628,N_9604,N_9876);
nor U13629 (N_13629,N_9478,N_9809);
or U13630 (N_13630,N_11595,N_10870);
xnor U13631 (N_13631,N_10074,N_11746);
and U13632 (N_13632,N_11045,N_11373);
xnor U13633 (N_13633,N_10412,N_10602);
nor U13634 (N_13634,N_11404,N_9711);
and U13635 (N_13635,N_10367,N_10930);
xor U13636 (N_13636,N_9061,N_9481);
and U13637 (N_13637,N_9063,N_9017);
xor U13638 (N_13638,N_10312,N_11843);
nor U13639 (N_13639,N_10890,N_9387);
nor U13640 (N_13640,N_10600,N_9967);
nand U13641 (N_13641,N_11390,N_11881);
nand U13642 (N_13642,N_11859,N_11654);
xnor U13643 (N_13643,N_9483,N_10100);
nand U13644 (N_13644,N_10498,N_10627);
xnor U13645 (N_13645,N_10682,N_11657);
or U13646 (N_13646,N_11093,N_11371);
nand U13647 (N_13647,N_10508,N_9778);
and U13648 (N_13648,N_9334,N_10431);
nand U13649 (N_13649,N_9897,N_9213);
nor U13650 (N_13650,N_9494,N_9004);
or U13651 (N_13651,N_9715,N_10434);
and U13652 (N_13652,N_11948,N_10124);
and U13653 (N_13653,N_11219,N_11118);
nor U13654 (N_13654,N_10410,N_9650);
nor U13655 (N_13655,N_11260,N_11602);
nor U13656 (N_13656,N_9517,N_9185);
nand U13657 (N_13657,N_9119,N_10875);
and U13658 (N_13658,N_9248,N_9463);
xnor U13659 (N_13659,N_10126,N_9167);
or U13660 (N_13660,N_10830,N_11004);
and U13661 (N_13661,N_9984,N_10886);
and U13662 (N_13662,N_10062,N_11591);
and U13663 (N_13663,N_10597,N_11196);
xor U13664 (N_13664,N_11469,N_10766);
and U13665 (N_13665,N_10633,N_9402);
xnor U13666 (N_13666,N_10893,N_11900);
and U13667 (N_13667,N_10631,N_11687);
nand U13668 (N_13668,N_11680,N_10180);
or U13669 (N_13669,N_10887,N_9985);
xnor U13670 (N_13670,N_9435,N_9764);
or U13671 (N_13671,N_11585,N_10664);
xor U13672 (N_13672,N_11850,N_10825);
or U13673 (N_13673,N_9184,N_10595);
or U13674 (N_13674,N_9282,N_9567);
nand U13675 (N_13675,N_9622,N_9193);
xor U13676 (N_13676,N_11000,N_11115);
nand U13677 (N_13677,N_10049,N_9679);
xnor U13678 (N_13678,N_10173,N_9598);
and U13679 (N_13679,N_11971,N_10428);
and U13680 (N_13680,N_9729,N_9534);
nor U13681 (N_13681,N_10707,N_10236);
nor U13682 (N_13682,N_11733,N_11631);
or U13683 (N_13683,N_9986,N_10882);
or U13684 (N_13684,N_9119,N_10685);
nand U13685 (N_13685,N_10331,N_9750);
nor U13686 (N_13686,N_10420,N_10847);
or U13687 (N_13687,N_11521,N_9714);
nand U13688 (N_13688,N_11942,N_9664);
xor U13689 (N_13689,N_10940,N_9226);
xnor U13690 (N_13690,N_9303,N_9951);
xor U13691 (N_13691,N_10012,N_10044);
and U13692 (N_13692,N_10968,N_9422);
or U13693 (N_13693,N_10549,N_10022);
or U13694 (N_13694,N_11996,N_9942);
and U13695 (N_13695,N_10864,N_10557);
and U13696 (N_13696,N_10471,N_11016);
and U13697 (N_13697,N_11518,N_9299);
nor U13698 (N_13698,N_9977,N_9335);
nand U13699 (N_13699,N_10775,N_10900);
xor U13700 (N_13700,N_10382,N_9843);
and U13701 (N_13701,N_9920,N_10763);
and U13702 (N_13702,N_11025,N_11010);
nor U13703 (N_13703,N_9052,N_11705);
nand U13704 (N_13704,N_10502,N_11586);
nor U13705 (N_13705,N_9176,N_9287);
or U13706 (N_13706,N_11812,N_9878);
xnor U13707 (N_13707,N_9902,N_9635);
or U13708 (N_13708,N_11011,N_11543);
or U13709 (N_13709,N_11158,N_9425);
xnor U13710 (N_13710,N_9746,N_11294);
and U13711 (N_13711,N_11196,N_9188);
nor U13712 (N_13712,N_11291,N_11808);
nor U13713 (N_13713,N_11030,N_9894);
and U13714 (N_13714,N_9500,N_9841);
nand U13715 (N_13715,N_11214,N_10056);
nor U13716 (N_13716,N_10194,N_9191);
nor U13717 (N_13717,N_9520,N_11792);
or U13718 (N_13718,N_10948,N_9976);
nor U13719 (N_13719,N_10504,N_11354);
xor U13720 (N_13720,N_9030,N_10736);
nand U13721 (N_13721,N_10723,N_11400);
nor U13722 (N_13722,N_11077,N_10920);
and U13723 (N_13723,N_10917,N_11169);
nor U13724 (N_13724,N_9946,N_10886);
nor U13725 (N_13725,N_10560,N_11750);
and U13726 (N_13726,N_11605,N_10852);
nor U13727 (N_13727,N_11696,N_11719);
or U13728 (N_13728,N_11614,N_10994);
or U13729 (N_13729,N_11686,N_11229);
nand U13730 (N_13730,N_9300,N_9741);
xor U13731 (N_13731,N_10489,N_9604);
nor U13732 (N_13732,N_9043,N_9271);
nor U13733 (N_13733,N_10825,N_11482);
and U13734 (N_13734,N_9587,N_10641);
or U13735 (N_13735,N_9143,N_10960);
nand U13736 (N_13736,N_10889,N_10549);
xnor U13737 (N_13737,N_11379,N_10526);
xor U13738 (N_13738,N_11772,N_10502);
and U13739 (N_13739,N_10760,N_11319);
xor U13740 (N_13740,N_11809,N_11895);
or U13741 (N_13741,N_10068,N_10513);
xor U13742 (N_13742,N_11950,N_11525);
and U13743 (N_13743,N_9400,N_9443);
nand U13744 (N_13744,N_10252,N_11794);
nor U13745 (N_13745,N_9988,N_10063);
nand U13746 (N_13746,N_10169,N_9032);
nor U13747 (N_13747,N_9520,N_10573);
xor U13748 (N_13748,N_10366,N_10745);
nand U13749 (N_13749,N_9759,N_11525);
nor U13750 (N_13750,N_9670,N_9070);
nand U13751 (N_13751,N_9695,N_11896);
or U13752 (N_13752,N_11895,N_10362);
nand U13753 (N_13753,N_11695,N_11643);
and U13754 (N_13754,N_10511,N_10738);
or U13755 (N_13755,N_9368,N_10998);
nor U13756 (N_13756,N_10575,N_9739);
nor U13757 (N_13757,N_10229,N_9989);
and U13758 (N_13758,N_11454,N_10853);
nand U13759 (N_13759,N_10944,N_11131);
nor U13760 (N_13760,N_9189,N_10870);
xor U13761 (N_13761,N_9189,N_9370);
and U13762 (N_13762,N_10044,N_10589);
nor U13763 (N_13763,N_9609,N_10602);
nor U13764 (N_13764,N_11991,N_11324);
nor U13765 (N_13765,N_11789,N_11290);
nor U13766 (N_13766,N_11551,N_11930);
and U13767 (N_13767,N_10528,N_10722);
nor U13768 (N_13768,N_9545,N_10783);
nand U13769 (N_13769,N_11849,N_10094);
and U13770 (N_13770,N_10379,N_11897);
nand U13771 (N_13771,N_10598,N_11632);
nor U13772 (N_13772,N_11536,N_9014);
nand U13773 (N_13773,N_11556,N_11331);
xor U13774 (N_13774,N_10591,N_11779);
nor U13775 (N_13775,N_11176,N_10300);
xnor U13776 (N_13776,N_11897,N_9161);
and U13777 (N_13777,N_9061,N_10652);
xnor U13778 (N_13778,N_11549,N_9732);
or U13779 (N_13779,N_10829,N_10687);
nand U13780 (N_13780,N_11377,N_9437);
nor U13781 (N_13781,N_9899,N_9588);
or U13782 (N_13782,N_9949,N_9922);
or U13783 (N_13783,N_9856,N_10803);
nand U13784 (N_13784,N_11329,N_11754);
xor U13785 (N_13785,N_10569,N_11949);
and U13786 (N_13786,N_11922,N_9541);
nor U13787 (N_13787,N_10489,N_11827);
or U13788 (N_13788,N_11698,N_10035);
or U13789 (N_13789,N_9755,N_9656);
xor U13790 (N_13790,N_11347,N_11586);
nor U13791 (N_13791,N_11451,N_11197);
nor U13792 (N_13792,N_10630,N_9522);
nand U13793 (N_13793,N_10227,N_9102);
xnor U13794 (N_13794,N_11685,N_11872);
and U13795 (N_13795,N_9865,N_10788);
and U13796 (N_13796,N_10504,N_10689);
xnor U13797 (N_13797,N_9587,N_9469);
xor U13798 (N_13798,N_10864,N_11931);
xnor U13799 (N_13799,N_9911,N_9378);
or U13800 (N_13800,N_10482,N_10677);
xnor U13801 (N_13801,N_10681,N_11680);
nand U13802 (N_13802,N_11950,N_11447);
or U13803 (N_13803,N_10656,N_10225);
and U13804 (N_13804,N_10673,N_9915);
and U13805 (N_13805,N_10517,N_9708);
nand U13806 (N_13806,N_10144,N_10322);
nand U13807 (N_13807,N_9914,N_11124);
xnor U13808 (N_13808,N_9378,N_9309);
nand U13809 (N_13809,N_10909,N_10192);
nor U13810 (N_13810,N_11406,N_10108);
or U13811 (N_13811,N_9765,N_9192);
and U13812 (N_13812,N_10994,N_10821);
or U13813 (N_13813,N_10455,N_11332);
xor U13814 (N_13814,N_10608,N_11870);
xnor U13815 (N_13815,N_10113,N_11038);
or U13816 (N_13816,N_11034,N_9819);
or U13817 (N_13817,N_9912,N_10892);
xor U13818 (N_13818,N_9466,N_9861);
and U13819 (N_13819,N_10195,N_11251);
and U13820 (N_13820,N_9808,N_9341);
nand U13821 (N_13821,N_11637,N_10518);
nor U13822 (N_13822,N_11964,N_11238);
nor U13823 (N_13823,N_10664,N_9240);
nand U13824 (N_13824,N_10233,N_11998);
nand U13825 (N_13825,N_9681,N_10990);
or U13826 (N_13826,N_11280,N_10057);
and U13827 (N_13827,N_11887,N_10768);
nand U13828 (N_13828,N_10376,N_9230);
nor U13829 (N_13829,N_9599,N_9713);
xnor U13830 (N_13830,N_11809,N_9711);
nand U13831 (N_13831,N_11597,N_9716);
xor U13832 (N_13832,N_10477,N_10457);
or U13833 (N_13833,N_10178,N_10460);
nand U13834 (N_13834,N_9759,N_11880);
and U13835 (N_13835,N_9030,N_9543);
xnor U13836 (N_13836,N_9306,N_11734);
nor U13837 (N_13837,N_10251,N_11082);
or U13838 (N_13838,N_9668,N_10144);
and U13839 (N_13839,N_10490,N_10219);
nor U13840 (N_13840,N_10784,N_11337);
or U13841 (N_13841,N_10312,N_10339);
or U13842 (N_13842,N_9531,N_9355);
nand U13843 (N_13843,N_10194,N_10154);
nand U13844 (N_13844,N_10943,N_9879);
nand U13845 (N_13845,N_9049,N_10084);
nand U13846 (N_13846,N_10614,N_9367);
nand U13847 (N_13847,N_9409,N_10783);
and U13848 (N_13848,N_10406,N_11074);
nand U13849 (N_13849,N_9899,N_11890);
and U13850 (N_13850,N_9064,N_9285);
or U13851 (N_13851,N_10496,N_10341);
xnor U13852 (N_13852,N_9375,N_10447);
nand U13853 (N_13853,N_10403,N_10663);
xnor U13854 (N_13854,N_10343,N_10539);
or U13855 (N_13855,N_10326,N_11789);
nand U13856 (N_13856,N_9274,N_9962);
and U13857 (N_13857,N_11225,N_9268);
nand U13858 (N_13858,N_11959,N_9266);
or U13859 (N_13859,N_10083,N_9182);
and U13860 (N_13860,N_11551,N_11920);
or U13861 (N_13861,N_9487,N_9356);
xnor U13862 (N_13862,N_10706,N_11619);
nor U13863 (N_13863,N_11652,N_9410);
xnor U13864 (N_13864,N_10763,N_9106);
xor U13865 (N_13865,N_10105,N_9192);
nor U13866 (N_13866,N_11403,N_10835);
xnor U13867 (N_13867,N_11620,N_9895);
nor U13868 (N_13868,N_9995,N_10807);
or U13869 (N_13869,N_9501,N_9259);
nor U13870 (N_13870,N_9546,N_10847);
nand U13871 (N_13871,N_9072,N_9836);
nand U13872 (N_13872,N_10128,N_11243);
xor U13873 (N_13873,N_9810,N_11630);
and U13874 (N_13874,N_11278,N_10183);
nand U13875 (N_13875,N_9602,N_11524);
and U13876 (N_13876,N_11398,N_9608);
nor U13877 (N_13877,N_11698,N_10784);
nor U13878 (N_13878,N_9624,N_10505);
xnor U13879 (N_13879,N_11387,N_9243);
nor U13880 (N_13880,N_10396,N_11922);
nor U13881 (N_13881,N_11345,N_9775);
or U13882 (N_13882,N_9940,N_11982);
and U13883 (N_13883,N_10359,N_10922);
or U13884 (N_13884,N_9925,N_11997);
and U13885 (N_13885,N_10038,N_9519);
nand U13886 (N_13886,N_11136,N_10927);
nor U13887 (N_13887,N_9800,N_11645);
nor U13888 (N_13888,N_11160,N_11962);
and U13889 (N_13889,N_11487,N_9056);
nand U13890 (N_13890,N_9918,N_9868);
or U13891 (N_13891,N_11308,N_11990);
and U13892 (N_13892,N_9368,N_9741);
and U13893 (N_13893,N_11293,N_11488);
xnor U13894 (N_13894,N_9343,N_9561);
nand U13895 (N_13895,N_10160,N_11465);
nand U13896 (N_13896,N_9956,N_10693);
and U13897 (N_13897,N_9097,N_11460);
nand U13898 (N_13898,N_11407,N_9449);
nand U13899 (N_13899,N_10616,N_10720);
nor U13900 (N_13900,N_10618,N_10283);
nand U13901 (N_13901,N_11078,N_9657);
nor U13902 (N_13902,N_10746,N_9483);
xor U13903 (N_13903,N_9767,N_9510);
xor U13904 (N_13904,N_11303,N_10658);
nor U13905 (N_13905,N_9140,N_11520);
nand U13906 (N_13906,N_10230,N_11121);
nor U13907 (N_13907,N_11550,N_9428);
nand U13908 (N_13908,N_11362,N_10704);
and U13909 (N_13909,N_9146,N_11336);
nor U13910 (N_13910,N_10704,N_9717);
nor U13911 (N_13911,N_10737,N_10532);
nand U13912 (N_13912,N_9226,N_10720);
nand U13913 (N_13913,N_9034,N_11163);
nand U13914 (N_13914,N_11493,N_11025);
nand U13915 (N_13915,N_10866,N_9904);
nand U13916 (N_13916,N_9644,N_9168);
or U13917 (N_13917,N_11297,N_9964);
nor U13918 (N_13918,N_11665,N_11028);
or U13919 (N_13919,N_11196,N_11302);
xnor U13920 (N_13920,N_10815,N_10621);
nand U13921 (N_13921,N_11619,N_9561);
and U13922 (N_13922,N_10498,N_10976);
or U13923 (N_13923,N_10184,N_11123);
or U13924 (N_13924,N_10568,N_10062);
nor U13925 (N_13925,N_9994,N_9263);
nand U13926 (N_13926,N_11804,N_10891);
and U13927 (N_13927,N_11388,N_11390);
or U13928 (N_13928,N_11833,N_9048);
or U13929 (N_13929,N_10431,N_11004);
or U13930 (N_13930,N_10150,N_9443);
xor U13931 (N_13931,N_9578,N_10292);
xnor U13932 (N_13932,N_11883,N_10947);
nor U13933 (N_13933,N_10531,N_10012);
nand U13934 (N_13934,N_11297,N_11900);
nand U13935 (N_13935,N_10073,N_10367);
or U13936 (N_13936,N_9147,N_11768);
and U13937 (N_13937,N_11372,N_11751);
xor U13938 (N_13938,N_9442,N_10524);
nor U13939 (N_13939,N_10448,N_10554);
nand U13940 (N_13940,N_9936,N_10154);
nor U13941 (N_13941,N_9338,N_9083);
nand U13942 (N_13942,N_10249,N_11366);
xor U13943 (N_13943,N_9452,N_11925);
nor U13944 (N_13944,N_9505,N_11312);
and U13945 (N_13945,N_10978,N_9642);
xor U13946 (N_13946,N_10141,N_11189);
or U13947 (N_13947,N_9556,N_10582);
nand U13948 (N_13948,N_11130,N_11345);
xnor U13949 (N_13949,N_10163,N_10315);
nand U13950 (N_13950,N_10270,N_11488);
xor U13951 (N_13951,N_11051,N_10993);
xor U13952 (N_13952,N_11553,N_10359);
nor U13953 (N_13953,N_11718,N_9290);
nand U13954 (N_13954,N_10679,N_11472);
and U13955 (N_13955,N_11093,N_10843);
nand U13956 (N_13956,N_10961,N_11291);
nor U13957 (N_13957,N_9420,N_9907);
and U13958 (N_13958,N_9484,N_11226);
and U13959 (N_13959,N_10025,N_9153);
and U13960 (N_13960,N_9876,N_10000);
and U13961 (N_13961,N_11111,N_10482);
nand U13962 (N_13962,N_9615,N_10781);
nor U13963 (N_13963,N_11712,N_9843);
or U13964 (N_13964,N_11420,N_9381);
xnor U13965 (N_13965,N_9991,N_11809);
nand U13966 (N_13966,N_10072,N_11942);
or U13967 (N_13967,N_11681,N_11252);
nor U13968 (N_13968,N_10733,N_10699);
or U13969 (N_13969,N_10808,N_11506);
nor U13970 (N_13970,N_11663,N_11368);
xnor U13971 (N_13971,N_11939,N_9437);
and U13972 (N_13972,N_9378,N_11037);
or U13973 (N_13973,N_9677,N_9053);
nand U13974 (N_13974,N_10026,N_10913);
and U13975 (N_13975,N_9791,N_10989);
nand U13976 (N_13976,N_9385,N_9088);
nand U13977 (N_13977,N_9180,N_9315);
nand U13978 (N_13978,N_10437,N_9585);
and U13979 (N_13979,N_11234,N_10482);
nand U13980 (N_13980,N_9905,N_11707);
and U13981 (N_13981,N_10920,N_11431);
xnor U13982 (N_13982,N_10621,N_9177);
xor U13983 (N_13983,N_9448,N_11223);
nand U13984 (N_13984,N_9763,N_11211);
or U13985 (N_13985,N_11379,N_10895);
nand U13986 (N_13986,N_9022,N_10894);
nor U13987 (N_13987,N_10392,N_10012);
or U13988 (N_13988,N_9673,N_11278);
xor U13989 (N_13989,N_11966,N_11858);
or U13990 (N_13990,N_9809,N_9894);
and U13991 (N_13991,N_10118,N_10404);
nand U13992 (N_13992,N_10860,N_10435);
nand U13993 (N_13993,N_9915,N_10263);
or U13994 (N_13994,N_10295,N_11322);
nor U13995 (N_13995,N_9475,N_10678);
nor U13996 (N_13996,N_10035,N_9596);
or U13997 (N_13997,N_11755,N_11420);
nand U13998 (N_13998,N_11607,N_11513);
and U13999 (N_13999,N_11091,N_11535);
xnor U14000 (N_14000,N_9627,N_9765);
nand U14001 (N_14001,N_10129,N_11368);
nand U14002 (N_14002,N_11010,N_10575);
xnor U14003 (N_14003,N_9238,N_11225);
nand U14004 (N_14004,N_9310,N_11006);
xor U14005 (N_14005,N_11450,N_11542);
and U14006 (N_14006,N_10026,N_10984);
nand U14007 (N_14007,N_10531,N_10151);
nand U14008 (N_14008,N_9919,N_11134);
or U14009 (N_14009,N_9367,N_10506);
or U14010 (N_14010,N_9927,N_9858);
nand U14011 (N_14011,N_10658,N_9377);
and U14012 (N_14012,N_11071,N_10321);
nor U14013 (N_14013,N_9757,N_11045);
nand U14014 (N_14014,N_10262,N_11830);
or U14015 (N_14015,N_10459,N_9880);
or U14016 (N_14016,N_11445,N_9518);
and U14017 (N_14017,N_9138,N_10212);
xnor U14018 (N_14018,N_10367,N_11801);
xor U14019 (N_14019,N_11346,N_9367);
nor U14020 (N_14020,N_10167,N_11907);
xnor U14021 (N_14021,N_9941,N_10388);
nand U14022 (N_14022,N_11165,N_11199);
or U14023 (N_14023,N_10995,N_9730);
nor U14024 (N_14024,N_10698,N_9688);
xnor U14025 (N_14025,N_9836,N_11523);
nor U14026 (N_14026,N_10559,N_9823);
and U14027 (N_14027,N_11284,N_11081);
nand U14028 (N_14028,N_11767,N_10313);
nor U14029 (N_14029,N_11139,N_9356);
or U14030 (N_14030,N_11398,N_10973);
nor U14031 (N_14031,N_11344,N_10144);
or U14032 (N_14032,N_10555,N_10562);
nor U14033 (N_14033,N_9851,N_9270);
nand U14034 (N_14034,N_11369,N_11532);
or U14035 (N_14035,N_9474,N_10180);
nor U14036 (N_14036,N_9135,N_11595);
nand U14037 (N_14037,N_11520,N_9439);
nand U14038 (N_14038,N_11769,N_10554);
nor U14039 (N_14039,N_10409,N_11439);
xor U14040 (N_14040,N_10268,N_10174);
xnor U14041 (N_14041,N_9881,N_10622);
xnor U14042 (N_14042,N_11123,N_9083);
xnor U14043 (N_14043,N_9739,N_10879);
or U14044 (N_14044,N_11497,N_11158);
or U14045 (N_14045,N_9719,N_9721);
and U14046 (N_14046,N_10644,N_10416);
or U14047 (N_14047,N_9621,N_11511);
xor U14048 (N_14048,N_10244,N_9975);
nor U14049 (N_14049,N_11557,N_10753);
nand U14050 (N_14050,N_10276,N_11771);
and U14051 (N_14051,N_10898,N_11760);
nor U14052 (N_14052,N_9096,N_9194);
nand U14053 (N_14053,N_10313,N_10626);
nand U14054 (N_14054,N_10483,N_9883);
and U14055 (N_14055,N_11028,N_10214);
or U14056 (N_14056,N_10553,N_10010);
nor U14057 (N_14057,N_10621,N_9868);
nand U14058 (N_14058,N_11770,N_10597);
nand U14059 (N_14059,N_9619,N_11877);
nor U14060 (N_14060,N_10381,N_11317);
or U14061 (N_14061,N_11713,N_10435);
or U14062 (N_14062,N_11367,N_9515);
xnor U14063 (N_14063,N_9449,N_10221);
or U14064 (N_14064,N_11863,N_10491);
nand U14065 (N_14065,N_9318,N_10800);
and U14066 (N_14066,N_9120,N_11493);
and U14067 (N_14067,N_10202,N_9203);
nor U14068 (N_14068,N_10073,N_10340);
or U14069 (N_14069,N_10507,N_9329);
or U14070 (N_14070,N_11690,N_10694);
or U14071 (N_14071,N_11798,N_9973);
xnor U14072 (N_14072,N_9593,N_9582);
or U14073 (N_14073,N_10119,N_9551);
and U14074 (N_14074,N_11626,N_10302);
and U14075 (N_14075,N_10479,N_9332);
nand U14076 (N_14076,N_10579,N_11998);
xor U14077 (N_14077,N_10971,N_9005);
nor U14078 (N_14078,N_9763,N_9409);
xor U14079 (N_14079,N_10114,N_9946);
and U14080 (N_14080,N_11782,N_9627);
xor U14081 (N_14081,N_11927,N_10668);
and U14082 (N_14082,N_11500,N_9568);
nand U14083 (N_14083,N_9976,N_10339);
nand U14084 (N_14084,N_11802,N_10544);
and U14085 (N_14085,N_11608,N_10120);
and U14086 (N_14086,N_11561,N_10713);
nand U14087 (N_14087,N_10005,N_9954);
xnor U14088 (N_14088,N_10452,N_10125);
xor U14089 (N_14089,N_9038,N_11250);
nor U14090 (N_14090,N_10973,N_11445);
nand U14091 (N_14091,N_10626,N_11355);
xnor U14092 (N_14092,N_10880,N_9152);
nor U14093 (N_14093,N_11109,N_10839);
nor U14094 (N_14094,N_9620,N_9357);
or U14095 (N_14095,N_10979,N_9895);
nor U14096 (N_14096,N_9988,N_11527);
nor U14097 (N_14097,N_11186,N_9627);
and U14098 (N_14098,N_11462,N_11658);
xnor U14099 (N_14099,N_10869,N_11726);
and U14100 (N_14100,N_10700,N_10490);
or U14101 (N_14101,N_11834,N_11663);
xnor U14102 (N_14102,N_11866,N_10664);
nand U14103 (N_14103,N_9210,N_10582);
xnor U14104 (N_14104,N_11502,N_10534);
and U14105 (N_14105,N_11895,N_11885);
xor U14106 (N_14106,N_11794,N_11329);
and U14107 (N_14107,N_10164,N_10840);
and U14108 (N_14108,N_9534,N_11266);
or U14109 (N_14109,N_9841,N_10006);
and U14110 (N_14110,N_11303,N_9337);
xnor U14111 (N_14111,N_9383,N_11810);
nand U14112 (N_14112,N_9723,N_10960);
xnor U14113 (N_14113,N_11415,N_9567);
nor U14114 (N_14114,N_10999,N_9278);
and U14115 (N_14115,N_10420,N_10548);
xnor U14116 (N_14116,N_11094,N_10126);
or U14117 (N_14117,N_10569,N_9763);
or U14118 (N_14118,N_10032,N_9134);
and U14119 (N_14119,N_11965,N_10813);
nand U14120 (N_14120,N_11108,N_10954);
nor U14121 (N_14121,N_10161,N_10653);
and U14122 (N_14122,N_9922,N_11224);
nand U14123 (N_14123,N_9462,N_9497);
nand U14124 (N_14124,N_9115,N_10840);
xor U14125 (N_14125,N_9748,N_9713);
or U14126 (N_14126,N_10912,N_10825);
nand U14127 (N_14127,N_9910,N_10757);
nand U14128 (N_14128,N_11703,N_9618);
nand U14129 (N_14129,N_11836,N_10784);
nor U14130 (N_14130,N_11487,N_10805);
nor U14131 (N_14131,N_11384,N_9980);
or U14132 (N_14132,N_9982,N_10978);
and U14133 (N_14133,N_11689,N_11405);
nor U14134 (N_14134,N_10343,N_9841);
or U14135 (N_14135,N_10176,N_9748);
and U14136 (N_14136,N_11656,N_9715);
or U14137 (N_14137,N_9430,N_10496);
nor U14138 (N_14138,N_9368,N_10549);
or U14139 (N_14139,N_11684,N_10862);
xnor U14140 (N_14140,N_9284,N_11443);
nand U14141 (N_14141,N_10631,N_9216);
nand U14142 (N_14142,N_11617,N_9666);
or U14143 (N_14143,N_11874,N_11242);
nor U14144 (N_14144,N_9433,N_9186);
nand U14145 (N_14145,N_11461,N_11388);
nor U14146 (N_14146,N_11157,N_9436);
and U14147 (N_14147,N_10197,N_9808);
or U14148 (N_14148,N_11535,N_10595);
nor U14149 (N_14149,N_10491,N_11118);
nor U14150 (N_14150,N_9950,N_11768);
nor U14151 (N_14151,N_10024,N_10544);
xnor U14152 (N_14152,N_9090,N_10759);
nor U14153 (N_14153,N_11442,N_9151);
nand U14154 (N_14154,N_11472,N_9972);
and U14155 (N_14155,N_11424,N_10964);
nor U14156 (N_14156,N_10976,N_9747);
or U14157 (N_14157,N_11939,N_9330);
or U14158 (N_14158,N_11724,N_11537);
or U14159 (N_14159,N_9816,N_9771);
and U14160 (N_14160,N_11788,N_11439);
xor U14161 (N_14161,N_10453,N_11803);
and U14162 (N_14162,N_11669,N_10665);
and U14163 (N_14163,N_11391,N_11494);
nor U14164 (N_14164,N_9631,N_11471);
xnor U14165 (N_14165,N_9081,N_10414);
nor U14166 (N_14166,N_11059,N_10866);
xor U14167 (N_14167,N_11193,N_11620);
nor U14168 (N_14168,N_11205,N_11626);
xor U14169 (N_14169,N_9898,N_9672);
nor U14170 (N_14170,N_11450,N_10688);
nand U14171 (N_14171,N_10690,N_9222);
nand U14172 (N_14172,N_10366,N_11832);
xnor U14173 (N_14173,N_10248,N_11806);
xnor U14174 (N_14174,N_11978,N_11208);
nor U14175 (N_14175,N_11149,N_10827);
nand U14176 (N_14176,N_9696,N_11657);
nand U14177 (N_14177,N_9601,N_11863);
nand U14178 (N_14178,N_11148,N_9603);
or U14179 (N_14179,N_10931,N_9659);
xnor U14180 (N_14180,N_10459,N_10747);
nand U14181 (N_14181,N_10072,N_10743);
or U14182 (N_14182,N_9103,N_11065);
and U14183 (N_14183,N_11816,N_11041);
or U14184 (N_14184,N_10175,N_10652);
nand U14185 (N_14185,N_9949,N_10488);
nand U14186 (N_14186,N_10311,N_10233);
or U14187 (N_14187,N_9378,N_10997);
xnor U14188 (N_14188,N_10984,N_11855);
or U14189 (N_14189,N_9775,N_10431);
xnor U14190 (N_14190,N_11181,N_10313);
xnor U14191 (N_14191,N_11586,N_11307);
nand U14192 (N_14192,N_10102,N_10288);
or U14193 (N_14193,N_11815,N_11066);
and U14194 (N_14194,N_9710,N_9371);
nor U14195 (N_14195,N_11385,N_9942);
nor U14196 (N_14196,N_9849,N_9918);
xor U14197 (N_14197,N_11829,N_10990);
or U14198 (N_14198,N_10968,N_9908);
nor U14199 (N_14199,N_11625,N_9760);
nand U14200 (N_14200,N_10191,N_11992);
xor U14201 (N_14201,N_11503,N_10924);
xor U14202 (N_14202,N_10985,N_9950);
nor U14203 (N_14203,N_9637,N_11350);
or U14204 (N_14204,N_10689,N_10010);
xnor U14205 (N_14205,N_9945,N_10508);
nand U14206 (N_14206,N_11562,N_9615);
or U14207 (N_14207,N_10690,N_10993);
or U14208 (N_14208,N_9063,N_10748);
nor U14209 (N_14209,N_9539,N_11834);
nand U14210 (N_14210,N_9268,N_11513);
nor U14211 (N_14211,N_10724,N_11178);
or U14212 (N_14212,N_11919,N_10431);
xor U14213 (N_14213,N_11463,N_11705);
or U14214 (N_14214,N_10096,N_9264);
or U14215 (N_14215,N_9570,N_10126);
nor U14216 (N_14216,N_11891,N_10214);
or U14217 (N_14217,N_9750,N_10982);
nand U14218 (N_14218,N_11848,N_11637);
and U14219 (N_14219,N_11392,N_9387);
or U14220 (N_14220,N_9241,N_10260);
nand U14221 (N_14221,N_10772,N_11272);
and U14222 (N_14222,N_9868,N_9213);
xor U14223 (N_14223,N_10052,N_9233);
nor U14224 (N_14224,N_11209,N_11758);
and U14225 (N_14225,N_9971,N_9460);
or U14226 (N_14226,N_11509,N_11655);
nor U14227 (N_14227,N_9473,N_10483);
or U14228 (N_14228,N_10721,N_11553);
xor U14229 (N_14229,N_9873,N_11161);
or U14230 (N_14230,N_10618,N_10477);
nor U14231 (N_14231,N_9239,N_11556);
nor U14232 (N_14232,N_11703,N_11063);
and U14233 (N_14233,N_10749,N_11422);
and U14234 (N_14234,N_10984,N_11269);
or U14235 (N_14235,N_10972,N_11058);
or U14236 (N_14236,N_11630,N_11433);
or U14237 (N_14237,N_11462,N_11389);
and U14238 (N_14238,N_11295,N_10933);
nor U14239 (N_14239,N_11934,N_10805);
or U14240 (N_14240,N_11972,N_9202);
or U14241 (N_14241,N_11797,N_11881);
or U14242 (N_14242,N_10460,N_9183);
nor U14243 (N_14243,N_10814,N_11359);
or U14244 (N_14244,N_11816,N_9254);
or U14245 (N_14245,N_9271,N_11271);
and U14246 (N_14246,N_11937,N_10780);
xor U14247 (N_14247,N_11223,N_9789);
or U14248 (N_14248,N_9397,N_11091);
nor U14249 (N_14249,N_10365,N_11950);
xor U14250 (N_14250,N_11489,N_11848);
nand U14251 (N_14251,N_11959,N_9375);
and U14252 (N_14252,N_10063,N_11253);
and U14253 (N_14253,N_11322,N_10222);
or U14254 (N_14254,N_9456,N_9502);
or U14255 (N_14255,N_10460,N_9179);
xor U14256 (N_14256,N_10576,N_9378);
xnor U14257 (N_14257,N_9634,N_9368);
or U14258 (N_14258,N_10324,N_9460);
or U14259 (N_14259,N_11604,N_10626);
nand U14260 (N_14260,N_11916,N_11065);
nor U14261 (N_14261,N_9449,N_10862);
nand U14262 (N_14262,N_10933,N_11851);
xor U14263 (N_14263,N_9764,N_9802);
or U14264 (N_14264,N_9407,N_11254);
xnor U14265 (N_14265,N_11171,N_10786);
or U14266 (N_14266,N_9784,N_9462);
nand U14267 (N_14267,N_11002,N_11513);
nand U14268 (N_14268,N_11214,N_11840);
xor U14269 (N_14269,N_9328,N_9745);
xor U14270 (N_14270,N_10123,N_10795);
and U14271 (N_14271,N_10043,N_11365);
nand U14272 (N_14272,N_10452,N_10922);
nand U14273 (N_14273,N_11477,N_10170);
xor U14274 (N_14274,N_10243,N_11540);
xnor U14275 (N_14275,N_11323,N_9560);
or U14276 (N_14276,N_10649,N_9249);
nand U14277 (N_14277,N_11715,N_10121);
or U14278 (N_14278,N_10733,N_10135);
nand U14279 (N_14279,N_9695,N_9791);
nor U14280 (N_14280,N_11736,N_11094);
xor U14281 (N_14281,N_9798,N_11302);
xnor U14282 (N_14282,N_11668,N_9906);
or U14283 (N_14283,N_9371,N_10249);
xor U14284 (N_14284,N_10681,N_9573);
nor U14285 (N_14285,N_10188,N_10780);
nor U14286 (N_14286,N_10703,N_9447);
or U14287 (N_14287,N_11871,N_10538);
and U14288 (N_14288,N_9930,N_10281);
and U14289 (N_14289,N_11312,N_11879);
nor U14290 (N_14290,N_11910,N_9397);
or U14291 (N_14291,N_9293,N_9828);
and U14292 (N_14292,N_9381,N_11091);
nor U14293 (N_14293,N_10575,N_11439);
or U14294 (N_14294,N_11065,N_9208);
or U14295 (N_14295,N_10102,N_11301);
or U14296 (N_14296,N_10012,N_9702);
nor U14297 (N_14297,N_11556,N_11195);
and U14298 (N_14298,N_9875,N_9252);
xnor U14299 (N_14299,N_10030,N_11028);
nor U14300 (N_14300,N_11934,N_10095);
xor U14301 (N_14301,N_11670,N_10718);
nand U14302 (N_14302,N_10488,N_9843);
nor U14303 (N_14303,N_11619,N_10154);
nor U14304 (N_14304,N_11772,N_9931);
xor U14305 (N_14305,N_9430,N_9262);
nand U14306 (N_14306,N_9314,N_10069);
xnor U14307 (N_14307,N_11260,N_10756);
and U14308 (N_14308,N_9727,N_10897);
nor U14309 (N_14309,N_9357,N_11619);
xnor U14310 (N_14310,N_11296,N_10040);
nand U14311 (N_14311,N_9956,N_10586);
and U14312 (N_14312,N_11036,N_9365);
nor U14313 (N_14313,N_9551,N_9184);
nor U14314 (N_14314,N_10858,N_9034);
and U14315 (N_14315,N_10650,N_9366);
nand U14316 (N_14316,N_10820,N_10725);
xnor U14317 (N_14317,N_11870,N_9223);
nand U14318 (N_14318,N_10939,N_9608);
or U14319 (N_14319,N_9771,N_10183);
or U14320 (N_14320,N_9849,N_10509);
or U14321 (N_14321,N_11133,N_10225);
nor U14322 (N_14322,N_9054,N_11328);
nor U14323 (N_14323,N_9057,N_11206);
nand U14324 (N_14324,N_11770,N_11418);
xnor U14325 (N_14325,N_9236,N_9868);
or U14326 (N_14326,N_9922,N_9391);
and U14327 (N_14327,N_9287,N_11798);
xnor U14328 (N_14328,N_10820,N_9481);
nand U14329 (N_14329,N_10575,N_10843);
xnor U14330 (N_14330,N_10710,N_10012);
or U14331 (N_14331,N_10922,N_10328);
or U14332 (N_14332,N_11129,N_9021);
nor U14333 (N_14333,N_10152,N_9703);
or U14334 (N_14334,N_11301,N_10429);
or U14335 (N_14335,N_9167,N_11218);
or U14336 (N_14336,N_10460,N_11778);
and U14337 (N_14337,N_11279,N_11837);
and U14338 (N_14338,N_10354,N_11607);
nor U14339 (N_14339,N_10191,N_9651);
nand U14340 (N_14340,N_9158,N_10823);
xor U14341 (N_14341,N_9993,N_10919);
or U14342 (N_14342,N_11133,N_10080);
nor U14343 (N_14343,N_11291,N_11005);
or U14344 (N_14344,N_9933,N_10422);
or U14345 (N_14345,N_11103,N_9097);
and U14346 (N_14346,N_10783,N_10158);
or U14347 (N_14347,N_9730,N_11737);
xnor U14348 (N_14348,N_10662,N_9674);
xnor U14349 (N_14349,N_11584,N_11184);
xnor U14350 (N_14350,N_11898,N_10340);
nor U14351 (N_14351,N_11193,N_11823);
nor U14352 (N_14352,N_10289,N_9286);
or U14353 (N_14353,N_10775,N_10888);
and U14354 (N_14354,N_10957,N_10628);
xor U14355 (N_14355,N_9882,N_11418);
and U14356 (N_14356,N_9570,N_10769);
nand U14357 (N_14357,N_9783,N_10957);
nand U14358 (N_14358,N_9832,N_11754);
nand U14359 (N_14359,N_10113,N_11565);
or U14360 (N_14360,N_10886,N_10749);
xnor U14361 (N_14361,N_11974,N_11256);
and U14362 (N_14362,N_11298,N_9315);
nand U14363 (N_14363,N_10900,N_11349);
and U14364 (N_14364,N_10111,N_9218);
xnor U14365 (N_14365,N_9142,N_9507);
nor U14366 (N_14366,N_10038,N_11623);
and U14367 (N_14367,N_11219,N_10739);
xnor U14368 (N_14368,N_10459,N_11641);
nand U14369 (N_14369,N_11466,N_11289);
nand U14370 (N_14370,N_10961,N_11966);
xor U14371 (N_14371,N_10209,N_9161);
nor U14372 (N_14372,N_10483,N_10618);
nand U14373 (N_14373,N_10702,N_11547);
or U14374 (N_14374,N_11669,N_9261);
or U14375 (N_14375,N_9088,N_9160);
and U14376 (N_14376,N_11711,N_10988);
nand U14377 (N_14377,N_11244,N_9291);
nand U14378 (N_14378,N_11140,N_10742);
or U14379 (N_14379,N_11259,N_9993);
xor U14380 (N_14380,N_10926,N_9517);
or U14381 (N_14381,N_10120,N_9527);
xor U14382 (N_14382,N_10258,N_10281);
and U14383 (N_14383,N_9838,N_10226);
or U14384 (N_14384,N_9882,N_11842);
nor U14385 (N_14385,N_10041,N_10694);
or U14386 (N_14386,N_9527,N_9192);
xor U14387 (N_14387,N_11298,N_11365);
or U14388 (N_14388,N_11177,N_10969);
nand U14389 (N_14389,N_11982,N_11221);
nor U14390 (N_14390,N_11517,N_9141);
nor U14391 (N_14391,N_10789,N_11329);
and U14392 (N_14392,N_11978,N_9439);
or U14393 (N_14393,N_10679,N_10422);
or U14394 (N_14394,N_9295,N_9032);
nor U14395 (N_14395,N_10647,N_11278);
and U14396 (N_14396,N_9110,N_10736);
and U14397 (N_14397,N_10797,N_11792);
or U14398 (N_14398,N_9245,N_10583);
xor U14399 (N_14399,N_11307,N_11022);
or U14400 (N_14400,N_10630,N_11183);
xor U14401 (N_14401,N_10342,N_11869);
nor U14402 (N_14402,N_10195,N_11513);
xnor U14403 (N_14403,N_11549,N_10812);
xor U14404 (N_14404,N_11050,N_9426);
and U14405 (N_14405,N_11774,N_10481);
and U14406 (N_14406,N_11365,N_11145);
or U14407 (N_14407,N_11345,N_9786);
nor U14408 (N_14408,N_10071,N_9497);
nand U14409 (N_14409,N_10219,N_9746);
xor U14410 (N_14410,N_11860,N_10917);
and U14411 (N_14411,N_10191,N_11889);
and U14412 (N_14412,N_10235,N_9427);
nor U14413 (N_14413,N_9730,N_9364);
and U14414 (N_14414,N_10374,N_11161);
nor U14415 (N_14415,N_9644,N_10761);
and U14416 (N_14416,N_9019,N_10114);
nor U14417 (N_14417,N_9001,N_10821);
or U14418 (N_14418,N_11919,N_11746);
xor U14419 (N_14419,N_10167,N_9728);
nor U14420 (N_14420,N_9111,N_10055);
nand U14421 (N_14421,N_10488,N_11095);
nor U14422 (N_14422,N_9907,N_11693);
or U14423 (N_14423,N_11359,N_10433);
nor U14424 (N_14424,N_11316,N_9967);
nand U14425 (N_14425,N_9595,N_9242);
or U14426 (N_14426,N_11184,N_9132);
or U14427 (N_14427,N_10749,N_11904);
nor U14428 (N_14428,N_11924,N_11378);
and U14429 (N_14429,N_10016,N_9708);
nand U14430 (N_14430,N_9574,N_9803);
or U14431 (N_14431,N_9951,N_9405);
nand U14432 (N_14432,N_9406,N_10460);
and U14433 (N_14433,N_9352,N_11299);
and U14434 (N_14434,N_11504,N_9469);
nor U14435 (N_14435,N_9785,N_10060);
or U14436 (N_14436,N_10393,N_11612);
or U14437 (N_14437,N_11599,N_11161);
nor U14438 (N_14438,N_9043,N_11839);
and U14439 (N_14439,N_9475,N_11538);
and U14440 (N_14440,N_9767,N_9074);
nand U14441 (N_14441,N_11610,N_10599);
nand U14442 (N_14442,N_10788,N_10272);
xor U14443 (N_14443,N_11482,N_10987);
xor U14444 (N_14444,N_11060,N_9576);
nor U14445 (N_14445,N_11767,N_9921);
and U14446 (N_14446,N_11749,N_11316);
xor U14447 (N_14447,N_9448,N_11494);
xnor U14448 (N_14448,N_9406,N_9116);
or U14449 (N_14449,N_9447,N_11359);
nand U14450 (N_14450,N_10261,N_9635);
nor U14451 (N_14451,N_10547,N_10740);
or U14452 (N_14452,N_9698,N_10636);
nor U14453 (N_14453,N_9642,N_11232);
xnor U14454 (N_14454,N_10889,N_11733);
nor U14455 (N_14455,N_11914,N_11348);
nor U14456 (N_14456,N_10175,N_9251);
or U14457 (N_14457,N_11633,N_10801);
nor U14458 (N_14458,N_10174,N_11948);
nor U14459 (N_14459,N_9392,N_10812);
nand U14460 (N_14460,N_10577,N_10399);
xnor U14461 (N_14461,N_9122,N_9334);
xnor U14462 (N_14462,N_11088,N_10282);
or U14463 (N_14463,N_9114,N_11621);
and U14464 (N_14464,N_11963,N_11172);
nand U14465 (N_14465,N_10180,N_10957);
and U14466 (N_14466,N_11129,N_11554);
nor U14467 (N_14467,N_9613,N_11100);
xor U14468 (N_14468,N_9316,N_9679);
nand U14469 (N_14469,N_9410,N_9164);
nand U14470 (N_14470,N_10953,N_11429);
xnor U14471 (N_14471,N_10410,N_9386);
nand U14472 (N_14472,N_11532,N_11018);
nor U14473 (N_14473,N_11754,N_11815);
xnor U14474 (N_14474,N_9141,N_9928);
or U14475 (N_14475,N_10496,N_10193);
and U14476 (N_14476,N_9294,N_11621);
nor U14477 (N_14477,N_10656,N_10264);
or U14478 (N_14478,N_11614,N_9967);
nor U14479 (N_14479,N_10924,N_11104);
or U14480 (N_14480,N_10155,N_9084);
nor U14481 (N_14481,N_10607,N_9468);
nand U14482 (N_14482,N_11040,N_11479);
nand U14483 (N_14483,N_10291,N_10311);
xor U14484 (N_14484,N_9041,N_10134);
nor U14485 (N_14485,N_10169,N_11517);
nor U14486 (N_14486,N_9050,N_11473);
nand U14487 (N_14487,N_10663,N_9715);
nor U14488 (N_14488,N_9159,N_11859);
or U14489 (N_14489,N_9132,N_10369);
nor U14490 (N_14490,N_10796,N_10802);
xnor U14491 (N_14491,N_9688,N_9684);
nor U14492 (N_14492,N_11285,N_10192);
xor U14493 (N_14493,N_9634,N_10288);
nand U14494 (N_14494,N_9464,N_11530);
or U14495 (N_14495,N_11432,N_9047);
and U14496 (N_14496,N_11110,N_10482);
xnor U14497 (N_14497,N_9252,N_9800);
or U14498 (N_14498,N_9271,N_9848);
xor U14499 (N_14499,N_10711,N_11742);
xor U14500 (N_14500,N_9151,N_9691);
and U14501 (N_14501,N_9164,N_9258);
and U14502 (N_14502,N_10646,N_10112);
or U14503 (N_14503,N_9171,N_11555);
nand U14504 (N_14504,N_11095,N_11885);
and U14505 (N_14505,N_10171,N_10193);
xor U14506 (N_14506,N_9999,N_11572);
or U14507 (N_14507,N_9722,N_10563);
nand U14508 (N_14508,N_11199,N_10873);
or U14509 (N_14509,N_10655,N_9188);
and U14510 (N_14510,N_11342,N_10409);
or U14511 (N_14511,N_11233,N_10502);
and U14512 (N_14512,N_10044,N_9143);
or U14513 (N_14513,N_10522,N_11730);
nand U14514 (N_14514,N_10359,N_10781);
or U14515 (N_14515,N_9477,N_10206);
nor U14516 (N_14516,N_9670,N_10395);
nor U14517 (N_14517,N_10266,N_10779);
and U14518 (N_14518,N_9034,N_11879);
and U14519 (N_14519,N_11248,N_11195);
or U14520 (N_14520,N_10968,N_11071);
and U14521 (N_14521,N_10949,N_9020);
nand U14522 (N_14522,N_9721,N_11689);
nand U14523 (N_14523,N_10409,N_9153);
and U14524 (N_14524,N_10050,N_10953);
nor U14525 (N_14525,N_11901,N_10993);
nand U14526 (N_14526,N_10840,N_9206);
nand U14527 (N_14527,N_10164,N_11360);
and U14528 (N_14528,N_11804,N_9407);
xnor U14529 (N_14529,N_11675,N_9174);
and U14530 (N_14530,N_9117,N_10262);
nor U14531 (N_14531,N_9914,N_10106);
xor U14532 (N_14532,N_11036,N_9130);
nor U14533 (N_14533,N_10811,N_10572);
xor U14534 (N_14534,N_11932,N_9699);
and U14535 (N_14535,N_10573,N_9853);
nand U14536 (N_14536,N_10139,N_11585);
nor U14537 (N_14537,N_9664,N_10489);
nand U14538 (N_14538,N_10431,N_9573);
or U14539 (N_14539,N_9761,N_9990);
or U14540 (N_14540,N_10794,N_10259);
xor U14541 (N_14541,N_11102,N_9483);
nand U14542 (N_14542,N_11832,N_11264);
nor U14543 (N_14543,N_9094,N_9041);
xor U14544 (N_14544,N_11932,N_10106);
and U14545 (N_14545,N_11193,N_10317);
or U14546 (N_14546,N_11135,N_9859);
or U14547 (N_14547,N_9565,N_10015);
or U14548 (N_14548,N_11337,N_11593);
or U14549 (N_14549,N_11591,N_11678);
and U14550 (N_14550,N_10652,N_9743);
and U14551 (N_14551,N_10586,N_11145);
and U14552 (N_14552,N_9974,N_9208);
and U14553 (N_14553,N_10566,N_9540);
or U14554 (N_14554,N_10160,N_9908);
and U14555 (N_14555,N_9694,N_9005);
nor U14556 (N_14556,N_9821,N_11542);
nor U14557 (N_14557,N_10735,N_10674);
xnor U14558 (N_14558,N_10947,N_9109);
xnor U14559 (N_14559,N_9644,N_9208);
nand U14560 (N_14560,N_11389,N_9358);
nand U14561 (N_14561,N_10486,N_9831);
or U14562 (N_14562,N_9956,N_9740);
nand U14563 (N_14563,N_9066,N_11909);
and U14564 (N_14564,N_11721,N_9278);
and U14565 (N_14565,N_10873,N_11440);
and U14566 (N_14566,N_10235,N_10028);
or U14567 (N_14567,N_11629,N_11404);
nand U14568 (N_14568,N_11992,N_11392);
and U14569 (N_14569,N_10233,N_11374);
and U14570 (N_14570,N_10980,N_9487);
or U14571 (N_14571,N_11447,N_11338);
nand U14572 (N_14572,N_10049,N_10119);
nand U14573 (N_14573,N_10090,N_9882);
and U14574 (N_14574,N_11259,N_11832);
and U14575 (N_14575,N_9211,N_10696);
and U14576 (N_14576,N_9018,N_11514);
nor U14577 (N_14577,N_9251,N_11688);
xnor U14578 (N_14578,N_11239,N_11803);
or U14579 (N_14579,N_9463,N_10090);
and U14580 (N_14580,N_11212,N_11893);
and U14581 (N_14581,N_11317,N_10262);
or U14582 (N_14582,N_9588,N_9668);
or U14583 (N_14583,N_11007,N_9205);
or U14584 (N_14584,N_9945,N_11856);
nor U14585 (N_14585,N_10950,N_9625);
nand U14586 (N_14586,N_9462,N_9049);
or U14587 (N_14587,N_10087,N_11818);
xor U14588 (N_14588,N_11136,N_9229);
and U14589 (N_14589,N_11491,N_10237);
nand U14590 (N_14590,N_11280,N_10103);
nor U14591 (N_14591,N_11988,N_9745);
xnor U14592 (N_14592,N_10522,N_10800);
nor U14593 (N_14593,N_11964,N_9702);
xor U14594 (N_14594,N_10277,N_10955);
and U14595 (N_14595,N_9423,N_9673);
and U14596 (N_14596,N_11821,N_9207);
or U14597 (N_14597,N_9165,N_9442);
nand U14598 (N_14598,N_10377,N_9780);
nor U14599 (N_14599,N_9923,N_11708);
or U14600 (N_14600,N_11997,N_9614);
or U14601 (N_14601,N_10867,N_9653);
nand U14602 (N_14602,N_10937,N_9537);
nor U14603 (N_14603,N_10407,N_11238);
and U14604 (N_14604,N_11296,N_11833);
xnor U14605 (N_14605,N_10260,N_10803);
nand U14606 (N_14606,N_11988,N_10470);
xnor U14607 (N_14607,N_10051,N_10845);
nor U14608 (N_14608,N_11036,N_10315);
nor U14609 (N_14609,N_9049,N_11598);
and U14610 (N_14610,N_10970,N_10729);
and U14611 (N_14611,N_9299,N_10401);
and U14612 (N_14612,N_11071,N_9938);
xnor U14613 (N_14613,N_9319,N_10818);
nand U14614 (N_14614,N_11033,N_11283);
nor U14615 (N_14615,N_9885,N_11441);
nand U14616 (N_14616,N_11307,N_11638);
xor U14617 (N_14617,N_10644,N_10012);
and U14618 (N_14618,N_11012,N_11238);
or U14619 (N_14619,N_9244,N_11736);
nand U14620 (N_14620,N_11687,N_9074);
nor U14621 (N_14621,N_9162,N_10007);
xor U14622 (N_14622,N_10934,N_11008);
or U14623 (N_14623,N_9154,N_11057);
nand U14624 (N_14624,N_9315,N_11354);
nand U14625 (N_14625,N_10009,N_9361);
or U14626 (N_14626,N_11980,N_11662);
or U14627 (N_14627,N_9062,N_11044);
nor U14628 (N_14628,N_10351,N_10846);
nand U14629 (N_14629,N_11561,N_10148);
nor U14630 (N_14630,N_10849,N_9177);
and U14631 (N_14631,N_10065,N_9706);
or U14632 (N_14632,N_9247,N_10148);
nand U14633 (N_14633,N_9325,N_9976);
nand U14634 (N_14634,N_10713,N_9326);
and U14635 (N_14635,N_10717,N_10545);
or U14636 (N_14636,N_10571,N_11481);
nor U14637 (N_14637,N_11012,N_11355);
nand U14638 (N_14638,N_11445,N_10758);
xor U14639 (N_14639,N_10795,N_9210);
nand U14640 (N_14640,N_11951,N_10639);
and U14641 (N_14641,N_11033,N_9583);
xnor U14642 (N_14642,N_11827,N_11790);
and U14643 (N_14643,N_9353,N_9051);
xnor U14644 (N_14644,N_10613,N_11293);
and U14645 (N_14645,N_9574,N_11932);
nor U14646 (N_14646,N_11873,N_10509);
and U14647 (N_14647,N_11886,N_10058);
or U14648 (N_14648,N_11702,N_10977);
and U14649 (N_14649,N_10181,N_11710);
nand U14650 (N_14650,N_9575,N_9865);
xnor U14651 (N_14651,N_11002,N_11108);
nand U14652 (N_14652,N_10006,N_11713);
nor U14653 (N_14653,N_10855,N_11169);
and U14654 (N_14654,N_10686,N_10812);
xnor U14655 (N_14655,N_10022,N_11700);
or U14656 (N_14656,N_10172,N_9037);
or U14657 (N_14657,N_9722,N_9240);
nand U14658 (N_14658,N_9065,N_9101);
nor U14659 (N_14659,N_11781,N_10700);
xnor U14660 (N_14660,N_10756,N_10487);
nand U14661 (N_14661,N_9085,N_9081);
nor U14662 (N_14662,N_10875,N_11846);
or U14663 (N_14663,N_11780,N_10885);
and U14664 (N_14664,N_11791,N_11698);
and U14665 (N_14665,N_9698,N_9883);
or U14666 (N_14666,N_10952,N_11695);
and U14667 (N_14667,N_10539,N_10374);
xor U14668 (N_14668,N_10718,N_9954);
nand U14669 (N_14669,N_9560,N_11102);
nor U14670 (N_14670,N_10454,N_9975);
and U14671 (N_14671,N_10842,N_9148);
nor U14672 (N_14672,N_11327,N_9893);
or U14673 (N_14673,N_9819,N_10038);
xor U14674 (N_14674,N_11768,N_10134);
or U14675 (N_14675,N_10542,N_10732);
nor U14676 (N_14676,N_9202,N_10071);
nand U14677 (N_14677,N_9514,N_9831);
nor U14678 (N_14678,N_9764,N_10604);
or U14679 (N_14679,N_11814,N_10488);
xnor U14680 (N_14680,N_9978,N_9733);
or U14681 (N_14681,N_10943,N_11022);
and U14682 (N_14682,N_9417,N_9477);
nor U14683 (N_14683,N_10600,N_11301);
or U14684 (N_14684,N_10151,N_9563);
xor U14685 (N_14685,N_9138,N_10662);
xnor U14686 (N_14686,N_11171,N_9433);
xnor U14687 (N_14687,N_10194,N_9272);
xnor U14688 (N_14688,N_11202,N_9251);
nor U14689 (N_14689,N_11879,N_11931);
nor U14690 (N_14690,N_10395,N_11538);
and U14691 (N_14691,N_10904,N_10814);
nor U14692 (N_14692,N_10737,N_10953);
xor U14693 (N_14693,N_9299,N_9521);
nor U14694 (N_14694,N_11113,N_9697);
nand U14695 (N_14695,N_9925,N_11663);
and U14696 (N_14696,N_9931,N_9655);
nor U14697 (N_14697,N_10558,N_9277);
and U14698 (N_14698,N_10275,N_10083);
nand U14699 (N_14699,N_9905,N_9409);
xor U14700 (N_14700,N_9545,N_10469);
xor U14701 (N_14701,N_9186,N_11280);
and U14702 (N_14702,N_10289,N_9157);
and U14703 (N_14703,N_9531,N_9156);
nor U14704 (N_14704,N_11892,N_11494);
or U14705 (N_14705,N_9941,N_10936);
and U14706 (N_14706,N_11843,N_10818);
or U14707 (N_14707,N_9850,N_9471);
or U14708 (N_14708,N_10744,N_10029);
xor U14709 (N_14709,N_11471,N_11684);
or U14710 (N_14710,N_10369,N_11781);
or U14711 (N_14711,N_10366,N_9711);
and U14712 (N_14712,N_10386,N_11643);
nor U14713 (N_14713,N_9516,N_11576);
or U14714 (N_14714,N_10310,N_10670);
xor U14715 (N_14715,N_10554,N_10537);
nor U14716 (N_14716,N_10175,N_9725);
or U14717 (N_14717,N_9186,N_11473);
and U14718 (N_14718,N_10882,N_9602);
or U14719 (N_14719,N_11472,N_9907);
xnor U14720 (N_14720,N_9831,N_9378);
xnor U14721 (N_14721,N_9656,N_10996);
or U14722 (N_14722,N_10968,N_10826);
or U14723 (N_14723,N_11292,N_11539);
or U14724 (N_14724,N_10720,N_11865);
or U14725 (N_14725,N_9866,N_11770);
xor U14726 (N_14726,N_9065,N_10712);
or U14727 (N_14727,N_11832,N_9751);
and U14728 (N_14728,N_10473,N_11550);
and U14729 (N_14729,N_9884,N_11399);
nand U14730 (N_14730,N_10664,N_10040);
nand U14731 (N_14731,N_11985,N_10893);
nand U14732 (N_14732,N_10327,N_11124);
or U14733 (N_14733,N_11810,N_9102);
xnor U14734 (N_14734,N_9293,N_10566);
nand U14735 (N_14735,N_11661,N_11893);
or U14736 (N_14736,N_9526,N_10889);
nor U14737 (N_14737,N_11425,N_9117);
nand U14738 (N_14738,N_11270,N_11861);
xnor U14739 (N_14739,N_9855,N_11982);
and U14740 (N_14740,N_9161,N_11387);
or U14741 (N_14741,N_9135,N_9871);
nand U14742 (N_14742,N_9109,N_11051);
nand U14743 (N_14743,N_10719,N_10289);
and U14744 (N_14744,N_11407,N_11510);
nand U14745 (N_14745,N_10245,N_11284);
and U14746 (N_14746,N_10910,N_10202);
nand U14747 (N_14747,N_10825,N_10242);
nor U14748 (N_14748,N_11569,N_10295);
and U14749 (N_14749,N_11116,N_11254);
nor U14750 (N_14750,N_9728,N_11714);
nor U14751 (N_14751,N_9177,N_10680);
xnor U14752 (N_14752,N_11346,N_11355);
xor U14753 (N_14753,N_10285,N_10166);
and U14754 (N_14754,N_11292,N_9648);
and U14755 (N_14755,N_9688,N_10380);
or U14756 (N_14756,N_10409,N_11814);
xnor U14757 (N_14757,N_10589,N_10264);
nor U14758 (N_14758,N_11451,N_11030);
nor U14759 (N_14759,N_10967,N_11156);
or U14760 (N_14760,N_10366,N_11612);
nor U14761 (N_14761,N_10537,N_10222);
nand U14762 (N_14762,N_9681,N_9243);
and U14763 (N_14763,N_9736,N_10069);
nor U14764 (N_14764,N_10655,N_11065);
nor U14765 (N_14765,N_11477,N_11619);
nand U14766 (N_14766,N_9361,N_9688);
nor U14767 (N_14767,N_10127,N_9575);
nor U14768 (N_14768,N_11134,N_11551);
and U14769 (N_14769,N_10669,N_9809);
nor U14770 (N_14770,N_9716,N_9851);
or U14771 (N_14771,N_10053,N_10168);
and U14772 (N_14772,N_9062,N_10084);
and U14773 (N_14773,N_10769,N_10385);
xnor U14774 (N_14774,N_11495,N_10576);
or U14775 (N_14775,N_11075,N_9214);
xnor U14776 (N_14776,N_9864,N_10331);
and U14777 (N_14777,N_9249,N_9143);
or U14778 (N_14778,N_11841,N_10456);
nand U14779 (N_14779,N_11347,N_10079);
or U14780 (N_14780,N_11910,N_11626);
and U14781 (N_14781,N_9918,N_10380);
xnor U14782 (N_14782,N_9244,N_9786);
or U14783 (N_14783,N_10069,N_10228);
and U14784 (N_14784,N_10322,N_10873);
xnor U14785 (N_14785,N_9456,N_10921);
nor U14786 (N_14786,N_11182,N_11014);
nor U14787 (N_14787,N_11989,N_10408);
nor U14788 (N_14788,N_11473,N_9925);
nand U14789 (N_14789,N_11512,N_11609);
and U14790 (N_14790,N_11203,N_9656);
nand U14791 (N_14791,N_10440,N_9379);
nor U14792 (N_14792,N_11999,N_10261);
and U14793 (N_14793,N_11923,N_9794);
or U14794 (N_14794,N_9872,N_9231);
and U14795 (N_14795,N_11178,N_9150);
or U14796 (N_14796,N_11495,N_10021);
and U14797 (N_14797,N_9064,N_11955);
xnor U14798 (N_14798,N_11530,N_9697);
or U14799 (N_14799,N_11591,N_11524);
nor U14800 (N_14800,N_9996,N_10936);
xnor U14801 (N_14801,N_11972,N_9184);
and U14802 (N_14802,N_9613,N_10069);
nand U14803 (N_14803,N_10441,N_10462);
nor U14804 (N_14804,N_9467,N_11515);
or U14805 (N_14805,N_9932,N_11353);
or U14806 (N_14806,N_9815,N_11219);
or U14807 (N_14807,N_11702,N_10935);
nand U14808 (N_14808,N_9136,N_10825);
and U14809 (N_14809,N_11299,N_9612);
and U14810 (N_14810,N_11461,N_9397);
nand U14811 (N_14811,N_11471,N_10555);
xnor U14812 (N_14812,N_11762,N_9710);
and U14813 (N_14813,N_11831,N_9020);
nand U14814 (N_14814,N_10689,N_10535);
and U14815 (N_14815,N_10315,N_11660);
xnor U14816 (N_14816,N_10351,N_11923);
xor U14817 (N_14817,N_11496,N_10613);
or U14818 (N_14818,N_9591,N_10860);
nor U14819 (N_14819,N_10747,N_10501);
or U14820 (N_14820,N_11153,N_9991);
or U14821 (N_14821,N_10910,N_10541);
or U14822 (N_14822,N_9237,N_10476);
xor U14823 (N_14823,N_9098,N_10757);
nor U14824 (N_14824,N_9702,N_10389);
or U14825 (N_14825,N_9421,N_10421);
nor U14826 (N_14826,N_10346,N_10557);
nor U14827 (N_14827,N_9301,N_11429);
xor U14828 (N_14828,N_9579,N_10316);
nor U14829 (N_14829,N_11493,N_11759);
xor U14830 (N_14830,N_10009,N_10662);
nand U14831 (N_14831,N_10053,N_10771);
nand U14832 (N_14832,N_9874,N_11524);
xnor U14833 (N_14833,N_9680,N_9541);
nor U14834 (N_14834,N_11516,N_10672);
nand U14835 (N_14835,N_9674,N_9526);
xor U14836 (N_14836,N_10827,N_11742);
xnor U14837 (N_14837,N_11103,N_10674);
nor U14838 (N_14838,N_10669,N_11724);
xnor U14839 (N_14839,N_10577,N_11837);
nor U14840 (N_14840,N_9255,N_10617);
nand U14841 (N_14841,N_10900,N_11871);
xor U14842 (N_14842,N_10223,N_9789);
or U14843 (N_14843,N_11786,N_11124);
and U14844 (N_14844,N_10596,N_11499);
and U14845 (N_14845,N_9469,N_10276);
and U14846 (N_14846,N_11918,N_9328);
xnor U14847 (N_14847,N_9860,N_9233);
nand U14848 (N_14848,N_9590,N_11046);
nand U14849 (N_14849,N_11439,N_9970);
xnor U14850 (N_14850,N_9556,N_11281);
xnor U14851 (N_14851,N_9363,N_11428);
nand U14852 (N_14852,N_10156,N_9231);
and U14853 (N_14853,N_11185,N_9259);
nand U14854 (N_14854,N_11322,N_9359);
nor U14855 (N_14855,N_9708,N_9745);
nor U14856 (N_14856,N_9438,N_9640);
xor U14857 (N_14857,N_10406,N_11995);
nand U14858 (N_14858,N_11388,N_11686);
xor U14859 (N_14859,N_9557,N_11647);
nor U14860 (N_14860,N_11862,N_10766);
and U14861 (N_14861,N_9328,N_11368);
nor U14862 (N_14862,N_10094,N_10962);
and U14863 (N_14863,N_10653,N_9102);
xnor U14864 (N_14864,N_9278,N_11936);
nand U14865 (N_14865,N_11470,N_10602);
or U14866 (N_14866,N_11727,N_9881);
nor U14867 (N_14867,N_10455,N_9563);
xor U14868 (N_14868,N_9313,N_11795);
and U14869 (N_14869,N_9171,N_9834);
xor U14870 (N_14870,N_10453,N_9770);
xor U14871 (N_14871,N_9189,N_10790);
xnor U14872 (N_14872,N_9528,N_10987);
or U14873 (N_14873,N_11092,N_11781);
xnor U14874 (N_14874,N_11045,N_11016);
xor U14875 (N_14875,N_9437,N_9039);
or U14876 (N_14876,N_9638,N_11948);
and U14877 (N_14877,N_9033,N_11545);
nand U14878 (N_14878,N_11744,N_11156);
or U14879 (N_14879,N_11125,N_9227);
nor U14880 (N_14880,N_9741,N_10843);
nand U14881 (N_14881,N_10824,N_11846);
nor U14882 (N_14882,N_11250,N_10091);
or U14883 (N_14883,N_10049,N_9850);
nand U14884 (N_14884,N_11051,N_9563);
and U14885 (N_14885,N_10876,N_9081);
xor U14886 (N_14886,N_10892,N_10131);
or U14887 (N_14887,N_10901,N_10895);
or U14888 (N_14888,N_10081,N_11728);
nor U14889 (N_14889,N_10032,N_10577);
or U14890 (N_14890,N_10302,N_9152);
nand U14891 (N_14891,N_11217,N_9018);
and U14892 (N_14892,N_9742,N_10141);
or U14893 (N_14893,N_10047,N_9568);
or U14894 (N_14894,N_9133,N_10650);
xor U14895 (N_14895,N_11089,N_9718);
nor U14896 (N_14896,N_10034,N_9536);
xnor U14897 (N_14897,N_9636,N_10318);
xnor U14898 (N_14898,N_10579,N_9028);
nor U14899 (N_14899,N_11605,N_10795);
xor U14900 (N_14900,N_9399,N_9930);
or U14901 (N_14901,N_10700,N_10515);
and U14902 (N_14902,N_9997,N_11304);
xor U14903 (N_14903,N_10837,N_10465);
and U14904 (N_14904,N_11446,N_11841);
or U14905 (N_14905,N_11347,N_10738);
nand U14906 (N_14906,N_9578,N_11206);
and U14907 (N_14907,N_10739,N_11654);
nand U14908 (N_14908,N_10910,N_10583);
nand U14909 (N_14909,N_10227,N_10262);
and U14910 (N_14910,N_11514,N_11193);
nor U14911 (N_14911,N_11649,N_9640);
nor U14912 (N_14912,N_9616,N_9789);
nor U14913 (N_14913,N_9924,N_10494);
nand U14914 (N_14914,N_10635,N_10885);
nor U14915 (N_14915,N_11223,N_11097);
and U14916 (N_14916,N_10340,N_11913);
nand U14917 (N_14917,N_10855,N_10777);
nor U14918 (N_14918,N_9796,N_11118);
xnor U14919 (N_14919,N_11762,N_9085);
and U14920 (N_14920,N_11686,N_10018);
or U14921 (N_14921,N_9380,N_11034);
xnor U14922 (N_14922,N_10157,N_11848);
and U14923 (N_14923,N_10377,N_11272);
nor U14924 (N_14924,N_10905,N_9909);
or U14925 (N_14925,N_10725,N_11114);
and U14926 (N_14926,N_9143,N_10266);
nand U14927 (N_14927,N_11252,N_9626);
nand U14928 (N_14928,N_9991,N_10679);
nand U14929 (N_14929,N_10793,N_9159);
xnor U14930 (N_14930,N_10136,N_9425);
or U14931 (N_14931,N_11409,N_11896);
nand U14932 (N_14932,N_9830,N_9478);
nor U14933 (N_14933,N_9084,N_9643);
or U14934 (N_14934,N_11340,N_10272);
nor U14935 (N_14935,N_11821,N_10368);
or U14936 (N_14936,N_9909,N_11900);
nand U14937 (N_14937,N_10948,N_9623);
nor U14938 (N_14938,N_10170,N_9087);
nand U14939 (N_14939,N_9496,N_10812);
and U14940 (N_14940,N_9186,N_9313);
xor U14941 (N_14941,N_11216,N_10050);
nand U14942 (N_14942,N_9444,N_11573);
or U14943 (N_14943,N_11348,N_9701);
xnor U14944 (N_14944,N_10457,N_10934);
nand U14945 (N_14945,N_9931,N_11038);
nand U14946 (N_14946,N_10320,N_11648);
xnor U14947 (N_14947,N_10886,N_9435);
and U14948 (N_14948,N_10637,N_11498);
and U14949 (N_14949,N_11144,N_9376);
nor U14950 (N_14950,N_10418,N_11191);
nor U14951 (N_14951,N_11858,N_11004);
xor U14952 (N_14952,N_9723,N_9053);
or U14953 (N_14953,N_9287,N_10213);
nand U14954 (N_14954,N_11693,N_9448);
and U14955 (N_14955,N_11430,N_9904);
or U14956 (N_14956,N_9972,N_10333);
or U14957 (N_14957,N_11457,N_11166);
xor U14958 (N_14958,N_9291,N_9646);
nor U14959 (N_14959,N_9370,N_9228);
xor U14960 (N_14960,N_11870,N_10761);
xnor U14961 (N_14961,N_9567,N_11368);
or U14962 (N_14962,N_9788,N_10782);
nor U14963 (N_14963,N_11147,N_10360);
nor U14964 (N_14964,N_10111,N_11601);
nand U14965 (N_14965,N_11846,N_9181);
nor U14966 (N_14966,N_11830,N_11904);
and U14967 (N_14967,N_10321,N_10162);
nor U14968 (N_14968,N_11718,N_10938);
xnor U14969 (N_14969,N_11063,N_11300);
nor U14970 (N_14970,N_10787,N_11663);
nand U14971 (N_14971,N_10911,N_11045);
nor U14972 (N_14972,N_9644,N_9974);
xnor U14973 (N_14973,N_9116,N_9681);
nand U14974 (N_14974,N_11642,N_9296);
or U14975 (N_14975,N_11360,N_10658);
nand U14976 (N_14976,N_10898,N_10915);
or U14977 (N_14977,N_9251,N_9313);
xor U14978 (N_14978,N_9434,N_11369);
xor U14979 (N_14979,N_10459,N_10855);
xor U14980 (N_14980,N_9083,N_9115);
or U14981 (N_14981,N_11118,N_10769);
nor U14982 (N_14982,N_9225,N_9421);
or U14983 (N_14983,N_11866,N_10494);
or U14984 (N_14984,N_10963,N_10329);
nand U14985 (N_14985,N_9402,N_11348);
or U14986 (N_14986,N_11950,N_9672);
xor U14987 (N_14987,N_11663,N_11517);
nor U14988 (N_14988,N_9589,N_11618);
nor U14989 (N_14989,N_9587,N_10873);
nor U14990 (N_14990,N_10084,N_10702);
and U14991 (N_14991,N_9784,N_10477);
xnor U14992 (N_14992,N_11629,N_11024);
xnor U14993 (N_14993,N_11356,N_11432);
nand U14994 (N_14994,N_9977,N_10439);
and U14995 (N_14995,N_9973,N_11489);
nor U14996 (N_14996,N_11310,N_10409);
nand U14997 (N_14997,N_10955,N_11367);
xnor U14998 (N_14998,N_11146,N_11451);
xnor U14999 (N_14999,N_9405,N_9561);
xnor U15000 (N_15000,N_12469,N_12592);
xor U15001 (N_15001,N_14676,N_12556);
nor U15002 (N_15002,N_14820,N_14880);
xor U15003 (N_15003,N_14411,N_14690);
or U15004 (N_15004,N_14841,N_13231);
xor U15005 (N_15005,N_13342,N_14060);
and U15006 (N_15006,N_14849,N_12240);
and U15007 (N_15007,N_13379,N_13163);
nor U15008 (N_15008,N_12279,N_14585);
nor U15009 (N_15009,N_13911,N_12905);
and U15010 (N_15010,N_14210,N_13384);
xor U15011 (N_15011,N_13353,N_13781);
xor U15012 (N_15012,N_14409,N_13704);
nor U15013 (N_15013,N_14954,N_12071);
nand U15014 (N_15014,N_12521,N_14757);
or U15015 (N_15015,N_12290,N_12120);
xor U15016 (N_15016,N_14012,N_14176);
nand U15017 (N_15017,N_14451,N_12941);
xnor U15018 (N_15018,N_12891,N_13573);
and U15019 (N_15019,N_13796,N_12808);
and U15020 (N_15020,N_14425,N_12403);
and U15021 (N_15021,N_13184,N_12079);
or U15022 (N_15022,N_12273,N_13482);
nor U15023 (N_15023,N_12777,N_14090);
and U15024 (N_15024,N_14037,N_14550);
or U15025 (N_15025,N_13111,N_12125);
nand U15026 (N_15026,N_13443,N_14271);
nand U15027 (N_15027,N_12118,N_12813);
xnor U15028 (N_15028,N_13851,N_12321);
or U15029 (N_15029,N_14462,N_12585);
and U15030 (N_15030,N_14034,N_14081);
nor U15031 (N_15031,N_12928,N_13800);
nand U15032 (N_15032,N_14931,N_13229);
or U15033 (N_15033,N_13833,N_13901);
nand U15034 (N_15034,N_13164,N_13354);
nor U15035 (N_15035,N_14016,N_12881);
and U15036 (N_15036,N_13021,N_13110);
and U15037 (N_15037,N_13621,N_14123);
xnor U15038 (N_15038,N_13351,N_12685);
nor U15039 (N_15039,N_14388,N_13271);
or U15040 (N_15040,N_14990,N_14414);
or U15041 (N_15041,N_12242,N_13128);
xnor U15042 (N_15042,N_12130,N_14423);
or U15043 (N_15043,N_14069,N_14241);
xnor U15044 (N_15044,N_14493,N_12773);
or U15045 (N_15045,N_13070,N_14167);
nand U15046 (N_15046,N_12363,N_13727);
nand U15047 (N_15047,N_13780,N_14084);
or U15048 (N_15048,N_13948,N_14994);
xnor U15049 (N_15049,N_14989,N_14879);
and U15050 (N_15050,N_12305,N_14041);
and U15051 (N_15051,N_13199,N_14042);
and U15052 (N_15052,N_12088,N_14453);
nor U15053 (N_15053,N_14431,N_13468);
or U15054 (N_15054,N_12869,N_14186);
xor U15055 (N_15055,N_12925,N_12107);
nor U15056 (N_15056,N_14712,N_12593);
nand U15057 (N_15057,N_13042,N_13358);
xor U15058 (N_15058,N_12366,N_12989);
or U15059 (N_15059,N_13740,N_14352);
xor U15060 (N_15060,N_13606,N_13862);
and U15061 (N_15061,N_12570,N_12659);
and U15062 (N_15062,N_13926,N_13333);
and U15063 (N_15063,N_14429,N_12539);
and U15064 (N_15064,N_12186,N_14103);
or U15065 (N_15065,N_14303,N_12298);
or U15066 (N_15066,N_12329,N_13630);
nand U15067 (N_15067,N_14104,N_12051);
xor U15068 (N_15068,N_12829,N_14056);
nor U15069 (N_15069,N_13041,N_13334);
xnor U15070 (N_15070,N_12849,N_13052);
nand U15071 (N_15071,N_13015,N_12189);
nand U15072 (N_15072,N_14524,N_13298);
nor U15073 (N_15073,N_12776,N_12901);
nand U15074 (N_15074,N_12992,N_12575);
nor U15075 (N_15075,N_13832,N_13132);
and U15076 (N_15076,N_13520,N_13966);
nand U15077 (N_15077,N_13531,N_14952);
and U15078 (N_15078,N_13922,N_13994);
nor U15079 (N_15079,N_14937,N_14615);
nor U15080 (N_15080,N_14969,N_12048);
nand U15081 (N_15081,N_13667,N_12175);
nand U15082 (N_15082,N_14513,N_13393);
xor U15083 (N_15083,N_13425,N_13102);
nand U15084 (N_15084,N_12263,N_12655);
nand U15085 (N_15085,N_12357,N_12606);
nand U15086 (N_15086,N_12880,N_14201);
and U15087 (N_15087,N_13762,N_12373);
or U15088 (N_15088,N_12170,N_14775);
xor U15089 (N_15089,N_13161,N_12875);
and U15090 (N_15090,N_12984,N_13859);
nand U15091 (N_15091,N_12047,N_14560);
or U15092 (N_15092,N_14895,N_14175);
nor U15093 (N_15093,N_13527,N_12024);
xor U15094 (N_15094,N_12212,N_13089);
nand U15095 (N_15095,N_12015,N_13261);
nand U15096 (N_15096,N_14733,N_14074);
xnor U15097 (N_15097,N_14465,N_13129);
nor U15098 (N_15098,N_13297,N_12225);
nand U15099 (N_15099,N_13441,N_12818);
nand U15100 (N_15100,N_14227,N_14758);
nand U15101 (N_15101,N_13471,N_13495);
and U15102 (N_15102,N_12464,N_13462);
nand U15103 (N_15103,N_13653,N_14569);
and U15104 (N_15104,N_14883,N_13338);
nand U15105 (N_15105,N_12326,N_12716);
or U15106 (N_15106,N_12266,N_12749);
or U15107 (N_15107,N_13293,N_14025);
xnor U15108 (N_15108,N_13294,N_14778);
or U15109 (N_15109,N_14053,N_14939);
nor U15110 (N_15110,N_13241,N_14221);
nor U15111 (N_15111,N_14089,N_12924);
nand U15112 (N_15112,N_12293,N_12319);
xnor U15113 (N_15113,N_13005,N_14334);
and U15114 (N_15114,N_13248,N_13602);
or U15115 (N_15115,N_12261,N_14728);
nor U15116 (N_15116,N_13319,N_13550);
xnor U15117 (N_15117,N_14756,N_12392);
xnor U15118 (N_15118,N_14310,N_14947);
and U15119 (N_15119,N_14397,N_13802);
and U15120 (N_15120,N_14270,N_14920);
nor U15121 (N_15121,N_14450,N_13494);
or U15122 (N_15122,N_14643,N_13839);
and U15123 (N_15123,N_13515,N_12661);
or U15124 (N_15124,N_14396,N_13399);
and U15125 (N_15125,N_12280,N_14054);
nor U15126 (N_15126,N_12632,N_13541);
nor U15127 (N_15127,N_13153,N_12448);
xor U15128 (N_15128,N_13291,N_12017);
xnor U15129 (N_15129,N_13883,N_12304);
nand U15130 (N_15130,N_13478,N_13688);
and U15131 (N_15131,N_12315,N_13265);
or U15132 (N_15132,N_14108,N_14032);
or U15133 (N_15133,N_12437,N_13917);
or U15134 (N_15134,N_14911,N_14761);
nor U15135 (N_15135,N_14696,N_12620);
or U15136 (N_15136,N_13871,N_14184);
and U15137 (N_15137,N_12757,N_13296);
and U15138 (N_15138,N_14634,N_12059);
xor U15139 (N_15139,N_13924,N_14861);
xor U15140 (N_15140,N_13061,N_12731);
nor U15141 (N_15141,N_12191,N_14516);
nor U15142 (N_15142,N_12098,N_14407);
and U15143 (N_15143,N_14022,N_14116);
and U15144 (N_15144,N_12911,N_14073);
xnor U15145 (N_15145,N_14460,N_12312);
nand U15146 (N_15146,N_13992,N_12255);
or U15147 (N_15147,N_12486,N_14926);
and U15148 (N_15148,N_12528,N_12381);
xor U15149 (N_15149,N_12221,N_14348);
or U15150 (N_15150,N_13475,N_14638);
nand U15151 (N_15151,N_13073,N_12308);
nor U15152 (N_15152,N_14114,N_13240);
nand U15153 (N_15153,N_12549,N_12504);
xor U15154 (N_15154,N_12588,N_13730);
xnor U15155 (N_15155,N_14412,N_14654);
and U15156 (N_15156,N_14913,N_12826);
or U15157 (N_15157,N_14943,N_12270);
nor U15158 (N_15158,N_12489,N_14050);
nand U15159 (N_15159,N_13956,N_13100);
and U15160 (N_15160,N_13996,N_13618);
or U15161 (N_15161,N_12996,N_13173);
nor U15162 (N_15162,N_13880,N_14632);
and U15163 (N_15163,N_12733,N_13689);
nand U15164 (N_15164,N_12820,N_13914);
nand U15165 (N_15165,N_14824,N_14802);
nand U15166 (N_15166,N_13349,N_13577);
and U15167 (N_15167,N_14660,N_12190);
or U15168 (N_15168,N_12384,N_14614);
nand U15169 (N_15169,N_14823,N_13801);
or U15170 (N_15170,N_12760,N_13193);
xnor U15171 (N_15171,N_14498,N_14147);
nor U15172 (N_15172,N_13784,N_13836);
or U15173 (N_15173,N_14933,N_13558);
xnor U15174 (N_15174,N_13510,N_13838);
nor U15175 (N_15175,N_12827,N_12081);
nor U15176 (N_15176,N_12722,N_12472);
xnor U15177 (N_15177,N_12837,N_13029);
or U15178 (N_15178,N_14700,N_12424);
and U15179 (N_15179,N_12004,N_13025);
nand U15180 (N_15180,N_14278,N_12307);
nand U15181 (N_15181,N_13869,N_13691);
nand U15182 (N_15182,N_14902,N_12960);
nor U15183 (N_15183,N_12287,N_14653);
or U15184 (N_15184,N_14096,N_13043);
nand U15185 (N_15185,N_12557,N_14991);
or U15186 (N_15186,N_13305,N_14571);
nor U15187 (N_15187,N_12336,N_12184);
nand U15188 (N_15188,N_14827,N_13844);
and U15189 (N_15189,N_14805,N_12822);
xnor U15190 (N_15190,N_14449,N_14680);
or U15191 (N_15191,N_14027,N_13736);
xor U15192 (N_15192,N_13818,N_13097);
xor U15193 (N_15193,N_13207,N_14871);
or U15194 (N_15194,N_12920,N_14415);
nor U15195 (N_15195,N_14283,N_12997);
nor U15196 (N_15196,N_12897,N_12168);
nor U15197 (N_15197,N_12903,N_14767);
or U15198 (N_15198,N_13642,N_14098);
nor U15199 (N_15199,N_13747,N_13710);
xor U15200 (N_15200,N_14521,N_12511);
xor U15201 (N_15201,N_12387,N_12738);
nor U15202 (N_15202,N_12207,N_12018);
xor U15203 (N_15203,N_14727,N_12815);
and U15204 (N_15204,N_14275,N_14608);
nor U15205 (N_15205,N_12149,N_12096);
nand U15206 (N_15206,N_12094,N_12551);
nor U15207 (N_15207,N_12823,N_12188);
or U15208 (N_15208,N_13392,N_14936);
xnor U15209 (N_15209,N_13212,N_13071);
xnor U15210 (N_15210,N_12629,N_13596);
or U15211 (N_15211,N_13079,N_12852);
nor U15212 (N_15212,N_13063,N_13921);
and U15213 (N_15213,N_13687,N_13247);
or U15214 (N_15214,N_12938,N_14635);
xor U15215 (N_15215,N_13017,N_13939);
nor U15216 (N_15216,N_13067,N_13320);
nor U15217 (N_15217,N_12419,N_12176);
and U15218 (N_15218,N_12954,N_14265);
xor U15219 (N_15219,N_14488,N_12861);
nand U15220 (N_15220,N_12534,N_12223);
nor U15221 (N_15221,N_12995,N_12604);
nor U15222 (N_15222,N_12112,N_12093);
nor U15223 (N_15223,N_12998,N_14086);
nand U15224 (N_15224,N_14329,N_13881);
nand U15225 (N_15225,N_13717,N_14385);
nor U15226 (N_15226,N_14229,N_14904);
nand U15227 (N_15227,N_13623,N_13563);
nor U15228 (N_15228,N_14185,N_14381);
xor U15229 (N_15229,N_13278,N_13284);
nor U15230 (N_15230,N_14255,N_14049);
xor U15231 (N_15231,N_14940,N_12099);
nand U15232 (N_15232,N_13729,N_12691);
nor U15233 (N_15233,N_12517,N_13485);
nand U15234 (N_15234,N_14187,N_13543);
nand U15235 (N_15235,N_14137,N_14238);
nor U15236 (N_15236,N_14522,N_12396);
or U15237 (N_15237,N_12509,N_13607);
nand U15238 (N_15238,N_12062,N_14673);
nor U15239 (N_15239,N_13064,N_12976);
nor U15240 (N_15240,N_13407,N_13656);
or U15241 (N_15241,N_13215,N_13086);
or U15242 (N_15242,N_13401,N_13321);
nor U15243 (N_15243,N_13908,N_14699);
or U15244 (N_15244,N_14979,N_14629);
nor U15245 (N_15245,N_12353,N_14068);
nor U15246 (N_15246,N_13146,N_13739);
nand U15247 (N_15247,N_14268,N_13394);
and U15248 (N_15248,N_12092,N_13898);
or U15249 (N_15249,N_12939,N_13503);
and U15250 (N_15250,N_14036,N_12423);
xor U15251 (N_15251,N_12598,N_13260);
nor U15252 (N_15252,N_12919,N_14956);
nand U15253 (N_15253,N_13157,N_12166);
nor U15254 (N_15254,N_13388,N_12249);
or U15255 (N_15255,N_12725,N_14655);
xnor U15256 (N_15256,N_13581,N_14142);
or U15257 (N_15257,N_12145,N_14769);
xnor U15258 (N_15258,N_13303,N_14173);
and U15259 (N_15259,N_12003,N_13032);
nor U15260 (N_15260,N_13929,N_13882);
xnor U15261 (N_15261,N_14203,N_13222);
and U15262 (N_15262,N_12378,N_12036);
xor U15263 (N_15263,N_12153,N_12838);
nand U15264 (N_15264,N_13951,N_14717);
nor U15265 (N_15265,N_13977,N_13777);
xnor U15266 (N_15266,N_12752,N_12426);
and U15267 (N_15267,N_13117,N_13179);
nor U15268 (N_15268,N_14720,N_13564);
xor U15269 (N_15269,N_13744,N_13533);
nand U15270 (N_15270,N_12370,N_13398);
nand U15271 (N_15271,N_14289,N_14531);
xnor U15272 (N_15272,N_13972,N_13373);
or U15273 (N_15273,N_14239,N_14064);
xnor U15274 (N_15274,N_14514,N_13118);
nor U15275 (N_15275,N_12172,N_14921);
nand U15276 (N_15276,N_13714,N_13845);
nand U15277 (N_15277,N_13909,N_12612);
nand U15278 (N_15278,N_14970,N_12558);
and U15279 (N_15279,N_12006,N_13509);
and U15280 (N_15280,N_12127,N_13336);
and U15281 (N_15281,N_12768,N_12202);
xor U15282 (N_15282,N_14293,N_14287);
nand U15283 (N_15283,N_13142,N_13657);
nor U15284 (N_15284,N_12203,N_13022);
or U15285 (N_15285,N_14924,N_13020);
nor U15286 (N_15286,N_12070,N_13715);
or U15287 (N_15287,N_14434,N_14166);
nor U15288 (N_15288,N_14770,N_12871);
nand U15289 (N_15289,N_14882,N_13574);
nand U15290 (N_15290,N_14836,N_12335);
and U15291 (N_15291,N_12433,N_14714);
or U15292 (N_15292,N_14974,N_14961);
xnor U15293 (N_15293,N_12354,N_12721);
and U15294 (N_15294,N_13371,N_14118);
or U15295 (N_15295,N_14009,N_13890);
nor U15296 (N_15296,N_12301,N_14332);
or U15297 (N_15297,N_14566,N_14981);
nand U15298 (N_15298,N_14214,N_12497);
nand U15299 (N_15299,N_13937,N_13290);
nor U15300 (N_15300,N_12247,N_14015);
and U15301 (N_15301,N_13819,N_14688);
nand U15302 (N_15302,N_12325,N_12117);
nor U15303 (N_15303,N_13962,N_14602);
xnor U15304 (N_15304,N_12602,N_12498);
or U15305 (N_15305,N_13650,N_13292);
xnor U15306 (N_15306,N_12578,N_13915);
or U15307 (N_15307,N_13137,N_14294);
xnor U15308 (N_15308,N_13706,N_14914);
and U15309 (N_15309,N_13344,N_12964);
nor U15310 (N_15310,N_13723,N_14484);
or U15311 (N_15311,N_14162,N_12200);
or U15312 (N_15312,N_12552,N_14427);
xnor U15313 (N_15313,N_12689,N_12488);
nand U15314 (N_15314,N_13410,N_14178);
or U15315 (N_15315,N_14206,N_14734);
xor U15316 (N_15316,N_13442,N_13788);
nor U15317 (N_15317,N_14151,N_14896);
nand U15318 (N_15318,N_14744,N_12567);
nand U15319 (N_15319,N_14748,N_14826);
or U15320 (N_15320,N_12148,N_13332);
nand U15321 (N_15321,N_14577,N_12978);
or U15322 (N_15322,N_14010,N_14563);
and U15323 (N_15323,N_14280,N_14356);
or U15324 (N_15324,N_12443,N_14259);
xnor U15325 (N_15325,N_12324,N_12688);
or U15326 (N_15326,N_12044,N_14842);
xnor U15327 (N_15327,N_12991,N_13178);
and U15328 (N_15328,N_13255,N_14469);
nand U15329 (N_15329,N_14612,N_12968);
nand U15330 (N_15330,N_13428,N_14636);
or U15331 (N_15331,N_13634,N_14244);
nand U15332 (N_15332,N_12475,N_13287);
and U15333 (N_15333,N_14859,N_13473);
nand U15334 (N_15334,N_14260,N_14648);
xnor U15335 (N_15335,N_12455,N_12365);
xnor U15336 (N_15336,N_12643,N_13006);
nor U15337 (N_15337,N_12058,N_14305);
xor U15338 (N_15338,N_14856,N_12398);
nand U15339 (N_15339,N_12320,N_13799);
and U15340 (N_15340,N_12653,N_13369);
nand U15341 (N_15341,N_14026,N_13920);
and U15342 (N_15342,N_14209,N_13814);
nor U15343 (N_15343,N_14708,N_12333);
nor U15344 (N_15344,N_14134,N_12719);
and U15345 (N_15345,N_13805,N_13539);
nand U15346 (N_15346,N_12197,N_13872);
xnor U15347 (N_15347,N_13242,N_13504);
nand U15348 (N_15348,N_13195,N_13430);
nand U15349 (N_15349,N_13434,N_12732);
nand U15350 (N_15350,N_14799,N_12297);
xnor U15351 (N_15351,N_13340,N_12883);
and U15352 (N_15352,N_13050,N_12582);
nand U15353 (N_15353,N_13794,N_13775);
xor U15354 (N_15354,N_13049,N_14078);
or U15355 (N_15355,N_13044,N_13980);
xor U15356 (N_15356,N_12817,N_13448);
or U15357 (N_15357,N_12702,N_13923);
and U15358 (N_15358,N_14567,N_13346);
nand U15359 (N_15359,N_12783,N_14962);
nor U15360 (N_15360,N_14852,N_14177);
nand U15361 (N_15361,N_13521,N_12364);
or U15362 (N_15362,N_14606,N_12930);
nand U15363 (N_15363,N_12114,N_14527);
and U15364 (N_15364,N_12239,N_13266);
nand U15365 (N_15365,N_12876,N_12779);
and U15366 (N_15366,N_13182,N_12569);
xnor U15367 (N_15367,N_13582,N_12229);
nand U15368 (N_15368,N_13580,N_13586);
nand U15369 (N_15369,N_12866,N_12041);
xor U15370 (N_15370,N_14377,N_14963);
nor U15371 (N_15371,N_13451,N_13474);
xor U15372 (N_15372,N_12709,N_14800);
nand U15373 (N_15373,N_13892,N_12670);
and U15374 (N_15374,N_13605,N_12123);
nand U15375 (N_15375,N_14532,N_13548);
nor U15376 (N_15376,N_12935,N_12595);
nor U15377 (N_15377,N_12181,N_14843);
nor U15378 (N_15378,N_14507,N_12420);
and U15379 (N_15379,N_12609,N_14325);
nor U15380 (N_15380,N_14006,N_14383);
or U15381 (N_15381,N_12260,N_13652);
xnor U15382 (N_15382,N_14452,N_12970);
nor U15383 (N_15383,N_12596,N_14245);
or U15384 (N_15384,N_13726,N_14277);
and U15385 (N_15385,N_13221,N_13300);
nor U15386 (N_15386,N_12660,N_14941);
nor U15387 (N_15387,N_12135,N_13684);
and U15388 (N_15388,N_14821,N_12167);
nor U15389 (N_15389,N_13860,N_13792);
nor U15390 (N_15390,N_13854,N_14951);
or U15391 (N_15391,N_14038,N_13660);
nand U15392 (N_15392,N_13771,N_13716);
nor U15393 (N_15393,N_13405,N_14393);
and U15394 (N_15394,N_14299,N_12262);
nand U15395 (N_15395,N_14059,N_14152);
nand U15396 (N_15396,N_14763,N_14341);
nand U15397 (N_15397,N_14487,N_14490);
or U15398 (N_15398,N_13617,N_14247);
and U15399 (N_15399,N_13786,N_14335);
xor U15400 (N_15400,N_14447,N_12216);
xnor U15401 (N_15401,N_14467,N_13542);
nor U15402 (N_15402,N_14645,N_12814);
nand U15403 (N_15403,N_14626,N_13846);
nand U15404 (N_15404,N_12737,N_12990);
xor U15405 (N_15405,N_13680,N_13331);
and U15406 (N_15406,N_13134,N_14605);
or U15407 (N_15407,N_12183,N_14682);
nor U15408 (N_15408,N_12182,N_12224);
or U15409 (N_15409,N_14338,N_14538);
nor U15410 (N_15410,N_14117,N_12295);
nor U15411 (N_15411,N_13252,N_13516);
or U15412 (N_15412,N_14344,N_14495);
nand U15413 (N_15413,N_12724,N_13325);
or U15414 (N_15414,N_14120,N_14342);
or U15415 (N_15415,N_13156,N_12980);
or U15416 (N_15416,N_13375,N_13066);
and U15417 (N_15417,N_14121,N_14753);
nor U15418 (N_15418,N_13057,N_14650);
or U15419 (N_15419,N_12401,N_12973);
or U15420 (N_15420,N_12965,N_14623);
nor U15421 (N_15421,N_12360,N_12434);
and U15422 (N_15422,N_14985,N_12402);
nor U15423 (N_15423,N_13651,N_12812);
nor U15424 (N_15424,N_13518,N_12801);
or U15425 (N_15425,N_14130,N_13497);
nand U15426 (N_15426,N_14755,N_12016);
xnor U15427 (N_15427,N_13416,N_14683);
and U15428 (N_15428,N_13763,N_12102);
nor U15429 (N_15429,N_14321,N_12522);
or U15430 (N_15430,N_13946,N_13733);
nor U15431 (N_15431,N_13938,N_14047);
nor U15432 (N_15432,N_12043,N_14458);
nand U15433 (N_15433,N_14301,N_12083);
nand U15434 (N_15434,N_13328,N_12507);
nor U15435 (N_15435,N_13357,N_12975);
nand U15436 (N_15436,N_12617,N_14466);
or U15437 (N_15437,N_13175,N_12037);
nor U15438 (N_15438,N_14212,N_12429);
nand U15439 (N_15439,N_12180,N_14122);
nor U15440 (N_15440,N_12907,N_13483);
or U15441 (N_15441,N_12514,N_14424);
nor U15442 (N_15442,N_14071,N_14033);
or U15443 (N_15443,N_12178,N_14472);
xnor U15444 (N_15444,N_12103,N_13314);
nor U15445 (N_15445,N_13830,N_13812);
nand U15446 (N_15446,N_12303,N_12759);
nor U15447 (N_15447,N_13529,N_14530);
xor U15448 (N_15448,N_12065,N_14723);
nor U15449 (N_15449,N_12872,N_13389);
nor U15450 (N_15450,N_14099,N_12476);
or U15451 (N_15451,N_14661,N_13815);
nand U15452 (N_15452,N_14331,N_14535);
or U15453 (N_15453,N_13850,N_13464);
nor U15454 (N_15454,N_12850,N_12805);
nor U15455 (N_15455,N_12131,N_12674);
or U15456 (N_15456,N_13906,N_13644);
xor U15457 (N_15457,N_13214,N_12825);
and U15458 (N_15458,N_14886,N_12900);
nor U15459 (N_15459,N_14950,N_14274);
nor U15460 (N_15460,N_14812,N_14292);
nor U15461 (N_15461,N_14809,N_13010);
or U15462 (N_15462,N_13234,N_14958);
xnor U15463 (N_15463,N_12339,N_14480);
or U15464 (N_15464,N_14853,N_13514);
and U15465 (N_15465,N_12481,N_13659);
or U15466 (N_15466,N_14219,N_13633);
xnor U15467 (N_15467,N_13545,N_14630);
nand U15468 (N_15468,N_13589,N_13082);
nand U15469 (N_15469,N_13481,N_13289);
nor U15470 (N_15470,N_14998,N_14156);
or U15471 (N_15471,N_13707,N_14833);
or U15472 (N_15472,N_14249,N_13899);
xor U15473 (N_15473,N_12028,N_12832);
xnor U15474 (N_15474,N_14432,N_14387);
nand U15475 (N_15475,N_12914,N_14316);
and U15476 (N_15476,N_14868,N_14603);
or U15477 (N_15477,N_13991,N_13455);
nor U15478 (N_15478,N_13286,N_12014);
nor U15479 (N_15479,N_14980,N_13382);
and U15480 (N_15480,N_14044,N_13059);
nand U15481 (N_15481,N_14438,N_13821);
or U15482 (N_15482,N_14506,N_14581);
nor U15483 (N_15483,N_14909,N_14562);
or U15484 (N_15484,N_13218,N_12132);
nor U15485 (N_15485,N_12068,N_14529);
or U15486 (N_15486,N_13643,N_12138);
nand U15487 (N_15487,N_12256,N_14782);
nand U15488 (N_15488,N_12050,N_14004);
or U15489 (N_15489,N_13348,N_12179);
nand U15490 (N_15490,N_12344,N_13795);
nor U15491 (N_15491,N_14906,N_13459);
and U15492 (N_15492,N_13722,N_14373);
nor U15493 (N_15493,N_14464,N_13963);
nor U15494 (N_15494,N_12807,N_14866);
and U15495 (N_15495,N_13989,N_12950);
xnor U15496 (N_15496,N_13578,N_13768);
nand U15497 (N_15497,N_12603,N_12579);
xor U15498 (N_15498,N_14618,N_13597);
nor U15499 (N_15499,N_13014,N_14158);
xnor U15500 (N_15500,N_12794,N_13562);
or U15501 (N_15501,N_14216,N_13620);
xnor U15502 (N_15502,N_12023,N_12728);
nor U15503 (N_15503,N_14399,N_14435);
nand U15504 (N_15504,N_13381,N_14253);
or U15505 (N_15505,N_14202,N_12663);
nand U15506 (N_15506,N_12893,N_12870);
and U15507 (N_15507,N_12146,N_14097);
nor U15508 (N_15508,N_14746,N_14364);
xnor U15509 (N_15509,N_12390,N_13330);
nor U15510 (N_15510,N_14391,N_13840);
xnor U15511 (N_15511,N_12929,N_12128);
or U15512 (N_15512,N_12244,N_13018);
or U15513 (N_15513,N_14595,N_12590);
nor U15514 (N_15514,N_13524,N_14317);
nand U15515 (N_15515,N_13506,N_12809);
nand U15516 (N_15516,N_13378,N_12034);
nand U15517 (N_15517,N_13932,N_12341);
xor U15518 (N_15518,N_12463,N_13551);
or U15519 (N_15519,N_13372,N_12775);
xor U15520 (N_15520,N_14599,N_14668);
nand U15521 (N_15521,N_14324,N_12126);
or U15522 (N_15522,N_13879,N_12008);
nor U15523 (N_15523,N_12896,N_12222);
nor U15524 (N_15524,N_13060,N_14865);
nand U15525 (N_15525,N_13600,N_13933);
nor U15526 (N_15526,N_13213,N_12432);
nand U15527 (N_15527,N_13793,N_13109);
xnor U15528 (N_15528,N_14314,N_13191);
xnor U15529 (N_15529,N_12459,N_14095);
xor U15530 (N_15530,N_12703,N_13194);
nor U15531 (N_15531,N_13499,N_12736);
or U15532 (N_15532,N_13817,N_13546);
and U15533 (N_15533,N_12999,N_12494);
nor U15534 (N_15534,N_14327,N_14213);
nor U15535 (N_15535,N_13352,N_13200);
and U15536 (N_15536,N_12252,N_12198);
nand U15537 (N_15537,N_13444,N_13120);
nand U15538 (N_15538,N_13902,N_14248);
nor U15539 (N_15539,N_14298,N_12994);
nor U15540 (N_15540,N_12981,N_12505);
or U15541 (N_15541,N_14918,N_14922);
or U15542 (N_15542,N_13188,N_12013);
nor U15543 (N_15543,N_13955,N_14172);
and U15544 (N_15544,N_13635,N_13149);
nor U15545 (N_15545,N_14061,N_13208);
xnor U15546 (N_15546,N_14035,N_14446);
xor U15547 (N_15547,N_12797,N_13610);
nand U15548 (N_15548,N_13148,N_13806);
xnor U15549 (N_15549,N_14076,N_14613);
or U15550 (N_15550,N_13493,N_12506);
or U15551 (N_15551,N_13317,N_13268);
and U15552 (N_15552,N_13811,N_13971);
xnor U15553 (N_15553,N_12956,N_12698);
xor U15554 (N_15554,N_14444,N_12458);
nand U15555 (N_15555,N_12931,N_12410);
or U15556 (N_15556,N_12194,N_14976);
and U15557 (N_15557,N_14242,N_12348);
xor U15558 (N_15558,N_13339,N_12072);
and U15559 (N_15559,N_13983,N_13984);
and U15560 (N_15560,N_13072,N_13944);
and U15561 (N_15561,N_13682,N_14360);
or U15562 (N_15562,N_14942,N_12144);
and U15563 (N_15563,N_13907,N_14021);
xor U15564 (N_15564,N_12792,N_12535);
xor U15565 (N_15565,N_13568,N_12097);
xor U15566 (N_15566,N_13960,N_14830);
nor U15567 (N_15567,N_13614,N_13904);
or U15568 (N_15568,N_12676,N_12701);
nand U15569 (N_15569,N_12063,N_14126);
or U15570 (N_15570,N_14029,N_13671);
nand U15571 (N_15571,N_13700,N_13105);
nand U15572 (N_15572,N_12678,N_12967);
xnor U15573 (N_15573,N_14528,N_12854);
xnor U15574 (N_15574,N_14777,N_14817);
nor U15575 (N_15575,N_14787,N_14232);
nor U15576 (N_15576,N_12226,N_13807);
xor U15577 (N_15577,N_13169,N_12734);
nand U15578 (N_15578,N_12525,N_12033);
or U15579 (N_15579,N_14199,N_13439);
nor U15580 (N_15580,N_14504,N_13608);
xor U15581 (N_15581,N_13738,N_14557);
nor U15582 (N_15582,N_12786,N_14011);
nand U15583 (N_15583,N_12031,N_13662);
nand U15584 (N_15584,N_12251,N_12345);
or U15585 (N_15585,N_14776,N_13387);
nand U15586 (N_15586,N_12680,N_12199);
nand U15587 (N_15587,N_14982,N_14666);
nand U15588 (N_15588,N_13828,N_13857);
nor U15589 (N_15589,N_13259,N_14211);
and U15590 (N_15590,N_14105,N_14109);
and U15591 (N_15591,N_12292,N_12542);
xor U15592 (N_15592,N_14246,N_13613);
xor U15593 (N_15593,N_14647,N_14138);
nor U15594 (N_15594,N_14588,N_14276);
nor U15595 (N_15595,N_14808,N_13302);
or U15596 (N_15596,N_14518,N_14740);
nand U15597 (N_15597,N_13162,N_13876);
and U15598 (N_15598,N_13365,N_13437);
nor U15599 (N_15599,N_13335,N_13456);
xor U15600 (N_15600,N_14129,N_13639);
or U15601 (N_15601,N_13609,N_12462);
nand U15602 (N_15602,N_13279,N_12564);
and U15603 (N_15603,N_12969,N_12165);
nand U15604 (N_15604,N_12057,N_12508);
and U15605 (N_15605,N_13856,N_12751);
and U15606 (N_15606,N_13502,N_13954);
and U15607 (N_15607,N_13092,N_12436);
and U15608 (N_15608,N_12115,N_13570);
xnor U15609 (N_15609,N_12468,N_14290);
or U15610 (N_15610,N_12641,N_12649);
nor U15611 (N_15611,N_12000,N_12784);
and U15612 (N_15612,N_12215,N_13627);
and U15613 (N_15613,N_14363,N_13827);
and U15614 (N_15614,N_12946,N_13101);
or U15615 (N_15615,N_13649,N_12347);
xor U15616 (N_15616,N_14701,N_12597);
and U15617 (N_15617,N_13058,N_12143);
and U15618 (N_15618,N_14890,N_14470);
nand U15619 (N_15619,N_12841,N_13673);
nand U15620 (N_15620,N_12232,N_14023);
nand U15621 (N_15621,N_14386,N_12192);
xnor U15622 (N_15622,N_12758,N_14226);
nor U15623 (N_15623,N_13804,N_13364);
nor U15624 (N_15624,N_14544,N_12136);
or U15625 (N_15625,N_13486,N_13891);
or U15626 (N_15626,N_12485,N_14311);
nand U15627 (N_15627,N_12627,N_12399);
xor U15628 (N_15628,N_14308,N_13224);
and U15629 (N_15629,N_13874,N_12095);
and U15630 (N_15630,N_13237,N_12141);
or U15631 (N_15631,N_13243,N_13076);
nand U15632 (N_15632,N_14794,N_13949);
xnor U15633 (N_15633,N_13492,N_12972);
or U15634 (N_15634,N_14168,N_13591);
nor U15635 (N_15635,N_12452,N_14917);
xnor U15636 (N_15636,N_14371,N_12235);
xor U15637 (N_15637,N_13576,N_13601);
and U15638 (N_15638,N_12408,N_12963);
or U15639 (N_15639,N_12471,N_13239);
and U15640 (N_15640,N_12780,N_12159);
and U15641 (N_15641,N_14536,N_13085);
xnor U15642 (N_15642,N_12447,N_14785);
or U15643 (N_15643,N_13028,N_14441);
and U15644 (N_15644,N_14675,N_12619);
and U15645 (N_15645,N_12400,N_14159);
or U15646 (N_15646,N_13698,N_13068);
nor U15647 (N_15647,N_14315,N_13735);
nor U15648 (N_15648,N_14288,N_12879);
nor U15649 (N_15649,N_14190,N_13625);
or U15650 (N_15650,N_14693,N_14113);
or U15651 (N_15651,N_14367,N_14234);
and U15652 (N_15652,N_12543,N_14771);
nor U15653 (N_15653,N_12090,N_13177);
nor U15654 (N_15654,N_14899,N_12106);
xor U15655 (N_15655,N_13469,N_14900);
nor U15656 (N_15656,N_14834,N_14741);
xor U15657 (N_15657,N_12358,N_13374);
xnor U15658 (N_15658,N_12637,N_14553);
xnor U15659 (N_15659,N_13282,N_12346);
nor U15660 (N_15660,N_14473,N_14732);
or U15661 (N_15661,N_13803,N_12743);
xnor U15662 (N_15662,N_14534,N_12484);
nand U15663 (N_15663,N_14160,N_14164);
nand U15664 (N_15664,N_14706,N_14401);
nor U15665 (N_15665,N_14687,N_13995);
nor U15666 (N_15666,N_12022,N_14598);
nor U15667 (N_15667,N_14389,N_12208);
nand U15668 (N_15668,N_14996,N_14910);
nor U15669 (N_15669,N_13843,N_14583);
or U15670 (N_15670,N_12040,N_12431);
nor U15671 (N_15671,N_14392,N_14124);
and U15672 (N_15672,N_14555,N_14191);
nor U15673 (N_15673,N_12726,N_13791);
nand U15674 (N_15674,N_14551,N_14003);
and U15675 (N_15675,N_12671,N_14838);
xor U15676 (N_15676,N_13104,N_14867);
nand U15677 (N_15677,N_12654,N_12035);
nand U15678 (N_15678,N_12799,N_13611);
and U15679 (N_15679,N_13587,N_13183);
and U15680 (N_15680,N_12651,N_12966);
nor U15681 (N_15681,N_12005,N_13201);
or U15682 (N_15682,N_13413,N_14561);
or U15683 (N_15683,N_12533,N_12406);
nand U15684 (N_15684,N_14254,N_12158);
or U15685 (N_15685,N_14616,N_12441);
xnor U15686 (N_15686,N_13720,N_12334);
and U15687 (N_15687,N_13196,N_13604);
and U15688 (N_15688,N_12248,N_12479);
xor U15689 (N_15689,N_12456,N_13790);
nor U15690 (N_15690,N_13235,N_14031);
or U15691 (N_15691,N_12611,N_14368);
xor U15692 (N_15692,N_13942,N_12108);
and U15693 (N_15693,N_12393,N_12926);
or U15694 (N_15694,N_12742,N_14045);
xnor U15695 (N_15695,N_14455,N_14702);
and U15696 (N_15696,N_12411,N_13145);
and U15697 (N_15697,N_13062,N_12754);
and U15698 (N_15698,N_14256,N_12451);
or U15699 (N_15699,N_14983,N_13476);
or U15700 (N_15700,N_13007,N_13685);
nor U15701 (N_15701,N_13080,N_13553);
nor U15702 (N_15702,N_14180,N_14765);
xnor U15703 (N_15703,N_13366,N_12902);
nor U15704 (N_15704,N_14862,N_12407);
and U15705 (N_15705,N_13701,N_12583);
xor U15706 (N_15706,N_12195,N_14801);
nor U15707 (N_15707,N_13590,N_14218);
xor U15708 (N_15708,N_12686,N_14851);
or U15709 (N_15709,N_14062,N_12842);
nor U15710 (N_15710,N_13523,N_13878);
xnor U15711 (N_15711,N_12412,N_13048);
nand U15712 (N_15712,N_14428,N_13310);
or U15713 (N_15713,N_13276,N_14876);
or U15714 (N_15714,N_13254,N_13979);
or U15715 (N_15715,N_12238,N_13534);
nand U15716 (N_15716,N_13910,N_12409);
and U15717 (N_15717,N_12388,N_13705);
nand U15718 (N_15718,N_13345,N_12302);
and U15719 (N_15719,N_14163,N_12473);
xnor U15720 (N_15720,N_14789,N_12706);
and U15721 (N_15721,N_13174,N_13295);
and U15722 (N_15722,N_14145,N_14609);
or U15723 (N_15723,N_12770,N_13816);
or U15724 (N_15724,N_14365,N_12527);
nor U15725 (N_15725,N_12089,N_13250);
nor U15726 (N_15726,N_13767,N_14584);
nand U15727 (N_15727,N_12753,N_12888);
nor U15728 (N_15728,N_14540,N_12756);
xor U15729 (N_15729,N_14426,N_12499);
or U15730 (N_15730,N_14832,N_14328);
nor U15731 (N_15731,N_14711,N_14681);
and U15732 (N_15732,N_12264,N_13186);
nand U15733 (N_15733,N_13488,N_12129);
xor U15734 (N_15734,N_14610,N_14217);
or U15735 (N_15735,N_13829,N_13665);
nor U15736 (N_15736,N_12580,N_13769);
xnor U15737 (N_15737,N_12121,N_14510);
nor U15738 (N_15738,N_12943,N_13719);
xor U15739 (N_15739,N_13166,N_13031);
and U15740 (N_15740,N_13536,N_13941);
nand U15741 (N_15741,N_12945,N_13094);
nor U15742 (N_15742,N_13069,N_12512);
xnor U15743 (N_15743,N_14872,N_14948);
nor U15744 (N_15744,N_13640,N_12778);
nor U15745 (N_15745,N_13056,N_14482);
nor U15746 (N_15746,N_12524,N_14067);
and U15747 (N_15747,N_13170,N_13216);
xnor U15748 (N_15748,N_14949,N_12648);
and U15749 (N_15749,N_12531,N_14320);
xnor U15750 (N_15750,N_14975,N_12091);
xnor U15751 (N_15751,N_14878,N_14671);
nand U15752 (N_15752,N_12633,N_12550);
nor U15753 (N_15753,N_12739,N_14815);
xor U15754 (N_15754,N_12246,N_12591);
nand U15755 (N_15755,N_14875,N_13429);
and U15756 (N_15756,N_13842,N_13547);
nand U15757 (N_15757,N_14930,N_13115);
xor U15758 (N_15758,N_14541,N_14684);
xor U15759 (N_15759,N_13419,N_13197);
xor U15760 (N_15760,N_13970,N_14471);
nor U15761 (N_15761,N_14726,N_14844);
nand U15762 (N_15762,N_14101,N_13151);
and U15763 (N_15763,N_12001,N_13893);
xnor U15764 (N_15764,N_12311,N_14542);
or U15765 (N_15765,N_14092,N_14459);
nor U15766 (N_15766,N_13112,N_14905);
or U15767 (N_15767,N_14578,N_12667);
nand U15768 (N_15768,N_12936,N_12705);
nor U15769 (N_15769,N_12142,N_14492);
or U15770 (N_15770,N_13415,N_12478);
and U15771 (N_15771,N_14257,N_13327);
nand U15772 (N_15772,N_14075,N_14443);
nand U15773 (N_15773,N_12214,N_14088);
and U15774 (N_15774,N_13124,N_14169);
and U15775 (N_15775,N_14421,N_14715);
xor U15776 (N_15776,N_13619,N_14552);
or U15777 (N_15777,N_14828,N_14468);
nand U15778 (N_15778,N_13123,N_12510);
and U15779 (N_15779,N_12196,N_12343);
xor U15780 (N_15780,N_12831,N_12833);
and U15781 (N_15781,N_12934,N_12555);
or U15782 (N_15782,N_14208,N_12821);
or U15783 (N_15783,N_14766,N_12565);
xor U15784 (N_15784,N_14272,N_14988);
and U15785 (N_15785,N_14002,N_12030);
xnor U15786 (N_15786,N_14330,N_14573);
xnor U15787 (N_15787,N_14887,N_12119);
or U15788 (N_15788,N_13631,N_13884);
nand U15789 (N_15789,N_14445,N_12615);
nor U15790 (N_15790,N_13304,N_13233);
and U15791 (N_15791,N_12064,N_13993);
nand U15792 (N_15792,N_12927,N_14873);
xor U15793 (N_15793,N_13787,N_12669);
nor U15794 (N_15794,N_13226,N_14179);
or U15795 (N_15795,N_12523,N_14582);
nor U15796 (N_15796,N_12630,N_14651);
or U15797 (N_15797,N_14346,N_13695);
nor U15798 (N_15798,N_12211,N_12460);
or U15799 (N_15799,N_13283,N_13081);
xnor U15800 (N_15800,N_14822,N_13426);
xnor U15801 (N_15801,N_12982,N_14405);
nor U15802 (N_15802,N_14323,N_13699);
nor U15803 (N_15803,N_14587,N_12394);
nor U15804 (N_15804,N_13889,N_12414);
or U15805 (N_15805,N_13065,N_12490);
and U15806 (N_15806,N_14559,N_14695);
or U15807 (N_15807,N_14174,N_14442);
nor U15808 (N_15808,N_14282,N_13624);
xnor U15809 (N_15809,N_14997,N_13894);
or U15810 (N_15810,N_13238,N_12272);
or U15811 (N_15811,N_12417,N_13711);
nand U15812 (N_15812,N_14197,N_13272);
and U15813 (N_15813,N_14747,N_12421);
nor U15814 (N_15814,N_13013,N_12340);
nand U15815 (N_15815,N_13864,N_13764);
nand U15816 (N_15816,N_13395,N_14863);
nand U15817 (N_15817,N_12906,N_14263);
or U15818 (N_15818,N_12532,N_13549);
xor U15819 (N_15819,N_12501,N_12230);
nand U15820 (N_15820,N_12614,N_12650);
and U15821 (N_15821,N_12234,N_14143);
and U15822 (N_15822,N_12921,N_13916);
xnor U15823 (N_15823,N_13831,N_13206);
and U15824 (N_15824,N_12816,N_12913);
and U15825 (N_15825,N_14354,N_13491);
nand U15826 (N_15826,N_12530,N_14261);
nand U15827 (N_15827,N_14721,N_14028);
nand U15828 (N_15828,N_12819,N_14013);
nand U15829 (N_15829,N_14580,N_13537);
nor U15830 (N_15830,N_12623,N_12772);
and U15831 (N_15831,N_12177,N_13603);
or U15832 (N_15832,N_13034,N_12568);
xnor U15833 (N_15833,N_13046,N_13150);
nor U15834 (N_15834,N_13135,N_14677);
and U15835 (N_15835,N_14858,N_12449);
nand U15836 (N_15836,N_12133,N_13508);
nand U15837 (N_15837,N_12684,N_12559);
xor U15838 (N_15838,N_13823,N_14546);
xor U15839 (N_15839,N_14627,N_13390);
nand U15840 (N_15840,N_12415,N_14537);
xor U15841 (N_15841,N_13036,N_13666);
or U15842 (N_15842,N_12741,N_14107);
nand U15843 (N_15843,N_14705,N_14891);
nor U15844 (N_15844,N_12474,N_13686);
or U15845 (N_15845,N_14416,N_12026);
nor U15846 (N_15846,N_13406,N_12642);
nor U15847 (N_15847,N_14230,N_14198);
xor U15848 (N_15848,N_13919,N_13051);
nand U15849 (N_15849,N_13986,N_12811);
xnor U15850 (N_15850,N_12056,N_14607);
nor U15851 (N_15851,N_14642,N_12717);
or U15852 (N_15852,N_13965,N_13552);
xnor U15853 (N_15853,N_12418,N_14266);
xor U15854 (N_15854,N_13778,N_12546);
or U15855 (N_15855,N_12086,N_12561);
or U15856 (N_15856,N_12454,N_14014);
nor U15857 (N_15857,N_14479,N_12713);
xor U15858 (N_15858,N_13055,N_14710);
and U15859 (N_15859,N_12744,N_12723);
xor U15860 (N_15860,N_12300,N_13223);
or U15861 (N_15861,N_14703,N_13967);
nand U15862 (N_15862,N_12077,N_14474);
xor U15863 (N_15863,N_14394,N_12577);
nor U15864 (N_15864,N_12276,N_13567);
and U15865 (N_15865,N_13825,N_12953);
nor U15866 (N_15866,N_14020,N_13077);
or U15867 (N_15867,N_14590,N_13420);
nor U15868 (N_15868,N_13858,N_12275);
nor U15869 (N_15869,N_12267,N_13192);
nor U15870 (N_15870,N_13913,N_12236);
or U15871 (N_15871,N_14704,N_13853);
or U15872 (N_15872,N_13985,N_13964);
and U15873 (N_15873,N_12600,N_14083);
nor U15874 (N_15874,N_12477,N_14678);
or U15875 (N_15875,N_12862,N_12587);
nor U15876 (N_15876,N_13810,N_14509);
nor U15877 (N_15877,N_13012,N_14549);
or U15878 (N_15878,N_12101,N_13773);
nor U15879 (N_15879,N_13538,N_12066);
nor U15880 (N_15880,N_12957,N_12318);
nand U15881 (N_15881,N_14485,N_13953);
nand U15882 (N_15882,N_14973,N_13168);
xor U15883 (N_15883,N_12002,N_14903);
nor U15884 (N_15884,N_12586,N_13143);
xor U15885 (N_15885,N_12574,N_13424);
and U15886 (N_15886,N_12453,N_14094);
or U15887 (N_15887,N_13359,N_14058);
nor U15888 (N_15888,N_13108,N_13952);
nor U15889 (N_15889,N_12782,N_14085);
and U15890 (N_15890,N_12500,N_14267);
nand U15891 (N_15891,N_13797,N_13530);
or U15892 (N_15892,N_13106,N_13599);
nand U15893 (N_15893,N_14503,N_14709);
or U15894 (N_15894,N_13848,N_14189);
and U15895 (N_15895,N_13209,N_14183);
nor U15896 (N_15896,N_13447,N_13697);
or U15897 (N_15897,N_14395,N_12425);
nor U15898 (N_15898,N_13672,N_12918);
or U15899 (N_15899,N_14640,N_13421);
nand U15900 (N_15900,N_12774,N_14749);
nand U15901 (N_15901,N_14731,N_12193);
nor U15902 (N_15902,N_13875,N_12067);
and U15903 (N_15903,N_14336,N_12520);
xor U15904 (N_15904,N_12483,N_12122);
xnor U15905 (N_15905,N_12039,N_13190);
and U15906 (N_15906,N_12470,N_13431);
or U15907 (N_15907,N_12882,N_13557);
nor U15908 (N_15908,N_12547,N_12220);
nor U15909 (N_15909,N_14894,N_12909);
or U15910 (N_15910,N_12764,N_12012);
nand U15911 (N_15911,N_12105,N_12205);
and U15912 (N_15912,N_14091,N_12638);
or U15913 (N_15913,N_14915,N_14508);
or U15914 (N_15914,N_12032,N_13927);
xor U15915 (N_15915,N_14908,N_12988);
nand U15916 (N_15916,N_13083,N_14960);
or U15917 (N_15917,N_14008,N_14874);
xor U15918 (N_15918,N_14525,N_14548);
xor U15919 (N_15919,N_12853,N_13479);
xnor U15920 (N_15920,N_14264,N_13355);
or U15921 (N_15921,N_12154,N_13973);
or U15922 (N_15922,N_12084,N_14885);
xnor U15923 (N_15923,N_13350,N_12284);
nor U15924 (N_15924,N_14840,N_13306);
or U15925 (N_15925,N_13205,N_14797);
and U15926 (N_15926,N_13127,N_12152);
or U15927 (N_15927,N_14007,N_12860);
xnor U15928 (N_15928,N_14351,N_12286);
nand U15929 (N_15929,N_13824,N_12594);
nand U15930 (N_15930,N_12695,N_12830);
xor U15931 (N_15931,N_14692,N_14302);
or U15932 (N_15932,N_12450,N_14570);
nor U15933 (N_15933,N_13131,N_13114);
nand U15934 (N_15934,N_14437,N_14357);
or U15935 (N_15935,N_13755,N_13312);
or U15936 (N_15936,N_14102,N_13776);
nor U15937 (N_15937,N_14359,N_12544);
or U15938 (N_15938,N_12529,N_12666);
and U15939 (N_15939,N_14228,N_13847);
xor U15940 (N_15940,N_13525,N_14478);
and U15941 (N_15941,N_13522,N_13280);
nor U15942 (N_15942,N_13870,N_12961);
xnor U15943 (N_15943,N_14754,N_14240);
nor U15944 (N_15944,N_13752,N_12683);
nor U15945 (N_15945,N_13918,N_13211);
and U15946 (N_15946,N_13566,N_14417);
xor U15947 (N_15947,N_13959,N_12082);
xor U15948 (N_15948,N_13141,N_13692);
and U15949 (N_15949,N_14125,N_13467);
or U15950 (N_15950,N_12806,N_12283);
nand U15951 (N_15951,N_12428,N_13742);
and U15952 (N_15952,N_12958,N_13363);
nor U15953 (N_15953,N_12218,N_13002);
and U15954 (N_15954,N_13313,N_14456);
xor U15955 (N_15955,N_14205,N_12209);
nor U15956 (N_15956,N_12201,N_13766);
nand U15957 (N_15957,N_13988,N_13935);
xor U15958 (N_15958,N_12278,N_13203);
or U15959 (N_15959,N_13422,N_12796);
xor U15960 (N_15960,N_13185,N_14554);
nor U15961 (N_15961,N_13721,N_14999);
or U15962 (N_15962,N_12060,N_14762);
nor U15963 (N_15963,N_13749,N_14165);
nor U15964 (N_15964,N_12804,N_14796);
nand U15965 (N_15965,N_14063,N_13356);
xnor U15966 (N_15966,N_13016,N_13511);
xnor U15967 (N_15967,N_13311,N_12720);
nor U15968 (N_15968,N_13024,N_12657);
or U15969 (N_15969,N_13391,N_13622);
or U15970 (N_15970,N_12947,N_12157);
or U15971 (N_15971,N_14589,N_13849);
nor U15972 (N_15972,N_13176,N_13757);
nor U15973 (N_15973,N_13045,N_12445);
nand U15974 (N_15974,N_14972,N_13003);
or U15975 (N_15975,N_13750,N_13267);
nand U15976 (N_15976,N_14181,N_14043);
and U15977 (N_15977,N_12316,N_12376);
xor U15978 (N_15978,N_13885,N_14024);
nor U15979 (N_15979,N_12268,N_14945);
or U15980 (N_15980,N_12581,N_13343);
and U15981 (N_15981,N_14353,N_12156);
nand U15982 (N_15982,N_14350,N_13925);
or U15983 (N_15983,N_13038,N_14694);
and U15984 (N_15984,N_13053,N_13554);
nand U15985 (N_15985,N_14093,N_13400);
and U15986 (N_15986,N_13253,N_13674);
nand U15987 (N_15987,N_12912,N_12887);
xnor U15988 (N_15988,N_14161,N_14925);
xor U15989 (N_15989,N_12640,N_13998);
nor U15990 (N_15990,N_12865,N_14200);
xor U15991 (N_15991,N_12791,N_12715);
or U15992 (N_15992,N_13758,N_13974);
xnor U15993 (N_15993,N_13575,N_14376);
nand U15994 (N_15994,N_12607,N_12798);
and U15995 (N_15995,N_12518,N_13277);
nand U15996 (N_15996,N_12355,N_14825);
or U15997 (N_15997,N_12185,N_13981);
or U15998 (N_15998,N_14786,N_14977);
or U15999 (N_15999,N_14362,N_13708);
or U16000 (N_16000,N_12802,N_14000);
nand U16001 (N_16001,N_12296,N_13154);
nand U16002 (N_16002,N_14430,N_13037);
nand U16003 (N_16003,N_14791,N_13122);
nand U16004 (N_16004,N_13809,N_13172);
and U16005 (N_16005,N_13262,N_14898);
nand U16006 (N_16006,N_12886,N_14337);
or U16007 (N_16007,N_12338,N_14759);
xor U16008 (N_16008,N_12873,N_12572);
xor U16009 (N_16009,N_12250,N_14380);
nand U16010 (N_16010,N_13559,N_12227);
or U16011 (N_16011,N_12933,N_12993);
xor U16012 (N_16012,N_14066,N_13318);
xnor U16013 (N_16013,N_14927,N_14716);
xnor U16014 (N_16014,N_13760,N_12730);
nand U16015 (N_16015,N_12851,N_14803);
and U16016 (N_16016,N_13968,N_13756);
nand U16017 (N_16017,N_12104,N_14119);
and U16018 (N_16018,N_14231,N_12495);
and U16019 (N_16019,N_12874,N_14220);
nor U16020 (N_16020,N_13873,N_12369);
and U16021 (N_16021,N_12541,N_13453);
or U16022 (N_16022,N_14774,N_12482);
and U16023 (N_16023,N_13655,N_14128);
xnor U16024 (N_16024,N_14656,N_12986);
and U16025 (N_16025,N_12781,N_12332);
nor U16026 (N_16026,N_13386,N_13896);
nand U16027 (N_16027,N_12857,N_12951);
and U16028 (N_16028,N_12625,N_13745);
xnor U16029 (N_16029,N_14486,N_12915);
xor U16030 (N_16030,N_14526,N_14850);
nor U16031 (N_16031,N_12672,N_14739);
xnor U16032 (N_16032,N_13930,N_13772);
or U16033 (N_16033,N_13337,N_12940);
nor U16034 (N_16034,N_12697,N_12763);
or U16035 (N_16035,N_13360,N_14436);
or U16036 (N_16036,N_14463,N_13087);
xnor U16037 (N_16037,N_13912,N_12053);
or U16038 (N_16038,N_12027,N_13454);
xnor U16039 (N_16039,N_13370,N_13661);
nand U16040 (N_16040,N_13561,N_12323);
xnor U16041 (N_16041,N_14984,N_14250);
xor U16042 (N_16042,N_12848,N_14155);
nand U16043 (N_16043,N_14965,N_13039);
and U16044 (N_16044,N_12923,N_13808);
nor U16045 (N_16045,N_14361,N_12747);
nor U16046 (N_16046,N_13084,N_12761);
nand U16047 (N_16047,N_12087,N_14686);
nand U16048 (N_16048,N_14611,N_13887);
nand U16049 (N_16049,N_12635,N_13834);
and U16050 (N_16050,N_13099,N_14339);
nand U16051 (N_16051,N_12299,N_13480);
or U16052 (N_16052,N_13274,N_14127);
or U16053 (N_16053,N_13136,N_14318);
or U16054 (N_16054,N_14743,N_14622);
xnor U16055 (N_16055,N_14968,N_14500);
nand U16056 (N_16056,N_12895,N_13326);
nand U16057 (N_16057,N_14533,N_12560);
nor U16058 (N_16058,N_12438,N_12711);
xnor U16059 (N_16059,N_14768,N_13116);
nand U16060 (N_16060,N_14652,N_13628);
xnor U16061 (N_16061,N_14284,N_13647);
nand U16062 (N_16062,N_12892,N_12313);
nor U16063 (N_16063,N_13646,N_12554);
or U16064 (N_16064,N_12377,N_14286);
nor U16065 (N_16065,N_12908,N_12750);
and U16066 (N_16066,N_13696,N_14601);
nor U16067 (N_16067,N_12052,N_14779);
nor U16068 (N_16068,N_12844,N_12219);
nor U16069 (N_16069,N_13498,N_12658);
xnor U16070 (N_16070,N_14079,N_12959);
nand U16071 (N_16071,N_14340,N_14491);
and U16072 (N_16072,N_12217,N_13501);
and U16073 (N_16073,N_13945,N_12492);
nand U16074 (N_16074,N_13288,N_14420);
and U16075 (N_16075,N_12435,N_12917);
nand U16076 (N_16076,N_14594,N_14413);
nand U16077 (N_16077,N_13432,N_14619);
nor U16078 (N_16078,N_14959,N_12694);
or U16079 (N_16079,N_13943,N_14750);
nor U16080 (N_16080,N_14273,N_12708);
nor U16081 (N_16081,N_13445,N_14691);
xor U16082 (N_16082,N_12427,N_12328);
or U16083 (N_16083,N_13227,N_12080);
xor U16084 (N_16084,N_12681,N_14955);
nand U16085 (N_16085,N_13822,N_12466);
nor U16086 (N_16086,N_14502,N_12493);
xnor U16087 (N_16087,N_14628,N_14604);
xnor U16088 (N_16088,N_14810,N_12624);
or U16089 (N_16089,N_12314,N_13886);
and U16090 (N_16090,N_12692,N_12952);
xnor U16091 (N_16091,N_14322,N_12884);
or U16092 (N_16092,N_13789,N_12834);
nor U16093 (N_16093,N_13487,N_12540);
nor U16094 (N_16094,N_13269,N_13457);
nor U16095 (N_16095,N_14192,N_12610);
xor U16096 (N_16096,N_12289,N_12974);
and U16097 (N_16097,N_13417,N_14132);
nand U16098 (N_16098,N_14792,N_13560);
and U16099 (N_16099,N_12054,N_14251);
nor U16100 (N_16100,N_13668,N_14100);
and U16101 (N_16101,N_12673,N_13198);
xor U16102 (N_16102,N_13329,N_14258);
or U16103 (N_16103,N_14593,N_13837);
or U16104 (N_16104,N_12322,N_14547);
nand U16105 (N_16105,N_12359,N_14236);
or U16106 (N_16106,N_12155,N_14773);
xnor U16107 (N_16107,N_14953,N_14576);
xor U16108 (N_16108,N_13376,N_12137);
nor U16109 (N_16109,N_12309,N_14662);
xnor U16110 (N_16110,N_13931,N_14005);
xnor U16111 (N_16111,N_12889,N_13470);
nor U16112 (N_16112,N_14829,N_14461);
nor U16113 (N_16113,N_13171,N_13728);
nor U16114 (N_16114,N_14689,N_13090);
nand U16115 (N_16115,N_14864,N_14139);
xnor U16116 (N_16116,N_13978,N_14140);
nor U16117 (N_16117,N_13158,N_13677);
or U16118 (N_16118,N_14928,N_14475);
or U16119 (N_16119,N_12245,N_13380);
nand U16120 (N_16120,N_13133,N_14837);
and U16121 (N_16121,N_14505,N_14738);
or U16122 (N_16122,N_13512,N_12162);
or U16123 (N_16123,N_14343,N_13251);
nand U16124 (N_16124,N_14592,N_13645);
nor U16125 (N_16125,N_12228,N_12075);
and U16126 (N_16126,N_13155,N_12538);
and U16127 (N_16127,N_14304,N_13011);
or U16128 (N_16128,N_13466,N_13638);
and U16129 (N_16129,N_12553,N_12397);
or U16130 (N_16130,N_14297,N_12187);
and U16131 (N_16131,N_13236,N_14347);
or U16132 (N_16132,N_13693,N_12038);
xor U16133 (N_16133,N_13897,N_13219);
nor U16134 (N_16134,N_13681,N_13556);
nor U16135 (N_16135,N_12971,N_13324);
xor U16136 (N_16136,N_14971,N_13347);
nand U16137 (N_16137,N_14499,N_12562);
nor U16138 (N_16138,N_12074,N_14620);
xnor U16139 (N_16139,N_12011,N_14400);
or U16140 (N_16140,N_14279,N_12766);
xnor U16141 (N_16141,N_13999,N_12584);
and U16142 (N_16142,N_12771,N_13569);
xor U16143 (N_16143,N_12932,N_14659);
nor U16144 (N_16144,N_13450,N_13047);
and U16145 (N_16145,N_12337,N_12987);
or U16146 (N_16146,N_14422,N_14848);
xnor U16147 (N_16147,N_14685,N_13404);
and U16148 (N_16148,N_12677,N_14892);
nand U16149 (N_16149,N_14987,N_12174);
nand U16150 (N_16150,N_14564,N_14665);
xor U16151 (N_16151,N_12789,N_13095);
or U16152 (N_16152,N_14204,N_12352);
or U16153 (N_16153,N_14664,N_12294);
nand U16154 (N_16154,N_14539,N_14798);
and U16155 (N_16155,N_13477,N_14597);
xor U16156 (N_16156,N_14929,N_12465);
or U16157 (N_16157,N_12237,N_14030);
xor U16158 (N_16158,N_13670,N_13958);
or U16159 (N_16159,N_14224,N_13113);
nand U16160 (N_16160,N_14110,N_14375);
nand U16161 (N_16161,N_13160,N_14501);
and U16162 (N_16162,N_13463,N_13641);
xnor U16163 (N_16163,N_12839,N_14454);
xnor U16164 (N_16164,N_12285,N_14309);
xnor U16165 (N_16165,N_14333,N_13592);
xnor U16166 (N_16166,N_14440,N_12696);
or U16167 (N_16167,N_14877,N_14141);
or U16168 (N_16168,N_14082,N_13957);
or U16169 (N_16169,N_13676,N_13734);
nor U16170 (N_16170,N_13987,N_12164);
nand U16171 (N_16171,N_12824,N_12675);
or U16172 (N_16172,N_12362,N_14398);
nand U16173 (N_16173,N_12439,N_13632);
or U16174 (N_16174,N_13435,N_14923);
or U16175 (N_16175,N_12652,N_14658);
and U16176 (N_16176,N_12350,N_12748);
nor U16177 (N_16177,N_12007,N_14637);
nand U16178 (N_16178,N_14992,N_12111);
or U16179 (N_16179,N_12868,N_12647);
nand U16180 (N_16180,N_12856,N_12793);
and U16181 (N_16181,N_13125,N_12480);
nand U16182 (N_16182,N_14055,N_13367);
nor U16183 (N_16183,N_14195,N_14772);
and U16184 (N_16184,N_13098,N_13460);
nor U16185 (N_16185,N_13867,N_14418);
xnor U16186 (N_16186,N_13612,N_14707);
and U16187 (N_16187,N_14669,N_14646);
or U16188 (N_16188,N_13779,N_12942);
xor U16189 (N_16189,N_13841,N_14133);
or U16190 (N_16190,N_14404,N_12124);
nand U16191 (N_16191,N_13275,N_13147);
or U16192 (N_16192,N_12160,N_14517);
and U16193 (N_16193,N_14146,N_14784);
nand U16194 (N_16194,N_12845,N_13936);
xor U16195 (N_16195,N_14157,N_12785);
and U16196 (N_16196,N_12843,N_14312);
nor U16197 (N_16197,N_13519,N_13140);
or U16198 (N_16198,N_12171,N_14639);
xor U16199 (N_16199,N_13461,N_14072);
or U16200 (N_16200,N_12327,N_13663);
nor U16201 (N_16201,N_13078,N_14233);
or U16202 (N_16202,N_14845,N_13517);
xor U16203 (N_16203,N_12977,N_13244);
xor U16204 (N_16204,N_12021,N_13368);
nor U16205 (N_16205,N_13446,N_13427);
and U16206 (N_16206,N_13866,N_14237);
nor U16207 (N_16207,N_12835,N_12386);
xor U16208 (N_16208,N_13702,N_13713);
or U16209 (N_16209,N_13270,N_13583);
xnor U16210 (N_16210,N_14345,N_14144);
or U16211 (N_16211,N_14938,N_12253);
xor U16212 (N_16212,N_12762,N_14631);
or U16213 (N_16213,N_13571,N_14149);
nor U16214 (N_16214,N_13027,N_13019);
and U16215 (N_16215,N_13555,N_12864);
or U16216 (N_16216,N_13658,N_13230);
xor U16217 (N_16217,N_14182,N_12413);
xnor U16218 (N_16218,N_12046,N_13126);
and U16219 (N_16219,N_14148,N_13598);
xor U16220 (N_16220,N_13905,N_14888);
nor U16221 (N_16221,N_12885,N_13855);
xor U16222 (N_16222,N_13301,N_12380);
or U16223 (N_16223,N_14934,N_12487);
nand U16224 (N_16224,N_12140,N_13362);
or U16225 (N_16225,N_13718,N_12042);
or U16226 (N_16226,N_12788,N_13436);
or U16227 (N_16227,N_13863,N_13397);
or U16228 (N_16228,N_12707,N_13540);
or U16229 (N_16229,N_13449,N_14788);
and U16230 (N_16230,N_12269,N_13074);
and U16231 (N_16231,N_13532,N_14378);
and U16232 (N_16232,N_12745,N_14575);
xor U16233 (N_16233,N_13637,N_12605);
or U16234 (N_16234,N_12233,N_12877);
or U16235 (N_16235,N_13396,N_12491);
nor U16236 (N_16236,N_13088,N_13458);
and U16237 (N_16237,N_14847,N_12664);
and U16238 (N_16238,N_12150,N_13228);
and U16239 (N_16239,N_13648,N_12291);
and U16240 (N_16240,N_12955,N_14819);
xor U16241 (N_16241,N_12025,N_13751);
or U16242 (N_16242,N_14207,N_14806);
or U16243 (N_16243,N_14591,N_13030);
nand U16244 (N_16244,N_14986,N_13544);
xnor U16245 (N_16245,N_12765,N_14048);
and U16246 (N_16246,N_12621,N_13217);
nor U16247 (N_16247,N_13753,N_12545);
xor U16248 (N_16248,N_12496,N_14269);
nand U16249 (N_16249,N_12282,N_12622);
and U16250 (N_16250,N_12828,N_14745);
xor U16251 (N_16251,N_12800,N_12257);
and U16252 (N_16252,N_12740,N_13167);
or U16253 (N_16253,N_12646,N_14572);
xnor U16254 (N_16254,N_12029,N_12277);
nor U16255 (N_16255,N_14433,N_14001);
nand U16256 (N_16256,N_12254,N_12878);
nor U16257 (N_16257,N_13496,N_12519);
or U16258 (N_16258,N_13513,N_12069);
or U16259 (N_16259,N_14077,N_12317);
nand U16260 (N_16260,N_12693,N_13263);
or U16261 (N_16261,N_14558,N_12243);
xor U16262 (N_16262,N_13414,N_14831);
nor U16263 (N_16263,N_14285,N_14783);
nor U16264 (N_16264,N_13026,N_12899);
nand U16265 (N_16265,N_12863,N_13748);
xor U16266 (N_16266,N_12631,N_13595);
and U16267 (N_16267,N_14319,N_12710);
nand U16268 (N_16268,N_13308,N_13654);
nor U16269 (N_16269,N_12442,N_12385);
and U16270 (N_16270,N_13770,N_12213);
or U16271 (N_16271,N_12395,N_12767);
and U16272 (N_16272,N_14957,N_14196);
nand U16273 (N_16273,N_14477,N_13361);
xor U16274 (N_16274,N_12161,N_14390);
or U16275 (N_16275,N_12704,N_13579);
and U16276 (N_16276,N_13119,N_13507);
nor U16277 (N_16277,N_12516,N_12206);
or U16278 (N_16278,N_14964,N_14919);
nor U16279 (N_16279,N_14621,N_13040);
or U16280 (N_16280,N_13593,N_13000);
nand U16281 (N_16281,N_12281,N_14568);
nor U16282 (N_16282,N_13826,N_12571);
nand U16283 (N_16283,N_14993,N_13565);
or U16284 (N_16284,N_13528,N_13256);
and U16285 (N_16285,N_14300,N_12113);
nand U16286 (N_16286,N_14476,N_13418);
nor U16287 (N_16287,N_14106,N_14374);
nand U16288 (N_16288,N_13895,N_12265);
xor U16289 (N_16289,N_12349,N_14046);
nor U16290 (N_16290,N_12169,N_12416);
nor U16291 (N_16291,N_13225,N_13615);
nor U16292 (N_16292,N_14052,N_14855);
and U16293 (N_16293,N_14087,N_13675);
nand U16294 (N_16294,N_12446,N_12537);
xor U16295 (N_16295,N_13152,N_12045);
nand U16296 (N_16296,N_13629,N_14901);
and U16297 (N_16297,N_14225,N_14811);
and U16298 (N_16298,N_14718,N_14519);
or U16299 (N_16299,N_14281,N_14171);
nand U16300 (N_16300,N_13928,N_14402);
xor U16301 (N_16301,N_14355,N_14408);
or U16302 (N_16302,N_13411,N_12055);
or U16303 (N_16303,N_13096,N_13761);
and U16304 (N_16304,N_12259,N_12019);
or U16305 (N_16305,N_14296,N_12665);
xnor U16306 (N_16306,N_12049,N_12746);
and U16307 (N_16307,N_12687,N_12690);
or U16308 (N_16308,N_14813,N_14722);
nand U16309 (N_16309,N_14816,N_12810);
xor U16310 (N_16310,N_14719,N_12983);
xor U16311 (N_16311,N_14846,N_12457);
nor U16312 (N_16312,N_13594,N_14781);
nand U16313 (N_16313,N_14995,N_12644);
xor U16314 (N_16314,N_12948,N_14349);
nand U16315 (N_16315,N_14679,N_13159);
or U16316 (N_16316,N_12009,N_14663);
and U16317 (N_16317,N_14136,N_14967);
and U16318 (N_16318,N_14793,N_13264);
nand U16319 (N_16319,N_12116,N_13694);
xnor U16320 (N_16320,N_13976,N_14907);
xnor U16321 (N_16321,N_12526,N_13075);
nand U16322 (N_16322,N_13054,N_14860);
nor U16323 (N_16323,N_14369,N_13683);
or U16324 (N_16324,N_14556,N_14881);
nand U16325 (N_16325,N_12204,N_13257);
or U16326 (N_16326,N_14978,N_14419);
nor U16327 (N_16327,N_12573,N_14170);
and U16328 (N_16328,N_12682,N_12949);
and U16329 (N_16329,N_13877,N_12576);
nand U16330 (N_16330,N_14496,N_13585);
xnor U16331 (N_16331,N_14600,N_14112);
or U16332 (N_16332,N_12375,N_12718);
or U16333 (N_16333,N_14235,N_13626);
or U16334 (N_16334,N_13865,N_14751);
or U16335 (N_16335,N_12110,N_14818);
nand U16336 (N_16336,N_13189,N_13180);
or U16337 (N_16337,N_13281,N_13433);
and U16338 (N_16338,N_12645,N_13472);
and U16339 (N_16339,N_13934,N_14884);
nor U16340 (N_16340,N_12085,N_14131);
or U16341 (N_16341,N_13712,N_14641);
nor U16342 (N_16342,N_12548,N_12714);
nand U16343 (N_16343,N_13035,N_14857);
nand U16344 (N_16344,N_12729,N_13505);
xor U16345 (N_16345,N_13490,N_14039);
or U16346 (N_16346,N_12636,N_14326);
xor U16347 (N_16347,N_13315,N_14215);
and U16348 (N_16348,N_13746,N_12634);
and U16349 (N_16349,N_14111,N_14649);
nor U16350 (N_16350,N_14018,N_13273);
xnor U16351 (N_16351,N_13900,N_12836);
or U16352 (N_16352,N_14307,N_14403);
and U16353 (N_16353,N_13835,N_14511);
or U16354 (N_16354,N_12288,N_13249);
nor U16355 (N_16355,N_14932,N_12147);
nor U16356 (N_16356,N_13033,N_12922);
nand U16357 (N_16357,N_12662,N_14814);
and U16358 (N_16358,N_14448,N_13465);
and U16359 (N_16359,N_12700,N_13299);
nor U16360 (N_16360,N_13130,N_14410);
xnor U16361 (N_16361,N_13690,N_13782);
or U16362 (N_16362,N_14520,N_12010);
xor U16363 (N_16363,N_13724,N_13572);
nor U16364 (N_16364,N_13868,N_13774);
and U16365 (N_16365,N_12258,N_13785);
xnor U16366 (N_16366,N_12368,N_12790);
xnor U16367 (N_16367,N_14017,N_13412);
nor U16368 (N_16368,N_12563,N_14194);
and U16369 (N_16369,N_14935,N_14497);
nand U16370 (N_16370,N_13210,N_13975);
nand U16371 (N_16371,N_13004,N_14135);
nor U16372 (N_16372,N_12803,N_13535);
and U16373 (N_16373,N_14839,N_14795);
xor U16374 (N_16374,N_13489,N_14724);
nand U16375 (N_16375,N_14869,N_12139);
or U16376 (N_16376,N_14633,N_14040);
nor U16377 (N_16377,N_13669,N_13220);
and U16378 (N_16378,N_14481,N_12656);
nor U16379 (N_16379,N_12840,N_14713);
nor U16380 (N_16380,N_12846,N_12639);
nand U16381 (N_16381,N_12608,N_14295);
and U16382 (N_16382,N_13107,N_12858);
nand U16383 (N_16383,N_13741,N_13950);
or U16384 (N_16384,N_12566,N_12210);
and U16385 (N_16385,N_12699,N_13664);
xnor U16386 (N_16386,N_14889,N_12847);
xor U16387 (N_16387,N_12894,N_14291);
nand U16388 (N_16388,N_14725,N_13187);
and U16389 (N_16389,N_13144,N_14262);
nor U16390 (N_16390,N_14752,N_12513);
nand U16391 (N_16391,N_12628,N_12613);
and U16392 (N_16392,N_13023,N_12440);
nor U16393 (N_16393,N_13990,N_12616);
xor U16394 (N_16394,N_13246,N_13969);
and U16395 (N_16395,N_12502,N_12430);
nor U16396 (N_16396,N_13423,N_12769);
or U16397 (N_16397,N_13377,N_12461);
nand U16398 (N_16398,N_12444,N_14657);
xor U16399 (N_16399,N_12371,N_13322);
or U16400 (N_16400,N_13961,N_13783);
nor U16401 (N_16401,N_12916,N_12020);
and U16402 (N_16402,N_14366,N_13138);
nand U16403 (N_16403,N_13165,N_12405);
xnor U16404 (N_16404,N_14358,N_14574);
nand U16405 (N_16405,N_13408,N_13409);
or U16406 (N_16406,N_14153,N_12076);
or U16407 (N_16407,N_14737,N_14897);
nor U16408 (N_16408,N_12330,N_12601);
nand U16409 (N_16409,N_14854,N_13258);
or U16410 (N_16410,N_12073,N_14372);
and U16411 (N_16411,N_13861,N_13813);
or U16412 (N_16412,N_13743,N_12109);
and U16413 (N_16413,N_13725,N_13307);
and U16414 (N_16414,N_14439,N_12735);
xor U16415 (N_16415,N_13103,N_13903);
xnor U16416 (N_16416,N_13204,N_14057);
xnor U16417 (N_16417,N_14672,N_14483);
xor U16418 (N_16418,N_13636,N_12890);
nand U16419 (N_16419,N_12589,N_14252);
nor U16420 (N_16420,N_12599,N_13008);
or U16421 (N_16421,N_12404,N_14736);
nor U16422 (N_16422,N_12342,N_14698);
nor U16423 (N_16423,N_12712,N_13232);
or U16424 (N_16424,N_13500,N_12979);
nand U16425 (N_16425,N_14624,N_14804);
and U16426 (N_16426,N_13731,N_14764);
nor U16427 (N_16427,N_13678,N_12361);
nor U16428 (N_16428,N_14625,N_12626);
and U16429 (N_16429,N_12374,N_14313);
nor U16430 (N_16430,N_13323,N_14697);
xnor U16431 (N_16431,N_13309,N_12910);
nand U16432 (N_16432,N_12904,N_13732);
and U16433 (N_16433,N_13679,N_14565);
or U16434 (N_16434,N_12100,N_14188);
or U16435 (N_16435,N_13947,N_13093);
or U16436 (N_16436,N_13245,N_12859);
or U16437 (N_16437,N_13009,N_13316);
xor U16438 (N_16438,N_14667,N_13403);
or U16439 (N_16439,N_12306,N_12937);
nand U16440 (N_16440,N_12467,N_14512);
nor U16441 (N_16441,N_14916,N_14893);
or U16442 (N_16442,N_14912,N_13709);
and U16443 (N_16443,N_13584,N_13754);
and U16444 (N_16444,N_12944,N_13888);
or U16445 (N_16445,N_14729,N_13997);
nor U16446 (N_16446,N_14384,N_14382);
and U16447 (N_16447,N_14222,N_12962);
nand U16448 (N_16448,N_14545,N_13759);
nor U16449 (N_16449,N_13526,N_14835);
nand U16450 (N_16450,N_14457,N_12061);
nor U16451 (N_16451,N_14070,N_12310);
nor U16452 (N_16452,N_14051,N_14379);
and U16453 (N_16453,N_13484,N_12134);
nand U16454 (N_16454,N_12503,N_13940);
and U16455 (N_16455,N_12173,N_13765);
nand U16456 (N_16456,N_14115,N_12755);
xor U16457 (N_16457,N_14019,N_14515);
or U16458 (N_16458,N_13852,N_13181);
nor U16459 (N_16459,N_14760,N_12787);
nor U16460 (N_16460,N_14523,N_12422);
xnor U16461 (N_16461,N_12389,N_14807);
and U16462 (N_16462,N_12367,N_12331);
nor U16463 (N_16463,N_12241,N_14644);
nor U16464 (N_16464,N_14579,N_12618);
or U16465 (N_16465,N_13402,N_13385);
nor U16466 (N_16466,N_12382,N_12855);
nand U16467 (N_16467,N_12231,N_14489);
and U16468 (N_16468,N_12898,N_12985);
nor U16469 (N_16469,N_14306,N_13452);
and U16470 (N_16470,N_12679,N_14780);
nand U16471 (N_16471,N_14966,N_12867);
nor U16472 (N_16472,N_14944,N_12515);
nor U16473 (N_16473,N_14730,N_14617);
nand U16474 (N_16474,N_13139,N_14406);
or U16475 (N_16475,N_12078,N_14494);
and U16476 (N_16476,N_14946,N_13001);
nor U16477 (N_16477,N_14065,N_14670);
nand U16478 (N_16478,N_12391,N_12274);
nor U16479 (N_16479,N_13616,N_13285);
xor U16480 (N_16480,N_14735,N_14586);
or U16481 (N_16481,N_13588,N_14080);
or U16482 (N_16482,N_13121,N_12668);
and U16483 (N_16483,N_14742,N_13383);
and U16484 (N_16484,N_12383,N_14790);
nor U16485 (N_16485,N_14223,N_13438);
or U16486 (N_16486,N_14870,N_13982);
nor U16487 (N_16487,N_12151,N_12163);
and U16488 (N_16488,N_13440,N_12379);
nand U16489 (N_16489,N_14154,N_14543);
nor U16490 (N_16490,N_13091,N_12536);
or U16491 (N_16491,N_12372,N_12271);
nor U16492 (N_16492,N_14150,N_14596);
and U16493 (N_16493,N_13202,N_14674);
and U16494 (N_16494,N_13820,N_13798);
and U16495 (N_16495,N_12351,N_12727);
and U16496 (N_16496,N_13737,N_12356);
and U16497 (N_16497,N_14243,N_14193);
xnor U16498 (N_16498,N_13341,N_14370);
nor U16499 (N_16499,N_12795,N_13703);
nor U16500 (N_16500,N_12698,N_12605);
xor U16501 (N_16501,N_13272,N_12509);
nand U16502 (N_16502,N_12220,N_13895);
or U16503 (N_16503,N_13344,N_12185);
or U16504 (N_16504,N_12424,N_13663);
or U16505 (N_16505,N_14190,N_13984);
or U16506 (N_16506,N_14226,N_13073);
xor U16507 (N_16507,N_12996,N_14724);
or U16508 (N_16508,N_14343,N_13555);
nor U16509 (N_16509,N_13874,N_13267);
nor U16510 (N_16510,N_14000,N_12081);
and U16511 (N_16511,N_12734,N_13121);
nand U16512 (N_16512,N_14808,N_13149);
nand U16513 (N_16513,N_14576,N_13417);
xnor U16514 (N_16514,N_13099,N_14562);
xnor U16515 (N_16515,N_13919,N_13715);
xor U16516 (N_16516,N_12740,N_13266);
nor U16517 (N_16517,N_12139,N_14620);
xor U16518 (N_16518,N_12736,N_12405);
xor U16519 (N_16519,N_13900,N_12848);
nand U16520 (N_16520,N_14396,N_14778);
and U16521 (N_16521,N_14047,N_12939);
or U16522 (N_16522,N_12168,N_13882);
nand U16523 (N_16523,N_13651,N_12698);
xor U16524 (N_16524,N_12327,N_14738);
and U16525 (N_16525,N_14428,N_12249);
xor U16526 (N_16526,N_13995,N_13143);
nor U16527 (N_16527,N_14852,N_12600);
nor U16528 (N_16528,N_13360,N_13833);
and U16529 (N_16529,N_14531,N_12970);
or U16530 (N_16530,N_12982,N_12415);
or U16531 (N_16531,N_14175,N_14190);
xnor U16532 (N_16532,N_14689,N_13262);
nand U16533 (N_16533,N_12139,N_12225);
and U16534 (N_16534,N_13756,N_12073);
xor U16535 (N_16535,N_14763,N_13515);
and U16536 (N_16536,N_12163,N_13286);
and U16537 (N_16537,N_14763,N_13013);
and U16538 (N_16538,N_14965,N_14609);
or U16539 (N_16539,N_14532,N_13960);
and U16540 (N_16540,N_14443,N_12837);
nand U16541 (N_16541,N_14278,N_13421);
and U16542 (N_16542,N_13288,N_12024);
or U16543 (N_16543,N_14087,N_13522);
or U16544 (N_16544,N_13582,N_12732);
xor U16545 (N_16545,N_12337,N_13126);
nand U16546 (N_16546,N_12216,N_13314);
xor U16547 (N_16547,N_14317,N_13258);
or U16548 (N_16548,N_13814,N_12804);
and U16549 (N_16549,N_13586,N_14058);
xor U16550 (N_16550,N_13461,N_14486);
xor U16551 (N_16551,N_13707,N_12684);
and U16552 (N_16552,N_12465,N_12859);
or U16553 (N_16553,N_13180,N_13139);
and U16554 (N_16554,N_12060,N_13874);
or U16555 (N_16555,N_14786,N_13215);
nor U16556 (N_16556,N_12155,N_12400);
nor U16557 (N_16557,N_13673,N_14427);
or U16558 (N_16558,N_12245,N_13778);
xor U16559 (N_16559,N_14531,N_13257);
or U16560 (N_16560,N_14005,N_14262);
nor U16561 (N_16561,N_12668,N_14334);
xnor U16562 (N_16562,N_12408,N_14572);
xor U16563 (N_16563,N_14735,N_12345);
and U16564 (N_16564,N_13744,N_12809);
nand U16565 (N_16565,N_13430,N_13410);
and U16566 (N_16566,N_12014,N_14816);
nor U16567 (N_16567,N_12604,N_13781);
nor U16568 (N_16568,N_12260,N_12419);
xnor U16569 (N_16569,N_13865,N_12841);
xnor U16570 (N_16570,N_14990,N_14718);
and U16571 (N_16571,N_13643,N_12595);
nand U16572 (N_16572,N_14612,N_12817);
nand U16573 (N_16573,N_13915,N_14536);
xnor U16574 (N_16574,N_13062,N_13502);
or U16575 (N_16575,N_13008,N_13435);
xnor U16576 (N_16576,N_12224,N_14220);
xor U16577 (N_16577,N_14328,N_13885);
nor U16578 (N_16578,N_14420,N_12492);
nand U16579 (N_16579,N_12551,N_14436);
nand U16580 (N_16580,N_13358,N_13328);
nor U16581 (N_16581,N_13249,N_12435);
and U16582 (N_16582,N_14208,N_13247);
nor U16583 (N_16583,N_13890,N_14185);
nand U16584 (N_16584,N_13804,N_12155);
and U16585 (N_16585,N_12942,N_12865);
xnor U16586 (N_16586,N_14399,N_14795);
or U16587 (N_16587,N_13240,N_13899);
and U16588 (N_16588,N_14809,N_12827);
nand U16589 (N_16589,N_12303,N_13820);
xnor U16590 (N_16590,N_12810,N_13050);
or U16591 (N_16591,N_14098,N_12037);
or U16592 (N_16592,N_13785,N_13963);
or U16593 (N_16593,N_13114,N_14970);
or U16594 (N_16594,N_13645,N_14491);
and U16595 (N_16595,N_13228,N_14829);
xnor U16596 (N_16596,N_14977,N_12637);
nor U16597 (N_16597,N_14747,N_13930);
nor U16598 (N_16598,N_12189,N_14700);
or U16599 (N_16599,N_13691,N_13138);
and U16600 (N_16600,N_13340,N_13341);
and U16601 (N_16601,N_14632,N_14401);
or U16602 (N_16602,N_12292,N_14131);
or U16603 (N_16603,N_12851,N_14596);
xnor U16604 (N_16604,N_14573,N_13423);
nand U16605 (N_16605,N_13902,N_13869);
and U16606 (N_16606,N_12990,N_14518);
or U16607 (N_16607,N_13970,N_14847);
nand U16608 (N_16608,N_12730,N_12193);
or U16609 (N_16609,N_12797,N_13534);
xnor U16610 (N_16610,N_13701,N_12162);
xor U16611 (N_16611,N_12405,N_14684);
nand U16612 (N_16612,N_12993,N_14301);
or U16613 (N_16613,N_14135,N_14084);
xor U16614 (N_16614,N_13011,N_12019);
nor U16615 (N_16615,N_14069,N_14655);
nand U16616 (N_16616,N_14856,N_12412);
nor U16617 (N_16617,N_14776,N_13946);
or U16618 (N_16618,N_13725,N_14159);
and U16619 (N_16619,N_13774,N_14440);
nor U16620 (N_16620,N_14752,N_14126);
and U16621 (N_16621,N_13958,N_14934);
or U16622 (N_16622,N_14657,N_14242);
xor U16623 (N_16623,N_12389,N_14270);
nand U16624 (N_16624,N_13187,N_12264);
and U16625 (N_16625,N_14534,N_13395);
nor U16626 (N_16626,N_14227,N_13654);
xnor U16627 (N_16627,N_14042,N_13038);
and U16628 (N_16628,N_13299,N_13066);
or U16629 (N_16629,N_12467,N_14701);
or U16630 (N_16630,N_13958,N_13759);
nand U16631 (N_16631,N_12672,N_14443);
or U16632 (N_16632,N_14889,N_12096);
nand U16633 (N_16633,N_12331,N_14040);
nand U16634 (N_16634,N_12759,N_12670);
nand U16635 (N_16635,N_12732,N_13526);
xor U16636 (N_16636,N_12979,N_12607);
xnor U16637 (N_16637,N_13043,N_13214);
nor U16638 (N_16638,N_12083,N_12175);
nand U16639 (N_16639,N_13028,N_12353);
nor U16640 (N_16640,N_13838,N_14930);
nand U16641 (N_16641,N_12166,N_12413);
or U16642 (N_16642,N_12563,N_14723);
nand U16643 (N_16643,N_14886,N_13453);
or U16644 (N_16644,N_13998,N_12731);
nor U16645 (N_16645,N_14282,N_14246);
nor U16646 (N_16646,N_12957,N_14228);
or U16647 (N_16647,N_13023,N_12391);
and U16648 (N_16648,N_14521,N_12860);
nor U16649 (N_16649,N_14728,N_12465);
and U16650 (N_16650,N_13881,N_12796);
or U16651 (N_16651,N_13495,N_14519);
nor U16652 (N_16652,N_13567,N_12046);
nor U16653 (N_16653,N_13141,N_14727);
nor U16654 (N_16654,N_12536,N_12975);
nor U16655 (N_16655,N_14516,N_13340);
nor U16656 (N_16656,N_13971,N_13869);
nand U16657 (N_16657,N_14945,N_12515);
nand U16658 (N_16658,N_14133,N_14442);
nor U16659 (N_16659,N_13001,N_12481);
nor U16660 (N_16660,N_14976,N_14268);
or U16661 (N_16661,N_13852,N_12881);
nor U16662 (N_16662,N_13744,N_14238);
or U16663 (N_16663,N_12532,N_14641);
nor U16664 (N_16664,N_12568,N_13673);
nor U16665 (N_16665,N_14373,N_12040);
and U16666 (N_16666,N_14665,N_12174);
nor U16667 (N_16667,N_13033,N_12562);
or U16668 (N_16668,N_12199,N_12441);
nand U16669 (N_16669,N_12945,N_12666);
or U16670 (N_16670,N_13010,N_12898);
and U16671 (N_16671,N_14100,N_12370);
nor U16672 (N_16672,N_12606,N_12047);
xor U16673 (N_16673,N_14321,N_12462);
and U16674 (N_16674,N_12311,N_14397);
and U16675 (N_16675,N_13569,N_14335);
nand U16676 (N_16676,N_12525,N_12581);
and U16677 (N_16677,N_14110,N_14244);
and U16678 (N_16678,N_13057,N_13148);
nor U16679 (N_16679,N_13132,N_13093);
xnor U16680 (N_16680,N_14486,N_13180);
nor U16681 (N_16681,N_12176,N_12516);
and U16682 (N_16682,N_14680,N_12537);
xnor U16683 (N_16683,N_13022,N_13621);
xor U16684 (N_16684,N_12975,N_13565);
nor U16685 (N_16685,N_14530,N_12543);
nand U16686 (N_16686,N_14471,N_13437);
nor U16687 (N_16687,N_13881,N_14845);
nor U16688 (N_16688,N_13337,N_12822);
or U16689 (N_16689,N_13896,N_14075);
or U16690 (N_16690,N_14354,N_13580);
nor U16691 (N_16691,N_13414,N_14029);
or U16692 (N_16692,N_13934,N_13268);
and U16693 (N_16693,N_14221,N_13758);
nand U16694 (N_16694,N_14831,N_12458);
nand U16695 (N_16695,N_14676,N_14370);
nand U16696 (N_16696,N_13597,N_14942);
and U16697 (N_16697,N_13977,N_14190);
or U16698 (N_16698,N_12525,N_14465);
and U16699 (N_16699,N_13615,N_13018);
or U16700 (N_16700,N_12548,N_14183);
xnor U16701 (N_16701,N_12008,N_14895);
or U16702 (N_16702,N_12832,N_13098);
or U16703 (N_16703,N_14532,N_14112);
nor U16704 (N_16704,N_13960,N_13181);
nor U16705 (N_16705,N_13231,N_12097);
or U16706 (N_16706,N_13429,N_12721);
xnor U16707 (N_16707,N_13626,N_14837);
xor U16708 (N_16708,N_13416,N_14634);
nor U16709 (N_16709,N_13527,N_13890);
nor U16710 (N_16710,N_13941,N_13237);
xor U16711 (N_16711,N_13252,N_13012);
nand U16712 (N_16712,N_12612,N_14451);
or U16713 (N_16713,N_14350,N_14094);
xnor U16714 (N_16714,N_13277,N_12270);
or U16715 (N_16715,N_12669,N_13486);
or U16716 (N_16716,N_12207,N_12632);
nor U16717 (N_16717,N_13697,N_12330);
xor U16718 (N_16718,N_13595,N_13592);
or U16719 (N_16719,N_14315,N_14365);
xor U16720 (N_16720,N_14814,N_14460);
and U16721 (N_16721,N_13330,N_12550);
and U16722 (N_16722,N_12735,N_14480);
nor U16723 (N_16723,N_12253,N_13037);
xnor U16724 (N_16724,N_12505,N_12543);
xnor U16725 (N_16725,N_13236,N_12036);
nand U16726 (N_16726,N_14416,N_13199);
or U16727 (N_16727,N_13539,N_14719);
xor U16728 (N_16728,N_12244,N_14302);
and U16729 (N_16729,N_14160,N_12579);
nand U16730 (N_16730,N_12802,N_14509);
and U16731 (N_16731,N_14455,N_14488);
nand U16732 (N_16732,N_13194,N_12316);
xor U16733 (N_16733,N_13103,N_14790);
and U16734 (N_16734,N_14504,N_12184);
nor U16735 (N_16735,N_14005,N_12945);
nand U16736 (N_16736,N_12105,N_12872);
or U16737 (N_16737,N_14341,N_13526);
nand U16738 (N_16738,N_12328,N_12052);
and U16739 (N_16739,N_13581,N_13520);
and U16740 (N_16740,N_13264,N_12414);
and U16741 (N_16741,N_12418,N_13027);
or U16742 (N_16742,N_13414,N_12722);
and U16743 (N_16743,N_12838,N_12541);
nor U16744 (N_16744,N_12745,N_13064);
or U16745 (N_16745,N_12652,N_13431);
and U16746 (N_16746,N_12611,N_12606);
xnor U16747 (N_16747,N_12206,N_12211);
nor U16748 (N_16748,N_14528,N_13954);
nor U16749 (N_16749,N_13867,N_13829);
nor U16750 (N_16750,N_12401,N_14699);
nand U16751 (N_16751,N_13513,N_13500);
nor U16752 (N_16752,N_12524,N_13343);
and U16753 (N_16753,N_13911,N_14659);
nand U16754 (N_16754,N_12815,N_14414);
or U16755 (N_16755,N_13450,N_12445);
nand U16756 (N_16756,N_14907,N_12144);
nand U16757 (N_16757,N_14664,N_14086);
and U16758 (N_16758,N_14109,N_12631);
nand U16759 (N_16759,N_13284,N_14687);
or U16760 (N_16760,N_14434,N_14107);
xor U16761 (N_16761,N_14016,N_13697);
or U16762 (N_16762,N_14613,N_12750);
nand U16763 (N_16763,N_14663,N_12240);
or U16764 (N_16764,N_14389,N_13750);
or U16765 (N_16765,N_14194,N_14445);
nand U16766 (N_16766,N_14423,N_12767);
and U16767 (N_16767,N_13417,N_14009);
nand U16768 (N_16768,N_13862,N_13900);
xor U16769 (N_16769,N_14408,N_13134);
nor U16770 (N_16770,N_13778,N_14205);
and U16771 (N_16771,N_12239,N_12679);
nand U16772 (N_16772,N_13067,N_14709);
xor U16773 (N_16773,N_13439,N_14921);
nor U16774 (N_16774,N_12062,N_12738);
or U16775 (N_16775,N_12409,N_14804);
nor U16776 (N_16776,N_12926,N_14376);
and U16777 (N_16777,N_12898,N_14217);
nand U16778 (N_16778,N_14042,N_12213);
and U16779 (N_16779,N_13007,N_12021);
nor U16780 (N_16780,N_13462,N_13443);
or U16781 (N_16781,N_12089,N_13160);
nor U16782 (N_16782,N_13363,N_12364);
nand U16783 (N_16783,N_13798,N_12349);
nor U16784 (N_16784,N_12304,N_12395);
nor U16785 (N_16785,N_12281,N_13087);
nor U16786 (N_16786,N_13126,N_14446);
xnor U16787 (N_16787,N_13138,N_12918);
nand U16788 (N_16788,N_14833,N_12411);
and U16789 (N_16789,N_14188,N_13766);
nand U16790 (N_16790,N_14294,N_12427);
or U16791 (N_16791,N_13231,N_13814);
and U16792 (N_16792,N_12589,N_13915);
and U16793 (N_16793,N_13349,N_12575);
xor U16794 (N_16794,N_14567,N_14246);
or U16795 (N_16795,N_14838,N_12211);
or U16796 (N_16796,N_14270,N_12911);
and U16797 (N_16797,N_12154,N_13335);
xor U16798 (N_16798,N_13664,N_14218);
xor U16799 (N_16799,N_13315,N_12403);
xor U16800 (N_16800,N_14208,N_14127);
nand U16801 (N_16801,N_14226,N_13961);
or U16802 (N_16802,N_13565,N_14874);
nand U16803 (N_16803,N_13756,N_12225);
nand U16804 (N_16804,N_14049,N_12937);
xor U16805 (N_16805,N_12051,N_12061);
nand U16806 (N_16806,N_12354,N_13695);
nor U16807 (N_16807,N_14564,N_14288);
nand U16808 (N_16808,N_13421,N_14625);
nor U16809 (N_16809,N_14051,N_14758);
xnor U16810 (N_16810,N_14928,N_14191);
xor U16811 (N_16811,N_14697,N_12074);
or U16812 (N_16812,N_12391,N_14496);
xnor U16813 (N_16813,N_12458,N_12206);
nand U16814 (N_16814,N_14579,N_14715);
nand U16815 (N_16815,N_12643,N_14680);
nor U16816 (N_16816,N_14582,N_13600);
nand U16817 (N_16817,N_12872,N_13810);
xor U16818 (N_16818,N_14119,N_13812);
nand U16819 (N_16819,N_14347,N_13050);
and U16820 (N_16820,N_12250,N_12172);
nand U16821 (N_16821,N_13122,N_12005);
nor U16822 (N_16822,N_13798,N_14927);
nand U16823 (N_16823,N_12845,N_13516);
or U16824 (N_16824,N_13130,N_12610);
or U16825 (N_16825,N_13500,N_13265);
nor U16826 (N_16826,N_13772,N_14332);
xor U16827 (N_16827,N_14089,N_14324);
or U16828 (N_16828,N_14233,N_13743);
or U16829 (N_16829,N_14856,N_14913);
nor U16830 (N_16830,N_13618,N_13177);
or U16831 (N_16831,N_14204,N_12604);
or U16832 (N_16832,N_12071,N_12556);
nor U16833 (N_16833,N_12951,N_12993);
and U16834 (N_16834,N_13041,N_14245);
nor U16835 (N_16835,N_12443,N_12053);
or U16836 (N_16836,N_12681,N_14576);
nand U16837 (N_16837,N_14436,N_13063);
nand U16838 (N_16838,N_12954,N_13444);
nor U16839 (N_16839,N_14824,N_12539);
nor U16840 (N_16840,N_12709,N_14983);
nand U16841 (N_16841,N_13517,N_13683);
and U16842 (N_16842,N_12284,N_12983);
nor U16843 (N_16843,N_14772,N_13693);
xor U16844 (N_16844,N_13695,N_13991);
and U16845 (N_16845,N_13078,N_12080);
nor U16846 (N_16846,N_14101,N_14726);
nor U16847 (N_16847,N_13381,N_13700);
nand U16848 (N_16848,N_13689,N_14474);
nor U16849 (N_16849,N_14711,N_14137);
and U16850 (N_16850,N_13184,N_13120);
nand U16851 (N_16851,N_13357,N_14995);
nor U16852 (N_16852,N_13668,N_12812);
nor U16853 (N_16853,N_13782,N_14376);
nor U16854 (N_16854,N_13630,N_13824);
nor U16855 (N_16855,N_12815,N_13438);
nand U16856 (N_16856,N_14630,N_12756);
and U16857 (N_16857,N_14876,N_13780);
nand U16858 (N_16858,N_14107,N_14761);
xor U16859 (N_16859,N_12365,N_13091);
nand U16860 (N_16860,N_13092,N_12487);
xor U16861 (N_16861,N_14691,N_13039);
nor U16862 (N_16862,N_13126,N_12356);
nand U16863 (N_16863,N_13594,N_13454);
and U16864 (N_16864,N_13511,N_13402);
and U16865 (N_16865,N_14228,N_12563);
xnor U16866 (N_16866,N_12153,N_14016);
and U16867 (N_16867,N_13076,N_14831);
nand U16868 (N_16868,N_13485,N_13830);
and U16869 (N_16869,N_12156,N_13342);
or U16870 (N_16870,N_14734,N_12367);
nand U16871 (N_16871,N_13732,N_14563);
xor U16872 (N_16872,N_13285,N_14036);
and U16873 (N_16873,N_14287,N_12856);
or U16874 (N_16874,N_12666,N_14023);
and U16875 (N_16875,N_14040,N_13722);
and U16876 (N_16876,N_14331,N_12100);
nor U16877 (N_16877,N_13823,N_14850);
nor U16878 (N_16878,N_13323,N_14087);
and U16879 (N_16879,N_14753,N_13218);
and U16880 (N_16880,N_14139,N_14171);
or U16881 (N_16881,N_14390,N_12295);
nand U16882 (N_16882,N_13664,N_12530);
or U16883 (N_16883,N_12780,N_14867);
and U16884 (N_16884,N_13543,N_14768);
nand U16885 (N_16885,N_14743,N_12801);
and U16886 (N_16886,N_14225,N_14390);
nor U16887 (N_16887,N_13085,N_13819);
nand U16888 (N_16888,N_14048,N_14712);
and U16889 (N_16889,N_14971,N_12043);
or U16890 (N_16890,N_12042,N_13461);
and U16891 (N_16891,N_14794,N_12078);
and U16892 (N_16892,N_12116,N_12658);
xor U16893 (N_16893,N_14068,N_13173);
nand U16894 (N_16894,N_12757,N_13033);
and U16895 (N_16895,N_12776,N_12911);
nand U16896 (N_16896,N_14957,N_13535);
and U16897 (N_16897,N_14754,N_12614);
nand U16898 (N_16898,N_13437,N_14155);
nor U16899 (N_16899,N_14302,N_14358);
nor U16900 (N_16900,N_13967,N_14820);
nor U16901 (N_16901,N_13363,N_14360);
nand U16902 (N_16902,N_13043,N_14838);
and U16903 (N_16903,N_13505,N_14106);
xor U16904 (N_16904,N_14951,N_13738);
and U16905 (N_16905,N_12518,N_13307);
nand U16906 (N_16906,N_14151,N_13453);
and U16907 (N_16907,N_12106,N_14225);
and U16908 (N_16908,N_13049,N_12496);
or U16909 (N_16909,N_13416,N_13215);
and U16910 (N_16910,N_13018,N_14157);
nand U16911 (N_16911,N_12865,N_13035);
or U16912 (N_16912,N_14454,N_13485);
xnor U16913 (N_16913,N_12592,N_13391);
and U16914 (N_16914,N_13237,N_12788);
or U16915 (N_16915,N_12045,N_13318);
or U16916 (N_16916,N_13536,N_14143);
nand U16917 (N_16917,N_12772,N_13209);
or U16918 (N_16918,N_12288,N_14557);
nand U16919 (N_16919,N_13752,N_14122);
xnor U16920 (N_16920,N_13716,N_12456);
or U16921 (N_16921,N_12215,N_13478);
xor U16922 (N_16922,N_14663,N_14794);
nor U16923 (N_16923,N_13808,N_13174);
xor U16924 (N_16924,N_12383,N_13463);
xnor U16925 (N_16925,N_13746,N_13119);
and U16926 (N_16926,N_13018,N_13748);
or U16927 (N_16927,N_13541,N_13113);
or U16928 (N_16928,N_14412,N_13321);
or U16929 (N_16929,N_14236,N_12536);
nand U16930 (N_16930,N_14710,N_12262);
nor U16931 (N_16931,N_14521,N_12409);
and U16932 (N_16932,N_12558,N_12780);
nor U16933 (N_16933,N_14522,N_14806);
or U16934 (N_16934,N_13872,N_13538);
and U16935 (N_16935,N_12829,N_12871);
or U16936 (N_16936,N_14801,N_13731);
nor U16937 (N_16937,N_13237,N_12547);
nor U16938 (N_16938,N_14666,N_13423);
nand U16939 (N_16939,N_13667,N_13811);
nor U16940 (N_16940,N_14784,N_12700);
xor U16941 (N_16941,N_12325,N_12475);
and U16942 (N_16942,N_12744,N_14397);
xor U16943 (N_16943,N_12118,N_12195);
nor U16944 (N_16944,N_13609,N_14659);
or U16945 (N_16945,N_12855,N_13107);
nor U16946 (N_16946,N_14858,N_13080);
nor U16947 (N_16947,N_12001,N_12209);
and U16948 (N_16948,N_12869,N_12248);
or U16949 (N_16949,N_14994,N_14871);
nor U16950 (N_16950,N_13671,N_12866);
nor U16951 (N_16951,N_12293,N_14767);
or U16952 (N_16952,N_12100,N_13166);
or U16953 (N_16953,N_14792,N_14712);
or U16954 (N_16954,N_13989,N_13467);
nand U16955 (N_16955,N_13752,N_14082);
or U16956 (N_16956,N_13643,N_14810);
nand U16957 (N_16957,N_12654,N_14842);
xor U16958 (N_16958,N_13388,N_13242);
and U16959 (N_16959,N_12647,N_12708);
nand U16960 (N_16960,N_12877,N_13080);
or U16961 (N_16961,N_12268,N_13704);
nor U16962 (N_16962,N_12826,N_12999);
xor U16963 (N_16963,N_14141,N_13085);
or U16964 (N_16964,N_12960,N_13982);
nor U16965 (N_16965,N_13450,N_13598);
or U16966 (N_16966,N_14331,N_14644);
nand U16967 (N_16967,N_14874,N_14830);
and U16968 (N_16968,N_13249,N_12032);
nor U16969 (N_16969,N_12082,N_12216);
nand U16970 (N_16970,N_12324,N_14841);
xor U16971 (N_16971,N_13075,N_13936);
nor U16972 (N_16972,N_13972,N_13652);
nor U16973 (N_16973,N_14830,N_13206);
and U16974 (N_16974,N_13397,N_12616);
or U16975 (N_16975,N_14867,N_13830);
and U16976 (N_16976,N_14472,N_13272);
nand U16977 (N_16977,N_14767,N_13255);
and U16978 (N_16978,N_12795,N_14978);
or U16979 (N_16979,N_12690,N_13573);
nor U16980 (N_16980,N_14569,N_14716);
nand U16981 (N_16981,N_12391,N_14849);
and U16982 (N_16982,N_14245,N_12875);
nand U16983 (N_16983,N_12011,N_12465);
nor U16984 (N_16984,N_12221,N_14034);
or U16985 (N_16985,N_14382,N_13825);
or U16986 (N_16986,N_14133,N_13465);
and U16987 (N_16987,N_12833,N_14237);
nor U16988 (N_16988,N_13245,N_14362);
xnor U16989 (N_16989,N_13660,N_14683);
nand U16990 (N_16990,N_12916,N_14816);
xnor U16991 (N_16991,N_14994,N_13201);
or U16992 (N_16992,N_13353,N_12361);
nand U16993 (N_16993,N_14378,N_13783);
or U16994 (N_16994,N_13204,N_12159);
and U16995 (N_16995,N_13969,N_12841);
nand U16996 (N_16996,N_13605,N_13254);
and U16997 (N_16997,N_13404,N_13822);
nor U16998 (N_16998,N_12385,N_13655);
or U16999 (N_16999,N_13668,N_13263);
nand U17000 (N_17000,N_13931,N_14441);
xor U17001 (N_17001,N_12621,N_14093);
and U17002 (N_17002,N_14082,N_12183);
nor U17003 (N_17003,N_13326,N_14360);
nor U17004 (N_17004,N_12894,N_13555);
or U17005 (N_17005,N_14294,N_12284);
or U17006 (N_17006,N_14725,N_12431);
xnor U17007 (N_17007,N_12208,N_12548);
and U17008 (N_17008,N_13797,N_13511);
nor U17009 (N_17009,N_13422,N_13438);
nand U17010 (N_17010,N_13999,N_12799);
nor U17011 (N_17011,N_13096,N_13919);
xnor U17012 (N_17012,N_13220,N_14814);
or U17013 (N_17013,N_12307,N_13393);
nor U17014 (N_17014,N_13173,N_12969);
xor U17015 (N_17015,N_14336,N_14834);
or U17016 (N_17016,N_12585,N_12928);
nor U17017 (N_17017,N_14878,N_14731);
nand U17018 (N_17018,N_14526,N_14000);
xor U17019 (N_17019,N_13282,N_12599);
xnor U17020 (N_17020,N_13231,N_12350);
or U17021 (N_17021,N_12887,N_12763);
or U17022 (N_17022,N_13847,N_12960);
nand U17023 (N_17023,N_13651,N_14763);
and U17024 (N_17024,N_14228,N_12666);
xor U17025 (N_17025,N_13204,N_14724);
xnor U17026 (N_17026,N_13249,N_12970);
xor U17027 (N_17027,N_12576,N_14776);
and U17028 (N_17028,N_14897,N_14209);
nand U17029 (N_17029,N_14502,N_12455);
or U17030 (N_17030,N_13064,N_12943);
or U17031 (N_17031,N_14454,N_13126);
nand U17032 (N_17032,N_13213,N_14469);
and U17033 (N_17033,N_14678,N_14896);
or U17034 (N_17034,N_12997,N_12150);
nor U17035 (N_17035,N_13721,N_12272);
and U17036 (N_17036,N_12039,N_13117);
nor U17037 (N_17037,N_12787,N_13325);
nand U17038 (N_17038,N_14913,N_14873);
or U17039 (N_17039,N_14943,N_14241);
and U17040 (N_17040,N_12311,N_14395);
and U17041 (N_17041,N_14424,N_12290);
nand U17042 (N_17042,N_14539,N_13278);
nor U17043 (N_17043,N_12547,N_13856);
xnor U17044 (N_17044,N_12107,N_13117);
or U17045 (N_17045,N_14844,N_13299);
xnor U17046 (N_17046,N_13421,N_13457);
nor U17047 (N_17047,N_14174,N_13232);
xnor U17048 (N_17048,N_12167,N_13516);
nor U17049 (N_17049,N_13816,N_14476);
xor U17050 (N_17050,N_14719,N_13354);
xor U17051 (N_17051,N_13980,N_13847);
xnor U17052 (N_17052,N_13376,N_14592);
xor U17053 (N_17053,N_14536,N_13673);
nand U17054 (N_17054,N_13025,N_14705);
and U17055 (N_17055,N_14422,N_12643);
and U17056 (N_17056,N_13530,N_13508);
nand U17057 (N_17057,N_12926,N_14739);
nor U17058 (N_17058,N_13745,N_13543);
and U17059 (N_17059,N_14015,N_13089);
nor U17060 (N_17060,N_13707,N_14308);
nand U17061 (N_17061,N_12057,N_14402);
or U17062 (N_17062,N_14957,N_14146);
xnor U17063 (N_17063,N_13184,N_13791);
xnor U17064 (N_17064,N_13310,N_13278);
or U17065 (N_17065,N_12226,N_12865);
or U17066 (N_17066,N_13063,N_14172);
nand U17067 (N_17067,N_12741,N_12259);
nand U17068 (N_17068,N_13336,N_14927);
nand U17069 (N_17069,N_12321,N_12822);
or U17070 (N_17070,N_14216,N_13850);
xnor U17071 (N_17071,N_14931,N_14704);
xnor U17072 (N_17072,N_13048,N_13822);
nor U17073 (N_17073,N_14704,N_12469);
nand U17074 (N_17074,N_12106,N_14103);
and U17075 (N_17075,N_14429,N_14079);
xor U17076 (N_17076,N_12272,N_14414);
or U17077 (N_17077,N_12949,N_12040);
and U17078 (N_17078,N_14946,N_14489);
or U17079 (N_17079,N_12201,N_14436);
nand U17080 (N_17080,N_12398,N_13888);
and U17081 (N_17081,N_12868,N_13736);
xnor U17082 (N_17082,N_13862,N_12473);
nor U17083 (N_17083,N_12460,N_13578);
or U17084 (N_17084,N_13120,N_12432);
or U17085 (N_17085,N_13331,N_12619);
nor U17086 (N_17086,N_14372,N_14284);
nor U17087 (N_17087,N_14423,N_14510);
xnor U17088 (N_17088,N_14871,N_12486);
or U17089 (N_17089,N_14019,N_12304);
xnor U17090 (N_17090,N_12452,N_12731);
nor U17091 (N_17091,N_12509,N_14326);
nand U17092 (N_17092,N_13169,N_13102);
nor U17093 (N_17093,N_13883,N_14730);
nor U17094 (N_17094,N_12550,N_14130);
nor U17095 (N_17095,N_13112,N_14317);
nor U17096 (N_17096,N_12376,N_14962);
xor U17097 (N_17097,N_13206,N_12014);
xnor U17098 (N_17098,N_14109,N_13989);
and U17099 (N_17099,N_12370,N_13685);
nor U17100 (N_17100,N_12455,N_14645);
nor U17101 (N_17101,N_12635,N_13641);
or U17102 (N_17102,N_13240,N_13636);
nor U17103 (N_17103,N_13771,N_12411);
and U17104 (N_17104,N_13740,N_14260);
and U17105 (N_17105,N_12585,N_13079);
nand U17106 (N_17106,N_13940,N_13963);
and U17107 (N_17107,N_12472,N_14415);
xnor U17108 (N_17108,N_14748,N_14137);
and U17109 (N_17109,N_12903,N_14307);
or U17110 (N_17110,N_13832,N_13508);
nand U17111 (N_17111,N_12038,N_13437);
nand U17112 (N_17112,N_13247,N_14204);
and U17113 (N_17113,N_13986,N_12823);
xnor U17114 (N_17114,N_14766,N_12446);
nor U17115 (N_17115,N_12113,N_14270);
and U17116 (N_17116,N_13326,N_12077);
nand U17117 (N_17117,N_14475,N_13883);
or U17118 (N_17118,N_13614,N_12648);
or U17119 (N_17119,N_14209,N_14891);
or U17120 (N_17120,N_12306,N_12620);
and U17121 (N_17121,N_12152,N_14652);
and U17122 (N_17122,N_13808,N_12375);
and U17123 (N_17123,N_14988,N_12697);
and U17124 (N_17124,N_13817,N_13658);
nor U17125 (N_17125,N_12893,N_14826);
nand U17126 (N_17126,N_14497,N_13027);
xor U17127 (N_17127,N_13276,N_12534);
nor U17128 (N_17128,N_12362,N_13578);
and U17129 (N_17129,N_14373,N_13173);
xnor U17130 (N_17130,N_13696,N_13015);
nor U17131 (N_17131,N_14517,N_13357);
and U17132 (N_17132,N_12513,N_14988);
xor U17133 (N_17133,N_12690,N_12314);
xor U17134 (N_17134,N_12216,N_13651);
nor U17135 (N_17135,N_13143,N_12907);
xor U17136 (N_17136,N_13403,N_13569);
xor U17137 (N_17137,N_13678,N_14983);
nor U17138 (N_17138,N_13474,N_14771);
and U17139 (N_17139,N_13500,N_14377);
nand U17140 (N_17140,N_13037,N_13015);
and U17141 (N_17141,N_14365,N_12012);
nand U17142 (N_17142,N_12212,N_14603);
nor U17143 (N_17143,N_14943,N_12567);
and U17144 (N_17144,N_13244,N_13267);
nor U17145 (N_17145,N_14527,N_12163);
xnor U17146 (N_17146,N_13931,N_14199);
xor U17147 (N_17147,N_12553,N_14001);
and U17148 (N_17148,N_14459,N_13036);
or U17149 (N_17149,N_12402,N_13429);
nand U17150 (N_17150,N_14555,N_14135);
xnor U17151 (N_17151,N_14471,N_14974);
and U17152 (N_17152,N_13149,N_14073);
xor U17153 (N_17153,N_14955,N_14186);
nor U17154 (N_17154,N_14385,N_13537);
or U17155 (N_17155,N_13208,N_12118);
or U17156 (N_17156,N_12382,N_13407);
and U17157 (N_17157,N_13834,N_12918);
and U17158 (N_17158,N_14111,N_13549);
or U17159 (N_17159,N_13484,N_13958);
and U17160 (N_17160,N_14247,N_13545);
nor U17161 (N_17161,N_14511,N_14336);
nand U17162 (N_17162,N_14952,N_12637);
xnor U17163 (N_17163,N_14758,N_13800);
xor U17164 (N_17164,N_13178,N_12208);
and U17165 (N_17165,N_13574,N_12328);
or U17166 (N_17166,N_13306,N_12155);
nand U17167 (N_17167,N_14797,N_13479);
xor U17168 (N_17168,N_13144,N_14218);
and U17169 (N_17169,N_12339,N_14441);
nor U17170 (N_17170,N_13996,N_13185);
and U17171 (N_17171,N_12957,N_12237);
and U17172 (N_17172,N_12390,N_13682);
nor U17173 (N_17173,N_14512,N_13900);
or U17174 (N_17174,N_13538,N_13186);
nor U17175 (N_17175,N_12244,N_13949);
and U17176 (N_17176,N_14485,N_13506);
xor U17177 (N_17177,N_14133,N_14583);
or U17178 (N_17178,N_13382,N_12486);
and U17179 (N_17179,N_12571,N_14796);
or U17180 (N_17180,N_13630,N_14029);
xor U17181 (N_17181,N_13933,N_12237);
or U17182 (N_17182,N_14096,N_12288);
nor U17183 (N_17183,N_14477,N_12837);
nand U17184 (N_17184,N_13224,N_12424);
nand U17185 (N_17185,N_14419,N_12834);
xor U17186 (N_17186,N_13689,N_13091);
nand U17187 (N_17187,N_13085,N_14182);
nor U17188 (N_17188,N_14421,N_12145);
or U17189 (N_17189,N_12100,N_14151);
and U17190 (N_17190,N_13772,N_14534);
nand U17191 (N_17191,N_14012,N_14513);
nand U17192 (N_17192,N_14323,N_12585);
and U17193 (N_17193,N_14052,N_14782);
nand U17194 (N_17194,N_12988,N_14653);
and U17195 (N_17195,N_12873,N_14482);
and U17196 (N_17196,N_12919,N_14023);
and U17197 (N_17197,N_13244,N_12959);
nor U17198 (N_17198,N_12302,N_12280);
or U17199 (N_17199,N_14852,N_14076);
and U17200 (N_17200,N_13526,N_13816);
xnor U17201 (N_17201,N_13029,N_13108);
nor U17202 (N_17202,N_14031,N_14463);
nor U17203 (N_17203,N_12374,N_13290);
xor U17204 (N_17204,N_13056,N_12732);
nor U17205 (N_17205,N_12207,N_12794);
xor U17206 (N_17206,N_13349,N_12456);
nor U17207 (N_17207,N_12925,N_13394);
nor U17208 (N_17208,N_13163,N_14290);
or U17209 (N_17209,N_12279,N_14094);
or U17210 (N_17210,N_12162,N_13729);
or U17211 (N_17211,N_13955,N_12186);
nor U17212 (N_17212,N_12903,N_13955);
or U17213 (N_17213,N_12099,N_13172);
xnor U17214 (N_17214,N_12031,N_12958);
nand U17215 (N_17215,N_14905,N_13255);
nand U17216 (N_17216,N_13516,N_14565);
xnor U17217 (N_17217,N_12469,N_12152);
xnor U17218 (N_17218,N_14184,N_13002);
nand U17219 (N_17219,N_12517,N_12059);
and U17220 (N_17220,N_12215,N_13743);
xnor U17221 (N_17221,N_14267,N_14248);
or U17222 (N_17222,N_12279,N_13993);
xor U17223 (N_17223,N_13199,N_12278);
xor U17224 (N_17224,N_14172,N_13965);
nand U17225 (N_17225,N_13625,N_14875);
nor U17226 (N_17226,N_12428,N_12337);
xnor U17227 (N_17227,N_12312,N_14875);
nand U17228 (N_17228,N_14539,N_14131);
and U17229 (N_17229,N_13997,N_12110);
or U17230 (N_17230,N_13840,N_14854);
or U17231 (N_17231,N_12375,N_12341);
nand U17232 (N_17232,N_12513,N_13886);
xor U17233 (N_17233,N_12563,N_12905);
or U17234 (N_17234,N_14927,N_14893);
or U17235 (N_17235,N_13913,N_13933);
nor U17236 (N_17236,N_14644,N_13785);
nand U17237 (N_17237,N_13369,N_13315);
nor U17238 (N_17238,N_14282,N_12509);
or U17239 (N_17239,N_14581,N_12386);
or U17240 (N_17240,N_13452,N_13236);
or U17241 (N_17241,N_12758,N_14358);
nand U17242 (N_17242,N_14450,N_13172);
xor U17243 (N_17243,N_13735,N_12829);
or U17244 (N_17244,N_14144,N_12000);
nor U17245 (N_17245,N_14279,N_14562);
xnor U17246 (N_17246,N_14199,N_13496);
or U17247 (N_17247,N_14047,N_13787);
xnor U17248 (N_17248,N_14121,N_14661);
nor U17249 (N_17249,N_14237,N_13316);
nor U17250 (N_17250,N_14986,N_12968);
xor U17251 (N_17251,N_12216,N_12622);
nor U17252 (N_17252,N_13678,N_13025);
and U17253 (N_17253,N_14126,N_13323);
or U17254 (N_17254,N_14179,N_14910);
xor U17255 (N_17255,N_12019,N_13203);
or U17256 (N_17256,N_14292,N_13001);
nor U17257 (N_17257,N_14831,N_14143);
nor U17258 (N_17258,N_12945,N_14276);
nand U17259 (N_17259,N_13074,N_12206);
or U17260 (N_17260,N_12593,N_14619);
and U17261 (N_17261,N_13900,N_13359);
nand U17262 (N_17262,N_12466,N_13127);
and U17263 (N_17263,N_14330,N_13373);
nand U17264 (N_17264,N_14359,N_13409);
nor U17265 (N_17265,N_14250,N_14160);
or U17266 (N_17266,N_14363,N_13721);
or U17267 (N_17267,N_12704,N_12486);
and U17268 (N_17268,N_13846,N_13248);
nand U17269 (N_17269,N_12064,N_12688);
and U17270 (N_17270,N_13383,N_12510);
or U17271 (N_17271,N_12854,N_12600);
nand U17272 (N_17272,N_12804,N_14212);
xnor U17273 (N_17273,N_13938,N_13760);
nand U17274 (N_17274,N_14924,N_13806);
or U17275 (N_17275,N_13709,N_13253);
or U17276 (N_17276,N_13643,N_12954);
and U17277 (N_17277,N_13122,N_13280);
or U17278 (N_17278,N_12355,N_14331);
nand U17279 (N_17279,N_12768,N_13740);
nand U17280 (N_17280,N_13296,N_14716);
or U17281 (N_17281,N_13199,N_13354);
nand U17282 (N_17282,N_14745,N_14475);
nand U17283 (N_17283,N_13917,N_12792);
or U17284 (N_17284,N_13633,N_13653);
xor U17285 (N_17285,N_12855,N_14846);
nor U17286 (N_17286,N_14555,N_13535);
or U17287 (N_17287,N_14897,N_14821);
nor U17288 (N_17288,N_12225,N_12495);
and U17289 (N_17289,N_14765,N_12569);
nor U17290 (N_17290,N_14349,N_14635);
and U17291 (N_17291,N_12163,N_13180);
nand U17292 (N_17292,N_12371,N_12417);
nor U17293 (N_17293,N_13025,N_14569);
nand U17294 (N_17294,N_13751,N_14231);
or U17295 (N_17295,N_13610,N_14399);
xnor U17296 (N_17296,N_14649,N_14923);
nor U17297 (N_17297,N_13386,N_13658);
nand U17298 (N_17298,N_13318,N_14571);
nor U17299 (N_17299,N_13714,N_12206);
and U17300 (N_17300,N_13770,N_13132);
xnor U17301 (N_17301,N_13567,N_14798);
nor U17302 (N_17302,N_13443,N_12710);
nand U17303 (N_17303,N_12361,N_12620);
nand U17304 (N_17304,N_12415,N_13416);
xnor U17305 (N_17305,N_13975,N_13279);
nor U17306 (N_17306,N_14673,N_12208);
xor U17307 (N_17307,N_12702,N_13617);
nor U17308 (N_17308,N_14024,N_14440);
nand U17309 (N_17309,N_13052,N_14210);
nand U17310 (N_17310,N_13101,N_13383);
or U17311 (N_17311,N_13826,N_12449);
and U17312 (N_17312,N_12995,N_13073);
or U17313 (N_17313,N_13343,N_12430);
nand U17314 (N_17314,N_12129,N_13490);
nand U17315 (N_17315,N_14862,N_12561);
xnor U17316 (N_17316,N_13342,N_14079);
or U17317 (N_17317,N_12316,N_14668);
nor U17318 (N_17318,N_12013,N_13077);
xnor U17319 (N_17319,N_13884,N_13513);
nor U17320 (N_17320,N_12726,N_12345);
and U17321 (N_17321,N_12794,N_12610);
nor U17322 (N_17322,N_14927,N_12521);
nor U17323 (N_17323,N_13869,N_13580);
xnor U17324 (N_17324,N_12316,N_12462);
or U17325 (N_17325,N_12841,N_12059);
and U17326 (N_17326,N_13110,N_13092);
xor U17327 (N_17327,N_12830,N_14249);
xor U17328 (N_17328,N_14274,N_13855);
and U17329 (N_17329,N_12162,N_12910);
nand U17330 (N_17330,N_12605,N_13310);
and U17331 (N_17331,N_13535,N_14656);
nand U17332 (N_17332,N_13418,N_13875);
xnor U17333 (N_17333,N_12405,N_12099);
xor U17334 (N_17334,N_14318,N_12621);
and U17335 (N_17335,N_14666,N_12967);
nor U17336 (N_17336,N_13460,N_14904);
or U17337 (N_17337,N_12139,N_12979);
nor U17338 (N_17338,N_13481,N_13998);
xor U17339 (N_17339,N_14521,N_14414);
nor U17340 (N_17340,N_13666,N_13446);
or U17341 (N_17341,N_14520,N_13871);
and U17342 (N_17342,N_14003,N_14956);
nand U17343 (N_17343,N_14349,N_12900);
or U17344 (N_17344,N_12431,N_14844);
and U17345 (N_17345,N_12003,N_13760);
nand U17346 (N_17346,N_13856,N_14642);
xor U17347 (N_17347,N_13202,N_14672);
and U17348 (N_17348,N_13483,N_13503);
and U17349 (N_17349,N_14213,N_12608);
nand U17350 (N_17350,N_12023,N_13894);
or U17351 (N_17351,N_13564,N_12508);
nand U17352 (N_17352,N_12739,N_14832);
nor U17353 (N_17353,N_14842,N_14717);
or U17354 (N_17354,N_13140,N_14323);
nand U17355 (N_17355,N_13708,N_13190);
and U17356 (N_17356,N_12010,N_14896);
nand U17357 (N_17357,N_13756,N_14862);
nor U17358 (N_17358,N_13039,N_14267);
and U17359 (N_17359,N_14797,N_13889);
or U17360 (N_17360,N_12854,N_14336);
or U17361 (N_17361,N_13236,N_13434);
nor U17362 (N_17362,N_14611,N_13326);
xor U17363 (N_17363,N_12796,N_13277);
nor U17364 (N_17364,N_14158,N_13034);
or U17365 (N_17365,N_13017,N_14187);
xnor U17366 (N_17366,N_14072,N_14410);
xnor U17367 (N_17367,N_12055,N_13674);
and U17368 (N_17368,N_12859,N_14718);
nand U17369 (N_17369,N_14913,N_13417);
nand U17370 (N_17370,N_12717,N_13982);
and U17371 (N_17371,N_14075,N_14723);
or U17372 (N_17372,N_12931,N_12605);
xnor U17373 (N_17373,N_13328,N_12678);
xor U17374 (N_17374,N_14842,N_13890);
xor U17375 (N_17375,N_12577,N_13538);
and U17376 (N_17376,N_12363,N_12521);
nor U17377 (N_17377,N_12997,N_14427);
and U17378 (N_17378,N_14213,N_12150);
or U17379 (N_17379,N_14987,N_12657);
xnor U17380 (N_17380,N_12333,N_12289);
nor U17381 (N_17381,N_13613,N_13650);
and U17382 (N_17382,N_13451,N_12958);
xor U17383 (N_17383,N_12712,N_14800);
nor U17384 (N_17384,N_14719,N_12128);
or U17385 (N_17385,N_12220,N_13091);
and U17386 (N_17386,N_13749,N_13477);
xnor U17387 (N_17387,N_13042,N_13600);
nand U17388 (N_17388,N_12699,N_12603);
xnor U17389 (N_17389,N_14795,N_12512);
xnor U17390 (N_17390,N_13098,N_13713);
nor U17391 (N_17391,N_14661,N_14122);
xor U17392 (N_17392,N_12193,N_12150);
nor U17393 (N_17393,N_13009,N_13039);
xnor U17394 (N_17394,N_14577,N_12848);
nor U17395 (N_17395,N_13678,N_13717);
nor U17396 (N_17396,N_12971,N_13494);
or U17397 (N_17397,N_12011,N_14579);
nor U17398 (N_17398,N_13168,N_14123);
nand U17399 (N_17399,N_13912,N_12278);
xnor U17400 (N_17400,N_13603,N_12058);
nand U17401 (N_17401,N_14371,N_14000);
xor U17402 (N_17402,N_12472,N_14236);
xnor U17403 (N_17403,N_13863,N_14173);
and U17404 (N_17404,N_12717,N_13367);
or U17405 (N_17405,N_14105,N_14872);
xnor U17406 (N_17406,N_14573,N_14271);
xor U17407 (N_17407,N_13498,N_12064);
xnor U17408 (N_17408,N_12465,N_14412);
xnor U17409 (N_17409,N_12718,N_12357);
nor U17410 (N_17410,N_13995,N_13380);
or U17411 (N_17411,N_13317,N_12105);
or U17412 (N_17412,N_12222,N_13090);
and U17413 (N_17413,N_13584,N_13490);
xnor U17414 (N_17414,N_14740,N_12866);
nor U17415 (N_17415,N_12521,N_14833);
nand U17416 (N_17416,N_12535,N_12132);
and U17417 (N_17417,N_14072,N_14899);
xor U17418 (N_17418,N_12638,N_13916);
xor U17419 (N_17419,N_14728,N_12053);
and U17420 (N_17420,N_14858,N_12601);
nand U17421 (N_17421,N_13369,N_14053);
nor U17422 (N_17422,N_13411,N_14649);
and U17423 (N_17423,N_12779,N_12419);
xor U17424 (N_17424,N_13995,N_14976);
or U17425 (N_17425,N_12230,N_14781);
xnor U17426 (N_17426,N_13263,N_12744);
and U17427 (N_17427,N_13608,N_12685);
nand U17428 (N_17428,N_13783,N_13065);
nor U17429 (N_17429,N_12829,N_12328);
xnor U17430 (N_17430,N_13383,N_14479);
xor U17431 (N_17431,N_12441,N_13057);
nand U17432 (N_17432,N_13325,N_12141);
xnor U17433 (N_17433,N_14651,N_12947);
nand U17434 (N_17434,N_12089,N_12046);
xor U17435 (N_17435,N_13753,N_14074);
and U17436 (N_17436,N_12710,N_14682);
or U17437 (N_17437,N_12679,N_13312);
nor U17438 (N_17438,N_13192,N_14367);
or U17439 (N_17439,N_12525,N_14014);
nand U17440 (N_17440,N_12637,N_13271);
or U17441 (N_17441,N_13863,N_13297);
or U17442 (N_17442,N_14139,N_14745);
xnor U17443 (N_17443,N_12245,N_12543);
and U17444 (N_17444,N_12217,N_14934);
and U17445 (N_17445,N_12430,N_13731);
and U17446 (N_17446,N_13784,N_13357);
and U17447 (N_17447,N_14990,N_12248);
nor U17448 (N_17448,N_14411,N_13416);
and U17449 (N_17449,N_13354,N_14933);
nor U17450 (N_17450,N_14562,N_14094);
and U17451 (N_17451,N_14999,N_13979);
nor U17452 (N_17452,N_14504,N_13425);
and U17453 (N_17453,N_13229,N_12722);
and U17454 (N_17454,N_13394,N_14573);
xnor U17455 (N_17455,N_14102,N_12744);
nor U17456 (N_17456,N_12013,N_12166);
nand U17457 (N_17457,N_14511,N_14460);
or U17458 (N_17458,N_14150,N_12779);
xnor U17459 (N_17459,N_13135,N_14635);
nor U17460 (N_17460,N_14885,N_12404);
and U17461 (N_17461,N_12780,N_14209);
or U17462 (N_17462,N_13760,N_14527);
nor U17463 (N_17463,N_12303,N_12473);
xor U17464 (N_17464,N_14498,N_14497);
nand U17465 (N_17465,N_12221,N_14567);
nor U17466 (N_17466,N_13129,N_12586);
and U17467 (N_17467,N_13305,N_14910);
xnor U17468 (N_17468,N_14705,N_14592);
nand U17469 (N_17469,N_14925,N_13825);
nand U17470 (N_17470,N_12798,N_12327);
xnor U17471 (N_17471,N_12826,N_13475);
nand U17472 (N_17472,N_13465,N_14807);
xnor U17473 (N_17473,N_12788,N_14408);
nand U17474 (N_17474,N_13725,N_12277);
xor U17475 (N_17475,N_14890,N_14823);
and U17476 (N_17476,N_12036,N_13290);
and U17477 (N_17477,N_14440,N_14140);
nand U17478 (N_17478,N_12693,N_12971);
nand U17479 (N_17479,N_13192,N_13662);
nor U17480 (N_17480,N_12887,N_13818);
nor U17481 (N_17481,N_13374,N_12466);
xnor U17482 (N_17482,N_13249,N_13062);
and U17483 (N_17483,N_12217,N_12285);
nor U17484 (N_17484,N_13698,N_13287);
nand U17485 (N_17485,N_13919,N_14557);
xor U17486 (N_17486,N_12787,N_13374);
xor U17487 (N_17487,N_14545,N_12958);
or U17488 (N_17488,N_12116,N_14197);
or U17489 (N_17489,N_14358,N_12878);
nor U17490 (N_17490,N_12408,N_12604);
or U17491 (N_17491,N_12958,N_13786);
nand U17492 (N_17492,N_13451,N_14025);
xnor U17493 (N_17493,N_12293,N_14689);
and U17494 (N_17494,N_12031,N_12369);
nor U17495 (N_17495,N_14236,N_14184);
xor U17496 (N_17496,N_14076,N_12957);
nand U17497 (N_17497,N_14341,N_12935);
nor U17498 (N_17498,N_14061,N_12956);
nor U17499 (N_17499,N_13541,N_13176);
nor U17500 (N_17500,N_12730,N_13335);
nand U17501 (N_17501,N_13537,N_12194);
nand U17502 (N_17502,N_13978,N_14736);
xor U17503 (N_17503,N_14858,N_14901);
nand U17504 (N_17504,N_14834,N_14673);
nand U17505 (N_17505,N_12338,N_13521);
nor U17506 (N_17506,N_12956,N_13003);
or U17507 (N_17507,N_13526,N_12924);
nor U17508 (N_17508,N_12256,N_13163);
or U17509 (N_17509,N_13105,N_12393);
nor U17510 (N_17510,N_14267,N_12145);
and U17511 (N_17511,N_14783,N_14532);
nor U17512 (N_17512,N_13086,N_13276);
xor U17513 (N_17513,N_12782,N_14757);
nor U17514 (N_17514,N_13377,N_13681);
nor U17515 (N_17515,N_12290,N_14205);
nor U17516 (N_17516,N_13937,N_14204);
and U17517 (N_17517,N_13808,N_13203);
xor U17518 (N_17518,N_14865,N_12835);
xor U17519 (N_17519,N_13445,N_14056);
xnor U17520 (N_17520,N_12362,N_12929);
and U17521 (N_17521,N_12200,N_14404);
or U17522 (N_17522,N_12259,N_14581);
or U17523 (N_17523,N_13780,N_14943);
xnor U17524 (N_17524,N_14493,N_13755);
and U17525 (N_17525,N_12867,N_13191);
nor U17526 (N_17526,N_12139,N_14441);
xnor U17527 (N_17527,N_14633,N_12348);
nand U17528 (N_17528,N_14826,N_13516);
or U17529 (N_17529,N_14739,N_13613);
or U17530 (N_17530,N_12836,N_12928);
and U17531 (N_17531,N_13207,N_14098);
xor U17532 (N_17532,N_13014,N_12601);
and U17533 (N_17533,N_12171,N_14245);
and U17534 (N_17534,N_14631,N_13068);
nor U17535 (N_17535,N_14801,N_13161);
or U17536 (N_17536,N_13664,N_12034);
nand U17537 (N_17537,N_14162,N_13500);
and U17538 (N_17538,N_14438,N_14548);
and U17539 (N_17539,N_12130,N_14638);
nor U17540 (N_17540,N_14652,N_14103);
nor U17541 (N_17541,N_14687,N_12797);
nand U17542 (N_17542,N_13850,N_14587);
and U17543 (N_17543,N_14923,N_13219);
or U17544 (N_17544,N_13523,N_13691);
nand U17545 (N_17545,N_14890,N_13116);
nand U17546 (N_17546,N_14774,N_13835);
nand U17547 (N_17547,N_13410,N_14385);
nor U17548 (N_17548,N_13049,N_12183);
or U17549 (N_17549,N_14806,N_12626);
xnor U17550 (N_17550,N_12740,N_14313);
or U17551 (N_17551,N_12281,N_12345);
and U17552 (N_17552,N_13596,N_14815);
xor U17553 (N_17553,N_12781,N_13142);
nor U17554 (N_17554,N_14983,N_14844);
nand U17555 (N_17555,N_13222,N_12554);
or U17556 (N_17556,N_13241,N_12624);
xnor U17557 (N_17557,N_13510,N_12499);
xor U17558 (N_17558,N_12222,N_13357);
or U17559 (N_17559,N_14959,N_14124);
and U17560 (N_17560,N_13091,N_12274);
and U17561 (N_17561,N_12052,N_14370);
nand U17562 (N_17562,N_12698,N_13412);
nor U17563 (N_17563,N_12656,N_14527);
nor U17564 (N_17564,N_12372,N_13353);
nand U17565 (N_17565,N_14410,N_13163);
or U17566 (N_17566,N_12296,N_12476);
nand U17567 (N_17567,N_12273,N_12165);
or U17568 (N_17568,N_14392,N_12087);
or U17569 (N_17569,N_14232,N_13914);
nor U17570 (N_17570,N_13362,N_12859);
and U17571 (N_17571,N_13750,N_14701);
nor U17572 (N_17572,N_14302,N_12885);
and U17573 (N_17573,N_14662,N_14624);
nor U17574 (N_17574,N_12107,N_13334);
nand U17575 (N_17575,N_13619,N_14826);
and U17576 (N_17576,N_14701,N_12109);
xor U17577 (N_17577,N_12717,N_13580);
nand U17578 (N_17578,N_14587,N_12963);
or U17579 (N_17579,N_14112,N_13275);
nand U17580 (N_17580,N_13594,N_14331);
and U17581 (N_17581,N_14971,N_14874);
nor U17582 (N_17582,N_13953,N_12090);
xnor U17583 (N_17583,N_13427,N_12048);
or U17584 (N_17584,N_14734,N_14291);
and U17585 (N_17585,N_13333,N_13566);
nand U17586 (N_17586,N_14604,N_14126);
or U17587 (N_17587,N_14176,N_13078);
nor U17588 (N_17588,N_12894,N_13562);
nand U17589 (N_17589,N_14521,N_12907);
nand U17590 (N_17590,N_12071,N_14614);
xnor U17591 (N_17591,N_12611,N_13422);
nand U17592 (N_17592,N_14611,N_12250);
or U17593 (N_17593,N_12331,N_13175);
xnor U17594 (N_17594,N_13651,N_14172);
xor U17595 (N_17595,N_12944,N_13797);
and U17596 (N_17596,N_12998,N_13104);
xor U17597 (N_17597,N_12334,N_13014);
xnor U17598 (N_17598,N_13532,N_12094);
nor U17599 (N_17599,N_13361,N_13619);
nand U17600 (N_17600,N_13466,N_14781);
nor U17601 (N_17601,N_13686,N_13415);
nand U17602 (N_17602,N_14884,N_12830);
xor U17603 (N_17603,N_12433,N_13276);
nor U17604 (N_17604,N_13128,N_13823);
nor U17605 (N_17605,N_13509,N_12878);
nand U17606 (N_17606,N_14008,N_12143);
xor U17607 (N_17607,N_13472,N_14297);
xnor U17608 (N_17608,N_12788,N_14347);
xor U17609 (N_17609,N_13363,N_14793);
nand U17610 (N_17610,N_14816,N_14939);
xnor U17611 (N_17611,N_14979,N_12045);
or U17612 (N_17612,N_12803,N_13317);
and U17613 (N_17613,N_13296,N_13183);
and U17614 (N_17614,N_13413,N_13542);
and U17615 (N_17615,N_12259,N_12015);
nand U17616 (N_17616,N_14369,N_13936);
xor U17617 (N_17617,N_13112,N_14063);
nor U17618 (N_17618,N_14762,N_13612);
or U17619 (N_17619,N_13185,N_14232);
nor U17620 (N_17620,N_14386,N_14174);
or U17621 (N_17621,N_13049,N_14228);
nand U17622 (N_17622,N_13591,N_13930);
and U17623 (N_17623,N_13086,N_13160);
nor U17624 (N_17624,N_14113,N_14341);
xor U17625 (N_17625,N_14025,N_12658);
and U17626 (N_17626,N_14405,N_14138);
nand U17627 (N_17627,N_14107,N_13304);
xnor U17628 (N_17628,N_12876,N_14458);
nand U17629 (N_17629,N_14760,N_13491);
xor U17630 (N_17630,N_13931,N_13892);
and U17631 (N_17631,N_13806,N_13101);
nor U17632 (N_17632,N_12196,N_13786);
or U17633 (N_17633,N_12780,N_12546);
nand U17634 (N_17634,N_13270,N_14075);
nand U17635 (N_17635,N_14173,N_14687);
and U17636 (N_17636,N_14305,N_12788);
nand U17637 (N_17637,N_12517,N_12087);
or U17638 (N_17638,N_14930,N_13950);
xnor U17639 (N_17639,N_14486,N_14516);
or U17640 (N_17640,N_12661,N_12886);
xnor U17641 (N_17641,N_14945,N_12060);
or U17642 (N_17642,N_13219,N_12939);
xor U17643 (N_17643,N_14895,N_12178);
and U17644 (N_17644,N_14918,N_13670);
nand U17645 (N_17645,N_13592,N_12903);
nand U17646 (N_17646,N_14868,N_12986);
nor U17647 (N_17647,N_12301,N_13292);
nand U17648 (N_17648,N_14656,N_14521);
and U17649 (N_17649,N_12110,N_14232);
xor U17650 (N_17650,N_13731,N_14950);
or U17651 (N_17651,N_14607,N_12492);
nand U17652 (N_17652,N_12552,N_12741);
nand U17653 (N_17653,N_13470,N_12813);
nor U17654 (N_17654,N_13910,N_13937);
nor U17655 (N_17655,N_12772,N_13116);
nor U17656 (N_17656,N_12988,N_12334);
xor U17657 (N_17657,N_13358,N_12032);
nand U17658 (N_17658,N_13393,N_14192);
nor U17659 (N_17659,N_12926,N_13083);
and U17660 (N_17660,N_14986,N_13890);
and U17661 (N_17661,N_12456,N_12667);
nand U17662 (N_17662,N_14320,N_14950);
xor U17663 (N_17663,N_13941,N_12385);
xnor U17664 (N_17664,N_14215,N_13102);
or U17665 (N_17665,N_13706,N_12697);
or U17666 (N_17666,N_14794,N_14902);
or U17667 (N_17667,N_14289,N_12209);
nand U17668 (N_17668,N_14868,N_13914);
nand U17669 (N_17669,N_12508,N_14600);
xor U17670 (N_17670,N_12761,N_12766);
nand U17671 (N_17671,N_12676,N_14149);
nor U17672 (N_17672,N_14235,N_12633);
xor U17673 (N_17673,N_13240,N_12904);
nand U17674 (N_17674,N_14289,N_14072);
xnor U17675 (N_17675,N_14348,N_13846);
and U17676 (N_17676,N_14494,N_14073);
and U17677 (N_17677,N_12612,N_14304);
xor U17678 (N_17678,N_12208,N_13083);
xnor U17679 (N_17679,N_12295,N_14486);
nand U17680 (N_17680,N_12986,N_13373);
and U17681 (N_17681,N_14561,N_14741);
xnor U17682 (N_17682,N_12333,N_12719);
nor U17683 (N_17683,N_12737,N_12147);
nor U17684 (N_17684,N_14812,N_12857);
or U17685 (N_17685,N_13057,N_13804);
nand U17686 (N_17686,N_12123,N_14816);
and U17687 (N_17687,N_13139,N_14988);
nor U17688 (N_17688,N_14016,N_14102);
or U17689 (N_17689,N_12289,N_12304);
nand U17690 (N_17690,N_12931,N_14867);
xnor U17691 (N_17691,N_12448,N_12638);
xnor U17692 (N_17692,N_14348,N_12979);
or U17693 (N_17693,N_13955,N_14834);
nor U17694 (N_17694,N_14356,N_14644);
xor U17695 (N_17695,N_12163,N_13186);
or U17696 (N_17696,N_13014,N_13098);
or U17697 (N_17697,N_13830,N_14611);
or U17698 (N_17698,N_13089,N_13683);
and U17699 (N_17699,N_13381,N_12014);
nor U17700 (N_17700,N_13220,N_12687);
nor U17701 (N_17701,N_14021,N_13324);
and U17702 (N_17702,N_13109,N_13166);
and U17703 (N_17703,N_12220,N_13007);
and U17704 (N_17704,N_12837,N_12597);
or U17705 (N_17705,N_14122,N_14882);
xnor U17706 (N_17706,N_13371,N_13432);
or U17707 (N_17707,N_12862,N_13160);
and U17708 (N_17708,N_13484,N_12858);
or U17709 (N_17709,N_13198,N_12720);
xor U17710 (N_17710,N_14122,N_12733);
or U17711 (N_17711,N_14649,N_12906);
nor U17712 (N_17712,N_12278,N_14093);
nand U17713 (N_17713,N_13377,N_14689);
or U17714 (N_17714,N_14046,N_14502);
nand U17715 (N_17715,N_13458,N_14491);
xor U17716 (N_17716,N_14971,N_14503);
nand U17717 (N_17717,N_12783,N_12323);
or U17718 (N_17718,N_14570,N_13680);
or U17719 (N_17719,N_14741,N_12350);
nor U17720 (N_17720,N_12130,N_12610);
nor U17721 (N_17721,N_12612,N_14612);
and U17722 (N_17722,N_14459,N_13475);
and U17723 (N_17723,N_12973,N_12668);
nand U17724 (N_17724,N_14353,N_14538);
nand U17725 (N_17725,N_13994,N_14586);
nor U17726 (N_17726,N_12208,N_13527);
and U17727 (N_17727,N_12959,N_12215);
and U17728 (N_17728,N_13713,N_14498);
and U17729 (N_17729,N_13359,N_14379);
xnor U17730 (N_17730,N_12435,N_13310);
nand U17731 (N_17731,N_12579,N_14436);
nand U17732 (N_17732,N_12157,N_13710);
nor U17733 (N_17733,N_14475,N_14387);
nor U17734 (N_17734,N_13370,N_13595);
nor U17735 (N_17735,N_14340,N_14421);
nor U17736 (N_17736,N_14553,N_14199);
xor U17737 (N_17737,N_13226,N_12959);
xnor U17738 (N_17738,N_13614,N_12834);
xor U17739 (N_17739,N_14064,N_13475);
xnor U17740 (N_17740,N_12112,N_12014);
xnor U17741 (N_17741,N_12122,N_14733);
or U17742 (N_17742,N_12837,N_12129);
nand U17743 (N_17743,N_13648,N_13569);
xnor U17744 (N_17744,N_14308,N_12586);
or U17745 (N_17745,N_14917,N_12835);
nor U17746 (N_17746,N_14743,N_14491);
or U17747 (N_17747,N_13901,N_14448);
nor U17748 (N_17748,N_12576,N_13518);
xor U17749 (N_17749,N_13511,N_12225);
nand U17750 (N_17750,N_14732,N_13727);
xor U17751 (N_17751,N_12546,N_14828);
nand U17752 (N_17752,N_12118,N_14204);
nand U17753 (N_17753,N_12715,N_12776);
or U17754 (N_17754,N_12428,N_13001);
nor U17755 (N_17755,N_13119,N_12394);
nor U17756 (N_17756,N_14109,N_12489);
and U17757 (N_17757,N_13488,N_12886);
and U17758 (N_17758,N_12834,N_12659);
nor U17759 (N_17759,N_13946,N_13413);
or U17760 (N_17760,N_13330,N_13019);
or U17761 (N_17761,N_12525,N_12409);
nor U17762 (N_17762,N_14453,N_12026);
and U17763 (N_17763,N_12850,N_13607);
nor U17764 (N_17764,N_14122,N_12392);
nor U17765 (N_17765,N_14210,N_12148);
and U17766 (N_17766,N_12921,N_13772);
nand U17767 (N_17767,N_13892,N_13089);
and U17768 (N_17768,N_14131,N_14931);
nor U17769 (N_17769,N_12584,N_12783);
nand U17770 (N_17770,N_12825,N_13683);
and U17771 (N_17771,N_13431,N_12570);
nor U17772 (N_17772,N_12100,N_13693);
and U17773 (N_17773,N_12919,N_13721);
and U17774 (N_17774,N_13246,N_12142);
nand U17775 (N_17775,N_14810,N_14945);
nor U17776 (N_17776,N_14655,N_14320);
nor U17777 (N_17777,N_14311,N_12164);
and U17778 (N_17778,N_14680,N_13436);
xnor U17779 (N_17779,N_12119,N_12272);
xnor U17780 (N_17780,N_14255,N_13567);
or U17781 (N_17781,N_13049,N_14186);
xnor U17782 (N_17782,N_13455,N_14733);
nor U17783 (N_17783,N_12844,N_13031);
or U17784 (N_17784,N_12210,N_13447);
nand U17785 (N_17785,N_13484,N_13583);
xor U17786 (N_17786,N_12861,N_13479);
nor U17787 (N_17787,N_13816,N_12636);
nand U17788 (N_17788,N_14199,N_14154);
and U17789 (N_17789,N_12986,N_13216);
and U17790 (N_17790,N_13112,N_12783);
nand U17791 (N_17791,N_13503,N_14994);
nor U17792 (N_17792,N_13392,N_14672);
nand U17793 (N_17793,N_13564,N_12101);
nand U17794 (N_17794,N_14243,N_12619);
or U17795 (N_17795,N_14957,N_13612);
and U17796 (N_17796,N_14275,N_12642);
nor U17797 (N_17797,N_12729,N_13446);
or U17798 (N_17798,N_12292,N_14422);
nand U17799 (N_17799,N_13216,N_13683);
xor U17800 (N_17800,N_14342,N_13038);
or U17801 (N_17801,N_14548,N_12886);
or U17802 (N_17802,N_13902,N_13627);
nor U17803 (N_17803,N_12067,N_12206);
nand U17804 (N_17804,N_13983,N_13904);
nand U17805 (N_17805,N_13211,N_13478);
and U17806 (N_17806,N_13128,N_12422);
and U17807 (N_17807,N_13383,N_13200);
nand U17808 (N_17808,N_12774,N_13834);
nor U17809 (N_17809,N_14269,N_14883);
nand U17810 (N_17810,N_14653,N_12542);
xnor U17811 (N_17811,N_12502,N_13209);
nor U17812 (N_17812,N_14105,N_12933);
or U17813 (N_17813,N_13859,N_12834);
and U17814 (N_17814,N_13705,N_13270);
nand U17815 (N_17815,N_13719,N_13471);
nand U17816 (N_17816,N_12180,N_13364);
and U17817 (N_17817,N_14921,N_14838);
nand U17818 (N_17818,N_12998,N_13174);
and U17819 (N_17819,N_13274,N_13961);
or U17820 (N_17820,N_12192,N_14926);
xor U17821 (N_17821,N_13495,N_13519);
xor U17822 (N_17822,N_13062,N_12886);
nand U17823 (N_17823,N_13696,N_12888);
xor U17824 (N_17824,N_13909,N_12988);
or U17825 (N_17825,N_13624,N_13580);
nor U17826 (N_17826,N_13738,N_12253);
xnor U17827 (N_17827,N_12988,N_13005);
xor U17828 (N_17828,N_13742,N_13725);
and U17829 (N_17829,N_12949,N_13803);
nor U17830 (N_17830,N_12117,N_13945);
and U17831 (N_17831,N_13358,N_12397);
xnor U17832 (N_17832,N_13586,N_13993);
and U17833 (N_17833,N_14558,N_12610);
or U17834 (N_17834,N_14383,N_14425);
nor U17835 (N_17835,N_14090,N_13998);
nor U17836 (N_17836,N_14031,N_13243);
and U17837 (N_17837,N_12724,N_13560);
or U17838 (N_17838,N_12527,N_13505);
nand U17839 (N_17839,N_13215,N_14211);
nor U17840 (N_17840,N_12259,N_12548);
or U17841 (N_17841,N_13157,N_12046);
and U17842 (N_17842,N_13245,N_13360);
and U17843 (N_17843,N_13178,N_12218);
and U17844 (N_17844,N_13449,N_14142);
nand U17845 (N_17845,N_13964,N_12759);
nand U17846 (N_17846,N_12496,N_14746);
nor U17847 (N_17847,N_13388,N_12241);
or U17848 (N_17848,N_14560,N_13882);
nor U17849 (N_17849,N_13016,N_13528);
nor U17850 (N_17850,N_14150,N_13264);
and U17851 (N_17851,N_14596,N_14268);
nand U17852 (N_17852,N_13266,N_12502);
or U17853 (N_17853,N_13800,N_13075);
or U17854 (N_17854,N_13413,N_14906);
or U17855 (N_17855,N_12419,N_13345);
and U17856 (N_17856,N_13019,N_13560);
nand U17857 (N_17857,N_14177,N_12669);
xor U17858 (N_17858,N_13734,N_14471);
xnor U17859 (N_17859,N_14853,N_14447);
xor U17860 (N_17860,N_14060,N_13420);
nand U17861 (N_17861,N_12433,N_13031);
nor U17862 (N_17862,N_14368,N_13010);
xor U17863 (N_17863,N_12776,N_13766);
nor U17864 (N_17864,N_14023,N_14483);
and U17865 (N_17865,N_12940,N_14420);
xor U17866 (N_17866,N_13232,N_14048);
xor U17867 (N_17867,N_12005,N_14295);
nand U17868 (N_17868,N_13657,N_13959);
or U17869 (N_17869,N_14612,N_14914);
nand U17870 (N_17870,N_14595,N_14744);
and U17871 (N_17871,N_12850,N_14707);
xnor U17872 (N_17872,N_14923,N_13622);
nor U17873 (N_17873,N_13083,N_12224);
or U17874 (N_17874,N_12529,N_12709);
nand U17875 (N_17875,N_12353,N_13835);
nor U17876 (N_17876,N_14455,N_14484);
or U17877 (N_17877,N_12490,N_13678);
nand U17878 (N_17878,N_13842,N_14146);
nor U17879 (N_17879,N_12595,N_14888);
xor U17880 (N_17880,N_14486,N_14059);
nor U17881 (N_17881,N_12711,N_12697);
nor U17882 (N_17882,N_13287,N_12296);
or U17883 (N_17883,N_14053,N_12793);
nor U17884 (N_17884,N_12378,N_14543);
xor U17885 (N_17885,N_13535,N_12943);
or U17886 (N_17886,N_14032,N_14298);
nand U17887 (N_17887,N_12629,N_14417);
and U17888 (N_17888,N_13013,N_12152);
xor U17889 (N_17889,N_12111,N_12635);
nand U17890 (N_17890,N_13387,N_14261);
xnor U17891 (N_17891,N_13965,N_14735);
nand U17892 (N_17892,N_12060,N_13973);
xor U17893 (N_17893,N_12073,N_14015);
nand U17894 (N_17894,N_14950,N_14993);
nand U17895 (N_17895,N_14603,N_12312);
nor U17896 (N_17896,N_13023,N_13409);
or U17897 (N_17897,N_12353,N_14652);
or U17898 (N_17898,N_14950,N_14187);
or U17899 (N_17899,N_12813,N_14136);
or U17900 (N_17900,N_12716,N_13813);
xnor U17901 (N_17901,N_12602,N_14344);
xnor U17902 (N_17902,N_13345,N_14193);
and U17903 (N_17903,N_12353,N_14460);
and U17904 (N_17904,N_13216,N_12070);
xnor U17905 (N_17905,N_12546,N_14493);
or U17906 (N_17906,N_13143,N_12546);
nor U17907 (N_17907,N_12281,N_12079);
and U17908 (N_17908,N_13373,N_12911);
or U17909 (N_17909,N_12721,N_12287);
xnor U17910 (N_17910,N_12078,N_14457);
nand U17911 (N_17911,N_12223,N_12697);
nand U17912 (N_17912,N_14921,N_14073);
xor U17913 (N_17913,N_13210,N_14907);
nor U17914 (N_17914,N_13891,N_13225);
nor U17915 (N_17915,N_12580,N_12712);
nor U17916 (N_17916,N_13215,N_13042);
or U17917 (N_17917,N_12680,N_14513);
nand U17918 (N_17918,N_12111,N_14332);
nor U17919 (N_17919,N_13562,N_13454);
xor U17920 (N_17920,N_14016,N_12621);
nand U17921 (N_17921,N_13971,N_14460);
xnor U17922 (N_17922,N_12455,N_13621);
xor U17923 (N_17923,N_12538,N_12361);
nand U17924 (N_17924,N_13995,N_14899);
nand U17925 (N_17925,N_14314,N_12709);
nor U17926 (N_17926,N_14212,N_13511);
or U17927 (N_17927,N_13188,N_14453);
and U17928 (N_17928,N_14798,N_12286);
nand U17929 (N_17929,N_12298,N_13375);
nor U17930 (N_17930,N_14268,N_14946);
nand U17931 (N_17931,N_14003,N_12868);
and U17932 (N_17932,N_13850,N_13029);
and U17933 (N_17933,N_13704,N_13461);
or U17934 (N_17934,N_12914,N_12353);
or U17935 (N_17935,N_14484,N_14774);
nor U17936 (N_17936,N_14652,N_13667);
nor U17937 (N_17937,N_14833,N_12302);
nor U17938 (N_17938,N_14917,N_12229);
or U17939 (N_17939,N_14349,N_13093);
nor U17940 (N_17940,N_12820,N_13126);
xor U17941 (N_17941,N_14200,N_13905);
nand U17942 (N_17942,N_12803,N_12820);
xnor U17943 (N_17943,N_13020,N_12635);
or U17944 (N_17944,N_12061,N_13252);
nand U17945 (N_17945,N_14132,N_12349);
and U17946 (N_17946,N_13721,N_13551);
nor U17947 (N_17947,N_14220,N_13420);
xnor U17948 (N_17948,N_14587,N_14818);
or U17949 (N_17949,N_13490,N_12210);
and U17950 (N_17950,N_13396,N_14326);
nand U17951 (N_17951,N_14346,N_13757);
xnor U17952 (N_17952,N_14064,N_12635);
or U17953 (N_17953,N_12325,N_12136);
and U17954 (N_17954,N_13844,N_14776);
or U17955 (N_17955,N_14687,N_12293);
and U17956 (N_17956,N_14695,N_12653);
and U17957 (N_17957,N_13545,N_14816);
nor U17958 (N_17958,N_14792,N_13528);
nor U17959 (N_17959,N_13365,N_12145);
or U17960 (N_17960,N_12797,N_12722);
nand U17961 (N_17961,N_12190,N_14679);
xnor U17962 (N_17962,N_14587,N_13899);
nand U17963 (N_17963,N_14762,N_13502);
nor U17964 (N_17964,N_14859,N_13410);
or U17965 (N_17965,N_12060,N_14129);
or U17966 (N_17966,N_12316,N_12681);
xor U17967 (N_17967,N_14839,N_14677);
or U17968 (N_17968,N_13827,N_13411);
nor U17969 (N_17969,N_13251,N_14273);
nor U17970 (N_17970,N_13901,N_12234);
or U17971 (N_17971,N_13413,N_14849);
nor U17972 (N_17972,N_13403,N_14915);
xor U17973 (N_17973,N_14384,N_12169);
nand U17974 (N_17974,N_12042,N_13825);
or U17975 (N_17975,N_14957,N_12607);
and U17976 (N_17976,N_13259,N_14188);
nand U17977 (N_17977,N_14965,N_13657);
nand U17978 (N_17978,N_13445,N_14644);
nor U17979 (N_17979,N_13142,N_13366);
or U17980 (N_17980,N_14567,N_12476);
and U17981 (N_17981,N_14040,N_14045);
nor U17982 (N_17982,N_14894,N_13018);
and U17983 (N_17983,N_14962,N_14242);
nor U17984 (N_17984,N_12537,N_12631);
and U17985 (N_17985,N_13603,N_13229);
or U17986 (N_17986,N_14200,N_12653);
and U17987 (N_17987,N_14635,N_12257);
and U17988 (N_17988,N_12562,N_14282);
and U17989 (N_17989,N_12655,N_14934);
nor U17990 (N_17990,N_13066,N_12596);
nor U17991 (N_17991,N_12897,N_12378);
and U17992 (N_17992,N_13363,N_14447);
and U17993 (N_17993,N_14077,N_12081);
xnor U17994 (N_17994,N_13847,N_14661);
nor U17995 (N_17995,N_13802,N_13800);
nand U17996 (N_17996,N_14898,N_14363);
xor U17997 (N_17997,N_13296,N_13478);
xor U17998 (N_17998,N_12962,N_14654);
nor U17999 (N_17999,N_14664,N_12242);
nand U18000 (N_18000,N_15624,N_15124);
nor U18001 (N_18001,N_15632,N_16055);
nand U18002 (N_18002,N_15305,N_15725);
and U18003 (N_18003,N_16105,N_15369);
xnor U18004 (N_18004,N_17799,N_17607);
or U18005 (N_18005,N_17075,N_17735);
nor U18006 (N_18006,N_15067,N_15488);
nand U18007 (N_18007,N_17967,N_15247);
nor U18008 (N_18008,N_17141,N_16126);
nor U18009 (N_18009,N_16262,N_17055);
nand U18010 (N_18010,N_15717,N_15393);
or U18011 (N_18011,N_17618,N_15076);
or U18012 (N_18012,N_17479,N_16030);
nor U18013 (N_18013,N_15586,N_15354);
and U18014 (N_18014,N_17155,N_15244);
and U18015 (N_18015,N_17498,N_15157);
nand U18016 (N_18016,N_15591,N_17530);
nor U18017 (N_18017,N_15439,N_16177);
nor U18018 (N_18018,N_15196,N_15803);
or U18019 (N_18019,N_16928,N_16589);
and U18020 (N_18020,N_17388,N_17246);
xor U18021 (N_18021,N_17980,N_16781);
and U18022 (N_18022,N_17296,N_16595);
xnor U18023 (N_18023,N_16682,N_16077);
nand U18024 (N_18024,N_15538,N_15818);
or U18025 (N_18025,N_15722,N_15989);
or U18026 (N_18026,N_17177,N_17825);
nand U18027 (N_18027,N_16817,N_17098);
nor U18028 (N_18028,N_17109,N_17727);
nor U18029 (N_18029,N_17092,N_15576);
nand U18030 (N_18030,N_17969,N_15512);
nand U18031 (N_18031,N_17736,N_17630);
and U18032 (N_18032,N_16993,N_15901);
and U18033 (N_18033,N_16675,N_17335);
nand U18034 (N_18034,N_16558,N_17781);
nor U18035 (N_18035,N_17250,N_15056);
xor U18036 (N_18036,N_17370,N_17993);
xnor U18037 (N_18037,N_17175,N_15492);
or U18038 (N_18038,N_16364,N_16261);
nand U18039 (N_18039,N_16286,N_16205);
xnor U18040 (N_18040,N_16348,N_17280);
and U18041 (N_18041,N_17531,N_15893);
nand U18042 (N_18042,N_16918,N_17716);
and U18043 (N_18043,N_15548,N_17183);
nand U18044 (N_18044,N_16838,N_15353);
nor U18045 (N_18045,N_16629,N_16909);
and U18046 (N_18046,N_16999,N_16665);
xor U18047 (N_18047,N_17744,N_15294);
and U18048 (N_18048,N_17963,N_15690);
and U18049 (N_18049,N_17649,N_17096);
xor U18050 (N_18050,N_15404,N_17095);
nand U18051 (N_18051,N_17717,N_17546);
nor U18052 (N_18052,N_16094,N_15060);
nand U18053 (N_18053,N_17356,N_15590);
nand U18054 (N_18054,N_17263,N_16718);
xnor U18055 (N_18055,N_15934,N_15481);
nand U18056 (N_18056,N_15832,N_17686);
nand U18057 (N_18057,N_16810,N_17934);
or U18058 (N_18058,N_16988,N_15317);
nor U18059 (N_18059,N_16995,N_15553);
or U18060 (N_18060,N_15332,N_16465);
xnor U18061 (N_18061,N_17537,N_15847);
xor U18062 (N_18062,N_15065,N_17099);
xor U18063 (N_18063,N_16968,N_15231);
nor U18064 (N_18064,N_15707,N_15057);
nor U18065 (N_18065,N_16901,N_15559);
nand U18066 (N_18066,N_15688,N_15092);
or U18067 (N_18067,N_15098,N_17289);
and U18068 (N_18068,N_15631,N_17854);
and U18069 (N_18069,N_16756,N_16827);
xnor U18070 (N_18070,N_17170,N_17880);
nand U18071 (N_18071,N_15461,N_17711);
nand U18072 (N_18072,N_17154,N_16764);
and U18073 (N_18073,N_15437,N_17312);
or U18074 (N_18074,N_17371,N_16564);
xnor U18075 (N_18075,N_17331,N_17938);
nor U18076 (N_18076,N_15568,N_16867);
xor U18077 (N_18077,N_15849,N_15822);
xor U18078 (N_18078,N_15851,N_16463);
nand U18079 (N_18079,N_17857,N_15699);
or U18080 (N_18080,N_16899,N_16639);
nand U18081 (N_18081,N_16972,N_15216);
xor U18082 (N_18082,N_16248,N_15182);
nand U18083 (N_18083,N_17569,N_15623);
and U18084 (N_18084,N_17150,N_15450);
and U18085 (N_18085,N_17439,N_17016);
nand U18086 (N_18086,N_17683,N_15258);
nand U18087 (N_18087,N_16686,N_17084);
nand U18088 (N_18088,N_17604,N_16638);
nor U18089 (N_18089,N_17281,N_15173);
nor U18090 (N_18090,N_16232,N_17153);
xnor U18091 (N_18091,N_16888,N_15636);
xor U18092 (N_18092,N_15443,N_16402);
nor U18093 (N_18093,N_17750,N_16976);
and U18094 (N_18094,N_15121,N_15563);
nand U18095 (N_18095,N_16354,N_15694);
xor U18096 (N_18096,N_17412,N_15455);
or U18097 (N_18097,N_16302,N_17087);
nor U18098 (N_18098,N_16869,N_16893);
xnor U18099 (N_18099,N_17243,N_17036);
nor U18100 (N_18100,N_16914,N_15695);
nor U18101 (N_18101,N_17915,N_16255);
nand U18102 (N_18102,N_15544,N_17533);
and U18103 (N_18103,N_16074,N_17071);
nor U18104 (N_18104,N_16678,N_16046);
xor U18105 (N_18105,N_16554,N_17186);
or U18106 (N_18106,N_15178,N_17432);
or U18107 (N_18107,N_17529,N_16852);
and U18108 (N_18108,N_15673,N_15606);
xnor U18109 (N_18109,N_15096,N_16712);
xnor U18110 (N_18110,N_17396,N_17078);
xor U18111 (N_18111,N_15165,N_15295);
nand U18112 (N_18112,N_16331,N_16966);
nor U18113 (N_18113,N_16104,N_17540);
xnor U18114 (N_18114,N_15891,N_15167);
nand U18115 (N_18115,N_17849,N_16184);
nand U18116 (N_18116,N_16380,N_16506);
nor U18117 (N_18117,N_16920,N_17167);
nand U18118 (N_18118,N_15184,N_15614);
or U18119 (N_18119,N_16053,N_16394);
xnor U18120 (N_18120,N_16926,N_17433);
nand U18121 (N_18121,N_16752,N_16258);
or U18122 (N_18122,N_17741,N_16509);
and U18123 (N_18123,N_15719,N_15028);
or U18124 (N_18124,N_15616,N_17062);
xor U18125 (N_18125,N_16118,N_15651);
nor U18126 (N_18126,N_16950,N_16193);
nor U18127 (N_18127,N_16359,N_17176);
xor U18128 (N_18128,N_16736,N_17444);
or U18129 (N_18129,N_16524,N_17000);
or U18130 (N_18130,N_17635,N_15844);
xnor U18131 (N_18131,N_16809,N_15612);
nor U18132 (N_18132,N_17621,N_15886);
xnor U18133 (N_18133,N_17774,N_16617);
and U18134 (N_18134,N_15012,N_16056);
nand U18135 (N_18135,N_15030,N_15865);
and U18136 (N_18136,N_17764,N_17509);
nor U18137 (N_18137,N_15147,N_16553);
and U18138 (N_18138,N_17605,N_15392);
nor U18139 (N_18139,N_17572,N_15206);
and U18140 (N_18140,N_16494,N_16883);
or U18141 (N_18141,N_15903,N_17279);
nor U18142 (N_18142,N_15997,N_17989);
and U18143 (N_18143,N_15641,N_16314);
nand U18144 (N_18144,N_15984,N_17020);
and U18145 (N_18145,N_15086,N_17470);
xnor U18146 (N_18146,N_17222,N_17972);
nor U18147 (N_18147,N_15445,N_16823);
xnor U18148 (N_18148,N_15728,N_16991);
nand U18149 (N_18149,N_16338,N_16604);
nand U18150 (N_18150,N_15644,N_15667);
and U18151 (N_18151,N_16133,N_15554);
nand U18152 (N_18152,N_16640,N_16796);
nand U18153 (N_18153,N_17401,N_15136);
nand U18154 (N_18154,N_16176,N_15780);
nand U18155 (N_18155,N_16215,N_17364);
nor U18156 (N_18156,N_15960,N_15050);
xnor U18157 (N_18157,N_15221,N_16711);
or U18158 (N_18158,N_16708,N_17395);
nand U18159 (N_18159,N_17687,N_15407);
nor U18160 (N_18160,N_15600,N_17107);
nor U18161 (N_18161,N_15267,N_16769);
xnor U18162 (N_18162,N_15465,N_16908);
xor U18163 (N_18163,N_17464,N_15498);
nand U18164 (N_18164,N_15877,N_17903);
and U18165 (N_18165,N_17944,N_15558);
and U18166 (N_18166,N_16260,N_15471);
or U18167 (N_18167,N_16361,N_15916);
or U18168 (N_18168,N_16814,N_15045);
xnor U18169 (N_18169,N_16275,N_15210);
nand U18170 (N_18170,N_16556,N_16862);
xnor U18171 (N_18171,N_16543,N_17112);
nor U18172 (N_18172,N_17860,N_16477);
or U18173 (N_18173,N_15000,N_16868);
nand U18174 (N_18174,N_15078,N_16825);
or U18175 (N_18175,N_16378,N_17419);
nor U18176 (N_18176,N_16561,N_15079);
and U18177 (N_18177,N_15489,N_15467);
xnor U18178 (N_18178,N_17230,N_16481);
or U18179 (N_18179,N_15827,N_16643);
xnor U18180 (N_18180,N_15841,N_15930);
nand U18181 (N_18181,N_17088,N_16609);
xor U18182 (N_18182,N_15052,N_16854);
or U18183 (N_18183,N_15625,N_16967);
nor U18184 (N_18184,N_17874,N_17643);
nor U18185 (N_18185,N_15910,N_16186);
nor U18186 (N_18186,N_15309,N_16947);
nor U18187 (N_18187,N_15145,N_16312);
nor U18188 (N_18188,N_15497,N_15806);
nor U18189 (N_18189,N_17747,N_16132);
nor U18190 (N_18190,N_17213,N_17157);
or U18191 (N_18191,N_17592,N_16803);
and U18192 (N_18192,N_16971,N_15172);
and U18193 (N_18193,N_17424,N_17478);
xor U18194 (N_18194,N_16033,N_15581);
nand U18195 (N_18195,N_15004,N_15589);
or U18196 (N_18196,N_16771,N_16086);
or U18197 (N_18197,N_17757,N_16517);
or U18198 (N_18198,N_15368,N_15863);
nand U18199 (N_18199,N_15367,N_15560);
and U18200 (N_18200,N_16801,N_16401);
or U18201 (N_18201,N_16614,N_17366);
and U18202 (N_18202,N_15618,N_15550);
nor U18203 (N_18203,N_15103,N_16171);
nor U18204 (N_18204,N_17159,N_17974);
nor U18205 (N_18205,N_15441,N_17120);
and U18206 (N_18206,N_17059,N_16121);
xor U18207 (N_18207,N_15879,N_17876);
xor U18208 (N_18208,N_17057,N_17228);
xnor U18209 (N_18209,N_16329,N_17574);
or U18210 (N_18210,N_16376,N_17952);
xnor U18211 (N_18211,N_17818,N_17805);
nor U18212 (N_18212,N_15420,N_15639);
and U18213 (N_18213,N_17698,N_15338);
and U18214 (N_18214,N_15015,N_15998);
and U18215 (N_18215,N_17066,N_16478);
and U18216 (N_18216,N_17520,N_17129);
or U18217 (N_18217,N_17385,N_16479);
xor U18218 (N_18218,N_15737,N_15711);
nor U18219 (N_18219,N_16324,N_17301);
nand U18220 (N_18220,N_17955,N_15684);
nand U18221 (N_18221,N_17442,N_17169);
xor U18222 (N_18222,N_15671,N_16052);
and U18223 (N_18223,N_17060,N_16588);
xnor U18224 (N_18224,N_17966,N_16570);
and U18225 (N_18225,N_16243,N_15941);
nand U18226 (N_18226,N_15784,N_17551);
nor U18227 (N_18227,N_15449,N_15205);
nand U18228 (N_18228,N_17914,N_15867);
nand U18229 (N_18229,N_16894,N_15494);
nor U18230 (N_18230,N_17429,N_17708);
xnor U18231 (N_18231,N_16034,N_15245);
nor U18232 (N_18232,N_15848,N_15238);
or U18233 (N_18233,N_15773,N_16577);
or U18234 (N_18234,N_16419,N_17068);
nor U18235 (N_18235,N_16473,N_15705);
xnor U18236 (N_18236,N_16565,N_15055);
and U18237 (N_18237,N_17695,N_16377);
and U18238 (N_18238,N_15232,N_17143);
and U18239 (N_18239,N_15111,N_17227);
nor U18240 (N_18240,N_16502,N_16946);
nand U18241 (N_18241,N_16226,N_15209);
or U18242 (N_18242,N_16089,N_16310);
and U18243 (N_18243,N_17270,N_17146);
nor U18244 (N_18244,N_17160,N_15168);
or U18245 (N_18245,N_16891,N_17072);
xnor U18246 (N_18246,N_17488,N_15575);
or U18247 (N_18247,N_15970,N_15036);
and U18248 (N_18248,N_15809,N_16169);
or U18249 (N_18249,N_16684,N_15657);
or U18250 (N_18250,N_17471,N_16211);
xor U18251 (N_18251,N_17856,N_17158);
nor U18252 (N_18252,N_16602,N_15552);
and U18253 (N_18253,N_17802,N_17156);
or U18254 (N_18254,N_15402,N_16592);
nand U18255 (N_18255,N_17130,N_15643);
or U18256 (N_18256,N_15220,N_16351);
and U18257 (N_18257,N_16871,N_16621);
nor U18258 (N_18258,N_17988,N_17767);
nand U18259 (N_18259,N_16192,N_15536);
nand U18260 (N_18260,N_15509,N_15307);
nor U18261 (N_18261,N_16627,N_16811);
xor U18262 (N_18262,N_16141,N_17584);
nand U18263 (N_18263,N_16548,N_16283);
and U18264 (N_18264,N_17714,N_17796);
nor U18265 (N_18265,N_15514,N_17642);
or U18266 (N_18266,N_17204,N_17305);
or U18267 (N_18267,N_17571,N_15740);
or U18268 (N_18268,N_16043,N_17188);
xnor U18269 (N_18269,N_17221,N_17600);
or U18270 (N_18270,N_17115,N_16196);
nand U18271 (N_18271,N_16280,N_17956);
and U18272 (N_18272,N_17885,N_16008);
or U18273 (N_18273,N_17996,N_16016);
or U18274 (N_18274,N_16953,N_17503);
or U18275 (N_18275,N_15426,N_15693);
nor U18276 (N_18276,N_16398,N_17214);
and U18277 (N_18277,N_16486,N_15284);
and U18278 (N_18278,N_15807,N_16415);
xor U18279 (N_18279,N_16751,N_17045);
nand U18280 (N_18280,N_15106,N_16674);
or U18281 (N_18281,N_17191,N_17873);
nand U18282 (N_18282,N_17768,N_15381);
nor U18283 (N_18283,N_17677,N_17065);
or U18284 (N_18284,N_15943,N_16204);
or U18285 (N_18285,N_17931,N_16453);
nor U18286 (N_18286,N_15878,N_17233);
xor U18287 (N_18287,N_15491,N_17933);
and U18288 (N_18288,N_15597,N_16225);
nand U18289 (N_18289,N_16601,N_15107);
and U18290 (N_18290,N_17042,N_16484);
nand U18291 (N_18291,N_17784,N_16590);
or U18292 (N_18292,N_16145,N_16518);
nand U18293 (N_18293,N_16689,N_15174);
nand U18294 (N_18294,N_16531,N_15884);
or U18295 (N_18295,N_17399,N_17467);
and U18296 (N_18296,N_17542,N_16207);
nor U18297 (N_18297,N_15403,N_15649);
or U18298 (N_18298,N_17681,N_17426);
nor U18299 (N_18299,N_17679,N_16285);
nand U18300 (N_18300,N_17434,N_16358);
nor U18301 (N_18301,N_17947,N_16071);
nand U18302 (N_18302,N_17653,N_17423);
nor U18303 (N_18303,N_15490,N_15023);
xnor U18304 (N_18304,N_16786,N_15897);
nand U18305 (N_18305,N_15311,N_15274);
and U18306 (N_18306,N_16010,N_15314);
xnor U18307 (N_18307,N_16519,N_17127);
xor U18308 (N_18308,N_15090,N_17164);
nand U18309 (N_18309,N_17178,N_16392);
xor U18310 (N_18310,N_16696,N_17553);
xor U18311 (N_18311,N_16581,N_15918);
nor U18312 (N_18312,N_15059,N_16902);
or U18313 (N_18313,N_16470,N_16699);
or U18314 (N_18314,N_17319,N_17459);
xnor U18315 (N_18315,N_15042,N_16450);
nand U18316 (N_18316,N_17665,N_15885);
nand U18317 (N_18317,N_15953,N_17329);
nand U18318 (N_18318,N_16001,N_15919);
and U18319 (N_18319,N_16093,N_15308);
nand U18320 (N_18320,N_16005,N_16713);
and U18321 (N_18321,N_15962,N_17007);
nor U18322 (N_18322,N_16998,N_16220);
xor U18323 (N_18323,N_16679,N_15801);
xnor U18324 (N_18324,N_15881,N_17916);
nor U18325 (N_18325,N_17050,N_15828);
or U18326 (N_18326,N_16218,N_15120);
or U18327 (N_18327,N_17678,N_15040);
nand U18328 (N_18328,N_15158,N_15333);
xnor U18329 (N_18329,N_16580,N_17124);
nor U18330 (N_18330,N_15224,N_16746);
nor U18331 (N_18331,N_17234,N_16963);
xnor U18332 (N_18332,N_15845,N_15902);
and U18333 (N_18333,N_15790,N_16791);
nor U18334 (N_18334,N_16961,N_17843);
nor U18335 (N_18335,N_15169,N_15565);
or U18336 (N_18336,N_15080,N_16240);
or U18337 (N_18337,N_15676,N_16870);
xor U18338 (N_18338,N_16701,N_15975);
xnor U18339 (N_18339,N_17094,N_15410);
nand U18340 (N_18340,N_15593,N_17220);
xnor U18341 (N_18341,N_17456,N_17252);
and U18342 (N_18342,N_16641,N_16740);
and U18343 (N_18343,N_15003,N_15947);
or U18344 (N_18344,N_16722,N_15914);
nand U18345 (N_18345,N_15416,N_15925);
and U18346 (N_18346,N_15540,N_15142);
and U18347 (N_18347,N_15131,N_16514);
nand U18348 (N_18348,N_16308,N_15044);
nand U18349 (N_18349,N_16793,N_16692);
xor U18350 (N_18350,N_15992,N_15104);
nor U18351 (N_18351,N_16539,N_17773);
xor U18352 (N_18352,N_15689,N_16384);
or U18353 (N_18353,N_17726,N_17122);
and U18354 (N_18354,N_17499,N_16977);
nor U18355 (N_18355,N_16299,N_17704);
and U18356 (N_18356,N_15150,N_17593);
and U18357 (N_18357,N_16198,N_15379);
and U18358 (N_18358,N_16457,N_16025);
nand U18359 (N_18359,N_16270,N_16824);
xor U18360 (N_18360,N_15061,N_17077);
and U18361 (N_18361,N_15990,N_15789);
or U18362 (N_18362,N_17877,N_15039);
or U18363 (N_18363,N_17591,N_15634);
or U18364 (N_18364,N_17882,N_15459);
and U18365 (N_18365,N_15742,N_17920);
and U18366 (N_18366,N_15419,N_15802);
nor U18367 (N_18367,N_17121,N_15460);
xor U18368 (N_18368,N_15001,N_16122);
nor U18369 (N_18369,N_15500,N_15347);
xnor U18370 (N_18370,N_16172,N_16974);
nor U18371 (N_18371,N_17589,N_17923);
nand U18372 (N_18372,N_16944,N_17082);
and U18373 (N_18373,N_15999,N_16488);
and U18374 (N_18374,N_16167,N_16440);
and U18375 (N_18375,N_17336,N_16181);
nor U18376 (N_18376,N_16252,N_16128);
nand U18377 (N_18377,N_17063,N_17842);
nor U18378 (N_18378,N_16654,N_17615);
xnor U18379 (N_18379,N_15718,N_17291);
or U18380 (N_18380,N_17514,N_16097);
or U18381 (N_18381,N_17494,N_16098);
or U18382 (N_18382,N_16800,N_17673);
and U18383 (N_18383,N_17196,N_17637);
or U18384 (N_18384,N_17868,N_16476);
xor U18385 (N_18385,N_15273,N_17561);
xnor U18386 (N_18386,N_15607,N_16960);
nor U18387 (N_18387,N_15937,N_15991);
nand U18388 (N_18388,N_17205,N_16731);
xor U18389 (N_18389,N_17184,N_17041);
nor U18390 (N_18390,N_15127,N_15513);
nand U18391 (N_18391,N_16087,N_16247);
xor U18392 (N_18392,N_17583,N_15799);
nand U18393 (N_18393,N_15763,N_16085);
or U18394 (N_18394,N_15720,N_15432);
and U18395 (N_18395,N_17602,N_17131);
xnor U18396 (N_18396,N_16497,N_16028);
nor U18397 (N_18397,N_16289,N_15954);
xnor U18398 (N_18398,N_15447,N_15924);
or U18399 (N_18399,N_17634,N_16075);
nand U18400 (N_18400,N_17976,N_17534);
nor U18401 (N_18401,N_16015,N_15895);
and U18402 (N_18402,N_16815,N_17435);
and U18403 (N_18403,N_15939,N_15415);
nand U18404 (N_18404,N_17443,N_16630);
and U18405 (N_18405,N_16103,N_17705);
nor U18406 (N_18406,N_15986,N_16691);
xor U18407 (N_18407,N_15977,N_15279);
xor U18408 (N_18408,N_15980,N_16620);
xor U18409 (N_18409,N_16668,N_16549);
nor U18410 (N_18410,N_16720,N_17828);
xnor U18411 (N_18411,N_15280,N_15824);
xnor U18412 (N_18412,N_16843,N_17853);
nand U18413 (N_18413,N_15268,N_15647);
nand U18414 (N_18414,N_16848,N_16572);
xnor U18415 (N_18415,N_16356,N_16491);
or U18416 (N_18416,N_16582,N_17431);
or U18417 (N_18417,N_15176,N_17939);
nand U18418 (N_18418,N_16131,N_15423);
nand U18419 (N_18419,N_15709,N_15088);
nand U18420 (N_18420,N_15013,N_15582);
nand U18421 (N_18421,N_16109,N_16726);
nor U18422 (N_18422,N_17053,N_17556);
xnor U18423 (N_18423,N_17611,N_17804);
nor U18424 (N_18424,N_15222,N_16608);
xnor U18425 (N_18425,N_17626,N_16102);
and U18426 (N_18426,N_15208,N_16236);
or U18427 (N_18427,N_17617,N_15382);
or U18428 (N_18428,N_16265,N_17133);
or U18429 (N_18429,N_16185,N_16858);
nand U18430 (N_18430,N_15219,N_16945);
nor U18431 (N_18431,N_15331,N_15746);
xor U18432 (N_18432,N_17249,N_15094);
and U18433 (N_18433,N_16231,N_17965);
and U18434 (N_18434,N_15633,N_17667);
nand U18435 (N_18435,N_17766,N_15257);
nand U18436 (N_18436,N_15965,N_17943);
nor U18437 (N_18437,N_16168,N_15336);
or U18438 (N_18438,N_16606,N_16301);
and U18439 (N_18439,N_17565,N_17048);
xor U18440 (N_18440,N_17547,N_15906);
nor U18441 (N_18441,N_15783,N_17454);
nand U18442 (N_18442,N_15805,N_16940);
nor U18443 (N_18443,N_15434,N_17447);
xor U18444 (N_18444,N_16532,N_15371);
and U18445 (N_18445,N_17732,N_17921);
nand U18446 (N_18446,N_16831,N_16957);
nor U18447 (N_18447,N_15285,N_16778);
and U18448 (N_18448,N_17614,N_15089);
nor U18449 (N_18449,N_16566,N_16253);
nand U18450 (N_18450,N_16449,N_15189);
nor U18451 (N_18451,N_16395,N_16545);
or U18452 (N_18452,N_15363,N_16335);
nand U18453 (N_18453,N_17723,N_16472);
nand U18454 (N_18454,N_15923,N_15656);
and U18455 (N_18455,N_17746,N_17603);
and U18456 (N_18456,N_17363,N_15674);
nor U18457 (N_18457,N_16146,N_15862);
and U18458 (N_18458,N_16559,N_15944);
or U18459 (N_18459,N_17719,N_17646);
nand U18460 (N_18460,N_17881,N_16941);
or U18461 (N_18461,N_17421,N_17526);
or U18462 (N_18462,N_15681,N_15396);
nand U18463 (N_18463,N_15532,N_17525);
and U18464 (N_18464,N_17508,N_17599);
and U18465 (N_18465,N_15502,N_17638);
and U18466 (N_18466,N_15611,N_17919);
xor U18467 (N_18467,N_16124,N_15712);
nand U18468 (N_18468,N_17625,N_16644);
and U18469 (N_18469,N_16607,N_15011);
or U18470 (N_18470,N_15974,N_16078);
nand U18471 (N_18471,N_15302,N_16383);
and U18472 (N_18472,N_16400,N_17765);
and U18473 (N_18473,N_15242,N_17436);
or U18474 (N_18474,N_16673,N_16422);
nor U18475 (N_18475,N_17061,N_17536);
nand U18476 (N_18476,N_17307,N_17986);
nor U18477 (N_18477,N_16323,N_15894);
xnor U18478 (N_18478,N_15635,N_16845);
and U18479 (N_18479,N_17003,N_16563);
and U18480 (N_18480,N_17393,N_17497);
xor U18481 (N_18481,N_17144,N_15515);
nand U18482 (N_18482,N_15567,N_17418);
nor U18483 (N_18483,N_16203,N_16035);
or U18484 (N_18484,N_15981,N_17693);
nand U18485 (N_18485,N_17240,N_16032);
xnor U18486 (N_18486,N_15064,N_15156);
or U18487 (N_18487,N_16738,N_15017);
or U18488 (N_18488,N_16975,N_15829);
or U18489 (N_18489,N_16355,N_16004);
and U18490 (N_18490,N_15495,N_15774);
or U18491 (N_18491,N_16886,N_17247);
xor U18492 (N_18492,N_17725,N_15475);
xnor U18493 (N_18493,N_15324,N_16520);
xnor U18494 (N_18494,N_17703,N_15759);
or U18495 (N_18495,N_17215,N_17317);
xnor U18496 (N_18496,N_15234,N_16487);
and U18497 (N_18497,N_16292,N_17851);
or U18498 (N_18498,N_17025,N_15431);
nor U18499 (N_18499,N_16774,N_16325);
or U18500 (N_18500,N_16705,N_17680);
nand U18501 (N_18501,N_17244,N_17970);
or U18502 (N_18502,N_16863,N_15063);
nand U18503 (N_18503,N_17272,N_16856);
nor U18504 (N_18504,N_16057,N_17869);
nor U18505 (N_18505,N_17422,N_15508);
or U18506 (N_18506,N_15398,N_17720);
nand U18507 (N_18507,N_17290,N_17081);
or U18508 (N_18508,N_16081,N_16239);
nand U18509 (N_18509,N_17787,N_17946);
nand U18510 (N_18510,N_15504,N_16567);
xor U18511 (N_18511,N_17002,N_17913);
and U18512 (N_18512,N_15610,N_16223);
or U18513 (N_18513,N_15665,N_17912);
or U18514 (N_18514,N_15670,N_17192);
nand U18515 (N_18515,N_16651,N_16388);
nand U18516 (N_18516,N_16938,N_15605);
nand U18517 (N_18517,N_16861,N_15282);
nand U18518 (N_18518,N_16061,N_16140);
nor U18519 (N_18519,N_17866,N_17341);
or U18520 (N_18520,N_17559,N_15648);
or U18521 (N_18521,N_17554,N_16147);
or U18522 (N_18522,N_16522,N_16763);
or U18523 (N_18523,N_16733,N_17566);
nand U18524 (N_18524,N_16294,N_16983);
xnor U18525 (N_18525,N_15679,N_15892);
xor U18526 (N_18526,N_17269,N_16943);
xor U18527 (N_18527,N_16284,N_17871);
xor U18528 (N_18528,N_17438,N_15171);
nor U18529 (N_18529,N_17266,N_16024);
and U18530 (N_18530,N_16955,N_16904);
nor U18531 (N_18531,N_17231,N_15794);
nor U18532 (N_18532,N_15020,N_17809);
or U18533 (N_18533,N_15692,N_15573);
or U18534 (N_18534,N_16139,N_17445);
or U18535 (N_18535,N_17962,N_17051);
xor U18536 (N_18536,N_15561,N_15866);
nand U18537 (N_18537,N_17959,N_15503);
nor U18538 (N_18538,N_17430,N_17119);
nor U18539 (N_18539,N_17031,N_15109);
or U18540 (N_18540,N_16156,N_15372);
nor U18541 (N_18541,N_16949,N_15519);
and U18542 (N_18542,N_16962,N_15510);
nand U18543 (N_18543,N_15797,N_15162);
xor U18544 (N_18544,N_17772,N_16633);
or U18545 (N_18545,N_17046,N_15915);
nand U18546 (N_18546,N_15430,N_16163);
and U18547 (N_18547,N_15723,N_17343);
nand U18548 (N_18548,N_16427,N_17300);
nand U18549 (N_18549,N_17174,N_17878);
or U18550 (N_18550,N_15596,N_16836);
nand U18551 (N_18551,N_17694,N_16346);
nor U18552 (N_18552,N_16064,N_17032);
nand U18553 (N_18553,N_16026,N_17052);
nand U18554 (N_18554,N_15298,N_16221);
nor U18555 (N_18555,N_15959,N_16397);
nor U18556 (N_18556,N_16505,N_16271);
xor U18557 (N_18557,N_15254,N_15026);
nand U18558 (N_18558,N_16038,N_17648);
and U18559 (N_18559,N_16027,N_17058);
nand U18560 (N_18560,N_17811,N_16144);
xnor U18561 (N_18561,N_16729,N_15444);
nand U18562 (N_18562,N_17511,N_17391);
xor U18563 (N_18563,N_16175,N_15956);
and U18564 (N_18564,N_17889,N_16461);
or U18565 (N_18565,N_16528,N_17461);
xor U18566 (N_18566,N_15541,N_15047);
or U18567 (N_18567,N_17203,N_17954);
xnor U18568 (N_18568,N_17163,N_15873);
nor U18569 (N_18569,N_15710,N_15485);
or U18570 (N_18570,N_15457,N_17575);
xnor U18571 (N_18571,N_16490,N_16723);
nand U18572 (N_18572,N_15243,N_15091);
and U18573 (N_18573,N_15726,N_15227);
xor U18574 (N_18574,N_17786,N_15170);
nand U18575 (N_18575,N_16922,N_16613);
nor U18576 (N_18576,N_15842,N_15875);
nor U18577 (N_18577,N_17753,N_16772);
or U18578 (N_18578,N_15337,N_15413);
nand U18579 (N_18579,N_17612,N_15778);
xnor U18580 (N_18580,N_16658,N_15128);
nor U18581 (N_18581,N_16768,N_16321);
xor U18582 (N_18582,N_15380,N_15961);
xnor U18583 (N_18583,N_17864,N_15889);
and U18584 (N_18584,N_17998,N_17613);
nand U18585 (N_18585,N_15530,N_15101);
or U18586 (N_18586,N_17728,N_17911);
or U18587 (N_18587,N_15537,N_17794);
nor U18588 (N_18588,N_15249,N_17006);
nor U18589 (N_18589,N_16919,N_15239);
nand U18590 (N_18590,N_16882,N_16948);
nor U18591 (N_18591,N_15191,N_15230);
xor U18592 (N_18592,N_16448,N_16534);
xor U18593 (N_18593,N_16363,N_16443);
xor U18594 (N_18594,N_16915,N_16821);
xnor U18595 (N_18595,N_15518,N_15228);
nor U18596 (N_18596,N_16138,N_16158);
or U18597 (N_18597,N_16157,N_15539);
nor U18598 (N_18598,N_16896,N_15062);
xnor U18599 (N_18599,N_17594,N_16719);
nor U18600 (N_18600,N_16822,N_15976);
nor U18601 (N_18601,N_17606,N_17659);
xor U18602 (N_18602,N_17629,N_16040);
and U18603 (N_18603,N_17790,N_16773);
or U18604 (N_18604,N_17839,N_17644);
xnor U18605 (N_18605,N_15328,N_16964);
and U18606 (N_18606,N_17951,N_16724);
nor U18607 (N_18607,N_17983,N_17372);
or U18608 (N_18608,N_17162,N_16523);
and U18609 (N_18609,N_15580,N_17776);
nor U18610 (N_18610,N_17754,N_17014);
nand U18611 (N_18611,N_15009,N_16859);
xor U18612 (N_18612,N_15422,N_15179);
and U18613 (N_18613,N_16788,N_15303);
xor U18614 (N_18614,N_17579,N_17785);
or U18615 (N_18615,N_17101,N_17033);
and U18616 (N_18616,N_16182,N_17715);
nand U18617 (N_18617,N_16217,N_17779);
or U18618 (N_18618,N_15043,N_15927);
and U18619 (N_18619,N_16413,N_16041);
xor U18620 (N_18620,N_17090,N_17278);
nor U18621 (N_18621,N_16195,N_15830);
nand U18622 (N_18622,N_16464,N_16533);
and U18623 (N_18623,N_15034,N_16076);
and U18624 (N_18624,N_17513,N_15350);
or U18625 (N_18625,N_16288,N_17495);
nor U18626 (N_18626,N_15342,N_15768);
xnor U18627 (N_18627,N_15387,N_16757);
nand U18628 (N_18628,N_17932,N_15700);
nand U18629 (N_18629,N_16212,N_17858);
nor U18630 (N_18630,N_16535,N_15817);
and U18631 (N_18631,N_17654,N_15329);
and U18632 (N_18632,N_17535,N_16642);
or U18633 (N_18633,N_17179,N_17892);
nor U18634 (N_18634,N_16269,N_15263);
nor U18635 (N_18635,N_16615,N_16066);
nand U18636 (N_18636,N_17697,N_17484);
nand U18637 (N_18637,N_15277,N_17550);
nor U18638 (N_18638,N_16311,N_15972);
and U18639 (N_18639,N_17440,N_15199);
nor U18640 (N_18640,N_15856,N_16462);
xnor U18641 (N_18641,N_15148,N_16127);
nor U18642 (N_18642,N_16625,N_17492);
or U18643 (N_18643,N_16409,N_17895);
and U18644 (N_18644,N_17548,N_16853);
and U18645 (N_18645,N_16222,N_17845);
or U18646 (N_18646,N_17867,N_16447);
nand U18647 (N_18647,N_16530,N_17709);
nand U18648 (N_18648,N_16767,N_17729);
and U18649 (N_18649,N_15758,N_17831);
and U18650 (N_18650,N_15033,N_17333);
or U18651 (N_18651,N_15429,N_17523);
xnor U18652 (N_18652,N_16703,N_17769);
nand U18653 (N_18653,N_17807,N_15203);
xnor U18654 (N_18654,N_17926,N_16337);
and U18655 (N_18655,N_16250,N_17700);
nand U18656 (N_18656,N_15246,N_17350);
nand U18657 (N_18657,N_16734,N_15815);
and U18658 (N_18658,N_17267,N_16550);
or U18659 (N_18659,N_16753,N_15472);
or U18660 (N_18660,N_16515,N_16107);
and U18661 (N_18661,N_16847,N_16605);
or U18662 (N_18662,N_16194,N_15291);
or U18663 (N_18663,N_17834,N_17658);
xnor U18664 (N_18664,N_15283,N_15453);
or U18665 (N_18665,N_16319,N_16579);
xor U18666 (N_18666,N_15792,N_15666);
xnor U18667 (N_18667,N_15855,N_17690);
xor U18668 (N_18668,N_16333,N_16460);
and U18669 (N_18669,N_15564,N_17539);
or U18670 (N_18670,N_16835,N_15900);
or U18671 (N_18671,N_16423,N_16411);
nand U18672 (N_18672,N_17379,N_16467);
nand U18673 (N_18673,N_17225,N_15322);
nand U18674 (N_18674,N_17724,N_17165);
xor U18675 (N_18675,N_17500,N_15340);
or U18676 (N_18676,N_16744,N_17684);
xor U18677 (N_18677,N_15272,N_16159);
xnor U18678 (N_18678,N_15181,N_15370);
nand U18679 (N_18679,N_17285,N_16655);
or U18680 (N_18680,N_16197,N_17288);
nor U18681 (N_18681,N_15438,N_15912);
nor U18682 (N_18682,N_17469,N_15187);
xor U18683 (N_18683,N_16150,N_15201);
xnor U18684 (N_18684,N_15755,N_15253);
and U18685 (N_18685,N_16200,N_16990);
or U18686 (N_18686,N_16952,N_17894);
nand U18687 (N_18687,N_16295,N_17852);
nand U18688 (N_18688,N_15810,N_16037);
or U18689 (N_18689,N_15072,N_17788);
nor U18690 (N_18690,N_17410,N_16510);
and U18691 (N_18691,N_16715,N_15290);
xor U18692 (N_18692,N_15764,N_17778);
xor U18693 (N_18693,N_17472,N_17010);
nor U18694 (N_18694,N_16973,N_16277);
and U18695 (N_18695,N_17749,N_15376);
nand U18696 (N_18696,N_15555,N_15917);
xnor U18697 (N_18697,N_16069,N_17636);
nand U18698 (N_18698,N_15037,N_16575);
nand U18699 (N_18699,N_16263,N_15706);
or U18700 (N_18700,N_15113,N_15535);
xor U18701 (N_18701,N_16166,N_16784);
nand U18702 (N_18702,N_17997,N_15770);
xnor U18703 (N_18703,N_15418,N_15852);
or U18704 (N_18704,N_16492,N_15574);
or U18705 (N_18705,N_17664,N_15193);
xnor U18706 (N_18706,N_17666,N_17688);
and U18707 (N_18707,N_15192,N_15860);
nor U18708 (N_18708,N_16939,N_16246);
or U18709 (N_18709,N_16251,N_17237);
or U18710 (N_18710,N_17206,N_17380);
xnor U18711 (N_18711,N_16916,N_17103);
nand U18712 (N_18712,N_15798,N_17324);
or U18713 (N_18713,N_16136,N_15383);
and U18714 (N_18714,N_17458,N_17202);
nand U18715 (N_18715,N_16698,N_15074);
and U18716 (N_18716,N_16344,N_17655);
nand U18717 (N_18717,N_15602,N_17258);
and U18718 (N_18718,N_17597,N_15983);
nand U18719 (N_18719,N_15456,N_15621);
or U18720 (N_18720,N_15482,N_16597);
and U18721 (N_18721,N_17378,N_15185);
nand U18722 (N_18722,N_17668,N_15138);
nand U18723 (N_18723,N_17522,N_17675);
or U18724 (N_18724,N_15327,N_16622);
nand U18725 (N_18725,N_15880,N_16160);
nor U18726 (N_18726,N_15466,N_16276);
or U18727 (N_18727,N_16979,N_16273);
and U18728 (N_18728,N_15743,N_15365);
xnor U18729 (N_18729,N_15839,N_16790);
or U18730 (N_18730,N_16504,N_16659);
nand U18731 (N_18731,N_17906,N_15926);
nor U18732 (N_18732,N_16282,N_16187);
nor U18733 (N_18733,N_17813,N_17491);
nor U18734 (N_18734,N_15351,N_16014);
nand U18735 (N_18735,N_15412,N_16002);
nand U18736 (N_18736,N_16370,N_16683);
and U18737 (N_18737,N_16956,N_15301);
and U18738 (N_18738,N_17619,N_16671);
nor U18739 (N_18739,N_17320,N_17935);
or U18740 (N_18740,N_15240,N_15745);
nand U18741 (N_18741,N_16892,N_17928);
or U18742 (N_18742,N_17755,N_17573);
xor U18743 (N_18743,N_17581,N_17587);
xor U18744 (N_18744,N_15252,N_15968);
nor U18745 (N_18745,N_15344,N_17822);
nand U18746 (N_18746,N_17453,N_15097);
and U18747 (N_18747,N_17255,N_17855);
nor U18748 (N_18748,N_17441,N_15545);
or U18749 (N_18749,N_17979,N_15619);
or U18750 (N_18750,N_17219,N_17079);
or U18751 (N_18751,N_15077,N_15319);
nand U18752 (N_18752,N_15428,N_15186);
nand U18753 (N_18753,N_15793,N_17731);
or U18754 (N_18754,N_17056,N_15967);
or U18755 (N_18755,N_16309,N_17901);
or U18756 (N_18756,N_16072,N_16485);
and U18757 (N_18757,N_17427,N_17816);
nand U18758 (N_18758,N_17999,N_17721);
xor U18759 (N_18759,N_17013,N_17770);
nor U18760 (N_18760,N_16540,N_17762);
nand U18761 (N_18761,N_16876,N_17359);
nand U18762 (N_18762,N_17128,N_15938);
nand U18763 (N_18763,N_15112,N_17792);
nand U18764 (N_18764,N_16937,N_15276);
and U18765 (N_18765,N_16190,N_17420);
nor U18766 (N_18766,N_15049,N_15084);
xnor U18767 (N_18767,N_15310,N_16741);
or U18768 (N_18768,N_16700,N_15935);
xor U18769 (N_18769,N_17982,N_16587);
nand U18770 (N_18770,N_17413,N_15397);
or U18771 (N_18771,N_17846,N_17995);
nand U18772 (N_18772,N_17315,N_15102);
and U18773 (N_18773,N_17351,N_15598);
xnor U18774 (N_18774,N_16603,N_17030);
nand U18775 (N_18775,N_17806,N_16249);
nand U18776 (N_18776,N_16134,N_17925);
nand U18777 (N_18777,N_17936,N_17891);
or U18778 (N_18778,N_15006,N_15791);
nand U18779 (N_18779,N_17171,N_17620);
nand U18780 (N_18780,N_17287,N_17114);
nand U18781 (N_18781,N_15682,N_17022);
nor U18782 (N_18782,N_17468,N_15942);
nor U18783 (N_18783,N_15008,N_16386);
nand U18784 (N_18784,N_15226,N_15506);
nor U18785 (N_18785,N_15528,N_17113);
xor U18786 (N_18786,N_16842,N_16611);
xnor U18787 (N_18787,N_15587,N_15027);
and U18788 (N_18788,N_17908,N_16739);
and U18789 (N_18789,N_15570,N_16645);
nand U18790 (N_18790,N_16866,N_17416);
nand U18791 (N_18791,N_16594,N_15390);
and U18792 (N_18792,N_16917,N_16278);
nand U18793 (N_18793,N_16923,N_16164);
or U18794 (N_18794,N_16954,N_16884);
nor U18795 (N_18795,N_16857,N_17623);
nand U18796 (N_18796,N_17463,N_17026);
nand U18797 (N_18797,N_15164,N_17309);
or U18798 (N_18798,N_15075,N_15908);
nand U18799 (N_18799,N_16636,N_17166);
and U18800 (N_18800,N_15896,N_16442);
xor U18801 (N_18801,N_17091,N_16501);
xor U18802 (N_18802,N_15480,N_16214);
or U18803 (N_18803,N_16474,N_17819);
nand U18804 (N_18804,N_16578,N_16439);
or U18805 (N_18805,N_16366,N_15031);
and U18806 (N_18806,N_16500,N_17223);
xnor U18807 (N_18807,N_16406,N_17859);
xor U18808 (N_18808,N_16706,N_17283);
nor U18809 (N_18809,N_16599,N_15010);
or U18810 (N_18810,N_16770,N_15479);
nor U18811 (N_18811,N_17557,N_15595);
nor U18812 (N_18812,N_16758,N_17841);
and U18813 (N_18813,N_16327,N_15739);
nor U18814 (N_18814,N_15549,N_17624);
nand U18815 (N_18815,N_16129,N_17872);
nor U18816 (N_18816,N_15775,N_16343);
nand U18817 (N_18817,N_16807,N_15025);
and U18818 (N_18818,N_17824,N_15716);
and U18819 (N_18819,N_17691,N_17820);
or U18820 (N_18820,N_16924,N_16108);
nand U18821 (N_18821,N_17450,N_17490);
or U18822 (N_18822,N_15260,N_15604);
nand U18823 (N_18823,N_16503,N_15787);
nand U18824 (N_18824,N_16912,N_15470);
nor U18825 (N_18825,N_16837,N_15630);
nand U18826 (N_18826,N_16552,N_17722);
and U18827 (N_18827,N_15334,N_15198);
and U18828 (N_18828,N_15408,N_15588);
nor U18829 (N_18829,N_17609,N_17218);
or U18830 (N_18830,N_17394,N_15913);
nand U18831 (N_18831,N_16084,N_17631);
nand U18832 (N_18832,N_15293,N_16511);
xnor U18833 (N_18833,N_16290,N_16374);
or U18834 (N_18834,N_15868,N_16889);
and U18835 (N_18835,N_15265,N_17685);
or U18836 (N_18836,N_17743,N_16352);
nor U18837 (N_18837,N_16897,N_17740);
nand U18838 (N_18838,N_16281,N_16981);
and U18839 (N_18839,N_16456,N_17641);
nand U18840 (N_18840,N_15638,N_15093);
nand U18841 (N_18841,N_16073,N_15225);
xor U18842 (N_18842,N_17987,N_17409);
nor U18843 (N_18843,N_17564,N_15478);
or U18844 (N_18844,N_15757,N_15271);
nor U18845 (N_18845,N_15499,N_15748);
nor U18846 (N_18846,N_16063,N_15414);
and U18847 (N_18847,N_15727,N_15753);
nor U18848 (N_18848,N_16111,N_15177);
and U18849 (N_18849,N_15105,N_16666);
nand U18850 (N_18850,N_17004,N_16931);
and U18851 (N_18851,N_15326,N_16410);
or U18852 (N_18852,N_15921,N_17376);
nor U18853 (N_18853,N_16537,N_15373);
nand U18854 (N_18854,N_17200,N_16885);
nor U18855 (N_18855,N_16090,N_15462);
and U18856 (N_18856,N_15928,N_16544);
and U18857 (N_18857,N_16789,N_15874);
and U18858 (N_18858,N_15680,N_15207);
nor U18859 (N_18859,N_16527,N_17660);
nor U18860 (N_18860,N_17292,N_16454);
nand U18861 (N_18861,N_16637,N_16446);
xor U18862 (N_18862,N_16162,N_16268);
nand U18863 (N_18863,N_16101,N_17977);
xnor U18864 (N_18864,N_15577,N_16507);
and U18865 (N_18865,N_16913,N_17850);
and U18866 (N_18866,N_17168,N_16012);
nand U18867 (N_18867,N_15389,N_15658);
nor U18868 (N_18868,N_17884,N_15433);
nor U18869 (N_18869,N_17039,N_15235);
nand U18870 (N_18870,N_17672,N_15734);
and U18871 (N_18871,N_16898,N_15115);
nand U18872 (N_18872,N_15123,N_17875);
and U18873 (N_18873,N_17145,N_15132);
xnor U18874 (N_18874,N_16783,N_17482);
nor U18875 (N_18875,N_16199,N_15645);
and U18876 (N_18876,N_16927,N_17322);
and U18877 (N_18877,N_16997,N_15315);
and U18878 (N_18878,N_17510,N_16435);
xnor U18879 (N_18879,N_16088,N_17560);
and U18880 (N_18880,N_16300,N_16583);
xnor U18881 (N_18881,N_17224,N_17507);
nor U18882 (N_18882,N_16541,N_15653);
nor U18883 (N_18883,N_16499,N_15007);
or U18884 (N_18884,N_17264,N_16880);
and U18885 (N_18885,N_17254,N_16936);
and U18886 (N_18886,N_16023,N_16313);
or U18887 (N_18887,N_15871,N_15153);
nor U18888 (N_18888,N_16765,N_15987);
or U18889 (N_18889,N_15487,N_15870);
xnor U18890 (N_18890,N_17148,N_17590);
nand U18891 (N_18891,N_16680,N_17374);
or U18892 (N_18892,N_17833,N_16512);
nor U18893 (N_18893,N_17306,N_15951);
xnor U18894 (N_18894,N_15019,N_15384);
and U18895 (N_18895,N_15399,N_15356);
and U18896 (N_18896,N_16804,N_16695);
and U18897 (N_18897,N_16340,N_16020);
xnor U18898 (N_18898,N_15081,N_16256);
and U18899 (N_18899,N_15516,N_15562);
or U18900 (N_18900,N_15677,N_16690);
or U18901 (N_18901,N_15622,N_15070);
nor U18902 (N_18902,N_17486,N_16483);
nor U18903 (N_18903,N_17256,N_15804);
nand U18904 (N_18904,N_16900,N_16851);
nor U18905 (N_18905,N_15835,N_16036);
nand U18906 (N_18906,N_16387,N_15831);
xnor U18907 (N_18907,N_16873,N_15741);
xnor U18908 (N_18908,N_15982,N_15335);
nor U18909 (N_18909,N_16452,N_17652);
nand U18910 (N_18910,N_16466,N_16381);
nor U18911 (N_18911,N_17532,N_16989);
xnor U18912 (N_18912,N_17890,N_15135);
nor U18913 (N_18913,N_17348,N_16067);
xor U18914 (N_18914,N_16982,N_15752);
and U18915 (N_18915,N_16287,N_16018);
xor U18916 (N_18916,N_16910,N_17902);
xor U18917 (N_18917,N_17702,N_15800);
xnor U18918 (N_18918,N_16065,N_17446);
nor U18919 (N_18919,N_17152,N_17242);
or U18920 (N_18920,N_17147,N_15520);
and U18921 (N_18921,N_15730,N_15675);
xnor U18922 (N_18922,N_15275,N_17984);
or U18923 (N_18923,N_17151,N_15642);
nor U18924 (N_18924,N_15446,N_16022);
xnor U18925 (N_18925,N_17361,N_16669);
or U18926 (N_18926,N_17835,N_15569);
or U18927 (N_18927,N_17274,N_16850);
nor U18928 (N_18928,N_16555,N_15463);
nor U18929 (N_18929,N_16403,N_17752);
nand U18930 (N_18930,N_16598,N_15729);
nor U18931 (N_18931,N_15887,N_17325);
xnor U18932 (N_18932,N_15160,N_16432);
xnor U18933 (N_18933,N_15255,N_15816);
nand U18934 (N_18934,N_15183,N_17707);
or U18935 (N_18935,N_17021,N_17217);
xor U18936 (N_18936,N_15292,N_17465);
or U18937 (N_18937,N_15858,N_16808);
and U18938 (N_18938,N_17387,N_16529);
xnor U18939 (N_18939,N_15640,N_15762);
nor U18940 (N_18940,N_16391,N_15306);
xor U18941 (N_18941,N_15534,N_16191);
nand U18942 (N_18942,N_17949,N_16750);
xor U18943 (N_18943,N_16573,N_16306);
or U18944 (N_18944,N_15812,N_15110);
or U18945 (N_18945,N_15703,N_17330);
nand U18946 (N_18946,N_15161,N_17303);
nand U18947 (N_18947,N_15250,N_15904);
or U18948 (N_18948,N_16372,N_16357);
nor U18949 (N_18949,N_16820,N_16766);
or U18950 (N_18950,N_17404,N_15655);
xnor U18951 (N_18951,N_17742,N_16887);
nor U18952 (N_18952,N_15343,N_15696);
nand U18953 (N_18953,N_15300,N_17149);
xnor U18954 (N_18954,N_17460,N_16408);
and U18955 (N_18955,N_15269,N_15473);
nand U18956 (N_18956,N_15996,N_17595);
xnor U18957 (N_18957,N_15911,N_15736);
or U18958 (N_18958,N_17760,N_16244);
nor U18959 (N_18959,N_15701,N_16202);
or U18960 (N_18960,N_17342,N_17670);
nor U18961 (N_18961,N_16727,N_17137);
or U18962 (N_18962,N_16137,N_17236);
xor U18963 (N_18963,N_16782,N_15629);
nor U18964 (N_18964,N_16428,N_15374);
nand U18965 (N_18965,N_17358,N_17990);
nand U18966 (N_18966,N_17474,N_16650);
nand U18967 (N_18967,N_16396,N_17968);
nand U18968 (N_18968,N_17402,N_16878);
and U18969 (N_18969,N_16693,N_17029);
and U18970 (N_18970,N_17210,N_17382);
xor U18971 (N_18971,N_16694,N_16775);
or U18972 (N_18972,N_15771,N_17037);
nor U18973 (N_18973,N_16958,N_17226);
or U18974 (N_18974,N_17297,N_16059);
nor U18975 (N_18975,N_17893,N_17318);
nor U18976 (N_18976,N_17260,N_15592);
and U18977 (N_18977,N_16426,N_17383);
nor U18978 (N_18978,N_17181,N_17355);
nand U18979 (N_18979,N_16471,N_17922);
or U18980 (N_18980,N_16165,N_15756);
and U18981 (N_18981,N_16206,N_17973);
nor U18982 (N_18982,N_16216,N_15005);
or U18983 (N_18983,N_16596,N_16242);
or U18984 (N_18984,N_17519,N_17538);
or U18985 (N_18985,N_15814,N_15151);
xnor U18986 (N_18986,N_16560,N_17710);
xor U18987 (N_18987,N_16365,N_15261);
nand U18988 (N_18988,N_16279,N_15159);
or U18989 (N_18989,N_17326,N_15339);
and U18990 (N_18990,N_16795,N_16369);
or U18991 (N_18991,N_15950,N_15346);
and U18992 (N_18992,N_15511,N_16670);
nor U18993 (N_18993,N_17428,N_17105);
xnor U18994 (N_18994,N_17904,N_15628);
or U18995 (N_18995,N_15119,N_15296);
xnor U18996 (N_18996,N_15521,N_16759);
nor U18997 (N_18997,N_17847,N_16969);
nand U18998 (N_18998,N_16714,N_16864);
or U18999 (N_18999,N_16303,N_17814);
and U19000 (N_19000,N_16013,N_17918);
or U19001 (N_19001,N_16349,N_16070);
nand U19002 (N_19002,N_16007,N_17232);
nor U19003 (N_19003,N_15761,N_17261);
or U19004 (N_19004,N_17992,N_16526);
nor U19005 (N_19005,N_17528,N_16430);
xnor U19006 (N_19006,N_15323,N_16798);
or U19007 (N_19007,N_17661,N_16091);
nand U19008 (N_19008,N_16732,N_16322);
nand U19009 (N_19009,N_16624,N_16779);
or U19010 (N_19010,N_16235,N_17328);
and U19011 (N_19011,N_15751,N_16315);
nand U19012 (N_19012,N_17451,N_17110);
and U19013 (N_19013,N_16521,N_15214);
or U19014 (N_19014,N_17001,N_17945);
or U19015 (N_19015,N_15352,N_17692);
or U19016 (N_19016,N_15421,N_16480);
xor U19017 (N_19017,N_15882,N_17437);
xor U19018 (N_19018,N_15278,N_16688);
and U19019 (N_19019,N_17777,N_16860);
nor U19020 (N_19020,N_17940,N_17311);
nand U19021 (N_19021,N_16634,N_15853);
and U19022 (N_19022,N_17209,N_17793);
or U19023 (N_19023,N_16932,N_17481);
or U19024 (N_19024,N_17848,N_17504);
nand U19025 (N_19025,N_17929,N_16120);
nor U19026 (N_19026,N_17917,N_16367);
nand U19027 (N_19027,N_17212,N_17795);
and U19028 (N_19028,N_15217,N_15425);
and U19029 (N_19029,N_17193,N_15117);
nand U19030 (N_19030,N_16113,N_17034);
or U19031 (N_19031,N_15687,N_17761);
nand U19032 (N_19032,N_17505,N_15405);
nand U19033 (N_19033,N_16009,N_15836);
and U19034 (N_19034,N_15905,N_16702);
or U19035 (N_19035,N_17076,N_15958);
nor U19036 (N_19036,N_16986,N_15212);
and U19037 (N_19037,N_15348,N_16437);
xnor U19038 (N_19038,N_16849,N_15584);
nor U19039 (N_19039,N_16631,N_16562);
xnor U19040 (N_19040,N_17338,N_15313);
nand U19041 (N_19041,N_16068,N_16353);
nor U19042 (N_19042,N_16267,N_15714);
nor U19043 (N_19043,N_15476,N_15731);
xor U19044 (N_19044,N_15524,N_16000);
xor U19045 (N_19045,N_15678,N_15531);
and U19046 (N_19046,N_15417,N_15724);
nand U19047 (N_19047,N_17194,N_17570);
nor U19048 (N_19048,N_15821,N_15738);
or U19049 (N_19049,N_15360,N_17207);
and U19050 (N_19050,N_15813,N_16547);
or U19051 (N_19051,N_16051,N_16965);
nor U19052 (N_19052,N_15400,N_16149);
nor U19053 (N_19053,N_15082,N_16985);
nor U19054 (N_19054,N_16234,N_16039);
nand U19055 (N_19055,N_16806,N_15899);
nand U19056 (N_19056,N_17093,N_15318);
xor U19057 (N_19057,N_17898,N_16569);
and U19058 (N_19058,N_15195,N_17298);
xnor U19059 (N_19059,N_17734,N_15411);
xor U19060 (N_19060,N_16441,N_16538);
or U19061 (N_19061,N_17524,N_15837);
nor U19062 (N_19062,N_16879,N_17552);
nor U19063 (N_19063,N_17142,N_15155);
or U19064 (N_19064,N_15068,N_17125);
nor U19065 (N_19065,N_17699,N_17844);
nand U19066 (N_19066,N_16050,N_16099);
or U19067 (N_19067,N_16420,N_17123);
or U19068 (N_19068,N_15095,N_15361);
and U19069 (N_19069,N_15788,N_16709);
nand U19070 (N_19070,N_15496,N_15850);
and U19071 (N_19071,N_16116,N_15304);
nand U19072 (N_19072,N_17627,N_15697);
and U19073 (N_19073,N_17403,N_16368);
nor U19074 (N_19074,N_16429,N_16029);
nand U19075 (N_19075,N_16855,N_16725);
xnor U19076 (N_19076,N_17862,N_16787);
nand U19077 (N_19077,N_15359,N_17887);
and U19078 (N_19078,N_17950,N_17909);
and U19079 (N_19079,N_15872,N_15248);
or U19080 (N_19080,N_15585,N_17896);
and U19081 (N_19081,N_15256,N_17502);
xor U19082 (N_19082,N_15603,N_17262);
or U19083 (N_19083,N_15152,N_15615);
and U19084 (N_19084,N_17832,N_17135);
nand U19085 (N_19085,N_16003,N_16125);
nand U19086 (N_19086,N_16047,N_15819);
nand U19087 (N_19087,N_17035,N_17838);
nor U19088 (N_19088,N_15826,N_17302);
nor U19089 (N_19089,N_17836,N_16626);
xnor U19090 (N_19090,N_15202,N_16846);
or U19091 (N_19091,N_15978,N_16316);
and U19092 (N_19092,N_15122,N_15137);
nand U19093 (N_19093,N_16151,N_16755);
nor U19094 (N_19094,N_15200,N_15188);
nor U19095 (N_19095,N_17512,N_16339);
xor U19096 (N_19096,N_17344,N_17924);
and U19097 (N_19097,N_17994,N_15366);
xor U19098 (N_19098,N_16749,N_16385);
xnor U19099 (N_19099,N_15241,N_15594);
xnor U19100 (N_19100,N_16652,N_17558);
or U19101 (N_19101,N_15952,N_16697);
xor U19102 (N_19102,N_17930,N_16841);
or U19103 (N_19103,N_16130,N_16716);
nor U19104 (N_19104,N_16148,N_17663);
and U19105 (N_19105,N_15287,N_15557);
xnor U19106 (N_19106,N_17789,N_15702);
or U19107 (N_19107,N_17189,N_16721);
nand U19108 (N_19108,N_15663,N_17840);
nor U19109 (N_19109,N_17047,N_16345);
nor U19110 (N_19110,N_17040,N_15442);
nand U19111 (N_19111,N_17377,N_16011);
xnor U19112 (N_19112,N_15406,N_15299);
or U19113 (N_19113,N_15652,N_16728);
nand U19114 (N_19114,N_15133,N_17622);
nor U19115 (N_19115,N_17199,N_15617);
xor U19116 (N_19116,N_17308,N_17455);
nor U19117 (N_19117,N_17339,N_16183);
nand U19118 (N_19118,N_16761,N_16320);
xnor U19119 (N_19119,N_15069,N_17390);
nor U19120 (N_19120,N_16042,N_17730);
and U19121 (N_19121,N_16828,N_17265);
and U19122 (N_19122,N_17562,N_15190);
nor U19123 (N_19123,N_17235,N_17518);
and U19124 (N_19124,N_16777,N_17398);
or U19125 (N_19125,N_17900,N_17282);
nor U19126 (N_19126,N_16568,N_17515);
xor U19127 (N_19127,N_15861,N_15547);
xnor U19128 (N_19128,N_16100,N_15321);
or U19129 (N_19129,N_17116,N_17696);
or U19130 (N_19130,N_15529,N_16760);
or U19131 (N_19131,N_16153,N_16717);
or U19132 (N_19132,N_17830,N_16451);
nand U19133 (N_19133,N_15236,N_17132);
nor U19134 (N_19134,N_17701,N_15375);
xnor U19135 (N_19135,N_16390,N_15785);
or U19136 (N_19136,N_15140,N_17927);
and U19137 (N_19137,N_15556,N_17313);
or U19138 (N_19138,N_15715,N_15840);
nor U19139 (N_19139,N_17367,N_15859);
nor U19140 (N_19140,N_15669,N_16341);
xnor U19141 (N_19141,N_16154,N_15071);
and U19142 (N_19142,N_15262,N_17829);
and U19143 (N_19143,N_16475,N_16405);
nor U19144 (N_19144,N_17745,N_15213);
and U19145 (N_19145,N_15320,N_17106);
or U19146 (N_19146,N_16840,N_16834);
or U19147 (N_19147,N_16228,N_17400);
xor U19148 (N_19148,N_17173,N_15708);
nor U19149 (N_19149,N_15964,N_17899);
and U19150 (N_19150,N_17425,N_15566);
nor U19151 (N_19151,N_15501,N_17118);
or U19152 (N_19152,N_16662,N_17563);
xnor U19153 (N_19153,N_15890,N_17545);
or U19154 (N_19154,N_17069,N_16350);
xnor U19155 (N_19155,N_15087,N_17245);
nand U19156 (N_19156,N_15571,N_15664);
or U19157 (N_19157,N_16660,N_15601);
xnor U19158 (N_19158,N_16342,N_15766);
or U19159 (N_19159,N_17011,N_16663);
nand U19160 (N_19160,N_17085,N_15377);
nor U19161 (N_19161,N_16844,N_17601);
or U19162 (N_19162,N_17080,N_17517);
and U19163 (N_19163,N_16425,N_17549);
or U19164 (N_19164,N_15833,N_16444);
or U19165 (N_19165,N_15533,N_15330);
or U19166 (N_19166,N_15627,N_17598);
xnor U19167 (N_19167,N_16881,N_15769);
or U19168 (N_19168,N_17293,N_17712);
and U19169 (N_19169,N_17541,N_16667);
and U19170 (N_19170,N_17375,N_17070);
nor U19171 (N_19171,N_17662,N_16748);
or U19172 (N_19172,N_16045,N_16903);
nand U19173 (N_19173,N_17981,N_16482);
or U19174 (N_19174,N_17360,N_16245);
and U19175 (N_19175,N_16635,N_16375);
and U19176 (N_19176,N_15932,N_17964);
nand U19177 (N_19177,N_15325,N_17568);
xor U19178 (N_19178,N_15713,N_15126);
and U19179 (N_19179,N_17314,N_16776);
xor U19180 (N_19180,N_16970,N_17406);
nand U19181 (N_19181,N_17044,N_16872);
or U19182 (N_19182,N_16616,N_15613);
or U19183 (N_19183,N_16819,N_16044);
and U19184 (N_19184,N_16096,N_15474);
and U19185 (N_19185,N_15626,N_15876);
nand U19186 (N_19186,N_17216,N_16591);
nand U19187 (N_19187,N_15909,N_15945);
or U19188 (N_19188,N_17737,N_16161);
xnor U19189 (N_19189,N_17043,N_15021);
nand U19190 (N_19190,N_17015,N_17483);
and U19191 (N_19191,N_15144,N_17136);
or U19192 (N_19192,N_16546,N_15907);
nand U19193 (N_19193,N_16906,N_15685);
nand U19194 (N_19194,N_17870,N_17633);
nand U19195 (N_19195,N_16935,N_17397);
xor U19196 (N_19196,N_17023,N_15229);
xnor U19197 (N_19197,N_15051,N_17365);
or U19198 (N_19198,N_17975,N_17354);
and U19199 (N_19199,N_15022,N_16762);
xor U19200 (N_19200,N_17211,N_17580);
and U19201 (N_19201,N_16083,N_15838);
xor U19202 (N_19202,N_16227,N_17271);
nand U19203 (N_19203,N_16495,N_15744);
or U19204 (N_19204,N_17782,N_17012);
xor U19205 (N_19205,N_16661,N_17555);
nor U19206 (N_19206,N_17682,N_16416);
nor U19207 (N_19207,N_16557,N_16925);
nand U19208 (N_19208,N_16237,N_17706);
xor U19209 (N_19209,N_16254,N_15922);
xor U19210 (N_19210,N_17576,N_15654);
xnor U19211 (N_19211,N_16813,N_16619);
and U19212 (N_19212,N_17089,N_15358);
nand U19213 (N_19213,N_15166,N_15424);
and U19214 (N_19214,N_17185,N_16298);
nand U19215 (N_19215,N_17369,N_17067);
nand U19216 (N_19216,N_16170,N_17273);
nand U19217 (N_19217,N_16832,N_15130);
xor U19218 (N_19218,N_16585,N_17596);
nand U19219 (N_19219,N_16336,N_16006);
xor U19220 (N_19220,N_16934,N_17527);
or U19221 (N_19221,N_15659,N_15264);
xor U19222 (N_19222,N_17368,N_15259);
and U19223 (N_19223,N_17414,N_17187);
xnor U19224 (N_19224,N_17251,N_17897);
and U19225 (N_19225,N_16334,N_16459);
nor U19226 (N_19226,N_16513,N_17763);
xor U19227 (N_19227,N_17208,N_15223);
nor U19228 (N_19228,N_15864,N_17009);
nand U19229 (N_19229,N_16996,N_16095);
or U19230 (N_19230,N_15668,N_15637);
xor U19231 (N_19231,N_16677,N_16516);
and U19232 (N_19232,N_17104,N_17487);
or U19233 (N_19233,N_16421,N_17405);
nor U19234 (N_19234,N_15854,N_17190);
nor U19235 (N_19235,N_16830,N_16110);
or U19236 (N_19236,N_16656,N_16930);
and U19237 (N_19237,N_17991,N_15782);
xnor U19238 (N_19238,N_17689,N_16911);
nand U19239 (N_19239,N_16431,N_16241);
nor U19240 (N_19240,N_17628,N_17506);
or U19241 (N_19241,N_16117,N_15963);
xor U19242 (N_19242,N_15747,N_15289);
xor U19243 (N_19243,N_16978,N_17905);
xnor U19244 (N_19244,N_17978,N_15542);
and U19245 (N_19245,N_17610,N_16115);
nor U19246 (N_19246,N_16360,N_15451);
and U19247 (N_19247,N_17826,N_15134);
nor U19248 (N_19248,N_16379,N_16414);
nand U19249 (N_19249,N_15931,N_17304);
xor U19250 (N_19250,N_17140,N_15777);
xnor U19251 (N_19251,N_15660,N_15364);
and U19252 (N_19252,N_16536,N_17650);
xor U19253 (N_19253,N_16994,N_16082);
or U19254 (N_19254,N_16079,N_17676);
or U19255 (N_19255,N_17284,N_15215);
and U19256 (N_19256,N_16326,N_17585);
or U19257 (N_19257,N_15427,N_17275);
and U19258 (N_19258,N_17475,N_15578);
and U19259 (N_19259,N_15477,N_15484);
and U19260 (N_19260,N_17798,N_16551);
and U19261 (N_19261,N_17008,N_17201);
or U19262 (N_19262,N_16707,N_17337);
xnor U19263 (N_19263,N_16687,N_17134);
and U19264 (N_19264,N_16875,N_17466);
xor U19265 (N_19265,N_17239,N_17086);
nand U19266 (N_19266,N_15988,N_16921);
and U19267 (N_19267,N_15469,N_15843);
xor U19268 (N_19268,N_15971,N_15139);
and U19269 (N_19269,N_16143,N_16833);
nand U19270 (N_19270,N_15957,N_17019);
nor U19271 (N_19271,N_17024,N_16649);
or U19272 (N_19272,N_16455,N_17138);
nand U19273 (N_19273,N_15823,N_15546);
nor U19274 (N_19274,N_15776,N_16407);
or U19275 (N_19275,N_16586,N_15995);
xnor U19276 (N_19276,N_17791,N_15579);
nand U19277 (N_19277,N_15041,N_17812);
nor U19278 (N_19278,N_16676,N_16305);
or U19279 (N_19279,N_16119,N_17321);
and U19280 (N_19280,N_17054,N_17651);
and U19281 (N_19281,N_16593,N_15357);
nor U19282 (N_19282,N_16874,N_17349);
or U19283 (N_19283,N_16681,N_17448);
and U19284 (N_19284,N_17480,N_17640);
nand U19285 (N_19285,N_17253,N_16433);
or U19286 (N_19286,N_17415,N_17117);
and U19287 (N_19287,N_15355,N_17942);
or U19288 (N_19288,N_15749,N_17543);
xor U19289 (N_19289,N_15054,N_17863);
xor U19290 (N_19290,N_16393,N_16213);
and U19291 (N_19291,N_15386,N_15046);
nor U19292 (N_19292,N_15341,N_15735);
and U19293 (N_19293,N_16017,N_17647);
nand U19294 (N_19294,N_17907,N_17738);
nand U19295 (N_19295,N_16060,N_15825);
nand U19296 (N_19296,N_15733,N_16259);
nor U19297 (N_19297,N_17759,N_16799);
nand U19298 (N_19298,N_17808,N_16304);
and U19299 (N_19299,N_16291,N_17748);
xnor U19300 (N_19300,N_16600,N_15029);
and U19301 (N_19301,N_16745,N_17457);
nand U19302 (N_19302,N_15032,N_15388);
nor U19303 (N_19303,N_16653,N_15750);
nor U19304 (N_19304,N_17713,N_15786);
and U19305 (N_19305,N_17669,N_17386);
and U19306 (N_19306,N_16434,N_15149);
nor U19307 (N_19307,N_17888,N_15129);
nor U19308 (N_19308,N_17452,N_15811);
and U19309 (N_19309,N_16208,N_17948);
and U19310 (N_19310,N_17111,N_15846);
xnor U19311 (N_19311,N_15781,N_15486);
xor U19312 (N_19312,N_15869,N_16571);
and U19313 (N_19313,N_16664,N_17299);
and U19314 (N_19314,N_17657,N_15118);
nor U19315 (N_19315,N_16238,N_15058);
xnor U19316 (N_19316,N_15349,N_16992);
and U19317 (N_19317,N_16233,N_16092);
or U19318 (N_19318,N_17886,N_17389);
xnor U19319 (N_19319,N_16317,N_16058);
or U19320 (N_19320,N_15888,N_15002);
and U19321 (N_19321,N_17373,N_16438);
or U19322 (N_19322,N_16019,N_17961);
xnor U19323 (N_19323,N_16418,N_15312);
and U19324 (N_19324,N_15973,N_17473);
or U19325 (N_19325,N_17100,N_16373);
or U19326 (N_19326,N_17810,N_15936);
or U19327 (N_19327,N_16584,N_16890);
xnor U19328 (N_19328,N_16951,N_15527);
xor U19329 (N_19329,N_15194,N_17718);
nor U19330 (N_19330,N_15507,N_16328);
nand U19331 (N_19331,N_16612,N_16412);
or U19332 (N_19332,N_17516,N_15754);
or U19333 (N_19333,N_15505,N_16743);
nor U19334 (N_19334,N_17310,N_15316);
nand U19335 (N_19335,N_15448,N_17327);
nor U19336 (N_19336,N_16048,N_16257);
nand U19337 (N_19337,N_15085,N_17259);
nor U19338 (N_19338,N_17353,N_17801);
or U19339 (N_19339,N_17316,N_15808);
and U19340 (N_19340,N_16610,N_17049);
nand U19341 (N_19341,N_17449,N_17384);
or U19342 (N_19342,N_16829,N_16272);
nor U19343 (N_19343,N_16672,N_15048);
and U19344 (N_19344,N_15883,N_17018);
nor U19345 (N_19345,N_15378,N_17241);
nand U19346 (N_19346,N_15857,N_15251);
xor U19347 (N_19347,N_15732,N_15018);
nor U19348 (N_19348,N_15620,N_16907);
nand U19349 (N_19349,N_15125,N_16347);
nand U19350 (N_19350,N_15266,N_16742);
nand U19351 (N_19351,N_15038,N_16785);
xor U19352 (N_19352,N_15646,N_17108);
nand U19353 (N_19353,N_16399,N_17771);
xor U19354 (N_19354,N_17953,N_15053);
xnor U19355 (N_19355,N_17340,N_16574);
and U19356 (N_19356,N_17739,N_16797);
nor U19357 (N_19357,N_16424,N_15288);
and U19358 (N_19358,N_15281,N_15114);
nand U19359 (N_19359,N_15517,N_15940);
xnor U19360 (N_19360,N_15270,N_15362);
or U19361 (N_19361,N_15083,N_17797);
xor U19362 (N_19362,N_15108,N_15385);
and U19363 (N_19363,N_16135,N_15572);
nor U19364 (N_19364,N_16632,N_17817);
nor U19365 (N_19365,N_16493,N_17489);
nor U19366 (N_19366,N_17493,N_17017);
and U19367 (N_19367,N_15767,N_16685);
xor U19368 (N_19368,N_17028,N_15211);
or U19369 (N_19369,N_16628,N_16623);
and U19370 (N_19370,N_15233,N_15985);
nand U19371 (N_19371,N_16839,N_17608);
nand U19372 (N_19372,N_17238,N_15395);
xor U19373 (N_19373,N_17161,N_16021);
nand U19374 (N_19374,N_16307,N_17332);
xnor U19375 (N_19375,N_15760,N_16188);
nand U19376 (N_19376,N_15949,N_15772);
nor U19377 (N_19377,N_16618,N_16794);
and U19378 (N_19378,N_17577,N_15468);
or U19379 (N_19379,N_15672,N_17097);
or U19380 (N_19380,N_15073,N_16123);
nor U19381 (N_19381,N_17346,N_16865);
xor U19382 (N_19382,N_17567,N_15704);
xor U19383 (N_19383,N_16180,N_17960);
and U19384 (N_19384,N_15175,N_15599);
nand U19385 (N_19385,N_15401,N_15143);
nand U19386 (N_19386,N_15898,N_15721);
nor U19387 (N_19387,N_15583,N_16816);
nand U19388 (N_19388,N_15197,N_15969);
nor U19389 (N_19389,N_15237,N_16508);
nor U19390 (N_19390,N_17496,N_16297);
or U19391 (N_19391,N_16293,N_17588);
and U19392 (N_19392,N_15024,N_16826);
nand U19393 (N_19393,N_16933,N_16735);
xor U19394 (N_19394,N_17879,N_15933);
nand U19395 (N_19395,N_15483,N_17582);
or U19396 (N_19396,N_16704,N_17775);
nor U19397 (N_19397,N_15683,N_16264);
or U19398 (N_19398,N_17971,N_15779);
nor U19399 (N_19399,N_15066,N_16576);
xor U19400 (N_19400,N_15686,N_15946);
or U19401 (N_19401,N_17408,N_17345);
or U19402 (N_19402,N_16469,N_15609);
or U19403 (N_19403,N_16178,N_15523);
nand U19404 (N_19404,N_16054,N_15154);
xor U19405 (N_19405,N_16382,N_17632);
nor U19406 (N_19406,N_17411,N_16371);
xor U19407 (N_19407,N_15966,N_15662);
xnor U19408 (N_19408,N_15551,N_16648);
or U19409 (N_19409,N_15163,N_17733);
nor U19410 (N_19410,N_17083,N_17883);
or U19411 (N_19411,N_15458,N_17198);
nor U19412 (N_19412,N_17286,N_16942);
xor U19413 (N_19413,N_17578,N_17005);
nor U19414 (N_19414,N_17139,N_16031);
or U19415 (N_19415,N_16112,N_16959);
nor U19416 (N_19416,N_17485,N_17257);
nand U19417 (N_19417,N_16905,N_17865);
nor U19418 (N_19418,N_16080,N_15141);
nand U19419 (N_19419,N_17800,N_17295);
nand U19420 (N_19420,N_17674,N_17586);
and U19421 (N_19421,N_16201,N_15920);
nor U19422 (N_19422,N_17751,N_16174);
nand U19423 (N_19423,N_17645,N_17073);
and U19424 (N_19424,N_16389,N_17126);
or U19425 (N_19425,N_15016,N_17783);
or U19426 (N_19426,N_16266,N_17276);
nand U19427 (N_19427,N_17027,N_15525);
xnor U19428 (N_19428,N_15698,N_17277);
xor U19429 (N_19429,N_16155,N_17229);
nor U19430 (N_19430,N_15014,N_15765);
nor U19431 (N_19431,N_15180,N_15650);
xor U19432 (N_19432,N_17462,N_16647);
xor U19433 (N_19433,N_17268,N_17407);
nand U19434 (N_19434,N_16224,N_16189);
xnor U19435 (N_19435,N_15955,N_16802);
xor U19436 (N_19436,N_16274,N_15409);
xor U19437 (N_19437,N_17064,N_16812);
and U19438 (N_19438,N_15436,N_16468);
or U19439 (N_19439,N_17195,N_17323);
or U19440 (N_19440,N_17347,N_17837);
and U19441 (N_19441,N_15454,N_15608);
nor U19442 (N_19442,N_15522,N_15526);
nand U19443 (N_19443,N_17910,N_16404);
nor U19444 (N_19444,N_16710,N_15929);
xnor U19445 (N_19445,N_16229,N_17656);
or U19446 (N_19446,N_17941,N_15464);
nor U19447 (N_19447,N_17803,N_16754);
nor U19448 (N_19448,N_16737,N_16987);
xor U19449 (N_19449,N_17780,N_16792);
xor U19450 (N_19450,N_15391,N_15116);
and U19451 (N_19451,N_15218,N_17102);
or U19452 (N_19452,N_16489,N_16230);
xor U19453 (N_19453,N_17381,N_16106);
nor U19454 (N_19454,N_15834,N_15394);
nor U19455 (N_19455,N_17958,N_16210);
or U19456 (N_19456,N_15146,N_16114);
and U19457 (N_19457,N_16318,N_15440);
or U19458 (N_19458,N_16646,N_16929);
or U19459 (N_19459,N_17985,N_16458);
xor U19460 (N_19460,N_16436,N_17827);
or U19461 (N_19461,N_15661,N_16417);
and U19462 (N_19462,N_17074,N_15543);
nand U19463 (N_19463,N_17815,N_17521);
and U19464 (N_19464,N_15795,N_17639);
and U19465 (N_19465,N_16498,N_16296);
nand U19466 (N_19466,N_16525,N_16332);
or U19467 (N_19467,N_16877,N_16984);
nand U19468 (N_19468,N_15493,N_16173);
nand U19469 (N_19469,N_17182,N_17671);
nor U19470 (N_19470,N_16152,N_17172);
and U19471 (N_19471,N_17821,N_17501);
nand U19472 (N_19472,N_15100,N_17248);
nor U19473 (N_19473,N_16747,N_15297);
and U19474 (N_19474,N_16730,N_15452);
or U19475 (N_19475,N_17544,N_17861);
nor U19476 (N_19476,N_17937,N_17362);
xnor U19477 (N_19477,N_15994,N_15993);
or U19478 (N_19478,N_17197,N_16980);
or U19479 (N_19479,N_15204,N_17417);
nand U19480 (N_19480,N_15979,N_17334);
or U19481 (N_19481,N_17823,N_15435);
and U19482 (N_19482,N_15099,N_16209);
and U19483 (N_19483,N_16657,N_16330);
or U19484 (N_19484,N_16818,N_17038);
and U19485 (N_19485,N_16496,N_17477);
and U19486 (N_19486,N_15691,N_17616);
or U19487 (N_19487,N_17957,N_17756);
nand U19488 (N_19488,N_17352,N_16219);
and U19489 (N_19489,N_15035,N_16780);
xor U19490 (N_19490,N_16062,N_16445);
or U19491 (N_19491,N_17476,N_16049);
or U19492 (N_19492,N_15820,N_17294);
or U19493 (N_19493,N_16362,N_15286);
and U19494 (N_19494,N_15796,N_15345);
xor U19495 (N_19495,N_16805,N_16142);
or U19496 (N_19496,N_15948,N_17180);
or U19497 (N_19497,N_16895,N_17357);
nor U19498 (N_19498,N_17392,N_16179);
or U19499 (N_19499,N_16542,N_17758);
or U19500 (N_19500,N_15168,N_16811);
xor U19501 (N_19501,N_15566,N_17403);
or U19502 (N_19502,N_15096,N_16780);
or U19503 (N_19503,N_16439,N_15601);
xnor U19504 (N_19504,N_15380,N_17165);
xor U19505 (N_19505,N_16500,N_17315);
or U19506 (N_19506,N_15828,N_16192);
nand U19507 (N_19507,N_15690,N_16363);
nand U19508 (N_19508,N_15511,N_15900);
nor U19509 (N_19509,N_16289,N_17201);
or U19510 (N_19510,N_17849,N_17254);
nand U19511 (N_19511,N_16282,N_16952);
nand U19512 (N_19512,N_16844,N_17456);
and U19513 (N_19513,N_17077,N_17593);
xnor U19514 (N_19514,N_15677,N_15131);
nor U19515 (N_19515,N_16743,N_17458);
xor U19516 (N_19516,N_15100,N_17159);
and U19517 (N_19517,N_17993,N_17173);
nor U19518 (N_19518,N_17056,N_15475);
xor U19519 (N_19519,N_16516,N_16468);
and U19520 (N_19520,N_15610,N_16373);
nor U19521 (N_19521,N_17061,N_17142);
nor U19522 (N_19522,N_17693,N_17171);
xnor U19523 (N_19523,N_16479,N_15106);
nor U19524 (N_19524,N_16377,N_15940);
or U19525 (N_19525,N_15951,N_15425);
and U19526 (N_19526,N_16242,N_16096);
and U19527 (N_19527,N_16347,N_15180);
and U19528 (N_19528,N_17257,N_17660);
and U19529 (N_19529,N_17405,N_16041);
xnor U19530 (N_19530,N_15385,N_16671);
nand U19531 (N_19531,N_17256,N_17774);
nand U19532 (N_19532,N_16206,N_17244);
or U19533 (N_19533,N_17996,N_17738);
xnor U19534 (N_19534,N_16126,N_16722);
or U19535 (N_19535,N_16067,N_17456);
or U19536 (N_19536,N_15709,N_17134);
xor U19537 (N_19537,N_16957,N_17352);
nand U19538 (N_19538,N_16532,N_15045);
and U19539 (N_19539,N_15077,N_16814);
and U19540 (N_19540,N_15614,N_17001);
and U19541 (N_19541,N_15831,N_17959);
nand U19542 (N_19542,N_15628,N_17895);
and U19543 (N_19543,N_16512,N_15655);
nand U19544 (N_19544,N_17285,N_16089);
or U19545 (N_19545,N_17267,N_17438);
nand U19546 (N_19546,N_16754,N_15459);
and U19547 (N_19547,N_15989,N_16700);
nor U19548 (N_19548,N_17823,N_15969);
and U19549 (N_19549,N_17574,N_17371);
nor U19550 (N_19550,N_15057,N_17419);
and U19551 (N_19551,N_16744,N_15371);
xnor U19552 (N_19552,N_17162,N_15848);
and U19553 (N_19553,N_15291,N_17577);
or U19554 (N_19554,N_16900,N_16450);
and U19555 (N_19555,N_17396,N_17288);
and U19556 (N_19556,N_15637,N_17075);
xor U19557 (N_19557,N_16436,N_16090);
nand U19558 (N_19558,N_17876,N_15335);
nand U19559 (N_19559,N_15953,N_15646);
or U19560 (N_19560,N_15490,N_16545);
or U19561 (N_19561,N_16468,N_17588);
and U19562 (N_19562,N_15579,N_17369);
xor U19563 (N_19563,N_17351,N_17589);
nand U19564 (N_19564,N_17946,N_16608);
and U19565 (N_19565,N_16881,N_15015);
xnor U19566 (N_19566,N_16121,N_15340);
nand U19567 (N_19567,N_17697,N_16192);
xor U19568 (N_19568,N_15512,N_16416);
and U19569 (N_19569,N_15070,N_15379);
nand U19570 (N_19570,N_15545,N_17571);
and U19571 (N_19571,N_15447,N_17780);
and U19572 (N_19572,N_17730,N_17152);
nand U19573 (N_19573,N_15404,N_16920);
nand U19574 (N_19574,N_16761,N_15420);
nand U19575 (N_19575,N_16343,N_16883);
or U19576 (N_19576,N_17128,N_16609);
nor U19577 (N_19577,N_16720,N_17590);
or U19578 (N_19578,N_17570,N_16427);
and U19579 (N_19579,N_16705,N_16840);
nand U19580 (N_19580,N_17180,N_15644);
nand U19581 (N_19581,N_16929,N_16651);
xor U19582 (N_19582,N_17905,N_16476);
and U19583 (N_19583,N_17522,N_16988);
nor U19584 (N_19584,N_17841,N_15752);
nand U19585 (N_19585,N_17173,N_16328);
and U19586 (N_19586,N_15405,N_16983);
xnor U19587 (N_19587,N_17086,N_17842);
nor U19588 (N_19588,N_17478,N_16352);
nor U19589 (N_19589,N_17831,N_17564);
or U19590 (N_19590,N_16731,N_17226);
or U19591 (N_19591,N_15489,N_17166);
nand U19592 (N_19592,N_17115,N_17297);
nand U19593 (N_19593,N_15794,N_16225);
nor U19594 (N_19594,N_16127,N_17056);
nor U19595 (N_19595,N_16075,N_17540);
and U19596 (N_19596,N_17202,N_16271);
nor U19597 (N_19597,N_17569,N_15812);
nor U19598 (N_19598,N_16085,N_17686);
nand U19599 (N_19599,N_15633,N_15378);
nand U19600 (N_19600,N_16553,N_15605);
nor U19601 (N_19601,N_17759,N_16049);
and U19602 (N_19602,N_16162,N_17026);
nor U19603 (N_19603,N_16406,N_16896);
xnor U19604 (N_19604,N_15176,N_17866);
xor U19605 (N_19605,N_16092,N_16613);
nor U19606 (N_19606,N_15746,N_17668);
nor U19607 (N_19607,N_16683,N_15281);
nor U19608 (N_19608,N_17765,N_15722);
nor U19609 (N_19609,N_17631,N_17604);
xor U19610 (N_19610,N_15092,N_17329);
nor U19611 (N_19611,N_17496,N_17251);
xor U19612 (N_19612,N_15357,N_16475);
nand U19613 (N_19613,N_15647,N_16524);
nor U19614 (N_19614,N_16017,N_17050);
and U19615 (N_19615,N_16064,N_17384);
or U19616 (N_19616,N_15891,N_16226);
nor U19617 (N_19617,N_16298,N_17481);
nor U19618 (N_19618,N_17875,N_17957);
nand U19619 (N_19619,N_15010,N_16253);
and U19620 (N_19620,N_16452,N_17061);
and U19621 (N_19621,N_17126,N_17373);
nor U19622 (N_19622,N_17339,N_15964);
nor U19623 (N_19623,N_16726,N_15840);
or U19624 (N_19624,N_17184,N_17796);
and U19625 (N_19625,N_16088,N_17592);
or U19626 (N_19626,N_17442,N_16771);
nor U19627 (N_19627,N_16246,N_15508);
nor U19628 (N_19628,N_16277,N_15319);
or U19629 (N_19629,N_17134,N_16825);
or U19630 (N_19630,N_16212,N_16900);
xnor U19631 (N_19631,N_16696,N_16745);
nor U19632 (N_19632,N_17403,N_17463);
nand U19633 (N_19633,N_16575,N_17545);
nand U19634 (N_19634,N_17389,N_16778);
xor U19635 (N_19635,N_16464,N_15158);
nor U19636 (N_19636,N_17864,N_17167);
nor U19637 (N_19637,N_15262,N_17661);
nand U19638 (N_19638,N_16296,N_15166);
and U19639 (N_19639,N_16837,N_17068);
nand U19640 (N_19640,N_17257,N_17695);
xor U19641 (N_19641,N_16878,N_16345);
or U19642 (N_19642,N_16382,N_17333);
xnor U19643 (N_19643,N_15832,N_15969);
nor U19644 (N_19644,N_16125,N_16839);
nand U19645 (N_19645,N_16882,N_16219);
and U19646 (N_19646,N_16471,N_17770);
xnor U19647 (N_19647,N_15260,N_17955);
or U19648 (N_19648,N_17961,N_15797);
nor U19649 (N_19649,N_17658,N_16531);
nor U19650 (N_19650,N_16453,N_16708);
nor U19651 (N_19651,N_17863,N_17053);
and U19652 (N_19652,N_15285,N_16196);
and U19653 (N_19653,N_16365,N_15616);
and U19654 (N_19654,N_16649,N_17862);
xor U19655 (N_19655,N_15367,N_16266);
or U19656 (N_19656,N_16243,N_16203);
xor U19657 (N_19657,N_16874,N_16273);
xnor U19658 (N_19658,N_15384,N_16402);
nor U19659 (N_19659,N_16391,N_17307);
or U19660 (N_19660,N_15744,N_15727);
or U19661 (N_19661,N_15732,N_15749);
and U19662 (N_19662,N_16411,N_17389);
nand U19663 (N_19663,N_15340,N_17265);
or U19664 (N_19664,N_15834,N_17382);
nor U19665 (N_19665,N_16769,N_16422);
and U19666 (N_19666,N_16346,N_16701);
xnor U19667 (N_19667,N_17770,N_15835);
nand U19668 (N_19668,N_15824,N_17256);
nand U19669 (N_19669,N_16210,N_16377);
nor U19670 (N_19670,N_15538,N_15910);
nand U19671 (N_19671,N_16003,N_15356);
or U19672 (N_19672,N_16804,N_17204);
and U19673 (N_19673,N_17609,N_15354);
and U19674 (N_19674,N_17089,N_17610);
and U19675 (N_19675,N_15921,N_16224);
nand U19676 (N_19676,N_17695,N_15304);
or U19677 (N_19677,N_15663,N_15783);
nand U19678 (N_19678,N_15545,N_16344);
nand U19679 (N_19679,N_16583,N_16276);
xnor U19680 (N_19680,N_15431,N_17584);
nand U19681 (N_19681,N_17578,N_16162);
and U19682 (N_19682,N_15869,N_17075);
nor U19683 (N_19683,N_16061,N_16393);
xor U19684 (N_19684,N_15657,N_16900);
xor U19685 (N_19685,N_15268,N_15279);
nor U19686 (N_19686,N_15690,N_15043);
nand U19687 (N_19687,N_15321,N_15645);
nand U19688 (N_19688,N_15878,N_15372);
nand U19689 (N_19689,N_16972,N_16105);
nand U19690 (N_19690,N_15327,N_15818);
or U19691 (N_19691,N_16648,N_16863);
xor U19692 (N_19692,N_17739,N_17224);
and U19693 (N_19693,N_17186,N_16500);
nand U19694 (N_19694,N_15683,N_17550);
nor U19695 (N_19695,N_15607,N_16115);
nor U19696 (N_19696,N_16244,N_16197);
xnor U19697 (N_19697,N_17282,N_15136);
xnor U19698 (N_19698,N_16510,N_16511);
or U19699 (N_19699,N_17685,N_16282);
or U19700 (N_19700,N_17003,N_17480);
nand U19701 (N_19701,N_17440,N_17510);
and U19702 (N_19702,N_16844,N_15425);
and U19703 (N_19703,N_17603,N_16820);
nand U19704 (N_19704,N_15580,N_16962);
nand U19705 (N_19705,N_17010,N_17529);
nand U19706 (N_19706,N_15798,N_17800);
and U19707 (N_19707,N_16659,N_16709);
or U19708 (N_19708,N_17564,N_16190);
or U19709 (N_19709,N_17664,N_15615);
nand U19710 (N_19710,N_15348,N_15534);
and U19711 (N_19711,N_15333,N_17058);
and U19712 (N_19712,N_15762,N_16905);
nand U19713 (N_19713,N_15677,N_15069);
and U19714 (N_19714,N_15810,N_15799);
xnor U19715 (N_19715,N_16273,N_15976);
and U19716 (N_19716,N_16756,N_16925);
and U19717 (N_19717,N_15529,N_16240);
and U19718 (N_19718,N_16771,N_16072);
xor U19719 (N_19719,N_17610,N_16895);
and U19720 (N_19720,N_16173,N_15957);
xnor U19721 (N_19721,N_17685,N_16102);
nor U19722 (N_19722,N_15189,N_15139);
nor U19723 (N_19723,N_15344,N_16815);
xor U19724 (N_19724,N_16998,N_17522);
xnor U19725 (N_19725,N_15478,N_17503);
xnor U19726 (N_19726,N_15973,N_15782);
or U19727 (N_19727,N_15803,N_17097);
xnor U19728 (N_19728,N_16469,N_17969);
xor U19729 (N_19729,N_17117,N_17572);
and U19730 (N_19730,N_17970,N_17091);
nand U19731 (N_19731,N_16812,N_17235);
and U19732 (N_19732,N_17459,N_15949);
nor U19733 (N_19733,N_17573,N_16731);
or U19734 (N_19734,N_17599,N_17971);
nor U19735 (N_19735,N_17784,N_17498);
nand U19736 (N_19736,N_17444,N_15519);
and U19737 (N_19737,N_17682,N_15761);
nand U19738 (N_19738,N_17571,N_15961);
xnor U19739 (N_19739,N_17725,N_15292);
and U19740 (N_19740,N_17725,N_16470);
and U19741 (N_19741,N_15647,N_15108);
and U19742 (N_19742,N_15736,N_15456);
nor U19743 (N_19743,N_17947,N_15421);
or U19744 (N_19744,N_15573,N_15982);
or U19745 (N_19745,N_16929,N_15376);
xor U19746 (N_19746,N_17845,N_15318);
nand U19747 (N_19747,N_15100,N_15062);
nand U19748 (N_19748,N_17922,N_15067);
nand U19749 (N_19749,N_17362,N_15327);
xor U19750 (N_19750,N_16457,N_16138);
and U19751 (N_19751,N_17912,N_16888);
xor U19752 (N_19752,N_17425,N_17804);
or U19753 (N_19753,N_16511,N_17516);
nand U19754 (N_19754,N_15817,N_16718);
nor U19755 (N_19755,N_15862,N_16087);
or U19756 (N_19756,N_16607,N_15943);
nand U19757 (N_19757,N_15799,N_17242);
and U19758 (N_19758,N_17857,N_15081);
and U19759 (N_19759,N_16387,N_15169);
nor U19760 (N_19760,N_16551,N_17533);
xnor U19761 (N_19761,N_15096,N_15684);
xor U19762 (N_19762,N_16122,N_15302);
and U19763 (N_19763,N_15900,N_16846);
nand U19764 (N_19764,N_15609,N_15391);
xnor U19765 (N_19765,N_17536,N_17740);
nand U19766 (N_19766,N_15815,N_17077);
and U19767 (N_19767,N_17444,N_17659);
xnor U19768 (N_19768,N_16883,N_17810);
and U19769 (N_19769,N_15654,N_17712);
or U19770 (N_19770,N_15152,N_16075);
xor U19771 (N_19771,N_17329,N_16946);
nand U19772 (N_19772,N_17912,N_15537);
xnor U19773 (N_19773,N_16606,N_15227);
and U19774 (N_19774,N_17186,N_15480);
or U19775 (N_19775,N_15692,N_17219);
xnor U19776 (N_19776,N_17350,N_17478);
nand U19777 (N_19777,N_17144,N_16838);
xnor U19778 (N_19778,N_15574,N_15765);
or U19779 (N_19779,N_16710,N_17648);
nand U19780 (N_19780,N_16954,N_16042);
nor U19781 (N_19781,N_17159,N_16756);
or U19782 (N_19782,N_16262,N_17723);
and U19783 (N_19783,N_17935,N_17707);
xnor U19784 (N_19784,N_16372,N_17409);
or U19785 (N_19785,N_16851,N_16439);
nor U19786 (N_19786,N_16307,N_16251);
or U19787 (N_19787,N_15784,N_16880);
nor U19788 (N_19788,N_17713,N_16783);
nand U19789 (N_19789,N_17625,N_16725);
nor U19790 (N_19790,N_16740,N_15557);
or U19791 (N_19791,N_15070,N_17757);
nand U19792 (N_19792,N_16775,N_15539);
nand U19793 (N_19793,N_16834,N_17681);
xor U19794 (N_19794,N_16283,N_15606);
or U19795 (N_19795,N_17490,N_17476);
and U19796 (N_19796,N_15661,N_15259);
or U19797 (N_19797,N_17758,N_17703);
or U19798 (N_19798,N_16824,N_17093);
xnor U19799 (N_19799,N_15555,N_15444);
or U19800 (N_19800,N_17294,N_16005);
or U19801 (N_19801,N_15127,N_17259);
nor U19802 (N_19802,N_15614,N_16465);
nand U19803 (N_19803,N_16414,N_15443);
xor U19804 (N_19804,N_16859,N_17945);
nand U19805 (N_19805,N_16523,N_16938);
and U19806 (N_19806,N_17086,N_17188);
and U19807 (N_19807,N_17949,N_16388);
nand U19808 (N_19808,N_15654,N_16487);
xnor U19809 (N_19809,N_15595,N_17501);
xor U19810 (N_19810,N_15717,N_17362);
xor U19811 (N_19811,N_16194,N_15577);
nor U19812 (N_19812,N_15333,N_15469);
or U19813 (N_19813,N_15933,N_15551);
xnor U19814 (N_19814,N_15505,N_17396);
xnor U19815 (N_19815,N_17866,N_16195);
nor U19816 (N_19816,N_16092,N_15924);
xor U19817 (N_19817,N_15008,N_15591);
nand U19818 (N_19818,N_15036,N_15939);
nand U19819 (N_19819,N_17968,N_17502);
xor U19820 (N_19820,N_15897,N_16118);
or U19821 (N_19821,N_16936,N_15306);
nor U19822 (N_19822,N_17344,N_17118);
xor U19823 (N_19823,N_15914,N_17620);
and U19824 (N_19824,N_16924,N_17499);
xnor U19825 (N_19825,N_17374,N_17029);
nand U19826 (N_19826,N_17485,N_15583);
nand U19827 (N_19827,N_17180,N_17305);
nor U19828 (N_19828,N_17880,N_16634);
nand U19829 (N_19829,N_15205,N_16698);
or U19830 (N_19830,N_17212,N_16607);
nand U19831 (N_19831,N_17678,N_17423);
nor U19832 (N_19832,N_16160,N_16864);
nand U19833 (N_19833,N_15843,N_17211);
or U19834 (N_19834,N_16164,N_17376);
and U19835 (N_19835,N_15721,N_15318);
or U19836 (N_19836,N_16852,N_15988);
nor U19837 (N_19837,N_17670,N_16230);
nand U19838 (N_19838,N_17481,N_17453);
xor U19839 (N_19839,N_16501,N_17860);
nor U19840 (N_19840,N_15939,N_16229);
or U19841 (N_19841,N_16633,N_15051);
xor U19842 (N_19842,N_16555,N_17462);
or U19843 (N_19843,N_16435,N_17750);
xor U19844 (N_19844,N_16961,N_17093);
or U19845 (N_19845,N_15067,N_16254);
nor U19846 (N_19846,N_15571,N_17288);
nor U19847 (N_19847,N_16279,N_17983);
or U19848 (N_19848,N_17439,N_15489);
nand U19849 (N_19849,N_15391,N_17494);
and U19850 (N_19850,N_15749,N_17858);
nor U19851 (N_19851,N_16860,N_16911);
nand U19852 (N_19852,N_17611,N_17186);
xnor U19853 (N_19853,N_15441,N_17093);
nand U19854 (N_19854,N_17766,N_16151);
nor U19855 (N_19855,N_15619,N_16666);
xor U19856 (N_19856,N_15918,N_17663);
nor U19857 (N_19857,N_16731,N_15865);
nand U19858 (N_19858,N_17485,N_16367);
xor U19859 (N_19859,N_15945,N_17936);
and U19860 (N_19860,N_17327,N_16515);
or U19861 (N_19861,N_15440,N_15575);
nor U19862 (N_19862,N_17385,N_17258);
xor U19863 (N_19863,N_15324,N_16944);
nand U19864 (N_19864,N_15292,N_16610);
or U19865 (N_19865,N_15397,N_17479);
and U19866 (N_19866,N_15458,N_15698);
and U19867 (N_19867,N_17073,N_17066);
nor U19868 (N_19868,N_17653,N_15397);
and U19869 (N_19869,N_16089,N_17464);
nand U19870 (N_19870,N_17372,N_16212);
xor U19871 (N_19871,N_15093,N_15387);
nand U19872 (N_19872,N_17797,N_16359);
or U19873 (N_19873,N_16663,N_15505);
or U19874 (N_19874,N_16858,N_16868);
or U19875 (N_19875,N_16517,N_15239);
nor U19876 (N_19876,N_16093,N_16541);
and U19877 (N_19877,N_17592,N_15294);
or U19878 (N_19878,N_15480,N_15980);
and U19879 (N_19879,N_17222,N_15696);
and U19880 (N_19880,N_17319,N_16462);
or U19881 (N_19881,N_17435,N_16310);
and U19882 (N_19882,N_15247,N_15246);
xor U19883 (N_19883,N_17688,N_17556);
and U19884 (N_19884,N_16416,N_17358);
and U19885 (N_19885,N_16014,N_16552);
nor U19886 (N_19886,N_15080,N_16445);
or U19887 (N_19887,N_15030,N_15069);
or U19888 (N_19888,N_16755,N_17575);
or U19889 (N_19889,N_17490,N_15531);
and U19890 (N_19890,N_16629,N_16524);
xor U19891 (N_19891,N_15342,N_15250);
nand U19892 (N_19892,N_16371,N_17228);
and U19893 (N_19893,N_17195,N_16973);
nand U19894 (N_19894,N_16754,N_16212);
and U19895 (N_19895,N_17680,N_16849);
xor U19896 (N_19896,N_16665,N_17441);
nor U19897 (N_19897,N_16137,N_15712);
nand U19898 (N_19898,N_17256,N_15684);
and U19899 (N_19899,N_16723,N_16300);
and U19900 (N_19900,N_16287,N_16373);
or U19901 (N_19901,N_16717,N_15809);
nor U19902 (N_19902,N_17275,N_15101);
nor U19903 (N_19903,N_17100,N_15953);
nor U19904 (N_19904,N_15215,N_15719);
and U19905 (N_19905,N_17391,N_16812);
and U19906 (N_19906,N_16188,N_17317);
and U19907 (N_19907,N_17287,N_15928);
nor U19908 (N_19908,N_15700,N_17149);
and U19909 (N_19909,N_17088,N_16915);
nand U19910 (N_19910,N_16588,N_16380);
nand U19911 (N_19911,N_17823,N_17530);
xnor U19912 (N_19912,N_15439,N_16705);
nand U19913 (N_19913,N_16733,N_17400);
nand U19914 (N_19914,N_17026,N_15674);
and U19915 (N_19915,N_16199,N_16257);
xnor U19916 (N_19916,N_16987,N_16218);
nand U19917 (N_19917,N_16072,N_17911);
nor U19918 (N_19918,N_15762,N_15867);
or U19919 (N_19919,N_16762,N_17409);
xor U19920 (N_19920,N_15438,N_17032);
and U19921 (N_19921,N_17484,N_17199);
and U19922 (N_19922,N_16786,N_15620);
or U19923 (N_19923,N_17053,N_17272);
nand U19924 (N_19924,N_16575,N_16421);
or U19925 (N_19925,N_15203,N_16616);
xor U19926 (N_19926,N_15666,N_15066);
or U19927 (N_19927,N_15612,N_16834);
nand U19928 (N_19928,N_15370,N_16618);
xnor U19929 (N_19929,N_17580,N_15639);
or U19930 (N_19930,N_17306,N_16832);
nand U19931 (N_19931,N_16651,N_16084);
or U19932 (N_19932,N_17701,N_15716);
nor U19933 (N_19933,N_16444,N_16031);
nand U19934 (N_19934,N_16636,N_17773);
or U19935 (N_19935,N_15328,N_17177);
or U19936 (N_19936,N_17904,N_16734);
nor U19937 (N_19937,N_16506,N_16864);
nand U19938 (N_19938,N_15979,N_17379);
nand U19939 (N_19939,N_17099,N_15862);
and U19940 (N_19940,N_15004,N_15871);
or U19941 (N_19941,N_15966,N_15707);
or U19942 (N_19942,N_16388,N_17610);
or U19943 (N_19943,N_16092,N_17488);
and U19944 (N_19944,N_16185,N_16119);
nor U19945 (N_19945,N_17894,N_17118);
or U19946 (N_19946,N_15900,N_17518);
and U19947 (N_19947,N_17182,N_15981);
and U19948 (N_19948,N_17987,N_17819);
xor U19949 (N_19949,N_16453,N_17297);
and U19950 (N_19950,N_16893,N_16134);
xor U19951 (N_19951,N_17902,N_17186);
nand U19952 (N_19952,N_17176,N_15965);
xnor U19953 (N_19953,N_15615,N_15876);
nor U19954 (N_19954,N_15231,N_15423);
or U19955 (N_19955,N_16321,N_15894);
nor U19956 (N_19956,N_16283,N_17537);
and U19957 (N_19957,N_15548,N_15495);
xnor U19958 (N_19958,N_17515,N_16733);
nand U19959 (N_19959,N_16230,N_16812);
nor U19960 (N_19960,N_16703,N_16883);
xor U19961 (N_19961,N_15738,N_15521);
or U19962 (N_19962,N_16808,N_15428);
nand U19963 (N_19963,N_16048,N_16489);
or U19964 (N_19964,N_17565,N_15823);
and U19965 (N_19965,N_15160,N_17519);
and U19966 (N_19966,N_16159,N_15048);
nand U19967 (N_19967,N_15044,N_15032);
and U19968 (N_19968,N_15237,N_15089);
nor U19969 (N_19969,N_17087,N_17646);
and U19970 (N_19970,N_17983,N_16490);
or U19971 (N_19971,N_17701,N_17615);
nand U19972 (N_19972,N_16014,N_15332);
or U19973 (N_19973,N_16642,N_16014);
or U19974 (N_19974,N_16289,N_17241);
nor U19975 (N_19975,N_15984,N_16817);
or U19976 (N_19976,N_15066,N_15876);
or U19977 (N_19977,N_17080,N_17351);
nor U19978 (N_19978,N_16074,N_15460);
and U19979 (N_19979,N_16935,N_16457);
or U19980 (N_19980,N_16316,N_16038);
nor U19981 (N_19981,N_16564,N_15855);
or U19982 (N_19982,N_15319,N_17951);
nor U19983 (N_19983,N_17790,N_16358);
nand U19984 (N_19984,N_15608,N_15308);
nand U19985 (N_19985,N_17102,N_17821);
nor U19986 (N_19986,N_15797,N_15736);
nand U19987 (N_19987,N_15548,N_17007);
nor U19988 (N_19988,N_16858,N_15574);
xnor U19989 (N_19989,N_15753,N_16522);
or U19990 (N_19990,N_16600,N_15314);
nand U19991 (N_19991,N_15084,N_15695);
and U19992 (N_19992,N_16558,N_16961);
nor U19993 (N_19993,N_17931,N_17371);
xor U19994 (N_19994,N_16936,N_15622);
and U19995 (N_19995,N_16608,N_16441);
and U19996 (N_19996,N_16840,N_15180);
xnor U19997 (N_19997,N_17697,N_17355);
nor U19998 (N_19998,N_16887,N_16739);
xor U19999 (N_19999,N_15792,N_16272);
and U20000 (N_20000,N_16570,N_17580);
nand U20001 (N_20001,N_16420,N_17879);
xnor U20002 (N_20002,N_15208,N_15290);
and U20003 (N_20003,N_17060,N_16467);
and U20004 (N_20004,N_16345,N_15688);
and U20005 (N_20005,N_16507,N_17277);
xor U20006 (N_20006,N_17903,N_17080);
or U20007 (N_20007,N_17853,N_15292);
and U20008 (N_20008,N_15224,N_17085);
xnor U20009 (N_20009,N_15245,N_16338);
and U20010 (N_20010,N_17656,N_17958);
xnor U20011 (N_20011,N_15989,N_17240);
xnor U20012 (N_20012,N_16392,N_15730);
or U20013 (N_20013,N_15255,N_17314);
nand U20014 (N_20014,N_16591,N_17662);
nand U20015 (N_20015,N_17332,N_16859);
nand U20016 (N_20016,N_15481,N_16048);
nand U20017 (N_20017,N_16312,N_15937);
nor U20018 (N_20018,N_15254,N_17980);
nand U20019 (N_20019,N_17948,N_17781);
and U20020 (N_20020,N_16042,N_15115);
nor U20021 (N_20021,N_15548,N_15552);
nand U20022 (N_20022,N_15748,N_17627);
nand U20023 (N_20023,N_15597,N_16418);
nor U20024 (N_20024,N_16774,N_16237);
nor U20025 (N_20025,N_15509,N_17008);
nand U20026 (N_20026,N_17042,N_17521);
nor U20027 (N_20027,N_16914,N_15710);
nand U20028 (N_20028,N_16758,N_17265);
xnor U20029 (N_20029,N_15733,N_17646);
nor U20030 (N_20030,N_15087,N_15447);
nand U20031 (N_20031,N_17041,N_17303);
xnor U20032 (N_20032,N_17632,N_15812);
nor U20033 (N_20033,N_15040,N_15518);
or U20034 (N_20034,N_17027,N_17959);
xor U20035 (N_20035,N_16272,N_16321);
nand U20036 (N_20036,N_15938,N_16940);
and U20037 (N_20037,N_15630,N_17075);
nor U20038 (N_20038,N_17026,N_16852);
and U20039 (N_20039,N_17158,N_16593);
nand U20040 (N_20040,N_17796,N_15430);
nor U20041 (N_20041,N_16261,N_17949);
and U20042 (N_20042,N_16718,N_15246);
or U20043 (N_20043,N_15051,N_16768);
and U20044 (N_20044,N_17724,N_15153);
nor U20045 (N_20045,N_16156,N_16930);
and U20046 (N_20046,N_16019,N_17295);
and U20047 (N_20047,N_15436,N_15492);
nand U20048 (N_20048,N_15986,N_16006);
or U20049 (N_20049,N_16969,N_15726);
nand U20050 (N_20050,N_15083,N_15023);
nor U20051 (N_20051,N_15365,N_15128);
nor U20052 (N_20052,N_16560,N_17701);
nor U20053 (N_20053,N_16755,N_17308);
and U20054 (N_20054,N_17288,N_15522);
nand U20055 (N_20055,N_16199,N_15277);
nor U20056 (N_20056,N_16295,N_15342);
or U20057 (N_20057,N_15367,N_15240);
xor U20058 (N_20058,N_15194,N_16719);
nand U20059 (N_20059,N_16137,N_16208);
nand U20060 (N_20060,N_17147,N_15568);
nand U20061 (N_20061,N_15296,N_16603);
xor U20062 (N_20062,N_15884,N_17202);
and U20063 (N_20063,N_16233,N_16937);
and U20064 (N_20064,N_16733,N_15385);
and U20065 (N_20065,N_17465,N_15225);
or U20066 (N_20066,N_16614,N_17177);
or U20067 (N_20067,N_17832,N_17012);
and U20068 (N_20068,N_17578,N_16223);
and U20069 (N_20069,N_17422,N_17599);
nand U20070 (N_20070,N_17294,N_17847);
xnor U20071 (N_20071,N_17123,N_15206);
xnor U20072 (N_20072,N_16785,N_16934);
nand U20073 (N_20073,N_16141,N_16463);
xnor U20074 (N_20074,N_15576,N_15906);
xor U20075 (N_20075,N_16098,N_16703);
or U20076 (N_20076,N_17750,N_15694);
or U20077 (N_20077,N_15879,N_17309);
xor U20078 (N_20078,N_15039,N_17535);
and U20079 (N_20079,N_15987,N_16486);
nand U20080 (N_20080,N_15745,N_16541);
xnor U20081 (N_20081,N_16601,N_17106);
xnor U20082 (N_20082,N_15564,N_15969);
or U20083 (N_20083,N_17569,N_17503);
nand U20084 (N_20084,N_17889,N_15275);
nand U20085 (N_20085,N_17756,N_15190);
or U20086 (N_20086,N_16927,N_17102);
or U20087 (N_20087,N_16099,N_16031);
nor U20088 (N_20088,N_17439,N_15947);
nor U20089 (N_20089,N_15161,N_15841);
nor U20090 (N_20090,N_15055,N_15456);
nor U20091 (N_20091,N_17724,N_17364);
nor U20092 (N_20092,N_17593,N_15044);
nor U20093 (N_20093,N_15879,N_17293);
and U20094 (N_20094,N_15885,N_15945);
nand U20095 (N_20095,N_15091,N_15828);
nand U20096 (N_20096,N_16807,N_16371);
xor U20097 (N_20097,N_15427,N_16779);
or U20098 (N_20098,N_16127,N_16595);
or U20099 (N_20099,N_15529,N_16296);
xnor U20100 (N_20100,N_17617,N_16879);
nor U20101 (N_20101,N_17322,N_16570);
and U20102 (N_20102,N_15977,N_15241);
nand U20103 (N_20103,N_15081,N_16072);
xor U20104 (N_20104,N_16354,N_17096);
nand U20105 (N_20105,N_16016,N_15659);
or U20106 (N_20106,N_15338,N_16811);
and U20107 (N_20107,N_15341,N_16305);
nor U20108 (N_20108,N_16916,N_17496);
nor U20109 (N_20109,N_15758,N_17725);
or U20110 (N_20110,N_17438,N_15513);
or U20111 (N_20111,N_16730,N_17064);
nand U20112 (N_20112,N_17129,N_16378);
or U20113 (N_20113,N_15774,N_17049);
and U20114 (N_20114,N_15795,N_16697);
nor U20115 (N_20115,N_17529,N_16489);
nand U20116 (N_20116,N_16703,N_16328);
nand U20117 (N_20117,N_15331,N_16202);
nand U20118 (N_20118,N_17602,N_15390);
or U20119 (N_20119,N_17372,N_15310);
or U20120 (N_20120,N_17669,N_16446);
nor U20121 (N_20121,N_15917,N_15967);
xnor U20122 (N_20122,N_16864,N_16335);
xnor U20123 (N_20123,N_15352,N_16303);
xnor U20124 (N_20124,N_16375,N_17072);
or U20125 (N_20125,N_15343,N_17558);
nor U20126 (N_20126,N_15952,N_16742);
and U20127 (N_20127,N_16847,N_15996);
or U20128 (N_20128,N_16815,N_16301);
or U20129 (N_20129,N_17270,N_17356);
or U20130 (N_20130,N_17629,N_16254);
and U20131 (N_20131,N_15125,N_15838);
nor U20132 (N_20132,N_16408,N_17696);
and U20133 (N_20133,N_16538,N_17230);
xor U20134 (N_20134,N_16514,N_17420);
nor U20135 (N_20135,N_17701,N_15398);
xor U20136 (N_20136,N_15470,N_15608);
nor U20137 (N_20137,N_16555,N_15834);
or U20138 (N_20138,N_15908,N_15752);
or U20139 (N_20139,N_15928,N_15576);
or U20140 (N_20140,N_17791,N_16147);
and U20141 (N_20141,N_16407,N_16165);
nand U20142 (N_20142,N_15442,N_15593);
xor U20143 (N_20143,N_15737,N_17881);
nor U20144 (N_20144,N_17787,N_17197);
nand U20145 (N_20145,N_15016,N_16166);
nor U20146 (N_20146,N_17206,N_17653);
nand U20147 (N_20147,N_15652,N_16544);
nand U20148 (N_20148,N_16824,N_15468);
or U20149 (N_20149,N_15161,N_17683);
or U20150 (N_20150,N_16086,N_15948);
or U20151 (N_20151,N_17919,N_15506);
nand U20152 (N_20152,N_17126,N_17908);
nand U20153 (N_20153,N_16648,N_16510);
xor U20154 (N_20154,N_15356,N_16450);
and U20155 (N_20155,N_16197,N_15255);
nor U20156 (N_20156,N_15577,N_17922);
xor U20157 (N_20157,N_17013,N_15683);
nand U20158 (N_20158,N_16737,N_17345);
and U20159 (N_20159,N_17843,N_17743);
nor U20160 (N_20160,N_15526,N_16548);
nor U20161 (N_20161,N_15343,N_15437);
xnor U20162 (N_20162,N_17132,N_17794);
or U20163 (N_20163,N_16113,N_16494);
nand U20164 (N_20164,N_17451,N_17326);
and U20165 (N_20165,N_15758,N_16192);
xnor U20166 (N_20166,N_16043,N_16412);
or U20167 (N_20167,N_16220,N_16707);
xor U20168 (N_20168,N_15765,N_16968);
xnor U20169 (N_20169,N_16109,N_17255);
or U20170 (N_20170,N_16494,N_15630);
nor U20171 (N_20171,N_15785,N_17114);
nand U20172 (N_20172,N_15077,N_15824);
or U20173 (N_20173,N_15216,N_15388);
or U20174 (N_20174,N_17529,N_17710);
nand U20175 (N_20175,N_15800,N_15972);
or U20176 (N_20176,N_16732,N_17035);
nand U20177 (N_20177,N_17548,N_16260);
nor U20178 (N_20178,N_15498,N_17908);
and U20179 (N_20179,N_16292,N_16549);
and U20180 (N_20180,N_15552,N_16143);
nand U20181 (N_20181,N_15259,N_15171);
and U20182 (N_20182,N_15823,N_16243);
or U20183 (N_20183,N_17165,N_17548);
and U20184 (N_20184,N_15987,N_17416);
or U20185 (N_20185,N_17490,N_15186);
nand U20186 (N_20186,N_15647,N_17329);
nand U20187 (N_20187,N_15495,N_17641);
or U20188 (N_20188,N_17130,N_17768);
or U20189 (N_20189,N_16597,N_17837);
or U20190 (N_20190,N_17434,N_16991);
nor U20191 (N_20191,N_16259,N_16998);
xor U20192 (N_20192,N_15488,N_15092);
xor U20193 (N_20193,N_16645,N_16890);
nor U20194 (N_20194,N_17940,N_17211);
nand U20195 (N_20195,N_15512,N_15366);
xnor U20196 (N_20196,N_15296,N_15373);
and U20197 (N_20197,N_15893,N_15024);
and U20198 (N_20198,N_17629,N_16581);
nor U20199 (N_20199,N_17933,N_15607);
nand U20200 (N_20200,N_17781,N_17659);
xnor U20201 (N_20201,N_15723,N_15191);
xnor U20202 (N_20202,N_15973,N_16053);
xnor U20203 (N_20203,N_15259,N_15773);
or U20204 (N_20204,N_17782,N_16017);
nor U20205 (N_20205,N_17162,N_17098);
nor U20206 (N_20206,N_15696,N_15701);
and U20207 (N_20207,N_17568,N_17562);
nor U20208 (N_20208,N_16329,N_15317);
or U20209 (N_20209,N_15919,N_16694);
and U20210 (N_20210,N_16679,N_17123);
nand U20211 (N_20211,N_17576,N_16530);
or U20212 (N_20212,N_17180,N_17312);
and U20213 (N_20213,N_17949,N_16183);
and U20214 (N_20214,N_16943,N_16897);
nand U20215 (N_20215,N_17189,N_17182);
nor U20216 (N_20216,N_15290,N_15137);
and U20217 (N_20217,N_17457,N_17731);
xor U20218 (N_20218,N_16424,N_15901);
nand U20219 (N_20219,N_15157,N_16366);
nor U20220 (N_20220,N_17430,N_15314);
nand U20221 (N_20221,N_16052,N_15008);
xor U20222 (N_20222,N_15778,N_15296);
or U20223 (N_20223,N_16284,N_15333);
nor U20224 (N_20224,N_16303,N_17571);
or U20225 (N_20225,N_17430,N_15838);
xnor U20226 (N_20226,N_17195,N_15634);
or U20227 (N_20227,N_17645,N_16411);
nor U20228 (N_20228,N_16913,N_16697);
nor U20229 (N_20229,N_16690,N_17233);
nand U20230 (N_20230,N_17683,N_16313);
or U20231 (N_20231,N_17246,N_17337);
and U20232 (N_20232,N_15288,N_17055);
xnor U20233 (N_20233,N_15176,N_16254);
and U20234 (N_20234,N_15652,N_15591);
or U20235 (N_20235,N_16901,N_15749);
nand U20236 (N_20236,N_17948,N_15663);
xnor U20237 (N_20237,N_17712,N_17416);
or U20238 (N_20238,N_15822,N_15550);
xnor U20239 (N_20239,N_15893,N_17635);
nor U20240 (N_20240,N_15536,N_15278);
nor U20241 (N_20241,N_16595,N_16303);
nand U20242 (N_20242,N_17153,N_15593);
and U20243 (N_20243,N_15356,N_16068);
or U20244 (N_20244,N_15180,N_17223);
nor U20245 (N_20245,N_16486,N_17592);
xor U20246 (N_20246,N_16710,N_17230);
or U20247 (N_20247,N_15989,N_17134);
or U20248 (N_20248,N_15563,N_16730);
and U20249 (N_20249,N_15757,N_15939);
and U20250 (N_20250,N_17657,N_16078);
nor U20251 (N_20251,N_15317,N_15445);
and U20252 (N_20252,N_17921,N_17298);
nor U20253 (N_20253,N_17552,N_16380);
xor U20254 (N_20254,N_17961,N_15404);
and U20255 (N_20255,N_17841,N_16866);
or U20256 (N_20256,N_15902,N_17566);
nor U20257 (N_20257,N_16068,N_16838);
nor U20258 (N_20258,N_16703,N_16187);
xor U20259 (N_20259,N_16273,N_16909);
or U20260 (N_20260,N_15919,N_16397);
and U20261 (N_20261,N_17425,N_17031);
and U20262 (N_20262,N_17551,N_17106);
xnor U20263 (N_20263,N_15830,N_15116);
nand U20264 (N_20264,N_15169,N_17343);
nand U20265 (N_20265,N_16423,N_16744);
nor U20266 (N_20266,N_15841,N_15238);
or U20267 (N_20267,N_16356,N_15869);
nor U20268 (N_20268,N_15017,N_16280);
and U20269 (N_20269,N_15603,N_17508);
or U20270 (N_20270,N_16283,N_16579);
xnor U20271 (N_20271,N_15976,N_17236);
or U20272 (N_20272,N_16098,N_17499);
nand U20273 (N_20273,N_15833,N_16522);
xor U20274 (N_20274,N_17150,N_17461);
nand U20275 (N_20275,N_15952,N_17221);
xnor U20276 (N_20276,N_16833,N_16509);
nor U20277 (N_20277,N_15768,N_15259);
or U20278 (N_20278,N_16692,N_15492);
nor U20279 (N_20279,N_16382,N_15427);
nand U20280 (N_20280,N_15858,N_16900);
xor U20281 (N_20281,N_15966,N_15198);
nand U20282 (N_20282,N_15431,N_17085);
xnor U20283 (N_20283,N_17904,N_15640);
nor U20284 (N_20284,N_17115,N_17119);
and U20285 (N_20285,N_17513,N_15379);
nor U20286 (N_20286,N_17567,N_15423);
xnor U20287 (N_20287,N_15874,N_16220);
and U20288 (N_20288,N_16319,N_17310);
nor U20289 (N_20289,N_15628,N_16798);
xor U20290 (N_20290,N_16521,N_15522);
nand U20291 (N_20291,N_17981,N_16945);
or U20292 (N_20292,N_17014,N_15032);
or U20293 (N_20293,N_17135,N_17124);
or U20294 (N_20294,N_17417,N_17267);
or U20295 (N_20295,N_17354,N_15944);
or U20296 (N_20296,N_16313,N_15840);
nor U20297 (N_20297,N_16601,N_16051);
nor U20298 (N_20298,N_16481,N_17613);
nand U20299 (N_20299,N_16459,N_16930);
nor U20300 (N_20300,N_17315,N_17692);
or U20301 (N_20301,N_15818,N_16725);
or U20302 (N_20302,N_17895,N_16734);
and U20303 (N_20303,N_15481,N_17692);
and U20304 (N_20304,N_16037,N_16791);
nor U20305 (N_20305,N_16892,N_17649);
nor U20306 (N_20306,N_15619,N_15879);
nand U20307 (N_20307,N_17984,N_16802);
nor U20308 (N_20308,N_15141,N_16290);
nor U20309 (N_20309,N_16990,N_17307);
or U20310 (N_20310,N_16570,N_15182);
and U20311 (N_20311,N_17501,N_17390);
nor U20312 (N_20312,N_17875,N_15563);
nand U20313 (N_20313,N_17343,N_16985);
nor U20314 (N_20314,N_15762,N_15372);
or U20315 (N_20315,N_15237,N_17836);
nor U20316 (N_20316,N_16376,N_15062);
xor U20317 (N_20317,N_16914,N_17282);
and U20318 (N_20318,N_16434,N_17254);
or U20319 (N_20319,N_16168,N_16122);
nor U20320 (N_20320,N_16995,N_15487);
nor U20321 (N_20321,N_17010,N_15546);
or U20322 (N_20322,N_15427,N_16447);
and U20323 (N_20323,N_17228,N_17921);
xor U20324 (N_20324,N_15637,N_17550);
or U20325 (N_20325,N_15098,N_15739);
nor U20326 (N_20326,N_17757,N_15363);
nor U20327 (N_20327,N_17883,N_17754);
and U20328 (N_20328,N_16910,N_17581);
nor U20329 (N_20329,N_17305,N_15531);
and U20330 (N_20330,N_17855,N_16920);
and U20331 (N_20331,N_15078,N_17305);
nor U20332 (N_20332,N_16309,N_16377);
nor U20333 (N_20333,N_16256,N_15301);
xor U20334 (N_20334,N_16899,N_17123);
nor U20335 (N_20335,N_15207,N_16326);
nor U20336 (N_20336,N_17817,N_15525);
xor U20337 (N_20337,N_15624,N_15294);
and U20338 (N_20338,N_17784,N_16579);
nor U20339 (N_20339,N_16534,N_15017);
nand U20340 (N_20340,N_15321,N_16199);
or U20341 (N_20341,N_16794,N_15247);
and U20342 (N_20342,N_15126,N_16433);
nor U20343 (N_20343,N_15941,N_16213);
and U20344 (N_20344,N_16397,N_15678);
nor U20345 (N_20345,N_15760,N_15541);
or U20346 (N_20346,N_16716,N_16413);
or U20347 (N_20347,N_17417,N_17643);
or U20348 (N_20348,N_17098,N_16021);
xnor U20349 (N_20349,N_17969,N_16347);
nand U20350 (N_20350,N_16442,N_15907);
nor U20351 (N_20351,N_17697,N_16184);
or U20352 (N_20352,N_16701,N_17658);
nor U20353 (N_20353,N_17389,N_17331);
xor U20354 (N_20354,N_15473,N_16515);
xor U20355 (N_20355,N_15322,N_16489);
and U20356 (N_20356,N_15349,N_15226);
or U20357 (N_20357,N_15807,N_17697);
nand U20358 (N_20358,N_15859,N_17874);
xor U20359 (N_20359,N_17947,N_17539);
nor U20360 (N_20360,N_15938,N_17896);
xor U20361 (N_20361,N_15592,N_16488);
or U20362 (N_20362,N_16425,N_17812);
or U20363 (N_20363,N_16665,N_16843);
or U20364 (N_20364,N_15447,N_16976);
xnor U20365 (N_20365,N_16580,N_17465);
xnor U20366 (N_20366,N_17321,N_15315);
xnor U20367 (N_20367,N_15678,N_17632);
nor U20368 (N_20368,N_17027,N_16846);
and U20369 (N_20369,N_16353,N_16269);
and U20370 (N_20370,N_15166,N_17471);
nand U20371 (N_20371,N_17037,N_15943);
or U20372 (N_20372,N_16833,N_15673);
xor U20373 (N_20373,N_15611,N_15121);
xnor U20374 (N_20374,N_17359,N_16299);
or U20375 (N_20375,N_15121,N_16217);
or U20376 (N_20376,N_17518,N_16696);
nor U20377 (N_20377,N_17378,N_16747);
nand U20378 (N_20378,N_17574,N_16737);
nand U20379 (N_20379,N_15423,N_15674);
or U20380 (N_20380,N_15751,N_17421);
nor U20381 (N_20381,N_15979,N_17387);
nor U20382 (N_20382,N_17083,N_15738);
nor U20383 (N_20383,N_15810,N_15599);
nor U20384 (N_20384,N_15949,N_15743);
nor U20385 (N_20385,N_16983,N_16806);
and U20386 (N_20386,N_15072,N_17363);
or U20387 (N_20387,N_15032,N_17483);
and U20388 (N_20388,N_15984,N_16088);
nand U20389 (N_20389,N_17191,N_17713);
or U20390 (N_20390,N_16100,N_17035);
nand U20391 (N_20391,N_15747,N_16273);
or U20392 (N_20392,N_15577,N_16096);
or U20393 (N_20393,N_15693,N_16197);
or U20394 (N_20394,N_17514,N_16783);
or U20395 (N_20395,N_17176,N_15747);
or U20396 (N_20396,N_15516,N_16661);
or U20397 (N_20397,N_16653,N_16661);
nand U20398 (N_20398,N_15259,N_17707);
nor U20399 (N_20399,N_16432,N_16641);
nor U20400 (N_20400,N_15287,N_17086);
and U20401 (N_20401,N_15383,N_17266);
and U20402 (N_20402,N_16229,N_17618);
or U20403 (N_20403,N_17602,N_16650);
nand U20404 (N_20404,N_17428,N_16616);
nand U20405 (N_20405,N_15406,N_17580);
and U20406 (N_20406,N_15694,N_17740);
xnor U20407 (N_20407,N_15489,N_16210);
or U20408 (N_20408,N_15622,N_15029);
or U20409 (N_20409,N_15252,N_17478);
or U20410 (N_20410,N_17860,N_15330);
or U20411 (N_20411,N_16924,N_16798);
xnor U20412 (N_20412,N_15365,N_17817);
xnor U20413 (N_20413,N_15623,N_17272);
nand U20414 (N_20414,N_17070,N_15867);
nor U20415 (N_20415,N_16192,N_15606);
and U20416 (N_20416,N_17712,N_16961);
nand U20417 (N_20417,N_15878,N_15560);
and U20418 (N_20418,N_15799,N_16600);
and U20419 (N_20419,N_17836,N_15734);
and U20420 (N_20420,N_15245,N_16372);
and U20421 (N_20421,N_17897,N_16393);
nand U20422 (N_20422,N_16715,N_17696);
nor U20423 (N_20423,N_16342,N_16934);
xnor U20424 (N_20424,N_17507,N_16589);
or U20425 (N_20425,N_15753,N_15871);
and U20426 (N_20426,N_15585,N_17574);
xor U20427 (N_20427,N_16201,N_17416);
nor U20428 (N_20428,N_15013,N_15739);
or U20429 (N_20429,N_15287,N_16589);
or U20430 (N_20430,N_15162,N_16889);
and U20431 (N_20431,N_17550,N_15661);
or U20432 (N_20432,N_16102,N_16418);
or U20433 (N_20433,N_15294,N_16784);
xor U20434 (N_20434,N_15781,N_16204);
or U20435 (N_20435,N_15920,N_16214);
nand U20436 (N_20436,N_15625,N_15484);
nor U20437 (N_20437,N_16479,N_17963);
nand U20438 (N_20438,N_15134,N_17857);
and U20439 (N_20439,N_15813,N_16327);
nor U20440 (N_20440,N_16578,N_16533);
or U20441 (N_20441,N_16286,N_15166);
nand U20442 (N_20442,N_17103,N_17665);
nand U20443 (N_20443,N_15257,N_15848);
nor U20444 (N_20444,N_16908,N_15722);
or U20445 (N_20445,N_15544,N_16497);
xnor U20446 (N_20446,N_17231,N_15924);
nand U20447 (N_20447,N_16786,N_15417);
nand U20448 (N_20448,N_16818,N_15849);
and U20449 (N_20449,N_17399,N_16246);
nor U20450 (N_20450,N_16477,N_17457);
nand U20451 (N_20451,N_17025,N_16881);
or U20452 (N_20452,N_17640,N_15778);
or U20453 (N_20453,N_17694,N_17931);
nor U20454 (N_20454,N_17080,N_16263);
and U20455 (N_20455,N_16010,N_15629);
and U20456 (N_20456,N_17171,N_16775);
nor U20457 (N_20457,N_17788,N_16145);
nor U20458 (N_20458,N_15336,N_15803);
nand U20459 (N_20459,N_15561,N_17416);
or U20460 (N_20460,N_15928,N_15194);
and U20461 (N_20461,N_17413,N_15750);
nor U20462 (N_20462,N_17368,N_16625);
and U20463 (N_20463,N_17547,N_17544);
and U20464 (N_20464,N_17248,N_17747);
or U20465 (N_20465,N_16549,N_16130);
and U20466 (N_20466,N_16832,N_16464);
nand U20467 (N_20467,N_17011,N_17000);
and U20468 (N_20468,N_15934,N_16345);
or U20469 (N_20469,N_17040,N_17932);
nor U20470 (N_20470,N_16757,N_17503);
and U20471 (N_20471,N_15970,N_15849);
and U20472 (N_20472,N_17607,N_15665);
nor U20473 (N_20473,N_15289,N_16717);
nor U20474 (N_20474,N_17710,N_15607);
nor U20475 (N_20475,N_15388,N_15335);
and U20476 (N_20476,N_15643,N_15771);
nand U20477 (N_20477,N_15089,N_17752);
nor U20478 (N_20478,N_15570,N_17845);
xor U20479 (N_20479,N_16399,N_15053);
and U20480 (N_20480,N_17562,N_16812);
nor U20481 (N_20481,N_17770,N_16122);
nand U20482 (N_20482,N_17301,N_15703);
and U20483 (N_20483,N_16526,N_15273);
and U20484 (N_20484,N_15839,N_15178);
xnor U20485 (N_20485,N_17784,N_15878);
xnor U20486 (N_20486,N_15138,N_17521);
xor U20487 (N_20487,N_15077,N_15404);
xor U20488 (N_20488,N_17151,N_15838);
xnor U20489 (N_20489,N_16720,N_15339);
nor U20490 (N_20490,N_17808,N_16742);
xnor U20491 (N_20491,N_17416,N_17123);
and U20492 (N_20492,N_16542,N_16868);
or U20493 (N_20493,N_16787,N_16670);
nor U20494 (N_20494,N_16556,N_17075);
nor U20495 (N_20495,N_15911,N_15916);
and U20496 (N_20496,N_15801,N_17647);
and U20497 (N_20497,N_15358,N_16299);
and U20498 (N_20498,N_17563,N_17632);
and U20499 (N_20499,N_16934,N_15334);
or U20500 (N_20500,N_16292,N_16051);
and U20501 (N_20501,N_16534,N_15029);
and U20502 (N_20502,N_16904,N_17181);
nor U20503 (N_20503,N_17720,N_16927);
nor U20504 (N_20504,N_16642,N_16462);
xor U20505 (N_20505,N_17316,N_16577);
and U20506 (N_20506,N_15150,N_16897);
nand U20507 (N_20507,N_15707,N_17306);
and U20508 (N_20508,N_17084,N_16188);
nor U20509 (N_20509,N_15967,N_17802);
nor U20510 (N_20510,N_17761,N_17902);
or U20511 (N_20511,N_15291,N_15509);
xnor U20512 (N_20512,N_16527,N_16158);
xnor U20513 (N_20513,N_15838,N_16746);
nor U20514 (N_20514,N_17986,N_17371);
nor U20515 (N_20515,N_16106,N_15598);
and U20516 (N_20516,N_16987,N_15251);
or U20517 (N_20517,N_15565,N_17332);
xnor U20518 (N_20518,N_17548,N_15636);
and U20519 (N_20519,N_16533,N_15047);
nand U20520 (N_20520,N_17117,N_16695);
nor U20521 (N_20521,N_16545,N_15688);
or U20522 (N_20522,N_17187,N_17435);
and U20523 (N_20523,N_17372,N_15780);
nor U20524 (N_20524,N_17429,N_16268);
and U20525 (N_20525,N_17366,N_17376);
xnor U20526 (N_20526,N_15372,N_15639);
nor U20527 (N_20527,N_15202,N_17645);
nand U20528 (N_20528,N_16162,N_17211);
nand U20529 (N_20529,N_15535,N_15543);
or U20530 (N_20530,N_15251,N_16947);
or U20531 (N_20531,N_16437,N_16335);
nand U20532 (N_20532,N_16611,N_16332);
and U20533 (N_20533,N_16933,N_16509);
or U20534 (N_20534,N_15222,N_15948);
nand U20535 (N_20535,N_17437,N_15107);
or U20536 (N_20536,N_15081,N_15992);
nand U20537 (N_20537,N_16866,N_15024);
xnor U20538 (N_20538,N_17355,N_15021);
nor U20539 (N_20539,N_16377,N_15423);
nor U20540 (N_20540,N_17825,N_17806);
and U20541 (N_20541,N_16989,N_16232);
and U20542 (N_20542,N_17900,N_17117);
and U20543 (N_20543,N_15309,N_17739);
or U20544 (N_20544,N_16687,N_15394);
or U20545 (N_20545,N_15443,N_17817);
nand U20546 (N_20546,N_16422,N_16208);
nand U20547 (N_20547,N_17350,N_16777);
nor U20548 (N_20548,N_16527,N_15295);
nand U20549 (N_20549,N_15937,N_17760);
nor U20550 (N_20550,N_16707,N_15003);
and U20551 (N_20551,N_17550,N_16471);
nand U20552 (N_20552,N_17129,N_17222);
nand U20553 (N_20553,N_17116,N_17777);
or U20554 (N_20554,N_15162,N_17686);
or U20555 (N_20555,N_17556,N_16871);
xnor U20556 (N_20556,N_17771,N_15645);
and U20557 (N_20557,N_17784,N_15208);
nor U20558 (N_20558,N_15121,N_15126);
or U20559 (N_20559,N_16578,N_15962);
and U20560 (N_20560,N_17831,N_16884);
nor U20561 (N_20561,N_17738,N_16866);
nand U20562 (N_20562,N_15748,N_17043);
xnor U20563 (N_20563,N_17621,N_17868);
nand U20564 (N_20564,N_17888,N_17013);
and U20565 (N_20565,N_15731,N_15838);
and U20566 (N_20566,N_15678,N_15400);
xor U20567 (N_20567,N_17523,N_17491);
xor U20568 (N_20568,N_16880,N_17566);
xnor U20569 (N_20569,N_15383,N_17845);
xnor U20570 (N_20570,N_16319,N_15883);
and U20571 (N_20571,N_16906,N_15954);
or U20572 (N_20572,N_16318,N_17429);
nor U20573 (N_20573,N_16005,N_17432);
or U20574 (N_20574,N_16500,N_15076);
xor U20575 (N_20575,N_16162,N_15088);
nand U20576 (N_20576,N_15174,N_17215);
and U20577 (N_20577,N_16014,N_16832);
or U20578 (N_20578,N_16644,N_16843);
xnor U20579 (N_20579,N_16945,N_15627);
and U20580 (N_20580,N_16450,N_16497);
and U20581 (N_20581,N_17688,N_17220);
or U20582 (N_20582,N_15365,N_15718);
nor U20583 (N_20583,N_17389,N_17415);
xor U20584 (N_20584,N_17150,N_16804);
or U20585 (N_20585,N_17090,N_17601);
or U20586 (N_20586,N_16601,N_16664);
nand U20587 (N_20587,N_17032,N_15325);
xor U20588 (N_20588,N_16986,N_16410);
xor U20589 (N_20589,N_15610,N_15345);
or U20590 (N_20590,N_17288,N_16410);
or U20591 (N_20591,N_16008,N_16631);
xor U20592 (N_20592,N_15830,N_16288);
or U20593 (N_20593,N_17414,N_17278);
or U20594 (N_20594,N_16002,N_17227);
and U20595 (N_20595,N_15460,N_16007);
nor U20596 (N_20596,N_16379,N_16193);
nand U20597 (N_20597,N_17918,N_16570);
nand U20598 (N_20598,N_15717,N_16555);
and U20599 (N_20599,N_15760,N_15117);
nor U20600 (N_20600,N_15245,N_16977);
nand U20601 (N_20601,N_16519,N_15842);
xor U20602 (N_20602,N_15875,N_17281);
xnor U20603 (N_20603,N_15498,N_17658);
or U20604 (N_20604,N_16150,N_15567);
xnor U20605 (N_20605,N_15786,N_16918);
xnor U20606 (N_20606,N_16804,N_17152);
nor U20607 (N_20607,N_16899,N_16378);
xor U20608 (N_20608,N_17367,N_16166);
nor U20609 (N_20609,N_15996,N_16860);
nand U20610 (N_20610,N_17400,N_15775);
xor U20611 (N_20611,N_15636,N_16493);
nor U20612 (N_20612,N_15632,N_15305);
nand U20613 (N_20613,N_17954,N_16882);
and U20614 (N_20614,N_15570,N_17651);
and U20615 (N_20615,N_16540,N_15699);
and U20616 (N_20616,N_17902,N_16183);
nand U20617 (N_20617,N_15062,N_17631);
xor U20618 (N_20618,N_15912,N_16888);
xor U20619 (N_20619,N_16077,N_15312);
or U20620 (N_20620,N_16883,N_16004);
nand U20621 (N_20621,N_15101,N_17645);
nand U20622 (N_20622,N_16678,N_15188);
and U20623 (N_20623,N_15398,N_17415);
and U20624 (N_20624,N_15447,N_16510);
nor U20625 (N_20625,N_15504,N_16095);
nand U20626 (N_20626,N_17612,N_17762);
nor U20627 (N_20627,N_16736,N_15098);
or U20628 (N_20628,N_17666,N_17608);
nand U20629 (N_20629,N_15955,N_15441);
xor U20630 (N_20630,N_15543,N_16799);
or U20631 (N_20631,N_16881,N_15796);
and U20632 (N_20632,N_16071,N_16076);
xnor U20633 (N_20633,N_15927,N_15002);
or U20634 (N_20634,N_16368,N_17709);
nand U20635 (N_20635,N_16847,N_17490);
xor U20636 (N_20636,N_17529,N_17922);
or U20637 (N_20637,N_16118,N_16363);
or U20638 (N_20638,N_17314,N_16414);
nand U20639 (N_20639,N_15598,N_17715);
or U20640 (N_20640,N_17810,N_17723);
nor U20641 (N_20641,N_16172,N_16490);
xor U20642 (N_20642,N_17397,N_16744);
nand U20643 (N_20643,N_17491,N_17356);
xnor U20644 (N_20644,N_17326,N_15744);
or U20645 (N_20645,N_17785,N_15406);
nand U20646 (N_20646,N_16579,N_16431);
nor U20647 (N_20647,N_17990,N_16334);
nand U20648 (N_20648,N_16700,N_15323);
nand U20649 (N_20649,N_16084,N_16021);
nor U20650 (N_20650,N_16992,N_16137);
nand U20651 (N_20651,N_16481,N_16722);
nor U20652 (N_20652,N_16331,N_15953);
or U20653 (N_20653,N_16753,N_17753);
nor U20654 (N_20654,N_15175,N_17360);
nand U20655 (N_20655,N_15824,N_16013);
or U20656 (N_20656,N_15051,N_16718);
nand U20657 (N_20657,N_16419,N_15674);
nor U20658 (N_20658,N_17004,N_15858);
nand U20659 (N_20659,N_15673,N_16658);
nor U20660 (N_20660,N_15231,N_17931);
or U20661 (N_20661,N_17857,N_17813);
or U20662 (N_20662,N_17234,N_16091);
nor U20663 (N_20663,N_15218,N_16047);
nand U20664 (N_20664,N_17639,N_16690);
xor U20665 (N_20665,N_15070,N_16886);
xor U20666 (N_20666,N_15541,N_15107);
or U20667 (N_20667,N_17833,N_17447);
or U20668 (N_20668,N_16896,N_17973);
and U20669 (N_20669,N_17534,N_16092);
nand U20670 (N_20670,N_16139,N_16075);
nand U20671 (N_20671,N_16409,N_15063);
nor U20672 (N_20672,N_17032,N_16449);
and U20673 (N_20673,N_16407,N_15000);
or U20674 (N_20674,N_17195,N_16971);
and U20675 (N_20675,N_16940,N_17849);
and U20676 (N_20676,N_16228,N_17200);
or U20677 (N_20677,N_15425,N_15370);
and U20678 (N_20678,N_17583,N_15258);
or U20679 (N_20679,N_15356,N_16403);
or U20680 (N_20680,N_15081,N_16951);
and U20681 (N_20681,N_15118,N_15842);
xor U20682 (N_20682,N_15225,N_17108);
xor U20683 (N_20683,N_15233,N_17615);
nand U20684 (N_20684,N_17167,N_15816);
nor U20685 (N_20685,N_15267,N_16960);
xor U20686 (N_20686,N_15098,N_15858);
nor U20687 (N_20687,N_17588,N_16801);
xor U20688 (N_20688,N_15946,N_16782);
xor U20689 (N_20689,N_17734,N_16779);
nor U20690 (N_20690,N_15982,N_16051);
and U20691 (N_20691,N_15814,N_15084);
nor U20692 (N_20692,N_16779,N_16479);
nor U20693 (N_20693,N_16624,N_17391);
xnor U20694 (N_20694,N_16394,N_16609);
or U20695 (N_20695,N_15233,N_16676);
xnor U20696 (N_20696,N_15722,N_15689);
xnor U20697 (N_20697,N_16421,N_16031);
nand U20698 (N_20698,N_15154,N_17941);
nand U20699 (N_20699,N_16237,N_16757);
and U20700 (N_20700,N_15878,N_17309);
xor U20701 (N_20701,N_17483,N_17232);
nor U20702 (N_20702,N_15352,N_15798);
or U20703 (N_20703,N_17335,N_15786);
nor U20704 (N_20704,N_17475,N_17772);
nand U20705 (N_20705,N_17708,N_16356);
xnor U20706 (N_20706,N_17118,N_17684);
nand U20707 (N_20707,N_15731,N_16459);
or U20708 (N_20708,N_16803,N_16826);
nand U20709 (N_20709,N_17400,N_17465);
and U20710 (N_20710,N_16375,N_17833);
or U20711 (N_20711,N_17784,N_16486);
xor U20712 (N_20712,N_16909,N_17013);
and U20713 (N_20713,N_16562,N_16155);
nand U20714 (N_20714,N_16876,N_16474);
nand U20715 (N_20715,N_15918,N_16333);
or U20716 (N_20716,N_17391,N_15242);
nand U20717 (N_20717,N_17743,N_16019);
nor U20718 (N_20718,N_15988,N_16978);
and U20719 (N_20719,N_17954,N_16260);
nor U20720 (N_20720,N_17265,N_17624);
nor U20721 (N_20721,N_15602,N_17099);
nor U20722 (N_20722,N_16627,N_15607);
and U20723 (N_20723,N_16025,N_15939);
nor U20724 (N_20724,N_15952,N_16892);
xor U20725 (N_20725,N_15977,N_15916);
xnor U20726 (N_20726,N_15216,N_15125);
or U20727 (N_20727,N_15718,N_15328);
xnor U20728 (N_20728,N_15421,N_16491);
nor U20729 (N_20729,N_17673,N_17275);
nor U20730 (N_20730,N_16547,N_15506);
and U20731 (N_20731,N_16154,N_16502);
and U20732 (N_20732,N_15862,N_17076);
xnor U20733 (N_20733,N_16124,N_16980);
and U20734 (N_20734,N_15573,N_15025);
or U20735 (N_20735,N_15660,N_17347);
nor U20736 (N_20736,N_17805,N_17265);
or U20737 (N_20737,N_15532,N_16192);
and U20738 (N_20738,N_17592,N_17698);
or U20739 (N_20739,N_17833,N_16731);
nand U20740 (N_20740,N_15252,N_16472);
nor U20741 (N_20741,N_17046,N_17176);
and U20742 (N_20742,N_17522,N_16489);
nand U20743 (N_20743,N_17422,N_17108);
nor U20744 (N_20744,N_15792,N_17776);
nor U20745 (N_20745,N_15721,N_17306);
nand U20746 (N_20746,N_16255,N_15466);
and U20747 (N_20747,N_17127,N_17642);
nor U20748 (N_20748,N_17239,N_16378);
and U20749 (N_20749,N_16392,N_15429);
xor U20750 (N_20750,N_17216,N_16320);
nor U20751 (N_20751,N_15512,N_15541);
xor U20752 (N_20752,N_16637,N_15564);
and U20753 (N_20753,N_17542,N_16283);
nand U20754 (N_20754,N_15038,N_16559);
nand U20755 (N_20755,N_17749,N_15194);
xnor U20756 (N_20756,N_15930,N_17604);
and U20757 (N_20757,N_17079,N_17736);
nor U20758 (N_20758,N_17577,N_16488);
and U20759 (N_20759,N_17853,N_17938);
nor U20760 (N_20760,N_15362,N_17406);
nand U20761 (N_20761,N_16886,N_17352);
or U20762 (N_20762,N_16054,N_17037);
and U20763 (N_20763,N_17844,N_16627);
nand U20764 (N_20764,N_16416,N_16234);
nand U20765 (N_20765,N_16162,N_16705);
nand U20766 (N_20766,N_15376,N_16188);
xnor U20767 (N_20767,N_17497,N_17388);
nand U20768 (N_20768,N_15684,N_15450);
nor U20769 (N_20769,N_16141,N_17222);
or U20770 (N_20770,N_16218,N_15422);
or U20771 (N_20771,N_15215,N_17391);
nand U20772 (N_20772,N_16189,N_17236);
xor U20773 (N_20773,N_15728,N_17077);
nor U20774 (N_20774,N_15354,N_15613);
or U20775 (N_20775,N_17615,N_17768);
nand U20776 (N_20776,N_15277,N_16257);
or U20777 (N_20777,N_15172,N_17482);
nor U20778 (N_20778,N_17372,N_16163);
or U20779 (N_20779,N_15801,N_17473);
or U20780 (N_20780,N_15919,N_16725);
xnor U20781 (N_20781,N_16643,N_17811);
and U20782 (N_20782,N_15921,N_17974);
nand U20783 (N_20783,N_16926,N_17258);
nor U20784 (N_20784,N_17051,N_17993);
nand U20785 (N_20785,N_17239,N_16987);
nor U20786 (N_20786,N_15719,N_16434);
nor U20787 (N_20787,N_17877,N_17383);
nand U20788 (N_20788,N_16724,N_16001);
xor U20789 (N_20789,N_17774,N_17754);
xnor U20790 (N_20790,N_16858,N_16909);
xor U20791 (N_20791,N_17703,N_17632);
nor U20792 (N_20792,N_16588,N_17172);
xor U20793 (N_20793,N_16038,N_17776);
nand U20794 (N_20794,N_15240,N_17238);
xnor U20795 (N_20795,N_17917,N_15322);
nor U20796 (N_20796,N_17704,N_16961);
or U20797 (N_20797,N_17682,N_15660);
and U20798 (N_20798,N_17317,N_17971);
nand U20799 (N_20799,N_15058,N_16585);
or U20800 (N_20800,N_17853,N_17016);
nand U20801 (N_20801,N_15875,N_16955);
nand U20802 (N_20802,N_15621,N_16109);
xor U20803 (N_20803,N_16685,N_16951);
nand U20804 (N_20804,N_15265,N_17612);
and U20805 (N_20805,N_16350,N_17788);
or U20806 (N_20806,N_16286,N_15700);
and U20807 (N_20807,N_17473,N_15226);
xnor U20808 (N_20808,N_15758,N_16368);
and U20809 (N_20809,N_17315,N_15448);
or U20810 (N_20810,N_16409,N_17978);
and U20811 (N_20811,N_16369,N_15048);
nor U20812 (N_20812,N_15801,N_16874);
and U20813 (N_20813,N_17949,N_16624);
and U20814 (N_20814,N_17862,N_17994);
or U20815 (N_20815,N_15922,N_17610);
and U20816 (N_20816,N_15229,N_17922);
nor U20817 (N_20817,N_17409,N_17232);
and U20818 (N_20818,N_15017,N_17124);
and U20819 (N_20819,N_17974,N_17615);
nand U20820 (N_20820,N_16632,N_16300);
and U20821 (N_20821,N_16839,N_16229);
nand U20822 (N_20822,N_15751,N_17376);
and U20823 (N_20823,N_15532,N_15349);
nand U20824 (N_20824,N_16982,N_17462);
or U20825 (N_20825,N_16230,N_15096);
or U20826 (N_20826,N_16761,N_15204);
or U20827 (N_20827,N_15896,N_17691);
xnor U20828 (N_20828,N_17051,N_16082);
nand U20829 (N_20829,N_16451,N_15875);
nand U20830 (N_20830,N_15017,N_17269);
xor U20831 (N_20831,N_17639,N_17128);
and U20832 (N_20832,N_17028,N_17824);
nor U20833 (N_20833,N_17887,N_15534);
nor U20834 (N_20834,N_17872,N_15837);
or U20835 (N_20835,N_16442,N_15287);
xor U20836 (N_20836,N_16642,N_16833);
nor U20837 (N_20837,N_16282,N_16726);
xnor U20838 (N_20838,N_15943,N_16991);
and U20839 (N_20839,N_16506,N_15527);
nand U20840 (N_20840,N_16620,N_16328);
and U20841 (N_20841,N_17782,N_15333);
nand U20842 (N_20842,N_16807,N_16607);
nand U20843 (N_20843,N_16064,N_15132);
and U20844 (N_20844,N_15480,N_15939);
or U20845 (N_20845,N_17585,N_17130);
and U20846 (N_20846,N_15588,N_15662);
xnor U20847 (N_20847,N_17753,N_15292);
nand U20848 (N_20848,N_16600,N_15592);
and U20849 (N_20849,N_16061,N_15914);
nand U20850 (N_20850,N_16342,N_16360);
and U20851 (N_20851,N_16040,N_17275);
and U20852 (N_20852,N_17070,N_17101);
nor U20853 (N_20853,N_15187,N_17850);
xnor U20854 (N_20854,N_17003,N_15848);
or U20855 (N_20855,N_17531,N_17159);
xor U20856 (N_20856,N_16200,N_17904);
nand U20857 (N_20857,N_16467,N_16295);
nor U20858 (N_20858,N_15746,N_15820);
and U20859 (N_20859,N_16203,N_17900);
or U20860 (N_20860,N_15408,N_16503);
nand U20861 (N_20861,N_17031,N_16144);
nand U20862 (N_20862,N_16783,N_16915);
nor U20863 (N_20863,N_15040,N_15390);
or U20864 (N_20864,N_15926,N_17199);
and U20865 (N_20865,N_15136,N_16827);
nand U20866 (N_20866,N_17223,N_17678);
nand U20867 (N_20867,N_15426,N_15286);
and U20868 (N_20868,N_16151,N_16261);
nand U20869 (N_20869,N_15789,N_17166);
nor U20870 (N_20870,N_15501,N_15880);
and U20871 (N_20871,N_16800,N_17067);
and U20872 (N_20872,N_17783,N_15652);
or U20873 (N_20873,N_15096,N_15067);
and U20874 (N_20874,N_15579,N_15021);
and U20875 (N_20875,N_16586,N_17832);
nand U20876 (N_20876,N_16838,N_15624);
nand U20877 (N_20877,N_16024,N_16409);
xor U20878 (N_20878,N_17232,N_17894);
and U20879 (N_20879,N_15220,N_15430);
and U20880 (N_20880,N_16764,N_16399);
nor U20881 (N_20881,N_15605,N_17304);
nor U20882 (N_20882,N_17190,N_15254);
nand U20883 (N_20883,N_17154,N_16989);
or U20884 (N_20884,N_17941,N_17416);
nor U20885 (N_20885,N_16058,N_15314);
nand U20886 (N_20886,N_16449,N_15177);
and U20887 (N_20887,N_16113,N_15648);
xor U20888 (N_20888,N_16788,N_17941);
xnor U20889 (N_20889,N_17702,N_17760);
xnor U20890 (N_20890,N_17529,N_17953);
nor U20891 (N_20891,N_17461,N_17010);
nor U20892 (N_20892,N_16539,N_17790);
xnor U20893 (N_20893,N_16216,N_15662);
or U20894 (N_20894,N_16765,N_15193);
or U20895 (N_20895,N_17970,N_15562);
or U20896 (N_20896,N_15445,N_17069);
nor U20897 (N_20897,N_15393,N_15359);
and U20898 (N_20898,N_16931,N_15161);
or U20899 (N_20899,N_15753,N_15603);
nand U20900 (N_20900,N_17545,N_16877);
and U20901 (N_20901,N_17902,N_16625);
and U20902 (N_20902,N_16590,N_17634);
xor U20903 (N_20903,N_15338,N_17080);
nor U20904 (N_20904,N_17428,N_16883);
nor U20905 (N_20905,N_16757,N_15594);
or U20906 (N_20906,N_15116,N_17825);
or U20907 (N_20907,N_17337,N_17137);
nor U20908 (N_20908,N_15736,N_17903);
nand U20909 (N_20909,N_16143,N_15948);
nor U20910 (N_20910,N_15814,N_17825);
nand U20911 (N_20911,N_15552,N_17056);
nor U20912 (N_20912,N_17578,N_17667);
nor U20913 (N_20913,N_17859,N_17569);
or U20914 (N_20914,N_16243,N_16376);
nand U20915 (N_20915,N_17460,N_15799);
or U20916 (N_20916,N_15250,N_15307);
xor U20917 (N_20917,N_15419,N_16624);
xor U20918 (N_20918,N_17402,N_16364);
or U20919 (N_20919,N_17719,N_16084);
nand U20920 (N_20920,N_15645,N_16750);
xor U20921 (N_20921,N_16466,N_17729);
nor U20922 (N_20922,N_16572,N_16786);
nor U20923 (N_20923,N_15644,N_15027);
xor U20924 (N_20924,N_17395,N_16849);
xor U20925 (N_20925,N_15738,N_15383);
or U20926 (N_20926,N_17835,N_15231);
and U20927 (N_20927,N_16508,N_17989);
nand U20928 (N_20928,N_15068,N_17105);
xor U20929 (N_20929,N_16363,N_16956);
and U20930 (N_20930,N_16445,N_16152);
nor U20931 (N_20931,N_16048,N_17590);
nor U20932 (N_20932,N_17617,N_17235);
or U20933 (N_20933,N_16311,N_16959);
or U20934 (N_20934,N_15482,N_15841);
and U20935 (N_20935,N_16860,N_15282);
nand U20936 (N_20936,N_15499,N_16129);
nor U20937 (N_20937,N_15841,N_17387);
or U20938 (N_20938,N_16204,N_16119);
xor U20939 (N_20939,N_16061,N_15501);
xor U20940 (N_20940,N_16054,N_17907);
and U20941 (N_20941,N_17578,N_15113);
xnor U20942 (N_20942,N_16175,N_15029);
and U20943 (N_20943,N_17866,N_17240);
xor U20944 (N_20944,N_17372,N_15183);
nor U20945 (N_20945,N_15376,N_15575);
nor U20946 (N_20946,N_17503,N_16318);
and U20947 (N_20947,N_16778,N_16781);
nand U20948 (N_20948,N_15505,N_16595);
or U20949 (N_20949,N_15849,N_16732);
nand U20950 (N_20950,N_16136,N_16361);
and U20951 (N_20951,N_17007,N_17704);
nor U20952 (N_20952,N_17996,N_17983);
or U20953 (N_20953,N_17225,N_16183);
nor U20954 (N_20954,N_15886,N_17442);
nand U20955 (N_20955,N_17994,N_17243);
and U20956 (N_20956,N_16591,N_16948);
nor U20957 (N_20957,N_16482,N_15951);
xor U20958 (N_20958,N_15653,N_15108);
and U20959 (N_20959,N_17268,N_17341);
and U20960 (N_20960,N_17718,N_15191);
or U20961 (N_20961,N_16101,N_16500);
or U20962 (N_20962,N_17359,N_16276);
nand U20963 (N_20963,N_16682,N_16175);
nand U20964 (N_20964,N_17073,N_17259);
nand U20965 (N_20965,N_17917,N_17617);
and U20966 (N_20966,N_17853,N_15958);
and U20967 (N_20967,N_16788,N_16695);
nor U20968 (N_20968,N_15855,N_16296);
xor U20969 (N_20969,N_16923,N_17951);
and U20970 (N_20970,N_17742,N_16335);
nor U20971 (N_20971,N_16168,N_17126);
nand U20972 (N_20972,N_15263,N_16704);
and U20973 (N_20973,N_15884,N_16754);
and U20974 (N_20974,N_16165,N_17115);
and U20975 (N_20975,N_15987,N_15242);
or U20976 (N_20976,N_17029,N_15377);
xnor U20977 (N_20977,N_16203,N_17353);
nor U20978 (N_20978,N_17876,N_17029);
nor U20979 (N_20979,N_16585,N_16662);
nand U20980 (N_20980,N_15255,N_16931);
nand U20981 (N_20981,N_16776,N_17123);
nor U20982 (N_20982,N_16191,N_16608);
or U20983 (N_20983,N_17833,N_15900);
or U20984 (N_20984,N_17867,N_17470);
nand U20985 (N_20985,N_17731,N_16695);
or U20986 (N_20986,N_17343,N_16178);
nor U20987 (N_20987,N_17241,N_15268);
and U20988 (N_20988,N_15753,N_17321);
and U20989 (N_20989,N_16941,N_17374);
nand U20990 (N_20990,N_15196,N_16252);
nor U20991 (N_20991,N_15549,N_17547);
and U20992 (N_20992,N_16847,N_17244);
and U20993 (N_20993,N_15055,N_16158);
nor U20994 (N_20994,N_16082,N_17490);
nand U20995 (N_20995,N_17189,N_15679);
xor U20996 (N_20996,N_16891,N_17007);
nor U20997 (N_20997,N_17999,N_15916);
or U20998 (N_20998,N_16033,N_16212);
xor U20999 (N_20999,N_16565,N_15310);
nor U21000 (N_21000,N_18987,N_19105);
xnor U21001 (N_21001,N_19329,N_19233);
nor U21002 (N_21002,N_19932,N_20149);
xnor U21003 (N_21003,N_18006,N_20771);
xor U21004 (N_21004,N_18822,N_19960);
and U21005 (N_21005,N_18063,N_18767);
or U21006 (N_21006,N_20978,N_18727);
and U21007 (N_21007,N_19617,N_20344);
nor U21008 (N_21008,N_18089,N_20377);
nand U21009 (N_21009,N_19686,N_19458);
xnor U21010 (N_21010,N_20274,N_20169);
nor U21011 (N_21011,N_20924,N_18653);
or U21012 (N_21012,N_20867,N_18944);
or U21013 (N_21013,N_19814,N_19575);
and U21014 (N_21014,N_18134,N_19839);
nor U21015 (N_21015,N_19530,N_19622);
xor U21016 (N_21016,N_20257,N_18425);
or U21017 (N_21017,N_18000,N_20234);
nand U21018 (N_21018,N_18235,N_19818);
nand U21019 (N_21019,N_20438,N_19920);
and U21020 (N_21020,N_20099,N_19115);
nor U21021 (N_21021,N_18773,N_18298);
nand U21022 (N_21022,N_18098,N_20028);
nand U21023 (N_21023,N_19768,N_20926);
and U21024 (N_21024,N_19051,N_18601);
and U21025 (N_21025,N_19971,N_19654);
nand U21026 (N_21026,N_20063,N_20853);
or U21027 (N_21027,N_18403,N_20158);
nand U21028 (N_21028,N_18287,N_20308);
and U21029 (N_21029,N_19807,N_20248);
nand U21030 (N_21030,N_18898,N_20921);
xnor U21031 (N_21031,N_20850,N_19714);
or U21032 (N_21032,N_19545,N_19604);
nor U21033 (N_21033,N_18528,N_20785);
nor U21034 (N_21034,N_18820,N_20493);
and U21035 (N_21035,N_18448,N_20076);
nand U21036 (N_21036,N_18470,N_18821);
xnor U21037 (N_21037,N_19940,N_18125);
nor U21038 (N_21038,N_19342,N_18884);
xnor U21039 (N_21039,N_20442,N_20016);
nand U21040 (N_21040,N_19741,N_20696);
nand U21041 (N_21041,N_19189,N_18569);
and U21042 (N_21042,N_20560,N_20622);
or U21043 (N_21043,N_19515,N_19528);
and U21044 (N_21044,N_20374,N_19255);
nand U21045 (N_21045,N_18738,N_19273);
and U21046 (N_21046,N_18906,N_20220);
nand U21047 (N_21047,N_18791,N_20406);
nor U21048 (N_21048,N_18223,N_20113);
xor U21049 (N_21049,N_20108,N_18829);
nor U21050 (N_21050,N_18921,N_20885);
nand U21051 (N_21051,N_18310,N_19759);
nor U21052 (N_21052,N_19757,N_20648);
nand U21053 (N_21053,N_19200,N_19346);
or U21054 (N_21054,N_19265,N_19711);
xor U21055 (N_21055,N_20386,N_18943);
xor U21056 (N_21056,N_19028,N_20711);
xor U21057 (N_21057,N_20665,N_19256);
nand U21058 (N_21058,N_20369,N_20598);
xor U21059 (N_21059,N_18260,N_18916);
xnor U21060 (N_21060,N_18766,N_19543);
xor U21061 (N_21061,N_18809,N_20186);
nand U21062 (N_21062,N_19375,N_20241);
nor U21063 (N_21063,N_20167,N_19999);
and U21064 (N_21064,N_19036,N_20574);
or U21065 (N_21065,N_20272,N_20769);
xor U21066 (N_21066,N_18564,N_20893);
xnor U21067 (N_21067,N_18212,N_18572);
and U21068 (N_21068,N_19328,N_19081);
and U21069 (N_21069,N_20196,N_18931);
nor U21070 (N_21070,N_19774,N_20048);
and U21071 (N_21071,N_20425,N_19896);
nand U21072 (N_21072,N_19534,N_20098);
nor U21073 (N_21073,N_19762,N_19518);
or U21074 (N_21074,N_20070,N_19562);
or U21075 (N_21075,N_20929,N_19516);
nor U21076 (N_21076,N_18256,N_20738);
or U21077 (N_21077,N_19345,N_20255);
nor U21078 (N_21078,N_19251,N_19602);
xor U21079 (N_21079,N_19882,N_20767);
and U21080 (N_21080,N_19208,N_19546);
nor U21081 (N_21081,N_18679,N_20403);
nor U21082 (N_21082,N_20841,N_20319);
nand U21083 (N_21083,N_18743,N_20716);
nand U21084 (N_21084,N_19552,N_18157);
nand U21085 (N_21085,N_18302,N_18228);
xnor U21086 (N_21086,N_20343,N_18656);
xor U21087 (N_21087,N_19531,N_18771);
or U21088 (N_21088,N_19243,N_19790);
or U21089 (N_21089,N_20195,N_18913);
nand U21090 (N_21090,N_20539,N_18507);
and U21091 (N_21091,N_18406,N_20170);
nor U21092 (N_21092,N_18051,N_20531);
nor U21093 (N_21093,N_18164,N_20602);
and U21094 (N_21094,N_20400,N_20592);
nand U21095 (N_21095,N_19108,N_19461);
and U21096 (N_21096,N_20429,N_19170);
xor U21097 (N_21097,N_20993,N_19568);
nor U21098 (N_21098,N_18495,N_19409);
nor U21099 (N_21099,N_19628,N_18345);
nand U21100 (N_21100,N_18057,N_18525);
or U21101 (N_21101,N_19596,N_19828);
xnor U21102 (N_21102,N_20032,N_19911);
nand U21103 (N_21103,N_19252,N_18816);
xnor U21104 (N_21104,N_20483,N_20965);
or U21105 (N_21105,N_20887,N_18012);
or U21106 (N_21106,N_18703,N_19067);
nor U21107 (N_21107,N_20776,N_20526);
nand U21108 (N_21108,N_18900,N_18749);
nand U21109 (N_21109,N_18591,N_20194);
nor U21110 (N_21110,N_18460,N_19389);
xnor U21111 (N_21111,N_19196,N_18934);
and U21112 (N_21112,N_18202,N_20511);
or U21113 (N_21113,N_20136,N_20258);
nand U21114 (N_21114,N_20768,N_18759);
xnor U21115 (N_21115,N_19647,N_19572);
and U21116 (N_21116,N_19061,N_19114);
nor U21117 (N_21117,N_20083,N_20759);
xor U21118 (N_21118,N_20705,N_20238);
nand U21119 (N_21119,N_20813,N_18067);
xor U21120 (N_21120,N_18390,N_19808);
xnor U21121 (N_21121,N_20570,N_20732);
and U21122 (N_21122,N_19749,N_19145);
nor U21123 (N_21123,N_20655,N_19627);
xor U21124 (N_21124,N_19047,N_18657);
and U21125 (N_21125,N_19742,N_19120);
or U21126 (N_21126,N_18387,N_20943);
or U21127 (N_21127,N_20524,N_18787);
xor U21128 (N_21128,N_18610,N_20634);
xnor U21129 (N_21129,N_20278,N_19897);
xor U21130 (N_21130,N_19154,N_18644);
nand U21131 (N_21131,N_20860,N_19140);
nand U21132 (N_21132,N_19169,N_18954);
and U21133 (N_21133,N_19282,N_20215);
xor U21134 (N_21134,N_19294,N_19886);
nor U21135 (N_21135,N_18339,N_20565);
nand U21136 (N_21136,N_19783,N_20073);
and U21137 (N_21137,N_19854,N_19758);
or U21138 (N_21138,N_20004,N_20187);
nor U21139 (N_21139,N_20722,N_18937);
or U21140 (N_21140,N_18247,N_18139);
nor U21141 (N_21141,N_18871,N_19365);
or U21142 (N_21142,N_20295,N_18094);
or U21143 (N_21143,N_20119,N_20142);
and U21144 (N_21144,N_19027,N_19476);
nand U21145 (N_21145,N_20065,N_19046);
nor U21146 (N_21146,N_19648,N_18293);
and U21147 (N_21147,N_18112,N_20132);
and U21148 (N_21148,N_19836,N_20733);
or U21149 (N_21149,N_19501,N_20348);
and U21150 (N_21150,N_18492,N_18505);
nand U21151 (N_21151,N_20820,N_19119);
xnor U21152 (N_21152,N_20695,N_19621);
or U21153 (N_21153,N_18803,N_19486);
xor U21154 (N_21154,N_20632,N_18581);
nor U21155 (N_21155,N_18690,N_18537);
and U21156 (N_21156,N_18253,N_19244);
nor U21157 (N_21157,N_18543,N_20506);
xor U21158 (N_21158,N_18945,N_18847);
nor U21159 (N_21159,N_19224,N_18153);
xor U21160 (N_21160,N_19474,N_20986);
and U21161 (N_21161,N_20322,N_19011);
or U21162 (N_21162,N_18694,N_18923);
and U21163 (N_21163,N_20401,N_20433);
nand U21164 (N_21164,N_18190,N_18558);
and U21165 (N_21165,N_19188,N_18734);
and U21166 (N_21166,N_20623,N_19964);
and U21167 (N_21167,N_18263,N_20989);
xnor U21168 (N_21168,N_18192,N_20082);
and U21169 (N_21169,N_18596,N_18480);
and U21170 (N_21170,N_19756,N_19743);
nor U21171 (N_21171,N_20456,N_20720);
nor U21172 (N_21172,N_19193,N_20479);
or U21173 (N_21173,N_19522,N_19553);
and U21174 (N_21174,N_19898,N_20210);
and U21175 (N_21175,N_18915,N_18503);
xnor U21176 (N_21176,N_20330,N_19107);
nor U21177 (N_21177,N_20678,N_20203);
nor U21178 (N_21178,N_18695,N_18385);
xnor U21179 (N_21179,N_19147,N_20532);
and U21180 (N_21180,N_20416,N_18476);
xnor U21181 (N_21181,N_18065,N_19348);
and U21182 (N_21182,N_20101,N_19595);
or U21183 (N_21183,N_18831,N_19677);
and U21184 (N_21184,N_20461,N_18963);
xnor U21185 (N_21185,N_18437,N_18785);
and U21186 (N_21186,N_18969,N_18418);
nand U21187 (N_21187,N_20277,N_19121);
nor U21188 (N_21188,N_20437,N_19434);
nand U21189 (N_21189,N_18401,N_18354);
or U21190 (N_21190,N_20999,N_20380);
or U21191 (N_21191,N_19205,N_20878);
and U21192 (N_21192,N_20795,N_19321);
and U21193 (N_21193,N_19704,N_18184);
nor U21194 (N_21194,N_18179,N_20638);
nor U21195 (N_21195,N_20939,N_20879);
xor U21196 (N_21196,N_19927,N_18824);
nor U21197 (N_21197,N_18928,N_20545);
and U21198 (N_21198,N_19934,N_19423);
nand U21199 (N_21199,N_18687,N_19701);
nor U21200 (N_21200,N_18022,N_18909);
or U21201 (N_21201,N_19418,N_18393);
nor U21202 (N_21202,N_19829,N_19526);
nor U21203 (N_21203,N_19088,N_19429);
xor U21204 (N_21204,N_19791,N_20579);
and U21205 (N_21205,N_20030,N_20452);
xor U21206 (N_21206,N_20951,N_18244);
nand U21207 (N_21207,N_18106,N_18623);
or U21208 (N_21208,N_18198,N_19833);
nor U21209 (N_21209,N_19978,N_20282);
xnor U21210 (N_21210,N_20928,N_20958);
nor U21211 (N_21211,N_19844,N_20530);
or U21212 (N_21212,N_19001,N_18286);
nor U21213 (N_21213,N_18185,N_20730);
nor U21214 (N_21214,N_19106,N_20973);
or U21215 (N_21215,N_20976,N_18872);
xnor U21216 (N_21216,N_18781,N_19715);
nand U21217 (N_21217,N_18011,N_18206);
and U21218 (N_21218,N_20141,N_19507);
and U21219 (N_21219,N_18194,N_18083);
nor U21220 (N_21220,N_18414,N_20882);
nor U21221 (N_21221,N_20902,N_20045);
and U21222 (N_21222,N_20575,N_20576);
nor U21223 (N_21223,N_19057,N_18031);
xnor U21224 (N_21224,N_20525,N_19894);
nand U21225 (N_21225,N_18541,N_18138);
nand U21226 (N_21226,N_20811,N_20129);
nand U21227 (N_21227,N_19161,N_18501);
or U21228 (N_21228,N_18918,N_19888);
xnor U21229 (N_21229,N_18283,N_20778);
or U21230 (N_21230,N_18967,N_18527);
or U21231 (N_21231,N_18182,N_19988);
nor U21232 (N_21232,N_19137,N_19491);
nand U21233 (N_21233,N_18469,N_18045);
or U21234 (N_21234,N_19951,N_18879);
or U21235 (N_21235,N_18713,N_20329);
or U21236 (N_21236,N_20494,N_18003);
and U21237 (N_21237,N_20895,N_20842);
xnor U21238 (N_21238,N_20823,N_19867);
or U21239 (N_21239,N_20341,N_19708);
xnor U21240 (N_21240,N_20447,N_18554);
xnor U21241 (N_21241,N_20420,N_18650);
and U21242 (N_21242,N_19010,N_19962);
xor U21243 (N_21243,N_18150,N_19449);
xor U21244 (N_21244,N_18688,N_20922);
nand U21245 (N_21245,N_18341,N_19338);
and U21246 (N_21246,N_20276,N_19662);
nand U21247 (N_21247,N_18578,N_20726);
nor U21248 (N_21248,N_19379,N_19102);
nor U21249 (N_21249,N_20517,N_18032);
xnor U21250 (N_21250,N_19696,N_20232);
and U21251 (N_21251,N_18976,N_18237);
nor U21252 (N_21252,N_18072,N_20012);
xnor U21253 (N_21253,N_18444,N_19240);
xor U21254 (N_21254,N_18236,N_19767);
or U21255 (N_21255,N_20488,N_20056);
and U21256 (N_21256,N_20037,N_19660);
nor U21257 (N_21257,N_18304,N_19250);
nor U21258 (N_21258,N_19019,N_18248);
nor U21259 (N_21259,N_19798,N_20743);
nor U21260 (N_21260,N_19915,N_20614);
xor U21261 (N_21261,N_18242,N_20050);
or U21262 (N_21262,N_18220,N_20868);
or U21263 (N_21263,N_20947,N_20968);
and U21264 (N_21264,N_20117,N_20584);
nor U21265 (N_21265,N_19733,N_18897);
nor U21266 (N_21266,N_19479,N_18196);
nand U21267 (N_21267,N_18948,N_19272);
nor U21268 (N_21268,N_20619,N_18901);
and U21269 (N_21269,N_19953,N_18896);
or U21270 (N_21270,N_19143,N_18782);
and U21271 (N_21271,N_20994,N_18582);
nand U21272 (N_21272,N_19664,N_20482);
xnor U21273 (N_21273,N_20651,N_19729);
nand U21274 (N_21274,N_18232,N_19269);
nor U21275 (N_21275,N_19573,N_20318);
nor U21276 (N_21276,N_19594,N_19500);
nand U21277 (N_21277,N_19679,N_18097);
and U21278 (N_21278,N_19916,N_18479);
nand U21279 (N_21279,N_19574,N_19626);
and U21280 (N_21280,N_19710,N_20446);
nand U21281 (N_21281,N_20847,N_20478);
nand U21282 (N_21282,N_19049,N_20959);
and U21283 (N_21283,N_19909,N_20345);
xnor U21284 (N_21284,N_20935,N_19416);
or U21285 (N_21285,N_18892,N_20225);
or U21286 (N_21286,N_18812,N_20706);
or U21287 (N_21287,N_19977,N_18477);
nor U21288 (N_21288,N_20957,N_18922);
xor U21289 (N_21289,N_20134,N_20802);
xnor U21290 (N_21290,N_20352,N_18524);
and U21291 (N_21291,N_18508,N_20873);
nand U21292 (N_21292,N_19678,N_19123);
and U21293 (N_21293,N_18736,N_19754);
or U21294 (N_21294,N_20918,N_18868);
and U21295 (N_21295,N_20321,N_18438);
nor U21296 (N_21296,N_19048,N_18994);
or U21297 (N_21297,N_20080,N_19017);
and U21298 (N_21298,N_19990,N_20475);
xnor U21299 (N_21299,N_20616,N_18409);
nor U21300 (N_21300,N_20297,N_20285);
and U21301 (N_21301,N_18561,N_20803);
or U21302 (N_21302,N_20643,N_19411);
xor U21303 (N_21303,N_18318,N_20671);
xor U21304 (N_21304,N_19376,N_19378);
xor U21305 (N_21305,N_18308,N_20801);
nor U21306 (N_21306,N_19773,N_18344);
xnor U21307 (N_21307,N_18323,N_20891);
and U21308 (N_21308,N_19052,N_19674);
nand U21309 (N_21309,N_19933,N_18129);
or U21310 (N_21310,N_20381,N_20500);
nand U21311 (N_21311,N_18268,N_20071);
and U21312 (N_21312,N_19619,N_20585);
nor U21313 (N_21313,N_18587,N_19153);
nor U21314 (N_21314,N_18951,N_19130);
or U21315 (N_21315,N_19457,N_20481);
nor U21316 (N_21316,N_18259,N_20115);
or U21317 (N_21317,N_18889,N_18442);
and U21318 (N_21318,N_19109,N_19373);
nor U21319 (N_21319,N_18911,N_19566);
xor U21320 (N_21320,N_19670,N_20428);
nor U21321 (N_21321,N_18002,N_19095);
nor U21322 (N_21322,N_18088,N_19618);
nor U21323 (N_21323,N_20411,N_20251);
nand U21324 (N_21324,N_19421,N_18481);
and U21325 (N_21325,N_18946,N_18311);
nor U21326 (N_21326,N_19204,N_18802);
and U21327 (N_21327,N_20875,N_20573);
nand U21328 (N_21328,N_19054,N_19825);
nor U21329 (N_21329,N_20349,N_20458);
xor U21330 (N_21330,N_19744,N_20181);
xnor U21331 (N_21331,N_18142,N_19948);
nand U21332 (N_21332,N_19085,N_20350);
or U21333 (N_21333,N_20824,N_19063);
and U21334 (N_21334,N_19709,N_19737);
nor U21335 (N_21335,N_19414,N_19673);
or U21336 (N_21336,N_19746,N_18163);
and U21337 (N_21337,N_20546,N_20736);
or U21338 (N_21338,N_18457,N_19863);
nor U21339 (N_21339,N_19353,N_19921);
xor U21340 (N_21340,N_18966,N_18941);
nor U21341 (N_21341,N_18685,N_20746);
nor U21342 (N_21342,N_20224,N_19687);
and U21343 (N_21343,N_20244,N_20826);
or U21344 (N_21344,N_18061,N_18441);
or U21345 (N_21345,N_19938,N_19195);
nand U21346 (N_21346,N_20703,N_18029);
xnor U21347 (N_21347,N_20764,N_20612);
xor U21348 (N_21348,N_19772,N_19959);
nand U21349 (N_21349,N_20120,N_20777);
nand U21350 (N_21350,N_19496,N_18701);
nor U21351 (N_21351,N_18178,N_20654);
nand U21352 (N_21352,N_19700,N_20618);
xor U21353 (N_21353,N_19974,N_18832);
nand U21354 (N_21354,N_19393,N_18938);
nor U21355 (N_21355,N_19487,N_19261);
nand U21356 (N_21356,N_19447,N_18104);
nor U21357 (N_21357,N_19337,N_20499);
and U21358 (N_21358,N_18914,N_18046);
or U21359 (N_21359,N_18254,N_18882);
xor U21360 (N_21360,N_18929,N_20629);
or U21361 (N_21361,N_20852,N_20932);
or U21362 (N_21362,N_19947,N_19313);
nor U21363 (N_21363,N_20476,N_20683);
nand U21364 (N_21364,N_19466,N_20264);
and U21365 (N_21365,N_20014,N_19502);
nand U21366 (N_21366,N_20301,N_18673);
nand U21367 (N_21367,N_18188,N_20581);
nand U21368 (N_21368,N_18936,N_20656);
nor U21369 (N_21369,N_20901,N_19796);
or U21370 (N_21370,N_20036,N_18282);
or U21371 (N_21371,N_18024,N_19937);
nand U21372 (N_21372,N_19035,N_18952);
nand U21373 (N_21373,N_20471,N_19066);
xnor U21374 (N_21374,N_20611,N_20085);
or U21375 (N_21375,N_19258,N_19363);
nand U21376 (N_21376,N_19381,N_20735);
nor U21377 (N_21377,N_18255,N_18777);
nand U21378 (N_21378,N_20024,N_18605);
xnor U21379 (N_21379,N_20122,N_19094);
nor U21380 (N_21380,N_18633,N_19603);
or U21381 (N_21381,N_18691,N_19952);
nand U21382 (N_21382,N_19523,N_20950);
and U21383 (N_21383,N_20010,N_20838);
xnor U21384 (N_21384,N_18806,N_19992);
nor U21385 (N_21385,N_19128,N_18484);
and U21386 (N_21386,N_18455,N_19593);
nand U21387 (N_21387,N_20909,N_18751);
and U21388 (N_21388,N_18458,N_19856);
nor U21389 (N_21389,N_18538,N_18189);
nor U21390 (N_21390,N_19537,N_20038);
or U21391 (N_21391,N_19467,N_20180);
nor U21392 (N_21392,N_18834,N_20306);
nand U21393 (N_21393,N_19478,N_20694);
xnor U21394 (N_21394,N_18565,N_18462);
and U21395 (N_21395,N_18102,N_19631);
or U21396 (N_21396,N_18810,N_20152);
and U21397 (N_21397,N_18725,N_20749);
and U21398 (N_21398,N_18843,N_20936);
nor U21399 (N_21399,N_20365,N_19922);
xnor U21400 (N_21400,N_20858,N_18026);
nor U21401 (N_21401,N_20514,N_18250);
nand U21402 (N_21402,N_20984,N_18711);
and U21403 (N_21403,N_20474,N_18126);
or U21404 (N_21404,N_19852,N_19083);
nor U21405 (N_21405,N_19675,N_20382);
nand U21406 (N_21406,N_18977,N_20834);
and U21407 (N_21407,N_20931,N_19433);
nor U21408 (N_21408,N_19386,N_20874);
and U21409 (N_21409,N_19972,N_18432);
xnor U21410 (N_21410,N_20586,N_20172);
nor U21411 (N_21411,N_19323,N_18549);
nor U21412 (N_21412,N_20833,N_19968);
xor U21413 (N_21413,N_18041,N_20661);
nor U21414 (N_21414,N_18225,N_18070);
xnor U21415 (N_21415,N_19374,N_19734);
or U21416 (N_21416,N_20940,N_19835);
nor U21417 (N_21417,N_19238,N_18135);
or U21418 (N_21418,N_20969,N_18612);
or U21419 (N_21419,N_19676,N_20967);
or U21420 (N_21420,N_19629,N_19246);
nand U21421 (N_21421,N_18100,N_18940);
or U21422 (N_21422,N_19324,N_18233);
nand U21423 (N_21423,N_20143,N_20913);
xor U21424 (N_21424,N_18165,N_20033);
or U21425 (N_21425,N_20304,N_19420);
nand U21426 (N_21426,N_19464,N_18170);
and U21427 (N_21427,N_19344,N_19497);
xnor U21428 (N_21428,N_19076,N_18262);
or U21429 (N_21429,N_18478,N_20385);
xnor U21430 (N_21430,N_18383,N_18526);
and U21431 (N_21431,N_19436,N_18400);
nand U21432 (N_21432,N_18209,N_20613);
xor U21433 (N_21433,N_18888,N_20398);
xor U21434 (N_21434,N_19688,N_20890);
nor U21435 (N_21435,N_20744,N_20324);
nand U21436 (N_21436,N_19804,N_19316);
and U21437 (N_21437,N_18919,N_18122);
nor U21438 (N_21438,N_20178,N_20639);
nand U21439 (N_21439,N_20491,N_18412);
or U21440 (N_21440,N_19391,N_20449);
and U21441 (N_21441,N_18842,N_18985);
or U21442 (N_21442,N_18839,N_20387);
and U21443 (N_21443,N_20674,N_19800);
nor U21444 (N_21444,N_20025,N_18891);
xor U21445 (N_21445,N_19451,N_18562);
nand U21446 (N_21446,N_19079,N_20246);
nor U21447 (N_21447,N_18023,N_19799);
and U21448 (N_21448,N_18552,N_19050);
nor U21449 (N_21449,N_18054,N_19215);
nor U21450 (N_21450,N_18085,N_18459);
nor U21451 (N_21451,N_19899,N_19900);
and U21452 (N_21452,N_20059,N_20808);
nand U21453 (N_21453,N_18325,N_19485);
and U21454 (N_21454,N_20392,N_19398);
nor U21455 (N_21455,N_20845,N_18855);
and U21456 (N_21456,N_19369,N_20923);
nand U21457 (N_21457,N_20357,N_18016);
nor U21458 (N_21458,N_18579,N_19350);
nor U21459 (N_21459,N_20621,N_19560);
xor U21460 (N_21460,N_19142,N_19330);
nor U21461 (N_21461,N_18485,N_18520);
nand U21462 (N_21462,N_20066,N_18887);
or U21463 (N_21463,N_20464,N_20829);
and U21464 (N_21464,N_20886,N_18502);
nor U21465 (N_21465,N_19382,N_18297);
xor U21466 (N_21466,N_18048,N_20409);
xnor U21467 (N_21467,N_20980,N_19957);
nand U21468 (N_21468,N_19422,N_19859);
or U21469 (N_21469,N_20571,N_19354);
nor U21470 (N_21470,N_19300,N_18510);
and U21471 (N_21471,N_19555,N_20757);
xor U21472 (N_21472,N_20992,N_18447);
nand U21473 (N_21473,N_18992,N_19958);
or U21474 (N_21474,N_20597,N_20556);
nor U21475 (N_21475,N_20528,N_18999);
nor U21476 (N_21476,N_19144,N_18518);
or U21477 (N_21477,N_18210,N_19625);
and U21478 (N_21478,N_20681,N_19455);
nand U21479 (N_21479,N_18631,N_18064);
nor U21480 (N_21480,N_20961,N_18301);
xor U21481 (N_21481,N_20985,N_19860);
or U21482 (N_21482,N_20088,N_19445);
or U21483 (N_21483,N_18768,N_19504);
nor U21484 (N_21484,N_20790,N_19459);
nand U21485 (N_21485,N_19878,N_20053);
or U21486 (N_21486,N_19007,N_18573);
nor U21487 (N_21487,N_19000,N_19841);
xnor U21488 (N_21488,N_20236,N_19441);
nor U21489 (N_21489,N_18880,N_18586);
or U21490 (N_21490,N_20434,N_19893);
nor U21491 (N_21491,N_18750,N_18156);
nor U21492 (N_21492,N_19462,N_18264);
or U21493 (N_21493,N_18517,N_20679);
xnor U21494 (N_21494,N_18647,N_18030);
nor U21495 (N_21495,N_20635,N_19851);
and U21496 (N_21496,N_18731,N_20388);
nor U21497 (N_21497,N_18143,N_20190);
xnor U21498 (N_21498,N_18551,N_20535);
nand U21499 (N_21499,N_20704,N_19302);
nor U21500 (N_21500,N_18300,N_20316);
nor U21501 (N_21501,N_19465,N_19018);
or U21502 (N_21502,N_18381,N_18266);
xnor U21503 (N_21503,N_19371,N_19339);
and U21504 (N_21504,N_19802,N_18227);
nor U21505 (N_21505,N_18111,N_18407);
or U21506 (N_21506,N_20871,N_19853);
xor U21507 (N_21507,N_20366,N_19172);
nor U21508 (N_21508,N_19716,N_18920);
or U21509 (N_21509,N_19489,N_20337);
xor U21510 (N_21510,N_20800,N_20064);
xor U21511 (N_21511,N_20783,N_19663);
nand U21512 (N_21512,N_18396,N_20102);
or U21513 (N_21513,N_19605,N_20417);
nand U21514 (N_21514,N_20515,N_18576);
xnor U21515 (N_21515,N_20497,N_20228);
and U21516 (N_21516,N_20455,N_19091);
xnor U21517 (N_21517,N_19437,N_20911);
nand U21518 (N_21518,N_20445,N_19834);
xnor U21519 (N_21519,N_19242,N_19110);
and U21520 (N_21520,N_20121,N_19745);
or U21521 (N_21521,N_19400,N_18451);
nand U21522 (N_21522,N_19980,N_18817);
nand U21523 (N_21523,N_20645,N_19029);
nand U21524 (N_21524,N_19059,N_20332);
xnor U21525 (N_21525,N_20907,N_20835);
and U21526 (N_21526,N_19862,N_18971);
or U21527 (N_21527,N_19288,N_20709);
or U21528 (N_21528,N_19089,N_20399);
nor U21529 (N_21529,N_19435,N_18613);
nand U21530 (N_21530,N_18790,N_20019);
xnor U21531 (N_21531,N_19275,N_19672);
and U21532 (N_21532,N_20084,N_19112);
and U21533 (N_21533,N_19838,N_19879);
or U21534 (N_21534,N_19241,N_20666);
nor U21535 (N_21535,N_18798,N_18532);
xor U21536 (N_21536,N_20396,N_20685);
xor U21537 (N_21537,N_18697,N_18515);
xor U21538 (N_21538,N_18546,N_19318);
nand U21539 (N_21539,N_20919,N_19148);
and U21540 (N_21540,N_19472,N_18595);
nor U21541 (N_21541,N_18278,N_19202);
nor U21542 (N_21542,N_19430,N_20168);
nor U21543 (N_21543,N_19319,N_18979);
or U21544 (N_21544,N_20739,N_18487);
nor U21545 (N_21545,N_20864,N_19370);
or U21546 (N_21546,N_19175,N_20899);
xnor U21547 (N_21547,N_18763,N_20116);
or U21548 (N_21548,N_19166,N_18539);
nand U21549 (N_21549,N_18754,N_20154);
xor U21550 (N_21550,N_20128,N_18904);
or U21551 (N_21551,N_20791,N_18616);
xnor U21552 (N_21552,N_19470,N_19989);
and U21553 (N_21553,N_20252,N_19405);
and U21554 (N_21554,N_19536,N_19887);
nor U21555 (N_21555,N_18394,N_20650);
nand U21556 (N_21556,N_18335,N_20092);
nor U21557 (N_21557,N_19902,N_19542);
xor U21558 (N_21558,N_20719,N_20536);
or U21559 (N_21559,N_20097,N_20162);
and U21560 (N_21560,N_19362,N_18548);
nand U21561 (N_21561,N_20112,N_18512);
or U21562 (N_21562,N_20825,N_18893);
nor U21563 (N_21563,N_19585,N_18739);
xor U21564 (N_21564,N_18903,N_18531);
nand U21565 (N_21565,N_19327,N_20897);
nand U21566 (N_21566,N_20311,N_18942);
xor U21567 (N_21567,N_20361,N_20595);
or U21568 (N_21568,N_19650,N_18663);
or U21569 (N_21569,N_20198,N_19134);
and U21570 (N_21570,N_18840,N_19579);
and U21571 (N_21571,N_19871,N_20789);
xnor U21572 (N_21572,N_19812,N_20317);
and U21573 (N_21573,N_20647,N_20233);
and U21574 (N_21574,N_19311,N_20211);
and U21575 (N_21575,N_20917,N_20782);
nand U21576 (N_21576,N_20990,N_20163);
nand U21577 (N_21577,N_18714,N_19192);
and U21578 (N_21578,N_20872,N_20009);
nor U21579 (N_21579,N_19498,N_19304);
nor U21580 (N_21580,N_19160,N_19310);
nor U21581 (N_21581,N_18846,N_19547);
nor U21582 (N_21582,N_18271,N_19614);
nand U21583 (N_21583,N_20781,N_20559);
and U21584 (N_21584,N_20331,N_20713);
nor U21585 (N_21585,N_18186,N_20755);
nand U21586 (N_21586,N_18413,N_20914);
nand U21587 (N_21587,N_18204,N_20139);
and U21588 (N_21588,N_18037,N_19443);
and U21589 (N_21589,N_18815,N_19357);
nand U21590 (N_21590,N_19864,N_19967);
xor U21591 (N_21591,N_20880,N_19100);
or U21592 (N_21592,N_19982,N_20127);
nand U21593 (N_21593,N_20356,N_20949);
and U21594 (N_21594,N_19750,N_18910);
or U21595 (N_21595,N_20590,N_18449);
or U21596 (N_21596,N_18705,N_19197);
xor U21597 (N_21597,N_19219,N_19453);
or U21598 (N_21598,N_20601,N_19020);
or U21599 (N_21599,N_18667,N_18723);
or U21600 (N_21600,N_19582,N_20057);
xor U21601 (N_21601,N_19093,N_19955);
and U21602 (N_21602,N_19577,N_19227);
nand U21603 (N_21603,N_20884,N_19446);
nor U21604 (N_21604,N_19116,N_18395);
nand U21605 (N_21605,N_20982,N_20315);
nor U21606 (N_21606,N_18599,N_20221);
nand U21607 (N_21607,N_19084,N_20199);
and U21608 (N_21608,N_18811,N_18103);
nand U21609 (N_21609,N_20631,N_19413);
and U21610 (N_21610,N_19006,N_20165);
xnor U21611 (N_21611,N_20373,N_18580);
nor U21612 (N_21612,N_18849,N_20933);
nand U21613 (N_21613,N_18463,N_19087);
or U21614 (N_21614,N_18215,N_20793);
xnor U21615 (N_21615,N_19524,N_19755);
nor U21616 (N_21616,N_20173,N_19099);
nor U21617 (N_21617,N_19905,N_20363);
nand U21618 (N_21618,N_20960,N_19070);
nor U21619 (N_21619,N_20988,N_18359);
xnor U21620 (N_21620,N_19763,N_19797);
and U21621 (N_21621,N_18075,N_19490);
nand U21622 (N_21622,N_19730,N_20908);
nor U21623 (N_21623,N_19881,N_18356);
nor U21624 (N_21624,N_20498,N_19789);
or U21625 (N_21625,N_19012,N_19125);
nor U21626 (N_21626,N_18246,N_18422);
or U21627 (N_21627,N_18778,N_19611);
nor U21628 (N_21628,N_19191,N_20269);
and U21629 (N_21629,N_20819,N_20140);
and U21630 (N_21630,N_18939,N_20354);
xnor U21631 (N_21631,N_18908,N_20692);
and U21632 (N_21632,N_18867,N_20840);
xor U21633 (N_21633,N_18597,N_18649);
nor U21634 (N_21634,N_20021,N_19301);
xnor U21635 (N_21635,N_20723,N_20408);
and U21636 (N_21636,N_20690,N_19141);
and U21637 (N_21637,N_20636,N_20395);
nor U21638 (N_21638,N_20107,N_20708);
xnor U21639 (N_21639,N_20489,N_19689);
or U21640 (N_21640,N_20495,N_20044);
nand U21641 (N_21641,N_19298,N_20309);
nand U21642 (N_21642,N_18632,N_19225);
or U21643 (N_21643,N_19877,N_19444);
xnor U21644 (N_21644,N_20176,N_20734);
or U21645 (N_21645,N_19239,N_20484);
nor U21646 (N_21646,N_18136,N_18292);
xor U21647 (N_21647,N_19512,N_19425);
xnor U21648 (N_21648,N_18424,N_19335);
xnor U21649 (N_21649,N_18681,N_19214);
and U21650 (N_21650,N_19460,N_18995);
and U21651 (N_21651,N_20553,N_18726);
nor U21652 (N_21652,N_19569,N_18472);
nor U21653 (N_21653,N_20519,N_18398);
xor U21654 (N_21654,N_19297,N_18523);
xor U21655 (N_21655,N_20979,N_20289);
xor U21656 (N_21656,N_20075,N_20351);
nand U21657 (N_21657,N_20393,N_20624);
xnor U21658 (N_21658,N_18757,N_19179);
or U21659 (N_21659,N_19030,N_19550);
and U21660 (N_21660,N_20662,N_19042);
or U21661 (N_21661,N_19403,N_18659);
xnor U21662 (N_21662,N_20725,N_18053);
or U21663 (N_21663,N_18742,N_18664);
xnor U21664 (N_21664,N_18646,N_19891);
nand U21665 (N_21665,N_20414,N_18245);
nor U21666 (N_21666,N_18575,N_18336);
or U21667 (N_21667,N_20644,N_18230);
nor U21668 (N_21668,N_19969,N_18683);
nand U21669 (N_21669,N_18071,N_18522);
or U21670 (N_21670,N_19133,N_19287);
xnor U21671 (N_21671,N_18131,N_19895);
xor U21672 (N_21672,N_19431,N_20610);
nor U21673 (N_21673,N_18724,N_18758);
xor U21674 (N_21674,N_18062,N_18808);
or U21675 (N_21675,N_20775,N_20527);
nand U21676 (N_21676,N_19210,N_18411);
nor U21677 (N_21677,N_20561,N_18346);
or U21678 (N_21678,N_18997,N_19493);
and U21679 (N_21679,N_19778,N_20175);
or U21680 (N_21680,N_19813,N_20389);
or U21681 (N_21681,N_18362,N_20379);
or U21682 (N_21682,N_18025,N_20432);
and U21683 (N_21683,N_19831,N_20218);
nor U21684 (N_21684,N_20780,N_18113);
xor U21685 (N_21685,N_19936,N_20805);
or U21686 (N_21686,N_18017,N_18201);
xor U21687 (N_21687,N_20663,N_19367);
and U21688 (N_21688,N_20667,N_20817);
nand U21689 (N_21689,N_18372,N_18590);
nor U21690 (N_21690,N_19024,N_19194);
nand U21691 (N_21691,N_19976,N_20836);
xnor U21692 (N_21692,N_20094,N_20370);
xnor U21693 (N_21693,N_18123,N_19452);
xnor U21694 (N_21694,N_20230,N_18547);
or U21695 (N_21695,N_19912,N_20353);
nor U21696 (N_21696,N_18974,N_18378);
xnor U21697 (N_21697,N_18643,N_18563);
and U21698 (N_21698,N_18792,N_20804);
nor U21699 (N_21699,N_20110,N_20888);
nand U21700 (N_21700,N_18217,N_20566);
nor U21701 (N_21701,N_19041,N_18670);
xor U21702 (N_21702,N_20718,N_18615);
nand U21703 (N_21703,N_18375,N_18275);
nand U21704 (N_21704,N_19942,N_18560);
or U21705 (N_21705,N_19685,N_19761);
xnor U21706 (N_21706,N_18086,N_20607);
and U21707 (N_21707,N_20837,N_19690);
nor U21708 (N_21708,N_18040,N_20827);
and U21709 (N_21709,N_18709,N_19875);
nor U21710 (N_21710,N_19695,N_19640);
xor U21711 (N_21711,N_20903,N_18177);
nand U21712 (N_21712,N_18972,N_18013);
nand U21713 (N_21713,N_20039,N_18567);
and U21714 (N_21714,N_18907,N_18600);
and U21715 (N_21715,N_19858,N_20970);
nand U21716 (N_21716,N_19392,N_20000);
xor U21717 (N_21717,N_18001,N_19257);
and U21718 (N_21718,N_18423,N_20422);
xnor U21719 (N_21719,N_18762,N_20061);
xor U21720 (N_21720,N_20552,N_20752);
or U21721 (N_21721,N_20861,N_20249);
or U21722 (N_21722,N_18468,N_19216);
xor U21723 (N_21723,N_19661,N_19118);
xnor U21724 (N_21724,N_20174,N_19349);
and U21725 (N_21725,N_18794,N_19359);
nor U21726 (N_21726,N_20854,N_18376);
and U21727 (N_21727,N_20023,N_19217);
nor U21728 (N_21728,N_19368,N_20910);
or U21729 (N_21729,N_19692,N_19914);
xor U21730 (N_21730,N_18028,N_18693);
and U21731 (N_21731,N_20192,N_19901);
or U21732 (N_21732,N_20453,N_19152);
or U21733 (N_21733,N_19669,N_19519);
and U21734 (N_21734,N_20201,N_20182);
nor U21735 (N_21735,N_18117,N_20450);
and U21736 (N_21736,N_20508,N_18321);
and U21737 (N_21737,N_18436,N_18555);
and U21738 (N_21738,N_18718,N_19997);
xor U21739 (N_21739,N_20340,N_19404);
or U21740 (N_21740,N_18793,N_18544);
xnor U21741 (N_21741,N_20035,N_18760);
nor U21742 (N_21742,N_18084,N_19164);
xnor U21743 (N_21743,N_19637,N_19532);
xor U21744 (N_21744,N_20809,N_18699);
nor U21745 (N_21745,N_18279,N_20216);
nand U21746 (N_21746,N_19571,N_20412);
nor U21747 (N_21747,N_19289,N_19206);
nor U21748 (N_21748,N_20753,N_18765);
nand U21749 (N_21749,N_19668,N_18243);
nor U21750 (N_21750,N_18288,N_18680);
nand U21751 (N_21751,N_19632,N_19609);
xor U21752 (N_21752,N_20254,N_20197);
or U21753 (N_21753,N_18147,N_18015);
or U21754 (N_21754,N_18774,N_20945);
xor U21755 (N_21755,N_18324,N_18453);
and U21756 (N_21756,N_19907,N_19473);
xor U21757 (N_21757,N_19983,N_18124);
xor U21758 (N_21758,N_18249,N_19383);
nand U21759 (N_21759,N_19521,N_19775);
or U21760 (N_21760,N_20051,N_19548);
nor U21761 (N_21761,N_20268,N_20843);
nand U21762 (N_21762,N_19561,N_18421);
xnor U21763 (N_21763,N_20439,N_20150);
xor U21764 (N_21764,N_20415,N_18095);
nand U21765 (N_21765,N_20470,N_20998);
or U21766 (N_21766,N_18729,N_18052);
xnor U21767 (N_21767,N_19401,N_19784);
and U21768 (N_21768,N_18678,N_19283);
and U21769 (N_21769,N_18584,N_18801);
nor U21770 (N_21770,N_18342,N_20855);
nand U21771 (N_21771,N_20818,N_18059);
xnor U21772 (N_21772,N_18187,N_18252);
xor U21773 (N_21773,N_18333,N_20578);
nor U21774 (N_21774,N_19222,N_20844);
and U21775 (N_21775,N_18866,N_18146);
xor U21776 (N_21776,N_18433,N_18752);
nand U21777 (N_21777,N_18044,N_18330);
nor U21778 (N_21778,N_18120,N_19612);
xnor U21779 (N_21779,N_18784,N_20737);
nand U21780 (N_21780,N_18010,N_18417);
xnor U21781 (N_21781,N_18956,N_19586);
xor U21782 (N_21782,N_19157,N_20558);
or U21783 (N_21783,N_18665,N_19424);
xor U21784 (N_21784,N_19442,N_19317);
or U21785 (N_21785,N_18039,N_20605);
or U21786 (N_21786,N_19597,N_19939);
nor U21787 (N_21787,N_20641,N_20292);
or U21788 (N_21788,N_19390,N_19698);
and U21789 (N_21789,N_18826,N_19454);
or U21790 (N_21790,N_19876,N_20490);
xor U21791 (N_21791,N_18619,N_19874);
and U21792 (N_21792,N_20302,N_18895);
nor U21793 (N_21793,N_18689,N_20007);
or U21794 (N_21794,N_18545,N_18686);
nor U21795 (N_21795,N_18732,N_19944);
xnor U21796 (N_21796,N_18392,N_20954);
nor U21797 (N_21797,N_19840,N_20096);
nor U21798 (N_21798,N_19760,N_19691);
xnor U21799 (N_21799,N_20513,N_19634);
xnor U21800 (N_21800,N_19364,N_20747);
xnor U21801 (N_21801,N_20240,N_20563);
and U21802 (N_21802,N_18009,N_20148);
xnor U21803 (N_21803,N_20849,N_18698);
and U21804 (N_21804,N_20589,N_20029);
xnor U21805 (N_21805,N_20894,N_18675);
or U21806 (N_21806,N_19267,N_20788);
xnor U21807 (N_21807,N_18998,N_20664);
and U21808 (N_21808,N_18885,N_20689);
nand U21809 (N_21809,N_20941,N_20283);
nand U21810 (N_21810,N_20687,N_19705);
nor U21811 (N_21811,N_20284,N_20741);
and U21812 (N_21812,N_18830,N_19003);
and U21813 (N_21813,N_19260,N_19266);
and U21814 (N_21814,N_18261,N_19395);
or U21815 (N_21815,N_18197,N_20856);
nor U21816 (N_21816,N_20288,N_20889);
nor U21817 (N_21817,N_19747,N_18014);
nor U21818 (N_21818,N_20360,N_18924);
and U21819 (N_21819,N_18490,N_20766);
nand U21820 (N_21820,N_18863,N_18047);
nand U21821 (N_21821,N_18874,N_19639);
nor U21822 (N_21822,N_20375,N_19058);
xor U21823 (N_21823,N_18671,N_18334);
or U21824 (N_21824,N_18927,N_19492);
xor U21825 (N_21825,N_19770,N_18257);
nor U21826 (N_21826,N_19245,N_19136);
or U21827 (N_21827,N_18764,N_18183);
nor U21828 (N_21828,N_19707,N_20516);
nand U21829 (N_21829,N_18241,N_20892);
or U21830 (N_21830,N_20468,N_20550);
or U21831 (N_21831,N_20786,N_19726);
nor U21832 (N_21832,N_19480,N_19706);
nand U21833 (N_21833,N_20477,N_18466);
or U21834 (N_21834,N_20955,N_20462);
and U21835 (N_21835,N_18899,N_18996);
or U21836 (N_21836,N_20538,N_20670);
or U21837 (N_21837,N_20742,N_20761);
or U21838 (N_21838,N_18949,N_18427);
xnor U21839 (N_21839,N_20567,N_20042);
nand U21840 (N_21840,N_18606,N_19174);
or U21841 (N_21841,N_18355,N_18796);
nor U21842 (N_21842,N_19387,N_20794);
and U21843 (N_21843,N_20569,N_19998);
nor U21844 (N_21844,N_20972,N_18961);
xnor U21845 (N_21845,N_18611,N_19150);
or U21846 (N_21846,N_18614,N_19725);
xor U21847 (N_21847,N_20626,N_18092);
nand U21848 (N_21848,N_18132,N_18875);
xor U21849 (N_21849,N_18007,N_18658);
nand U21850 (N_21850,N_18035,N_19970);
nor U21851 (N_21851,N_19987,N_18640);
and U21852 (N_21852,N_20259,N_19657);
and U21853 (N_21853,N_20814,N_18827);
and U21854 (N_21854,N_20305,N_19865);
xor U21855 (N_21855,N_18137,N_18837);
xor U21856 (N_21856,N_20523,N_20001);
nand U21857 (N_21857,N_19274,N_19751);
xnor U21858 (N_21858,N_19652,N_20454);
nand U21859 (N_21859,N_20189,N_20106);
and U21860 (N_21860,N_20011,N_19165);
and U21861 (N_21861,N_20591,N_19842);
and U21862 (N_21862,N_18682,N_19926);
and U21863 (N_21863,N_18119,N_18299);
or U21864 (N_21864,N_20124,N_19471);
nand U21865 (N_21865,N_18145,N_18101);
nand U21866 (N_21866,N_18629,N_20376);
and U21867 (N_21867,N_20534,N_19185);
and U21868 (N_21868,N_18415,N_19326);
nor U21869 (N_21869,N_19167,N_19132);
or U21870 (N_21870,N_18800,N_20603);
and U21871 (N_21871,N_20625,N_19576);
or U21872 (N_21872,N_18962,N_18668);
xnor U21873 (N_21873,N_20642,N_18004);
xor U21874 (N_21874,N_19665,N_20465);
nand U21875 (N_21875,N_18574,N_20596);
or U21876 (N_21876,N_20145,N_18327);
and U21877 (N_21877,N_20160,N_18981);
nor U21878 (N_21878,N_19078,N_20652);
nand U21879 (N_21879,N_20925,N_18224);
and U21880 (N_21880,N_18216,N_20334);
nor U21881 (N_21881,N_18930,N_18542);
xor U21882 (N_21882,N_20250,N_20660);
and U21883 (N_21883,N_19394,N_19043);
xnor U21884 (N_21884,N_20448,N_18716);
nor U21885 (N_21885,N_20237,N_19022);
xnor U21886 (N_21886,N_20095,N_18389);
nand U21887 (N_21887,N_18289,N_20877);
nor U21888 (N_21888,N_18175,N_20423);
nand U21889 (N_21889,N_20286,N_19633);
and U21890 (N_21890,N_19372,N_18303);
or U21891 (N_21891,N_18034,N_18155);
and U21892 (N_21892,N_20089,N_18169);
nor U21893 (N_21893,N_20740,N_19832);
nor U21894 (N_21894,N_18957,N_19380);
xnor U21895 (N_21895,N_20604,N_20522);
nand U21896 (N_21896,N_19124,N_19565);
xnor U21897 (N_21897,N_19538,N_19996);
nand U21898 (N_21898,N_18737,N_18434);
xor U21899 (N_21899,N_18494,N_18799);
nand U21900 (N_21900,N_20762,N_20503);
xor U21901 (N_21901,N_19979,N_18399);
or U21902 (N_21902,N_20046,N_20822);
or U21903 (N_21903,N_19351,N_20320);
xor U21904 (N_21904,N_20062,N_19090);
and U21905 (N_21905,N_20555,N_19008);
and U21906 (N_21906,N_18696,N_19658);
xnor U21907 (N_21907,N_19505,N_19883);
and U21908 (N_21908,N_18353,N_19483);
nand U21909 (N_21909,N_19945,N_19906);
xor U21910 (N_21910,N_19820,N_19268);
or U21911 (N_21911,N_18819,N_19264);
or U21912 (N_21912,N_19139,N_19540);
and U21913 (N_21913,N_19201,N_19607);
or U21914 (N_21914,N_20502,N_19040);
or U21915 (N_21915,N_19610,N_20707);
nor U21916 (N_21916,N_20815,N_19795);
nor U21917 (N_21917,N_18274,N_20784);
nor U21918 (N_21918,N_20242,N_19649);
and U21919 (N_21919,N_20916,N_20486);
nand U21920 (N_21920,N_19861,N_20657);
xor U21921 (N_21921,N_19417,N_20219);
nor U21922 (N_21922,N_18496,N_20314);
or U21923 (N_21923,N_20287,N_19608);
nor U21924 (N_21924,N_20157,N_18669);
xor U21925 (N_21925,N_20191,N_19693);
nor U21926 (N_21926,N_19299,N_18295);
xnor U21927 (N_21927,N_20587,N_19908);
or U21928 (N_21928,N_18058,N_20821);
nand U21929 (N_21929,N_18181,N_18592);
and U21930 (N_21930,N_18890,N_18367);
nand U21931 (N_21931,N_20328,N_18761);
nor U21932 (N_21932,N_18109,N_20047);
and U21933 (N_21933,N_18180,N_18702);
nor U21934 (N_21934,N_18873,N_19253);
xor U21935 (N_21935,N_19104,N_20394);
or U21936 (N_21936,N_18315,N_20799);
or U21937 (N_21937,N_18231,N_18309);
nand U21938 (N_21938,N_18211,N_18329);
or U21939 (N_21939,N_20693,N_18886);
xor U21940 (N_21940,N_19399,N_19315);
or U21941 (N_21941,N_19923,N_18797);
nor U21942 (N_21942,N_19954,N_19314);
and U21943 (N_21943,N_18008,N_18486);
nor U21944 (N_21944,N_18570,N_20672);
nor U21945 (N_21945,N_20133,N_20371);
or U21946 (N_21946,N_18684,N_20518);
xor U21947 (N_21947,N_20715,N_18540);
nand U21948 (N_21948,N_19056,N_20202);
and U21949 (N_21949,N_19080,N_20430);
or U21950 (N_21950,N_20077,N_20646);
nor U21951 (N_21951,N_19262,N_20946);
and U21952 (N_21952,N_18214,N_20751);
and U21953 (N_21953,N_18514,N_19681);
nor U21954 (N_21954,N_19075,N_19769);
or U21955 (N_21955,N_18328,N_19554);
and U21956 (N_21956,N_18081,N_19559);
and U21957 (N_21957,N_20870,N_19659);
and U21958 (N_21958,N_20405,N_20688);
xnor U21959 (N_21959,N_18205,N_20049);
nor U21960 (N_21960,N_19930,N_18869);
nor U21961 (N_21961,N_18779,N_19525);
xnor U21962 (N_21962,N_18654,N_18499);
nand U21963 (N_21963,N_20981,N_20273);
nand U21964 (N_21964,N_19722,N_19787);
or U21965 (N_21965,N_20333,N_18162);
xor U21966 (N_21966,N_20617,N_19925);
nand U21967 (N_21967,N_19181,N_20205);
nor U21968 (N_21968,N_20529,N_18050);
xnor U21969 (N_21969,N_18530,N_19731);
and U21970 (N_21970,N_19308,N_18571);
or U21971 (N_21971,N_20797,N_18604);
nand U21972 (N_21972,N_19279,N_20153);
or U21973 (N_21973,N_19295,N_18876);
xnor U21974 (N_21974,N_18450,N_19643);
xnor U21975 (N_21975,N_20123,N_20594);
nor U21976 (N_21976,N_20290,N_20303);
and U21977 (N_21977,N_18676,N_20859);
nand U21978 (N_21978,N_19803,N_19293);
and U21979 (N_21979,N_20130,N_18482);
xor U21980 (N_21980,N_19340,N_19280);
or U21981 (N_21981,N_18405,N_19816);
or U21982 (N_21982,N_18193,N_18497);
nor U21983 (N_21983,N_19384,N_19904);
nand U21984 (N_21984,N_19641,N_20003);
nand U21985 (N_21985,N_20034,N_19322);
and U21986 (N_21986,N_19332,N_19517);
or U21987 (N_21987,N_20200,N_18265);
nor U21988 (N_21988,N_19023,N_18340);
and U21989 (N_21989,N_19419,N_20963);
and U21990 (N_21990,N_19599,N_19341);
xnor U21991 (N_21991,N_19823,N_19903);
and U21992 (N_21992,N_19551,N_20125);
or U21993 (N_21993,N_19237,N_20052);
xor U21994 (N_21994,N_19025,N_19015);
nor U21995 (N_21995,N_18964,N_18608);
nand U21996 (N_21996,N_19683,N_18452);
nand U21997 (N_21997,N_19642,N_20291);
xnor U21998 (N_21998,N_19510,N_20577);
xnor U21999 (N_21999,N_20848,N_20367);
nand U22000 (N_22000,N_19786,N_20459);
nor U22001 (N_22001,N_20962,N_20668);
nand U22002 (N_22002,N_20724,N_18019);
and U22003 (N_22003,N_18322,N_20582);
nor U22004 (N_22004,N_20727,N_18783);
and U22005 (N_22005,N_18055,N_19333);
nor U22006 (N_22006,N_19535,N_18769);
or U22007 (N_22007,N_20072,N_18568);
xor U22008 (N_22008,N_19849,N_20391);
xnor U22009 (N_22009,N_19198,N_20137);
and U22010 (N_22010,N_20812,N_20562);
and U22011 (N_22011,N_20469,N_20266);
nor U22012 (N_22012,N_19053,N_20697);
xor U22013 (N_22013,N_18529,N_18553);
xor U22014 (N_22014,N_19033,N_19511);
nor U22015 (N_22015,N_20294,N_19872);
or U22016 (N_22016,N_18622,N_19666);
xor U22017 (N_22017,N_18240,N_20339);
or U22018 (N_22018,N_19870,N_19884);
xnor U22019 (N_22019,N_20710,N_18475);
xor U22020 (N_22020,N_20580,N_19822);
xnor U22021 (N_22021,N_20537,N_20905);
and U22022 (N_22022,N_20952,N_18141);
nand U22023 (N_22023,N_18078,N_18430);
xor U22024 (N_22024,N_18467,N_20701);
nor U22025 (N_22025,N_19163,N_18506);
nor U22026 (N_22026,N_20554,N_18173);
nor U22027 (N_22027,N_19578,N_18583);
and U22028 (N_22028,N_19717,N_20313);
and U22029 (N_22029,N_18069,N_20540);
nor U22030 (N_22030,N_19981,N_20544);
and U22031 (N_22031,N_19598,N_18602);
or U22032 (N_22032,N_20105,N_20135);
and U22033 (N_22033,N_20944,N_19765);
nand U22034 (N_22034,N_20920,N_20005);
or U22035 (N_22035,N_20851,N_20774);
or U22036 (N_22036,N_18352,N_18594);
or U22037 (N_22037,N_18439,N_18199);
xnor U22038 (N_22038,N_19151,N_20512);
or U22039 (N_22039,N_20900,N_19138);
or U22040 (N_22040,N_20179,N_18838);
and U22041 (N_22041,N_19117,N_18861);
nor U22042 (N_22042,N_19793,N_19290);
nor U22043 (N_22043,N_18087,N_18854);
nor U22044 (N_22044,N_19656,N_19739);
xor U22045 (N_22045,N_18912,N_18636);
or U22046 (N_22046,N_18471,N_18305);
and U22047 (N_22047,N_18077,N_18066);
or U22048 (N_22048,N_20857,N_18426);
and U22049 (N_22049,N_20185,N_19591);
nand U22050 (N_22050,N_20017,N_20896);
nor U22051 (N_22051,N_18428,N_19427);
xor U22052 (N_22052,N_18593,N_20229);
xor U22053 (N_22053,N_18982,N_19866);
or U22054 (N_22054,N_19616,N_20609);
and U22055 (N_22055,N_19320,N_18853);
nor U22056 (N_22056,N_20588,N_18805);
and U22057 (N_22057,N_19533,N_19062);
xor U22058 (N_22058,N_18755,N_18218);
nand U22059 (N_22059,N_20748,N_19469);
nand U22060 (N_22060,N_20549,N_18348);
nand U22061 (N_22061,N_18060,N_19740);
nand U22062 (N_22062,N_19975,N_19581);
and U22063 (N_22063,N_19355,N_20419);
xor U22064 (N_22064,N_18980,N_19600);
nand U22065 (N_22065,N_19276,N_19587);
and U22066 (N_22066,N_19966,N_18360);
xor U22067 (N_22067,N_20930,N_18195);
or U22068 (N_22068,N_20069,N_19509);
or U22069 (N_22069,N_19655,N_19183);
nand U22070 (N_22070,N_18079,N_19935);
or U22071 (N_22071,N_18960,N_18020);
xnor U22072 (N_22072,N_18027,N_18238);
nor U22073 (N_22073,N_18883,N_20253);
or U22074 (N_22074,N_18269,N_18272);
or U22075 (N_22075,N_20865,N_18140);
xnor U22076 (N_22076,N_20177,N_19111);
nor U22077 (N_22077,N_20564,N_18021);
nand U22078 (N_22078,N_20231,N_19720);
nor U22079 (N_22079,N_19014,N_18281);
or U22080 (N_22080,N_20298,N_20630);
or U22081 (N_22081,N_20807,N_18814);
nand U22082 (N_22082,N_18291,N_20676);
or U22083 (N_22083,N_18108,N_20754);
xor U22084 (N_22084,N_18959,N_20207);
and U22085 (N_22085,N_19514,N_18978);
or U22086 (N_22086,N_19636,N_20729);
nand U22087 (N_22087,N_20227,N_18740);
or U22088 (N_22088,N_20183,N_20310);
nand U22089 (N_22089,N_19218,N_18851);
and U22090 (N_22090,N_19103,N_18993);
or U22091 (N_22091,N_18114,N_20501);
nand U22092 (N_22092,N_19651,N_20040);
or U22093 (N_22093,N_20686,N_18391);
or U22094 (N_22094,N_19396,N_18965);
xnor U22095 (N_22095,N_20043,N_20606);
xor U22096 (N_22096,N_20473,N_18776);
nand U22097 (N_22097,N_18807,N_20041);
nor U22098 (N_22098,N_18159,N_19388);
and U22099 (N_22099,N_18521,N_19805);
nor U22100 (N_22100,N_18708,N_19097);
xnor U22101 (N_22101,N_20436,N_20760);
nor U22102 (N_22102,N_18504,N_20103);
xor U22103 (N_22103,N_18172,N_20342);
nor U22104 (N_22104,N_19026,N_19406);
nand U22105 (N_22105,N_19171,N_20443);
or U22106 (N_22106,N_19567,N_19810);
nand U22107 (N_22107,N_19077,N_20466);
xnor U22108 (N_22108,N_18307,N_20245);
and U22109 (N_22109,N_18655,N_19941);
and U22110 (N_22110,N_18519,N_19232);
nand U22111 (N_22111,N_19527,N_18203);
or U22112 (N_22112,N_18351,N_19635);
xnor U22113 (N_22113,N_19785,N_18770);
nand U22114 (N_22114,N_19703,N_20206);
nor U22115 (N_22115,N_20507,N_18416);
xnor U22116 (N_22116,N_19615,N_19291);
nor U22117 (N_22117,N_20533,N_19584);
and U22118 (N_22118,N_20927,N_20239);
and U22119 (N_22119,N_18589,N_19544);
nor U22120 (N_22120,N_19910,N_18692);
and U22121 (N_22121,N_18326,N_18712);
and U22122 (N_22122,N_18818,N_18473);
xor U22123 (N_22123,N_20078,N_18384);
xor U22124 (N_22124,N_19699,N_19360);
xor U22125 (N_22125,N_18635,N_20147);
xor U22126 (N_22126,N_18296,N_20658);
or U22127 (N_22127,N_20018,N_18618);
xnor U22128 (N_22128,N_19630,N_19792);
nor U22129 (N_22129,N_19821,N_19682);
nor U22130 (N_22130,N_18191,N_19415);
or U22131 (N_22131,N_18933,N_20384);
or U22132 (N_22132,N_18534,N_18639);
nand U22133 (N_22133,N_18435,N_18239);
nor U22134 (N_22134,N_18152,N_20378);
nand U22135 (N_22135,N_18642,N_19780);
or U22136 (N_22136,N_18042,N_18208);
and U22137 (N_22137,N_19771,N_18115);
nand U22138 (N_22138,N_20364,N_19843);
nand U22139 (N_22139,N_19230,N_19892);
xor U22140 (N_22140,N_18368,N_20444);
nand U22141 (N_22141,N_20557,N_18626);
xnor U22142 (N_22142,N_18337,N_18364);
xor U22143 (N_22143,N_19570,N_18357);
xor U22144 (N_22144,N_20472,N_20876);
nor U22145 (N_22145,N_20702,N_20467);
and U22146 (N_22146,N_20222,N_20008);
nor U22147 (N_22147,N_19919,N_18443);
and U22148 (N_22148,N_19806,N_20275);
nor U22149 (N_22149,N_19440,N_20964);
or U22150 (N_22150,N_19736,N_20093);
nand U22151 (N_22151,N_18780,N_18577);
nor U22152 (N_22152,N_20161,N_19231);
and U22153 (N_22153,N_18533,N_18917);
nor U22154 (N_22154,N_18365,N_18091);
and U22155 (N_22155,N_20355,N_20296);
and U22156 (N_22156,N_19044,N_19263);
xor U22157 (N_22157,N_19060,N_19827);
xor U22158 (N_22158,N_18149,N_18074);
and U22159 (N_22159,N_19620,N_20997);
and U22160 (N_22160,N_18018,N_20058);
or U22161 (N_22161,N_18775,N_19801);
nor U22162 (N_22162,N_20111,N_20779);
nand U22163 (N_22163,N_18379,N_19697);
nor U22164 (N_22164,N_19213,N_19645);
xnor U22165 (N_22165,N_19086,N_18772);
nand U22166 (N_22166,N_19065,N_18624);
nand U22167 (N_22167,N_18049,N_18535);
nor U22168 (N_22168,N_18076,N_19438);
nand U22169 (N_22169,N_19309,N_20583);
nand U22170 (N_22170,N_18313,N_20435);
and U22171 (N_22171,N_19869,N_18710);
or U22172 (N_22172,N_19723,N_18171);
xnor U22173 (N_22173,N_18717,N_20006);
nor U22174 (N_22174,N_18312,N_19494);
and U22175 (N_22175,N_19817,N_18270);
and U22176 (N_22176,N_20717,N_20013);
or U22177 (N_22177,N_19973,N_18090);
and U22178 (N_22178,N_18371,N_19450);
or U22179 (N_22179,N_18374,N_19448);
and U22180 (N_22180,N_19271,N_20144);
and U22181 (N_22181,N_19284,N_20074);
nand U22182 (N_22182,N_18719,N_18258);
nor U22183 (N_22183,N_18226,N_18073);
nor U22184 (N_22184,N_20299,N_19727);
nor U22185 (N_22185,N_19653,N_18674);
nor U22186 (N_22186,N_20265,N_19694);
nor U22187 (N_22187,N_18870,N_20700);
xnor U22188 (N_22188,N_19296,N_20915);
and U22189 (N_22189,N_20731,N_20390);
and U22190 (N_22190,N_19002,N_19752);
nor U22191 (N_22191,N_19644,N_20087);
nor U22192 (N_22192,N_19557,N_20457);
xnor U22193 (N_22193,N_18080,N_19815);
nand U22194 (N_22194,N_19031,N_18314);
or U22195 (N_22195,N_19336,N_20426);
or U22196 (N_22196,N_19146,N_19782);
xor U22197 (N_22197,N_18347,N_18661);
or U22198 (N_22198,N_20773,N_18666);
or U22199 (N_22199,N_19963,N_19994);
xnor U22200 (N_22200,N_18144,N_19847);
nand U22201 (N_22201,N_20055,N_19278);
nor U22202 (N_22202,N_19377,N_18557);
xnor U22203 (N_22203,N_19159,N_18968);
xnor U22204 (N_22204,N_19220,N_18788);
nor U22205 (N_22205,N_19564,N_18429);
and U22206 (N_22206,N_19126,N_19235);
nor U22207 (N_22207,N_18148,N_19211);
nand U22208 (N_22208,N_20649,N_18953);
or U22209 (N_22209,N_18509,N_19176);
xor U22210 (N_22210,N_19412,N_18410);
xor U22211 (N_22211,N_20828,N_20637);
nand U22212 (N_22212,N_20712,N_18641);
nor U22213 (N_22213,N_18234,N_20346);
or U22214 (N_22214,N_20912,N_20126);
xor U22215 (N_22215,N_19735,N_20953);
nor U22216 (N_22216,N_19943,N_19830);
and U22217 (N_22217,N_20060,N_20204);
nor U22218 (N_22218,N_18988,N_20714);
nand U22219 (N_22219,N_19009,N_18598);
and U22220 (N_22220,N_19732,N_19209);
nand U22221 (N_22221,N_20114,N_19259);
nor U22222 (N_22222,N_18005,N_19004);
or U22223 (N_22223,N_18116,N_18828);
nand U22224 (N_22224,N_18068,N_18128);
nor U22225 (N_22225,N_18733,N_20323);
nor U22226 (N_22226,N_18617,N_19092);
xnor U22227 (N_22227,N_18905,N_19286);
or U22228 (N_22228,N_19638,N_20728);
nor U22229 (N_22229,N_19809,N_20863);
nand U22230 (N_22230,N_20869,N_19719);
or U22231 (N_22231,N_18154,N_19129);
nor U22232 (N_22232,N_20217,N_18720);
xnor U22233 (N_22233,N_20347,N_20521);
nor U22234 (N_22234,N_20020,N_20281);
nand U22235 (N_22235,N_20541,N_19305);
nor U22236 (N_22236,N_20068,N_19432);
nor U22237 (N_22237,N_20983,N_18628);
or U22238 (N_22238,N_20608,N_20691);
or U22239 (N_22239,N_18878,N_19229);
xor U22240 (N_22240,N_19426,N_19397);
nand U22241 (N_22241,N_18176,N_19985);
or U22242 (N_22242,N_19187,N_20397);
nor U22243 (N_22243,N_20090,N_20031);
nand U22244 (N_22244,N_19016,N_20256);
nor U22245 (N_22245,N_19724,N_18857);
xor U22246 (N_22246,N_20002,N_20081);
or U22247 (N_22247,N_18160,N_20898);
xor U22248 (N_22248,N_19096,N_19753);
nand U22249 (N_22249,N_18446,N_19074);
or U22250 (N_22250,N_20086,N_20792);
nor U22251 (N_22251,N_19508,N_19468);
nand U22252 (N_22252,N_19098,N_18213);
and U22253 (N_22253,N_19055,N_18454);
or U22254 (N_22254,N_18276,N_18677);
nand U22255 (N_22255,N_19680,N_18516);
nor U22256 (N_22256,N_20721,N_18319);
and U22257 (N_22257,N_20684,N_20404);
and U22258 (N_22258,N_19277,N_19826);
nor U22259 (N_22259,N_19182,N_20948);
nor U22260 (N_22260,N_18862,N_18625);
nand U22261 (N_22261,N_18361,N_19221);
or U22262 (N_22262,N_18363,N_19495);
nand U22263 (N_22263,N_20300,N_20118);
or U22264 (N_22264,N_20485,N_18848);
and U22265 (N_22265,N_20327,N_18852);
nor U22266 (N_22266,N_18825,N_18343);
xnor U22267 (N_22267,N_19728,N_19880);
nand U22268 (N_22268,N_19292,N_19556);
or U22269 (N_22269,N_19212,N_18955);
nor U22270 (N_22270,N_19558,N_19303);
nor U22271 (N_22271,N_20335,N_19439);
nor U22272 (N_22272,N_19984,N_18096);
and U22273 (N_22273,N_19456,N_18556);
xnor U22274 (N_22274,N_18121,N_19503);
xnor U22275 (N_22275,N_18397,N_20325);
xor U22276 (N_22276,N_18493,N_20336);
and U22277 (N_22277,N_19794,N_19484);
and U22278 (N_22278,N_20839,N_19993);
nand U22279 (N_22279,N_18151,N_19819);
xor U22280 (N_22280,N_18461,N_19624);
nand U22281 (N_22281,N_18419,N_19162);
nand U22282 (N_22282,N_19158,N_18174);
xor U22283 (N_22283,N_20151,N_18366);
xor U22284 (N_22284,N_19965,N_19248);
xnor U22285 (N_22285,N_19352,N_19177);
and U22286 (N_22286,N_19082,N_19788);
or U22287 (N_22287,N_18056,N_18093);
nor U22288 (N_22288,N_20109,N_18973);
xnor U22289 (N_22289,N_18420,N_19101);
or U22290 (N_22290,N_18306,N_18652);
nor U22291 (N_22291,N_19890,N_18745);
nand U22292 (N_22292,N_19995,N_20698);
nor U22293 (N_22293,N_20209,N_19917);
and U22294 (N_22294,N_19889,N_18844);
nor U22295 (N_22295,N_20460,N_18388);
nor U22296 (N_22296,N_18370,N_18465);
nor U22297 (N_22297,N_18033,N_19588);
or U22298 (N_22298,N_20326,N_18222);
xor U22299 (N_22299,N_20383,N_20599);
xor U22300 (N_22300,N_18958,N_19366);
nor U22301 (N_22301,N_19779,N_20682);
xor U22302 (N_22302,N_19781,N_18741);
nand U22303 (N_22303,N_19184,N_19885);
or U22304 (N_22304,N_18408,N_20542);
nand U22305 (N_22305,N_18382,N_18634);
and U22306 (N_22306,N_19270,N_20463);
or U22307 (N_22307,N_20214,N_20653);
or U22308 (N_22308,N_20418,N_20816);
xor U22309 (N_22309,N_18789,N_20673);
and U22310 (N_22310,N_20487,N_20492);
or U22311 (N_22311,N_20881,N_19021);
nor U22312 (N_22312,N_19592,N_20271);
xor U22313 (N_22313,N_20441,N_20091);
nand U22314 (N_22314,N_19846,N_18513);
nor U22315 (N_22315,N_20756,N_20022);
nor U22316 (N_22316,N_19173,N_20188);
and U22317 (N_22317,N_19539,N_20402);
xor U22318 (N_22318,N_19928,N_18107);
and U22319 (N_22319,N_18630,N_20260);
nand U22320 (N_22320,N_19949,N_19149);
and U22321 (N_22321,N_18200,N_20407);
xor U22322 (N_22322,N_19848,N_20424);
and U22323 (N_22323,N_18221,N_20975);
xor U22324 (N_22324,N_20100,N_18280);
or U22325 (N_22325,N_20798,N_18856);
xnor U22326 (N_22326,N_18894,N_19045);
and U22327 (N_22327,N_19135,N_20772);
nor U22328 (N_22328,N_18331,N_20358);
and U22329 (N_22329,N_20810,N_19918);
and U22330 (N_22330,N_20440,N_18795);
xor U22331 (N_22331,N_19385,N_20568);
nand U22332 (N_22332,N_18099,N_18833);
nand U22333 (N_22333,N_18700,N_19541);
nand U22334 (N_22334,N_19580,N_20620);
or U22335 (N_22335,N_20421,N_19038);
and U22336 (N_22336,N_20359,N_19776);
and U22337 (N_22337,N_19857,N_18043);
nand U22338 (N_22338,N_19845,N_20496);
and U22339 (N_22339,N_19331,N_18445);
nor U22340 (N_22340,N_18835,N_20212);
xnor U22341 (N_22341,N_18748,N_18603);
nor U22342 (N_22342,N_20131,N_20312);
nand U22343 (N_22343,N_19488,N_20164);
nor U22344 (N_22344,N_19307,N_20208);
or U22345 (N_22345,N_19358,N_19131);
or U22346 (N_22346,N_19946,N_18845);
nor U22347 (N_22347,N_19873,N_18986);
or U22348 (N_22348,N_20243,N_18559);
xor U22349 (N_22349,N_18358,N_19991);
nand U22350 (N_22350,N_19667,N_19956);
and U22351 (N_22351,N_20338,N_19950);
nand U22352 (N_22352,N_19407,N_19064);
xor U22353 (N_22353,N_18369,N_18935);
nor U22354 (N_22354,N_19738,N_18627);
nor U22355 (N_22355,N_19684,N_18704);
nor U22356 (N_22356,N_20280,N_20368);
or U22357 (N_22357,N_20510,N_18158);
xor U22358 (N_22358,N_20372,N_20155);
nand U22359 (N_22359,N_18841,N_19764);
or U22360 (N_22360,N_19613,N_18607);
xor U22361 (N_22361,N_19199,N_19589);
nor U22362 (N_22362,N_18662,N_18161);
nor U22363 (N_22363,N_20758,N_19713);
or U22364 (N_22364,N_20966,N_20628);
or U22365 (N_22365,N_20806,N_18550);
xor U22366 (N_22366,N_20680,N_20846);
and U22367 (N_22367,N_18491,N_18349);
nor U22368 (N_22368,N_18925,N_19312);
nor U22369 (N_22369,N_19122,N_18648);
xor U22370 (N_22370,N_18277,N_20431);
nand U22371 (N_22371,N_19402,N_19929);
or U22372 (N_22372,N_18456,N_18859);
xnor U22373 (N_22373,N_19590,N_20787);
nor U22374 (N_22374,N_18786,N_20832);
xnor U22375 (N_22375,N_19986,N_20600);
xor U22376 (N_22376,N_19071,N_20362);
and U22377 (N_22377,N_20307,N_18804);
xor U22378 (N_22378,N_20548,N_20593);
nand U22379 (N_22379,N_20770,N_19513);
nor U22380 (N_22380,N_18989,N_18350);
or U22381 (N_22381,N_19482,N_18585);
and U22382 (N_22382,N_20293,N_19410);
nor U22383 (N_22383,N_20883,N_20627);
or U22384 (N_22384,N_20427,N_18511);
or U22385 (N_22385,N_18747,N_18715);
nor U22386 (N_22386,N_19073,N_18316);
or U22387 (N_22387,N_19712,N_18133);
or U22388 (N_22388,N_20906,N_18902);
xnor U22389 (N_22389,N_18620,N_18950);
or U22390 (N_22390,N_18645,N_18377);
or U22391 (N_22391,N_20079,N_18219);
or U22392 (N_22392,N_18621,N_18127);
nor U22393 (N_22393,N_18722,N_20996);
nor U22394 (N_22394,N_19186,N_18756);
nor U22395 (N_22395,N_19168,N_18651);
nand U22396 (N_22396,N_19347,N_18380);
nor U22397 (N_22397,N_18229,N_18294);
nand U22398 (N_22398,N_20904,N_20193);
nor U22399 (N_22399,N_18730,N_19428);
xnor U22400 (N_22400,N_20146,N_19646);
xor U22401 (N_22401,N_19529,N_18744);
and U22402 (N_22402,N_19037,N_18483);
or U22403 (N_22403,N_19811,N_18402);
nor U22404 (N_22404,N_19850,N_18588);
and U22405 (N_22405,N_20572,N_19855);
xnor U22406 (N_22406,N_19931,N_19343);
nand U22407 (N_22407,N_18983,N_20171);
nor U22408 (N_22408,N_20026,N_20971);
nand U22409 (N_22409,N_19601,N_20138);
xor U22410 (N_22410,N_19623,N_19285);
and U22411 (N_22411,N_19961,N_19824);
or U22412 (N_22412,N_20104,N_19325);
xnor U22413 (N_22413,N_20480,N_19190);
nor U22414 (N_22414,N_18166,N_18877);
nand U22415 (N_22415,N_19180,N_19520);
nand U22416 (N_22416,N_20675,N_18836);
nor U22417 (N_22417,N_19475,N_20669);
xnor U22418 (N_22418,N_18168,N_18672);
nor U22419 (N_22419,N_20934,N_19234);
nand U22420 (N_22420,N_19924,N_18317);
and U22421 (N_22421,N_20451,N_20223);
and U22422 (N_22422,N_20504,N_20831);
and U22423 (N_22423,N_20866,N_19039);
or U22424 (N_22424,N_18609,N_20027);
and U22425 (N_22425,N_18984,N_18991);
and U22426 (N_22426,N_20956,N_20267);
or U22427 (N_22427,N_18404,N_18320);
and U22428 (N_22428,N_19223,N_19506);
nand U22429 (N_22429,N_18498,N_18130);
nand U22430 (N_22430,N_18332,N_19777);
or U22431 (N_22431,N_18290,N_18251);
nor U22432 (N_22432,N_18284,N_18566);
and U22433 (N_22433,N_19583,N_19281);
nand U22434 (N_22434,N_18975,N_18536);
or U22435 (N_22435,N_19766,N_18440);
nor U22436 (N_22436,N_20166,N_19499);
nor U22437 (N_22437,N_19671,N_20862);
xnor U22438 (N_22438,N_20270,N_18990);
nor U22439 (N_22439,N_20995,N_19013);
nand U22440 (N_22440,N_20184,N_18728);
nor U22441 (N_22441,N_19356,N_18373);
nand U22442 (N_22442,N_19408,N_18285);
nor U22443 (N_22443,N_20977,N_20938);
and U22444 (N_22444,N_19207,N_20796);
nand U22445 (N_22445,N_19072,N_18638);
and U22446 (N_22446,N_18488,N_20410);
and U22447 (N_22447,N_20765,N_20015);
xor U22448 (N_22448,N_19155,N_19034);
and U22449 (N_22449,N_18823,N_18110);
and U22450 (N_22450,N_19254,N_19361);
nand U22451 (N_22451,N_18947,N_20763);
xor U22452 (N_22452,N_20551,N_18970);
or U22453 (N_22453,N_19606,N_18167);
or U22454 (N_22454,N_20615,N_19113);
nor U22455 (N_22455,N_18474,N_20156);
nor U22456 (N_22456,N_18500,N_20159);
and U22457 (N_22457,N_18746,N_19247);
or U22458 (N_22458,N_20247,N_20054);
nor U22459 (N_22459,N_18637,N_20235);
xor U22460 (N_22460,N_18813,N_20067);
nand U22461 (N_22461,N_18865,N_19228);
nor U22462 (N_22462,N_20745,N_20937);
and U22463 (N_22463,N_18707,N_19068);
nor U22464 (N_22464,N_18464,N_19005);
or U22465 (N_22465,N_18864,N_19236);
nor U22466 (N_22466,N_18932,N_18431);
nand U22467 (N_22467,N_20413,N_18860);
nor U22468 (N_22468,N_20942,N_20261);
and U22469 (N_22469,N_19306,N_18489);
or U22470 (N_22470,N_18105,N_19178);
and U22471 (N_22471,N_18706,N_20974);
or U22472 (N_22472,N_20505,N_20509);
nand U22473 (N_22473,N_18735,N_19226);
nand U22474 (N_22474,N_20750,N_20279);
xor U22475 (N_22475,N_19477,N_20991);
xnor U22476 (N_22476,N_20633,N_19913);
nor U22477 (N_22477,N_18660,N_20226);
or U22478 (N_22478,N_19249,N_20699);
or U22479 (N_22479,N_20659,N_19127);
and U22480 (N_22480,N_19069,N_19868);
or U22481 (N_22481,N_18207,N_19563);
nand U22482 (N_22482,N_18721,N_18753);
xnor U22483 (N_22483,N_19748,N_20263);
and U22484 (N_22484,N_18386,N_19702);
nor U22485 (N_22485,N_19481,N_19032);
and U22486 (N_22486,N_19203,N_20213);
xnor U22487 (N_22487,N_20987,N_18118);
nor U22488 (N_22488,N_18926,N_19718);
nor U22489 (N_22489,N_18858,N_18036);
and U22490 (N_22490,N_19721,N_20677);
or U22491 (N_22491,N_20640,N_18082);
xnor U22492 (N_22492,N_19463,N_18038);
or U22493 (N_22493,N_19156,N_19549);
and U22494 (N_22494,N_18267,N_20547);
xnor U22495 (N_22495,N_20830,N_19837);
and U22496 (N_22496,N_20520,N_20262);
or U22497 (N_22497,N_19334,N_18881);
xnor U22498 (N_22498,N_18273,N_18850);
or U22499 (N_22499,N_20543,N_18338);
or U22500 (N_22500,N_18716,N_19480);
and U22501 (N_22501,N_18378,N_19718);
or U22502 (N_22502,N_19553,N_19772);
xnor U22503 (N_22503,N_20274,N_18575);
and U22504 (N_22504,N_18869,N_18997);
nand U22505 (N_22505,N_19369,N_20342);
nor U22506 (N_22506,N_18189,N_20664);
and U22507 (N_22507,N_19024,N_19670);
xor U22508 (N_22508,N_20954,N_20809);
or U22509 (N_22509,N_18127,N_19068);
and U22510 (N_22510,N_20378,N_19880);
nor U22511 (N_22511,N_20577,N_20470);
and U22512 (N_22512,N_20813,N_19027);
nor U22513 (N_22513,N_20589,N_20517);
nand U22514 (N_22514,N_18350,N_18566);
and U22515 (N_22515,N_19662,N_19480);
or U22516 (N_22516,N_20406,N_20886);
nor U22517 (N_22517,N_19080,N_19309);
nand U22518 (N_22518,N_19889,N_18959);
nand U22519 (N_22519,N_18125,N_20591);
and U22520 (N_22520,N_19699,N_18928);
and U22521 (N_22521,N_19105,N_18728);
nor U22522 (N_22522,N_18047,N_18877);
nor U22523 (N_22523,N_20328,N_19618);
xnor U22524 (N_22524,N_19582,N_18770);
nor U22525 (N_22525,N_18204,N_18643);
nor U22526 (N_22526,N_18403,N_20960);
nand U22527 (N_22527,N_20011,N_20233);
nor U22528 (N_22528,N_19270,N_18220);
nor U22529 (N_22529,N_19188,N_19342);
nor U22530 (N_22530,N_20280,N_18620);
nand U22531 (N_22531,N_19384,N_19819);
or U22532 (N_22532,N_18862,N_20132);
or U22533 (N_22533,N_18935,N_19776);
or U22534 (N_22534,N_19592,N_18291);
nand U22535 (N_22535,N_20159,N_18643);
nand U22536 (N_22536,N_18679,N_20271);
or U22537 (N_22537,N_18410,N_20714);
nor U22538 (N_22538,N_19291,N_19940);
xor U22539 (N_22539,N_20512,N_20079);
and U22540 (N_22540,N_18132,N_18959);
nor U22541 (N_22541,N_20884,N_19929);
and U22542 (N_22542,N_18293,N_20228);
or U22543 (N_22543,N_19115,N_18687);
or U22544 (N_22544,N_20161,N_20203);
xor U22545 (N_22545,N_20815,N_18368);
and U22546 (N_22546,N_19375,N_19031);
or U22547 (N_22547,N_20393,N_18076);
xnor U22548 (N_22548,N_20530,N_18322);
xor U22549 (N_22549,N_18489,N_20771);
and U22550 (N_22550,N_18758,N_18046);
or U22551 (N_22551,N_19459,N_18665);
nand U22552 (N_22552,N_20179,N_20566);
and U22553 (N_22553,N_19425,N_19622);
or U22554 (N_22554,N_19800,N_20160);
nand U22555 (N_22555,N_18340,N_20780);
and U22556 (N_22556,N_18965,N_20551);
nand U22557 (N_22557,N_20485,N_20583);
nor U22558 (N_22558,N_18997,N_19109);
xnor U22559 (N_22559,N_19661,N_18103);
xor U22560 (N_22560,N_20790,N_20110);
or U22561 (N_22561,N_19613,N_20877);
or U22562 (N_22562,N_20157,N_18110);
nor U22563 (N_22563,N_19228,N_19473);
nand U22564 (N_22564,N_18080,N_20954);
or U22565 (N_22565,N_20637,N_20480);
or U22566 (N_22566,N_19834,N_19646);
nand U22567 (N_22567,N_18132,N_20623);
nor U22568 (N_22568,N_19229,N_20532);
and U22569 (N_22569,N_20508,N_20776);
nand U22570 (N_22570,N_20685,N_19681);
nand U22571 (N_22571,N_18063,N_18880);
or U22572 (N_22572,N_18000,N_19048);
or U22573 (N_22573,N_18932,N_19787);
and U22574 (N_22574,N_19096,N_19625);
and U22575 (N_22575,N_20124,N_18269);
nor U22576 (N_22576,N_18802,N_19187);
xnor U22577 (N_22577,N_19485,N_20990);
xnor U22578 (N_22578,N_20936,N_20057);
nor U22579 (N_22579,N_19281,N_18933);
nor U22580 (N_22580,N_18203,N_18248);
or U22581 (N_22581,N_20445,N_18243);
and U22582 (N_22582,N_19401,N_18483);
and U22583 (N_22583,N_18287,N_19297);
nor U22584 (N_22584,N_18666,N_20555);
nor U22585 (N_22585,N_20875,N_20646);
xor U22586 (N_22586,N_20767,N_20973);
nor U22587 (N_22587,N_19139,N_20426);
nand U22588 (N_22588,N_18485,N_18240);
nand U22589 (N_22589,N_19312,N_18980);
or U22590 (N_22590,N_20505,N_20567);
nor U22591 (N_22591,N_19608,N_18708);
nand U22592 (N_22592,N_20102,N_19011);
nand U22593 (N_22593,N_20601,N_18443);
and U22594 (N_22594,N_18558,N_18164);
nor U22595 (N_22595,N_19961,N_18737);
xor U22596 (N_22596,N_20579,N_19022);
and U22597 (N_22597,N_19999,N_18578);
nor U22598 (N_22598,N_19486,N_18189);
and U22599 (N_22599,N_19440,N_20513);
nor U22600 (N_22600,N_18972,N_19359);
xor U22601 (N_22601,N_19720,N_19162);
and U22602 (N_22602,N_19234,N_20242);
nor U22603 (N_22603,N_20899,N_19219);
nor U22604 (N_22604,N_19474,N_18329);
nor U22605 (N_22605,N_20380,N_20678);
nand U22606 (N_22606,N_19234,N_20486);
or U22607 (N_22607,N_19916,N_18602);
xor U22608 (N_22608,N_20167,N_18708);
and U22609 (N_22609,N_18512,N_20912);
or U22610 (N_22610,N_20968,N_18414);
nor U22611 (N_22611,N_18259,N_19360);
nand U22612 (N_22612,N_19297,N_18899);
and U22613 (N_22613,N_18535,N_19329);
nand U22614 (N_22614,N_18523,N_18385);
nor U22615 (N_22615,N_18501,N_19576);
nor U22616 (N_22616,N_18133,N_20686);
and U22617 (N_22617,N_20553,N_20776);
and U22618 (N_22618,N_18817,N_20390);
nand U22619 (N_22619,N_20833,N_18616);
nand U22620 (N_22620,N_18306,N_20708);
nor U22621 (N_22621,N_20129,N_20153);
or U22622 (N_22622,N_20833,N_20712);
nor U22623 (N_22623,N_19321,N_19240);
xor U22624 (N_22624,N_20415,N_19606);
xnor U22625 (N_22625,N_18605,N_18200);
nor U22626 (N_22626,N_20629,N_18939);
or U22627 (N_22627,N_20078,N_18675);
nand U22628 (N_22628,N_18504,N_18303);
nand U22629 (N_22629,N_19095,N_19283);
nor U22630 (N_22630,N_20342,N_19660);
or U22631 (N_22631,N_19958,N_18683);
xor U22632 (N_22632,N_20971,N_18339);
nand U22633 (N_22633,N_18241,N_20910);
or U22634 (N_22634,N_18355,N_20239);
or U22635 (N_22635,N_19796,N_18751);
xnor U22636 (N_22636,N_18449,N_18290);
xnor U22637 (N_22637,N_18406,N_19156);
xor U22638 (N_22638,N_18654,N_18063);
xnor U22639 (N_22639,N_20034,N_18050);
xnor U22640 (N_22640,N_20702,N_18416);
nand U22641 (N_22641,N_20615,N_19473);
or U22642 (N_22642,N_19396,N_20901);
nand U22643 (N_22643,N_19367,N_19720);
and U22644 (N_22644,N_19994,N_18411);
xnor U22645 (N_22645,N_18149,N_18847);
xor U22646 (N_22646,N_20044,N_20809);
nor U22647 (N_22647,N_19469,N_18235);
nand U22648 (N_22648,N_20324,N_19944);
or U22649 (N_22649,N_18902,N_19907);
nand U22650 (N_22650,N_18249,N_20394);
or U22651 (N_22651,N_19362,N_20586);
and U22652 (N_22652,N_20173,N_19734);
xor U22653 (N_22653,N_20598,N_20658);
and U22654 (N_22654,N_18878,N_20060);
nor U22655 (N_22655,N_20841,N_19834);
xnor U22656 (N_22656,N_19742,N_20247);
xnor U22657 (N_22657,N_20740,N_18753);
or U22658 (N_22658,N_20405,N_19166);
or U22659 (N_22659,N_20405,N_19606);
nand U22660 (N_22660,N_18102,N_19989);
and U22661 (N_22661,N_19452,N_18893);
or U22662 (N_22662,N_18437,N_19423);
nor U22663 (N_22663,N_20726,N_20177);
nand U22664 (N_22664,N_20965,N_19786);
and U22665 (N_22665,N_20558,N_19468);
or U22666 (N_22666,N_20873,N_19161);
xor U22667 (N_22667,N_20084,N_18891);
xnor U22668 (N_22668,N_19299,N_18638);
xor U22669 (N_22669,N_18859,N_19255);
nor U22670 (N_22670,N_20384,N_20306);
nand U22671 (N_22671,N_19560,N_19092);
xnor U22672 (N_22672,N_19015,N_20361);
nor U22673 (N_22673,N_19709,N_18131);
and U22674 (N_22674,N_19491,N_20631);
xnor U22675 (N_22675,N_19467,N_20574);
nor U22676 (N_22676,N_19495,N_19985);
nand U22677 (N_22677,N_19413,N_18465);
or U22678 (N_22678,N_20670,N_20589);
or U22679 (N_22679,N_20034,N_18709);
and U22680 (N_22680,N_19880,N_19551);
and U22681 (N_22681,N_18347,N_18537);
nand U22682 (N_22682,N_18384,N_20297);
nand U22683 (N_22683,N_20607,N_18722);
and U22684 (N_22684,N_19737,N_18063);
and U22685 (N_22685,N_18565,N_19958);
nand U22686 (N_22686,N_20232,N_19775);
nand U22687 (N_22687,N_18343,N_18679);
or U22688 (N_22688,N_18051,N_19535);
xnor U22689 (N_22689,N_18580,N_18597);
nor U22690 (N_22690,N_18511,N_19400);
and U22691 (N_22691,N_18595,N_19942);
and U22692 (N_22692,N_18487,N_20320);
and U22693 (N_22693,N_20008,N_19060);
nor U22694 (N_22694,N_18781,N_19090);
nor U22695 (N_22695,N_18632,N_20981);
xor U22696 (N_22696,N_20742,N_19446);
nand U22697 (N_22697,N_18195,N_20651);
or U22698 (N_22698,N_19465,N_20323);
or U22699 (N_22699,N_18392,N_18472);
or U22700 (N_22700,N_18837,N_18724);
and U22701 (N_22701,N_20934,N_18968);
nor U22702 (N_22702,N_20401,N_20864);
nor U22703 (N_22703,N_20210,N_20988);
and U22704 (N_22704,N_20736,N_20880);
nand U22705 (N_22705,N_20925,N_20213);
or U22706 (N_22706,N_19707,N_18332);
nor U22707 (N_22707,N_19417,N_18609);
and U22708 (N_22708,N_20339,N_18760);
nor U22709 (N_22709,N_20251,N_19677);
nand U22710 (N_22710,N_19450,N_18781);
nor U22711 (N_22711,N_18029,N_19256);
nor U22712 (N_22712,N_18793,N_18041);
nor U22713 (N_22713,N_18020,N_18348);
xnor U22714 (N_22714,N_18292,N_19738);
nor U22715 (N_22715,N_18412,N_18883);
or U22716 (N_22716,N_20647,N_19628);
or U22717 (N_22717,N_19756,N_20431);
and U22718 (N_22718,N_18709,N_18133);
or U22719 (N_22719,N_18456,N_19627);
xnor U22720 (N_22720,N_19999,N_20937);
xor U22721 (N_22721,N_19361,N_19983);
nor U22722 (N_22722,N_19363,N_20563);
or U22723 (N_22723,N_20650,N_19023);
and U22724 (N_22724,N_20381,N_19043);
xnor U22725 (N_22725,N_18701,N_19766);
nor U22726 (N_22726,N_19516,N_19730);
or U22727 (N_22727,N_18924,N_20721);
nand U22728 (N_22728,N_19122,N_19832);
or U22729 (N_22729,N_19630,N_18584);
xor U22730 (N_22730,N_19077,N_18406);
and U22731 (N_22731,N_19389,N_19113);
or U22732 (N_22732,N_19997,N_20315);
xnor U22733 (N_22733,N_19755,N_18366);
nand U22734 (N_22734,N_20582,N_18282);
xor U22735 (N_22735,N_19787,N_19774);
xor U22736 (N_22736,N_19848,N_20125);
nand U22737 (N_22737,N_18205,N_18474);
xor U22738 (N_22738,N_20142,N_18422);
nand U22739 (N_22739,N_18508,N_19998);
nand U22740 (N_22740,N_20165,N_20431);
xor U22741 (N_22741,N_19107,N_18968);
nor U22742 (N_22742,N_20377,N_18485);
nand U22743 (N_22743,N_18387,N_19577);
nor U22744 (N_22744,N_20740,N_20403);
xor U22745 (N_22745,N_19567,N_20152);
or U22746 (N_22746,N_20836,N_19222);
or U22747 (N_22747,N_19862,N_20280);
or U22748 (N_22748,N_18672,N_18491);
or U22749 (N_22749,N_18507,N_19856);
and U22750 (N_22750,N_19423,N_19047);
nor U22751 (N_22751,N_19101,N_19436);
or U22752 (N_22752,N_20381,N_20109);
or U22753 (N_22753,N_19839,N_19223);
nor U22754 (N_22754,N_19572,N_19795);
or U22755 (N_22755,N_19676,N_19054);
xor U22756 (N_22756,N_18801,N_18762);
nor U22757 (N_22757,N_18456,N_18903);
or U22758 (N_22758,N_19467,N_18870);
xnor U22759 (N_22759,N_18301,N_18202);
xor U22760 (N_22760,N_20599,N_19340);
nor U22761 (N_22761,N_19188,N_18449);
nor U22762 (N_22762,N_20702,N_18145);
and U22763 (N_22763,N_18711,N_19487);
xnor U22764 (N_22764,N_20570,N_18228);
and U22765 (N_22765,N_20397,N_20859);
or U22766 (N_22766,N_19886,N_19281);
and U22767 (N_22767,N_18438,N_18413);
or U22768 (N_22768,N_20426,N_18925);
nor U22769 (N_22769,N_19685,N_20971);
or U22770 (N_22770,N_19552,N_18027);
and U22771 (N_22771,N_20243,N_19729);
xnor U22772 (N_22772,N_20858,N_18537);
xnor U22773 (N_22773,N_20630,N_20524);
or U22774 (N_22774,N_19430,N_20571);
or U22775 (N_22775,N_20893,N_18687);
nor U22776 (N_22776,N_20969,N_18122);
or U22777 (N_22777,N_20426,N_19434);
or U22778 (N_22778,N_20091,N_20292);
nand U22779 (N_22779,N_18263,N_20631);
or U22780 (N_22780,N_18946,N_20968);
xor U22781 (N_22781,N_20217,N_20533);
nand U22782 (N_22782,N_20452,N_19898);
xor U22783 (N_22783,N_19403,N_18782);
xor U22784 (N_22784,N_18513,N_20895);
or U22785 (N_22785,N_18322,N_18529);
nand U22786 (N_22786,N_20075,N_20080);
xor U22787 (N_22787,N_19148,N_18135);
nand U22788 (N_22788,N_19513,N_20313);
nor U22789 (N_22789,N_18804,N_19365);
xor U22790 (N_22790,N_19157,N_20186);
nor U22791 (N_22791,N_20336,N_19741);
xor U22792 (N_22792,N_18786,N_19437);
and U22793 (N_22793,N_18272,N_19932);
nor U22794 (N_22794,N_19433,N_19938);
and U22795 (N_22795,N_18867,N_20732);
and U22796 (N_22796,N_19848,N_18938);
nor U22797 (N_22797,N_19970,N_20588);
xor U22798 (N_22798,N_18626,N_19026);
nor U22799 (N_22799,N_20166,N_18598);
and U22800 (N_22800,N_20977,N_20986);
and U22801 (N_22801,N_20857,N_18104);
nand U22802 (N_22802,N_20750,N_19846);
nor U22803 (N_22803,N_19018,N_18512);
nor U22804 (N_22804,N_18840,N_20855);
nand U22805 (N_22805,N_20852,N_20986);
nor U22806 (N_22806,N_18117,N_20072);
or U22807 (N_22807,N_18058,N_20616);
nor U22808 (N_22808,N_18504,N_19546);
nor U22809 (N_22809,N_18387,N_19040);
xnor U22810 (N_22810,N_18316,N_20081);
xor U22811 (N_22811,N_20632,N_20682);
nor U22812 (N_22812,N_19952,N_20481);
or U22813 (N_22813,N_19838,N_18013);
or U22814 (N_22814,N_20810,N_18340);
or U22815 (N_22815,N_20573,N_20407);
and U22816 (N_22816,N_19180,N_20969);
nand U22817 (N_22817,N_20825,N_19461);
nor U22818 (N_22818,N_20083,N_19116);
and U22819 (N_22819,N_20675,N_19433);
nor U22820 (N_22820,N_20590,N_18310);
and U22821 (N_22821,N_19721,N_18727);
xnor U22822 (N_22822,N_20541,N_19886);
xnor U22823 (N_22823,N_18111,N_20546);
nand U22824 (N_22824,N_18644,N_20699);
nand U22825 (N_22825,N_18094,N_18913);
or U22826 (N_22826,N_18588,N_18447);
and U22827 (N_22827,N_19132,N_20062);
or U22828 (N_22828,N_20840,N_18130);
xor U22829 (N_22829,N_18790,N_18483);
and U22830 (N_22830,N_18695,N_19736);
nor U22831 (N_22831,N_18539,N_19517);
or U22832 (N_22832,N_20680,N_19434);
or U22833 (N_22833,N_18001,N_18552);
nor U22834 (N_22834,N_18857,N_20909);
and U22835 (N_22835,N_18484,N_20616);
and U22836 (N_22836,N_19631,N_18088);
nand U22837 (N_22837,N_19094,N_20245);
or U22838 (N_22838,N_18869,N_18838);
nor U22839 (N_22839,N_18350,N_20249);
or U22840 (N_22840,N_18968,N_20696);
xor U22841 (N_22841,N_20929,N_18332);
nor U22842 (N_22842,N_18738,N_19792);
and U22843 (N_22843,N_20961,N_19993);
nor U22844 (N_22844,N_19647,N_18949);
or U22845 (N_22845,N_20116,N_19898);
and U22846 (N_22846,N_20057,N_20526);
nor U22847 (N_22847,N_18807,N_20678);
nor U22848 (N_22848,N_20095,N_20752);
or U22849 (N_22849,N_19567,N_20361);
and U22850 (N_22850,N_19906,N_18136);
nand U22851 (N_22851,N_20829,N_20838);
nand U22852 (N_22852,N_20676,N_19148);
nand U22853 (N_22853,N_18031,N_20755);
or U22854 (N_22854,N_19358,N_18565);
xnor U22855 (N_22855,N_19620,N_19543);
nand U22856 (N_22856,N_18987,N_20011);
nor U22857 (N_22857,N_20022,N_20596);
xnor U22858 (N_22858,N_19978,N_19213);
or U22859 (N_22859,N_19358,N_19799);
nand U22860 (N_22860,N_18356,N_20268);
nor U22861 (N_22861,N_18808,N_20156);
xnor U22862 (N_22862,N_19894,N_19918);
nor U22863 (N_22863,N_20693,N_18703);
nand U22864 (N_22864,N_20726,N_20568);
nor U22865 (N_22865,N_18898,N_18961);
nor U22866 (N_22866,N_19293,N_19419);
xnor U22867 (N_22867,N_20422,N_19513);
and U22868 (N_22868,N_18708,N_19813);
nor U22869 (N_22869,N_19555,N_19116);
xor U22870 (N_22870,N_18205,N_19454);
or U22871 (N_22871,N_18204,N_18891);
or U22872 (N_22872,N_18528,N_19363);
xnor U22873 (N_22873,N_18501,N_20893);
xor U22874 (N_22874,N_18652,N_18811);
and U22875 (N_22875,N_20191,N_18827);
nand U22876 (N_22876,N_19900,N_20780);
and U22877 (N_22877,N_20057,N_19144);
or U22878 (N_22878,N_18752,N_18908);
and U22879 (N_22879,N_18225,N_19246);
and U22880 (N_22880,N_20506,N_19026);
or U22881 (N_22881,N_19460,N_19429);
nor U22882 (N_22882,N_19574,N_18464);
and U22883 (N_22883,N_20399,N_20184);
and U22884 (N_22884,N_18635,N_19265);
xor U22885 (N_22885,N_19658,N_20892);
and U22886 (N_22886,N_20420,N_19505);
nand U22887 (N_22887,N_18019,N_18819);
xnor U22888 (N_22888,N_18461,N_20671);
nand U22889 (N_22889,N_19852,N_18450);
xor U22890 (N_22890,N_19781,N_19715);
and U22891 (N_22891,N_18401,N_18113);
nor U22892 (N_22892,N_20459,N_18985);
nor U22893 (N_22893,N_18243,N_20781);
xnor U22894 (N_22894,N_20201,N_18786);
or U22895 (N_22895,N_18922,N_20613);
or U22896 (N_22896,N_19782,N_18215);
nor U22897 (N_22897,N_20670,N_20327);
nand U22898 (N_22898,N_20104,N_18862);
nand U22899 (N_22899,N_18537,N_20322);
and U22900 (N_22900,N_19297,N_19700);
nand U22901 (N_22901,N_18711,N_19206);
nor U22902 (N_22902,N_20902,N_20052);
and U22903 (N_22903,N_20596,N_18617);
or U22904 (N_22904,N_19312,N_18539);
nor U22905 (N_22905,N_19416,N_20003);
and U22906 (N_22906,N_18595,N_18850);
and U22907 (N_22907,N_18799,N_18012);
nor U22908 (N_22908,N_20582,N_18080);
nand U22909 (N_22909,N_19655,N_20165);
nand U22910 (N_22910,N_19621,N_18896);
nor U22911 (N_22911,N_20130,N_18095);
nor U22912 (N_22912,N_19656,N_20429);
nor U22913 (N_22913,N_19288,N_18964);
nand U22914 (N_22914,N_20631,N_18743);
or U22915 (N_22915,N_18166,N_18181);
and U22916 (N_22916,N_18157,N_18348);
and U22917 (N_22917,N_20237,N_19228);
nand U22918 (N_22918,N_20403,N_19924);
or U22919 (N_22919,N_18840,N_19775);
nand U22920 (N_22920,N_19520,N_20757);
nand U22921 (N_22921,N_19679,N_19409);
nand U22922 (N_22922,N_19273,N_20716);
or U22923 (N_22923,N_19588,N_19943);
xor U22924 (N_22924,N_18126,N_20613);
nand U22925 (N_22925,N_20679,N_19591);
xnor U22926 (N_22926,N_18661,N_18418);
nor U22927 (N_22927,N_18711,N_20643);
or U22928 (N_22928,N_18663,N_19529);
xnor U22929 (N_22929,N_19108,N_18416);
and U22930 (N_22930,N_18710,N_19508);
or U22931 (N_22931,N_20566,N_18622);
and U22932 (N_22932,N_20654,N_19135);
xnor U22933 (N_22933,N_20511,N_19280);
nor U22934 (N_22934,N_19691,N_19271);
nand U22935 (N_22935,N_20579,N_19077);
and U22936 (N_22936,N_20401,N_20251);
nand U22937 (N_22937,N_18636,N_18695);
or U22938 (N_22938,N_20702,N_20669);
nor U22939 (N_22939,N_18854,N_18464);
nand U22940 (N_22940,N_20277,N_20825);
or U22941 (N_22941,N_20940,N_18670);
or U22942 (N_22942,N_18816,N_19150);
and U22943 (N_22943,N_20512,N_20137);
and U22944 (N_22944,N_18386,N_20747);
nor U22945 (N_22945,N_19561,N_20526);
and U22946 (N_22946,N_20789,N_18647);
nor U22947 (N_22947,N_18263,N_18735);
nand U22948 (N_22948,N_18726,N_20565);
xor U22949 (N_22949,N_18082,N_20494);
nand U22950 (N_22950,N_18360,N_18004);
or U22951 (N_22951,N_19670,N_18662);
xor U22952 (N_22952,N_19012,N_20938);
and U22953 (N_22953,N_18684,N_18551);
and U22954 (N_22954,N_20846,N_19345);
nor U22955 (N_22955,N_18275,N_20736);
nor U22956 (N_22956,N_19209,N_18979);
nor U22957 (N_22957,N_18196,N_18397);
and U22958 (N_22958,N_18129,N_19355);
nor U22959 (N_22959,N_18791,N_18569);
or U22960 (N_22960,N_20570,N_20035);
nor U22961 (N_22961,N_19232,N_20443);
and U22962 (N_22962,N_19102,N_18897);
nand U22963 (N_22963,N_20616,N_18527);
nor U22964 (N_22964,N_20797,N_19360);
nand U22965 (N_22965,N_18373,N_20413);
or U22966 (N_22966,N_18021,N_18576);
xnor U22967 (N_22967,N_19983,N_20037);
or U22968 (N_22968,N_20846,N_18373);
and U22969 (N_22969,N_19511,N_19637);
nor U22970 (N_22970,N_20391,N_20277);
nor U22971 (N_22971,N_20138,N_18933);
nand U22972 (N_22972,N_18559,N_20739);
or U22973 (N_22973,N_19316,N_20206);
nor U22974 (N_22974,N_20723,N_20128);
xnor U22975 (N_22975,N_18560,N_19336);
xor U22976 (N_22976,N_19024,N_18728);
and U22977 (N_22977,N_19904,N_19896);
and U22978 (N_22978,N_19914,N_18760);
or U22979 (N_22979,N_20939,N_20819);
nor U22980 (N_22980,N_18241,N_18842);
or U22981 (N_22981,N_20165,N_19689);
xor U22982 (N_22982,N_19214,N_20422);
and U22983 (N_22983,N_19673,N_18770);
nand U22984 (N_22984,N_19314,N_20174);
and U22985 (N_22985,N_18318,N_20067);
and U22986 (N_22986,N_18079,N_20933);
nor U22987 (N_22987,N_19429,N_19745);
or U22988 (N_22988,N_19264,N_20886);
nor U22989 (N_22989,N_18351,N_18969);
nand U22990 (N_22990,N_19250,N_19590);
nand U22991 (N_22991,N_18581,N_18808);
and U22992 (N_22992,N_19268,N_18359);
and U22993 (N_22993,N_18911,N_20772);
or U22994 (N_22994,N_20542,N_20879);
nand U22995 (N_22995,N_19028,N_19149);
or U22996 (N_22996,N_18047,N_18568);
or U22997 (N_22997,N_20204,N_18760);
or U22998 (N_22998,N_20472,N_18472);
and U22999 (N_22999,N_18541,N_20639);
nor U23000 (N_23000,N_20264,N_19970);
and U23001 (N_23001,N_19038,N_18893);
nand U23002 (N_23002,N_20063,N_18687);
xor U23003 (N_23003,N_19457,N_18448);
or U23004 (N_23004,N_19729,N_20714);
xor U23005 (N_23005,N_19017,N_18288);
nand U23006 (N_23006,N_20470,N_18563);
nor U23007 (N_23007,N_19125,N_19985);
xor U23008 (N_23008,N_20747,N_20794);
nor U23009 (N_23009,N_18946,N_19299);
nor U23010 (N_23010,N_18446,N_18105);
or U23011 (N_23011,N_20021,N_19784);
nand U23012 (N_23012,N_20168,N_19784);
nor U23013 (N_23013,N_18314,N_19975);
nand U23014 (N_23014,N_18397,N_19220);
nor U23015 (N_23015,N_19795,N_20321);
and U23016 (N_23016,N_20800,N_20080);
or U23017 (N_23017,N_18221,N_18012);
nor U23018 (N_23018,N_18077,N_19715);
or U23019 (N_23019,N_20671,N_18191);
xnor U23020 (N_23020,N_20481,N_18356);
or U23021 (N_23021,N_19051,N_19501);
nor U23022 (N_23022,N_19511,N_20492);
xor U23023 (N_23023,N_20664,N_20039);
or U23024 (N_23024,N_20995,N_20527);
and U23025 (N_23025,N_19812,N_20154);
nand U23026 (N_23026,N_20048,N_18218);
nand U23027 (N_23027,N_20408,N_19455);
nand U23028 (N_23028,N_19328,N_19097);
and U23029 (N_23029,N_19245,N_18687);
xnor U23030 (N_23030,N_20481,N_18725);
xor U23031 (N_23031,N_20917,N_18309);
and U23032 (N_23032,N_18956,N_18240);
xor U23033 (N_23033,N_19485,N_18908);
nand U23034 (N_23034,N_18924,N_20140);
xor U23035 (N_23035,N_18601,N_19241);
xnor U23036 (N_23036,N_19198,N_18232);
or U23037 (N_23037,N_18838,N_19767);
or U23038 (N_23038,N_18650,N_20692);
xor U23039 (N_23039,N_20160,N_19796);
or U23040 (N_23040,N_18936,N_18494);
and U23041 (N_23041,N_19673,N_19235);
nor U23042 (N_23042,N_18772,N_20921);
nor U23043 (N_23043,N_18966,N_18916);
xnor U23044 (N_23044,N_20940,N_19268);
nand U23045 (N_23045,N_18930,N_20459);
and U23046 (N_23046,N_18570,N_19011);
nor U23047 (N_23047,N_19841,N_18767);
xnor U23048 (N_23048,N_18328,N_18337);
and U23049 (N_23049,N_19387,N_19394);
or U23050 (N_23050,N_20572,N_18003);
nor U23051 (N_23051,N_19132,N_19524);
nand U23052 (N_23052,N_19371,N_18686);
nor U23053 (N_23053,N_18634,N_19763);
nand U23054 (N_23054,N_19976,N_19169);
xnor U23055 (N_23055,N_18617,N_18983);
xnor U23056 (N_23056,N_20909,N_19135);
nor U23057 (N_23057,N_18357,N_20954);
nand U23058 (N_23058,N_19038,N_20679);
xnor U23059 (N_23059,N_19613,N_19061);
nand U23060 (N_23060,N_18206,N_20564);
and U23061 (N_23061,N_19560,N_20730);
and U23062 (N_23062,N_19106,N_18390);
or U23063 (N_23063,N_18045,N_19928);
or U23064 (N_23064,N_19659,N_18173);
nor U23065 (N_23065,N_20404,N_19759);
nor U23066 (N_23066,N_18959,N_18666);
xnor U23067 (N_23067,N_19772,N_18638);
and U23068 (N_23068,N_18065,N_20729);
nor U23069 (N_23069,N_18478,N_19347);
and U23070 (N_23070,N_20274,N_19131);
or U23071 (N_23071,N_19938,N_19263);
nor U23072 (N_23072,N_20988,N_19814);
xor U23073 (N_23073,N_20194,N_20741);
nand U23074 (N_23074,N_20766,N_19526);
and U23075 (N_23075,N_18087,N_20593);
and U23076 (N_23076,N_19320,N_18913);
xor U23077 (N_23077,N_19856,N_19601);
or U23078 (N_23078,N_19741,N_19004);
and U23079 (N_23079,N_20030,N_19577);
xnor U23080 (N_23080,N_19370,N_19578);
nor U23081 (N_23081,N_20992,N_20035);
or U23082 (N_23082,N_19323,N_18858);
and U23083 (N_23083,N_19434,N_18638);
nor U23084 (N_23084,N_20741,N_19747);
nor U23085 (N_23085,N_18652,N_19202);
nand U23086 (N_23086,N_20585,N_20616);
and U23087 (N_23087,N_20315,N_18580);
or U23088 (N_23088,N_19788,N_18218);
xor U23089 (N_23089,N_20982,N_20593);
and U23090 (N_23090,N_18591,N_20165);
xor U23091 (N_23091,N_19584,N_19733);
xor U23092 (N_23092,N_20240,N_19242);
nand U23093 (N_23093,N_19068,N_18638);
nor U23094 (N_23094,N_20404,N_18320);
nand U23095 (N_23095,N_20064,N_18791);
nor U23096 (N_23096,N_20172,N_19271);
or U23097 (N_23097,N_18581,N_18792);
or U23098 (N_23098,N_20750,N_18494);
and U23099 (N_23099,N_19890,N_20641);
and U23100 (N_23100,N_20987,N_20941);
nor U23101 (N_23101,N_20573,N_19839);
and U23102 (N_23102,N_19498,N_19557);
nand U23103 (N_23103,N_20320,N_20046);
and U23104 (N_23104,N_20939,N_19062);
or U23105 (N_23105,N_19035,N_19424);
or U23106 (N_23106,N_19260,N_18710);
and U23107 (N_23107,N_19333,N_20306);
nor U23108 (N_23108,N_20800,N_18187);
xnor U23109 (N_23109,N_18375,N_20577);
xor U23110 (N_23110,N_19973,N_19790);
nand U23111 (N_23111,N_19334,N_18364);
nor U23112 (N_23112,N_20629,N_20333);
nor U23113 (N_23113,N_20795,N_19361);
and U23114 (N_23114,N_19515,N_18601);
nand U23115 (N_23115,N_19607,N_19955);
xor U23116 (N_23116,N_20698,N_20522);
nand U23117 (N_23117,N_18327,N_18119);
nor U23118 (N_23118,N_20781,N_20323);
and U23119 (N_23119,N_18258,N_20118);
nand U23120 (N_23120,N_19450,N_20714);
or U23121 (N_23121,N_19953,N_19021);
xor U23122 (N_23122,N_19454,N_19738);
or U23123 (N_23123,N_18421,N_18031);
xor U23124 (N_23124,N_18561,N_19015);
or U23125 (N_23125,N_18810,N_19789);
xnor U23126 (N_23126,N_20749,N_20865);
or U23127 (N_23127,N_19532,N_19668);
xnor U23128 (N_23128,N_19545,N_20259);
xnor U23129 (N_23129,N_19725,N_20698);
nand U23130 (N_23130,N_19088,N_19063);
or U23131 (N_23131,N_20191,N_19013);
or U23132 (N_23132,N_19081,N_18710);
xor U23133 (N_23133,N_20367,N_18996);
xor U23134 (N_23134,N_18798,N_20776);
xnor U23135 (N_23135,N_19213,N_19298);
xor U23136 (N_23136,N_19912,N_18983);
and U23137 (N_23137,N_19689,N_18096);
nand U23138 (N_23138,N_18622,N_19310);
and U23139 (N_23139,N_20489,N_20114);
xnor U23140 (N_23140,N_18034,N_18727);
nor U23141 (N_23141,N_20090,N_18517);
or U23142 (N_23142,N_19957,N_18653);
nand U23143 (N_23143,N_19513,N_19683);
or U23144 (N_23144,N_20516,N_20582);
xor U23145 (N_23145,N_19483,N_20093);
and U23146 (N_23146,N_18415,N_19564);
and U23147 (N_23147,N_20306,N_19581);
nand U23148 (N_23148,N_19118,N_19554);
or U23149 (N_23149,N_19084,N_18302);
nor U23150 (N_23150,N_20539,N_18882);
nand U23151 (N_23151,N_19125,N_18419);
xor U23152 (N_23152,N_18375,N_19102);
nand U23153 (N_23153,N_20402,N_19940);
nand U23154 (N_23154,N_18287,N_19032);
xnor U23155 (N_23155,N_19497,N_18882);
xnor U23156 (N_23156,N_18616,N_18872);
xnor U23157 (N_23157,N_20323,N_20891);
and U23158 (N_23158,N_20351,N_18496);
nand U23159 (N_23159,N_18623,N_19676);
xor U23160 (N_23160,N_19132,N_19398);
nor U23161 (N_23161,N_19924,N_18676);
and U23162 (N_23162,N_19202,N_18685);
or U23163 (N_23163,N_20920,N_20882);
nand U23164 (N_23164,N_20457,N_19353);
xor U23165 (N_23165,N_19121,N_19976);
xor U23166 (N_23166,N_19350,N_18577);
and U23167 (N_23167,N_20068,N_18304);
xor U23168 (N_23168,N_18747,N_18015);
or U23169 (N_23169,N_20365,N_20651);
xor U23170 (N_23170,N_20262,N_19578);
xor U23171 (N_23171,N_19454,N_20193);
nand U23172 (N_23172,N_18318,N_19742);
nand U23173 (N_23173,N_18218,N_20848);
or U23174 (N_23174,N_19108,N_19295);
nor U23175 (N_23175,N_19421,N_20654);
xnor U23176 (N_23176,N_18560,N_20823);
xnor U23177 (N_23177,N_20630,N_20571);
nand U23178 (N_23178,N_19931,N_19445);
nor U23179 (N_23179,N_20598,N_20486);
and U23180 (N_23180,N_18059,N_18430);
nand U23181 (N_23181,N_19019,N_18373);
nor U23182 (N_23182,N_19903,N_18160);
nand U23183 (N_23183,N_19107,N_20998);
and U23184 (N_23184,N_18554,N_18641);
nand U23185 (N_23185,N_18384,N_19641);
and U23186 (N_23186,N_19437,N_18390);
and U23187 (N_23187,N_20141,N_20340);
nor U23188 (N_23188,N_20160,N_18347);
xor U23189 (N_23189,N_19109,N_19952);
nand U23190 (N_23190,N_18306,N_18491);
xnor U23191 (N_23191,N_19810,N_20002);
nand U23192 (N_23192,N_20838,N_19229);
or U23193 (N_23193,N_19105,N_19319);
and U23194 (N_23194,N_20973,N_19418);
or U23195 (N_23195,N_19710,N_18079);
nor U23196 (N_23196,N_18279,N_19215);
xnor U23197 (N_23197,N_19829,N_18514);
xor U23198 (N_23198,N_18934,N_20889);
nand U23199 (N_23199,N_18894,N_19622);
nor U23200 (N_23200,N_19166,N_18433);
and U23201 (N_23201,N_18822,N_19324);
nand U23202 (N_23202,N_20304,N_19930);
or U23203 (N_23203,N_18809,N_18822);
nand U23204 (N_23204,N_19582,N_19414);
xor U23205 (N_23205,N_18934,N_19918);
xnor U23206 (N_23206,N_19904,N_20555);
nand U23207 (N_23207,N_19717,N_18899);
xnor U23208 (N_23208,N_18504,N_20443);
nor U23209 (N_23209,N_18331,N_20706);
and U23210 (N_23210,N_20296,N_19763);
or U23211 (N_23211,N_18766,N_18936);
and U23212 (N_23212,N_19656,N_20509);
xor U23213 (N_23213,N_19254,N_19918);
nor U23214 (N_23214,N_20723,N_18886);
nand U23215 (N_23215,N_18815,N_20670);
or U23216 (N_23216,N_19905,N_20430);
and U23217 (N_23217,N_18919,N_18108);
or U23218 (N_23218,N_19104,N_19948);
xnor U23219 (N_23219,N_19044,N_19824);
and U23220 (N_23220,N_18199,N_18926);
nor U23221 (N_23221,N_20754,N_19044);
and U23222 (N_23222,N_20936,N_18280);
xor U23223 (N_23223,N_20731,N_18136);
nand U23224 (N_23224,N_18257,N_18324);
and U23225 (N_23225,N_18174,N_19355);
nor U23226 (N_23226,N_20354,N_19361);
nand U23227 (N_23227,N_20619,N_20006);
and U23228 (N_23228,N_20097,N_18869);
nand U23229 (N_23229,N_20845,N_20685);
nand U23230 (N_23230,N_18937,N_18780);
and U23231 (N_23231,N_19727,N_19921);
or U23232 (N_23232,N_19523,N_18462);
nor U23233 (N_23233,N_18232,N_18497);
xnor U23234 (N_23234,N_19505,N_20747);
nand U23235 (N_23235,N_20172,N_18757);
and U23236 (N_23236,N_19254,N_20518);
nor U23237 (N_23237,N_19731,N_19237);
nand U23238 (N_23238,N_19228,N_20067);
nor U23239 (N_23239,N_20150,N_19327);
xnor U23240 (N_23240,N_18320,N_18096);
or U23241 (N_23241,N_19523,N_20923);
xor U23242 (N_23242,N_18645,N_18990);
nor U23243 (N_23243,N_18623,N_20170);
xor U23244 (N_23244,N_18419,N_19635);
or U23245 (N_23245,N_20493,N_18335);
nand U23246 (N_23246,N_19112,N_20786);
or U23247 (N_23247,N_20365,N_20920);
and U23248 (N_23248,N_20635,N_19741);
nand U23249 (N_23249,N_18166,N_20561);
nor U23250 (N_23250,N_20170,N_19630);
and U23251 (N_23251,N_19909,N_18761);
nand U23252 (N_23252,N_18129,N_19834);
or U23253 (N_23253,N_20981,N_19025);
nand U23254 (N_23254,N_20423,N_20620);
nand U23255 (N_23255,N_20698,N_19589);
nand U23256 (N_23256,N_18329,N_20850);
and U23257 (N_23257,N_18830,N_18541);
xor U23258 (N_23258,N_20079,N_19217);
nand U23259 (N_23259,N_18604,N_18737);
xor U23260 (N_23260,N_18943,N_18944);
nand U23261 (N_23261,N_20402,N_19228);
and U23262 (N_23262,N_18043,N_18581);
or U23263 (N_23263,N_20589,N_18613);
xnor U23264 (N_23264,N_19170,N_18975);
and U23265 (N_23265,N_19553,N_20181);
and U23266 (N_23266,N_18648,N_20200);
xnor U23267 (N_23267,N_20559,N_19387);
and U23268 (N_23268,N_19751,N_20475);
nand U23269 (N_23269,N_18151,N_20860);
nand U23270 (N_23270,N_20384,N_20507);
nor U23271 (N_23271,N_19823,N_18206);
or U23272 (N_23272,N_20205,N_19660);
xor U23273 (N_23273,N_18150,N_18218);
or U23274 (N_23274,N_20463,N_19141);
or U23275 (N_23275,N_19608,N_18000);
nor U23276 (N_23276,N_19611,N_20232);
and U23277 (N_23277,N_19957,N_18761);
nor U23278 (N_23278,N_19258,N_18871);
or U23279 (N_23279,N_19230,N_18355);
xnor U23280 (N_23280,N_20322,N_18181);
or U23281 (N_23281,N_19970,N_19748);
nand U23282 (N_23282,N_18203,N_20668);
nor U23283 (N_23283,N_19189,N_19492);
nand U23284 (N_23284,N_18841,N_19208);
nand U23285 (N_23285,N_19505,N_20404);
and U23286 (N_23286,N_20776,N_20095);
nor U23287 (N_23287,N_20497,N_20710);
nor U23288 (N_23288,N_19145,N_18049);
nand U23289 (N_23289,N_20089,N_20228);
or U23290 (N_23290,N_18190,N_19432);
nand U23291 (N_23291,N_18445,N_19932);
nor U23292 (N_23292,N_20453,N_19258);
or U23293 (N_23293,N_20757,N_20993);
xnor U23294 (N_23294,N_20439,N_20842);
or U23295 (N_23295,N_20742,N_19469);
nor U23296 (N_23296,N_18942,N_18425);
or U23297 (N_23297,N_20045,N_18090);
nand U23298 (N_23298,N_19627,N_18002);
and U23299 (N_23299,N_19817,N_18380);
nor U23300 (N_23300,N_20452,N_19383);
nor U23301 (N_23301,N_19432,N_20773);
nand U23302 (N_23302,N_19708,N_19436);
nor U23303 (N_23303,N_20431,N_20583);
nand U23304 (N_23304,N_20077,N_19524);
nor U23305 (N_23305,N_18577,N_19636);
xnor U23306 (N_23306,N_18934,N_19001);
or U23307 (N_23307,N_18472,N_18971);
and U23308 (N_23308,N_18404,N_19458);
and U23309 (N_23309,N_19479,N_18138);
or U23310 (N_23310,N_18628,N_20405);
or U23311 (N_23311,N_20678,N_18467);
nand U23312 (N_23312,N_18538,N_20619);
nand U23313 (N_23313,N_18966,N_19918);
and U23314 (N_23314,N_18742,N_20362);
or U23315 (N_23315,N_19738,N_19665);
xnor U23316 (N_23316,N_20624,N_19300);
xor U23317 (N_23317,N_18529,N_19973);
nor U23318 (N_23318,N_19257,N_19771);
nor U23319 (N_23319,N_20324,N_18268);
and U23320 (N_23320,N_20764,N_20394);
xnor U23321 (N_23321,N_20369,N_19862);
or U23322 (N_23322,N_20453,N_18260);
nand U23323 (N_23323,N_19168,N_20865);
or U23324 (N_23324,N_19893,N_20489);
or U23325 (N_23325,N_19213,N_20779);
nor U23326 (N_23326,N_20650,N_19217);
and U23327 (N_23327,N_19879,N_20572);
nor U23328 (N_23328,N_19078,N_19013);
nor U23329 (N_23329,N_18762,N_19278);
and U23330 (N_23330,N_20126,N_18734);
nand U23331 (N_23331,N_19885,N_19339);
nand U23332 (N_23332,N_20672,N_20933);
xor U23333 (N_23333,N_18769,N_18670);
nand U23334 (N_23334,N_20693,N_20120);
and U23335 (N_23335,N_18049,N_20677);
nand U23336 (N_23336,N_18384,N_20231);
nor U23337 (N_23337,N_19672,N_20610);
and U23338 (N_23338,N_19981,N_18128);
nor U23339 (N_23339,N_18684,N_20369);
nand U23340 (N_23340,N_20097,N_18866);
and U23341 (N_23341,N_18946,N_18789);
nand U23342 (N_23342,N_19811,N_20473);
nor U23343 (N_23343,N_20070,N_18030);
nor U23344 (N_23344,N_19701,N_18028);
xnor U23345 (N_23345,N_18550,N_19569);
xnor U23346 (N_23346,N_20813,N_19721);
or U23347 (N_23347,N_20232,N_18306);
nor U23348 (N_23348,N_19948,N_19307);
or U23349 (N_23349,N_20400,N_18276);
or U23350 (N_23350,N_20282,N_19663);
nor U23351 (N_23351,N_19319,N_19096);
nand U23352 (N_23352,N_20594,N_19429);
nor U23353 (N_23353,N_18480,N_18528);
nand U23354 (N_23354,N_19097,N_20961);
and U23355 (N_23355,N_20273,N_18899);
nor U23356 (N_23356,N_19094,N_19371);
xnor U23357 (N_23357,N_19437,N_18567);
nand U23358 (N_23358,N_19554,N_19083);
xor U23359 (N_23359,N_18208,N_20678);
nor U23360 (N_23360,N_19008,N_19780);
and U23361 (N_23361,N_20312,N_19546);
nor U23362 (N_23362,N_18898,N_20592);
and U23363 (N_23363,N_20601,N_20487);
xnor U23364 (N_23364,N_20101,N_18336);
or U23365 (N_23365,N_18953,N_20240);
nand U23366 (N_23366,N_18384,N_19454);
and U23367 (N_23367,N_18226,N_19247);
nor U23368 (N_23368,N_19824,N_18103);
nor U23369 (N_23369,N_18563,N_18279);
or U23370 (N_23370,N_18566,N_18989);
nor U23371 (N_23371,N_18109,N_20548);
nand U23372 (N_23372,N_20587,N_18148);
nor U23373 (N_23373,N_18109,N_19382);
xnor U23374 (N_23374,N_18119,N_18636);
xor U23375 (N_23375,N_19215,N_19078);
or U23376 (N_23376,N_20351,N_20741);
or U23377 (N_23377,N_20930,N_20598);
nand U23378 (N_23378,N_19151,N_19928);
and U23379 (N_23379,N_20233,N_18448);
nor U23380 (N_23380,N_20718,N_19957);
nor U23381 (N_23381,N_19721,N_18812);
nor U23382 (N_23382,N_18856,N_18447);
or U23383 (N_23383,N_19691,N_18068);
nand U23384 (N_23384,N_20106,N_19154);
nand U23385 (N_23385,N_18666,N_19490);
nor U23386 (N_23386,N_19571,N_19677);
nor U23387 (N_23387,N_19075,N_19403);
and U23388 (N_23388,N_20199,N_20248);
xnor U23389 (N_23389,N_18743,N_18095);
and U23390 (N_23390,N_18194,N_18698);
nor U23391 (N_23391,N_18346,N_20283);
and U23392 (N_23392,N_19629,N_18345);
and U23393 (N_23393,N_20490,N_20469);
nor U23394 (N_23394,N_19712,N_18676);
or U23395 (N_23395,N_19363,N_20900);
xor U23396 (N_23396,N_18295,N_20995);
xor U23397 (N_23397,N_19992,N_18529);
or U23398 (N_23398,N_19054,N_18972);
nor U23399 (N_23399,N_20937,N_18299);
nand U23400 (N_23400,N_20391,N_20175);
nor U23401 (N_23401,N_19616,N_18202);
xor U23402 (N_23402,N_20311,N_18644);
and U23403 (N_23403,N_18621,N_18292);
xor U23404 (N_23404,N_20947,N_20717);
nand U23405 (N_23405,N_18167,N_18473);
or U23406 (N_23406,N_19338,N_19327);
xnor U23407 (N_23407,N_18533,N_20465);
xor U23408 (N_23408,N_20268,N_18991);
and U23409 (N_23409,N_20738,N_18432);
nor U23410 (N_23410,N_18059,N_19409);
nand U23411 (N_23411,N_18858,N_18022);
xnor U23412 (N_23412,N_19378,N_19097);
nand U23413 (N_23413,N_18424,N_18964);
or U23414 (N_23414,N_20944,N_19578);
xor U23415 (N_23415,N_18415,N_19138);
or U23416 (N_23416,N_20802,N_20306);
xor U23417 (N_23417,N_20529,N_20430);
xor U23418 (N_23418,N_20857,N_19919);
or U23419 (N_23419,N_18772,N_18939);
nand U23420 (N_23420,N_20491,N_19302);
nor U23421 (N_23421,N_20350,N_19828);
and U23422 (N_23422,N_19476,N_19396);
or U23423 (N_23423,N_20089,N_19151);
xnor U23424 (N_23424,N_18954,N_19439);
nor U23425 (N_23425,N_19334,N_19397);
xnor U23426 (N_23426,N_20016,N_19009);
and U23427 (N_23427,N_19621,N_18194);
or U23428 (N_23428,N_18526,N_20604);
and U23429 (N_23429,N_20450,N_18433);
nand U23430 (N_23430,N_20475,N_18713);
or U23431 (N_23431,N_19825,N_18073);
xor U23432 (N_23432,N_18624,N_19782);
nand U23433 (N_23433,N_19421,N_20586);
and U23434 (N_23434,N_19123,N_19259);
nor U23435 (N_23435,N_20267,N_18620);
and U23436 (N_23436,N_18494,N_20059);
nand U23437 (N_23437,N_20433,N_18215);
nand U23438 (N_23438,N_20796,N_20811);
nand U23439 (N_23439,N_18295,N_19361);
and U23440 (N_23440,N_20729,N_20659);
or U23441 (N_23441,N_19301,N_18955);
nor U23442 (N_23442,N_19728,N_19013);
or U23443 (N_23443,N_18538,N_18257);
xnor U23444 (N_23444,N_20395,N_20957);
and U23445 (N_23445,N_20226,N_19675);
xnor U23446 (N_23446,N_19978,N_18956);
nor U23447 (N_23447,N_20325,N_19926);
nor U23448 (N_23448,N_19196,N_18010);
nor U23449 (N_23449,N_18680,N_18218);
nor U23450 (N_23450,N_20678,N_20802);
or U23451 (N_23451,N_20729,N_19403);
nand U23452 (N_23452,N_19960,N_18613);
or U23453 (N_23453,N_19531,N_20155);
and U23454 (N_23454,N_20959,N_20698);
or U23455 (N_23455,N_19251,N_20116);
and U23456 (N_23456,N_20860,N_18507);
nor U23457 (N_23457,N_20461,N_20404);
xor U23458 (N_23458,N_19806,N_18362);
nand U23459 (N_23459,N_18646,N_20561);
nand U23460 (N_23460,N_20644,N_19339);
xnor U23461 (N_23461,N_19732,N_20587);
and U23462 (N_23462,N_20290,N_19305);
and U23463 (N_23463,N_20729,N_19577);
and U23464 (N_23464,N_20339,N_18219);
nor U23465 (N_23465,N_18941,N_19764);
and U23466 (N_23466,N_18453,N_19940);
xnor U23467 (N_23467,N_20455,N_18579);
nor U23468 (N_23468,N_19916,N_20290);
nand U23469 (N_23469,N_18948,N_18773);
xnor U23470 (N_23470,N_19565,N_19864);
and U23471 (N_23471,N_19598,N_20763);
nand U23472 (N_23472,N_19930,N_18979);
nor U23473 (N_23473,N_20012,N_18256);
or U23474 (N_23474,N_20960,N_19378);
nor U23475 (N_23475,N_18851,N_18781);
xnor U23476 (N_23476,N_18685,N_19880);
and U23477 (N_23477,N_20431,N_19491);
xor U23478 (N_23478,N_20490,N_20392);
or U23479 (N_23479,N_20171,N_19724);
xnor U23480 (N_23480,N_19711,N_19069);
and U23481 (N_23481,N_19936,N_20630);
nor U23482 (N_23482,N_19062,N_20066);
nand U23483 (N_23483,N_19116,N_19882);
nand U23484 (N_23484,N_20068,N_18871);
nor U23485 (N_23485,N_20593,N_20985);
nand U23486 (N_23486,N_19354,N_20720);
nor U23487 (N_23487,N_20410,N_18517);
xor U23488 (N_23488,N_20140,N_19745);
and U23489 (N_23489,N_18247,N_18647);
xor U23490 (N_23490,N_20254,N_19597);
nor U23491 (N_23491,N_20885,N_20417);
and U23492 (N_23492,N_18831,N_19600);
nor U23493 (N_23493,N_20409,N_18309);
and U23494 (N_23494,N_20341,N_18728);
and U23495 (N_23495,N_18039,N_18063);
and U23496 (N_23496,N_20742,N_19483);
and U23497 (N_23497,N_18620,N_20995);
and U23498 (N_23498,N_19224,N_18851);
nand U23499 (N_23499,N_20073,N_20579);
and U23500 (N_23500,N_20145,N_19345);
or U23501 (N_23501,N_19865,N_18490);
xor U23502 (N_23502,N_20351,N_18943);
nand U23503 (N_23503,N_20002,N_19918);
nand U23504 (N_23504,N_20925,N_18954);
or U23505 (N_23505,N_19708,N_18964);
nor U23506 (N_23506,N_19707,N_18796);
nand U23507 (N_23507,N_19880,N_20601);
nand U23508 (N_23508,N_20565,N_20489);
xnor U23509 (N_23509,N_19140,N_19882);
or U23510 (N_23510,N_19880,N_19963);
xnor U23511 (N_23511,N_19216,N_20846);
or U23512 (N_23512,N_20813,N_20772);
nand U23513 (N_23513,N_19325,N_19451);
xnor U23514 (N_23514,N_19833,N_20220);
and U23515 (N_23515,N_19370,N_18076);
or U23516 (N_23516,N_18803,N_19330);
or U23517 (N_23517,N_18623,N_19837);
or U23518 (N_23518,N_19954,N_20597);
xnor U23519 (N_23519,N_19755,N_18182);
xnor U23520 (N_23520,N_18353,N_18036);
or U23521 (N_23521,N_19461,N_18378);
or U23522 (N_23522,N_20432,N_19992);
and U23523 (N_23523,N_19569,N_20809);
nor U23524 (N_23524,N_19067,N_18734);
nand U23525 (N_23525,N_18426,N_19613);
nor U23526 (N_23526,N_20541,N_20871);
nand U23527 (N_23527,N_18591,N_19444);
nand U23528 (N_23528,N_18420,N_18054);
nand U23529 (N_23529,N_20316,N_19030);
nor U23530 (N_23530,N_20563,N_18207);
xor U23531 (N_23531,N_20714,N_20320);
or U23532 (N_23532,N_18534,N_18707);
nor U23533 (N_23533,N_19308,N_19509);
nand U23534 (N_23534,N_18628,N_19512);
and U23535 (N_23535,N_18903,N_18447);
and U23536 (N_23536,N_18388,N_18600);
nor U23537 (N_23537,N_19722,N_18011);
nor U23538 (N_23538,N_19210,N_20204);
xnor U23539 (N_23539,N_19036,N_20413);
or U23540 (N_23540,N_19190,N_19073);
and U23541 (N_23541,N_19411,N_18607);
xnor U23542 (N_23542,N_20955,N_20078);
or U23543 (N_23543,N_19766,N_18827);
nand U23544 (N_23544,N_19574,N_20825);
and U23545 (N_23545,N_18642,N_20387);
or U23546 (N_23546,N_19033,N_18594);
and U23547 (N_23547,N_20730,N_19215);
nand U23548 (N_23548,N_19789,N_18408);
xor U23549 (N_23549,N_19402,N_18415);
nand U23550 (N_23550,N_20646,N_19007);
and U23551 (N_23551,N_18903,N_20838);
xnor U23552 (N_23552,N_18986,N_18450);
xor U23553 (N_23553,N_20726,N_19906);
xor U23554 (N_23554,N_20241,N_20570);
and U23555 (N_23555,N_18387,N_18053);
xnor U23556 (N_23556,N_20678,N_18406);
or U23557 (N_23557,N_20642,N_18382);
and U23558 (N_23558,N_18839,N_19576);
and U23559 (N_23559,N_20839,N_18408);
and U23560 (N_23560,N_18054,N_18632);
or U23561 (N_23561,N_19254,N_19037);
xnor U23562 (N_23562,N_19947,N_18525);
or U23563 (N_23563,N_19978,N_18044);
nor U23564 (N_23564,N_20005,N_20342);
nand U23565 (N_23565,N_19757,N_20698);
nand U23566 (N_23566,N_19641,N_19666);
nor U23567 (N_23567,N_18812,N_20290);
nand U23568 (N_23568,N_19899,N_20857);
and U23569 (N_23569,N_19967,N_20840);
and U23570 (N_23570,N_20504,N_19013);
and U23571 (N_23571,N_19872,N_19323);
or U23572 (N_23572,N_20600,N_18455);
xor U23573 (N_23573,N_20611,N_19328);
nand U23574 (N_23574,N_20324,N_18451);
nand U23575 (N_23575,N_18994,N_19968);
xnor U23576 (N_23576,N_20685,N_18155);
or U23577 (N_23577,N_20531,N_20737);
xor U23578 (N_23578,N_20875,N_20882);
nand U23579 (N_23579,N_20010,N_18299);
nand U23580 (N_23580,N_18058,N_20825);
xor U23581 (N_23581,N_19123,N_20104);
or U23582 (N_23582,N_18518,N_20376);
nor U23583 (N_23583,N_19330,N_18343);
nor U23584 (N_23584,N_20356,N_18686);
xor U23585 (N_23585,N_19396,N_19985);
nor U23586 (N_23586,N_20941,N_19484);
nand U23587 (N_23587,N_19440,N_18928);
and U23588 (N_23588,N_18699,N_18068);
nor U23589 (N_23589,N_18233,N_19166);
nand U23590 (N_23590,N_20402,N_18494);
and U23591 (N_23591,N_19537,N_20885);
nand U23592 (N_23592,N_18515,N_20851);
or U23593 (N_23593,N_18278,N_19732);
nor U23594 (N_23594,N_20004,N_19182);
and U23595 (N_23595,N_19706,N_20344);
nor U23596 (N_23596,N_18049,N_20399);
xor U23597 (N_23597,N_19622,N_18722);
nor U23598 (N_23598,N_20036,N_19235);
xor U23599 (N_23599,N_18178,N_20363);
nand U23600 (N_23600,N_20972,N_18500);
xor U23601 (N_23601,N_20202,N_19736);
and U23602 (N_23602,N_20017,N_18655);
nor U23603 (N_23603,N_19726,N_18220);
nand U23604 (N_23604,N_19370,N_18088);
nand U23605 (N_23605,N_20223,N_18379);
nor U23606 (N_23606,N_20297,N_19699);
nand U23607 (N_23607,N_18679,N_20997);
nor U23608 (N_23608,N_20427,N_20396);
nand U23609 (N_23609,N_18101,N_19073);
xnor U23610 (N_23610,N_19422,N_18226);
or U23611 (N_23611,N_20419,N_18365);
nand U23612 (N_23612,N_19565,N_19589);
nand U23613 (N_23613,N_19177,N_20609);
nor U23614 (N_23614,N_18019,N_19786);
or U23615 (N_23615,N_18894,N_20503);
and U23616 (N_23616,N_18493,N_18484);
or U23617 (N_23617,N_19668,N_18288);
nand U23618 (N_23618,N_20544,N_20164);
nor U23619 (N_23619,N_18948,N_20814);
and U23620 (N_23620,N_18313,N_19397);
xnor U23621 (N_23621,N_19550,N_18917);
xor U23622 (N_23622,N_20051,N_18368);
nand U23623 (N_23623,N_18045,N_20997);
and U23624 (N_23624,N_20467,N_20882);
xnor U23625 (N_23625,N_19383,N_19444);
xnor U23626 (N_23626,N_18815,N_20258);
xor U23627 (N_23627,N_18083,N_20713);
xor U23628 (N_23628,N_18747,N_20820);
nand U23629 (N_23629,N_19495,N_20119);
and U23630 (N_23630,N_20420,N_18467);
xnor U23631 (N_23631,N_18102,N_18381);
xor U23632 (N_23632,N_20888,N_18923);
nor U23633 (N_23633,N_20989,N_20428);
or U23634 (N_23634,N_18032,N_19620);
nand U23635 (N_23635,N_19172,N_20896);
or U23636 (N_23636,N_20229,N_20998);
or U23637 (N_23637,N_20203,N_18980);
xor U23638 (N_23638,N_19331,N_20986);
or U23639 (N_23639,N_19294,N_18824);
xor U23640 (N_23640,N_19666,N_18760);
nor U23641 (N_23641,N_19523,N_18922);
or U23642 (N_23642,N_20088,N_20291);
nor U23643 (N_23643,N_18256,N_18938);
nand U23644 (N_23644,N_20412,N_20972);
or U23645 (N_23645,N_18153,N_18811);
or U23646 (N_23646,N_18343,N_20635);
nor U23647 (N_23647,N_19559,N_19394);
nand U23648 (N_23648,N_20685,N_20887);
and U23649 (N_23649,N_19787,N_20637);
or U23650 (N_23650,N_20980,N_19858);
nor U23651 (N_23651,N_19372,N_18715);
nand U23652 (N_23652,N_18112,N_20882);
or U23653 (N_23653,N_19423,N_20218);
nor U23654 (N_23654,N_19969,N_18221);
nor U23655 (N_23655,N_18960,N_18505);
and U23656 (N_23656,N_19037,N_18539);
xnor U23657 (N_23657,N_20964,N_18843);
nand U23658 (N_23658,N_20323,N_19767);
nand U23659 (N_23659,N_18206,N_18010);
nor U23660 (N_23660,N_19677,N_18196);
and U23661 (N_23661,N_18279,N_19191);
nor U23662 (N_23662,N_18625,N_18356);
and U23663 (N_23663,N_19348,N_18375);
nand U23664 (N_23664,N_19980,N_18354);
and U23665 (N_23665,N_19797,N_18538);
nand U23666 (N_23666,N_18051,N_20915);
nand U23667 (N_23667,N_18264,N_20839);
or U23668 (N_23668,N_20165,N_20895);
nand U23669 (N_23669,N_20848,N_18978);
and U23670 (N_23670,N_20914,N_20751);
nor U23671 (N_23671,N_18009,N_20179);
nor U23672 (N_23672,N_19656,N_19354);
xnor U23673 (N_23673,N_18290,N_20702);
nand U23674 (N_23674,N_18265,N_20590);
and U23675 (N_23675,N_20552,N_19273);
and U23676 (N_23676,N_19253,N_19901);
or U23677 (N_23677,N_19654,N_19559);
xor U23678 (N_23678,N_20111,N_18584);
nand U23679 (N_23679,N_18169,N_19112);
or U23680 (N_23680,N_19447,N_18479);
xnor U23681 (N_23681,N_20753,N_20878);
xnor U23682 (N_23682,N_18482,N_19356);
nor U23683 (N_23683,N_20556,N_18668);
xor U23684 (N_23684,N_20745,N_19258);
nand U23685 (N_23685,N_19952,N_18563);
and U23686 (N_23686,N_20651,N_18242);
nand U23687 (N_23687,N_19072,N_18192);
and U23688 (N_23688,N_19174,N_19367);
nor U23689 (N_23689,N_18409,N_19032);
nor U23690 (N_23690,N_20109,N_20709);
xnor U23691 (N_23691,N_19075,N_20124);
nor U23692 (N_23692,N_19848,N_18387);
and U23693 (N_23693,N_19689,N_18978);
or U23694 (N_23694,N_18539,N_20031);
and U23695 (N_23695,N_18526,N_20569);
nor U23696 (N_23696,N_20602,N_18417);
xnor U23697 (N_23697,N_20709,N_19265);
or U23698 (N_23698,N_18583,N_19533);
or U23699 (N_23699,N_18389,N_19733);
nand U23700 (N_23700,N_18351,N_20584);
nor U23701 (N_23701,N_19225,N_20109);
nor U23702 (N_23702,N_20286,N_18759);
and U23703 (N_23703,N_20525,N_20625);
nor U23704 (N_23704,N_19336,N_19073);
or U23705 (N_23705,N_18255,N_20809);
or U23706 (N_23706,N_20314,N_20052);
and U23707 (N_23707,N_19366,N_20335);
or U23708 (N_23708,N_20526,N_19366);
nand U23709 (N_23709,N_20579,N_19001);
xor U23710 (N_23710,N_19085,N_20862);
or U23711 (N_23711,N_20424,N_18820);
nor U23712 (N_23712,N_18225,N_20430);
nor U23713 (N_23713,N_19992,N_18731);
or U23714 (N_23714,N_19987,N_18218);
nor U23715 (N_23715,N_19052,N_18451);
xor U23716 (N_23716,N_20719,N_19384);
nand U23717 (N_23717,N_19884,N_19454);
nand U23718 (N_23718,N_19621,N_18528);
and U23719 (N_23719,N_19429,N_20631);
or U23720 (N_23720,N_18006,N_20783);
or U23721 (N_23721,N_19829,N_19071);
nand U23722 (N_23722,N_20012,N_19681);
or U23723 (N_23723,N_20921,N_18122);
nand U23724 (N_23724,N_18785,N_18213);
nor U23725 (N_23725,N_19875,N_18914);
xnor U23726 (N_23726,N_19554,N_19393);
nor U23727 (N_23727,N_19068,N_18797);
or U23728 (N_23728,N_18082,N_20383);
nor U23729 (N_23729,N_20721,N_20334);
and U23730 (N_23730,N_18708,N_19178);
or U23731 (N_23731,N_20645,N_20230);
nand U23732 (N_23732,N_19569,N_19263);
and U23733 (N_23733,N_20597,N_18009);
nand U23734 (N_23734,N_18349,N_20944);
and U23735 (N_23735,N_18850,N_19032);
and U23736 (N_23736,N_20302,N_20363);
nor U23737 (N_23737,N_20257,N_18313);
or U23738 (N_23738,N_19995,N_18600);
xor U23739 (N_23739,N_20445,N_18944);
xor U23740 (N_23740,N_18130,N_19183);
nand U23741 (N_23741,N_20849,N_18628);
and U23742 (N_23742,N_20493,N_18372);
xor U23743 (N_23743,N_20802,N_18393);
xor U23744 (N_23744,N_18759,N_20112);
or U23745 (N_23745,N_19799,N_20045);
nand U23746 (N_23746,N_20866,N_19161);
xnor U23747 (N_23747,N_20269,N_19552);
xor U23748 (N_23748,N_20406,N_18685);
nand U23749 (N_23749,N_20497,N_20605);
nor U23750 (N_23750,N_18559,N_19472);
or U23751 (N_23751,N_18175,N_19881);
or U23752 (N_23752,N_20968,N_18278);
nor U23753 (N_23753,N_20097,N_19280);
or U23754 (N_23754,N_20830,N_20505);
and U23755 (N_23755,N_19212,N_18241);
nand U23756 (N_23756,N_19915,N_19725);
nor U23757 (N_23757,N_20258,N_18308);
xnor U23758 (N_23758,N_20285,N_20034);
xor U23759 (N_23759,N_20103,N_19801);
nor U23760 (N_23760,N_18780,N_20341);
nand U23761 (N_23761,N_20612,N_19290);
and U23762 (N_23762,N_18989,N_20645);
xor U23763 (N_23763,N_19523,N_18652);
and U23764 (N_23764,N_20441,N_20274);
nand U23765 (N_23765,N_18584,N_19480);
nand U23766 (N_23766,N_20793,N_20405);
or U23767 (N_23767,N_19528,N_19343);
and U23768 (N_23768,N_18515,N_19197);
or U23769 (N_23769,N_20644,N_18572);
nor U23770 (N_23770,N_18023,N_20480);
xnor U23771 (N_23771,N_18501,N_20364);
or U23772 (N_23772,N_18049,N_20854);
xor U23773 (N_23773,N_20242,N_18727);
nor U23774 (N_23774,N_20441,N_18758);
nor U23775 (N_23775,N_18990,N_20014);
and U23776 (N_23776,N_19781,N_19554);
nand U23777 (N_23777,N_18006,N_18066);
or U23778 (N_23778,N_20382,N_19356);
or U23779 (N_23779,N_18493,N_20876);
and U23780 (N_23780,N_19037,N_20157);
and U23781 (N_23781,N_19791,N_20641);
nand U23782 (N_23782,N_18753,N_20996);
xnor U23783 (N_23783,N_18560,N_19787);
or U23784 (N_23784,N_18170,N_18526);
xor U23785 (N_23785,N_19161,N_18109);
and U23786 (N_23786,N_18860,N_19585);
nand U23787 (N_23787,N_19754,N_20317);
nand U23788 (N_23788,N_19089,N_18641);
nor U23789 (N_23789,N_19027,N_20887);
and U23790 (N_23790,N_18375,N_18972);
and U23791 (N_23791,N_19642,N_18298);
and U23792 (N_23792,N_20301,N_19782);
nand U23793 (N_23793,N_20943,N_20808);
nand U23794 (N_23794,N_18642,N_20186);
nand U23795 (N_23795,N_20689,N_18556);
nand U23796 (N_23796,N_19999,N_20768);
nor U23797 (N_23797,N_19079,N_20827);
nor U23798 (N_23798,N_18268,N_18704);
nor U23799 (N_23799,N_20234,N_19384);
or U23800 (N_23800,N_19615,N_18584);
and U23801 (N_23801,N_18085,N_20340);
or U23802 (N_23802,N_20149,N_20036);
nand U23803 (N_23803,N_18590,N_18940);
nand U23804 (N_23804,N_19236,N_20535);
and U23805 (N_23805,N_19606,N_18431);
and U23806 (N_23806,N_20364,N_20939);
xor U23807 (N_23807,N_19028,N_18294);
nand U23808 (N_23808,N_19642,N_18314);
or U23809 (N_23809,N_19308,N_19420);
nor U23810 (N_23810,N_18209,N_20342);
xnor U23811 (N_23811,N_20633,N_20249);
nor U23812 (N_23812,N_20448,N_20860);
nor U23813 (N_23813,N_18844,N_20088);
nor U23814 (N_23814,N_19984,N_19881);
xor U23815 (N_23815,N_19683,N_19936);
and U23816 (N_23816,N_18831,N_19669);
and U23817 (N_23817,N_19445,N_18731);
xnor U23818 (N_23818,N_19377,N_18890);
xor U23819 (N_23819,N_20932,N_20715);
xor U23820 (N_23820,N_19422,N_20221);
nor U23821 (N_23821,N_20611,N_18327);
xnor U23822 (N_23822,N_19417,N_20484);
or U23823 (N_23823,N_20541,N_19893);
nand U23824 (N_23824,N_18748,N_19426);
and U23825 (N_23825,N_20944,N_18179);
xnor U23826 (N_23826,N_19371,N_19722);
or U23827 (N_23827,N_19371,N_18328);
nor U23828 (N_23828,N_18606,N_18621);
nor U23829 (N_23829,N_19695,N_19714);
and U23830 (N_23830,N_18726,N_18414);
or U23831 (N_23831,N_19096,N_19766);
nand U23832 (N_23832,N_19851,N_19871);
xor U23833 (N_23833,N_18352,N_19387);
nor U23834 (N_23834,N_20633,N_20737);
or U23835 (N_23835,N_19575,N_20295);
xor U23836 (N_23836,N_19151,N_20917);
or U23837 (N_23837,N_19825,N_20562);
nor U23838 (N_23838,N_19424,N_20109);
or U23839 (N_23839,N_20186,N_18444);
xnor U23840 (N_23840,N_18730,N_20101);
and U23841 (N_23841,N_20335,N_19594);
or U23842 (N_23842,N_20895,N_20864);
or U23843 (N_23843,N_19153,N_19218);
nor U23844 (N_23844,N_19016,N_18531);
xor U23845 (N_23845,N_18574,N_19327);
xor U23846 (N_23846,N_19664,N_20161);
and U23847 (N_23847,N_18357,N_18575);
or U23848 (N_23848,N_18053,N_20638);
nand U23849 (N_23849,N_20289,N_19472);
nor U23850 (N_23850,N_18419,N_20059);
or U23851 (N_23851,N_20526,N_18520);
nor U23852 (N_23852,N_20481,N_19934);
nor U23853 (N_23853,N_20454,N_20802);
nor U23854 (N_23854,N_20966,N_20761);
or U23855 (N_23855,N_18910,N_19418);
nand U23856 (N_23856,N_19946,N_19822);
or U23857 (N_23857,N_18181,N_20577);
nand U23858 (N_23858,N_19795,N_20636);
and U23859 (N_23859,N_18386,N_19609);
or U23860 (N_23860,N_18282,N_19767);
and U23861 (N_23861,N_18132,N_19358);
nor U23862 (N_23862,N_20400,N_20296);
nor U23863 (N_23863,N_20372,N_19230);
and U23864 (N_23864,N_20139,N_20838);
xnor U23865 (N_23865,N_18367,N_20544);
xnor U23866 (N_23866,N_19393,N_20910);
nor U23867 (N_23867,N_20712,N_18182);
or U23868 (N_23868,N_19010,N_20699);
nand U23869 (N_23869,N_20471,N_20145);
nor U23870 (N_23870,N_20294,N_18201);
xor U23871 (N_23871,N_20579,N_20159);
nor U23872 (N_23872,N_18767,N_18586);
and U23873 (N_23873,N_18608,N_20503);
or U23874 (N_23874,N_18449,N_18606);
nor U23875 (N_23875,N_18340,N_20746);
or U23876 (N_23876,N_18422,N_18939);
nand U23877 (N_23877,N_20895,N_19761);
or U23878 (N_23878,N_19492,N_18572);
nor U23879 (N_23879,N_19184,N_19923);
nor U23880 (N_23880,N_19520,N_20246);
or U23881 (N_23881,N_19650,N_18130);
or U23882 (N_23882,N_18296,N_18891);
xnor U23883 (N_23883,N_19023,N_20446);
and U23884 (N_23884,N_19301,N_18948);
or U23885 (N_23885,N_18578,N_20343);
nor U23886 (N_23886,N_20388,N_20158);
xor U23887 (N_23887,N_19082,N_19707);
nor U23888 (N_23888,N_18826,N_18393);
nor U23889 (N_23889,N_20656,N_18005);
or U23890 (N_23890,N_18331,N_18611);
nand U23891 (N_23891,N_20431,N_20146);
and U23892 (N_23892,N_19119,N_20892);
nor U23893 (N_23893,N_19867,N_19935);
nand U23894 (N_23894,N_18945,N_20259);
nor U23895 (N_23895,N_20368,N_20153);
nor U23896 (N_23896,N_19377,N_20732);
nor U23897 (N_23897,N_18243,N_20268);
or U23898 (N_23898,N_20051,N_19819);
and U23899 (N_23899,N_20053,N_20792);
nand U23900 (N_23900,N_18417,N_20290);
and U23901 (N_23901,N_19140,N_18274);
or U23902 (N_23902,N_20963,N_18681);
or U23903 (N_23903,N_19208,N_18466);
xnor U23904 (N_23904,N_19662,N_20159);
nor U23905 (N_23905,N_18503,N_19819);
or U23906 (N_23906,N_20774,N_20764);
xor U23907 (N_23907,N_18588,N_20613);
nor U23908 (N_23908,N_19339,N_20042);
and U23909 (N_23909,N_18727,N_19971);
xnor U23910 (N_23910,N_20625,N_20819);
xor U23911 (N_23911,N_19085,N_18152);
nor U23912 (N_23912,N_19299,N_18512);
or U23913 (N_23913,N_20436,N_18041);
xor U23914 (N_23914,N_20108,N_18005);
and U23915 (N_23915,N_20849,N_19342);
or U23916 (N_23916,N_20474,N_20147);
and U23917 (N_23917,N_19933,N_18178);
or U23918 (N_23918,N_20082,N_18620);
or U23919 (N_23919,N_20439,N_20914);
nand U23920 (N_23920,N_18179,N_18979);
nand U23921 (N_23921,N_19656,N_19838);
and U23922 (N_23922,N_20785,N_18109);
nor U23923 (N_23923,N_19498,N_20441);
and U23924 (N_23924,N_20567,N_19723);
xnor U23925 (N_23925,N_18601,N_18743);
and U23926 (N_23926,N_20612,N_19224);
xor U23927 (N_23927,N_19286,N_20879);
and U23928 (N_23928,N_19603,N_18496);
nand U23929 (N_23929,N_19763,N_20696);
and U23930 (N_23930,N_19917,N_20365);
and U23931 (N_23931,N_20422,N_18770);
xor U23932 (N_23932,N_19702,N_20839);
nor U23933 (N_23933,N_20729,N_18342);
nor U23934 (N_23934,N_20858,N_19735);
and U23935 (N_23935,N_18555,N_20115);
xnor U23936 (N_23936,N_20554,N_19805);
or U23937 (N_23937,N_18752,N_18397);
or U23938 (N_23938,N_20207,N_19624);
xnor U23939 (N_23939,N_19656,N_20036);
nor U23940 (N_23940,N_18955,N_20299);
xnor U23941 (N_23941,N_19904,N_18544);
nand U23942 (N_23942,N_18378,N_20037);
xnor U23943 (N_23943,N_18528,N_18337);
and U23944 (N_23944,N_19588,N_19566);
and U23945 (N_23945,N_18282,N_18502);
or U23946 (N_23946,N_19493,N_18654);
nor U23947 (N_23947,N_18003,N_18548);
nand U23948 (N_23948,N_20599,N_18585);
xor U23949 (N_23949,N_18508,N_18143);
and U23950 (N_23950,N_18951,N_20433);
and U23951 (N_23951,N_20059,N_18281);
and U23952 (N_23952,N_20292,N_19656);
and U23953 (N_23953,N_18724,N_19187);
or U23954 (N_23954,N_20588,N_18702);
and U23955 (N_23955,N_19575,N_20565);
nor U23956 (N_23956,N_18548,N_19087);
or U23957 (N_23957,N_19427,N_20331);
and U23958 (N_23958,N_19723,N_20908);
or U23959 (N_23959,N_19110,N_19759);
nor U23960 (N_23960,N_20937,N_20311);
or U23961 (N_23961,N_18571,N_18787);
xor U23962 (N_23962,N_20978,N_19944);
and U23963 (N_23963,N_19166,N_18096);
and U23964 (N_23964,N_18498,N_19133);
or U23965 (N_23965,N_19951,N_20020);
xnor U23966 (N_23966,N_19315,N_18868);
nand U23967 (N_23967,N_19548,N_19986);
xnor U23968 (N_23968,N_18594,N_20330);
and U23969 (N_23969,N_20447,N_18768);
nand U23970 (N_23970,N_19468,N_18975);
xnor U23971 (N_23971,N_19717,N_20430);
nand U23972 (N_23972,N_20966,N_18353);
or U23973 (N_23973,N_19347,N_18081);
xnor U23974 (N_23974,N_19468,N_18268);
nand U23975 (N_23975,N_19149,N_20661);
nor U23976 (N_23976,N_18211,N_19867);
and U23977 (N_23977,N_20511,N_19712);
xnor U23978 (N_23978,N_20608,N_20876);
and U23979 (N_23979,N_20090,N_19714);
nand U23980 (N_23980,N_18039,N_20277);
nor U23981 (N_23981,N_20909,N_18210);
nor U23982 (N_23982,N_20293,N_18934);
or U23983 (N_23983,N_19930,N_20349);
and U23984 (N_23984,N_18913,N_20480);
or U23985 (N_23985,N_19651,N_20095);
and U23986 (N_23986,N_18538,N_20458);
xor U23987 (N_23987,N_18631,N_19797);
xor U23988 (N_23988,N_20895,N_18734);
or U23989 (N_23989,N_19912,N_20016);
and U23990 (N_23990,N_20286,N_20151);
nor U23991 (N_23991,N_20055,N_18691);
xor U23992 (N_23992,N_19598,N_20482);
nand U23993 (N_23993,N_19384,N_19421);
or U23994 (N_23994,N_19478,N_19446);
or U23995 (N_23995,N_20987,N_19345);
nor U23996 (N_23996,N_19848,N_20467);
nand U23997 (N_23997,N_20177,N_19076);
or U23998 (N_23998,N_20375,N_20217);
nor U23999 (N_23999,N_20178,N_19366);
nand U24000 (N_24000,N_21479,N_21811);
or U24001 (N_24001,N_21313,N_23790);
nor U24002 (N_24002,N_21102,N_23555);
or U24003 (N_24003,N_23257,N_22359);
or U24004 (N_24004,N_22994,N_23446);
and U24005 (N_24005,N_21756,N_21550);
and U24006 (N_24006,N_23601,N_22225);
nor U24007 (N_24007,N_22832,N_22816);
xnor U24008 (N_24008,N_22744,N_23030);
xor U24009 (N_24009,N_21019,N_23920);
or U24010 (N_24010,N_21521,N_23178);
and U24011 (N_24011,N_22356,N_22047);
and U24012 (N_24012,N_21123,N_22797);
or U24013 (N_24013,N_21600,N_22191);
xor U24014 (N_24014,N_23591,N_21296);
nand U24015 (N_24015,N_23630,N_23162);
xor U24016 (N_24016,N_22414,N_22272);
nand U24017 (N_24017,N_23596,N_23725);
xnor U24018 (N_24018,N_23055,N_21404);
or U24019 (N_24019,N_21833,N_23411);
or U24020 (N_24020,N_22656,N_23231);
nor U24021 (N_24021,N_23091,N_22624);
nor U24022 (N_24022,N_22062,N_22567);
nand U24023 (N_24023,N_21819,N_22973);
or U24024 (N_24024,N_23509,N_23093);
or U24025 (N_24025,N_21297,N_22422);
or U24026 (N_24026,N_21801,N_23439);
xnor U24027 (N_24027,N_21006,N_23215);
or U24028 (N_24028,N_23943,N_21930);
or U24029 (N_24029,N_21568,N_21117);
xor U24030 (N_24030,N_23043,N_21229);
and U24031 (N_24031,N_22507,N_21596);
nand U24032 (N_24032,N_22837,N_23075);
nor U24033 (N_24033,N_22545,N_23615);
or U24034 (N_24034,N_22658,N_22049);
nor U24035 (N_24035,N_21320,N_22565);
nor U24036 (N_24036,N_22826,N_21058);
and U24037 (N_24037,N_22841,N_21465);
or U24038 (N_24038,N_21468,N_22100);
or U24039 (N_24039,N_22636,N_23638);
nor U24040 (N_24040,N_23239,N_23900);
xnor U24041 (N_24041,N_23792,N_23424);
nor U24042 (N_24042,N_21597,N_23549);
nor U24043 (N_24043,N_23760,N_21182);
nor U24044 (N_24044,N_22364,N_23425);
xnor U24045 (N_24045,N_22587,N_23081);
nor U24046 (N_24046,N_23757,N_23076);
nor U24047 (N_24047,N_23886,N_21451);
nor U24048 (N_24048,N_21629,N_22423);
xnor U24049 (N_24049,N_22207,N_22774);
nand U24050 (N_24050,N_23336,N_22103);
nor U24051 (N_24051,N_23082,N_21408);
nor U24052 (N_24052,N_22186,N_21707);
nor U24053 (N_24053,N_21696,N_21984);
nand U24054 (N_24054,N_22685,N_21884);
or U24055 (N_24055,N_21288,N_23260);
xor U24056 (N_24056,N_23933,N_21178);
or U24057 (N_24057,N_21129,N_21033);
or U24058 (N_24058,N_22120,N_23583);
xor U24059 (N_24059,N_21350,N_23947);
and U24060 (N_24060,N_21116,N_22426);
and U24061 (N_24061,N_21781,N_23230);
nand U24062 (N_24062,N_21137,N_23267);
nor U24063 (N_24063,N_21767,N_21007);
or U24064 (N_24064,N_21131,N_21220);
nor U24065 (N_24065,N_21736,N_22132);
nand U24066 (N_24066,N_23308,N_21735);
nand U24067 (N_24067,N_22676,N_23589);
nand U24068 (N_24068,N_23536,N_21263);
nand U24069 (N_24069,N_21854,N_21349);
nand U24070 (N_24070,N_22267,N_23448);
nor U24071 (N_24071,N_22410,N_23212);
xor U24072 (N_24072,N_21905,N_22287);
xor U24073 (N_24073,N_23149,N_22501);
nand U24074 (N_24074,N_23941,N_22704);
xnor U24075 (N_24075,N_21776,N_21495);
nand U24076 (N_24076,N_22038,N_22335);
xnor U24077 (N_24077,N_22833,N_23586);
nor U24078 (N_24078,N_22851,N_21308);
or U24079 (N_24079,N_23558,N_23667);
and U24080 (N_24080,N_21954,N_23880);
and U24081 (N_24081,N_23687,N_22889);
and U24082 (N_24082,N_22828,N_23343);
or U24083 (N_24083,N_22705,N_22105);
and U24084 (N_24084,N_21793,N_21660);
and U24085 (N_24085,N_23373,N_22042);
or U24086 (N_24086,N_21744,N_23070);
nor U24087 (N_24087,N_23529,N_22275);
and U24088 (N_24088,N_22854,N_21402);
and U24089 (N_24089,N_23608,N_22714);
nor U24090 (N_24090,N_23401,N_23441);
nand U24091 (N_24091,N_23817,N_23606);
nand U24092 (N_24092,N_21725,N_21952);
and U24093 (N_24093,N_23191,N_23797);
xnor U24094 (N_24094,N_22664,N_23090);
or U24095 (N_24095,N_23501,N_21418);
nor U24096 (N_24096,N_21647,N_21514);
and U24097 (N_24097,N_23644,N_22963);
nor U24098 (N_24098,N_22790,N_21192);
nor U24099 (N_24099,N_23845,N_23242);
or U24100 (N_24100,N_22546,N_23612);
or U24101 (N_24101,N_23525,N_23289);
xor U24102 (N_24102,N_23171,N_22382);
and U24103 (N_24103,N_23557,N_23831);
nand U24104 (N_24104,N_21300,N_23154);
nand U24105 (N_24105,N_21061,N_21407);
nor U24106 (N_24106,N_22892,N_21098);
nor U24107 (N_24107,N_23695,N_23940);
nand U24108 (N_24108,N_21101,N_21574);
and U24109 (N_24109,N_23629,N_21513);
nand U24110 (N_24110,N_22617,N_23392);
and U24111 (N_24111,N_21012,N_23570);
nand U24112 (N_24112,N_21284,N_21403);
nand U24113 (N_24113,N_21005,N_23617);
xor U24114 (N_24114,N_22712,N_23318);
and U24115 (N_24115,N_22291,N_23374);
nor U24116 (N_24116,N_23378,N_22032);
and U24117 (N_24117,N_22210,N_22593);
nand U24118 (N_24118,N_21991,N_23859);
nor U24119 (N_24119,N_22258,N_21561);
or U24120 (N_24120,N_23164,N_23674);
nand U24121 (N_24121,N_22852,N_23377);
nand U24122 (N_24122,N_23944,N_23530);
nand U24123 (N_24123,N_21232,N_21648);
nor U24124 (N_24124,N_22491,N_23434);
xor U24125 (N_24125,N_21084,N_23681);
and U24126 (N_24126,N_23042,N_21873);
and U24127 (N_24127,N_22557,N_21920);
nand U24128 (N_24128,N_21569,N_21955);
or U24129 (N_24129,N_21614,N_21671);
nand U24130 (N_24130,N_23213,N_22281);
and U24131 (N_24131,N_22689,N_21014);
nor U24132 (N_24132,N_22997,N_21193);
and U24133 (N_24133,N_21380,N_23320);
nand U24134 (N_24134,N_23496,N_21079);
nor U24135 (N_24135,N_22875,N_22159);
or U24136 (N_24136,N_22900,N_22845);
nor U24137 (N_24137,N_21974,N_23243);
and U24138 (N_24138,N_21471,N_21162);
nand U24139 (N_24139,N_21743,N_22128);
nor U24140 (N_24140,N_21312,N_22820);
and U24141 (N_24141,N_21967,N_22453);
xnor U24142 (N_24142,N_22162,N_21372);
nor U24143 (N_24143,N_23670,N_22427);
or U24144 (N_24144,N_23346,N_21335);
or U24145 (N_24145,N_22778,N_23729);
and U24146 (N_24146,N_23008,N_22288);
and U24147 (N_24147,N_23906,N_23255);
xnor U24148 (N_24148,N_22663,N_22072);
nor U24149 (N_24149,N_22048,N_23568);
or U24150 (N_24150,N_22583,N_22381);
or U24151 (N_24151,N_21053,N_23172);
and U24152 (N_24152,N_21925,N_23420);
or U24153 (N_24153,N_21806,N_23248);
xor U24154 (N_24154,N_22164,N_23018);
nand U24155 (N_24155,N_21849,N_22295);
nor U24156 (N_24156,N_23651,N_21551);
and U24157 (N_24157,N_21760,N_21616);
nor U24158 (N_24158,N_21982,N_23347);
nor U24159 (N_24159,N_22595,N_22838);
xnor U24160 (N_24160,N_23510,N_23551);
nand U24161 (N_24161,N_23761,N_22400);
nor U24162 (N_24162,N_21367,N_22532);
xnor U24163 (N_24163,N_23106,N_21280);
xnor U24164 (N_24164,N_22622,N_23655);
xnor U24165 (N_24165,N_21938,N_23607);
nand U24166 (N_24166,N_23362,N_22781);
nand U24167 (N_24167,N_22987,N_23550);
or U24168 (N_24168,N_22978,N_22493);
nor U24169 (N_24169,N_21532,N_22630);
and U24170 (N_24170,N_21640,N_22478);
and U24171 (N_24171,N_22680,N_22513);
and U24172 (N_24172,N_22659,N_21695);
xnor U24173 (N_24173,N_21196,N_21037);
nand U24174 (N_24174,N_22026,N_23388);
nor U24175 (N_24175,N_22355,N_22388);
and U24176 (N_24176,N_22366,N_22347);
nor U24177 (N_24177,N_22122,N_21382);
or U24178 (N_24178,N_21893,N_22958);
nand U24179 (N_24179,N_21573,N_23495);
nand U24180 (N_24180,N_23396,N_23968);
nand U24181 (N_24181,N_23706,N_21439);
nor U24182 (N_24182,N_23581,N_22050);
and U24183 (N_24183,N_22830,N_21700);
nor U24184 (N_24184,N_21430,N_23507);
nor U24185 (N_24185,N_23497,N_21915);
nor U24186 (N_24186,N_21539,N_21771);
and U24187 (N_24187,N_21166,N_23447);
xnor U24188 (N_24188,N_21831,N_21881);
or U24189 (N_24189,N_23627,N_21322);
and U24190 (N_24190,N_23143,N_23768);
xor U24191 (N_24191,N_23486,N_21822);
xnor U24192 (N_24192,N_21840,N_22662);
nor U24193 (N_24193,N_23515,N_21205);
xor U24194 (N_24194,N_23155,N_22697);
xnor U24195 (N_24195,N_22383,N_23833);
nor U24196 (N_24196,N_21699,N_23882);
nand U24197 (N_24197,N_21655,N_23433);
nor U24198 (N_24198,N_23650,N_21935);
nand U24199 (N_24199,N_23680,N_21879);
nand U24200 (N_24200,N_22696,N_21487);
xnor U24201 (N_24201,N_22632,N_23039);
xor U24202 (N_24202,N_23460,N_22443);
or U24203 (N_24203,N_21612,N_22880);
or U24204 (N_24204,N_22971,N_23641);
nor U24205 (N_24205,N_22849,N_23244);
nand U24206 (N_24206,N_22134,N_23220);
or U24207 (N_24207,N_23827,N_22448);
and U24208 (N_24208,N_22019,N_21936);
nand U24209 (N_24209,N_22486,N_21444);
nor U24210 (N_24210,N_23288,N_21533);
nor U24211 (N_24211,N_21497,N_22435);
or U24212 (N_24212,N_23254,N_23223);
nor U24213 (N_24213,N_21460,N_22176);
and U24214 (N_24214,N_21553,N_22495);
and U24215 (N_24215,N_23986,N_21163);
nand U24216 (N_24216,N_21168,N_23079);
xor U24217 (N_24217,N_21684,N_21828);
xnor U24218 (N_24218,N_21644,N_22602);
xor U24219 (N_24219,N_22130,N_23393);
nand U24220 (N_24220,N_23562,N_22842);
nor U24221 (N_24221,N_23214,N_21804);
and U24222 (N_24222,N_22929,N_23110);
and U24223 (N_24223,N_22730,N_21637);
nor U24224 (N_24224,N_21557,N_22938);
nand U24225 (N_24225,N_23368,N_22044);
and U24226 (N_24226,N_23286,N_21703);
and U24227 (N_24227,N_22984,N_22677);
or U24228 (N_24228,N_23523,N_22165);
xnor U24229 (N_24229,N_23746,N_22279);
or U24230 (N_24230,N_21317,N_21999);
or U24231 (N_24231,N_22885,N_23716);
xnor U24232 (N_24232,N_22732,N_22957);
xor U24233 (N_24233,N_22661,N_21475);
nand U24234 (N_24234,N_21476,N_21638);
xnor U24235 (N_24235,N_22133,N_22764);
nand U24236 (N_24236,N_21266,N_23521);
nand U24237 (N_24237,N_21080,N_23022);
xnor U24238 (N_24238,N_21292,N_23619);
nor U24239 (N_24239,N_22651,N_22727);
xor U24240 (N_24240,N_23526,N_23170);
or U24241 (N_24241,N_23846,N_22319);
nand U24242 (N_24242,N_23636,N_21496);
or U24243 (N_24243,N_22761,N_23633);
nand U24244 (N_24244,N_23999,N_23634);
or U24245 (N_24245,N_22251,N_21285);
or U24246 (N_24246,N_22736,N_22910);
or U24247 (N_24247,N_22966,N_21441);
nor U24248 (N_24248,N_22488,N_23314);
nor U24249 (N_24249,N_23556,N_23136);
nor U24250 (N_24250,N_22389,N_21797);
nor U24251 (N_24251,N_22652,N_23522);
and U24252 (N_24252,N_23590,N_22175);
or U24253 (N_24253,N_22979,N_22728);
nor U24254 (N_24254,N_22230,N_21906);
xor U24255 (N_24255,N_23682,N_22215);
and U24256 (N_24256,N_23616,N_21352);
or U24257 (N_24257,N_22070,N_22882);
nand U24258 (N_24258,N_23878,N_21094);
and U24259 (N_24259,N_22260,N_23356);
nand U24260 (N_24260,N_21347,N_23796);
nand U24261 (N_24261,N_23176,N_21103);
and U24262 (N_24262,N_23594,N_22522);
nand U24263 (N_24263,N_23078,N_21040);
nor U24264 (N_24264,N_22339,N_23744);
and U24265 (N_24265,N_21179,N_22594);
and U24266 (N_24266,N_23157,N_21913);
and U24267 (N_24267,N_23868,N_21184);
and U24268 (N_24268,N_22065,N_22104);
and U24269 (N_24269,N_23531,N_23580);
nand U24270 (N_24270,N_21165,N_22850);
xor U24271 (N_24271,N_22323,N_21358);
and U24272 (N_24272,N_21555,N_23147);
nor U24273 (N_24273,N_23766,N_21688);
nor U24274 (N_24274,N_23185,N_22217);
nand U24275 (N_24275,N_22615,N_22223);
nor U24276 (N_24276,N_22596,N_22030);
xor U24277 (N_24277,N_22980,N_23745);
and U24278 (N_24278,N_22445,N_22582);
and U24279 (N_24279,N_21310,N_21332);
and U24280 (N_24280,N_21770,N_22723);
and U24281 (N_24281,N_21398,N_22800);
nor U24282 (N_24282,N_21830,N_23726);
nor U24283 (N_24283,N_21556,N_21500);
or U24284 (N_24284,N_21060,N_23552);
nand U24285 (N_24285,N_22812,N_22303);
xor U24286 (N_24286,N_22046,N_21421);
nand U24287 (N_24287,N_22311,N_22218);
nand U24288 (N_24288,N_22305,N_23351);
and U24289 (N_24289,N_21081,N_21257);
xnor U24290 (N_24290,N_21845,N_23101);
nand U24291 (N_24291,N_21966,N_22528);
nand U24292 (N_24292,N_22618,N_22671);
or U24293 (N_24293,N_22004,N_22190);
nor U24294 (N_24294,N_21151,N_21096);
xnor U24295 (N_24295,N_23739,N_23488);
nand U24296 (N_24296,N_23820,N_22406);
xnor U24297 (N_24297,N_21473,N_23696);
nand U24298 (N_24298,N_21029,N_23282);
nand U24299 (N_24299,N_23049,N_21683);
nand U24300 (N_24300,N_22243,N_23359);
or U24301 (N_24301,N_22413,N_22462);
nor U24302 (N_24302,N_21200,N_22621);
or U24303 (N_24303,N_22377,N_23537);
nor U24304 (N_24304,N_23137,N_22234);
xor U24305 (N_24305,N_21467,N_22809);
or U24306 (N_24306,N_21512,N_21715);
nand U24307 (N_24307,N_21113,N_21846);
nand U24308 (N_24308,N_22579,N_21331);
nand U24309 (N_24309,N_21713,N_23863);
and U24310 (N_24310,N_23002,N_23891);
nand U24311 (N_24311,N_22695,N_23319);
or U24312 (N_24312,N_23924,N_22315);
and U24313 (N_24313,N_22558,N_23077);
and U24314 (N_24314,N_22536,N_23724);
nor U24315 (N_24315,N_22117,N_21369);
and U24316 (N_24316,N_23112,N_21027);
and U24317 (N_24317,N_21851,N_21388);
nor U24318 (N_24318,N_21386,N_22722);
or U24319 (N_24319,N_22193,N_21134);
and U24320 (N_24320,N_23847,N_21714);
nor U24321 (N_24321,N_22642,N_23427);
xor U24322 (N_24322,N_23321,N_23543);
or U24323 (N_24323,N_23258,N_21552);
xnor U24324 (N_24324,N_23970,N_23698);
xor U24325 (N_24325,N_23186,N_21721);
xor U24326 (N_24326,N_23150,N_23436);
or U24327 (N_24327,N_23793,N_23794);
and U24328 (N_24328,N_21883,N_21021);
or U24329 (N_24329,N_21939,N_22163);
nor U24330 (N_24330,N_23519,N_22570);
and U24331 (N_24331,N_22361,N_21406);
and U24332 (N_24332,N_21252,N_23548);
xor U24333 (N_24333,N_22574,N_22917);
nor U24334 (N_24334,N_22936,N_21039);
nand U24335 (N_24335,N_22535,N_21097);
and U24336 (N_24336,N_23332,N_22846);
and U24337 (N_24337,N_23100,N_23909);
xor U24338 (N_24338,N_21273,N_23003);
or U24339 (N_24339,N_22914,N_21885);
xnor U24340 (N_24340,N_22989,N_22201);
xnor U24341 (N_24341,N_22109,N_21927);
nand U24342 (N_24342,N_22726,N_21942);
and U24343 (N_24343,N_21563,N_22282);
or U24344 (N_24344,N_23216,N_22566);
and U24345 (N_24345,N_22187,N_22221);
xnor U24346 (N_24346,N_22578,N_21302);
xor U24347 (N_24347,N_22280,N_21590);
nand U24348 (N_24348,N_22992,N_21052);
nor U24349 (N_24349,N_23104,N_23235);
xnor U24350 (N_24350,N_21669,N_22471);
xnor U24351 (N_24351,N_23652,N_22773);
nand U24352 (N_24352,N_22185,N_21436);
xor U24353 (N_24353,N_22033,N_22896);
or U24354 (N_24354,N_21412,N_23587);
or U24355 (N_24355,N_22083,N_21914);
and U24356 (N_24356,N_23065,N_23544);
xnor U24357 (N_24357,N_23457,N_22902);
nand U24358 (N_24358,N_21070,N_21236);
xnor U24359 (N_24359,N_23367,N_22371);
or U24360 (N_24360,N_23639,N_21717);
and U24361 (N_24361,N_21454,N_23249);
xor U24362 (N_24362,N_23857,N_21869);
nor U24363 (N_24363,N_23097,N_22603);
and U24364 (N_24364,N_22283,N_23038);
or U24365 (N_24365,N_22073,N_21843);
xor U24366 (N_24366,N_22296,N_21216);
nand U24367 (N_24367,N_22467,N_23099);
and U24368 (N_24368,N_21839,N_21405);
or U24369 (N_24369,N_21803,N_21578);
and U24370 (N_24370,N_22153,N_22150);
and U24371 (N_24371,N_22748,N_23115);
nand U24372 (N_24372,N_22052,N_21209);
xor U24373 (N_24373,N_23264,N_23747);
xor U24374 (N_24374,N_23754,N_22156);
nand U24375 (N_24375,N_22344,N_22506);
and U24376 (N_24376,N_21321,N_22612);
xor U24377 (N_24377,N_21316,N_23822);
nor U24378 (N_24378,N_22893,N_23413);
and U24379 (N_24379,N_21022,N_22148);
nor U24380 (N_24380,N_23429,N_23265);
and U24381 (N_24381,N_21900,N_23340);
nand U24382 (N_24382,N_23490,N_23858);
and U24383 (N_24383,N_22224,N_23094);
xnor U24384 (N_24384,N_23764,N_21259);
nor U24385 (N_24385,N_22666,N_23089);
or U24386 (N_24386,N_21836,N_23598);
nand U24387 (N_24387,N_22657,N_23168);
and U24388 (N_24388,N_21718,N_22941);
or U24389 (N_24389,N_22804,N_23603);
xnor U24390 (N_24390,N_22235,N_21445);
xnor U24391 (N_24391,N_23435,N_22365);
or U24392 (N_24392,N_21706,N_21904);
or U24393 (N_24393,N_23997,N_23454);
xnor U24394 (N_24394,N_23275,N_22729);
nor U24395 (N_24395,N_23132,N_21924);
and U24396 (N_24396,N_23114,N_21780);
nor U24397 (N_24397,N_22840,N_23232);
nand U24398 (N_24398,N_21946,N_22379);
xnor U24399 (N_24399,N_23421,N_22953);
or U24400 (N_24400,N_21132,N_22908);
and U24401 (N_24401,N_23417,N_23190);
nand U24402 (N_24402,N_23934,N_23158);
nor U24403 (N_24403,N_21197,N_21493);
nand U24404 (N_24404,N_22437,N_22808);
nand U24405 (N_24405,N_22449,N_23410);
and U24406 (N_24406,N_21384,N_21633);
nand U24407 (N_24407,N_21230,N_21888);
or U24408 (N_24408,N_23668,N_22484);
and U24409 (N_24409,N_21844,N_23012);
nand U24410 (N_24410,N_23160,N_23966);
nand U24411 (N_24411,N_23678,N_21664);
nand U24412 (N_24412,N_21701,N_23217);
or U24413 (N_24413,N_22742,N_22029);
nand U24414 (N_24414,N_22394,N_23708);
xnor U24415 (N_24415,N_21339,N_21581);
or U24416 (N_24416,N_21459,N_23498);
or U24417 (N_24417,N_23161,N_22325);
xor U24418 (N_24418,N_21621,N_21566);
nor U24419 (N_24419,N_22068,N_21492);
and U24420 (N_24420,N_21741,N_23414);
nand U24421 (N_24421,N_21376,N_22274);
nand U24422 (N_24422,N_22644,N_21737);
nand U24423 (N_24423,N_22784,N_22789);
and U24424 (N_24424,N_22011,N_23480);
or U24425 (N_24425,N_23034,N_23053);
and U24426 (N_24426,N_21413,N_21035);
nand U24427 (N_24427,N_23928,N_22015);
xor U24428 (N_24428,N_21792,N_21753);
and U24429 (N_24429,N_21242,N_22829);
nand U24430 (N_24430,N_22711,N_23957);
nand U24431 (N_24431,N_23426,N_23506);
and U24432 (N_24432,N_23218,N_22554);
xnor U24433 (N_24433,N_22972,N_23602);
nor U24434 (N_24434,N_23409,N_21528);
or U24435 (N_24435,N_21976,N_23663);
nor U24436 (N_24436,N_21447,N_22160);
xnor U24437 (N_24437,N_21054,N_22779);
nor U24438 (N_24438,N_22475,N_22360);
or U24439 (N_24439,N_23743,N_23348);
or U24440 (N_24440,N_23202,N_23107);
nand U24441 (N_24441,N_22860,N_22031);
xnor U24442 (N_24442,N_21450,N_22678);
xor U24443 (N_24443,N_22284,N_22597);
or U24444 (N_24444,N_23534,N_21545);
nand U24445 (N_24445,N_21586,N_23406);
nand U24446 (N_24446,N_21774,N_22805);
and U24447 (N_24447,N_23415,N_23326);
nand U24448 (N_24448,N_21902,N_22839);
and U24449 (N_24449,N_22527,N_21003);
or U24450 (N_24450,N_21505,N_22127);
nand U24451 (N_24451,N_21141,N_21702);
nand U24452 (N_24452,N_22990,N_21298);
nor U24453 (N_24453,N_21301,N_23705);
and U24454 (N_24454,N_23948,N_22718);
xnor U24455 (N_24455,N_21896,N_22584);
or U24456 (N_24456,N_23983,N_22205);
or U24457 (N_24457,N_23227,N_21758);
nor U24458 (N_24458,N_22036,N_22197);
and U24459 (N_24459,N_22158,N_23801);
and U24460 (N_24460,N_21368,N_22009);
xnor U24461 (N_24461,N_23103,N_21120);
or U24462 (N_24462,N_21728,N_22717);
or U24463 (N_24463,N_22928,N_23390);
xor U24464 (N_24464,N_23786,N_23124);
or U24465 (N_24465,N_23799,N_21944);
and U24466 (N_24466,N_23956,N_23753);
nor U24467 (N_24467,N_22312,N_22329);
nand U24468 (N_24468,N_23328,N_22873);
xor U24469 (N_24469,N_23016,N_22749);
xor U24470 (N_24470,N_21517,N_22906);
and U24471 (N_24471,N_21279,N_21289);
or U24472 (N_24472,N_22460,N_21891);
nor U24473 (N_24473,N_23198,N_23571);
xnor U24474 (N_24474,N_21338,N_21150);
xor U24475 (N_24475,N_21329,N_23814);
and U24476 (N_24476,N_23085,N_23330);
nand U24477 (N_24477,N_22257,N_23095);
or U24478 (N_24478,N_21112,N_23350);
nand U24479 (N_24479,N_22376,N_22681);
xor U24480 (N_24480,N_21693,N_22635);
and U24481 (N_24481,N_22517,N_21678);
and U24482 (N_24482,N_22701,N_23502);
and U24483 (N_24483,N_23385,N_23324);
and U24484 (N_24484,N_22226,N_22599);
nand U24485 (N_24485,N_23818,N_21853);
xnor U24486 (N_24486,N_22866,N_23762);
or U24487 (N_24487,N_21139,N_21463);
or U24488 (N_24488,N_22682,N_21727);
or U24489 (N_24489,N_23383,N_23669);
nor U24490 (N_24490,N_22813,N_22183);
nand U24491 (N_24491,N_21618,N_23062);
or U24492 (N_24492,N_22440,N_23665);
nand U24493 (N_24493,N_21625,N_21950);
or U24494 (N_24494,N_22300,N_23399);
xor U24495 (N_24495,N_23666,N_22707);
nand U24496 (N_24496,N_22920,N_23808);
nand U24497 (N_24497,N_23684,N_21227);
nor U24498 (N_24498,N_21363,N_23785);
or U24499 (N_24499,N_21195,N_22687);
or U24500 (N_24500,N_21941,N_21820);
nand U24501 (N_24501,N_22821,N_22057);
xnor U24502 (N_24502,N_23823,N_21158);
nand U24503 (N_24503,N_22559,N_21656);
and U24504 (N_24504,N_22182,N_21865);
xor U24505 (N_24505,N_23844,N_23481);
or U24506 (N_24506,N_22619,N_23713);
or U24507 (N_24507,N_23930,N_23397);
or U24508 (N_24508,N_23691,N_22328);
nand U24509 (N_24509,N_23423,N_21142);
and U24510 (N_24510,N_23758,N_22686);
or U24511 (N_24511,N_21940,N_23896);
xor U24512 (N_24512,N_23365,N_23912);
xnor U24513 (N_24513,N_21639,N_21658);
xor U24514 (N_24514,N_21958,N_22337);
xor U24515 (N_24515,N_22084,N_21087);
nor U24516 (N_24516,N_21215,N_21127);
or U24517 (N_24517,N_23233,N_22350);
nand U24518 (N_24518,N_22262,N_22306);
nor U24519 (N_24519,N_22434,N_22149);
xor U24520 (N_24520,N_21272,N_22095);
nor U24521 (N_24521,N_21387,N_23123);
nand U24522 (N_24522,N_23125,N_21580);
nand U24523 (N_24523,N_23102,N_21603);
or U24524 (N_24524,N_22118,N_21378);
or U24525 (N_24525,N_22188,N_23752);
nor U24526 (N_24526,N_21038,N_23297);
xor U24527 (N_24527,N_21417,N_21410);
and U24528 (N_24528,N_23440,N_22420);
and U24529 (N_24529,N_22320,N_22169);
xnor U24530 (N_24530,N_23019,N_23499);
nand U24531 (N_24531,N_23969,N_21542);
nor U24532 (N_24532,N_21558,N_22219);
and U24533 (N_24533,N_23174,N_21013);
or U24534 (N_24534,N_22757,N_21211);
nor U24535 (N_24535,N_21244,N_22646);
nand U24536 (N_24536,N_21825,N_21504);
xnor U24537 (N_24537,N_22913,N_21892);
nor U24538 (N_24538,N_21208,N_23564);
and U24539 (N_24539,N_23628,N_23058);
xnor U24540 (N_24540,N_23211,N_22497);
or U24541 (N_24541,N_21969,N_23777);
or U24542 (N_24542,N_23253,N_22867);
and U24543 (N_24543,N_21399,N_22534);
or U24544 (N_24544,N_23711,N_21499);
nor U24545 (N_24545,N_23138,N_23001);
xor U24546 (N_24546,N_23166,N_23841);
or U24547 (N_24547,N_22968,N_21996);
or U24548 (N_24548,N_23395,N_22631);
and U24549 (N_24549,N_21795,N_23563);
nand U24550 (N_24550,N_23806,N_23927);
nor U24551 (N_24551,N_21235,N_21929);
nand U24552 (N_24552,N_23904,N_23925);
nand U24553 (N_24553,N_23072,N_22314);
and U24554 (N_24554,N_21325,N_21130);
nand U24555 (N_24555,N_21243,N_21485);
or U24556 (N_24556,N_22012,N_21138);
or U24557 (N_24557,N_21796,N_21359);
or U24558 (N_24558,N_22823,N_23482);
and U24559 (N_24559,N_21095,N_23492);
nand U24560 (N_24560,N_23014,N_21253);
and U24561 (N_24561,N_23236,N_23259);
or U24562 (N_24562,N_23572,N_21354);
or U24563 (N_24563,N_23988,N_23825);
xnor U24564 (N_24564,N_23671,N_22514);
nor U24565 (N_24565,N_22798,N_21972);
and U24566 (N_24566,N_23241,N_21870);
nand U24567 (N_24567,N_23991,N_23702);
nor U24568 (N_24568,N_21501,N_21198);
or U24569 (N_24569,N_22576,N_22321);
or U24570 (N_24570,N_21690,N_21309);
nand U24571 (N_24571,N_21419,N_21240);
nand U24572 (N_24572,N_22111,N_23251);
nor U24573 (N_24573,N_22088,N_22604);
or U24574 (N_24574,N_21383,N_23875);
nor U24575 (N_24575,N_22611,N_22137);
and U24576 (N_24576,N_22556,N_21149);
xnor U24577 (N_24577,N_22451,N_21990);
nor U24578 (N_24578,N_21304,N_23914);
nor U24579 (N_24579,N_22709,N_22327);
nor U24580 (N_24580,N_23605,N_22396);
nand U24581 (N_24581,N_21788,N_21278);
nand U24582 (N_24582,N_22212,N_21085);
xor U24583 (N_24583,N_21281,N_21871);
nand U24584 (N_24584,N_22463,N_21508);
nand U24585 (N_24585,N_23366,N_22930);
or U24586 (N_24586,N_22770,N_23372);
xor U24587 (N_24587,N_23701,N_22096);
nor U24588 (N_24588,N_23913,N_22285);
or U24589 (N_24589,N_23000,N_23048);
nand U24590 (N_24590,N_23197,N_21008);
nor U24591 (N_24591,N_21857,N_22214);
nand U24592 (N_24592,N_21221,N_22367);
nand U24593 (N_24593,N_21837,N_22575);
nand U24594 (N_24594,N_22452,N_22056);
nand U24595 (N_24595,N_22123,N_23391);
or U24596 (N_24596,N_23011,N_22259);
nand U24597 (N_24597,N_21004,N_22871);
nand U24598 (N_24598,N_21609,N_22179);
nand U24599 (N_24599,N_22154,N_21047);
nor U24600 (N_24600,N_22375,N_21663);
and U24601 (N_24601,N_22572,N_23907);
and U24602 (N_24602,N_22907,N_22060);
and U24603 (N_24603,N_23290,N_23092);
and U24604 (N_24604,N_22625,N_22023);
and U24605 (N_24605,N_21453,N_21104);
nand U24606 (N_24606,N_23119,N_23405);
and U24607 (N_24607,N_22549,N_23040);
or U24608 (N_24608,N_23505,N_23748);
nand U24609 (N_24609,N_21228,N_22919);
and U24610 (N_24610,N_21147,N_23029);
nor U24611 (N_24611,N_23033,N_21143);
nand U24612 (N_24612,N_21790,N_22981);
or U24613 (N_24613,N_21549,N_22020);
nand U24614 (N_24614,N_21456,N_21234);
or U24615 (N_24615,N_21370,N_21634);
nor U24616 (N_24616,N_22933,N_23542);
xor U24617 (N_24617,N_23310,N_21978);
nand U24618 (N_24618,N_22945,N_22141);
and U24619 (N_24619,N_23998,N_23193);
and U24620 (N_24620,N_21423,N_21897);
xor U24621 (N_24621,N_21903,N_22759);
nor U24622 (N_24622,N_21011,N_21159);
and U24623 (N_24623,N_22144,N_23201);
and U24624 (N_24624,N_21814,N_22824);
and U24625 (N_24625,N_21623,N_23296);
nor U24626 (N_24626,N_23990,N_23730);
and U24627 (N_24627,N_21214,N_22660);
xnor U24628 (N_24628,N_23838,N_23915);
and U24629 (N_24629,N_21344,N_22151);
nor U24630 (N_24630,N_22270,N_23645);
nor U24631 (N_24631,N_21617,N_23276);
nor U24632 (N_24632,N_22035,N_23658);
nand U24633 (N_24633,N_23341,N_21435);
xnor U24634 (N_24634,N_22338,N_21020);
or U24635 (N_24635,N_23908,N_22904);
and U24636 (N_24636,N_22131,N_22857);
or U24637 (N_24637,N_22861,N_21583);
nor U24638 (N_24638,N_23697,N_23309);
nor U24639 (N_24639,N_21443,N_21821);
xor U24640 (N_24640,N_22702,N_21348);
nor U24641 (N_24641,N_21507,N_21478);
or U24642 (N_24642,N_23980,N_21125);
nor U24643 (N_24643,N_23905,N_23673);
or U24644 (N_24644,N_21691,N_21917);
xor U24645 (N_24645,N_23520,N_23533);
or U24646 (N_24646,N_21224,N_21815);
or U24647 (N_24647,N_23010,N_22793);
and U24648 (N_24648,N_21685,N_23659);
nand U24649 (N_24649,N_23451,N_23491);
xor U24650 (N_24650,N_23006,N_21682);
or U24651 (N_24651,N_23210,N_22949);
or U24652 (N_24652,N_23398,N_23717);
nor U24653 (N_24653,N_21567,N_21028);
nand U24654 (N_24654,N_22878,N_22962);
nand U24655 (N_24655,N_22606,N_22518);
and U24656 (N_24656,N_22806,N_21074);
and U24657 (N_24657,N_23361,N_22627);
and U24658 (N_24658,N_22431,N_22553);
or U24659 (N_24659,N_21654,N_23953);
nand U24660 (N_24660,N_23584,N_21745);
nand U24661 (N_24661,N_22353,N_21470);
nor U24662 (N_24662,N_21661,N_23830);
nand U24663 (N_24663,N_23338,N_23349);
nor U24664 (N_24664,N_22129,N_21140);
and U24665 (N_24665,N_21631,N_21286);
nand U24666 (N_24666,N_21863,N_22927);
and U24667 (N_24667,N_22265,N_21250);
nand U24668 (N_24668,N_23977,N_21480);
and U24669 (N_24669,N_22340,N_21816);
nand U24670 (N_24670,N_23237,N_21522);
nor U24671 (N_24671,N_23005,N_22231);
nor U24672 (N_24672,N_21615,N_22373);
xor U24673 (N_24673,N_23849,N_23778);
and U24674 (N_24674,N_22061,N_23899);
nor U24675 (N_24675,N_23850,N_23751);
nor U24676 (N_24676,N_21254,N_22716);
or U24677 (N_24677,N_21088,N_22537);
and U24678 (N_24678,N_22037,N_23122);
nor U24679 (N_24679,N_21813,N_23069);
xnor U24680 (N_24680,N_22147,N_23204);
and U24681 (N_24681,N_22316,N_22836);
nand U24682 (N_24682,N_22161,N_23809);
or U24683 (N_24683,N_21315,N_23113);
nand U24684 (N_24684,N_21687,N_23574);
xnor U24685 (N_24685,N_22903,N_21506);
nor U24686 (N_24686,N_23560,N_23445);
xnor U24687 (N_24687,N_22509,N_23653);
or U24688 (N_24688,N_21210,N_22357);
nand U24689 (N_24689,N_23517,N_23791);
nand U24690 (N_24690,N_22157,N_21798);
nor U24691 (N_24691,N_23469,N_21241);
nor U24692 (N_24692,N_21345,N_22530);
or U24693 (N_24693,N_23503,N_23468);
nor U24694 (N_24694,N_22782,N_23493);
nand U24695 (N_24695,N_22034,N_21161);
nor U24696 (N_24696,N_22894,N_22418);
xnor U24697 (N_24697,N_21670,N_23450);
xnor U24698 (N_24698,N_23609,N_23299);
and U24699 (N_24699,N_22380,N_23699);
or U24700 (N_24700,N_22719,N_22093);
nor U24701 (N_24701,N_21356,N_21099);
xor U24702 (N_24702,N_21759,N_22074);
nor U24703 (N_24703,N_22001,N_22239);
nand U24704 (N_24704,N_22318,N_22482);
nor U24705 (N_24705,N_21544,N_22741);
and U24706 (N_24706,N_21630,N_22673);
or U24707 (N_24707,N_22645,N_23470);
and U24708 (N_24708,N_23461,N_23994);
nor U24709 (N_24709,N_21526,N_21303);
nand U24710 (N_24710,N_21858,N_21527);
nand U24711 (N_24711,N_23465,N_21748);
nor U24712 (N_24712,N_21739,N_22276);
nand U24713 (N_24713,N_21679,N_22054);
and U24714 (N_24714,N_23026,N_21752);
xor U24715 (N_24715,N_23832,N_22516);
nor U24716 (N_24716,N_21740,N_21694);
xor U24717 (N_24717,N_21337,N_22417);
xnor U24718 (N_24718,N_21992,N_23789);
nand U24719 (N_24719,N_21225,N_23293);
or U24720 (N_24720,N_21789,N_23487);
or U24721 (N_24721,N_21746,N_23304);
and U24722 (N_24722,N_21311,N_23610);
xor U24723 (N_24723,N_23200,N_23203);
xnor U24724 (N_24724,N_22058,N_22326);
and U24725 (N_24725,N_23834,N_23815);
and U24726 (N_24726,N_23626,N_23955);
nor U24727 (N_24727,N_23052,N_22633);
nand U24728 (N_24728,N_21653,N_23027);
nor U24729 (N_24729,N_22189,N_22924);
and U24730 (N_24730,N_21810,N_22346);
or U24731 (N_24731,N_23921,N_22762);
nand U24732 (N_24732,N_23061,N_22540);
or U24733 (N_24733,N_21852,N_21628);
nand U24734 (N_24734,N_21520,N_21391);
nand U24735 (N_24735,N_21959,N_21156);
or U24736 (N_24736,N_21726,N_23206);
or U24737 (N_24737,N_21698,N_21270);
and U24738 (N_24738,N_21983,N_22835);
nor U24739 (N_24739,N_23084,N_23950);
nor U24740 (N_24740,N_22521,N_22985);
or U24741 (N_24741,N_21981,N_22469);
and U24742 (N_24742,N_23518,N_21223);
nand U24743 (N_24743,N_22403,N_21203);
xnor U24744 (N_24744,N_23618,N_21173);
nor U24745 (N_24745,N_23611,N_22787);
and U24746 (N_24746,N_21750,N_23295);
xnor U24747 (N_24747,N_23889,N_23946);
xnor U24748 (N_24748,N_23494,N_22424);
or U24749 (N_24749,N_23938,N_22562);
or U24750 (N_24750,N_21856,N_22679);
nand U24751 (N_24751,N_22947,N_21861);
nor U24752 (N_24752,N_22825,N_23181);
nor U24753 (N_24753,N_23222,N_21091);
nor U24754 (N_24754,N_21207,N_21146);
nand U24755 (N_24755,N_21709,N_23238);
nor U24756 (N_24756,N_23353,N_23776);
xor U24757 (N_24757,N_22580,N_21779);
or U24758 (N_24758,N_21076,N_23041);
nand U24759 (N_24759,N_21961,N_23898);
and U24760 (N_24760,N_21167,N_23428);
xnor U24761 (N_24761,N_22703,N_23298);
nand U24762 (N_24762,N_21360,N_21488);
nor U24763 (N_24763,N_23245,N_22724);
nand U24764 (N_24764,N_22006,N_23767);
and U24765 (N_24765,N_21264,N_21923);
nand U24766 (N_24766,N_21199,N_23614);
xnor U24767 (N_24767,N_21876,N_21262);
nor U24768 (N_24768,N_23959,N_22253);
xnor U24769 (N_24769,N_23305,N_23207);
nor U24770 (N_24770,N_22766,N_21543);
nor U24771 (N_24771,N_23703,N_22745);
nand U24772 (N_24772,N_22801,N_23219);
or U24773 (N_24773,N_22476,N_23404);
nand U24774 (N_24774,N_23919,N_21608);
nor U24775 (N_24775,N_22483,N_23693);
nand U24776 (N_24776,N_23331,N_21775);
and U24777 (N_24777,N_21299,N_23578);
and U24778 (N_24778,N_23978,N_23810);
nor U24779 (N_24779,N_22236,N_23648);
nand U24780 (N_24780,N_23133,N_23828);
nand U24781 (N_24781,N_22609,N_21791);
and U24782 (N_24782,N_21114,N_21336);
and U24783 (N_24783,N_22733,N_21868);
xnor U24784 (N_24784,N_23325,N_22099);
or U24785 (N_24785,N_23992,N_22974);
nor U24786 (N_24786,N_22877,N_21484);
xnor U24787 (N_24787,N_23672,N_23861);
and U24788 (N_24788,N_22891,N_23782);
nor U24789 (N_24789,N_23452,N_21457);
and U24790 (N_24790,N_23853,N_23654);
xor U24791 (N_24791,N_21018,N_23117);
or U24792 (N_24792,N_21364,N_22087);
nand U24793 (N_24793,N_23159,N_23004);
nand U24794 (N_24794,N_22975,N_23271);
xnor U24795 (N_24795,N_22152,N_21841);
nand U24796 (N_24796,N_21710,N_21908);
or U24797 (N_24797,N_22097,N_23013);
xnor U24798 (N_24798,N_22456,N_23892);
or U24799 (N_24799,N_22459,N_22430);
xor U24800 (N_24800,N_22174,N_23683);
nand U24801 (N_24801,N_22264,N_22263);
or U24802 (N_24802,N_23842,N_21455);
or U24803 (N_24803,N_22415,N_22292);
or U24804 (N_24804,N_22102,N_21188);
xor U24805 (N_24805,N_22799,N_21073);
nand U24806 (N_24806,N_22412,N_22091);
or U24807 (N_24807,N_21000,N_23685);
and U24808 (N_24808,N_23922,N_21065);
xnor U24809 (N_24809,N_21763,N_23877);
xnor U24810 (N_24810,N_22693,N_21148);
and U24811 (N_24811,N_21483,N_23962);
xnor U24812 (N_24812,N_21922,N_21481);
and U24813 (N_24813,N_23187,N_23430);
and U24814 (N_24814,N_21847,N_23600);
xnor U24815 (N_24815,N_23513,N_23694);
nand U24816 (N_24816,N_23532,N_23156);
nor U24817 (N_24817,N_21078,N_23167);
xor U24818 (N_24818,N_23478,N_23036);
and U24819 (N_24819,N_23989,N_21559);
nor U24820 (N_24820,N_21732,N_23545);
xnor U24821 (N_24821,N_23649,N_21762);
xor U24822 (N_24822,N_22464,N_21420);
or U24823 (N_24823,N_22585,N_23128);
or U24824 (N_24824,N_23142,N_21046);
or U24825 (N_24825,N_23916,N_22785);
nand U24826 (N_24826,N_21170,N_23246);
or U24827 (N_24827,N_22811,N_21864);
and U24828 (N_24828,N_21659,N_23873);
and U24829 (N_24829,N_21716,N_22114);
nand U24830 (N_24830,N_21133,N_23982);
nand U24831 (N_24831,N_23588,N_23964);
nand U24832 (N_24832,N_23247,N_23677);
xor U24833 (N_24833,N_22746,N_22655);
xnor U24834 (N_24834,N_21626,N_22937);
xnor U24835 (N_24835,N_21850,N_22411);
nand U24836 (N_24836,N_23194,N_21987);
nor U24837 (N_24837,N_23432,N_22993);
nor U24838 (N_24838,N_22950,N_21307);
nor U24839 (N_24839,N_21995,N_21290);
nor U24840 (N_24840,N_23354,N_22868);
and U24841 (N_24841,N_22043,N_23234);
nor U24842 (N_24842,N_22195,N_22967);
xor U24843 (N_24843,N_23807,N_21515);
nor U24844 (N_24844,N_23508,N_23573);
or U24845 (N_24845,N_21239,N_23540);
and U24846 (N_24846,N_21276,N_21034);
and U24847 (N_24847,N_22803,N_22322);
nor U24848 (N_24848,N_22571,N_21206);
nand U24849 (N_24849,N_21466,N_22017);
or U24850 (N_24850,N_23418,N_21002);
and U24851 (N_24851,N_22756,N_22954);
xor U24852 (N_24852,N_22614,N_23139);
nand U24853 (N_24853,N_21887,N_21832);
xnor U24854 (N_24854,N_21547,N_23360);
xor U24855 (N_24855,N_22755,N_23675);
nor U24856 (N_24856,N_22751,N_22923);
and U24857 (N_24857,N_21189,N_21152);
xor U24858 (N_24858,N_21986,N_23826);
nor U24859 (N_24859,N_21202,N_22085);
or U24860 (N_24860,N_23145,N_21931);
xor U24861 (N_24861,N_22302,N_23559);
nor U24862 (N_24862,N_22921,N_23967);
nand U24863 (N_24863,N_23307,N_23582);
nor U24864 (N_24864,N_21009,N_21442);
nand U24865 (N_24865,N_22368,N_22960);
or U24866 (N_24866,N_22998,N_23303);
nand U24867 (N_24867,N_22266,N_21645);
nor U24868 (N_24868,N_23881,N_22405);
nor U24869 (N_24869,N_21169,N_21275);
nand U24870 (N_24870,N_21595,N_22063);
and U24871 (N_24871,N_22079,N_23449);
or U24872 (N_24872,N_22758,N_22252);
or U24873 (N_24873,N_22352,N_21247);
and U24874 (N_24874,N_23358,N_23848);
or U24875 (N_24875,N_22010,N_23431);
nand U24876 (N_24876,N_21599,N_21899);
and U24877 (N_24877,N_22441,N_23829);
and U24878 (N_24878,N_22818,N_21960);
and U24879 (N_24879,N_23784,N_21686);
or U24880 (N_24880,N_23802,N_23477);
xnor U24881 (N_24881,N_23466,N_21805);
nor U24882 (N_24882,N_23270,N_22249);
xnor U24883 (N_24883,N_21911,N_21268);
and U24884 (N_24884,N_22740,N_23083);
nand U24885 (N_24885,N_21346,N_23263);
nor U24886 (N_24886,N_21947,N_21800);
and U24887 (N_24887,N_22855,N_22988);
xnor U24888 (N_24888,N_22970,N_21049);
nor U24889 (N_24889,N_21673,N_21491);
nor U24890 (N_24890,N_21525,N_22592);
nor U24891 (N_24891,N_21464,N_22121);
nand U24892 (N_24892,N_23007,N_21531);
xor U24893 (N_24893,N_23071,N_23268);
or U24894 (N_24894,N_21026,N_22763);
nor U24895 (N_24895,N_22089,N_21829);
xor U24896 (N_24896,N_23592,N_21855);
or U24897 (N_24897,N_22641,N_21016);
and U24898 (N_24898,N_22308,N_23126);
nand U24899 (N_24899,N_22881,N_22783);
xor U24900 (N_24900,N_23208,N_21509);
nor U24901 (N_24901,N_23939,N_23118);
nand U24902 (N_24902,N_22108,N_23597);
nand U24903 (N_24903,N_23737,N_21882);
or U24904 (N_24904,N_22991,N_21564);
xnor U24905 (N_24905,N_21190,N_22241);
xnor U24906 (N_24906,N_23344,N_21666);
or U24907 (N_24907,N_23342,N_22203);
or U24908 (N_24908,N_22639,N_21646);
nor U24909 (N_24909,N_23472,N_21246);
nand U24910 (N_24910,N_22995,N_21622);
nand U24911 (N_24911,N_23316,N_23266);
nand U24912 (N_24912,N_23527,N_22391);
nand U24913 (N_24913,N_21571,N_22045);
nor U24914 (N_24914,N_21341,N_21396);
and U24915 (N_24915,N_23676,N_23273);
nor U24916 (N_24916,N_21063,N_23903);
xnor U24917 (N_24917,N_21069,N_21588);
nor U24918 (N_24918,N_22468,N_23444);
or U24919 (N_24919,N_23736,N_22699);
or U24920 (N_24920,N_22935,N_22568);
and U24921 (N_24921,N_21237,N_23804);
or U24922 (N_24922,N_22647,N_23951);
xor U24923 (N_24923,N_23144,N_21469);
nor U24924 (N_24924,N_23689,N_23108);
and U24925 (N_24925,N_23322,N_21649);
xor U24926 (N_24926,N_23954,N_23613);
nand U24927 (N_24927,N_22286,N_23819);
xor U24928 (N_24928,N_22387,N_23541);
or U24929 (N_24929,N_21541,N_21546);
or U24930 (N_24930,N_23661,N_23554);
xnor U24931 (N_24931,N_22028,N_21083);
xor U24932 (N_24932,N_23942,N_23524);
nand U24933 (N_24933,N_21962,N_21374);
xor U24934 (N_24934,N_22649,N_22027);
and U24935 (N_24935,N_23840,N_23895);
nand U24936 (N_24936,N_23787,N_21357);
nor U24937 (N_24937,N_22354,N_22909);
nor U24938 (N_24938,N_21570,N_21045);
xnor U24939 (N_24939,N_22481,N_22498);
xor U24940 (N_24940,N_23993,N_22080);
xnor U24941 (N_24941,N_22489,N_23750);
and U24942 (N_24942,N_21373,N_21267);
nand U24943 (N_24943,N_22858,N_21572);
nand U24944 (N_24944,N_21217,N_21916);
nand U24945 (N_24945,N_22713,N_21607);
or U24946 (N_24946,N_22330,N_22177);
nand U24947 (N_24947,N_21434,N_21201);
or U24948 (N_24948,N_23727,N_23473);
nor U24949 (N_24949,N_22238,N_22623);
or U24950 (N_24950,N_22003,N_22005);
and U24951 (N_24951,N_21901,N_23274);
nand U24952 (N_24952,N_23285,N_22555);
and U24953 (N_24953,N_23569,N_21089);
nor U24954 (N_24954,N_22772,N_23623);
nand U24955 (N_24955,N_22959,N_23824);
nor U24956 (N_24956,N_22390,N_21111);
xnor U24957 (N_24957,N_22884,N_23291);
xor U24958 (N_24958,N_22229,N_23096);
nor U24959 (N_24959,N_22817,N_21503);
nor U24960 (N_24960,N_22098,N_22654);
nand U24961 (N_24961,N_23874,N_21393);
or U24962 (N_24962,N_23302,N_23852);
or U24963 (N_24963,N_22171,N_21105);
nor U24964 (N_24964,N_21973,N_23375);
and U24965 (N_24965,N_22810,N_21965);
or U24966 (N_24966,N_21668,N_21970);
or U24967 (N_24967,N_23779,N_21400);
nor U24968 (N_24968,N_21024,N_21604);
nand U24969 (N_24969,N_23152,N_21511);
or U24970 (N_24970,N_23514,N_23884);
and U24971 (N_24971,N_22951,N_22216);
or U24972 (N_24972,N_23333,N_22538);
xnor U24973 (N_24973,N_21353,N_23734);
nor U24974 (N_24974,N_21385,N_21536);
or U24975 (N_24975,N_23839,N_21642);
nor U24976 (N_24976,N_21827,N_21429);
or U24977 (N_24977,N_21226,N_22106);
nand U24978 (N_24978,N_23585,N_22586);
and U24979 (N_24979,N_21953,N_23538);
nor U24980 (N_24980,N_22250,N_22242);
or U24981 (N_24981,N_21477,N_23419);
nand U24982 (N_24982,N_21537,N_21390);
nor U24983 (N_24983,N_23700,N_21422);
nand U24984 (N_24984,N_23788,N_23467);
or U24985 (N_24985,N_22533,N_23742);
xor U24986 (N_24986,N_21747,N_22466);
xnor U24987 (N_24987,N_23973,N_21784);
nand U24988 (N_24988,N_23604,N_23960);
nor U24989 (N_24989,N_22948,N_21050);
or U24990 (N_24990,N_22374,N_22940);
nand U24991 (N_24991,N_23576,N_23917);
xnor U24992 (N_24992,N_22244,N_21918);
xor U24993 (N_24993,N_23169,N_22393);
or U24994 (N_24994,N_23455,N_21183);
nand U24995 (N_24995,N_21090,N_23707);
xor U24996 (N_24996,N_23067,N_23996);
nor U24997 (N_24997,N_23890,N_23479);
or U24998 (N_24998,N_21665,N_23199);
xnor U24999 (N_24999,N_23769,N_23935);
xnor U25000 (N_25000,N_21562,N_21394);
and U25001 (N_25001,N_21001,N_22386);
nand U25002 (N_25002,N_22939,N_22688);
xnor U25003 (N_25003,N_23599,N_22931);
or U25004 (N_25004,N_22946,N_22996);
and U25005 (N_25005,N_22094,N_21397);
or U25006 (N_25006,N_21823,N_22569);
xnor U25007 (N_25007,N_23363,N_23883);
nor U25008 (N_25008,N_23105,N_22317);
nand U25009 (N_25009,N_22007,N_23625);
or U25010 (N_25010,N_22600,N_22547);
or U25011 (N_25011,N_21761,N_22181);
xnor U25012 (N_25012,N_22246,N_23539);
nand U25013 (N_25013,N_21565,N_23500);
and U25014 (N_25014,N_21176,N_22204);
nor U25015 (N_25015,N_21997,N_22304);
nand U25016 (N_25016,N_22601,N_21071);
nand U25017 (N_25017,N_23952,N_22055);
nor U25018 (N_25018,N_22454,N_21898);
and U25019 (N_25019,N_23312,N_23225);
or U25020 (N_25020,N_21323,N_22531);
or U25021 (N_25021,N_23647,N_22358);
and U25022 (N_25022,N_21977,N_23901);
nor U25023 (N_25023,N_22271,N_22299);
or U25024 (N_25024,N_23749,N_22669);
nand U25025 (N_25025,N_21769,N_23657);
nor U25026 (N_25026,N_22138,N_21157);
xnor U25027 (N_25027,N_22890,N_23885);
and U25028 (N_25028,N_23995,N_21213);
nand U25029 (N_25029,N_22145,N_21343);
nor U25030 (N_25030,N_21723,N_23192);
and U25031 (N_25031,N_23837,N_22348);
xnor U25032 (N_25032,N_23412,N_22613);
or U25033 (N_25033,N_23177,N_22863);
and U25034 (N_25034,N_22590,N_23183);
or U25035 (N_25035,N_22178,N_22500);
and U25036 (N_25036,N_21591,N_23153);
nor U25037 (N_25037,N_23715,N_21121);
xnor U25038 (N_25038,N_22474,N_21524);
xor U25039 (N_25039,N_23087,N_22384);
or U25040 (N_25040,N_23985,N_23054);
and U25041 (N_25041,N_22667,N_22765);
or U25042 (N_25042,N_21392,N_22458);
nand U25043 (N_25043,N_21416,N_23381);
or U25044 (N_25044,N_21218,N_21643);
nor U25045 (N_25045,N_23485,N_22429);
nand U25046 (N_25046,N_22273,N_22014);
and U25047 (N_25047,N_22983,N_22698);
and U25048 (N_25048,N_23821,N_21794);
xor U25049 (N_25049,N_23315,N_21587);
and U25050 (N_25050,N_21258,N_22192);
and U25051 (N_25051,N_21077,N_21154);
or U25052 (N_25052,N_22499,N_22629);
nand U25053 (N_25053,N_22233,N_23553);
nor U25054 (N_25054,N_21584,N_21366);
and U25055 (N_25055,N_22092,N_23116);
xnor U25056 (N_25056,N_22628,N_23660);
nor U25057 (N_25057,N_23387,N_23733);
nand U25058 (N_25058,N_23252,N_23963);
xnor U25059 (N_25059,N_22848,N_21260);
nor U25060 (N_25060,N_23780,N_23577);
or U25061 (N_25061,N_22220,N_22297);
xor U25062 (N_25062,N_22166,N_22544);
and U25063 (N_25063,N_23535,N_22490);
xor U25064 (N_25064,N_23283,N_21180);
or U25065 (N_25065,N_21389,N_22170);
xnor U25066 (N_25066,N_21048,N_23074);
xor U25067 (N_25067,N_21185,N_22041);
nor U25068 (N_25068,N_23961,N_23579);
nand U25069 (N_25069,N_23306,N_22025);
and U25070 (N_25070,N_23284,N_22425);
xnor U25071 (N_25071,N_23384,N_21650);
and U25072 (N_25072,N_22616,N_23050);
or U25073 (N_25073,N_22700,N_22926);
or U25074 (N_25074,N_22228,N_23416);
nand U25075 (N_25075,N_21632,N_21516);
xor U25076 (N_25076,N_21534,N_22675);
and U25077 (N_25077,N_21711,N_21817);
nor U25078 (N_25078,N_21486,N_21032);
nand U25079 (N_25079,N_22943,N_23109);
xor U25080 (N_25080,N_23855,N_22872);
or U25081 (N_25081,N_23772,N_23009);
nand U25082 (N_25082,N_21249,N_22409);
nand U25083 (N_25083,N_21107,N_23088);
and U25084 (N_25084,N_22334,N_23719);
nor U25085 (N_25085,N_21538,N_22261);
or U25086 (N_25086,N_22245,N_21601);
xor U25087 (N_25087,N_21880,N_23357);
nand U25088 (N_25088,N_21722,N_21171);
nor U25089 (N_25089,N_22529,N_21375);
nor U25090 (N_25090,N_22404,N_21611);
or U25091 (N_25091,N_21015,N_22232);
and U25092 (N_25092,N_23209,N_22795);
or U25093 (N_25093,N_21877,N_22760);
xor U25094 (N_25094,N_21956,N_23345);
or U25095 (N_25095,N_23965,N_22520);
xor U25096 (N_25096,N_21452,N_21030);
nor U25097 (N_25097,N_21174,N_21108);
nand U25098 (N_25098,N_22198,N_22897);
or U25099 (N_25099,N_21271,N_21306);
and U25100 (N_25100,N_23141,N_23146);
nor U25101 (N_25101,N_21319,N_22492);
and U25102 (N_25102,N_21494,N_22588);
nand U25103 (N_25103,N_22450,N_21594);
xor U25104 (N_25104,N_22791,N_22653);
nor U25105 (N_25105,N_22298,N_21401);
nor U25106 (N_25106,N_22777,N_23422);
and U25107 (N_25107,N_23407,N_21674);
nor U25108 (N_25108,N_21277,N_23025);
nor U25109 (N_25109,N_22735,N_22341);
nor U25110 (N_25110,N_22307,N_21867);
nand U25111 (N_25111,N_23864,N_23851);
and U25112 (N_25112,N_23364,N_22976);
or U25113 (N_25113,N_22392,N_21055);
or U25114 (N_25114,N_21261,N_23862);
and U25115 (N_25115,N_22792,N_21848);
nor U25116 (N_25116,N_21708,N_21676);
xor U25117 (N_25117,N_21835,N_23664);
nand U25118 (N_25118,N_21812,N_22146);
nand U25119 (N_25119,N_21677,N_21530);
xor U25120 (N_25120,N_22222,N_23643);
and U25121 (N_25121,N_22869,N_22753);
nor U25122 (N_25122,N_22000,N_23805);
nand U25123 (N_25123,N_21144,N_23394);
xor U25124 (N_25124,N_23317,N_21124);
or U25125 (N_25125,N_22208,N_23632);
nand U25126 (N_25126,N_21689,N_21933);
and U25127 (N_25127,N_23763,N_23865);
xor U25128 (N_25128,N_21577,N_21118);
nand U25129 (N_25129,N_22290,N_23269);
xor U25130 (N_25130,N_23972,N_22525);
nor U25131 (N_25131,N_21768,N_21119);
xnor U25132 (N_25132,N_23949,N_23262);
xor U25133 (N_25133,N_23974,N_22416);
nand U25134 (N_25134,N_22734,N_22505);
or U25135 (N_25135,N_21186,N_21765);
nor U25136 (N_25136,N_23292,N_22209);
or U25137 (N_25137,N_22107,N_22473);
nor U25138 (N_25138,N_22142,N_21802);
xor U25139 (N_25139,N_21461,N_21424);
nor U25140 (N_25140,N_21636,N_22502);
and U25141 (N_25141,N_22362,N_23511);
and U25142 (N_25142,N_21431,N_21064);
nor U25143 (N_25143,N_21993,N_23028);
xnor U25144 (N_25144,N_21274,N_23073);
xnor U25145 (N_25145,N_22438,N_23624);
nor U25146 (N_25146,N_23165,N_21245);
nand U25147 (N_25147,N_23710,N_23979);
or U25148 (N_25148,N_21086,N_23894);
and U25149 (N_25149,N_22870,N_23335);
nor U25150 (N_25150,N_22278,N_22240);
nand U25151 (N_25151,N_22563,N_23250);
or U25152 (N_25152,N_22886,N_22542);
nor U25153 (N_25153,N_22457,N_22932);
and U25154 (N_25154,N_22634,N_23188);
and U25155 (N_25155,N_23595,N_23180);
nor U25156 (N_25156,N_22883,N_22119);
nand U25157 (N_25157,N_23718,N_21787);
and U25158 (N_25158,N_22794,N_22548);
xnor U25159 (N_25159,N_22013,N_22780);
nor U25160 (N_25160,N_21989,N_23379);
nand U25161 (N_25161,N_21136,N_21610);
and U25162 (N_25162,N_23740,N_23835);
xnor U25163 (N_25163,N_23679,N_21160);
xnor U25164 (N_25164,N_23474,N_21248);
nand U25165 (N_25165,N_21371,N_21932);
xor U25166 (N_25166,N_23205,N_23888);
and U25167 (N_25167,N_22982,N_21283);
or U25168 (N_25168,N_23163,N_21128);
nor U25169 (N_25169,N_21921,N_22591);
nor U25170 (N_25170,N_22802,N_23032);
and U25171 (N_25171,N_22551,N_23945);
nor U25172 (N_25172,N_22796,N_22822);
and U25173 (N_25173,N_22643,N_23893);
nor U25174 (N_25174,N_21624,N_21502);
and U25175 (N_25175,N_23017,N_23910);
nor U25176 (N_25176,N_22508,N_23690);
nor U25177 (N_25177,N_23279,N_21017);
xor U25178 (N_25178,N_21256,N_22066);
or U25179 (N_25179,N_23704,N_21474);
xnor U25180 (N_25180,N_22077,N_23867);
nor U25181 (N_25181,N_21783,N_22301);
or U25182 (N_25182,N_22071,N_21172);
or U25183 (N_25183,N_21602,N_21949);
xnor U25184 (N_25184,N_23471,N_21362);
nor U25185 (N_25185,N_21204,N_21126);
and U25186 (N_25186,N_23646,N_22018);
or U25187 (N_25187,N_22725,N_21635);
nor U25188 (N_25188,N_22887,N_22332);
and U25189 (N_25189,N_21219,N_21540);
and U25190 (N_25190,N_22002,N_21291);
nand U25191 (N_25191,N_22255,N_22385);
nor U25192 (N_25192,N_22922,N_21523);
xor U25193 (N_25193,N_21328,N_21462);
nor U25194 (N_25194,N_21330,N_23327);
xnor U25195 (N_25195,N_23723,N_23774);
nand U25196 (N_25196,N_22638,N_21680);
nand U25197 (N_25197,N_22370,N_23370);
nand U25198 (N_25198,N_23756,N_22504);
xnor U25199 (N_25199,N_22372,N_23741);
nor U25200 (N_25200,N_21994,N_22256);
nor U25201 (N_25201,N_22560,N_21153);
and U25202 (N_25202,N_21334,N_23937);
nand U25203 (N_25203,N_22081,N_21092);
nand U25204 (N_25204,N_22343,N_21585);
xnor U25205 (N_25205,N_21177,N_22313);
nand U25206 (N_25206,N_21490,N_22738);
xor U25207 (N_25207,N_23462,N_23662);
nand U25208 (N_25208,N_23086,N_22419);
and U25209 (N_25209,N_21175,N_21681);
nand U25210 (N_25210,N_22853,N_23686);
nand U25211 (N_25211,N_23984,N_23593);
or U25212 (N_25212,N_23911,N_23064);
and U25213 (N_25213,N_23798,N_21411);
nand U25214 (N_25214,N_21082,N_23566);
and U25215 (N_25215,N_22672,N_23897);
and U25216 (N_25216,N_22912,N_21818);
nor U25217 (N_25217,N_21238,N_22776);
and U25218 (N_25218,N_22465,N_22648);
xor U25219 (N_25219,N_22421,N_23060);
or U25220 (N_25220,N_21212,N_22349);
nor U25221 (N_25221,N_21548,N_21866);
nand U25222 (N_25222,N_21409,N_21675);
xnor U25223 (N_25223,N_23722,N_23929);
and U25224 (N_25224,N_21742,N_21593);
or U25225 (N_25225,N_23023,N_22173);
nand U25226 (N_25226,N_22523,N_23575);
xnor U25227 (N_25227,N_23866,N_21874);
nor U25228 (N_25228,N_23311,N_23871);
and U25229 (N_25229,N_22064,N_22442);
or U25230 (N_25230,N_23173,N_21265);
nand U25231 (N_25231,N_21059,N_23800);
and U25232 (N_25232,N_23926,N_21449);
nor U25233 (N_25233,N_22856,N_22399);
nand U25234 (N_25234,N_22196,N_23121);
or U25235 (N_25235,N_23224,N_23622);
and U25236 (N_25236,N_23376,N_21934);
nor U25237 (N_25237,N_23773,N_22401);
and U25238 (N_25238,N_22247,N_21988);
nor U25239 (N_25239,N_23860,N_23051);
nor U25240 (N_25240,N_21909,N_22342);
xor U25241 (N_25241,N_22526,N_23442);
nand U25242 (N_25242,N_21518,N_23735);
or U25243 (N_25243,N_21068,N_22439);
and U25244 (N_25244,N_21878,N_21458);
and U25245 (N_25245,N_22254,N_21326);
nor U25246 (N_25246,N_22814,N_21998);
xnor U25247 (N_25247,N_21754,N_22543);
xnor U25248 (N_25248,N_23932,N_22864);
xor U25249 (N_25249,N_22428,N_21010);
nand U25250 (N_25250,N_21719,N_22879);
and U25251 (N_25251,N_22432,N_22771);
nand U25252 (N_25252,N_21324,N_22113);
or U25253 (N_25253,N_22874,N_21667);
nand U25254 (N_25254,N_22573,N_23389);
nand U25255 (N_25255,N_21926,N_22277);
and U25256 (N_25256,N_22843,N_21575);
nand U25257 (N_25257,N_23272,N_21025);
xnor U25258 (N_25258,N_21093,N_23765);
nor U25259 (N_25259,N_21437,N_22539);
nor U25260 (N_25260,N_21295,N_23887);
nor U25261 (N_25261,N_21231,N_21738);
or U25262 (N_25262,N_23135,N_23504);
nor U25263 (N_25263,N_23337,N_22747);
nor U25264 (N_25264,N_21778,N_21772);
xnor U25265 (N_25265,N_23453,N_23856);
nor U25266 (N_25266,N_22008,N_21187);
xor U25267 (N_25267,N_23621,N_22494);
nand U25268 (N_25268,N_22541,N_21652);
nand U25269 (N_25269,N_21066,N_21807);
or U25270 (N_25270,N_22710,N_21051);
nor U25271 (N_25271,N_21730,N_22815);
nand U25272 (N_25272,N_23720,N_23313);
nor U25273 (N_25273,N_21415,N_23056);
or U25274 (N_25274,N_21613,N_21605);
xnor U25275 (N_25275,N_21448,N_22378);
nor U25276 (N_25276,N_22561,N_21862);
nand U25277 (N_25277,N_22180,N_22739);
nand U25278 (N_25278,N_23475,N_22511);
xor U25279 (N_25279,N_22788,N_22754);
nor U25280 (N_25280,N_21510,N_23063);
or U25281 (N_25281,N_22668,N_22485);
xor U25282 (N_25282,N_23803,N_22310);
and U25283 (N_25283,N_22977,N_22827);
nand U25284 (N_25284,N_23976,N_21657);
nor U25285 (N_25285,N_23059,N_22519);
nand U25286 (N_25286,N_22899,N_23371);
or U25287 (N_25287,N_23812,N_23870);
nand U25288 (N_25288,N_23770,N_21377);
xor U25289 (N_25289,N_22743,N_21433);
and U25290 (N_25290,N_23294,N_23179);
or U25291 (N_25291,N_22684,N_22059);
or U25292 (N_25292,N_23854,N_23278);
nor U25293 (N_25293,N_22605,N_21724);
nor U25294 (N_25294,N_23816,N_23811);
nor U25295 (N_25295,N_21834,N_22397);
or U25296 (N_25296,N_23189,N_21340);
or U25297 (N_25297,N_21907,N_22202);
or U25298 (N_25298,N_23066,N_22200);
or U25299 (N_25299,N_22206,N_23656);
and U25300 (N_25300,N_23813,N_21110);
nor U25301 (N_25301,N_21432,N_21749);
and U25302 (N_25302,N_22184,N_21554);
nor U25303 (N_25303,N_21115,N_23714);
nand U25304 (N_25304,N_22692,N_22607);
and U25305 (N_25305,N_23561,N_23459);
xnor U25306 (N_25306,N_22915,N_23024);
nand U25307 (N_25307,N_22069,N_23546);
and U25308 (N_25308,N_22911,N_22455);
xnor U25309 (N_25309,N_23458,N_22640);
nand U25310 (N_25310,N_22112,N_23047);
and U25311 (N_25311,N_23721,N_22665);
xor U25312 (N_25312,N_21031,N_21294);
or U25313 (N_25313,N_23931,N_21428);
or U25314 (N_25314,N_21365,N_21498);
and U25315 (N_25315,N_22961,N_21890);
xnor U25316 (N_25316,N_23775,N_22289);
and U25317 (N_25317,N_22768,N_22691);
or U25318 (N_25318,N_21919,N_23732);
and U25319 (N_25319,N_23547,N_22834);
xnor U25320 (N_25320,N_21928,N_22918);
and U25321 (N_25321,N_22934,N_21826);
nor U25322 (N_25322,N_22496,N_23281);
and U25323 (N_25323,N_23484,N_22470);
xnor U25324 (N_25324,N_22598,N_23046);
xnor U25325 (N_25325,N_21589,N_22140);
nand U25326 (N_25326,N_21269,N_21255);
xnor U25327 (N_25327,N_22956,N_22136);
nand U25328 (N_25328,N_23712,N_22269);
nor U25329 (N_25329,N_21733,N_21044);
and U25330 (N_25330,N_21734,N_21606);
and U25331 (N_25331,N_22172,N_23709);
or U25332 (N_25332,N_22925,N_23781);
or U25333 (N_25333,N_23120,N_21318);
or U25334 (N_25334,N_22168,N_23688);
or U25335 (N_25335,N_22022,N_21957);
xnor U25336 (N_25336,N_22895,N_22116);
nor U25337 (N_25337,N_23037,N_22336);
or U25338 (N_25338,N_21109,N_22888);
or U25339 (N_25339,N_23184,N_21100);
nor U25340 (N_25340,N_22819,N_21251);
nor U25341 (N_25341,N_21489,N_22309);
and U25342 (N_25342,N_22402,N_21799);
xnor U25343 (N_25343,N_22564,N_21651);
nand U25344 (N_25344,N_22135,N_21482);
xor U25345 (N_25345,N_21945,N_23221);
nand U25346 (N_25346,N_23476,N_23031);
xnor U25347 (N_25347,N_23148,N_21519);
xor U25348 (N_25348,N_21427,N_22737);
or U25349 (N_25349,N_22477,N_23151);
xor U25350 (N_25350,N_22407,N_22720);
nand U25351 (N_25351,N_22472,N_21872);
xor U25352 (N_25352,N_22769,N_23287);
and U25353 (N_25353,N_22461,N_21057);
nor U25354 (N_25354,N_22859,N_22999);
or U25355 (N_25355,N_22775,N_23261);
xnor U25356 (N_25356,N_22844,N_23987);
xnor U25357 (N_25357,N_21786,N_23240);
or U25358 (N_25358,N_22395,N_23755);
nand U25359 (N_25359,N_21824,N_22901);
or U25360 (N_25360,N_23127,N_21889);
nor U25361 (N_25361,N_21808,N_21333);
or U25362 (N_25362,N_21975,N_22589);
xor U25363 (N_25363,N_23229,N_23483);
or U25364 (N_25364,N_22248,N_23020);
xnor U25365 (N_25365,N_22331,N_21438);
nand U25366 (N_25366,N_22510,N_22670);
nor U25367 (N_25367,N_21766,N_23771);
nand U25368 (N_25368,N_22581,N_21043);
nand U25369 (N_25369,N_22125,N_21579);
nand U25370 (N_25370,N_23182,N_21619);
xor U25371 (N_25371,N_21426,N_21620);
nor U25372 (N_25372,N_22964,N_23759);
or U25373 (N_25373,N_22708,N_23728);
or U25374 (N_25374,N_23456,N_23140);
nand U25375 (N_25375,N_23918,N_22865);
or U25376 (N_25376,N_23923,N_21838);
or U25377 (N_25377,N_21948,N_23175);
nand U25378 (N_25378,N_22552,N_22674);
nand U25379 (N_25379,N_21067,N_21446);
xnor U25380 (N_25380,N_22479,N_23463);
nand U25381 (N_25381,N_22847,N_23196);
and U25382 (N_25382,N_21425,N_22446);
nand U25383 (N_25383,N_23129,N_22905);
or U25384 (N_25384,N_22021,N_21314);
nand U25385 (N_25385,N_22101,N_23567);
or U25386 (N_25386,N_21627,N_23280);
and U25387 (N_25387,N_23300,N_22436);
nor U25388 (N_25388,N_21181,N_22268);
xor U25389 (N_25389,N_21968,N_22293);
and U25390 (N_25390,N_21985,N_22082);
nor U25391 (N_25391,N_22115,N_22124);
nand U25392 (N_25392,N_23876,N_22831);
nand U25393 (N_25393,N_22986,N_21582);
nand U25394 (N_25394,N_21672,N_21886);
or U25395 (N_25395,N_23035,N_22969);
nor U25396 (N_25396,N_22075,N_21751);
nand U25397 (N_25397,N_21875,N_21894);
and U25398 (N_25398,N_22345,N_22067);
and U25399 (N_25399,N_22408,N_22807);
and U25400 (N_25400,N_21712,N_22213);
nand U25401 (N_25401,N_21529,N_22952);
and U25402 (N_25402,N_21282,N_23400);
nand U25403 (N_25403,N_22369,N_22610);
nand U25404 (N_25404,N_21355,N_21592);
and U25405 (N_25405,N_23843,N_22876);
nor U25406 (N_25406,N_22199,N_21106);
and U25407 (N_25407,N_21705,N_21164);
and U25408 (N_25408,N_21731,N_23512);
or U25409 (N_25409,N_22786,N_23301);
and U25410 (N_25410,N_21535,N_23352);
nand U25411 (N_25411,N_21379,N_22143);
or U25412 (N_25412,N_23380,N_22750);
or U25413 (N_25413,N_22351,N_23528);
and U25414 (N_25414,N_23369,N_23256);
xor U25415 (N_25415,N_21222,N_22752);
and U25416 (N_25416,N_22690,N_21327);
and U25417 (N_25417,N_23195,N_21287);
xnor U25418 (N_25418,N_22237,N_22090);
nand U25419 (N_25419,N_21964,N_21757);
nand U25420 (N_25420,N_23044,N_22447);
and U25421 (N_25421,N_22524,N_21072);
or U25422 (N_25422,N_23277,N_22363);
and U25423 (N_25423,N_23902,N_23516);
nor U25424 (N_25424,N_21662,N_22650);
or U25425 (N_25425,N_22706,N_21729);
or U25426 (N_25426,N_23021,N_22126);
or U25427 (N_25427,N_22767,N_22078);
nand U25428 (N_25428,N_21697,N_22916);
nand U25429 (N_25429,N_22039,N_22626);
or U25430 (N_25430,N_21233,N_22731);
xnor U25431 (N_25431,N_21912,N_23131);
xnor U25432 (N_25432,N_23226,N_23958);
or U25433 (N_25433,N_21361,N_21155);
nand U25434 (N_25434,N_23872,N_23464);
and U25435 (N_25435,N_21937,N_21062);
xor U25436 (N_25436,N_21773,N_22333);
nand U25437 (N_25437,N_23443,N_22515);
nor U25438 (N_25438,N_23971,N_21041);
or U25439 (N_25439,N_21414,N_22211);
and U25440 (N_25440,N_23635,N_21704);
xnor U25441 (N_25441,N_23981,N_22480);
xor U25442 (N_25442,N_23738,N_22139);
xnor U25443 (N_25443,N_22862,N_22040);
or U25444 (N_25444,N_23080,N_22715);
nand U25445 (N_25445,N_23783,N_22503);
xnor U25446 (N_25446,N_21598,N_22942);
and U25447 (N_25447,N_22637,N_23015);
xnor U25448 (N_25448,N_21056,N_21145);
and U25449 (N_25449,N_21641,N_23228);
nor U25450 (N_25450,N_22944,N_21842);
nor U25451 (N_25451,N_23692,N_21342);
nor U25452 (N_25452,N_22577,N_22965);
or U25453 (N_25453,N_22683,N_21859);
nand U25454 (N_25454,N_23936,N_23637);
xnor U25455 (N_25455,N_21755,N_21042);
or U25456 (N_25456,N_21785,N_23045);
and U25457 (N_25457,N_21560,N_23489);
or U25458 (N_25458,N_21395,N_22227);
or U25459 (N_25459,N_23329,N_23382);
nand U25460 (N_25460,N_21293,N_22512);
xnor U25461 (N_25461,N_23068,N_22051);
nor U25462 (N_25462,N_21963,N_21351);
xor U25463 (N_25463,N_23323,N_23403);
and U25464 (N_25464,N_22194,N_22721);
or U25465 (N_25465,N_21381,N_21135);
nor U25466 (N_25466,N_23130,N_22086);
or U25467 (N_25467,N_21860,N_22487);
or U25468 (N_25468,N_23339,N_23836);
nand U25469 (N_25469,N_21122,N_21971);
nor U25470 (N_25470,N_21782,N_21764);
nor U25471 (N_25471,N_22110,N_22294);
xnor U25472 (N_25472,N_23869,N_22955);
nand U25473 (N_25473,N_23437,N_23134);
or U25474 (N_25474,N_23879,N_23795);
nor U25475 (N_25475,N_23098,N_22076);
and U25476 (N_25476,N_21692,N_21895);
or U25477 (N_25477,N_21036,N_21191);
nand U25478 (N_25478,N_22898,N_22694);
xnor U25479 (N_25479,N_21194,N_23975);
nor U25480 (N_25480,N_23642,N_21809);
and U25481 (N_25481,N_21720,N_21023);
nand U25482 (N_25482,N_22053,N_22608);
nor U25483 (N_25483,N_22433,N_21943);
xnor U25484 (N_25484,N_22444,N_23565);
xor U25485 (N_25485,N_21305,N_23408);
nor U25486 (N_25486,N_23620,N_21440);
nor U25487 (N_25487,N_22016,N_23640);
or U25488 (N_25488,N_23402,N_21979);
and U25489 (N_25489,N_21075,N_22620);
nor U25490 (N_25490,N_22167,N_21980);
and U25491 (N_25491,N_21472,N_23438);
nor U25492 (N_25492,N_23057,N_23111);
or U25493 (N_25493,N_22550,N_21910);
or U25494 (N_25494,N_23731,N_21576);
and U25495 (N_25495,N_23386,N_23631);
xor U25496 (N_25496,N_23355,N_23334);
nand U25497 (N_25497,N_22398,N_22324);
or U25498 (N_25498,N_21951,N_21777);
or U25499 (N_25499,N_22155,N_22024);
or U25500 (N_25500,N_23030,N_22412);
or U25501 (N_25501,N_23623,N_23412);
nor U25502 (N_25502,N_22799,N_22822);
nor U25503 (N_25503,N_21037,N_22559);
xnor U25504 (N_25504,N_21357,N_22980);
or U25505 (N_25505,N_22775,N_22262);
and U25506 (N_25506,N_21425,N_21371);
nand U25507 (N_25507,N_22799,N_23003);
and U25508 (N_25508,N_23859,N_21760);
or U25509 (N_25509,N_21184,N_23915);
xnor U25510 (N_25510,N_22996,N_23071);
nand U25511 (N_25511,N_23558,N_23832);
nor U25512 (N_25512,N_21213,N_23412);
nand U25513 (N_25513,N_21108,N_21379);
nand U25514 (N_25514,N_22343,N_21832);
nor U25515 (N_25515,N_23856,N_21605);
and U25516 (N_25516,N_21136,N_22496);
xnor U25517 (N_25517,N_23533,N_22043);
or U25518 (N_25518,N_21816,N_21527);
and U25519 (N_25519,N_21287,N_23975);
nor U25520 (N_25520,N_23522,N_21144);
xor U25521 (N_25521,N_22029,N_22109);
nor U25522 (N_25522,N_22986,N_21722);
or U25523 (N_25523,N_21473,N_21143);
and U25524 (N_25524,N_23136,N_22547);
xnor U25525 (N_25525,N_21717,N_22941);
or U25526 (N_25526,N_22401,N_22958);
nand U25527 (N_25527,N_21830,N_22215);
or U25528 (N_25528,N_23330,N_23991);
nor U25529 (N_25529,N_21636,N_21975);
xnor U25530 (N_25530,N_21430,N_23005);
xor U25531 (N_25531,N_21134,N_21076);
or U25532 (N_25532,N_23338,N_21845);
nor U25533 (N_25533,N_21479,N_23045);
and U25534 (N_25534,N_22956,N_23574);
nor U25535 (N_25535,N_23575,N_23918);
or U25536 (N_25536,N_22439,N_22554);
and U25537 (N_25537,N_23218,N_22409);
and U25538 (N_25538,N_22871,N_21988);
and U25539 (N_25539,N_21245,N_23556);
nor U25540 (N_25540,N_21890,N_23434);
xor U25541 (N_25541,N_21242,N_21021);
xnor U25542 (N_25542,N_21299,N_21531);
nand U25543 (N_25543,N_22728,N_21511);
xor U25544 (N_25544,N_21623,N_23330);
and U25545 (N_25545,N_21743,N_21672);
xnor U25546 (N_25546,N_21392,N_21849);
nor U25547 (N_25547,N_22366,N_23075);
nor U25548 (N_25548,N_23659,N_22461);
xnor U25549 (N_25549,N_22367,N_22978);
xnor U25550 (N_25550,N_22418,N_23372);
or U25551 (N_25551,N_22263,N_22005);
xnor U25552 (N_25552,N_23599,N_21294);
xor U25553 (N_25553,N_23910,N_21386);
nand U25554 (N_25554,N_23437,N_22879);
nand U25555 (N_25555,N_21391,N_23859);
or U25556 (N_25556,N_22006,N_23138);
nor U25557 (N_25557,N_21658,N_23004);
nand U25558 (N_25558,N_23040,N_21007);
nand U25559 (N_25559,N_22480,N_21465);
xor U25560 (N_25560,N_22000,N_21651);
and U25561 (N_25561,N_21309,N_23450);
nor U25562 (N_25562,N_23006,N_23494);
nand U25563 (N_25563,N_23368,N_21128);
nor U25564 (N_25564,N_23439,N_22304);
or U25565 (N_25565,N_21793,N_23250);
and U25566 (N_25566,N_22873,N_23399);
nor U25567 (N_25567,N_23016,N_23200);
nor U25568 (N_25568,N_22198,N_21389);
nor U25569 (N_25569,N_22414,N_21558);
or U25570 (N_25570,N_23989,N_21004);
xor U25571 (N_25571,N_22877,N_22875);
xor U25572 (N_25572,N_23058,N_22081);
nand U25573 (N_25573,N_23463,N_22560);
or U25574 (N_25574,N_21915,N_22150);
and U25575 (N_25575,N_21398,N_23533);
xor U25576 (N_25576,N_22539,N_21671);
and U25577 (N_25577,N_23718,N_23072);
xor U25578 (N_25578,N_21886,N_22222);
nor U25579 (N_25579,N_22598,N_23506);
nor U25580 (N_25580,N_21338,N_22609);
nor U25581 (N_25581,N_23292,N_21888);
nand U25582 (N_25582,N_22966,N_21866);
xnor U25583 (N_25583,N_21574,N_21505);
or U25584 (N_25584,N_21681,N_22831);
or U25585 (N_25585,N_22023,N_21694);
or U25586 (N_25586,N_23695,N_22762);
or U25587 (N_25587,N_22373,N_21868);
and U25588 (N_25588,N_21929,N_23527);
xnor U25589 (N_25589,N_22797,N_21665);
nand U25590 (N_25590,N_22459,N_21894);
nand U25591 (N_25591,N_23274,N_21969);
nor U25592 (N_25592,N_22009,N_21015);
xnor U25593 (N_25593,N_23414,N_21438);
nor U25594 (N_25594,N_23055,N_23381);
or U25595 (N_25595,N_21889,N_22101);
nand U25596 (N_25596,N_23624,N_21526);
xnor U25597 (N_25597,N_22613,N_21406);
xnor U25598 (N_25598,N_21153,N_21494);
nor U25599 (N_25599,N_23610,N_21413);
nand U25600 (N_25600,N_22115,N_21123);
or U25601 (N_25601,N_21235,N_23257);
and U25602 (N_25602,N_22036,N_21175);
nand U25603 (N_25603,N_23459,N_22176);
nand U25604 (N_25604,N_22453,N_22449);
nor U25605 (N_25605,N_23496,N_22999);
nand U25606 (N_25606,N_21888,N_21929);
xnor U25607 (N_25607,N_21786,N_23688);
or U25608 (N_25608,N_22961,N_21474);
nor U25609 (N_25609,N_21204,N_22250);
nor U25610 (N_25610,N_23956,N_21541);
and U25611 (N_25611,N_22903,N_23105);
and U25612 (N_25612,N_21244,N_23203);
xnor U25613 (N_25613,N_21280,N_23208);
xnor U25614 (N_25614,N_23485,N_21917);
nor U25615 (N_25615,N_23130,N_22982);
nand U25616 (N_25616,N_22854,N_23542);
nand U25617 (N_25617,N_23976,N_21986);
nand U25618 (N_25618,N_21865,N_21771);
nor U25619 (N_25619,N_23909,N_22135);
or U25620 (N_25620,N_22850,N_23316);
xor U25621 (N_25621,N_21749,N_22936);
xnor U25622 (N_25622,N_21748,N_22596);
xnor U25623 (N_25623,N_21422,N_23994);
nand U25624 (N_25624,N_22281,N_21431);
nor U25625 (N_25625,N_21843,N_22510);
and U25626 (N_25626,N_23077,N_22341);
nand U25627 (N_25627,N_22641,N_21317);
xnor U25628 (N_25628,N_23964,N_22215);
nor U25629 (N_25629,N_21000,N_22972);
nor U25630 (N_25630,N_23457,N_23020);
nand U25631 (N_25631,N_23237,N_21800);
and U25632 (N_25632,N_23164,N_23079);
or U25633 (N_25633,N_23126,N_23284);
nand U25634 (N_25634,N_21657,N_22963);
nand U25635 (N_25635,N_23118,N_21602);
and U25636 (N_25636,N_21255,N_23187);
nand U25637 (N_25637,N_23772,N_22009);
nand U25638 (N_25638,N_22985,N_21072);
nor U25639 (N_25639,N_21075,N_22932);
xor U25640 (N_25640,N_22743,N_23482);
or U25641 (N_25641,N_23193,N_21885);
nor U25642 (N_25642,N_23538,N_21884);
xnor U25643 (N_25643,N_22673,N_22386);
nor U25644 (N_25644,N_23604,N_23774);
nor U25645 (N_25645,N_22901,N_21992);
nor U25646 (N_25646,N_21556,N_23139);
nand U25647 (N_25647,N_21537,N_23977);
and U25648 (N_25648,N_22663,N_23598);
or U25649 (N_25649,N_21918,N_21752);
xnor U25650 (N_25650,N_23779,N_23794);
xor U25651 (N_25651,N_21183,N_22155);
and U25652 (N_25652,N_23024,N_22266);
nor U25653 (N_25653,N_23757,N_21454);
and U25654 (N_25654,N_21052,N_22639);
nand U25655 (N_25655,N_23440,N_22440);
nor U25656 (N_25656,N_22957,N_21854);
nor U25657 (N_25657,N_22247,N_23840);
or U25658 (N_25658,N_23063,N_23516);
nand U25659 (N_25659,N_22611,N_22897);
nand U25660 (N_25660,N_21228,N_23739);
nand U25661 (N_25661,N_22930,N_21373);
or U25662 (N_25662,N_23850,N_22071);
and U25663 (N_25663,N_23005,N_22173);
or U25664 (N_25664,N_22146,N_21212);
xnor U25665 (N_25665,N_23498,N_22980);
nand U25666 (N_25666,N_21052,N_22416);
nand U25667 (N_25667,N_22515,N_23807);
nand U25668 (N_25668,N_21904,N_22922);
nor U25669 (N_25669,N_21724,N_22294);
nand U25670 (N_25670,N_22347,N_23400);
nor U25671 (N_25671,N_22487,N_21631);
nand U25672 (N_25672,N_21536,N_22363);
xor U25673 (N_25673,N_21061,N_22626);
nand U25674 (N_25674,N_22541,N_22130);
nor U25675 (N_25675,N_21445,N_23473);
nand U25676 (N_25676,N_23515,N_22843);
and U25677 (N_25677,N_21552,N_22784);
or U25678 (N_25678,N_23506,N_22790);
nand U25679 (N_25679,N_22730,N_23070);
xor U25680 (N_25680,N_23813,N_21816);
nand U25681 (N_25681,N_21428,N_22206);
or U25682 (N_25682,N_22596,N_22491);
nor U25683 (N_25683,N_23813,N_23885);
and U25684 (N_25684,N_22399,N_23170);
and U25685 (N_25685,N_23885,N_23881);
or U25686 (N_25686,N_21441,N_22912);
xnor U25687 (N_25687,N_23909,N_23106);
nor U25688 (N_25688,N_21429,N_23625);
and U25689 (N_25689,N_22253,N_23551);
xor U25690 (N_25690,N_21364,N_21644);
nand U25691 (N_25691,N_21856,N_21639);
xor U25692 (N_25692,N_23056,N_22526);
nor U25693 (N_25693,N_21098,N_21947);
and U25694 (N_25694,N_21661,N_21972);
nand U25695 (N_25695,N_23713,N_22071);
xor U25696 (N_25696,N_21895,N_21035);
xor U25697 (N_25697,N_22762,N_21945);
and U25698 (N_25698,N_22008,N_21415);
nand U25699 (N_25699,N_21964,N_22721);
and U25700 (N_25700,N_23263,N_21169);
or U25701 (N_25701,N_23705,N_21005);
xor U25702 (N_25702,N_21489,N_21769);
nand U25703 (N_25703,N_22227,N_22898);
and U25704 (N_25704,N_23253,N_23942);
nand U25705 (N_25705,N_22289,N_22142);
nand U25706 (N_25706,N_22186,N_22365);
or U25707 (N_25707,N_21146,N_22471);
xor U25708 (N_25708,N_22972,N_23123);
and U25709 (N_25709,N_22744,N_21244);
nor U25710 (N_25710,N_23728,N_22162);
and U25711 (N_25711,N_22563,N_21002);
nand U25712 (N_25712,N_22057,N_21010);
or U25713 (N_25713,N_23515,N_21253);
and U25714 (N_25714,N_22015,N_23787);
and U25715 (N_25715,N_22547,N_23537);
or U25716 (N_25716,N_23925,N_23212);
or U25717 (N_25717,N_23787,N_22278);
and U25718 (N_25718,N_22494,N_21515);
or U25719 (N_25719,N_23265,N_23132);
and U25720 (N_25720,N_21252,N_23174);
and U25721 (N_25721,N_21339,N_21743);
xor U25722 (N_25722,N_23211,N_22468);
nor U25723 (N_25723,N_23353,N_21603);
or U25724 (N_25724,N_23616,N_22534);
nand U25725 (N_25725,N_21497,N_21449);
xor U25726 (N_25726,N_23824,N_21527);
or U25727 (N_25727,N_21780,N_22195);
and U25728 (N_25728,N_21680,N_23096);
nor U25729 (N_25729,N_21104,N_23132);
and U25730 (N_25730,N_22674,N_22560);
or U25731 (N_25731,N_23794,N_22239);
xnor U25732 (N_25732,N_23355,N_21874);
and U25733 (N_25733,N_23319,N_23751);
and U25734 (N_25734,N_22426,N_22475);
xnor U25735 (N_25735,N_22428,N_21158);
nor U25736 (N_25736,N_21230,N_22672);
nand U25737 (N_25737,N_23213,N_21359);
and U25738 (N_25738,N_21381,N_21588);
nand U25739 (N_25739,N_23525,N_22099);
and U25740 (N_25740,N_21223,N_23320);
and U25741 (N_25741,N_23011,N_22775);
nand U25742 (N_25742,N_23574,N_23011);
xor U25743 (N_25743,N_21435,N_21420);
xnor U25744 (N_25744,N_21004,N_23430);
or U25745 (N_25745,N_23667,N_23706);
xnor U25746 (N_25746,N_21446,N_23127);
nand U25747 (N_25747,N_22264,N_23905);
and U25748 (N_25748,N_21248,N_21134);
nor U25749 (N_25749,N_21152,N_21927);
and U25750 (N_25750,N_23387,N_23765);
xor U25751 (N_25751,N_23678,N_23858);
or U25752 (N_25752,N_22659,N_21388);
and U25753 (N_25753,N_23903,N_21718);
and U25754 (N_25754,N_23738,N_22770);
or U25755 (N_25755,N_22372,N_23544);
nand U25756 (N_25756,N_22474,N_21526);
nand U25757 (N_25757,N_21218,N_21973);
nor U25758 (N_25758,N_21535,N_22643);
and U25759 (N_25759,N_22833,N_23626);
nor U25760 (N_25760,N_23688,N_21268);
xor U25761 (N_25761,N_22892,N_21029);
xor U25762 (N_25762,N_22064,N_21173);
nand U25763 (N_25763,N_21164,N_23201);
xnor U25764 (N_25764,N_21028,N_22695);
nand U25765 (N_25765,N_23264,N_21604);
and U25766 (N_25766,N_22763,N_21035);
nor U25767 (N_25767,N_23035,N_21362);
or U25768 (N_25768,N_23026,N_23437);
xnor U25769 (N_25769,N_22511,N_21328);
nand U25770 (N_25770,N_23788,N_23641);
nor U25771 (N_25771,N_21202,N_21611);
nor U25772 (N_25772,N_22283,N_21677);
nand U25773 (N_25773,N_23553,N_22440);
and U25774 (N_25774,N_22369,N_22818);
or U25775 (N_25775,N_23212,N_23886);
nor U25776 (N_25776,N_21072,N_23003);
nand U25777 (N_25777,N_22418,N_21567);
nor U25778 (N_25778,N_23184,N_22346);
or U25779 (N_25779,N_23362,N_22454);
or U25780 (N_25780,N_22886,N_23135);
and U25781 (N_25781,N_21792,N_22637);
xor U25782 (N_25782,N_21893,N_23220);
nor U25783 (N_25783,N_21407,N_23430);
or U25784 (N_25784,N_23271,N_22287);
nand U25785 (N_25785,N_21710,N_23922);
nand U25786 (N_25786,N_22187,N_22983);
nand U25787 (N_25787,N_22556,N_23851);
nor U25788 (N_25788,N_23889,N_22151);
nand U25789 (N_25789,N_21436,N_23401);
nand U25790 (N_25790,N_23053,N_22615);
or U25791 (N_25791,N_22525,N_21615);
nand U25792 (N_25792,N_23923,N_23703);
or U25793 (N_25793,N_22825,N_22559);
nand U25794 (N_25794,N_21627,N_21935);
nor U25795 (N_25795,N_21633,N_22986);
nor U25796 (N_25796,N_21605,N_22219);
nand U25797 (N_25797,N_23858,N_22302);
nor U25798 (N_25798,N_21393,N_22409);
nor U25799 (N_25799,N_21695,N_22755);
nand U25800 (N_25800,N_23731,N_21406);
xnor U25801 (N_25801,N_21497,N_21269);
nor U25802 (N_25802,N_21639,N_21183);
and U25803 (N_25803,N_21535,N_22901);
xor U25804 (N_25804,N_23733,N_23047);
or U25805 (N_25805,N_23890,N_21396);
nand U25806 (N_25806,N_22153,N_22314);
nor U25807 (N_25807,N_23567,N_22582);
nor U25808 (N_25808,N_21359,N_21865);
xor U25809 (N_25809,N_21809,N_22180);
nand U25810 (N_25810,N_22897,N_22675);
xnor U25811 (N_25811,N_21573,N_22787);
nor U25812 (N_25812,N_23890,N_22240);
nand U25813 (N_25813,N_23220,N_23377);
or U25814 (N_25814,N_22206,N_22936);
or U25815 (N_25815,N_22669,N_21743);
nor U25816 (N_25816,N_23672,N_22590);
nand U25817 (N_25817,N_22546,N_22309);
or U25818 (N_25818,N_21181,N_22194);
nand U25819 (N_25819,N_22534,N_22579);
and U25820 (N_25820,N_22692,N_21514);
xnor U25821 (N_25821,N_23662,N_23513);
and U25822 (N_25822,N_21074,N_22819);
nand U25823 (N_25823,N_23104,N_21266);
nand U25824 (N_25824,N_21509,N_22959);
nand U25825 (N_25825,N_22815,N_22642);
xor U25826 (N_25826,N_22044,N_21295);
nor U25827 (N_25827,N_21927,N_23909);
or U25828 (N_25828,N_23096,N_21519);
nor U25829 (N_25829,N_23606,N_22478);
nor U25830 (N_25830,N_23896,N_22211);
or U25831 (N_25831,N_21002,N_21991);
xor U25832 (N_25832,N_22799,N_23979);
nand U25833 (N_25833,N_21548,N_22311);
xor U25834 (N_25834,N_21695,N_21563);
nand U25835 (N_25835,N_21903,N_21825);
or U25836 (N_25836,N_21791,N_23497);
or U25837 (N_25837,N_23764,N_21618);
or U25838 (N_25838,N_21396,N_21103);
or U25839 (N_25839,N_21404,N_21141);
nand U25840 (N_25840,N_23005,N_22328);
and U25841 (N_25841,N_21867,N_21921);
nand U25842 (N_25842,N_22132,N_22713);
nor U25843 (N_25843,N_21620,N_23894);
and U25844 (N_25844,N_22917,N_23454);
and U25845 (N_25845,N_21931,N_23101);
or U25846 (N_25846,N_21652,N_21561);
nand U25847 (N_25847,N_21124,N_21863);
nand U25848 (N_25848,N_23355,N_23785);
nor U25849 (N_25849,N_22322,N_22000);
xnor U25850 (N_25850,N_22047,N_23092);
xnor U25851 (N_25851,N_23088,N_22157);
or U25852 (N_25852,N_21103,N_21748);
nor U25853 (N_25853,N_22726,N_23807);
and U25854 (N_25854,N_23879,N_23218);
and U25855 (N_25855,N_21021,N_21933);
xor U25856 (N_25856,N_22660,N_22761);
and U25857 (N_25857,N_23768,N_21771);
nand U25858 (N_25858,N_21255,N_23345);
xnor U25859 (N_25859,N_22872,N_21067);
xnor U25860 (N_25860,N_21627,N_22429);
nor U25861 (N_25861,N_21326,N_22164);
and U25862 (N_25862,N_23298,N_21540);
xor U25863 (N_25863,N_21774,N_21335);
and U25864 (N_25864,N_22170,N_23469);
nand U25865 (N_25865,N_22323,N_22382);
nor U25866 (N_25866,N_23396,N_21450);
nor U25867 (N_25867,N_22215,N_21882);
nand U25868 (N_25868,N_21372,N_23869);
and U25869 (N_25869,N_21902,N_23425);
or U25870 (N_25870,N_23422,N_21633);
nand U25871 (N_25871,N_23761,N_21231);
nand U25872 (N_25872,N_23549,N_23291);
and U25873 (N_25873,N_23679,N_23123);
xor U25874 (N_25874,N_23251,N_23245);
and U25875 (N_25875,N_21106,N_23006);
or U25876 (N_25876,N_21390,N_23048);
and U25877 (N_25877,N_22459,N_21706);
and U25878 (N_25878,N_22562,N_21628);
nor U25879 (N_25879,N_21918,N_23501);
xor U25880 (N_25880,N_22042,N_23872);
and U25881 (N_25881,N_22525,N_22398);
or U25882 (N_25882,N_21286,N_21220);
or U25883 (N_25883,N_22102,N_22466);
nand U25884 (N_25884,N_22142,N_21477);
and U25885 (N_25885,N_23393,N_23823);
nand U25886 (N_25886,N_22037,N_22865);
xnor U25887 (N_25887,N_23253,N_22601);
nor U25888 (N_25888,N_22134,N_21153);
and U25889 (N_25889,N_22523,N_23731);
nor U25890 (N_25890,N_22679,N_21548);
nor U25891 (N_25891,N_22911,N_23208);
and U25892 (N_25892,N_21980,N_21505);
nor U25893 (N_25893,N_22641,N_22832);
xor U25894 (N_25894,N_23798,N_22204);
nor U25895 (N_25895,N_21907,N_22342);
xor U25896 (N_25896,N_23459,N_21432);
nand U25897 (N_25897,N_21238,N_21185);
and U25898 (N_25898,N_21295,N_22897);
nor U25899 (N_25899,N_21993,N_22858);
or U25900 (N_25900,N_21906,N_21680);
nor U25901 (N_25901,N_23251,N_21634);
and U25902 (N_25902,N_22639,N_22654);
and U25903 (N_25903,N_21562,N_23403);
nand U25904 (N_25904,N_23991,N_22174);
nor U25905 (N_25905,N_21174,N_23175);
xor U25906 (N_25906,N_21468,N_23787);
or U25907 (N_25907,N_23381,N_22540);
nand U25908 (N_25908,N_22489,N_21066);
and U25909 (N_25909,N_22962,N_22600);
nor U25910 (N_25910,N_22255,N_22303);
xor U25911 (N_25911,N_21501,N_23202);
or U25912 (N_25912,N_21671,N_23973);
or U25913 (N_25913,N_22125,N_22680);
and U25914 (N_25914,N_21060,N_21265);
nand U25915 (N_25915,N_21885,N_21249);
nand U25916 (N_25916,N_23624,N_23191);
or U25917 (N_25917,N_21859,N_23142);
and U25918 (N_25918,N_23947,N_21390);
and U25919 (N_25919,N_23023,N_22274);
nand U25920 (N_25920,N_23416,N_22476);
and U25921 (N_25921,N_23254,N_21454);
or U25922 (N_25922,N_21494,N_22434);
nand U25923 (N_25923,N_21975,N_22167);
or U25924 (N_25924,N_21801,N_21297);
or U25925 (N_25925,N_23846,N_23694);
nor U25926 (N_25926,N_21420,N_21362);
nor U25927 (N_25927,N_21154,N_23236);
nand U25928 (N_25928,N_21659,N_21988);
xor U25929 (N_25929,N_21471,N_22577);
xor U25930 (N_25930,N_23920,N_22027);
or U25931 (N_25931,N_23771,N_23296);
and U25932 (N_25932,N_22995,N_23421);
xnor U25933 (N_25933,N_22003,N_23434);
nor U25934 (N_25934,N_22935,N_23659);
nand U25935 (N_25935,N_22871,N_23090);
nand U25936 (N_25936,N_21340,N_23116);
or U25937 (N_25937,N_21547,N_21629);
nor U25938 (N_25938,N_21574,N_23114);
nor U25939 (N_25939,N_21988,N_23045);
and U25940 (N_25940,N_23811,N_22940);
xnor U25941 (N_25941,N_23808,N_21852);
and U25942 (N_25942,N_23646,N_21176);
nor U25943 (N_25943,N_22858,N_21862);
and U25944 (N_25944,N_23370,N_23854);
nand U25945 (N_25945,N_22408,N_22373);
nor U25946 (N_25946,N_23268,N_21899);
and U25947 (N_25947,N_21037,N_21341);
or U25948 (N_25948,N_21973,N_22548);
xor U25949 (N_25949,N_23491,N_21105);
and U25950 (N_25950,N_21098,N_23718);
nor U25951 (N_25951,N_22074,N_21002);
and U25952 (N_25952,N_23800,N_23671);
or U25953 (N_25953,N_23260,N_22880);
and U25954 (N_25954,N_22775,N_21874);
and U25955 (N_25955,N_23561,N_21804);
xnor U25956 (N_25956,N_22268,N_21905);
nand U25957 (N_25957,N_21990,N_21434);
or U25958 (N_25958,N_21302,N_21721);
nor U25959 (N_25959,N_23525,N_23976);
nand U25960 (N_25960,N_23463,N_23917);
and U25961 (N_25961,N_22873,N_22701);
and U25962 (N_25962,N_22313,N_21269);
nand U25963 (N_25963,N_22474,N_21623);
nand U25964 (N_25964,N_22343,N_21812);
and U25965 (N_25965,N_23144,N_23320);
nor U25966 (N_25966,N_21038,N_22089);
and U25967 (N_25967,N_21309,N_23279);
or U25968 (N_25968,N_21248,N_21301);
nand U25969 (N_25969,N_22955,N_22573);
and U25970 (N_25970,N_21269,N_22684);
nor U25971 (N_25971,N_21118,N_22886);
nor U25972 (N_25972,N_21851,N_21923);
xnor U25973 (N_25973,N_21452,N_23159);
and U25974 (N_25974,N_22097,N_22128);
nand U25975 (N_25975,N_23432,N_23772);
and U25976 (N_25976,N_23656,N_22302);
nand U25977 (N_25977,N_21886,N_23967);
nand U25978 (N_25978,N_22954,N_23786);
or U25979 (N_25979,N_22442,N_22960);
and U25980 (N_25980,N_23152,N_21655);
xnor U25981 (N_25981,N_21406,N_21711);
and U25982 (N_25982,N_23138,N_23387);
nand U25983 (N_25983,N_21834,N_23476);
or U25984 (N_25984,N_21462,N_23655);
or U25985 (N_25985,N_23025,N_23044);
xnor U25986 (N_25986,N_22956,N_21676);
nand U25987 (N_25987,N_23219,N_22829);
nand U25988 (N_25988,N_22720,N_22787);
or U25989 (N_25989,N_22124,N_23339);
or U25990 (N_25990,N_23544,N_22308);
xor U25991 (N_25991,N_22558,N_21504);
or U25992 (N_25992,N_23715,N_22964);
nand U25993 (N_25993,N_22647,N_21230);
xor U25994 (N_25994,N_22681,N_22041);
xnor U25995 (N_25995,N_21798,N_23716);
nor U25996 (N_25996,N_22098,N_21851);
nand U25997 (N_25997,N_23993,N_23517);
nor U25998 (N_25998,N_21152,N_22300);
nand U25999 (N_25999,N_22057,N_21065);
and U26000 (N_26000,N_23674,N_21628);
and U26001 (N_26001,N_22108,N_22153);
nor U26002 (N_26002,N_21895,N_23241);
or U26003 (N_26003,N_21192,N_22084);
xnor U26004 (N_26004,N_23416,N_22379);
xor U26005 (N_26005,N_21235,N_21838);
and U26006 (N_26006,N_21664,N_23464);
nor U26007 (N_26007,N_22474,N_21118);
xor U26008 (N_26008,N_23619,N_22404);
xnor U26009 (N_26009,N_21491,N_22095);
xnor U26010 (N_26010,N_22445,N_22004);
xor U26011 (N_26011,N_22939,N_23739);
or U26012 (N_26012,N_22540,N_21030);
and U26013 (N_26013,N_21511,N_23007);
nor U26014 (N_26014,N_21693,N_22839);
xor U26015 (N_26015,N_22125,N_23689);
nor U26016 (N_26016,N_21148,N_21754);
and U26017 (N_26017,N_21251,N_22341);
xor U26018 (N_26018,N_23032,N_22501);
nor U26019 (N_26019,N_21564,N_21834);
xnor U26020 (N_26020,N_21586,N_23724);
and U26021 (N_26021,N_22342,N_23864);
nand U26022 (N_26022,N_23431,N_21366);
nand U26023 (N_26023,N_22758,N_22194);
and U26024 (N_26024,N_22038,N_22187);
xnor U26025 (N_26025,N_21151,N_23908);
and U26026 (N_26026,N_23367,N_21469);
xor U26027 (N_26027,N_22826,N_22081);
and U26028 (N_26028,N_22608,N_22809);
nand U26029 (N_26029,N_21639,N_21400);
nand U26030 (N_26030,N_22854,N_22879);
xnor U26031 (N_26031,N_23405,N_21345);
or U26032 (N_26032,N_21925,N_23368);
xor U26033 (N_26033,N_21095,N_21998);
or U26034 (N_26034,N_21582,N_21193);
and U26035 (N_26035,N_22592,N_22166);
nor U26036 (N_26036,N_23763,N_22835);
nor U26037 (N_26037,N_21009,N_23722);
nand U26038 (N_26038,N_23047,N_23850);
nand U26039 (N_26039,N_22858,N_21130);
and U26040 (N_26040,N_21475,N_21848);
xor U26041 (N_26041,N_21215,N_23246);
and U26042 (N_26042,N_21391,N_21018);
nand U26043 (N_26043,N_21787,N_23971);
and U26044 (N_26044,N_22308,N_23641);
xor U26045 (N_26045,N_23141,N_23089);
xor U26046 (N_26046,N_22303,N_22968);
nand U26047 (N_26047,N_23884,N_21114);
or U26048 (N_26048,N_23109,N_21495);
xnor U26049 (N_26049,N_21238,N_23453);
nor U26050 (N_26050,N_23691,N_22395);
and U26051 (N_26051,N_23740,N_22034);
nand U26052 (N_26052,N_21167,N_22196);
or U26053 (N_26053,N_21296,N_22308);
and U26054 (N_26054,N_23535,N_23833);
nand U26055 (N_26055,N_21541,N_22291);
or U26056 (N_26056,N_23086,N_21176);
nand U26057 (N_26057,N_22001,N_23082);
xnor U26058 (N_26058,N_22561,N_22946);
and U26059 (N_26059,N_22906,N_22297);
nand U26060 (N_26060,N_22621,N_22237);
nand U26061 (N_26061,N_22804,N_22263);
or U26062 (N_26062,N_21032,N_23031);
nor U26063 (N_26063,N_21646,N_22758);
xor U26064 (N_26064,N_22653,N_22436);
nor U26065 (N_26065,N_21854,N_22014);
nor U26066 (N_26066,N_22929,N_21390);
or U26067 (N_26067,N_22067,N_23251);
xnor U26068 (N_26068,N_22316,N_23882);
nand U26069 (N_26069,N_21370,N_22776);
xnor U26070 (N_26070,N_23865,N_21778);
xnor U26071 (N_26071,N_23642,N_23980);
xnor U26072 (N_26072,N_22725,N_22086);
xor U26073 (N_26073,N_21686,N_21781);
nor U26074 (N_26074,N_21892,N_22963);
xor U26075 (N_26075,N_21330,N_22841);
or U26076 (N_26076,N_23115,N_23665);
and U26077 (N_26077,N_22106,N_23480);
nor U26078 (N_26078,N_21415,N_23236);
and U26079 (N_26079,N_23313,N_22865);
and U26080 (N_26080,N_21805,N_23949);
nor U26081 (N_26081,N_22124,N_22605);
or U26082 (N_26082,N_23034,N_23515);
nor U26083 (N_26083,N_23097,N_23829);
or U26084 (N_26084,N_23252,N_23647);
nand U26085 (N_26085,N_22319,N_22755);
or U26086 (N_26086,N_22455,N_21602);
xor U26087 (N_26087,N_23394,N_21296);
xnor U26088 (N_26088,N_21788,N_22768);
nand U26089 (N_26089,N_21093,N_21860);
or U26090 (N_26090,N_23422,N_23414);
nand U26091 (N_26091,N_23592,N_23284);
nand U26092 (N_26092,N_23998,N_23489);
or U26093 (N_26093,N_22384,N_22014);
and U26094 (N_26094,N_21731,N_23316);
nand U26095 (N_26095,N_23799,N_22594);
and U26096 (N_26096,N_23466,N_21261);
nand U26097 (N_26097,N_23063,N_23677);
and U26098 (N_26098,N_21736,N_22698);
xor U26099 (N_26099,N_23835,N_22695);
and U26100 (N_26100,N_22574,N_23727);
nor U26101 (N_26101,N_23571,N_22430);
nand U26102 (N_26102,N_22712,N_21594);
xnor U26103 (N_26103,N_22246,N_21049);
nor U26104 (N_26104,N_21888,N_23482);
nand U26105 (N_26105,N_21864,N_21746);
nor U26106 (N_26106,N_21714,N_22281);
or U26107 (N_26107,N_23778,N_23666);
nand U26108 (N_26108,N_21842,N_22267);
xnor U26109 (N_26109,N_21375,N_23567);
xnor U26110 (N_26110,N_23847,N_21172);
nor U26111 (N_26111,N_22527,N_23751);
nor U26112 (N_26112,N_21644,N_23847);
or U26113 (N_26113,N_23486,N_21149);
and U26114 (N_26114,N_21095,N_21368);
nand U26115 (N_26115,N_21747,N_22259);
nor U26116 (N_26116,N_21651,N_21145);
or U26117 (N_26117,N_23384,N_22147);
xnor U26118 (N_26118,N_22318,N_21702);
xnor U26119 (N_26119,N_22614,N_21839);
or U26120 (N_26120,N_22672,N_21778);
nand U26121 (N_26121,N_23307,N_23359);
nand U26122 (N_26122,N_22325,N_23112);
xor U26123 (N_26123,N_21825,N_22079);
or U26124 (N_26124,N_21207,N_23306);
xnor U26125 (N_26125,N_23998,N_23699);
and U26126 (N_26126,N_22294,N_22152);
xor U26127 (N_26127,N_23162,N_21073);
xor U26128 (N_26128,N_21951,N_21379);
and U26129 (N_26129,N_22326,N_23533);
or U26130 (N_26130,N_23266,N_23686);
or U26131 (N_26131,N_23079,N_23828);
or U26132 (N_26132,N_21405,N_23705);
nor U26133 (N_26133,N_23780,N_21849);
xor U26134 (N_26134,N_22516,N_21763);
or U26135 (N_26135,N_23998,N_22862);
and U26136 (N_26136,N_22633,N_21209);
nor U26137 (N_26137,N_22359,N_22945);
xnor U26138 (N_26138,N_23114,N_22362);
or U26139 (N_26139,N_23300,N_21216);
and U26140 (N_26140,N_22389,N_21860);
xnor U26141 (N_26141,N_23663,N_22341);
and U26142 (N_26142,N_23634,N_22375);
and U26143 (N_26143,N_21236,N_21864);
or U26144 (N_26144,N_22847,N_22706);
nor U26145 (N_26145,N_21528,N_22426);
nor U26146 (N_26146,N_23101,N_21096);
nand U26147 (N_26147,N_21773,N_22465);
xnor U26148 (N_26148,N_21359,N_22344);
nor U26149 (N_26149,N_21927,N_23991);
and U26150 (N_26150,N_23410,N_22709);
nor U26151 (N_26151,N_22183,N_21127);
or U26152 (N_26152,N_23722,N_21371);
nor U26153 (N_26153,N_22027,N_22406);
nor U26154 (N_26154,N_21402,N_21463);
xor U26155 (N_26155,N_22145,N_21333);
nor U26156 (N_26156,N_23210,N_23088);
xor U26157 (N_26157,N_21635,N_23845);
nor U26158 (N_26158,N_21004,N_22723);
nand U26159 (N_26159,N_23205,N_21350);
xor U26160 (N_26160,N_21692,N_22109);
or U26161 (N_26161,N_22559,N_21805);
xnor U26162 (N_26162,N_22028,N_23543);
nand U26163 (N_26163,N_22366,N_23948);
and U26164 (N_26164,N_21836,N_22001);
nand U26165 (N_26165,N_22018,N_22284);
nand U26166 (N_26166,N_22798,N_23041);
and U26167 (N_26167,N_22958,N_23231);
xor U26168 (N_26168,N_23734,N_22099);
and U26169 (N_26169,N_22792,N_23053);
or U26170 (N_26170,N_23133,N_21518);
xor U26171 (N_26171,N_21196,N_21843);
and U26172 (N_26172,N_22777,N_21231);
nor U26173 (N_26173,N_23159,N_23077);
xnor U26174 (N_26174,N_21268,N_22910);
nand U26175 (N_26175,N_21699,N_21899);
nand U26176 (N_26176,N_23716,N_23939);
nand U26177 (N_26177,N_21354,N_22410);
nor U26178 (N_26178,N_23567,N_23167);
nor U26179 (N_26179,N_22037,N_23824);
and U26180 (N_26180,N_23884,N_22281);
xor U26181 (N_26181,N_22698,N_22549);
and U26182 (N_26182,N_23147,N_23000);
nand U26183 (N_26183,N_21685,N_23261);
and U26184 (N_26184,N_23689,N_22858);
nor U26185 (N_26185,N_21111,N_22517);
and U26186 (N_26186,N_21795,N_22532);
nand U26187 (N_26187,N_23106,N_22895);
xor U26188 (N_26188,N_21316,N_23041);
xnor U26189 (N_26189,N_22992,N_23253);
nor U26190 (N_26190,N_23024,N_22388);
nor U26191 (N_26191,N_22789,N_21692);
nand U26192 (N_26192,N_23753,N_23125);
xor U26193 (N_26193,N_21711,N_21971);
and U26194 (N_26194,N_21903,N_22090);
nor U26195 (N_26195,N_22154,N_22122);
nand U26196 (N_26196,N_23916,N_22664);
nor U26197 (N_26197,N_23084,N_21939);
and U26198 (N_26198,N_23468,N_22192);
nor U26199 (N_26199,N_23775,N_23041);
xnor U26200 (N_26200,N_23286,N_21357);
nand U26201 (N_26201,N_22116,N_22226);
xor U26202 (N_26202,N_23630,N_21557);
nand U26203 (N_26203,N_22552,N_22044);
or U26204 (N_26204,N_21072,N_23934);
and U26205 (N_26205,N_23581,N_22858);
or U26206 (N_26206,N_21001,N_23223);
or U26207 (N_26207,N_22132,N_22847);
nand U26208 (N_26208,N_21078,N_21432);
and U26209 (N_26209,N_23870,N_22738);
xnor U26210 (N_26210,N_22406,N_21014);
nor U26211 (N_26211,N_21994,N_22985);
xor U26212 (N_26212,N_21032,N_23605);
xnor U26213 (N_26213,N_23057,N_22966);
and U26214 (N_26214,N_21144,N_22597);
nor U26215 (N_26215,N_21271,N_22485);
and U26216 (N_26216,N_22845,N_22857);
and U26217 (N_26217,N_21821,N_21603);
and U26218 (N_26218,N_23117,N_22113);
nand U26219 (N_26219,N_21373,N_21477);
or U26220 (N_26220,N_23291,N_21344);
nand U26221 (N_26221,N_21496,N_23393);
nand U26222 (N_26222,N_22281,N_21317);
nor U26223 (N_26223,N_21359,N_23631);
xnor U26224 (N_26224,N_23408,N_23542);
and U26225 (N_26225,N_23454,N_21474);
or U26226 (N_26226,N_21143,N_22253);
nor U26227 (N_26227,N_21728,N_21026);
nor U26228 (N_26228,N_22390,N_22981);
or U26229 (N_26229,N_22827,N_21064);
nor U26230 (N_26230,N_21678,N_22290);
and U26231 (N_26231,N_22513,N_23836);
nand U26232 (N_26232,N_23866,N_23498);
nand U26233 (N_26233,N_23849,N_22277);
xor U26234 (N_26234,N_23750,N_21955);
nand U26235 (N_26235,N_22623,N_22746);
and U26236 (N_26236,N_23949,N_21746);
nor U26237 (N_26237,N_23086,N_23350);
nand U26238 (N_26238,N_23636,N_23198);
nand U26239 (N_26239,N_22396,N_23692);
xor U26240 (N_26240,N_23205,N_22233);
or U26241 (N_26241,N_22921,N_22868);
xnor U26242 (N_26242,N_21085,N_23213);
or U26243 (N_26243,N_22102,N_22986);
and U26244 (N_26244,N_21167,N_21739);
xnor U26245 (N_26245,N_22034,N_21946);
xor U26246 (N_26246,N_23311,N_23358);
or U26247 (N_26247,N_21058,N_21811);
or U26248 (N_26248,N_21613,N_22687);
nor U26249 (N_26249,N_21293,N_23053);
nor U26250 (N_26250,N_23765,N_23805);
or U26251 (N_26251,N_21547,N_22786);
and U26252 (N_26252,N_22410,N_23047);
nand U26253 (N_26253,N_21597,N_23830);
xnor U26254 (N_26254,N_23873,N_21348);
and U26255 (N_26255,N_21063,N_22037);
and U26256 (N_26256,N_21311,N_22951);
xor U26257 (N_26257,N_21775,N_22190);
and U26258 (N_26258,N_22356,N_22748);
and U26259 (N_26259,N_21724,N_21873);
nand U26260 (N_26260,N_21528,N_21358);
nand U26261 (N_26261,N_23918,N_21827);
nor U26262 (N_26262,N_21771,N_21490);
and U26263 (N_26263,N_21033,N_22309);
or U26264 (N_26264,N_23499,N_22100);
nor U26265 (N_26265,N_22938,N_22745);
xor U26266 (N_26266,N_21819,N_22254);
nand U26267 (N_26267,N_23217,N_23546);
nor U26268 (N_26268,N_22044,N_23577);
and U26269 (N_26269,N_21901,N_23954);
nor U26270 (N_26270,N_22682,N_22573);
and U26271 (N_26271,N_21272,N_22052);
or U26272 (N_26272,N_23920,N_22374);
nand U26273 (N_26273,N_21657,N_22016);
and U26274 (N_26274,N_23269,N_23065);
xor U26275 (N_26275,N_22301,N_21229);
nor U26276 (N_26276,N_21684,N_23783);
and U26277 (N_26277,N_22551,N_22778);
and U26278 (N_26278,N_23005,N_21727);
xnor U26279 (N_26279,N_23849,N_22141);
xnor U26280 (N_26280,N_22118,N_21795);
and U26281 (N_26281,N_22233,N_23146);
xor U26282 (N_26282,N_22210,N_23781);
and U26283 (N_26283,N_21417,N_23494);
or U26284 (N_26284,N_23209,N_23974);
nand U26285 (N_26285,N_22911,N_23459);
or U26286 (N_26286,N_21700,N_22655);
nand U26287 (N_26287,N_23093,N_22344);
nor U26288 (N_26288,N_22705,N_22604);
nor U26289 (N_26289,N_22631,N_23495);
nor U26290 (N_26290,N_23332,N_21698);
and U26291 (N_26291,N_21036,N_23296);
nor U26292 (N_26292,N_22639,N_22052);
nand U26293 (N_26293,N_22109,N_23740);
or U26294 (N_26294,N_22257,N_23177);
xor U26295 (N_26295,N_23577,N_21320);
or U26296 (N_26296,N_23887,N_21243);
and U26297 (N_26297,N_21825,N_23737);
nand U26298 (N_26298,N_22182,N_21100);
nor U26299 (N_26299,N_22669,N_23045);
or U26300 (N_26300,N_23259,N_22054);
or U26301 (N_26301,N_21898,N_23013);
or U26302 (N_26302,N_22431,N_22196);
nor U26303 (N_26303,N_21910,N_21648);
nand U26304 (N_26304,N_22333,N_23422);
xor U26305 (N_26305,N_21002,N_23601);
nand U26306 (N_26306,N_23376,N_21250);
xor U26307 (N_26307,N_22796,N_22861);
xnor U26308 (N_26308,N_23634,N_21161);
nand U26309 (N_26309,N_23314,N_22074);
and U26310 (N_26310,N_22381,N_21032);
and U26311 (N_26311,N_21294,N_21172);
or U26312 (N_26312,N_23816,N_22411);
xor U26313 (N_26313,N_23600,N_23180);
nor U26314 (N_26314,N_21892,N_22794);
nand U26315 (N_26315,N_22906,N_23961);
xor U26316 (N_26316,N_22137,N_23194);
xor U26317 (N_26317,N_23631,N_23794);
nor U26318 (N_26318,N_21906,N_21429);
and U26319 (N_26319,N_22727,N_23273);
and U26320 (N_26320,N_22622,N_23937);
xnor U26321 (N_26321,N_21156,N_22143);
nor U26322 (N_26322,N_23652,N_23759);
and U26323 (N_26323,N_23428,N_21968);
or U26324 (N_26324,N_23709,N_22929);
xnor U26325 (N_26325,N_22024,N_23956);
and U26326 (N_26326,N_21052,N_22144);
nor U26327 (N_26327,N_21872,N_22631);
xor U26328 (N_26328,N_21814,N_22216);
or U26329 (N_26329,N_21842,N_21571);
or U26330 (N_26330,N_23790,N_23588);
xnor U26331 (N_26331,N_21632,N_21210);
nand U26332 (N_26332,N_23985,N_23803);
xor U26333 (N_26333,N_23243,N_23883);
nand U26334 (N_26334,N_22719,N_21562);
or U26335 (N_26335,N_22093,N_22884);
xnor U26336 (N_26336,N_23076,N_21331);
and U26337 (N_26337,N_22321,N_21107);
and U26338 (N_26338,N_23587,N_22323);
and U26339 (N_26339,N_22817,N_21670);
nor U26340 (N_26340,N_23626,N_21426);
nand U26341 (N_26341,N_21203,N_23601);
nor U26342 (N_26342,N_23226,N_23056);
nand U26343 (N_26343,N_21063,N_23571);
xor U26344 (N_26344,N_22528,N_21397);
nand U26345 (N_26345,N_21385,N_23436);
and U26346 (N_26346,N_21409,N_23333);
nand U26347 (N_26347,N_22868,N_23212);
nand U26348 (N_26348,N_23521,N_23745);
and U26349 (N_26349,N_23491,N_23570);
nand U26350 (N_26350,N_23011,N_23001);
nand U26351 (N_26351,N_23010,N_21641);
nor U26352 (N_26352,N_23367,N_23221);
xnor U26353 (N_26353,N_21738,N_21280);
or U26354 (N_26354,N_21891,N_22705);
nor U26355 (N_26355,N_23321,N_21335);
nor U26356 (N_26356,N_22116,N_21432);
xnor U26357 (N_26357,N_22912,N_21811);
or U26358 (N_26358,N_21518,N_22755);
or U26359 (N_26359,N_22735,N_21270);
or U26360 (N_26360,N_22878,N_21526);
nor U26361 (N_26361,N_21364,N_21331);
and U26362 (N_26362,N_23636,N_22947);
nand U26363 (N_26363,N_21528,N_23312);
xnor U26364 (N_26364,N_21316,N_23356);
nor U26365 (N_26365,N_23599,N_22722);
nand U26366 (N_26366,N_22805,N_21417);
nand U26367 (N_26367,N_23429,N_22496);
or U26368 (N_26368,N_23952,N_23014);
nand U26369 (N_26369,N_23648,N_23952);
xnor U26370 (N_26370,N_22809,N_22400);
and U26371 (N_26371,N_22105,N_21333);
and U26372 (N_26372,N_22839,N_21110);
xor U26373 (N_26373,N_21009,N_21043);
and U26374 (N_26374,N_23786,N_22886);
or U26375 (N_26375,N_23042,N_21664);
xnor U26376 (N_26376,N_23051,N_23969);
nor U26377 (N_26377,N_21733,N_22469);
xor U26378 (N_26378,N_23437,N_23482);
and U26379 (N_26379,N_22885,N_23642);
nand U26380 (N_26380,N_21715,N_21418);
or U26381 (N_26381,N_23485,N_22243);
nor U26382 (N_26382,N_21032,N_22715);
xor U26383 (N_26383,N_23695,N_21103);
or U26384 (N_26384,N_21174,N_21841);
nor U26385 (N_26385,N_22604,N_22501);
and U26386 (N_26386,N_21142,N_21680);
or U26387 (N_26387,N_22529,N_22708);
xor U26388 (N_26388,N_21231,N_23850);
xnor U26389 (N_26389,N_22231,N_21038);
xnor U26390 (N_26390,N_21975,N_22472);
or U26391 (N_26391,N_21320,N_23989);
and U26392 (N_26392,N_22570,N_22609);
or U26393 (N_26393,N_22832,N_22186);
xnor U26394 (N_26394,N_22854,N_21866);
nor U26395 (N_26395,N_22376,N_21969);
nand U26396 (N_26396,N_21384,N_23183);
xnor U26397 (N_26397,N_23899,N_21197);
nor U26398 (N_26398,N_22912,N_21551);
or U26399 (N_26399,N_21859,N_21368);
nor U26400 (N_26400,N_22874,N_22892);
nor U26401 (N_26401,N_23623,N_23245);
nand U26402 (N_26402,N_22352,N_22840);
xnor U26403 (N_26403,N_22726,N_21940);
or U26404 (N_26404,N_21910,N_22470);
or U26405 (N_26405,N_21936,N_22641);
nand U26406 (N_26406,N_22664,N_21020);
nand U26407 (N_26407,N_23326,N_23358);
nor U26408 (N_26408,N_21611,N_22786);
nor U26409 (N_26409,N_21391,N_23708);
nand U26410 (N_26410,N_23028,N_23532);
and U26411 (N_26411,N_22128,N_21453);
and U26412 (N_26412,N_21217,N_23937);
nand U26413 (N_26413,N_21312,N_22743);
and U26414 (N_26414,N_23632,N_22660);
nor U26415 (N_26415,N_23088,N_22329);
or U26416 (N_26416,N_21787,N_23987);
nand U26417 (N_26417,N_22282,N_23314);
nand U26418 (N_26418,N_21167,N_23243);
or U26419 (N_26419,N_22507,N_22413);
xor U26420 (N_26420,N_21140,N_22615);
xnor U26421 (N_26421,N_21657,N_23409);
nor U26422 (N_26422,N_21902,N_22556);
xor U26423 (N_26423,N_22297,N_22856);
and U26424 (N_26424,N_22766,N_23309);
and U26425 (N_26425,N_23017,N_23253);
nor U26426 (N_26426,N_21030,N_22120);
or U26427 (N_26427,N_21451,N_21181);
nand U26428 (N_26428,N_23894,N_22223);
and U26429 (N_26429,N_23258,N_21195);
and U26430 (N_26430,N_21004,N_22176);
nor U26431 (N_26431,N_21946,N_22800);
nor U26432 (N_26432,N_21192,N_21200);
or U26433 (N_26433,N_21999,N_21227);
or U26434 (N_26434,N_21323,N_21370);
nor U26435 (N_26435,N_23390,N_22937);
nand U26436 (N_26436,N_21317,N_21858);
nor U26437 (N_26437,N_22686,N_23740);
nand U26438 (N_26438,N_23120,N_22859);
and U26439 (N_26439,N_22767,N_21415);
and U26440 (N_26440,N_23625,N_22602);
nor U26441 (N_26441,N_23240,N_21821);
nor U26442 (N_26442,N_22514,N_23302);
or U26443 (N_26443,N_22513,N_21137);
and U26444 (N_26444,N_23079,N_23537);
or U26445 (N_26445,N_23738,N_22736);
nor U26446 (N_26446,N_23875,N_23524);
nand U26447 (N_26447,N_23953,N_22469);
nand U26448 (N_26448,N_23586,N_21090);
nand U26449 (N_26449,N_23950,N_22363);
nand U26450 (N_26450,N_23685,N_23287);
or U26451 (N_26451,N_22937,N_21533);
and U26452 (N_26452,N_22872,N_21833);
xor U26453 (N_26453,N_23438,N_23033);
xnor U26454 (N_26454,N_23797,N_23415);
and U26455 (N_26455,N_23317,N_22810);
nand U26456 (N_26456,N_21864,N_21833);
or U26457 (N_26457,N_23773,N_22201);
and U26458 (N_26458,N_23245,N_22705);
xnor U26459 (N_26459,N_23073,N_21280);
xor U26460 (N_26460,N_23314,N_21551);
and U26461 (N_26461,N_22306,N_22242);
and U26462 (N_26462,N_22491,N_23861);
and U26463 (N_26463,N_21238,N_23645);
and U26464 (N_26464,N_23869,N_21615);
or U26465 (N_26465,N_23337,N_21370);
or U26466 (N_26466,N_21921,N_22716);
xnor U26467 (N_26467,N_21811,N_23829);
or U26468 (N_26468,N_22630,N_21621);
nor U26469 (N_26469,N_22285,N_21920);
and U26470 (N_26470,N_21686,N_21516);
or U26471 (N_26471,N_22061,N_22594);
nor U26472 (N_26472,N_23470,N_23169);
nor U26473 (N_26473,N_21528,N_23314);
xnor U26474 (N_26474,N_23873,N_21356);
or U26475 (N_26475,N_22140,N_22801);
xnor U26476 (N_26476,N_21441,N_23703);
or U26477 (N_26477,N_22867,N_21959);
nor U26478 (N_26478,N_21273,N_22502);
nor U26479 (N_26479,N_23414,N_23195);
nor U26480 (N_26480,N_22016,N_21636);
and U26481 (N_26481,N_22049,N_21841);
or U26482 (N_26482,N_22689,N_22159);
and U26483 (N_26483,N_21989,N_22276);
xnor U26484 (N_26484,N_22373,N_22019);
and U26485 (N_26485,N_21244,N_21335);
xor U26486 (N_26486,N_23466,N_22176);
xor U26487 (N_26487,N_21216,N_23105);
nor U26488 (N_26488,N_22904,N_21936);
and U26489 (N_26489,N_23193,N_21270);
or U26490 (N_26490,N_23288,N_23979);
xnor U26491 (N_26491,N_21716,N_21462);
xnor U26492 (N_26492,N_21217,N_23624);
and U26493 (N_26493,N_22812,N_22830);
and U26494 (N_26494,N_22054,N_21094);
nand U26495 (N_26495,N_22678,N_23294);
xnor U26496 (N_26496,N_23575,N_21368);
and U26497 (N_26497,N_21359,N_21307);
nand U26498 (N_26498,N_21792,N_21910);
and U26499 (N_26499,N_22716,N_21739);
or U26500 (N_26500,N_22122,N_22381);
nor U26501 (N_26501,N_21326,N_23900);
or U26502 (N_26502,N_22107,N_22701);
nor U26503 (N_26503,N_23080,N_23756);
nand U26504 (N_26504,N_23055,N_21205);
and U26505 (N_26505,N_21750,N_23159);
or U26506 (N_26506,N_22486,N_23892);
or U26507 (N_26507,N_21821,N_21527);
nand U26508 (N_26508,N_21303,N_23317);
or U26509 (N_26509,N_23619,N_23864);
nand U26510 (N_26510,N_21148,N_22228);
xor U26511 (N_26511,N_23495,N_21720);
nor U26512 (N_26512,N_23617,N_22625);
nand U26513 (N_26513,N_23080,N_21032);
nor U26514 (N_26514,N_22641,N_23453);
nor U26515 (N_26515,N_22747,N_23736);
or U26516 (N_26516,N_22255,N_23999);
and U26517 (N_26517,N_21646,N_21866);
xor U26518 (N_26518,N_21962,N_22001);
or U26519 (N_26519,N_22688,N_23496);
nand U26520 (N_26520,N_21991,N_23182);
nand U26521 (N_26521,N_22200,N_22005);
or U26522 (N_26522,N_21206,N_21234);
and U26523 (N_26523,N_22855,N_22292);
nand U26524 (N_26524,N_22201,N_23307);
or U26525 (N_26525,N_23146,N_21397);
or U26526 (N_26526,N_21431,N_23795);
nand U26527 (N_26527,N_21431,N_23053);
or U26528 (N_26528,N_21712,N_21525);
nor U26529 (N_26529,N_21916,N_23366);
nor U26530 (N_26530,N_23828,N_22548);
nor U26531 (N_26531,N_21397,N_23174);
or U26532 (N_26532,N_22377,N_23823);
or U26533 (N_26533,N_23598,N_23366);
nand U26534 (N_26534,N_22734,N_22125);
xor U26535 (N_26535,N_23851,N_21372);
or U26536 (N_26536,N_21618,N_21783);
xor U26537 (N_26537,N_21680,N_23021);
or U26538 (N_26538,N_22771,N_21886);
and U26539 (N_26539,N_23143,N_22284);
or U26540 (N_26540,N_22398,N_21308);
xor U26541 (N_26541,N_21065,N_21726);
and U26542 (N_26542,N_22286,N_23328);
nor U26543 (N_26543,N_22670,N_21995);
or U26544 (N_26544,N_23149,N_23017);
nand U26545 (N_26545,N_22529,N_22220);
or U26546 (N_26546,N_23835,N_23607);
nor U26547 (N_26547,N_21674,N_23271);
xnor U26548 (N_26548,N_21467,N_22938);
nor U26549 (N_26549,N_21993,N_21834);
and U26550 (N_26550,N_21899,N_21341);
xor U26551 (N_26551,N_21847,N_22358);
nor U26552 (N_26552,N_23141,N_21040);
xnor U26553 (N_26553,N_21384,N_21967);
nand U26554 (N_26554,N_22318,N_22314);
nor U26555 (N_26555,N_22795,N_22455);
nor U26556 (N_26556,N_22108,N_22626);
xor U26557 (N_26557,N_21207,N_21047);
or U26558 (N_26558,N_21309,N_21505);
xor U26559 (N_26559,N_22683,N_21367);
nand U26560 (N_26560,N_22028,N_22505);
xor U26561 (N_26561,N_22991,N_23961);
and U26562 (N_26562,N_21324,N_22731);
xnor U26563 (N_26563,N_22560,N_21238);
nor U26564 (N_26564,N_23988,N_22077);
xnor U26565 (N_26565,N_23641,N_21707);
xnor U26566 (N_26566,N_21729,N_22988);
nand U26567 (N_26567,N_22615,N_23989);
xnor U26568 (N_26568,N_23728,N_21259);
and U26569 (N_26569,N_22449,N_23040);
nor U26570 (N_26570,N_21197,N_23905);
and U26571 (N_26571,N_23173,N_23284);
nor U26572 (N_26572,N_22637,N_22424);
xor U26573 (N_26573,N_22356,N_22988);
nor U26574 (N_26574,N_22349,N_22644);
nand U26575 (N_26575,N_22562,N_23705);
or U26576 (N_26576,N_23772,N_23442);
or U26577 (N_26577,N_21828,N_22572);
nand U26578 (N_26578,N_23299,N_21208);
xnor U26579 (N_26579,N_23912,N_21812);
and U26580 (N_26580,N_21803,N_23054);
or U26581 (N_26581,N_23066,N_21521);
or U26582 (N_26582,N_21636,N_22895);
nand U26583 (N_26583,N_21087,N_21211);
nor U26584 (N_26584,N_22156,N_22586);
nor U26585 (N_26585,N_22221,N_21484);
nand U26586 (N_26586,N_22967,N_23080);
and U26587 (N_26587,N_21875,N_22459);
nand U26588 (N_26588,N_23072,N_23290);
or U26589 (N_26589,N_21081,N_21926);
xor U26590 (N_26590,N_21217,N_21226);
nor U26591 (N_26591,N_21150,N_22661);
nor U26592 (N_26592,N_21676,N_23110);
or U26593 (N_26593,N_23030,N_22121);
xor U26594 (N_26594,N_23521,N_23869);
and U26595 (N_26595,N_23668,N_21433);
nor U26596 (N_26596,N_22101,N_23540);
nor U26597 (N_26597,N_23405,N_22833);
or U26598 (N_26598,N_23101,N_23047);
and U26599 (N_26599,N_21207,N_21623);
nand U26600 (N_26600,N_21951,N_21524);
xor U26601 (N_26601,N_23049,N_22065);
xnor U26602 (N_26602,N_21997,N_22927);
xnor U26603 (N_26603,N_21510,N_22111);
or U26604 (N_26604,N_22124,N_23354);
or U26605 (N_26605,N_21190,N_23503);
and U26606 (N_26606,N_21833,N_22667);
nand U26607 (N_26607,N_23256,N_22596);
xor U26608 (N_26608,N_22472,N_23327);
nor U26609 (N_26609,N_23913,N_21869);
and U26610 (N_26610,N_21108,N_23256);
xor U26611 (N_26611,N_21416,N_22034);
or U26612 (N_26612,N_22663,N_21236);
nand U26613 (N_26613,N_22107,N_21328);
nand U26614 (N_26614,N_23144,N_23480);
nand U26615 (N_26615,N_22453,N_21017);
xnor U26616 (N_26616,N_23847,N_21627);
and U26617 (N_26617,N_21188,N_23142);
and U26618 (N_26618,N_22501,N_23227);
nand U26619 (N_26619,N_22515,N_22670);
nand U26620 (N_26620,N_23698,N_22821);
or U26621 (N_26621,N_22771,N_22405);
nor U26622 (N_26622,N_22435,N_22349);
xnor U26623 (N_26623,N_22325,N_22445);
and U26624 (N_26624,N_23908,N_22770);
xor U26625 (N_26625,N_21270,N_23810);
and U26626 (N_26626,N_22594,N_21737);
xnor U26627 (N_26627,N_21980,N_21846);
nor U26628 (N_26628,N_22001,N_22680);
nand U26629 (N_26629,N_22167,N_23857);
or U26630 (N_26630,N_23758,N_23201);
xor U26631 (N_26631,N_21012,N_23498);
xnor U26632 (N_26632,N_22497,N_22185);
nand U26633 (N_26633,N_23580,N_23519);
and U26634 (N_26634,N_22216,N_23395);
nand U26635 (N_26635,N_23439,N_22993);
and U26636 (N_26636,N_23988,N_22605);
and U26637 (N_26637,N_22688,N_23944);
xor U26638 (N_26638,N_23952,N_21631);
or U26639 (N_26639,N_22614,N_21916);
or U26640 (N_26640,N_21405,N_23027);
or U26641 (N_26641,N_23431,N_22902);
xnor U26642 (N_26642,N_22858,N_22961);
or U26643 (N_26643,N_23996,N_22907);
xnor U26644 (N_26644,N_22071,N_21018);
xnor U26645 (N_26645,N_21600,N_21277);
or U26646 (N_26646,N_23700,N_23711);
or U26647 (N_26647,N_22750,N_22060);
nand U26648 (N_26648,N_21868,N_23707);
and U26649 (N_26649,N_22402,N_22974);
nor U26650 (N_26650,N_22183,N_23041);
nor U26651 (N_26651,N_23365,N_22250);
xor U26652 (N_26652,N_22477,N_22955);
xnor U26653 (N_26653,N_21897,N_22895);
xor U26654 (N_26654,N_23649,N_22871);
nand U26655 (N_26655,N_22413,N_21025);
nor U26656 (N_26656,N_21776,N_21254);
or U26657 (N_26657,N_21727,N_22246);
or U26658 (N_26658,N_23069,N_21685);
and U26659 (N_26659,N_22200,N_21969);
nand U26660 (N_26660,N_21319,N_23363);
nand U26661 (N_26661,N_22010,N_21713);
nor U26662 (N_26662,N_22297,N_22633);
nor U26663 (N_26663,N_22654,N_21086);
and U26664 (N_26664,N_23539,N_21973);
xor U26665 (N_26665,N_23281,N_21772);
and U26666 (N_26666,N_22231,N_23398);
and U26667 (N_26667,N_21995,N_22931);
or U26668 (N_26668,N_21986,N_22958);
and U26669 (N_26669,N_22143,N_22568);
or U26670 (N_26670,N_22599,N_21605);
and U26671 (N_26671,N_22304,N_23190);
or U26672 (N_26672,N_22843,N_23213);
xor U26673 (N_26673,N_22617,N_23313);
or U26674 (N_26674,N_23938,N_21994);
and U26675 (N_26675,N_22390,N_22895);
or U26676 (N_26676,N_22887,N_23417);
nor U26677 (N_26677,N_22529,N_22928);
xor U26678 (N_26678,N_21767,N_22686);
nand U26679 (N_26679,N_22460,N_23025);
xnor U26680 (N_26680,N_21584,N_21586);
and U26681 (N_26681,N_21418,N_21316);
nand U26682 (N_26682,N_21764,N_21031);
and U26683 (N_26683,N_23319,N_22387);
nand U26684 (N_26684,N_23182,N_21849);
nand U26685 (N_26685,N_23888,N_21166);
nor U26686 (N_26686,N_23045,N_22673);
nor U26687 (N_26687,N_22048,N_23983);
and U26688 (N_26688,N_22526,N_21358);
or U26689 (N_26689,N_22820,N_23576);
or U26690 (N_26690,N_23919,N_23140);
or U26691 (N_26691,N_21488,N_23145);
and U26692 (N_26692,N_22969,N_22013);
or U26693 (N_26693,N_21058,N_22498);
xor U26694 (N_26694,N_21498,N_21468);
xor U26695 (N_26695,N_22926,N_23422);
and U26696 (N_26696,N_23900,N_22119);
or U26697 (N_26697,N_21891,N_22235);
nand U26698 (N_26698,N_21844,N_22988);
xor U26699 (N_26699,N_22662,N_22811);
and U26700 (N_26700,N_21514,N_21834);
xnor U26701 (N_26701,N_21745,N_21310);
xnor U26702 (N_26702,N_22214,N_22053);
or U26703 (N_26703,N_21912,N_21087);
nor U26704 (N_26704,N_22147,N_22861);
and U26705 (N_26705,N_22702,N_22909);
xor U26706 (N_26706,N_23457,N_23059);
nand U26707 (N_26707,N_21470,N_23688);
nand U26708 (N_26708,N_22786,N_21668);
xnor U26709 (N_26709,N_22902,N_23490);
nand U26710 (N_26710,N_21215,N_21600);
and U26711 (N_26711,N_22822,N_22053);
nor U26712 (N_26712,N_22327,N_22469);
nor U26713 (N_26713,N_23152,N_22900);
xnor U26714 (N_26714,N_23622,N_21896);
or U26715 (N_26715,N_21188,N_23380);
nand U26716 (N_26716,N_23245,N_22841);
nor U26717 (N_26717,N_21763,N_21601);
nand U26718 (N_26718,N_23140,N_22538);
or U26719 (N_26719,N_23136,N_23300);
nand U26720 (N_26720,N_21093,N_23412);
and U26721 (N_26721,N_21836,N_23712);
nand U26722 (N_26722,N_22211,N_23373);
xnor U26723 (N_26723,N_21747,N_23370);
xor U26724 (N_26724,N_23340,N_21488);
xnor U26725 (N_26725,N_22828,N_21690);
and U26726 (N_26726,N_23627,N_21722);
nor U26727 (N_26727,N_22051,N_21440);
and U26728 (N_26728,N_23790,N_23781);
xnor U26729 (N_26729,N_23881,N_23752);
or U26730 (N_26730,N_21920,N_22877);
xnor U26731 (N_26731,N_23620,N_21818);
and U26732 (N_26732,N_23874,N_22407);
nand U26733 (N_26733,N_22633,N_21938);
and U26734 (N_26734,N_21495,N_22035);
nor U26735 (N_26735,N_22412,N_22112);
nor U26736 (N_26736,N_21201,N_22150);
or U26737 (N_26737,N_23409,N_23932);
nor U26738 (N_26738,N_23216,N_21808);
or U26739 (N_26739,N_21364,N_21979);
or U26740 (N_26740,N_22219,N_23344);
nor U26741 (N_26741,N_21473,N_23044);
and U26742 (N_26742,N_21870,N_21362);
xor U26743 (N_26743,N_23426,N_22560);
xnor U26744 (N_26744,N_22494,N_21763);
nand U26745 (N_26745,N_22851,N_21686);
nor U26746 (N_26746,N_21184,N_21707);
nor U26747 (N_26747,N_22244,N_21149);
xor U26748 (N_26748,N_22747,N_22235);
or U26749 (N_26749,N_22051,N_22837);
xor U26750 (N_26750,N_21181,N_22572);
or U26751 (N_26751,N_21861,N_22490);
or U26752 (N_26752,N_21792,N_22753);
xnor U26753 (N_26753,N_21880,N_21599);
nand U26754 (N_26754,N_21683,N_23787);
nand U26755 (N_26755,N_21063,N_23175);
nor U26756 (N_26756,N_22642,N_22469);
nand U26757 (N_26757,N_23387,N_23781);
and U26758 (N_26758,N_21389,N_21094);
and U26759 (N_26759,N_21142,N_23317);
nor U26760 (N_26760,N_23899,N_23002);
xnor U26761 (N_26761,N_23682,N_23796);
or U26762 (N_26762,N_23650,N_21854);
xor U26763 (N_26763,N_22819,N_23649);
and U26764 (N_26764,N_22541,N_23880);
nand U26765 (N_26765,N_22786,N_23464);
nand U26766 (N_26766,N_22842,N_21641);
nor U26767 (N_26767,N_22927,N_21735);
nand U26768 (N_26768,N_21390,N_23368);
or U26769 (N_26769,N_23346,N_21186);
xnor U26770 (N_26770,N_22547,N_22614);
xnor U26771 (N_26771,N_22599,N_23252);
nand U26772 (N_26772,N_21137,N_21871);
or U26773 (N_26773,N_22908,N_22633);
nor U26774 (N_26774,N_21237,N_23519);
nor U26775 (N_26775,N_22915,N_23407);
or U26776 (N_26776,N_23177,N_22859);
xor U26777 (N_26777,N_23328,N_22676);
and U26778 (N_26778,N_22612,N_23333);
xor U26779 (N_26779,N_22284,N_22389);
or U26780 (N_26780,N_21016,N_21335);
or U26781 (N_26781,N_23129,N_23698);
nand U26782 (N_26782,N_21354,N_21975);
and U26783 (N_26783,N_23619,N_23271);
and U26784 (N_26784,N_21479,N_23166);
xnor U26785 (N_26785,N_21157,N_21185);
nor U26786 (N_26786,N_23946,N_22829);
and U26787 (N_26787,N_22970,N_23393);
and U26788 (N_26788,N_21215,N_23282);
xnor U26789 (N_26789,N_23747,N_21751);
nand U26790 (N_26790,N_21433,N_23156);
nand U26791 (N_26791,N_22791,N_23885);
xor U26792 (N_26792,N_21391,N_23258);
xor U26793 (N_26793,N_23152,N_21245);
or U26794 (N_26794,N_21656,N_23247);
and U26795 (N_26795,N_21010,N_23150);
nor U26796 (N_26796,N_23544,N_23051);
or U26797 (N_26797,N_23123,N_21710);
xor U26798 (N_26798,N_23427,N_22120);
xor U26799 (N_26799,N_21500,N_23326);
nor U26800 (N_26800,N_23008,N_21654);
nor U26801 (N_26801,N_23459,N_22726);
or U26802 (N_26802,N_22924,N_22168);
or U26803 (N_26803,N_21427,N_21139);
or U26804 (N_26804,N_22941,N_23386);
nor U26805 (N_26805,N_23149,N_22695);
nand U26806 (N_26806,N_21849,N_21844);
nand U26807 (N_26807,N_22026,N_22219);
nor U26808 (N_26808,N_22458,N_22515);
nand U26809 (N_26809,N_23533,N_21813);
and U26810 (N_26810,N_22050,N_22642);
nand U26811 (N_26811,N_21034,N_22606);
nand U26812 (N_26812,N_22064,N_22688);
xnor U26813 (N_26813,N_23640,N_21868);
xnor U26814 (N_26814,N_21821,N_22216);
and U26815 (N_26815,N_21652,N_21371);
xnor U26816 (N_26816,N_21493,N_21743);
or U26817 (N_26817,N_21422,N_21718);
or U26818 (N_26818,N_21091,N_21540);
nor U26819 (N_26819,N_21234,N_22112);
nand U26820 (N_26820,N_22219,N_23430);
xor U26821 (N_26821,N_23736,N_23069);
nor U26822 (N_26822,N_21983,N_21306);
nand U26823 (N_26823,N_21476,N_21783);
xnor U26824 (N_26824,N_22109,N_22897);
and U26825 (N_26825,N_23137,N_22625);
nor U26826 (N_26826,N_21649,N_21417);
or U26827 (N_26827,N_23201,N_23520);
nand U26828 (N_26828,N_23240,N_22182);
and U26829 (N_26829,N_23998,N_22222);
or U26830 (N_26830,N_23944,N_21214);
and U26831 (N_26831,N_21536,N_23746);
or U26832 (N_26832,N_21449,N_21290);
nand U26833 (N_26833,N_22517,N_23321);
nand U26834 (N_26834,N_22779,N_22637);
and U26835 (N_26835,N_22989,N_21893);
nand U26836 (N_26836,N_22400,N_21434);
nor U26837 (N_26837,N_23192,N_23002);
xnor U26838 (N_26838,N_22787,N_22390);
xor U26839 (N_26839,N_23009,N_21807);
or U26840 (N_26840,N_21836,N_22790);
or U26841 (N_26841,N_21693,N_23519);
nand U26842 (N_26842,N_22286,N_22653);
nor U26843 (N_26843,N_22860,N_22942);
or U26844 (N_26844,N_21060,N_23308);
and U26845 (N_26845,N_23720,N_23578);
nor U26846 (N_26846,N_23819,N_23481);
or U26847 (N_26847,N_22552,N_21757);
or U26848 (N_26848,N_22708,N_22896);
nand U26849 (N_26849,N_23511,N_22663);
xor U26850 (N_26850,N_21467,N_22583);
or U26851 (N_26851,N_23848,N_21475);
xnor U26852 (N_26852,N_23514,N_21199);
nand U26853 (N_26853,N_23255,N_22816);
nor U26854 (N_26854,N_23519,N_23663);
and U26855 (N_26855,N_22399,N_22743);
nor U26856 (N_26856,N_23248,N_21117);
nor U26857 (N_26857,N_23214,N_22864);
nand U26858 (N_26858,N_21650,N_21400);
or U26859 (N_26859,N_23946,N_22723);
nor U26860 (N_26860,N_21359,N_23174);
nand U26861 (N_26861,N_22286,N_23423);
xor U26862 (N_26862,N_21814,N_21990);
nor U26863 (N_26863,N_21194,N_21604);
nand U26864 (N_26864,N_21306,N_23419);
xor U26865 (N_26865,N_21574,N_21078);
xor U26866 (N_26866,N_21424,N_21946);
nor U26867 (N_26867,N_21435,N_23486);
nand U26868 (N_26868,N_22172,N_22975);
and U26869 (N_26869,N_21145,N_22336);
nand U26870 (N_26870,N_22657,N_23211);
nor U26871 (N_26871,N_21542,N_23852);
nor U26872 (N_26872,N_21550,N_23707);
nor U26873 (N_26873,N_22415,N_22622);
or U26874 (N_26874,N_23192,N_22391);
nand U26875 (N_26875,N_22412,N_21576);
xor U26876 (N_26876,N_22815,N_22942);
or U26877 (N_26877,N_23435,N_21726);
xor U26878 (N_26878,N_21485,N_23303);
nor U26879 (N_26879,N_21184,N_21309);
nor U26880 (N_26880,N_23993,N_23808);
xnor U26881 (N_26881,N_21370,N_22720);
xnor U26882 (N_26882,N_22123,N_22156);
nor U26883 (N_26883,N_22242,N_22352);
nand U26884 (N_26884,N_21772,N_23843);
nand U26885 (N_26885,N_22969,N_21565);
or U26886 (N_26886,N_22694,N_21540);
or U26887 (N_26887,N_22985,N_21452);
and U26888 (N_26888,N_23395,N_23243);
and U26889 (N_26889,N_21108,N_21651);
nand U26890 (N_26890,N_21580,N_23209);
nor U26891 (N_26891,N_22670,N_21060);
and U26892 (N_26892,N_23347,N_22611);
xor U26893 (N_26893,N_21966,N_21793);
nand U26894 (N_26894,N_22449,N_21164);
or U26895 (N_26895,N_22975,N_21101);
xor U26896 (N_26896,N_21035,N_22377);
and U26897 (N_26897,N_23461,N_21289);
or U26898 (N_26898,N_22692,N_23836);
nand U26899 (N_26899,N_21665,N_22475);
nor U26900 (N_26900,N_22129,N_22867);
or U26901 (N_26901,N_21157,N_22368);
or U26902 (N_26902,N_22488,N_23396);
xor U26903 (N_26903,N_22651,N_22637);
nand U26904 (N_26904,N_22172,N_23872);
xor U26905 (N_26905,N_22388,N_22851);
nand U26906 (N_26906,N_23622,N_21338);
xor U26907 (N_26907,N_22194,N_22104);
xnor U26908 (N_26908,N_22892,N_23058);
nand U26909 (N_26909,N_22631,N_21648);
nand U26910 (N_26910,N_23699,N_23104);
xor U26911 (N_26911,N_22527,N_22834);
nor U26912 (N_26912,N_21937,N_23905);
or U26913 (N_26913,N_23933,N_21100);
nand U26914 (N_26914,N_21333,N_23626);
and U26915 (N_26915,N_22509,N_21046);
nand U26916 (N_26916,N_21344,N_22623);
and U26917 (N_26917,N_22309,N_23761);
or U26918 (N_26918,N_23847,N_22458);
xnor U26919 (N_26919,N_23617,N_21324);
xnor U26920 (N_26920,N_22890,N_23991);
nand U26921 (N_26921,N_23407,N_21722);
nand U26922 (N_26922,N_21538,N_21381);
or U26923 (N_26923,N_21051,N_22758);
and U26924 (N_26924,N_21264,N_21103);
nand U26925 (N_26925,N_22110,N_21216);
or U26926 (N_26926,N_23322,N_22122);
nand U26927 (N_26927,N_21656,N_22842);
or U26928 (N_26928,N_22556,N_22726);
and U26929 (N_26929,N_22269,N_23051);
nor U26930 (N_26930,N_21394,N_22310);
xor U26931 (N_26931,N_21507,N_21278);
and U26932 (N_26932,N_22151,N_21483);
or U26933 (N_26933,N_21099,N_23622);
xor U26934 (N_26934,N_21208,N_22944);
and U26935 (N_26935,N_23037,N_21468);
nor U26936 (N_26936,N_22263,N_22976);
nand U26937 (N_26937,N_23162,N_21482);
and U26938 (N_26938,N_22057,N_22453);
nor U26939 (N_26939,N_21817,N_21236);
or U26940 (N_26940,N_23850,N_22696);
nor U26941 (N_26941,N_23438,N_22045);
nand U26942 (N_26942,N_23561,N_22397);
and U26943 (N_26943,N_22466,N_22940);
nand U26944 (N_26944,N_22145,N_23812);
xor U26945 (N_26945,N_22600,N_22440);
nor U26946 (N_26946,N_23893,N_22256);
and U26947 (N_26947,N_21832,N_22032);
nor U26948 (N_26948,N_21561,N_22447);
nand U26949 (N_26949,N_23262,N_21890);
and U26950 (N_26950,N_23580,N_21007);
or U26951 (N_26951,N_21389,N_23127);
or U26952 (N_26952,N_21165,N_23022);
and U26953 (N_26953,N_23653,N_21429);
xor U26954 (N_26954,N_21248,N_21990);
xnor U26955 (N_26955,N_23360,N_21681);
and U26956 (N_26956,N_22408,N_21044);
nand U26957 (N_26957,N_23050,N_23482);
nand U26958 (N_26958,N_23184,N_21297);
xor U26959 (N_26959,N_22324,N_22499);
xnor U26960 (N_26960,N_22223,N_23501);
nor U26961 (N_26961,N_22879,N_22950);
nor U26962 (N_26962,N_22381,N_22793);
and U26963 (N_26963,N_23394,N_21442);
and U26964 (N_26964,N_23745,N_22603);
or U26965 (N_26965,N_22405,N_23850);
nor U26966 (N_26966,N_23333,N_21248);
or U26967 (N_26967,N_21162,N_23044);
xnor U26968 (N_26968,N_23404,N_22372);
or U26969 (N_26969,N_21909,N_22821);
xor U26970 (N_26970,N_21318,N_23506);
or U26971 (N_26971,N_21837,N_22691);
nor U26972 (N_26972,N_21100,N_23075);
nand U26973 (N_26973,N_22926,N_21317);
and U26974 (N_26974,N_21536,N_21460);
nor U26975 (N_26975,N_23713,N_21180);
nor U26976 (N_26976,N_23988,N_23663);
or U26977 (N_26977,N_22410,N_22058);
nor U26978 (N_26978,N_22706,N_21358);
nor U26979 (N_26979,N_22698,N_22077);
nand U26980 (N_26980,N_22772,N_21134);
nor U26981 (N_26981,N_22940,N_21066);
and U26982 (N_26982,N_23323,N_23542);
nand U26983 (N_26983,N_22335,N_23847);
xnor U26984 (N_26984,N_23927,N_21883);
nor U26985 (N_26985,N_23233,N_21367);
or U26986 (N_26986,N_22293,N_21405);
and U26987 (N_26987,N_22772,N_23050);
or U26988 (N_26988,N_21264,N_21006);
and U26989 (N_26989,N_21159,N_22796);
or U26990 (N_26990,N_22459,N_22857);
or U26991 (N_26991,N_21570,N_23037);
nor U26992 (N_26992,N_23271,N_22374);
nand U26993 (N_26993,N_23681,N_21253);
nand U26994 (N_26994,N_21790,N_21968);
xor U26995 (N_26995,N_21379,N_21739);
and U26996 (N_26996,N_22775,N_23030);
nor U26997 (N_26997,N_22600,N_21300);
xor U26998 (N_26998,N_21498,N_22010);
xor U26999 (N_26999,N_22394,N_22425);
nor U27000 (N_27000,N_25553,N_24937);
xnor U27001 (N_27001,N_26428,N_26028);
xnor U27002 (N_27002,N_25825,N_24096);
xnor U27003 (N_27003,N_25969,N_24837);
nand U27004 (N_27004,N_26116,N_25882);
nor U27005 (N_27005,N_25193,N_26823);
and U27006 (N_27006,N_25275,N_24359);
nand U27007 (N_27007,N_25594,N_25347);
nor U27008 (N_27008,N_26389,N_26250);
nand U27009 (N_27009,N_26984,N_25314);
nand U27010 (N_27010,N_26267,N_24465);
nor U27011 (N_27011,N_26064,N_25031);
nand U27012 (N_27012,N_26879,N_25616);
nor U27013 (N_27013,N_25294,N_25346);
and U27014 (N_27014,N_26927,N_25220);
xor U27015 (N_27015,N_26668,N_26466);
nand U27016 (N_27016,N_26171,N_26727);
xor U27017 (N_27017,N_25263,N_24865);
xor U27018 (N_27018,N_24866,N_26655);
or U27019 (N_27019,N_25608,N_26045);
xnor U27020 (N_27020,N_24755,N_24619);
or U27021 (N_27021,N_26806,N_24646);
xnor U27022 (N_27022,N_24233,N_26755);
xnor U27023 (N_27023,N_24612,N_26035);
and U27024 (N_27024,N_25269,N_25325);
nor U27025 (N_27025,N_26185,N_24297);
nand U27026 (N_27026,N_24103,N_25961);
nor U27027 (N_27027,N_24329,N_24182);
xnor U27028 (N_27028,N_25898,N_25261);
nor U27029 (N_27029,N_26646,N_24027);
or U27030 (N_27030,N_24768,N_24687);
and U27031 (N_27031,N_25692,N_26248);
xnor U27032 (N_27032,N_26381,N_26872);
or U27033 (N_27033,N_25104,N_25878);
nor U27034 (N_27034,N_24758,N_26593);
nand U27035 (N_27035,N_24430,N_25929);
nor U27036 (N_27036,N_24964,N_24533);
or U27037 (N_27037,N_24169,N_26538);
or U27038 (N_27038,N_26323,N_25589);
or U27039 (N_27039,N_25297,N_24886);
nor U27040 (N_27040,N_26326,N_24741);
or U27041 (N_27041,N_26475,N_25381);
or U27042 (N_27042,N_24236,N_24834);
and U27043 (N_27043,N_26373,N_25267);
and U27044 (N_27044,N_26976,N_24561);
and U27045 (N_27045,N_25207,N_26296);
nand U27046 (N_27046,N_25135,N_26314);
nor U27047 (N_27047,N_26693,N_25422);
nor U27048 (N_27048,N_26867,N_24318);
or U27049 (N_27049,N_26262,N_24677);
nand U27050 (N_27050,N_25130,N_25392);
or U27051 (N_27051,N_26610,N_25204);
xnor U27052 (N_27052,N_24116,N_25729);
nand U27053 (N_27053,N_26745,N_26397);
or U27054 (N_27054,N_26498,N_24547);
xnor U27055 (N_27055,N_26560,N_26406);
and U27056 (N_27056,N_24067,N_25040);
xor U27057 (N_27057,N_26127,N_25775);
and U27058 (N_27058,N_25056,N_26094);
and U27059 (N_27059,N_25361,N_25860);
or U27060 (N_27060,N_24152,N_24603);
nor U27061 (N_27061,N_25415,N_25554);
nor U27062 (N_27062,N_26187,N_24501);
xor U27063 (N_27063,N_25804,N_24638);
nor U27064 (N_27064,N_24023,N_25168);
nand U27065 (N_27065,N_26584,N_25542);
nor U27066 (N_27066,N_24172,N_24678);
or U27067 (N_27067,N_26905,N_26103);
and U27068 (N_27068,N_25694,N_26989);
nor U27069 (N_27069,N_25720,N_24796);
or U27070 (N_27070,N_24367,N_26704);
nor U27071 (N_27071,N_25476,N_26821);
nor U27072 (N_27072,N_26369,N_24826);
or U27073 (N_27073,N_24380,N_26735);
xnor U27074 (N_27074,N_26391,N_26939);
xor U27075 (N_27075,N_24611,N_24939);
nor U27076 (N_27076,N_26473,N_26677);
xor U27077 (N_27077,N_24061,N_25285);
xor U27078 (N_27078,N_25217,N_26804);
nand U27079 (N_27079,N_24774,N_25625);
and U27080 (N_27080,N_25763,N_26513);
xor U27081 (N_27081,N_24994,N_26639);
nor U27082 (N_27082,N_25592,N_24969);
or U27083 (N_27083,N_25344,N_25805);
xnor U27084 (N_27084,N_26069,N_25103);
nor U27085 (N_27085,N_24594,N_25971);
and U27086 (N_27086,N_24225,N_24180);
nor U27087 (N_27087,N_26449,N_25477);
xnor U27088 (N_27088,N_26364,N_26095);
nand U27089 (N_27089,N_26000,N_25189);
nor U27090 (N_27090,N_25844,N_26889);
and U27091 (N_27091,N_25219,N_24833);
nand U27092 (N_27092,N_25052,N_25364);
or U27093 (N_27093,N_25824,N_25367);
nor U27094 (N_27094,N_24398,N_24753);
or U27095 (N_27095,N_26793,N_24406);
or U27096 (N_27096,N_25153,N_25270);
or U27097 (N_27097,N_25790,N_26047);
nor U27098 (N_27098,N_26058,N_24376);
or U27099 (N_27099,N_24953,N_26025);
xnor U27100 (N_27100,N_24874,N_26690);
or U27101 (N_27101,N_26268,N_26149);
nand U27102 (N_27102,N_24066,N_25850);
and U27103 (N_27103,N_26606,N_26215);
xnor U27104 (N_27104,N_24975,N_24275);
nor U27105 (N_27105,N_26293,N_24720);
and U27106 (N_27106,N_24078,N_24106);
and U27107 (N_27107,N_24876,N_24868);
and U27108 (N_27108,N_24676,N_26730);
nor U27109 (N_27109,N_25619,N_26828);
xnor U27110 (N_27110,N_26357,N_26178);
or U27111 (N_27111,N_25107,N_25590);
nor U27112 (N_27112,N_26835,N_25760);
nand U27113 (N_27113,N_26315,N_26535);
and U27114 (N_27114,N_26600,N_25308);
and U27115 (N_27115,N_26067,N_26131);
or U27116 (N_27116,N_24656,N_26908);
xnor U27117 (N_27117,N_26285,N_24602);
and U27118 (N_27118,N_25584,N_25461);
xnor U27119 (N_27119,N_25491,N_25252);
or U27120 (N_27120,N_26403,N_26141);
and U27121 (N_27121,N_26348,N_24524);
and U27122 (N_27122,N_25093,N_26533);
and U27123 (N_27123,N_25456,N_25497);
nor U27124 (N_27124,N_24527,N_24265);
xor U27125 (N_27125,N_26492,N_24852);
nand U27126 (N_27126,N_24914,N_25813);
or U27127 (N_27127,N_25397,N_24467);
nand U27128 (N_27128,N_26532,N_25530);
and U27129 (N_27129,N_25567,N_24862);
or U27130 (N_27130,N_24728,N_24962);
and U27131 (N_27131,N_24489,N_24884);
xnor U27132 (N_27132,N_24610,N_25845);
nand U27133 (N_27133,N_26517,N_26259);
and U27134 (N_27134,N_26374,N_24186);
nor U27135 (N_27135,N_26156,N_25597);
and U27136 (N_27136,N_25051,N_26590);
and U27137 (N_27137,N_24437,N_24118);
nand U27138 (N_27138,N_24498,N_25280);
or U27139 (N_27139,N_26265,N_25287);
nor U27140 (N_27140,N_24452,N_25934);
or U27141 (N_27141,N_25890,N_26561);
nand U27142 (N_27142,N_26522,N_26436);
or U27143 (N_27143,N_25849,N_25469);
nor U27144 (N_27144,N_26578,N_26910);
and U27145 (N_27145,N_25770,N_26702);
and U27146 (N_27146,N_25740,N_26394);
nand U27147 (N_27147,N_24268,N_26765);
nor U27148 (N_27148,N_25241,N_25444);
or U27149 (N_27149,N_26799,N_24967);
or U27150 (N_27150,N_25336,N_24449);
or U27151 (N_27151,N_26551,N_26651);
nand U27152 (N_27152,N_25539,N_26950);
nor U27153 (N_27153,N_25666,N_24827);
xor U27154 (N_27154,N_26478,N_24840);
and U27155 (N_27155,N_25513,N_24222);
nand U27156 (N_27156,N_25631,N_26206);
nand U27157 (N_27157,N_24509,N_25575);
xnor U27158 (N_27158,N_25018,N_25895);
nor U27159 (N_27159,N_25232,N_24421);
or U27160 (N_27160,N_26949,N_26153);
and U27161 (N_27161,N_26916,N_26240);
or U27162 (N_27162,N_26819,N_25678);
nor U27163 (N_27163,N_25416,N_26662);
and U27164 (N_27164,N_24651,N_26831);
nor U27165 (N_27165,N_26633,N_26113);
nor U27166 (N_27166,N_24335,N_24490);
or U27167 (N_27167,N_24856,N_26219);
nor U27168 (N_27168,N_24013,N_25441);
xnor U27169 (N_27169,N_24574,N_24998);
xor U27170 (N_27170,N_26115,N_26712);
and U27171 (N_27171,N_24719,N_25266);
and U27172 (N_27172,N_25195,N_25281);
or U27173 (N_27173,N_25496,N_26506);
or U27174 (N_27174,N_24385,N_25810);
nand U27175 (N_27175,N_25739,N_24143);
and U27176 (N_27176,N_26818,N_25467);
nor U27177 (N_27177,N_25015,N_25373);
and U27178 (N_27178,N_26987,N_26553);
nor U27179 (N_27179,N_25029,N_24581);
or U27180 (N_27180,N_26824,N_26812);
and U27181 (N_27181,N_26965,N_24521);
nor U27182 (N_27182,N_24842,N_26907);
or U27183 (N_27183,N_25774,N_25809);
and U27184 (N_27184,N_25648,N_26895);
nor U27185 (N_27185,N_26981,N_25889);
nor U27186 (N_27186,N_26698,N_26866);
nand U27187 (N_27187,N_24759,N_26004);
nor U27188 (N_27188,N_26980,N_24871);
nor U27189 (N_27189,N_26174,N_26050);
nand U27190 (N_27190,N_24054,N_25600);
or U27191 (N_27191,N_24185,N_24160);
or U27192 (N_27192,N_24889,N_25348);
or U27193 (N_27193,N_26195,N_26288);
and U27194 (N_27194,N_24260,N_25559);
and U27195 (N_27195,N_26468,N_25134);
nor U27196 (N_27196,N_26795,N_26245);
xnor U27197 (N_27197,N_25372,N_26645);
xor U27198 (N_27198,N_24294,N_25613);
nand U27199 (N_27199,N_24822,N_25533);
nor U27200 (N_27200,N_24418,N_26112);
and U27201 (N_27201,N_25026,N_24769);
or U27202 (N_27202,N_26182,N_24203);
nand U27203 (N_27203,N_26597,N_24691);
or U27204 (N_27204,N_25827,N_25665);
nand U27205 (N_27205,N_26502,N_26827);
and U27206 (N_27206,N_24530,N_26362);
or U27207 (N_27207,N_25927,N_25120);
or U27208 (N_27208,N_24256,N_25393);
nand U27209 (N_27209,N_24906,N_24276);
and U27210 (N_27210,N_25187,N_26400);
or U27211 (N_27211,N_24861,N_26294);
nor U27212 (N_27212,N_25701,N_25924);
nand U27213 (N_27213,N_24240,N_26258);
xnor U27214 (N_27214,N_26343,N_24767);
nor U27215 (N_27215,N_24466,N_26683);
and U27216 (N_27216,N_25744,N_24790);
nor U27217 (N_27217,N_25198,N_24754);
xnor U27218 (N_27218,N_25106,N_24316);
xor U27219 (N_27219,N_24352,N_26931);
or U27220 (N_27220,N_26539,N_25888);
nor U27221 (N_27221,N_24776,N_24872);
nor U27222 (N_27222,N_26587,N_25815);
or U27223 (N_27223,N_24712,N_25464);
nand U27224 (N_27224,N_25006,N_24613);
and U27225 (N_27225,N_24296,N_24600);
nor U27226 (N_27226,N_24785,N_25011);
nor U27227 (N_27227,N_24420,N_24151);
or U27228 (N_27228,N_24623,N_25875);
or U27229 (N_27229,N_24925,N_24694);
nand U27230 (N_27230,N_26752,N_26233);
nand U27231 (N_27231,N_26536,N_25264);
nand U27232 (N_27232,N_24804,N_24496);
nand U27233 (N_27233,N_25487,N_25736);
nand U27234 (N_27234,N_24844,N_26380);
nand U27235 (N_27235,N_25150,N_25330);
nor U27236 (N_27236,N_25038,N_24371);
and U27237 (N_27237,N_25795,N_25622);
or U27238 (N_27238,N_26673,N_24351);
nand U27239 (N_27239,N_25812,N_26464);
nor U27240 (N_27240,N_25765,N_26163);
nand U27241 (N_27241,N_26179,N_24596);
or U27242 (N_27242,N_25118,N_24556);
xnor U27243 (N_27243,N_25033,N_25941);
nor U27244 (N_27244,N_26969,N_25494);
nor U27245 (N_27245,N_26516,N_24681);
or U27246 (N_27246,N_24789,N_26272);
nor U27247 (N_27247,N_26985,N_26589);
or U27248 (N_27248,N_25398,N_26221);
and U27249 (N_27249,N_26658,N_25645);
and U27250 (N_27250,N_26802,N_26604);
and U27251 (N_27251,N_25425,N_24113);
nand U27252 (N_27252,N_25377,N_26452);
nor U27253 (N_27253,N_25829,N_26845);
and U27254 (N_27254,N_26720,N_26148);
or U27255 (N_27255,N_24654,N_24551);
and U27256 (N_27256,N_26780,N_25798);
and U27257 (N_27257,N_24303,N_26489);
nand U27258 (N_27258,N_26279,N_24735);
or U27259 (N_27259,N_24693,N_25615);
nand U27260 (N_27260,N_25843,N_25483);
xnor U27261 (N_27261,N_26086,N_24195);
xnor U27262 (N_27262,N_25136,N_26722);
xnor U27263 (N_27263,N_25349,N_24104);
nand U27264 (N_27264,N_26507,N_26911);
and U27265 (N_27265,N_25634,N_25831);
nor U27266 (N_27266,N_26302,N_25089);
or U27267 (N_27267,N_26244,N_26543);
nor U27268 (N_27268,N_24554,N_25638);
and U27269 (N_27269,N_25112,N_25288);
and U27270 (N_27270,N_26569,N_26859);
or U27271 (N_27271,N_26942,N_25839);
and U27272 (N_27272,N_24636,N_26978);
nor U27273 (N_27273,N_25506,N_26929);
nor U27274 (N_27274,N_26694,N_26437);
nand U27275 (N_27275,N_26881,N_25711);
nand U27276 (N_27276,N_25920,N_24081);
or U27277 (N_27277,N_24570,N_25655);
and U27278 (N_27278,N_25556,N_25585);
xor U27279 (N_27279,N_26959,N_24954);
xnor U27280 (N_27280,N_26143,N_24518);
nand U27281 (N_27281,N_26986,N_26723);
nor U27282 (N_27282,N_24491,N_26497);
nand U27283 (N_27283,N_24716,N_24389);
xor U27284 (N_27284,N_24823,N_25328);
or U27285 (N_27285,N_25432,N_24536);
xnor U27286 (N_27286,N_25174,N_24976);
xnor U27287 (N_27287,N_24344,N_25936);
or U27288 (N_27288,N_26423,N_26708);
nand U27289 (N_27289,N_26807,N_26383);
and U27290 (N_27290,N_24053,N_26208);
nand U27291 (N_27291,N_24109,N_26764);
or U27292 (N_27292,N_26670,N_24848);
or U27293 (N_27293,N_26415,N_26736);
or U27294 (N_27294,N_26583,N_26334);
and U27295 (N_27295,N_25564,N_25001);
or U27296 (N_27296,N_25200,N_25327);
nor U27297 (N_27297,N_26659,N_26405);
xor U27298 (N_27298,N_24414,N_24133);
nor U27299 (N_27299,N_26124,N_25079);
or U27300 (N_27300,N_25909,N_26260);
or U27301 (N_27301,N_26384,N_24407);
xor U27302 (N_27302,N_26499,N_26038);
or U27303 (N_27303,N_24230,N_26619);
and U27304 (N_27304,N_26572,N_25523);
xor U27305 (N_27305,N_24448,N_25743);
and U27306 (N_27306,N_25532,N_24734);
nor U27307 (N_27307,N_24892,N_24704);
nand U27308 (N_27308,N_24269,N_26085);
nand U27309 (N_27309,N_24419,N_24773);
xor U27310 (N_27310,N_26176,N_24908);
nand U27311 (N_27311,N_24640,N_24642);
or U27312 (N_27312,N_25566,N_26170);
and U27313 (N_27313,N_26559,N_26070);
or U27314 (N_27314,N_24922,N_25166);
or U27315 (N_27315,N_24122,N_26919);
or U27316 (N_27316,N_25529,N_26494);
and U27317 (N_27317,N_25660,N_26505);
xnor U27318 (N_27318,N_25054,N_25379);
nor U27319 (N_27319,N_26836,N_24077);
xor U27320 (N_27320,N_26453,N_25642);
nor U27321 (N_27321,N_25209,N_26283);
nand U27322 (N_27322,N_25549,N_24913);
nand U27323 (N_27323,N_24666,N_24107);
xor U27324 (N_27324,N_25562,N_26579);
and U27325 (N_27325,N_24632,N_26351);
nand U27326 (N_27326,N_25338,N_26335);
and U27327 (N_27327,N_25593,N_26853);
xnor U27328 (N_27328,N_25687,N_24340);
or U27329 (N_27329,N_24038,N_26940);
and U27330 (N_27330,N_26700,N_25250);
nor U27331 (N_27331,N_26422,N_25706);
xor U27332 (N_27332,N_26042,N_24427);
and U27333 (N_27333,N_24628,N_24927);
and U27334 (N_27334,N_24806,N_24679);
xor U27335 (N_27335,N_24438,N_24464);
xor U27336 (N_27336,N_25061,N_26515);
and U27337 (N_27337,N_25108,N_26665);
xnor U27338 (N_27338,N_26225,N_25742);
and U27339 (N_27339,N_24382,N_25356);
or U27340 (N_27340,N_25696,N_24586);
nand U27341 (N_27341,N_24960,N_24649);
or U27342 (N_27342,N_25408,N_26734);
nor U27343 (N_27343,N_26439,N_26988);
nor U27344 (N_27344,N_25997,N_25389);
nor U27345 (N_27345,N_25673,N_26331);
or U27346 (N_27346,N_26903,N_26669);
or U27347 (N_27347,N_25251,N_25350);
or U27348 (N_27348,N_25465,N_25173);
xor U27349 (N_27349,N_24481,N_25842);
or U27350 (N_27350,N_26483,N_26787);
nand U27351 (N_27351,N_24912,N_26923);
and U27352 (N_27352,N_25664,N_25859);
and U27353 (N_27353,N_25921,N_26558);
nand U27354 (N_27354,N_24685,N_26706);
or U27355 (N_27355,N_25414,N_26541);
nor U27356 (N_27356,N_26459,N_25904);
or U27357 (N_27357,N_24086,N_26231);
nand U27358 (N_27358,N_24144,N_26705);
or U27359 (N_27359,N_24963,N_25947);
or U27360 (N_27360,N_26714,N_26945);
xor U27361 (N_27361,N_25587,N_24929);
xor U27362 (N_27362,N_24949,N_24919);
nor U27363 (N_27363,N_26242,N_25175);
or U27364 (N_27364,N_26748,N_25682);
xor U27365 (N_27365,N_24224,N_26834);
xor U27366 (N_27366,N_24319,N_25574);
or U27367 (N_27367,N_25916,N_26072);
nor U27368 (N_27368,N_26717,N_26904);
nand U27369 (N_27369,N_24950,N_26556);
nor U27370 (N_27370,N_26060,N_24161);
or U27371 (N_27371,N_25899,N_24812);
and U27372 (N_27372,N_25658,N_26462);
nor U27373 (N_27373,N_24641,N_25881);
and U27374 (N_27374,N_24644,N_25957);
nand U27375 (N_27375,N_25675,N_26966);
xor U27376 (N_27376,N_24620,N_24342);
nand U27377 (N_27377,N_24933,N_25272);
and U27378 (N_27378,N_25866,N_26421);
and U27379 (N_27379,N_26068,N_24097);
xor U27380 (N_27380,N_25403,N_24119);
nand U27381 (N_27381,N_26382,N_24936);
and U27382 (N_27382,N_25894,N_24718);
nor U27383 (N_27383,N_24601,N_25647);
nor U27384 (N_27384,N_25090,N_25546);
or U27385 (N_27385,N_25311,N_24267);
or U27386 (N_27386,N_24932,N_26774);
or U27387 (N_27387,N_24005,N_24670);
xor U27388 (N_27388,N_24567,N_24058);
and U27389 (N_27389,N_26571,N_26001);
nand U27390 (N_27390,N_24955,N_26210);
xor U27391 (N_27391,N_24791,N_24274);
and U27392 (N_27392,N_26059,N_25299);
xor U27393 (N_27393,N_25950,N_26740);
xnor U27394 (N_27394,N_24880,N_25213);
nor U27395 (N_27395,N_25792,N_25560);
nand U27396 (N_27396,N_24473,N_26295);
xnor U27397 (N_27397,N_26278,N_26598);
and U27398 (N_27398,N_24346,N_25139);
xor U27399 (N_27399,N_26350,N_26183);
or U27400 (N_27400,N_25510,N_26345);
or U27401 (N_27401,N_26220,N_24887);
nor U27402 (N_27402,N_24614,N_24637);
and U27403 (N_27403,N_25826,N_25194);
and U27404 (N_27404,N_26239,N_26692);
nand U27405 (N_27405,N_24504,N_26425);
and U27406 (N_27406,N_24703,N_25707);
and U27407 (N_27407,N_25224,N_24458);
or U27408 (N_27408,N_25309,N_24343);
xnor U27409 (N_27409,N_26349,N_26729);
or U27410 (N_27410,N_24037,N_24742);
and U27411 (N_27411,N_24212,N_24511);
nor U27412 (N_27412,N_25265,N_26914);
and U27413 (N_27413,N_26671,N_26953);
nor U27414 (N_27414,N_25502,N_26896);
xor U27415 (N_27415,N_25003,N_25872);
nor U27416 (N_27416,N_26631,N_24502);
nand U27417 (N_27417,N_24423,N_25643);
or U27418 (N_27418,N_26249,N_25363);
nand U27419 (N_27419,N_26891,N_24049);
or U27420 (N_27420,N_24453,N_24621);
nor U27421 (N_27421,N_24141,N_26749);
or U27422 (N_27422,N_25715,N_24746);
nor U27423 (N_27423,N_24065,N_24813);
xor U27424 (N_27424,N_25146,N_24470);
nor U27425 (N_27425,N_25479,N_24966);
nor U27426 (N_27426,N_24055,N_25390);
nor U27427 (N_27427,N_26932,N_25065);
xor U27428 (N_27428,N_25965,N_26681);
and U27429 (N_27429,N_26746,N_24948);
and U27430 (N_27430,N_25953,N_24270);
and U27431 (N_27431,N_26254,N_24545);
or U27432 (N_27432,N_26618,N_24337);
nor U27433 (N_27433,N_24730,N_24991);
nand U27434 (N_27434,N_25069,N_24043);
or U27435 (N_27435,N_24731,N_26300);
nand U27436 (N_27436,N_24845,N_24593);
nand U27437 (N_27437,N_25749,N_24263);
and U27438 (N_27438,N_26758,N_25588);
nand U27439 (N_27439,N_25852,N_25596);
xor U27440 (N_27440,N_24497,N_26679);
or U27441 (N_27441,N_26622,N_24197);
nand U27442 (N_27442,N_25395,N_26562);
or U27443 (N_27443,N_24618,N_25837);
nand U27444 (N_27444,N_25557,N_24830);
or U27445 (N_27445,N_25717,N_25055);
nor U27446 (N_27446,N_25923,N_26075);
xnor U27447 (N_27447,N_24246,N_25925);
and U27448 (N_27448,N_26930,N_26743);
and U27449 (N_27449,N_25536,N_24885);
xor U27450 (N_27450,N_26341,N_25334);
and U27451 (N_27451,N_26395,N_24129);
nand U27452 (N_27452,N_26031,N_24553);
or U27453 (N_27453,N_25507,N_24974);
or U27454 (N_27454,N_26119,N_26956);
nand U27455 (N_27455,N_25084,N_24176);
or U27456 (N_27456,N_25360,N_25745);
xnor U27457 (N_27457,N_25131,N_24445);
xnor U27458 (N_27458,N_26408,N_24820);
or U27459 (N_27459,N_25607,N_24859);
or U27460 (N_27460,N_25229,N_26125);
nand U27461 (N_27461,N_24870,N_24609);
xor U27462 (N_27462,N_24354,N_24305);
nor U27463 (N_27463,N_24643,N_26299);
and U27464 (N_27464,N_24639,N_25324);
xnor U27465 (N_27465,N_24391,N_26592);
or U27466 (N_27466,N_26892,N_25172);
or U27467 (N_27467,N_25214,N_25448);
or U27468 (N_27468,N_26656,N_24474);
nand U27469 (N_27469,N_25595,N_26747);
nor U27470 (N_27470,N_25092,N_26194);
or U27471 (N_27471,N_24818,N_26641);
xor U27472 (N_27472,N_26709,N_24672);
and U27473 (N_27473,N_26992,N_25887);
nand U27474 (N_27474,N_25042,N_25782);
xnor U27475 (N_27475,N_26108,N_26634);
nor U27476 (N_27476,N_25970,N_24523);
nand U27477 (N_27477,N_25238,N_24214);
and U27478 (N_27478,N_24472,N_24431);
nand U27479 (N_27479,N_25010,N_25186);
nand U27480 (N_27480,N_26317,N_26771);
nand U27481 (N_27481,N_24934,N_24108);
nand U27482 (N_27482,N_26401,N_26685);
or U27483 (N_27483,N_26454,N_24126);
and U27484 (N_27484,N_26833,N_26056);
nor U27485 (N_27485,N_24958,N_25504);
or U27486 (N_27486,N_26321,N_25726);
nand U27487 (N_27487,N_26570,N_24881);
and U27488 (N_27488,N_24894,N_24942);
nor U27489 (N_27489,N_26514,N_25738);
nor U27490 (N_27490,N_25439,N_26491);
nor U27491 (N_27491,N_24155,N_25591);
nand U27492 (N_27492,N_26887,N_26829);
xor U27493 (N_27493,N_24245,N_26432);
nand U27494 (N_27494,N_26797,N_26241);
or U27495 (N_27495,N_26044,N_24253);
xnor U27496 (N_27496,N_25035,N_24578);
nor U27497 (N_27497,N_26762,N_25569);
and U27498 (N_27498,N_26826,N_25544);
or U27499 (N_27499,N_26894,N_26476);
nand U27500 (N_27500,N_24543,N_24552);
xor U27501 (N_27501,N_24725,N_24189);
nor U27502 (N_27502,N_25948,N_26344);
or U27503 (N_27503,N_24447,N_26234);
nor U27504 (N_27504,N_24541,N_26277);
nor U27505 (N_27505,N_24665,N_24251);
and U27506 (N_27506,N_25180,N_25503);
and U27507 (N_27507,N_26637,N_25972);
and U27508 (N_27508,N_25190,N_24479);
nor U27509 (N_27509,N_25167,N_25621);
xnor U27510 (N_27510,N_26083,N_25672);
nor U27511 (N_27511,N_26875,N_26636);
nand U27512 (N_27512,N_26026,N_26577);
and U27513 (N_27513,N_25401,N_25988);
nand U27514 (N_27514,N_25919,N_26531);
nand U27515 (N_27515,N_25698,N_25515);
nand U27516 (N_27516,N_25735,N_25908);
or U27517 (N_27517,N_24387,N_25952);
nor U27518 (N_27518,N_24089,N_26504);
xor U27519 (N_27519,N_25024,N_25486);
nor U27520 (N_27520,N_26791,N_26145);
nand U27521 (N_27521,N_25629,N_26603);
nand U27522 (N_27522,N_24400,N_26548);
xnor U27523 (N_27523,N_25258,N_26202);
nand U27524 (N_27524,N_26608,N_24323);
xor U27525 (N_27525,N_26442,N_25677);
and U27526 (N_27526,N_26130,N_24882);
and U27527 (N_27527,N_24145,N_26189);
nand U27528 (N_27528,N_25359,N_25893);
and U27529 (N_27529,N_24436,N_24689);
xor U27530 (N_27530,N_25239,N_24358);
xor U27531 (N_27531,N_26624,N_26161);
and U27532 (N_27532,N_26664,N_24800);
nand U27533 (N_27533,N_26322,N_24215);
nor U27534 (N_27534,N_25705,N_26128);
xnor U27535 (N_27535,N_26617,N_26858);
and U27536 (N_27536,N_25342,N_24428);
xnor U27537 (N_27537,N_25047,N_26160);
or U27538 (N_27538,N_26520,N_24505);
nand U27539 (N_27539,N_25321,N_24317);
nor U27540 (N_27540,N_24223,N_25520);
or U27541 (N_27541,N_26566,N_24213);
and U27542 (N_27542,N_24984,N_26217);
nor U27543 (N_27543,N_26412,N_25446);
and U27544 (N_27544,N_25651,N_24015);
nor U27545 (N_27545,N_26667,N_25524);
and U27546 (N_27546,N_24443,N_25702);
and U27547 (N_27547,N_25212,N_24738);
xor U27548 (N_27548,N_24433,N_24048);
nand U27549 (N_27549,N_26114,N_25830);
nand U27550 (N_27550,N_25966,N_26918);
and U27551 (N_27551,N_24930,N_26154);
and U27552 (N_27552,N_25110,N_24007);
or U27553 (N_27553,N_25149,N_25602);
and U27554 (N_27554,N_24397,N_25246);
nand U27555 (N_27555,N_24020,N_26463);
nor U27556 (N_27556,N_25659,N_26544);
or U27557 (N_27557,N_26750,N_24508);
nand U27558 (N_27558,N_25746,N_26599);
nand U27559 (N_27559,N_25165,N_24658);
and U27560 (N_27560,N_26650,N_26638);
xor U27561 (N_27561,N_26991,N_25087);
nor U27562 (N_27562,N_25942,N_25979);
nor U27563 (N_27563,N_25085,N_24392);
xnor U27564 (N_27564,N_24989,N_25340);
or U27565 (N_27565,N_26785,N_24403);
nor U27566 (N_27566,N_24254,N_24999);
nand U27567 (N_27567,N_24257,N_26630);
xnor U27568 (N_27568,N_25855,N_24292);
and U27569 (N_27569,N_25159,N_24724);
xor U27570 (N_27570,N_25641,N_26184);
nand U27571 (N_27571,N_24205,N_25534);
nor U27572 (N_27572,N_26181,N_24750);
nand U27573 (N_27573,N_26777,N_24661);
or U27574 (N_27574,N_26205,N_26540);
or U27575 (N_27575,N_26198,N_25624);
and U27576 (N_27576,N_24854,N_26006);
or U27577 (N_27577,N_26446,N_24494);
and U27578 (N_27578,N_24432,N_26699);
nor U27579 (N_27579,N_24328,N_24739);
nand U27580 (N_27580,N_25780,N_25646);
nand U27581 (N_27581,N_24117,N_25183);
and U27582 (N_27582,N_24794,N_24009);
nand U27583 (N_27583,N_24817,N_26546);
or U27584 (N_27584,N_25796,N_24653);
xnor U27585 (N_27585,N_24082,N_26107);
and U27586 (N_27586,N_24749,N_25628);
or U27587 (N_27587,N_24990,N_26482);
and U27588 (N_27588,N_24850,N_25652);
nor U27589 (N_27589,N_26142,N_24307);
or U27590 (N_27590,N_26054,N_26256);
or U27591 (N_27591,N_24019,N_26393);
nand U27592 (N_27592,N_26865,N_25630);
xnor U27593 (N_27593,N_24674,N_26076);
xnor U27594 (N_27594,N_25277,N_26353);
and U27595 (N_27595,N_26716,N_25451);
nor U27596 (N_27596,N_25528,N_26954);
nand U27597 (N_27597,N_24783,N_25910);
or U27598 (N_27598,N_26055,N_25911);
nand U27599 (N_27599,N_26010,N_25365);
nand U27600 (N_27600,N_26191,N_24041);
and U27601 (N_27601,N_25984,N_25848);
nor U27602 (N_27602,N_25555,N_24532);
nor U27603 (N_27603,N_25847,N_24737);
nor U27604 (N_27604,N_26524,N_26093);
or U27605 (N_27605,N_26534,N_24171);
nor U27606 (N_27606,N_24478,N_25716);
xor U27607 (N_27607,N_26092,N_24146);
xnor U27608 (N_27608,N_25973,N_26340);
xnor U27609 (N_27609,N_24797,N_26274);
xnor U27610 (N_27610,N_26525,N_25077);
or U27611 (N_27611,N_24555,N_24560);
and U27612 (N_27612,N_26324,N_25599);
nor U27613 (N_27613,N_24896,N_24484);
xor U27614 (N_27614,N_24216,N_26620);
nor U27615 (N_27615,N_26082,N_24915);
nor U27616 (N_27616,N_26118,N_24147);
or U27617 (N_27617,N_26841,N_25436);
nor U27618 (N_27618,N_25148,N_24014);
and U27619 (N_27619,N_24190,N_24163);
and U27620 (N_27620,N_26920,N_26356);
nor U27621 (N_27621,N_26140,N_25633);
and U27622 (N_27622,N_24879,N_25109);
nand U27623 (N_27623,N_26022,N_26371);
nor U27624 (N_27624,N_26695,N_25216);
or U27625 (N_27625,N_25586,N_26573);
and U27626 (N_27626,N_25963,N_26595);
nand U27627 (N_27627,N_24604,N_26211);
xor U27628 (N_27628,N_26567,N_25306);
or U27629 (N_27629,N_25078,N_25091);
xor U27630 (N_27630,N_25757,N_24353);
nand U27631 (N_27631,N_25247,N_25192);
xnor U27632 (N_27632,N_26549,N_25059);
and U27633 (N_27633,N_24150,N_26860);
or U27634 (N_27634,N_26946,N_26438);
nand U27635 (N_27635,N_24650,N_26649);
and U27636 (N_27636,N_24517,N_26471);
nand U27637 (N_27637,N_25025,N_26810);
nand U27638 (N_27638,N_25699,N_24579);
nand U27639 (N_27639,N_24659,N_26168);
nor U27640 (N_27640,N_24682,N_25002);
or U27641 (N_27641,N_25005,N_26811);
nand U27642 (N_27642,N_24622,N_26429);
and U27643 (N_27643,N_25227,N_24379);
or U27644 (N_27644,N_24124,N_24943);
xor U27645 (N_27645,N_24313,N_24232);
xnor U27646 (N_27646,N_25044,N_25800);
and U27647 (N_27647,N_26269,N_25527);
and U27648 (N_27648,N_24137,N_24902);
or U27649 (N_27649,N_24194,N_25661);
or U27650 (N_27650,N_26696,N_25380);
or U27651 (N_27651,N_24394,N_26554);
or U27652 (N_27652,N_26311,N_26663);
or U27653 (N_27653,N_24384,N_24098);
and U27654 (N_27654,N_25351,N_24729);
nand U27655 (N_27655,N_25236,N_24935);
or U27656 (N_27656,N_25259,N_25243);
nand U27657 (N_27657,N_26313,N_24673);
xor U27658 (N_27658,N_24516,N_25097);
nor U27659 (N_27659,N_26413,N_24557);
or U27660 (N_27660,N_26805,N_24322);
xor U27661 (N_27661,N_24591,N_26838);
and U27662 (N_27662,N_25385,N_25293);
nor U27663 (N_27663,N_26922,N_25276);
or U27664 (N_27664,N_24572,N_26754);
xor U27665 (N_27665,N_25540,N_24959);
or U27666 (N_27666,N_26528,N_24064);
nand U27667 (N_27667,N_24462,N_25388);
and U27668 (N_27668,N_25598,N_25722);
xnor U27669 (N_27669,N_24634,N_25245);
nor U27670 (N_27670,N_25326,N_25996);
xor U27671 (N_27671,N_24193,N_26983);
nor U27672 (N_27672,N_25475,N_24947);
xnor U27673 (N_27673,N_24148,N_24063);
or U27674 (N_27674,N_25538,N_24805);
and U27675 (N_27675,N_25156,N_25188);
nand U27676 (N_27676,N_26943,N_25323);
and U27677 (N_27677,N_26048,N_26647);
and U27678 (N_27678,N_26510,N_25906);
xor U27679 (N_27679,N_25184,N_25472);
nor U27680 (N_27680,N_26456,N_26399);
nand U27681 (N_27681,N_24544,N_24252);
nor U27682 (N_27682,N_25828,N_26803);
nand U27683 (N_27683,N_25956,N_24429);
xor U27684 (N_27684,N_26995,N_26057);
nor U27685 (N_27685,N_24709,N_25951);
xor U27686 (N_27686,N_25164,N_25930);
nand U27687 (N_27687,N_25499,N_24520);
nand U27688 (N_27688,N_24584,N_26652);
and U27689 (N_27689,N_26721,N_26568);
nor U27690 (N_27690,N_24951,N_26366);
or U27691 (N_27691,N_25370,N_26332);
xnor U27692 (N_27692,N_25057,N_26675);
nand U27693 (N_27693,N_24751,N_25822);
xnor U27694 (N_27694,N_24334,N_25670);
xor U27695 (N_27695,N_24304,N_24016);
nor U27696 (N_27696,N_24849,N_24207);
or U27697 (N_27697,N_26273,N_25310);
or U27698 (N_27698,N_25418,N_24201);
nor U27699 (N_27699,N_24668,N_26150);
xnor U27700 (N_27700,N_24291,N_26512);
and U27701 (N_27701,N_26159,N_26760);
nand U27702 (N_27702,N_25974,N_24173);
xor U27703 (N_27703,N_24441,N_25773);
and U27704 (N_27704,N_24565,N_26602);
nand U27705 (N_27705,N_24030,N_24277);
nand U27706 (N_27706,N_26719,N_24700);
xor U27707 (N_27707,N_26862,N_26822);
and U27708 (N_27708,N_26545,N_25115);
or U27709 (N_27709,N_25723,N_26292);
or U27710 (N_27710,N_25712,N_24250);
nand U27711 (N_27711,N_25273,N_26264);
xnor U27712 (N_27712,N_24264,N_26870);
or U27713 (N_27713,N_26843,N_26960);
nor U27714 (N_27714,N_26733,N_24744);
nand U27715 (N_27715,N_24280,N_24891);
nor U27716 (N_27716,N_26015,N_26739);
nand U27717 (N_27717,N_24168,N_26337);
nor U27718 (N_27718,N_24829,N_24028);
and U27719 (N_27719,N_25147,N_24134);
nand U27720 (N_27720,N_26417,N_24564);
nor U27721 (N_27721,N_26186,N_25939);
or U27722 (N_27722,N_26238,N_26041);
nand U27723 (N_27723,N_25205,N_26065);
nand U27724 (N_27724,N_26088,N_25255);
and U27725 (N_27725,N_25201,N_24878);
xnor U27726 (N_27726,N_26697,N_26759);
nand U27727 (N_27727,N_26177,N_24309);
nor U27728 (N_27728,N_25649,N_26109);
nor U27729 (N_27729,N_26147,N_26090);
nor U27730 (N_27730,N_24615,N_24217);
xor U27731 (N_27731,N_26414,N_24924);
and U27732 (N_27732,N_24931,N_24977);
xor U27733 (N_27733,N_24012,N_25086);
and U27734 (N_27734,N_26019,N_26523);
or U27735 (N_27735,N_24229,N_26526);
or U27736 (N_27736,N_26372,N_26162);
xnor U27737 (N_27737,N_24996,N_26359);
xor U27738 (N_27738,N_24059,N_24952);
and U27739 (N_27739,N_24779,N_26416);
or U27740 (N_27740,N_25801,N_24191);
xnor U27741 (N_27741,N_25305,N_25318);
nand U27742 (N_27742,N_25857,N_25685);
nor U27743 (N_27743,N_24799,N_24200);
nand U27744 (N_27744,N_24981,N_25821);
or U27745 (N_27745,N_25867,N_24522);
and U27746 (N_27746,N_26715,N_25485);
and U27747 (N_27747,N_25834,N_25298);
nand U27748 (N_27748,N_26033,N_25714);
xor U27749 (N_27749,N_25222,N_26342);
or U27750 (N_27750,N_24372,N_24624);
nor U27751 (N_27751,N_26761,N_24390);
xnor U27752 (N_27752,N_25606,N_25283);
xnor U27753 (N_27753,N_24219,N_24945);
or U27754 (N_27754,N_25337,N_25656);
or U27755 (N_27755,N_24310,N_24788);
nor U27756 (N_27756,N_26365,N_25880);
xnor U27757 (N_27757,N_24425,N_26654);
and U27758 (N_27758,N_25786,N_24732);
nand U27759 (N_27759,N_25407,N_26358);
nand U27760 (N_27760,N_26855,N_25231);
and U27761 (N_27761,N_24595,N_25041);
and U27762 (N_27762,N_26770,N_24388);
nand U27763 (N_27763,N_24941,N_24153);
nor U27764 (N_27764,N_26973,N_26596);
nand U27765 (N_27765,N_26643,N_25064);
xnor U27766 (N_27766,N_25319,N_24542);
nand U27767 (N_27767,N_26888,N_24839);
and U27768 (N_27768,N_24784,N_25278);
or U27769 (N_27769,N_25522,N_24426);
nand U27770 (N_27770,N_25873,N_26846);
or U27771 (N_27771,N_26435,N_26947);
nor U27772 (N_27772,N_25353,N_26757);
nor U27773 (N_27773,N_24743,N_25060);
nand U27774 (N_27774,N_26110,N_26053);
nor U27775 (N_27775,N_26247,N_25579);
nand U27776 (N_27776,N_25937,N_25181);
nand U27777 (N_27777,N_26199,N_25955);
nand U27778 (N_27778,N_24393,N_24076);
xor U27779 (N_27779,N_24286,N_24987);
xor U27780 (N_27780,N_25650,N_25823);
nand U27781 (N_27781,N_24831,N_25358);
and U27782 (N_27782,N_24548,N_26360);
nor U27783 (N_27783,N_24079,N_25151);
and U27784 (N_27784,N_24910,N_25371);
nor U27785 (N_27785,N_25940,N_25237);
or U27786 (N_27786,N_24515,N_24378);
nand U27787 (N_27787,N_26557,N_25732);
nor U27788 (N_27788,N_25653,N_24285);
xor U27789 (N_27789,N_24460,N_26298);
xor U27790 (N_27790,N_25676,N_26925);
xor U27791 (N_27791,N_25179,N_26433);
xnor U27792 (N_27792,N_24373,N_26580);
or U27793 (N_27793,N_26227,N_25289);
or U27794 (N_27794,N_24052,N_24451);
and U27795 (N_27795,N_24381,N_25526);
and U27796 (N_27796,N_25450,N_25074);
or U27797 (N_27797,N_24302,N_25978);
xnor U27798 (N_27798,N_24539,N_25405);
nand U27799 (N_27799,N_26591,N_25819);
or U27800 (N_27800,N_25113,N_24782);
nand U27801 (N_27801,N_24444,N_25603);
xor U27802 (N_27802,N_26542,N_25071);
xor U27803 (N_27803,N_26825,N_25787);
nor U27804 (N_27804,N_26967,N_25945);
xnor U27805 (N_27805,N_26842,N_25474);
xnor U27806 (N_27806,N_26301,N_24034);
or U27807 (N_27807,N_26628,N_26601);
or U27808 (N_27808,N_26338,N_24244);
nor U27809 (N_27809,N_24809,N_25463);
xnor U27810 (N_27810,N_24100,N_26271);
nor U27811 (N_27811,N_26009,N_25161);
nor U27812 (N_27812,N_26120,N_26451);
nor U27813 (N_27813,N_24417,N_25462);
xor U27814 (N_27814,N_26607,N_24875);
nor U27815 (N_27815,N_26229,N_26613);
nand U27816 (N_27816,N_24660,N_24370);
or U27817 (N_27817,N_25954,N_25982);
nor U27818 (N_27818,N_24279,N_24781);
nor U27819 (N_27819,N_24811,N_24711);
nor U27820 (N_27820,N_24476,N_24587);
and U27821 (N_27821,N_26962,N_26347);
and U27822 (N_27822,N_24863,N_25689);
xnor U27823 (N_27823,N_24972,N_24904);
nor U27824 (N_27824,N_26495,N_26798);
nor U27825 (N_27825,N_25012,N_25411);
or U27826 (N_27826,N_26355,N_24795);
nor U27827 (N_27827,N_24956,N_24582);
xor U27828 (N_27828,N_26688,N_25437);
nand U27829 (N_27829,N_26710,N_25840);
and U27830 (N_27830,N_26850,N_24858);
or U27831 (N_27831,N_24123,N_26460);
xnor U27832 (N_27832,N_26594,N_24778);
xor U27833 (N_27833,N_25838,N_24938);
nor U27834 (N_27834,N_25021,N_26005);
nand U27835 (N_27835,N_25803,N_24736);
nor U27836 (N_27836,N_25695,N_24860);
nand U27837 (N_27837,N_24184,N_24228);
or U27838 (N_27838,N_24940,N_26135);
or U27839 (N_27839,N_26672,N_25731);
or U27840 (N_27840,N_25482,N_25576);
and U27841 (N_27841,N_26472,N_26073);
nor U27842 (N_27842,N_26325,N_24290);
or U27843 (N_27843,N_24071,N_26100);
nand U27844 (N_27844,N_25976,N_24320);
or U27845 (N_27845,N_26530,N_25088);
nor U27846 (N_27846,N_24971,N_26409);
nor U27847 (N_27847,N_24456,N_25864);
and U27848 (N_27848,N_26290,N_25058);
nand U27849 (N_27849,N_25424,N_24748);
nand U27850 (N_27850,N_25295,N_26678);
nand U27851 (N_27851,N_24590,N_24401);
nor U27852 (N_27852,N_26832,N_25291);
xor U27853 (N_27853,N_26096,N_25396);
and U27854 (N_27854,N_25654,N_25578);
nor U27855 (N_27855,N_24455,N_24271);
xor U27856 (N_27856,N_24042,N_25045);
nor U27857 (N_27857,N_26447,N_26284);
xnor U27858 (N_27858,N_25443,N_24810);
and U27859 (N_27859,N_26255,N_25686);
xor U27860 (N_27860,N_26640,N_26982);
or U27861 (N_27861,N_24625,N_24440);
and U27862 (N_27862,N_26040,N_25032);
nor U27863 (N_27863,N_25962,N_25755);
nand U27864 (N_27864,N_24110,N_24816);
nor U27865 (N_27865,N_26854,N_24488);
or U27866 (N_27866,N_26139,N_25868);
nor U27867 (N_27867,N_25421,N_25897);
xnor U27868 (N_27868,N_26329,N_25883);
and U27869 (N_27869,N_25680,N_24159);
or U27870 (N_27870,N_25037,N_26392);
nor U27871 (N_27871,N_24857,N_26781);
or U27872 (N_27872,N_26291,N_24662);
and U27873 (N_27873,N_24434,N_26511);
nor U27874 (N_27874,N_24916,N_26648);
nand U27875 (N_27875,N_24004,N_24339);
nor U27876 (N_27876,N_26964,N_26111);
nor U27877 (N_27877,N_25027,N_25697);
nand U27878 (N_27878,N_26848,N_25891);
xor U27879 (N_27879,N_25573,N_24763);
and U27880 (N_27880,N_24695,N_25143);
and U27881 (N_27881,N_24836,N_25007);
or U27882 (N_27882,N_24979,N_26496);
nor U27883 (N_27883,N_24627,N_25402);
nand U27884 (N_27884,N_24368,N_26467);
and U27885 (N_27885,N_25902,N_25674);
and U27886 (N_27886,N_24792,N_26420);
xor U27887 (N_27887,N_26212,N_26087);
and U27888 (N_27888,N_26955,N_24786);
xnor U27889 (N_27889,N_24366,N_25457);
xnor U27890 (N_27890,N_26327,N_26155);
nand U27891 (N_27891,N_26527,N_24926);
nand U27892 (N_27892,N_25818,N_24588);
and U27893 (N_27893,N_25171,N_24529);
or U27894 (N_27894,N_24550,N_25944);
or U27895 (N_27895,N_26201,N_26014);
nand U27896 (N_27896,N_24121,N_25879);
nand U27897 (N_27897,N_24068,N_24179);
or U27898 (N_27898,N_24350,N_25082);
nand U27899 (N_27899,N_25999,N_26144);
and U27900 (N_27900,N_26305,N_26479);
and U27901 (N_27901,N_24035,N_25387);
or U27902 (N_27902,N_25604,N_26232);
nand U27903 (N_27903,N_26487,N_25301);
xor U27904 (N_27904,N_24825,N_25121);
or U27905 (N_27905,N_25154,N_26703);
or U27906 (N_27906,N_24566,N_25249);
nand U27907 (N_27907,N_26691,N_24088);
nor U27908 (N_27908,N_26501,N_24714);
and U27909 (N_27909,N_25394,N_24242);
or U27910 (N_27910,N_24721,N_26844);
and U27911 (N_27911,N_25413,N_26078);
or U27912 (N_27912,N_24598,N_24487);
xnor U27913 (N_27913,N_25820,N_25772);
or U27914 (N_27914,N_24355,N_26051);
xnor U27915 (N_27915,N_25116,N_25230);
or U27916 (N_27916,N_26081,N_26316);
or U27917 (N_27917,N_26856,N_24558);
or U27918 (N_27918,N_26032,N_25419);
xor U27919 (N_27919,N_26661,N_25105);
nand U27920 (N_27920,N_25671,N_24503);
xor U27921 (N_27921,N_26897,N_26623);
or U27922 (N_27922,N_24918,N_24512);
or U27923 (N_27923,N_25098,N_25335);
or U27924 (N_27924,N_24761,N_24821);
xor U27925 (N_27925,N_24321,N_26857);
or U27926 (N_27926,N_26431,N_25282);
nand U27927 (N_27927,N_24568,N_24300);
xor U27928 (N_27928,N_24306,N_26612);
nor U27929 (N_27929,N_24690,N_24301);
nand U27930 (N_27930,N_25374,N_25133);
xnor U27931 (N_27931,N_26237,N_24299);
or U27932 (N_27932,N_25748,N_24697);
nor U27933 (N_27933,N_24204,N_24033);
nand U27934 (N_27934,N_25771,N_26071);
nand U27935 (N_27935,N_25417,N_26814);
or U27936 (N_27936,N_24630,N_26105);
nand U27937 (N_27937,N_25609,N_24362);
or U27938 (N_27938,N_26952,N_26726);
nor U27939 (N_27939,N_24177,N_26310);
and U27940 (N_27940,N_24995,N_24506);
nand U27941 (N_27941,N_24136,N_25558);
xnor U27942 (N_27942,N_26099,N_25663);
or U27943 (N_27943,N_24101,N_24835);
nor U27944 (N_27944,N_26368,N_26158);
nor U27945 (N_27945,N_26609,N_25501);
and U27946 (N_27946,N_24261,N_26097);
xnor U27947 (N_27947,N_26427,N_26008);
xnor U27948 (N_27948,N_24766,N_25583);
nand U27949 (N_27949,N_25981,N_24413);
nor U27950 (N_27950,N_25753,N_26074);
nor U27951 (N_27951,N_26027,N_26352);
nor U27952 (N_27952,N_26893,N_25315);
and U27953 (N_27953,N_26133,N_25762);
and U27954 (N_27954,N_26089,N_25892);
nand U27955 (N_27955,N_24315,N_24583);
or U27956 (N_27956,N_26402,N_25049);
nor U27957 (N_27957,N_24284,N_26077);
nand U27958 (N_27958,N_24569,N_25741);
xor U27959 (N_27959,N_24288,N_25455);
xor U27960 (N_27960,N_24493,N_25623);
nor U27961 (N_27961,N_26934,N_25582);
nor U27962 (N_27962,N_25612,N_25008);
and U27963 (N_27963,N_25215,N_25547);
and U27964 (N_27964,N_26419,N_26063);
or U27965 (N_27965,N_26635,N_24412);
and U27966 (N_27966,N_24699,N_25233);
or U27967 (N_27967,N_24198,N_25357);
and U27968 (N_27968,N_25070,N_25508);
or U27969 (N_27969,N_25332,N_24605);
xor U27970 (N_27970,N_24968,N_24514);
xor U27971 (N_27971,N_24127,N_26968);
and U27972 (N_27972,N_24648,N_24780);
nand U27973 (N_27973,N_24698,N_25111);
nor U27974 (N_27974,N_25196,N_24001);
xor U27975 (N_27975,N_24010,N_25493);
nor U27976 (N_27976,N_26386,N_24469);
xor U27977 (N_27977,N_24073,N_25449);
xnor U27978 (N_27978,N_26246,N_24111);
nand U27979 (N_27979,N_25856,N_24683);
or U27980 (N_27980,N_24409,N_25915);
nand U27981 (N_27981,N_26621,N_26485);
or U27982 (N_27982,N_24900,N_26666);
xnor U27983 (N_27983,N_24114,N_25203);
nor U27984 (N_27984,N_24471,N_24897);
nor U27985 (N_27985,N_24283,N_26304);
and U27986 (N_27986,N_25570,N_24580);
nor U27987 (N_27987,N_26164,N_25072);
nand U27988 (N_27988,N_25811,N_24446);
xor U27989 (N_27989,N_24314,N_26333);
and U27990 (N_27990,N_24247,N_25490);
or U27991 (N_27991,N_24752,N_26794);
xnor U27992 (N_27992,N_26957,N_25050);
nand U27993 (N_27993,N_24036,N_24680);
xnor U27994 (N_27994,N_24105,N_25257);
and U27995 (N_27995,N_24166,N_25481);
and U27996 (N_27996,N_25935,N_26029);
and U27997 (N_27997,N_25468,N_24702);
and U27998 (N_27998,N_26230,N_26555);
nand U27999 (N_27999,N_25752,N_25100);
nor U28000 (N_28000,N_24597,N_24327);
or U28001 (N_28001,N_26167,N_26574);
or U28002 (N_28002,N_25053,N_24843);
nand U28003 (N_28003,N_26477,N_24332);
or U28004 (N_28004,N_25572,N_24492);
xor U28005 (N_28005,N_26303,N_24227);
or U28006 (N_28006,N_24396,N_24404);
xor U28007 (N_28007,N_24895,N_24824);
nor U28008 (N_28008,N_24911,N_24909);
and U28009 (N_28009,N_25862,N_24347);
and U28010 (N_28010,N_26994,N_25635);
nand U28011 (N_28011,N_25794,N_26687);
xnor U28012 (N_28012,N_25152,N_25733);
and U28013 (N_28013,N_24486,N_24083);
nor U28014 (N_28014,N_25958,N_24360);
xor U28015 (N_28015,N_24312,N_25704);
nor U28016 (N_28016,N_26900,N_24298);
and U28017 (N_28017,N_25129,N_24798);
nor U28018 (N_28018,N_25498,N_26565);
or U28019 (N_28019,N_26684,N_26784);
xor U28020 (N_28020,N_26913,N_26307);
and U28021 (N_28021,N_24510,N_24424);
xor U28022 (N_28022,N_26280,N_25096);
or U28023 (N_28023,N_25737,N_25142);
nor U28024 (N_28024,N_25206,N_25185);
or U28025 (N_28025,N_24807,N_24961);
or U28026 (N_28026,N_26873,N_24710);
nor U28027 (N_28027,N_26586,N_24399);
and U28028 (N_28028,N_26308,N_25863);
nor U28029 (N_28029,N_24202,N_25208);
nand U28030 (N_28030,N_26788,N_25435);
and U28031 (N_28031,N_24234,N_24923);
or U28032 (N_28032,N_25639,N_26779);
or U28033 (N_28033,N_26776,N_24402);
xnor U28034 (N_28034,N_26039,N_25125);
xnor U28035 (N_28035,N_24415,N_24531);
nor U28036 (N_28036,N_24873,N_24538);
or U28037 (N_28037,N_26682,N_26016);
or U28038 (N_28038,N_25545,N_26769);
or U28039 (N_28039,N_24838,N_25580);
and U28040 (N_28040,N_25292,N_26938);
nand U28041 (N_28041,N_24282,N_25355);
and U28042 (N_28042,N_26611,N_26424);
xor U28043 (N_28043,N_26336,N_26328);
and U28044 (N_28044,N_25768,N_25710);
and U28045 (N_28045,N_26869,N_26204);
xor U28046 (N_28046,N_25218,N_26474);
and U28047 (N_28047,N_24917,N_25577);
xor U28048 (N_28048,N_26773,N_25478);
nand U28049 (N_28049,N_25119,N_26711);
nor U28050 (N_28050,N_25447,N_24983);
or U28051 (N_28051,N_25458,N_26226);
or U28052 (N_28052,N_25833,N_24722);
nand U28053 (N_28053,N_25440,N_26547);
nand U28054 (N_28054,N_24040,N_26196);
or U28055 (N_28055,N_25788,N_25369);
nand U28056 (N_28056,N_25202,N_25876);
nand U28057 (N_28057,N_26251,N_25176);
nand U28058 (N_28058,N_24295,N_26378);
nand U28059 (N_28059,N_25708,N_25412);
nor U28060 (N_28060,N_24156,N_25043);
and U28061 (N_28061,N_25989,N_24021);
or U28062 (N_28062,N_26737,N_25434);
or U28063 (N_28063,N_25571,N_24631);
or U28064 (N_28064,N_26370,N_24888);
nor U28065 (N_28065,N_24056,N_24154);
nand U28066 (N_28066,N_26724,N_24237);
or U28067 (N_28067,N_24477,N_26632);
and U28068 (N_28068,N_26886,N_26519);
nand U28069 (N_28069,N_24165,N_25797);
xnor U28070 (N_28070,N_25234,N_24408);
nor U28071 (N_28071,N_25352,N_26915);
nor U28072 (N_28072,N_25688,N_26576);
nand U28073 (N_28073,N_25662,N_25470);
or U28074 (N_28074,N_24793,N_24188);
xor U28075 (N_28075,N_25713,N_24369);
nand U28076 (N_28076,N_25922,N_26136);
and U28077 (N_28077,N_24361,N_26999);
nand U28078 (N_28078,N_25286,N_25793);
nor U28079 (N_28079,N_24395,N_24074);
or U28080 (N_28080,N_26117,N_24374);
or U28081 (N_28081,N_26871,N_24175);
nor U28082 (N_28082,N_24675,N_24633);
nor U28083 (N_28083,N_25480,N_25861);
xnor U28084 (N_28084,N_24980,N_25679);
nor U28085 (N_28085,N_24747,N_25262);
and U28086 (N_28086,N_24771,N_24032);
or U28087 (N_28087,N_26169,N_24726);
xnor U28088 (N_28088,N_26398,N_25048);
nand U28089 (N_28089,N_25211,N_25253);
or U28090 (N_28090,N_24324,N_24626);
and U28091 (N_28091,N_26190,N_24209);
nand U28092 (N_28092,N_24080,N_26529);
or U28093 (N_28093,N_26518,N_24957);
nor U28094 (N_28094,N_24255,N_26480);
or U28095 (N_28095,N_24869,N_24025);
nor U28096 (N_28096,N_25871,N_24562);
or U28097 (N_28097,N_25620,N_24717);
and U28098 (N_28098,N_24338,N_24363);
xnor U28099 (N_28099,N_26996,N_25516);
xor U28100 (N_28100,N_25601,N_25368);
or U28101 (N_28101,N_26469,N_26266);
and U28102 (N_28102,N_25123,N_26550);
xnor U28103 (N_28103,N_26052,N_25063);
nand U28104 (N_28104,N_24410,N_24657);
and U28105 (N_28105,N_25581,N_25865);
xnor U28106 (N_28106,N_24853,N_26500);
nor U28107 (N_28107,N_24715,N_25913);
or U28108 (N_28108,N_25693,N_24135);
or U28109 (N_28109,N_24519,N_25459);
xor U28110 (N_28110,N_24006,N_25004);
nand U28111 (N_28111,N_24008,N_24777);
and U28112 (N_28112,N_25075,N_26789);
nand U28113 (N_28113,N_26878,N_24364);
or U28114 (N_28114,N_24589,N_26756);
nor U28115 (N_28115,N_24093,N_24965);
and U28116 (N_28116,N_26629,N_25543);
nand U28117 (N_28117,N_24092,N_26738);
nand U28118 (N_28118,N_24051,N_24468);
or U28119 (N_28119,N_25322,N_25709);
nor U28120 (N_28120,N_26207,N_24241);
or U28121 (N_28121,N_26030,N_26653);
nand U28122 (N_28122,N_25126,N_25725);
and U28123 (N_28123,N_24326,N_26839);
and U28124 (N_28124,N_24062,N_25669);
nor U28125 (N_28125,N_25509,N_25552);
and U28126 (N_28126,N_26257,N_25290);
or U28127 (N_28127,N_24348,N_25307);
or U28128 (N_28128,N_24439,N_25983);
xor U28129 (N_28129,N_25343,N_25452);
xnor U28130 (N_28130,N_24102,N_25137);
xor U28131 (N_28131,N_24383,N_25492);
nor U28132 (N_28132,N_24740,N_26809);
or U28133 (N_28133,N_26837,N_25728);
xnor U28134 (N_28134,N_25430,N_26252);
xnor U28135 (N_28135,N_24696,N_24386);
and U28136 (N_28136,N_24803,N_24349);
or U28137 (N_28137,N_26782,N_25968);
xor U28138 (N_28138,N_24029,N_26104);
or U28139 (N_28139,N_26440,N_26906);
or U28140 (N_28140,N_25568,N_25870);
nor U28141 (N_28141,N_25145,N_26379);
xor U28142 (N_28142,N_24671,N_25158);
nor U28143 (N_28143,N_24208,N_24405);
and U28144 (N_28144,N_25117,N_25228);
or U28145 (N_28145,N_24599,N_24647);
nor U28146 (N_28146,N_26890,N_26817);
nor U28147 (N_28147,N_25378,N_26751);
or U28148 (N_28148,N_24692,N_26101);
and U28149 (N_28149,N_25128,N_26146);
or U28150 (N_28150,N_24664,N_24365);
xor U28151 (N_28151,N_24087,N_25014);
xor U28152 (N_28152,N_26783,N_25080);
xor U28153 (N_28153,N_25331,N_25700);
xnor U28154 (N_28154,N_26792,N_25248);
and U28155 (N_28155,N_24513,N_26674);
nand U28156 (N_28156,N_26800,N_26037);
and U28157 (N_28157,N_24617,N_24686);
and U28158 (N_28158,N_25409,N_26445);
and U28159 (N_28159,N_24480,N_24112);
or U28160 (N_28160,N_25016,N_26084);
nand U28161 (N_28161,N_24576,N_25313);
or U28162 (N_28162,N_25776,N_25514);
nor U28163 (N_28163,N_25747,N_24243);
nor U28164 (N_28164,N_24563,N_26289);
or U28165 (N_28165,N_25781,N_26043);
xor U28166 (N_28166,N_25766,N_24713);
nand U28167 (N_28167,N_26898,N_26444);
xnor U28168 (N_28168,N_25406,N_26883);
or U28169 (N_28169,N_24705,N_25244);
nand U28170 (N_28170,N_26152,N_26263);
nor U28171 (N_28171,N_26861,N_24039);
nor U28172 (N_28172,N_25317,N_26970);
nand U28173 (N_28173,N_26582,N_24311);
nor U28174 (N_28174,N_26689,N_24333);
or U28175 (N_28175,N_25668,N_25124);
nand U28176 (N_28176,N_25226,N_25427);
or U28177 (N_28177,N_25730,N_26129);
nor U28178 (N_28178,N_26509,N_25987);
xor U28179 (N_28179,N_26763,N_26686);
and U28180 (N_28180,N_26493,N_25657);
nand U28181 (N_28181,N_25525,N_25917);
or U28182 (N_28182,N_25998,N_26367);
nor U28183 (N_28183,N_25667,N_24024);
and U28184 (N_28184,N_25928,N_24723);
nand U28185 (N_28185,N_25802,N_26228);
or U28186 (N_28186,N_25959,N_24278);
or U28187 (N_28187,N_25611,N_26767);
nand U28188 (N_28188,N_25279,N_26046);
nand U28189 (N_28189,N_26614,N_25719);
nand U28190 (N_28190,N_26921,N_25518);
xor U28191 (N_28191,N_25399,N_26002);
or U28192 (N_28192,N_24920,N_24308);
nor U28193 (N_28193,N_26615,N_25816);
or U28194 (N_28194,N_24272,N_25832);
and U28195 (N_28195,N_26151,N_25114);
xnor U28196 (N_28196,N_26707,N_24072);
and U28197 (N_28197,N_26701,N_26320);
or U28198 (N_28198,N_26418,N_26725);
xnor U28199 (N_28199,N_26961,N_26276);
nand U28200 (N_28200,N_26448,N_26626);
or U28201 (N_28201,N_26286,N_26017);
nand U28202 (N_28202,N_26625,N_25758);
nor U28203 (N_28203,N_25426,N_26172);
or U28204 (N_28204,N_25030,N_24031);
xor U28205 (N_28205,N_25734,N_26924);
nor U28206 (N_28206,N_26236,N_26434);
xor U28207 (N_28207,N_24206,N_24162);
or U28208 (N_28208,N_24157,N_25274);
xor U28209 (N_28209,N_26137,N_24772);
nand U28210 (N_28210,N_26899,N_24526);
nor U28211 (N_28211,N_26020,N_26214);
or U28212 (N_28212,N_25767,N_25814);
nor U28213 (N_28213,N_25296,N_26808);
or U28214 (N_28214,N_25127,N_24540);
nand U28215 (N_28215,N_25946,N_25886);
nor U28216 (N_28216,N_25632,N_26874);
and U28217 (N_28217,N_24688,N_24422);
nor U28218 (N_28218,N_24192,N_24266);
xor U28219 (N_28219,N_24535,N_25519);
and U28220 (N_28220,N_24485,N_24046);
and U28221 (N_28221,N_24125,N_25268);
nor U28222 (N_28222,N_24482,N_26732);
nor U28223 (N_28223,N_26585,N_24158);
and U28224 (N_28224,N_26387,N_25727);
and U28225 (N_28225,N_25460,N_26470);
xor U28226 (N_28226,N_26197,N_26011);
or U28227 (N_28227,N_25605,N_25933);
nor U28228 (N_28228,N_24507,N_26318);
xor U28229 (N_28229,N_25284,N_26012);
nor U28230 (N_28230,N_25777,N_24094);
nor U28231 (N_28231,N_25420,N_26319);
and U28232 (N_28232,N_25531,N_25885);
or U28233 (N_28233,N_25471,N_24475);
xnor U28234 (N_28234,N_24289,N_24616);
or U28235 (N_28235,N_25320,N_25807);
and U28236 (N_28236,N_24592,N_25791);
nand U28237 (N_28237,N_25141,N_25271);
nor U28238 (N_28238,N_24607,N_24629);
or U28239 (N_28239,N_26778,N_26851);
nor U28240 (N_28240,N_25433,N_25808);
or U28241 (N_28241,N_25548,N_26411);
nor U28242 (N_28242,N_26933,N_24864);
xor U28243 (N_28243,N_26213,N_26790);
and U28244 (N_28244,N_26660,N_24187);
and U28245 (N_28245,N_25254,N_25541);
and U28246 (N_28246,N_25362,N_25993);
or U28247 (N_28247,N_25169,N_26868);
or U28248 (N_28248,N_26936,N_26948);
nand U28249 (N_28249,N_26192,N_25466);
or U28250 (N_28250,N_26998,N_24986);
nand U28251 (N_28251,N_25197,N_26902);
xnor U28252 (N_28252,N_26486,N_25905);
nor U28253 (N_28253,N_24457,N_24898);
or U28254 (N_28254,N_25068,N_26180);
or U28255 (N_28255,N_24982,N_26508);
xnor U28256 (N_28256,N_24525,N_25162);
xnor U28257 (N_28257,N_26224,N_26080);
or U28258 (N_28258,N_26731,N_24178);
xnor U28259 (N_28259,N_26091,N_24099);
or U28260 (N_28260,N_24669,N_24139);
and U28261 (N_28261,N_24706,N_26013);
xnor U28262 (N_28262,N_24727,N_24495);
xnor U28263 (N_28263,N_25099,N_24026);
nor U28264 (N_28264,N_25943,N_25977);
xor U28265 (N_28265,N_26481,N_25199);
nand U28266 (N_28266,N_24483,N_26884);
xnor U28267 (N_28267,N_24183,N_25428);
nor U28268 (N_28268,N_25841,N_26062);
nand U28269 (N_28269,N_25316,N_26235);
and U28270 (N_28270,N_24287,N_26563);
or U28271 (N_28271,N_24808,N_24069);
and U28272 (N_28272,N_25901,N_25690);
or U28273 (N_28273,N_24356,N_24928);
xor U28274 (N_28274,N_24411,N_24819);
nor U28275 (N_28275,N_26275,N_26282);
nor U28276 (N_28276,N_25565,N_26134);
nor U28277 (N_28277,N_26138,N_26388);
nand U28278 (N_28278,N_26375,N_26937);
nor U28279 (N_28279,N_25382,N_26297);
nand U28280 (N_28280,N_25836,N_24760);
and U28281 (N_28281,N_24461,N_26644);
xor U28282 (N_28282,N_24606,N_26488);
or U28283 (N_28283,N_26281,N_24442);
and U28284 (N_28284,N_26935,N_26270);
nor U28285 (N_28285,N_24336,N_26537);
and U28286 (N_28286,N_25914,N_24573);
or U28287 (N_28287,N_25769,N_26627);
or U28288 (N_28288,N_24325,N_25225);
or U28289 (N_28289,N_24331,N_24330);
xnor U28290 (N_28290,N_25454,N_24170);
and U28291 (N_28291,N_24528,N_24115);
nand U28292 (N_28292,N_25489,N_25858);
xor U28293 (N_28293,N_26287,N_26912);
or U28294 (N_28294,N_24855,N_25761);
nand U28295 (N_28295,N_26261,N_25938);
nand U28296 (N_28296,N_25333,N_24645);
and U28297 (N_28297,N_26021,N_26218);
or U28298 (N_28298,N_25779,N_24775);
nor U28299 (N_28299,N_24575,N_26958);
and U28300 (N_28300,N_24701,N_25806);
nor U28301 (N_28301,N_24585,N_24764);
nor U28302 (N_28302,N_26951,N_25681);
and U28303 (N_28303,N_25410,N_25964);
xor U28304 (N_28304,N_26363,N_26253);
xnor U28305 (N_28305,N_25191,N_26605);
and U28306 (N_28306,N_26106,N_24684);
and U28307 (N_28307,N_24549,N_25442);
nand U28308 (N_28308,N_25995,N_24847);
and U28309 (N_28309,N_26126,N_24828);
or U28310 (N_28310,N_26840,N_24708);
and U28311 (N_28311,N_25754,N_25724);
xnor U28312 (N_28312,N_26450,N_25345);
or U28313 (N_28313,N_24841,N_25511);
and U28314 (N_28314,N_25614,N_26306);
xor U28315 (N_28315,N_24003,N_25537);
and U28316 (N_28316,N_26971,N_25235);
nor U28317 (N_28317,N_24901,N_26997);
and U28318 (N_28318,N_24057,N_24877);
xor U28319 (N_28319,N_24635,N_26455);
or U28320 (N_28320,N_26066,N_24500);
xor U28321 (N_28321,N_25210,N_24357);
nor U28322 (N_28322,N_26852,N_26309);
and U28323 (N_28323,N_24273,N_24132);
nor U28324 (N_28324,N_25784,N_25985);
xor U28325 (N_28325,N_26680,N_26339);
xnor U28326 (N_28326,N_25094,N_26744);
xnor U28327 (N_28327,N_26173,N_25303);
nand U28328 (N_28328,N_25073,N_25517);
and U28329 (N_28329,N_25182,N_25178);
nor U28330 (N_28330,N_25256,N_25907);
nor U28331 (N_28331,N_24130,N_26813);
xor U28332 (N_28332,N_25240,N_25484);
nor U28333 (N_28333,N_25627,N_25260);
nand U28334 (N_28334,N_24435,N_25386);
nand U28335 (N_28335,N_26354,N_25144);
nand U28336 (N_28336,N_24050,N_26581);
nor U28337 (N_28337,N_24070,N_24832);
and U28338 (N_28338,N_25990,N_25404);
nor U28339 (N_28339,N_25163,N_24921);
xor U28340 (N_28340,N_25242,N_26457);
nand U28341 (N_28341,N_24846,N_26552);
or U28342 (N_28342,N_26880,N_25980);
and U28343 (N_28343,N_25618,N_26786);
nor U28344 (N_28344,N_25637,N_25718);
nor U28345 (N_28345,N_26963,N_24142);
nor U28346 (N_28346,N_26079,N_26977);
and U28347 (N_28347,N_25789,N_26796);
nor U28348 (N_28348,N_25177,N_25521);
xor U28349 (N_28349,N_26815,N_26166);
nor U28350 (N_28350,N_24258,N_26713);
or U28351 (N_28351,N_25960,N_24988);
or U28352 (N_28352,N_26816,N_25101);
nor U28353 (N_28353,N_26018,N_25036);
or U28354 (N_28354,N_24946,N_24867);
nor U28355 (N_28355,N_24757,N_25918);
and U28356 (N_28356,N_24174,N_24210);
xor U28357 (N_28357,N_26243,N_24220);
nand U28358 (N_28358,N_25354,N_25931);
nand U28359 (N_28359,N_26820,N_26426);
nor U28360 (N_28360,N_26847,N_24733);
nand U28361 (N_28361,N_25155,N_26944);
nor U28362 (N_28362,N_24235,N_26376);
and U28363 (N_28363,N_24281,N_26775);
and U28364 (N_28364,N_26132,N_26564);
and U28365 (N_28365,N_24022,N_25081);
and U28366 (N_28366,N_25992,N_25561);
or U28367 (N_28367,N_25066,N_26410);
and U28368 (N_28368,N_25896,N_25854);
and U28369 (N_28369,N_26876,N_26098);
nor U28370 (N_28370,N_25684,N_26830);
nand U28371 (N_28371,N_24140,N_25683);
nor U28372 (N_28372,N_25610,N_24450);
and U28373 (N_28373,N_26036,N_25869);
nand U28374 (N_28374,N_24973,N_24231);
nor U28375 (N_28375,N_24018,N_25009);
xor U28376 (N_28376,N_25994,N_26503);
or U28377 (N_28377,N_26575,N_24499);
and U28378 (N_28378,N_25785,N_26728);
nor U28379 (N_28379,N_26165,N_24120);
nand U28380 (N_28380,N_26346,N_25550);
nor U28381 (N_28381,N_26003,N_26864);
xor U28382 (N_28382,N_24262,N_26863);
and U28383 (N_28383,N_24238,N_25034);
xnor U28384 (N_28384,N_25473,N_24341);
or U28385 (N_28385,N_25846,N_25991);
or U28386 (N_28386,N_25488,N_25783);
xnor U28387 (N_28387,N_25495,N_25170);
nand U28388 (N_28388,N_24000,N_24787);
nor U28389 (N_28389,N_25551,N_24090);
and U28390 (N_28390,N_26007,N_24095);
nor U28391 (N_28391,N_24128,N_26768);
nand U28392 (N_28392,N_25926,N_24199);
nand U28393 (N_28393,N_24045,N_26616);
nor U28394 (N_28394,N_25636,N_26430);
xnor U28395 (N_28395,N_26979,N_24293);
or U28396 (N_28396,N_25563,N_25223);
nor U28397 (N_28397,N_25312,N_24978);
nor U28398 (N_28398,N_25900,N_26801);
or U28399 (N_28399,N_24259,N_25453);
and U28400 (N_28400,N_26990,N_24226);
xor U28401 (N_28401,N_25535,N_25341);
nand U28402 (N_28402,N_25039,N_26102);
and U28403 (N_28403,N_26465,N_26742);
xnor U28404 (N_28404,N_26917,N_26972);
nor U28405 (N_28405,N_26034,N_25339);
nor U28406 (N_28406,N_24663,N_24815);
or U28407 (N_28407,N_25000,N_24463);
and U28408 (N_28408,N_25076,N_25376);
xor U28409 (N_28409,N_26676,N_24546);
or U28410 (N_28410,N_24559,N_26642);
or U28411 (N_28411,N_25986,N_26521);
xor U28412 (N_28412,N_24211,N_24571);
nand U28413 (N_28413,N_26849,N_26404);
nand U28414 (N_28414,N_24075,N_25764);
and U28415 (N_28415,N_24745,N_24131);
nand U28416 (N_28416,N_26193,N_26484);
xnor U28417 (N_28417,N_24375,N_26941);
nor U28418 (N_28418,N_25751,N_25138);
xor U28419 (N_28419,N_26882,N_24416);
and U28420 (N_28420,N_24608,N_25384);
xnor U28421 (N_28421,N_25423,N_26993);
and U28422 (N_28422,N_26926,N_24756);
xor U28423 (N_28423,N_26049,N_26461);
nor U28424 (N_28424,N_25102,N_26718);
nor U28425 (N_28425,N_25375,N_26377);
or U28426 (N_28426,N_25157,N_24655);
nor U28427 (N_28427,N_26407,N_25023);
nor U28428 (N_28428,N_26123,N_26122);
xor U28429 (N_28429,N_24091,N_24770);
nor U28430 (N_28430,N_25028,N_24249);
xor U28431 (N_28431,N_24196,N_25932);
and U28432 (N_28432,N_24060,N_25020);
nand U28433 (N_28433,N_25903,N_24084);
and U28434 (N_28434,N_25756,N_24985);
and U28435 (N_28435,N_25366,N_26312);
xnor U28436 (N_28436,N_25400,N_24248);
nor U28437 (N_28437,N_26361,N_26330);
and U28438 (N_28438,N_25835,N_26588);
nand U28439 (N_28439,N_24851,N_26121);
or U28440 (N_28440,N_24992,N_25817);
nor U28441 (N_28441,N_26223,N_25302);
and U28442 (N_28442,N_24537,N_26772);
xnor U28443 (N_28443,N_24459,N_26975);
or U28444 (N_28444,N_25095,N_25300);
and U28445 (N_28445,N_26157,N_25975);
and U28446 (N_28446,N_24970,N_25778);
nand U28447 (N_28447,N_26061,N_25644);
nor U28448 (N_28448,N_25017,N_26441);
nor U28449 (N_28449,N_25799,N_26209);
nand U28450 (N_28450,N_25160,N_25691);
and U28451 (N_28451,N_24883,N_26385);
xor U28452 (N_28452,N_25445,N_25391);
xnor U28453 (N_28453,N_26928,N_24164);
nand U28454 (N_28454,N_24667,N_25438);
xnor U28455 (N_28455,N_24762,N_25877);
or U28456 (N_28456,N_26222,N_26203);
or U28457 (N_28457,N_24993,N_24221);
nor U28458 (N_28458,N_24814,N_25019);
and U28459 (N_28459,N_25874,N_25512);
or U28460 (N_28460,N_24181,N_24890);
xnor U28461 (N_28461,N_26909,N_24017);
or U28462 (N_28462,N_25122,N_25500);
nand U28463 (N_28463,N_24899,N_25140);
or U28464 (N_28464,N_26741,N_24802);
nand U28465 (N_28465,N_26657,N_25617);
xnor U28466 (N_28466,N_26974,N_25013);
or U28467 (N_28467,N_24085,N_25505);
nand U28468 (N_28468,N_24167,N_25067);
nor U28469 (N_28469,N_24047,N_24801);
nand U28470 (N_28470,N_26458,N_26200);
and U28471 (N_28471,N_24997,N_25221);
xnor U28472 (N_28472,N_24577,N_25046);
nor U28473 (N_28473,N_24002,N_24239);
and U28474 (N_28474,N_26175,N_24044);
xnor U28475 (N_28475,N_26877,N_25626);
or U28476 (N_28476,N_25967,N_24345);
xnor U28477 (N_28477,N_26443,N_24903);
nor U28478 (N_28478,N_25884,N_24149);
nand U28479 (N_28479,N_25750,N_24944);
and U28480 (N_28480,N_25304,N_25912);
and U28481 (N_28481,N_26023,N_26766);
and U28482 (N_28482,N_24765,N_26885);
xnor U28483 (N_28483,N_26024,N_25329);
or U28484 (N_28484,N_26901,N_25429);
xnor U28485 (N_28485,N_25083,N_25640);
nand U28486 (N_28486,N_25022,N_25431);
xor U28487 (N_28487,N_26490,N_24138);
nand U28488 (N_28488,N_25383,N_25759);
xnor U28489 (N_28489,N_26188,N_25853);
nand U28490 (N_28490,N_25851,N_24707);
nand U28491 (N_28491,N_25132,N_24652);
and U28492 (N_28492,N_26396,N_25949);
and U28493 (N_28493,N_24893,N_26390);
nand U28494 (N_28494,N_26753,N_25062);
nand U28495 (N_28495,N_24011,N_24907);
xnor U28496 (N_28496,N_26216,N_25721);
and U28497 (N_28497,N_24454,N_24377);
nand U28498 (N_28498,N_25703,N_24534);
nor U28499 (N_28499,N_24905,N_24218);
nand U28500 (N_28500,N_25939,N_26879);
nand U28501 (N_28501,N_24430,N_25913);
nand U28502 (N_28502,N_24325,N_26913);
nor U28503 (N_28503,N_24964,N_25730);
nor U28504 (N_28504,N_25259,N_26291);
or U28505 (N_28505,N_25701,N_25553);
and U28506 (N_28506,N_24037,N_26258);
nor U28507 (N_28507,N_25955,N_26049);
nand U28508 (N_28508,N_24862,N_24677);
nand U28509 (N_28509,N_25493,N_26233);
nand U28510 (N_28510,N_26619,N_25636);
xnor U28511 (N_28511,N_26780,N_25702);
nand U28512 (N_28512,N_25654,N_24922);
nand U28513 (N_28513,N_25157,N_24332);
nor U28514 (N_28514,N_24286,N_24225);
nand U28515 (N_28515,N_24548,N_26308);
nand U28516 (N_28516,N_25019,N_24263);
xor U28517 (N_28517,N_25646,N_25196);
or U28518 (N_28518,N_25325,N_26586);
nor U28519 (N_28519,N_24247,N_24604);
xnor U28520 (N_28520,N_25467,N_25302);
and U28521 (N_28521,N_24013,N_24207);
or U28522 (N_28522,N_25031,N_25923);
xor U28523 (N_28523,N_26283,N_25816);
nor U28524 (N_28524,N_26138,N_25780);
or U28525 (N_28525,N_24595,N_24353);
nand U28526 (N_28526,N_26075,N_24187);
or U28527 (N_28527,N_24415,N_25714);
or U28528 (N_28528,N_25198,N_24515);
nor U28529 (N_28529,N_25703,N_26186);
nand U28530 (N_28530,N_25865,N_24090);
nor U28531 (N_28531,N_25499,N_26685);
nor U28532 (N_28532,N_24072,N_25089);
and U28533 (N_28533,N_25789,N_26041);
or U28534 (N_28534,N_26733,N_24588);
nand U28535 (N_28535,N_26727,N_24509);
and U28536 (N_28536,N_26389,N_25508);
and U28537 (N_28537,N_26981,N_24709);
and U28538 (N_28538,N_26825,N_24084);
nor U28539 (N_28539,N_24849,N_25646);
nor U28540 (N_28540,N_26922,N_25008);
nand U28541 (N_28541,N_24541,N_24246);
nand U28542 (N_28542,N_26709,N_25252);
and U28543 (N_28543,N_25650,N_24928);
or U28544 (N_28544,N_26981,N_25913);
nand U28545 (N_28545,N_24151,N_26819);
nor U28546 (N_28546,N_26422,N_24509);
nor U28547 (N_28547,N_24247,N_24093);
and U28548 (N_28548,N_26875,N_24713);
nand U28549 (N_28549,N_26955,N_25188);
and U28550 (N_28550,N_25253,N_26111);
or U28551 (N_28551,N_26894,N_26060);
nand U28552 (N_28552,N_26131,N_26444);
nor U28553 (N_28553,N_24363,N_26770);
or U28554 (N_28554,N_24951,N_24733);
xor U28555 (N_28555,N_25456,N_26633);
nand U28556 (N_28556,N_26606,N_24528);
and U28557 (N_28557,N_24094,N_24754);
or U28558 (N_28558,N_25046,N_26989);
nand U28559 (N_28559,N_24117,N_25221);
or U28560 (N_28560,N_24825,N_26195);
or U28561 (N_28561,N_25782,N_24903);
or U28562 (N_28562,N_26638,N_26078);
or U28563 (N_28563,N_26789,N_26006);
nor U28564 (N_28564,N_25579,N_24388);
or U28565 (N_28565,N_26525,N_25758);
and U28566 (N_28566,N_26221,N_24883);
xor U28567 (N_28567,N_26292,N_24272);
nand U28568 (N_28568,N_25366,N_24621);
nor U28569 (N_28569,N_25410,N_25374);
and U28570 (N_28570,N_26549,N_25446);
xor U28571 (N_28571,N_24706,N_26384);
and U28572 (N_28572,N_24411,N_24548);
and U28573 (N_28573,N_24297,N_24396);
nor U28574 (N_28574,N_26672,N_25891);
nor U28575 (N_28575,N_26238,N_24337);
xnor U28576 (N_28576,N_24158,N_25099);
or U28577 (N_28577,N_26641,N_24807);
nor U28578 (N_28578,N_26590,N_26273);
nor U28579 (N_28579,N_25929,N_24889);
and U28580 (N_28580,N_25555,N_24984);
or U28581 (N_28581,N_26572,N_24588);
xnor U28582 (N_28582,N_26135,N_26782);
nor U28583 (N_28583,N_25691,N_24580);
or U28584 (N_28584,N_26864,N_25872);
nor U28585 (N_28585,N_26542,N_26647);
xnor U28586 (N_28586,N_26116,N_25227);
or U28587 (N_28587,N_24450,N_26645);
nor U28588 (N_28588,N_26931,N_26382);
and U28589 (N_28589,N_24842,N_25220);
nand U28590 (N_28590,N_25050,N_26971);
nor U28591 (N_28591,N_24000,N_26025);
xnor U28592 (N_28592,N_26312,N_24559);
nand U28593 (N_28593,N_25979,N_24421);
and U28594 (N_28594,N_24374,N_26392);
xnor U28595 (N_28595,N_26093,N_25175);
xor U28596 (N_28596,N_25763,N_26325);
nand U28597 (N_28597,N_25488,N_24821);
nand U28598 (N_28598,N_25469,N_25459);
and U28599 (N_28599,N_26321,N_24538);
and U28600 (N_28600,N_25137,N_24549);
or U28601 (N_28601,N_24629,N_26927);
nand U28602 (N_28602,N_25683,N_25006);
or U28603 (N_28603,N_26190,N_25150);
and U28604 (N_28604,N_26633,N_24308);
or U28605 (N_28605,N_25644,N_26616);
xor U28606 (N_28606,N_26667,N_26579);
or U28607 (N_28607,N_25941,N_26927);
nand U28608 (N_28608,N_24157,N_24790);
and U28609 (N_28609,N_26144,N_26497);
nor U28610 (N_28610,N_26924,N_26114);
nand U28611 (N_28611,N_26029,N_26395);
nand U28612 (N_28612,N_26804,N_26695);
nand U28613 (N_28613,N_26556,N_24767);
xnor U28614 (N_28614,N_26553,N_24484);
nor U28615 (N_28615,N_26848,N_24170);
and U28616 (N_28616,N_25737,N_25566);
xnor U28617 (N_28617,N_25719,N_24158);
nand U28618 (N_28618,N_26413,N_25476);
nor U28619 (N_28619,N_24560,N_26114);
or U28620 (N_28620,N_24375,N_24035);
xnor U28621 (N_28621,N_26316,N_25183);
and U28622 (N_28622,N_24632,N_24308);
or U28623 (N_28623,N_25639,N_26749);
nor U28624 (N_28624,N_25874,N_24754);
and U28625 (N_28625,N_24064,N_26817);
nand U28626 (N_28626,N_25481,N_24319);
or U28627 (N_28627,N_25732,N_25453);
or U28628 (N_28628,N_25255,N_24156);
or U28629 (N_28629,N_25956,N_25756);
nor U28630 (N_28630,N_26449,N_26615);
and U28631 (N_28631,N_26583,N_26998);
and U28632 (N_28632,N_26893,N_24273);
xor U28633 (N_28633,N_24737,N_26930);
nand U28634 (N_28634,N_24714,N_26927);
or U28635 (N_28635,N_25234,N_24018);
xnor U28636 (N_28636,N_24608,N_25561);
nand U28637 (N_28637,N_26521,N_25331);
xor U28638 (N_28638,N_24300,N_24496);
nand U28639 (N_28639,N_26766,N_24665);
or U28640 (N_28640,N_25048,N_24539);
xnor U28641 (N_28641,N_25960,N_25131);
nor U28642 (N_28642,N_25318,N_26022);
nor U28643 (N_28643,N_24321,N_26914);
nor U28644 (N_28644,N_26931,N_24033);
xor U28645 (N_28645,N_26867,N_25028);
or U28646 (N_28646,N_25319,N_24861);
and U28647 (N_28647,N_26145,N_25285);
xnor U28648 (N_28648,N_24254,N_24414);
xnor U28649 (N_28649,N_25080,N_26417);
and U28650 (N_28650,N_24783,N_26858);
and U28651 (N_28651,N_24961,N_26867);
or U28652 (N_28652,N_26864,N_25518);
or U28653 (N_28653,N_24261,N_24427);
or U28654 (N_28654,N_25339,N_26087);
nor U28655 (N_28655,N_25517,N_26317);
nand U28656 (N_28656,N_26209,N_24608);
nor U28657 (N_28657,N_26853,N_26646);
nor U28658 (N_28658,N_25854,N_25984);
and U28659 (N_28659,N_26547,N_26980);
and U28660 (N_28660,N_25737,N_24208);
xnor U28661 (N_28661,N_26413,N_26299);
or U28662 (N_28662,N_25200,N_25496);
nor U28663 (N_28663,N_25172,N_26583);
or U28664 (N_28664,N_26620,N_24567);
xnor U28665 (N_28665,N_26976,N_25017);
and U28666 (N_28666,N_26089,N_25426);
or U28667 (N_28667,N_26315,N_24630);
xnor U28668 (N_28668,N_26089,N_26120);
nand U28669 (N_28669,N_26476,N_26903);
nor U28670 (N_28670,N_25858,N_25872);
nand U28671 (N_28671,N_26362,N_24999);
nor U28672 (N_28672,N_24189,N_25839);
nor U28673 (N_28673,N_24611,N_26636);
and U28674 (N_28674,N_25308,N_25783);
and U28675 (N_28675,N_26492,N_24355);
xor U28676 (N_28676,N_26777,N_25263);
xnor U28677 (N_28677,N_24563,N_26399);
and U28678 (N_28678,N_26725,N_26621);
and U28679 (N_28679,N_25314,N_25687);
nand U28680 (N_28680,N_24819,N_25286);
and U28681 (N_28681,N_26198,N_24402);
or U28682 (N_28682,N_26927,N_25992);
nand U28683 (N_28683,N_26762,N_25855);
nor U28684 (N_28684,N_24560,N_25802);
nor U28685 (N_28685,N_26548,N_24765);
or U28686 (N_28686,N_25396,N_25809);
or U28687 (N_28687,N_26377,N_26794);
xnor U28688 (N_28688,N_24900,N_24214);
and U28689 (N_28689,N_26310,N_25353);
and U28690 (N_28690,N_25018,N_25590);
and U28691 (N_28691,N_24616,N_24822);
nor U28692 (N_28692,N_26215,N_24305);
or U28693 (N_28693,N_24498,N_26735);
or U28694 (N_28694,N_24858,N_25253);
xor U28695 (N_28695,N_25204,N_26021);
nand U28696 (N_28696,N_25045,N_24505);
and U28697 (N_28697,N_26217,N_26570);
and U28698 (N_28698,N_24001,N_24003);
or U28699 (N_28699,N_24847,N_25572);
or U28700 (N_28700,N_25905,N_25735);
xnor U28701 (N_28701,N_26889,N_24598);
or U28702 (N_28702,N_26146,N_26137);
or U28703 (N_28703,N_24224,N_25463);
xor U28704 (N_28704,N_24487,N_26038);
nand U28705 (N_28705,N_26417,N_24057);
xor U28706 (N_28706,N_26646,N_26520);
nor U28707 (N_28707,N_26750,N_26646);
or U28708 (N_28708,N_26072,N_25528);
nor U28709 (N_28709,N_24107,N_25021);
nand U28710 (N_28710,N_24929,N_25765);
or U28711 (N_28711,N_26489,N_25041);
or U28712 (N_28712,N_26187,N_26387);
or U28713 (N_28713,N_26944,N_25753);
xor U28714 (N_28714,N_24351,N_24874);
xnor U28715 (N_28715,N_24008,N_26014);
and U28716 (N_28716,N_26340,N_26747);
nor U28717 (N_28717,N_24512,N_24477);
xor U28718 (N_28718,N_24595,N_24872);
and U28719 (N_28719,N_26156,N_24545);
and U28720 (N_28720,N_26179,N_26689);
or U28721 (N_28721,N_24964,N_26337);
or U28722 (N_28722,N_25407,N_26902);
nand U28723 (N_28723,N_25057,N_24932);
nand U28724 (N_28724,N_26005,N_25451);
nor U28725 (N_28725,N_26148,N_24520);
nand U28726 (N_28726,N_26893,N_24845);
xnor U28727 (N_28727,N_24437,N_26059);
or U28728 (N_28728,N_24842,N_24609);
nand U28729 (N_28729,N_24746,N_25099);
nor U28730 (N_28730,N_26413,N_24247);
xnor U28731 (N_28731,N_25353,N_25346);
nand U28732 (N_28732,N_24923,N_26989);
nand U28733 (N_28733,N_26732,N_25373);
and U28734 (N_28734,N_25191,N_26646);
and U28735 (N_28735,N_26056,N_26570);
nand U28736 (N_28736,N_25006,N_26075);
and U28737 (N_28737,N_25375,N_24682);
or U28738 (N_28738,N_25738,N_26259);
nand U28739 (N_28739,N_26305,N_25127);
nand U28740 (N_28740,N_25172,N_24430);
nand U28741 (N_28741,N_26101,N_24770);
nor U28742 (N_28742,N_25606,N_25235);
and U28743 (N_28743,N_25410,N_24030);
or U28744 (N_28744,N_26810,N_25651);
xor U28745 (N_28745,N_24764,N_26799);
nand U28746 (N_28746,N_25114,N_25917);
and U28747 (N_28747,N_26126,N_25300);
nand U28748 (N_28748,N_26850,N_25772);
xnor U28749 (N_28749,N_26030,N_26312);
nand U28750 (N_28750,N_24337,N_24918);
and U28751 (N_28751,N_26351,N_26964);
and U28752 (N_28752,N_25903,N_26295);
and U28753 (N_28753,N_25690,N_25502);
nor U28754 (N_28754,N_26264,N_26256);
nor U28755 (N_28755,N_25619,N_24793);
and U28756 (N_28756,N_25658,N_25742);
nor U28757 (N_28757,N_25480,N_24273);
xor U28758 (N_28758,N_25487,N_25282);
and U28759 (N_28759,N_25906,N_26180);
nand U28760 (N_28760,N_26977,N_24637);
nor U28761 (N_28761,N_24307,N_26010);
nor U28762 (N_28762,N_26341,N_24342);
nor U28763 (N_28763,N_26018,N_24862);
and U28764 (N_28764,N_25475,N_25904);
xnor U28765 (N_28765,N_24859,N_24197);
xnor U28766 (N_28766,N_25843,N_26384);
xor U28767 (N_28767,N_24109,N_25293);
and U28768 (N_28768,N_25533,N_25519);
and U28769 (N_28769,N_25538,N_24308);
nor U28770 (N_28770,N_26906,N_24579);
and U28771 (N_28771,N_24704,N_25801);
or U28772 (N_28772,N_26472,N_24116);
xor U28773 (N_28773,N_24225,N_25816);
nor U28774 (N_28774,N_24500,N_24166);
nor U28775 (N_28775,N_25879,N_24665);
xor U28776 (N_28776,N_26646,N_24543);
xnor U28777 (N_28777,N_26929,N_25667);
nor U28778 (N_28778,N_26492,N_24735);
nand U28779 (N_28779,N_26759,N_25412);
nand U28780 (N_28780,N_24754,N_24299);
nor U28781 (N_28781,N_25521,N_24879);
nand U28782 (N_28782,N_25679,N_24211);
and U28783 (N_28783,N_26105,N_24748);
and U28784 (N_28784,N_25379,N_25150);
and U28785 (N_28785,N_24542,N_24620);
and U28786 (N_28786,N_26073,N_26017);
and U28787 (N_28787,N_25896,N_24489);
nand U28788 (N_28788,N_26465,N_25258);
xnor U28789 (N_28789,N_26006,N_24868);
xor U28790 (N_28790,N_25061,N_24214);
or U28791 (N_28791,N_25006,N_25626);
xnor U28792 (N_28792,N_25381,N_24884);
nor U28793 (N_28793,N_24206,N_26286);
or U28794 (N_28794,N_26580,N_25491);
nand U28795 (N_28795,N_26226,N_25539);
or U28796 (N_28796,N_25354,N_25457);
xor U28797 (N_28797,N_25106,N_26113);
nand U28798 (N_28798,N_26222,N_25862);
nand U28799 (N_28799,N_24900,N_24503);
and U28800 (N_28800,N_24118,N_26211);
or U28801 (N_28801,N_25422,N_24298);
nor U28802 (N_28802,N_24331,N_26436);
and U28803 (N_28803,N_26890,N_24890);
nor U28804 (N_28804,N_24856,N_24343);
nand U28805 (N_28805,N_26736,N_25456);
or U28806 (N_28806,N_25333,N_25049);
and U28807 (N_28807,N_26104,N_24843);
and U28808 (N_28808,N_25177,N_24271);
xor U28809 (N_28809,N_24700,N_24656);
and U28810 (N_28810,N_25481,N_25735);
xor U28811 (N_28811,N_24763,N_25914);
xnor U28812 (N_28812,N_25799,N_25007);
nor U28813 (N_28813,N_24858,N_25280);
nor U28814 (N_28814,N_26072,N_25487);
and U28815 (N_28815,N_26555,N_26492);
xor U28816 (N_28816,N_26386,N_25021);
nand U28817 (N_28817,N_26882,N_25734);
and U28818 (N_28818,N_25586,N_24282);
nor U28819 (N_28819,N_26996,N_24424);
and U28820 (N_28820,N_24106,N_24688);
nor U28821 (N_28821,N_25994,N_25005);
and U28822 (N_28822,N_26164,N_24198);
or U28823 (N_28823,N_25572,N_26316);
nand U28824 (N_28824,N_24197,N_25022);
nor U28825 (N_28825,N_24748,N_24267);
xnor U28826 (N_28826,N_26453,N_26125);
nand U28827 (N_28827,N_24741,N_25850);
nand U28828 (N_28828,N_24371,N_26055);
xnor U28829 (N_28829,N_24663,N_26501);
or U28830 (N_28830,N_25090,N_25944);
xor U28831 (N_28831,N_25262,N_25299);
and U28832 (N_28832,N_25978,N_26210);
and U28833 (N_28833,N_25470,N_26484);
or U28834 (N_28834,N_25988,N_25842);
nor U28835 (N_28835,N_24228,N_25279);
nor U28836 (N_28836,N_24670,N_25080);
nand U28837 (N_28837,N_24854,N_24906);
xor U28838 (N_28838,N_25026,N_25010);
nand U28839 (N_28839,N_24267,N_25133);
or U28840 (N_28840,N_24782,N_24054);
xor U28841 (N_28841,N_26801,N_25661);
nor U28842 (N_28842,N_25106,N_25777);
xor U28843 (N_28843,N_24393,N_25195);
nor U28844 (N_28844,N_25475,N_26285);
nand U28845 (N_28845,N_26515,N_25870);
and U28846 (N_28846,N_26936,N_26753);
and U28847 (N_28847,N_25463,N_26222);
or U28848 (N_28848,N_25038,N_25153);
nand U28849 (N_28849,N_25734,N_26382);
and U28850 (N_28850,N_25295,N_24552);
nor U28851 (N_28851,N_26885,N_25579);
nor U28852 (N_28852,N_24425,N_24320);
xnor U28853 (N_28853,N_25372,N_25216);
xor U28854 (N_28854,N_24502,N_24850);
and U28855 (N_28855,N_26418,N_25207);
and U28856 (N_28856,N_24679,N_26677);
nand U28857 (N_28857,N_26601,N_25490);
xnor U28858 (N_28858,N_26144,N_26644);
or U28859 (N_28859,N_25260,N_24421);
and U28860 (N_28860,N_25006,N_24381);
nand U28861 (N_28861,N_26479,N_26918);
and U28862 (N_28862,N_24012,N_24624);
or U28863 (N_28863,N_26316,N_25516);
nor U28864 (N_28864,N_26170,N_26311);
nand U28865 (N_28865,N_24377,N_26143);
xor U28866 (N_28866,N_26539,N_26796);
or U28867 (N_28867,N_26974,N_25769);
xnor U28868 (N_28868,N_26453,N_25729);
xnor U28869 (N_28869,N_24239,N_24707);
nor U28870 (N_28870,N_24040,N_25403);
xor U28871 (N_28871,N_26645,N_26261);
nand U28872 (N_28872,N_25489,N_25790);
nor U28873 (N_28873,N_26523,N_26110);
or U28874 (N_28874,N_24219,N_26234);
or U28875 (N_28875,N_25787,N_26524);
xnor U28876 (N_28876,N_25850,N_26969);
and U28877 (N_28877,N_24798,N_26882);
or U28878 (N_28878,N_25881,N_25158);
xor U28879 (N_28879,N_26159,N_25835);
nor U28880 (N_28880,N_25383,N_24159);
or U28881 (N_28881,N_26942,N_24918);
and U28882 (N_28882,N_24124,N_25202);
and U28883 (N_28883,N_25601,N_25102);
and U28884 (N_28884,N_26268,N_24268);
nand U28885 (N_28885,N_26981,N_26835);
or U28886 (N_28886,N_25461,N_24461);
or U28887 (N_28887,N_25937,N_26595);
xnor U28888 (N_28888,N_25002,N_24747);
or U28889 (N_28889,N_26014,N_24762);
nand U28890 (N_28890,N_26193,N_24728);
xnor U28891 (N_28891,N_26410,N_26994);
xnor U28892 (N_28892,N_26333,N_24113);
xnor U28893 (N_28893,N_25037,N_26298);
xnor U28894 (N_28894,N_25163,N_24498);
xor U28895 (N_28895,N_25999,N_24631);
or U28896 (N_28896,N_26317,N_25627);
xnor U28897 (N_28897,N_26281,N_25658);
nor U28898 (N_28898,N_25003,N_24084);
xnor U28899 (N_28899,N_25550,N_24376);
nand U28900 (N_28900,N_24803,N_26054);
xnor U28901 (N_28901,N_24729,N_25642);
xnor U28902 (N_28902,N_26329,N_26424);
xnor U28903 (N_28903,N_24184,N_24643);
nor U28904 (N_28904,N_24286,N_25983);
nor U28905 (N_28905,N_24245,N_25103);
and U28906 (N_28906,N_25382,N_24330);
nor U28907 (N_28907,N_25630,N_25611);
or U28908 (N_28908,N_26255,N_25641);
nor U28909 (N_28909,N_25455,N_25619);
nor U28910 (N_28910,N_26040,N_24465);
or U28911 (N_28911,N_26529,N_25343);
xor U28912 (N_28912,N_26776,N_25937);
and U28913 (N_28913,N_25182,N_26735);
or U28914 (N_28914,N_26200,N_24614);
or U28915 (N_28915,N_24898,N_26287);
or U28916 (N_28916,N_26243,N_25662);
nand U28917 (N_28917,N_26208,N_25284);
nand U28918 (N_28918,N_25206,N_24132);
or U28919 (N_28919,N_26094,N_24265);
or U28920 (N_28920,N_26915,N_26919);
nand U28921 (N_28921,N_24916,N_25314);
xnor U28922 (N_28922,N_24267,N_24883);
nand U28923 (N_28923,N_26469,N_26984);
and U28924 (N_28924,N_25707,N_24302);
nor U28925 (N_28925,N_26237,N_25279);
and U28926 (N_28926,N_25312,N_25776);
and U28927 (N_28927,N_26213,N_24369);
nand U28928 (N_28928,N_25589,N_25508);
or U28929 (N_28929,N_24249,N_26568);
or U28930 (N_28930,N_25375,N_24799);
nor U28931 (N_28931,N_24664,N_24527);
and U28932 (N_28932,N_26164,N_24540);
or U28933 (N_28933,N_24218,N_25762);
nor U28934 (N_28934,N_24519,N_26533);
and U28935 (N_28935,N_24791,N_24696);
and U28936 (N_28936,N_25426,N_24830);
xor U28937 (N_28937,N_25688,N_24721);
and U28938 (N_28938,N_25353,N_26618);
or U28939 (N_28939,N_24983,N_24389);
nand U28940 (N_28940,N_24227,N_25923);
and U28941 (N_28941,N_25664,N_26533);
or U28942 (N_28942,N_24886,N_26795);
nand U28943 (N_28943,N_24189,N_24904);
nor U28944 (N_28944,N_26697,N_24106);
nor U28945 (N_28945,N_26465,N_25126);
nand U28946 (N_28946,N_25722,N_26107);
nand U28947 (N_28947,N_26738,N_25341);
nand U28948 (N_28948,N_26105,N_26849);
and U28949 (N_28949,N_25672,N_24162);
or U28950 (N_28950,N_26892,N_26812);
nand U28951 (N_28951,N_26719,N_25030);
nor U28952 (N_28952,N_26474,N_26122);
or U28953 (N_28953,N_24490,N_25555);
xor U28954 (N_28954,N_25274,N_24982);
or U28955 (N_28955,N_24292,N_26396);
nand U28956 (N_28956,N_24493,N_25418);
or U28957 (N_28957,N_26324,N_26283);
nor U28958 (N_28958,N_25277,N_24287);
xnor U28959 (N_28959,N_24650,N_24265);
nand U28960 (N_28960,N_24346,N_25942);
nand U28961 (N_28961,N_26521,N_25896);
nor U28962 (N_28962,N_25247,N_24956);
or U28963 (N_28963,N_24993,N_24722);
nor U28964 (N_28964,N_26804,N_25561);
or U28965 (N_28965,N_25634,N_25808);
nand U28966 (N_28966,N_24908,N_26857);
xnor U28967 (N_28967,N_26122,N_24227);
nor U28968 (N_28968,N_24985,N_25798);
or U28969 (N_28969,N_25116,N_25702);
nand U28970 (N_28970,N_24866,N_25403);
xnor U28971 (N_28971,N_26209,N_24265);
and U28972 (N_28972,N_24863,N_26305);
and U28973 (N_28973,N_26475,N_24736);
and U28974 (N_28974,N_26111,N_24277);
nand U28975 (N_28975,N_25917,N_26304);
nor U28976 (N_28976,N_26500,N_26234);
xnor U28977 (N_28977,N_26031,N_26784);
nand U28978 (N_28978,N_25978,N_26496);
nor U28979 (N_28979,N_26030,N_25418);
nand U28980 (N_28980,N_25416,N_24869);
or U28981 (N_28981,N_24949,N_24158);
or U28982 (N_28982,N_24632,N_25657);
and U28983 (N_28983,N_25902,N_26117);
or U28984 (N_28984,N_25342,N_25380);
xnor U28985 (N_28985,N_26759,N_26417);
xnor U28986 (N_28986,N_26308,N_26304);
and U28987 (N_28987,N_25751,N_24563);
nand U28988 (N_28988,N_24965,N_24748);
xor U28989 (N_28989,N_26484,N_26338);
nor U28990 (N_28990,N_25788,N_24311);
or U28991 (N_28991,N_26768,N_25958);
xnor U28992 (N_28992,N_24626,N_25128);
xnor U28993 (N_28993,N_24602,N_24751);
or U28994 (N_28994,N_25154,N_25568);
or U28995 (N_28995,N_25704,N_26230);
or U28996 (N_28996,N_24915,N_25025);
nor U28997 (N_28997,N_26496,N_25343);
and U28998 (N_28998,N_26007,N_25344);
and U28999 (N_28999,N_26522,N_26489);
xnor U29000 (N_29000,N_26987,N_25404);
xor U29001 (N_29001,N_24651,N_25396);
nor U29002 (N_29002,N_25670,N_26645);
xnor U29003 (N_29003,N_25580,N_25681);
nor U29004 (N_29004,N_26194,N_24071);
or U29005 (N_29005,N_25311,N_25245);
nand U29006 (N_29006,N_24145,N_26047);
xor U29007 (N_29007,N_24765,N_24148);
nor U29008 (N_29008,N_25660,N_26528);
nand U29009 (N_29009,N_24620,N_24016);
nor U29010 (N_29010,N_26771,N_26607);
or U29011 (N_29011,N_25375,N_26049);
nor U29012 (N_29012,N_25001,N_24367);
or U29013 (N_29013,N_24208,N_24560);
xor U29014 (N_29014,N_26834,N_24236);
nor U29015 (N_29015,N_25861,N_26944);
and U29016 (N_29016,N_26781,N_25655);
xor U29017 (N_29017,N_24593,N_26534);
and U29018 (N_29018,N_24940,N_24434);
and U29019 (N_29019,N_25800,N_26892);
or U29020 (N_29020,N_24492,N_24797);
nor U29021 (N_29021,N_25248,N_25613);
nor U29022 (N_29022,N_25623,N_24668);
nor U29023 (N_29023,N_25364,N_25700);
nor U29024 (N_29024,N_24309,N_26303);
and U29025 (N_29025,N_26342,N_25149);
or U29026 (N_29026,N_25425,N_24393);
nor U29027 (N_29027,N_24400,N_24306);
or U29028 (N_29028,N_24100,N_25387);
and U29029 (N_29029,N_25992,N_25801);
xnor U29030 (N_29030,N_25492,N_26483);
xnor U29031 (N_29031,N_26937,N_25467);
nor U29032 (N_29032,N_25916,N_26200);
and U29033 (N_29033,N_26245,N_24850);
or U29034 (N_29034,N_25572,N_24549);
nor U29035 (N_29035,N_25964,N_26162);
nor U29036 (N_29036,N_25614,N_26068);
nor U29037 (N_29037,N_26234,N_24238);
nand U29038 (N_29038,N_26365,N_26517);
xnor U29039 (N_29039,N_24010,N_26308);
and U29040 (N_29040,N_24023,N_25251);
xor U29041 (N_29041,N_24661,N_25794);
nor U29042 (N_29042,N_26714,N_25986);
xor U29043 (N_29043,N_25116,N_25683);
nand U29044 (N_29044,N_25823,N_26365);
or U29045 (N_29045,N_25204,N_25162);
xnor U29046 (N_29046,N_24370,N_24293);
or U29047 (N_29047,N_24405,N_25972);
nor U29048 (N_29048,N_26473,N_26232);
nor U29049 (N_29049,N_25043,N_24852);
nand U29050 (N_29050,N_26029,N_24848);
nor U29051 (N_29051,N_25090,N_25357);
or U29052 (N_29052,N_24581,N_24436);
or U29053 (N_29053,N_24674,N_25218);
nand U29054 (N_29054,N_26172,N_25945);
xor U29055 (N_29055,N_25785,N_25913);
nand U29056 (N_29056,N_26723,N_25890);
nor U29057 (N_29057,N_24388,N_26198);
nor U29058 (N_29058,N_25527,N_24758);
xor U29059 (N_29059,N_24961,N_26321);
or U29060 (N_29060,N_25969,N_24199);
and U29061 (N_29061,N_26607,N_25288);
and U29062 (N_29062,N_25769,N_24813);
xor U29063 (N_29063,N_25635,N_26235);
nand U29064 (N_29064,N_26099,N_25359);
and U29065 (N_29065,N_24204,N_24460);
nor U29066 (N_29066,N_24152,N_25981);
xor U29067 (N_29067,N_24338,N_25603);
nor U29068 (N_29068,N_26182,N_26784);
xnor U29069 (N_29069,N_24833,N_25655);
nor U29070 (N_29070,N_26437,N_26416);
or U29071 (N_29071,N_24926,N_26751);
nand U29072 (N_29072,N_26728,N_24861);
or U29073 (N_29073,N_24537,N_26647);
xnor U29074 (N_29074,N_25296,N_24828);
nand U29075 (N_29075,N_26285,N_24478);
xor U29076 (N_29076,N_26508,N_26594);
nor U29077 (N_29077,N_26139,N_25953);
nor U29078 (N_29078,N_24871,N_25531);
xnor U29079 (N_29079,N_25518,N_24778);
nor U29080 (N_29080,N_26383,N_24068);
nor U29081 (N_29081,N_24916,N_25554);
and U29082 (N_29082,N_26272,N_24115);
or U29083 (N_29083,N_26484,N_24166);
or U29084 (N_29084,N_26911,N_26076);
nor U29085 (N_29085,N_24233,N_24127);
nand U29086 (N_29086,N_25017,N_26902);
and U29087 (N_29087,N_24816,N_26886);
nor U29088 (N_29088,N_26952,N_25352);
or U29089 (N_29089,N_25685,N_26222);
nor U29090 (N_29090,N_25389,N_26495);
nand U29091 (N_29091,N_25579,N_26021);
or U29092 (N_29092,N_24599,N_24125);
nor U29093 (N_29093,N_24802,N_24502);
nor U29094 (N_29094,N_24509,N_25900);
or U29095 (N_29095,N_25793,N_24574);
or U29096 (N_29096,N_26105,N_24272);
and U29097 (N_29097,N_24686,N_26022);
nor U29098 (N_29098,N_24688,N_25275);
or U29099 (N_29099,N_25029,N_25384);
and U29100 (N_29100,N_26394,N_24447);
nand U29101 (N_29101,N_25215,N_24868);
nor U29102 (N_29102,N_24112,N_25655);
nand U29103 (N_29103,N_26122,N_25324);
xor U29104 (N_29104,N_24669,N_26843);
or U29105 (N_29105,N_26303,N_26947);
nor U29106 (N_29106,N_26065,N_26796);
or U29107 (N_29107,N_24552,N_25342);
or U29108 (N_29108,N_26078,N_24006);
nor U29109 (N_29109,N_24945,N_26245);
nor U29110 (N_29110,N_25590,N_26216);
and U29111 (N_29111,N_25297,N_25978);
nor U29112 (N_29112,N_26354,N_24522);
nor U29113 (N_29113,N_25898,N_26291);
nand U29114 (N_29114,N_26016,N_24491);
nor U29115 (N_29115,N_26860,N_24333);
nand U29116 (N_29116,N_24444,N_26880);
xor U29117 (N_29117,N_26373,N_25885);
and U29118 (N_29118,N_25364,N_25831);
or U29119 (N_29119,N_24878,N_24106);
nand U29120 (N_29120,N_24690,N_26059);
or U29121 (N_29121,N_26066,N_25555);
nor U29122 (N_29122,N_26789,N_26892);
and U29123 (N_29123,N_25908,N_26369);
or U29124 (N_29124,N_26171,N_24745);
or U29125 (N_29125,N_26003,N_26030);
and U29126 (N_29126,N_26373,N_24061);
xnor U29127 (N_29127,N_24465,N_24826);
and U29128 (N_29128,N_26592,N_25835);
nand U29129 (N_29129,N_24988,N_25516);
xor U29130 (N_29130,N_25707,N_26175);
and U29131 (N_29131,N_26609,N_24778);
nor U29132 (N_29132,N_26944,N_24306);
xor U29133 (N_29133,N_26674,N_25935);
and U29134 (N_29134,N_24794,N_26113);
nand U29135 (N_29135,N_25184,N_24990);
nor U29136 (N_29136,N_25102,N_26365);
and U29137 (N_29137,N_25681,N_25267);
xor U29138 (N_29138,N_24550,N_25098);
nand U29139 (N_29139,N_25996,N_26994);
nor U29140 (N_29140,N_25186,N_26347);
nor U29141 (N_29141,N_26592,N_25053);
nand U29142 (N_29142,N_26221,N_25791);
nand U29143 (N_29143,N_24100,N_24424);
nor U29144 (N_29144,N_24379,N_25682);
nand U29145 (N_29145,N_26771,N_26499);
or U29146 (N_29146,N_24562,N_25823);
xnor U29147 (N_29147,N_26858,N_24411);
and U29148 (N_29148,N_25736,N_25297);
nand U29149 (N_29149,N_25288,N_25529);
xnor U29150 (N_29150,N_24832,N_24067);
nor U29151 (N_29151,N_26327,N_26220);
and U29152 (N_29152,N_26339,N_26629);
xor U29153 (N_29153,N_25891,N_24238);
xor U29154 (N_29154,N_25182,N_26519);
and U29155 (N_29155,N_26329,N_25864);
nor U29156 (N_29156,N_26695,N_24124);
and U29157 (N_29157,N_24489,N_24687);
nor U29158 (N_29158,N_26927,N_24344);
xnor U29159 (N_29159,N_24165,N_24486);
or U29160 (N_29160,N_24423,N_26201);
and U29161 (N_29161,N_24732,N_25900);
xnor U29162 (N_29162,N_25564,N_24252);
or U29163 (N_29163,N_26182,N_25284);
xor U29164 (N_29164,N_25705,N_24101);
and U29165 (N_29165,N_26572,N_24681);
nand U29166 (N_29166,N_25501,N_25241);
xor U29167 (N_29167,N_25328,N_25841);
nor U29168 (N_29168,N_25643,N_24831);
nand U29169 (N_29169,N_24296,N_24945);
nand U29170 (N_29170,N_25931,N_24830);
nor U29171 (N_29171,N_24984,N_25019);
and U29172 (N_29172,N_26317,N_24442);
and U29173 (N_29173,N_26851,N_26742);
nor U29174 (N_29174,N_25039,N_25105);
xnor U29175 (N_29175,N_25718,N_24858);
nor U29176 (N_29176,N_26560,N_25174);
xnor U29177 (N_29177,N_24019,N_26326);
and U29178 (N_29178,N_24484,N_26967);
xnor U29179 (N_29179,N_26512,N_25610);
and U29180 (N_29180,N_25222,N_26336);
or U29181 (N_29181,N_26522,N_26737);
xor U29182 (N_29182,N_26953,N_26701);
nor U29183 (N_29183,N_25420,N_26373);
and U29184 (N_29184,N_24703,N_24505);
nand U29185 (N_29185,N_24507,N_26258);
nor U29186 (N_29186,N_26040,N_25495);
and U29187 (N_29187,N_25304,N_26514);
nor U29188 (N_29188,N_26842,N_24011);
nor U29189 (N_29189,N_25655,N_24807);
and U29190 (N_29190,N_24032,N_24062);
nand U29191 (N_29191,N_25268,N_25039);
or U29192 (N_29192,N_25558,N_25185);
or U29193 (N_29193,N_24511,N_25658);
nor U29194 (N_29194,N_25785,N_26276);
and U29195 (N_29195,N_26974,N_26959);
nand U29196 (N_29196,N_26700,N_24004);
nand U29197 (N_29197,N_26718,N_24060);
or U29198 (N_29198,N_26939,N_25364);
xor U29199 (N_29199,N_26830,N_24433);
or U29200 (N_29200,N_24358,N_26181);
nor U29201 (N_29201,N_26359,N_24783);
or U29202 (N_29202,N_25536,N_24745);
or U29203 (N_29203,N_25765,N_25217);
or U29204 (N_29204,N_25840,N_26283);
and U29205 (N_29205,N_24926,N_24234);
nor U29206 (N_29206,N_24164,N_24388);
xor U29207 (N_29207,N_25938,N_24359);
nor U29208 (N_29208,N_25373,N_26413);
nand U29209 (N_29209,N_24116,N_25727);
nor U29210 (N_29210,N_26356,N_26522);
xor U29211 (N_29211,N_24452,N_26149);
xor U29212 (N_29212,N_25886,N_26113);
nor U29213 (N_29213,N_24359,N_25791);
nand U29214 (N_29214,N_24251,N_25030);
and U29215 (N_29215,N_26720,N_24495);
xnor U29216 (N_29216,N_24207,N_26561);
or U29217 (N_29217,N_24352,N_25337);
xnor U29218 (N_29218,N_25379,N_25047);
or U29219 (N_29219,N_24039,N_25793);
xor U29220 (N_29220,N_24040,N_25473);
nand U29221 (N_29221,N_25788,N_24143);
nand U29222 (N_29222,N_26651,N_26593);
or U29223 (N_29223,N_25308,N_26910);
or U29224 (N_29224,N_26556,N_26914);
nor U29225 (N_29225,N_25844,N_24251);
xnor U29226 (N_29226,N_24032,N_24313);
xor U29227 (N_29227,N_26999,N_25765);
xnor U29228 (N_29228,N_24221,N_26835);
or U29229 (N_29229,N_24125,N_24822);
nand U29230 (N_29230,N_26243,N_24715);
and U29231 (N_29231,N_25138,N_26800);
nor U29232 (N_29232,N_24452,N_25871);
nand U29233 (N_29233,N_26882,N_24612);
nand U29234 (N_29234,N_25402,N_26994);
nor U29235 (N_29235,N_24776,N_25285);
and U29236 (N_29236,N_25037,N_25265);
nand U29237 (N_29237,N_25489,N_24448);
or U29238 (N_29238,N_24882,N_26957);
or U29239 (N_29239,N_26003,N_24755);
nand U29240 (N_29240,N_25094,N_26514);
xor U29241 (N_29241,N_25585,N_25814);
xnor U29242 (N_29242,N_24533,N_26826);
and U29243 (N_29243,N_26125,N_25167);
nand U29244 (N_29244,N_25855,N_26932);
nor U29245 (N_29245,N_24580,N_26097);
nand U29246 (N_29246,N_25871,N_26498);
or U29247 (N_29247,N_26244,N_25598);
xnor U29248 (N_29248,N_24651,N_25669);
xnor U29249 (N_29249,N_24311,N_24918);
or U29250 (N_29250,N_24078,N_25549);
or U29251 (N_29251,N_26216,N_25925);
xnor U29252 (N_29252,N_24853,N_24715);
and U29253 (N_29253,N_24066,N_24280);
nor U29254 (N_29254,N_25609,N_25223);
or U29255 (N_29255,N_26843,N_26880);
xnor U29256 (N_29256,N_26019,N_24963);
nor U29257 (N_29257,N_26681,N_24501);
and U29258 (N_29258,N_24140,N_26467);
and U29259 (N_29259,N_26087,N_26175);
nand U29260 (N_29260,N_26104,N_24398);
nand U29261 (N_29261,N_26440,N_25730);
nor U29262 (N_29262,N_25536,N_26837);
nand U29263 (N_29263,N_26200,N_26146);
and U29264 (N_29264,N_26792,N_26492);
nand U29265 (N_29265,N_26676,N_26729);
nand U29266 (N_29266,N_24994,N_26989);
and U29267 (N_29267,N_26559,N_26051);
and U29268 (N_29268,N_24541,N_26614);
and U29269 (N_29269,N_24274,N_26357);
nor U29270 (N_29270,N_24378,N_26040);
nor U29271 (N_29271,N_26396,N_26188);
and U29272 (N_29272,N_24617,N_24277);
nor U29273 (N_29273,N_26909,N_26829);
xor U29274 (N_29274,N_25917,N_24441);
nand U29275 (N_29275,N_24898,N_25477);
nor U29276 (N_29276,N_26448,N_24070);
xnor U29277 (N_29277,N_24703,N_25087);
nor U29278 (N_29278,N_24484,N_26575);
nand U29279 (N_29279,N_26129,N_25010);
nor U29280 (N_29280,N_25658,N_25392);
and U29281 (N_29281,N_26839,N_24642);
nor U29282 (N_29282,N_24449,N_24752);
nor U29283 (N_29283,N_26185,N_24571);
xnor U29284 (N_29284,N_24219,N_25571);
nor U29285 (N_29285,N_25013,N_26350);
nand U29286 (N_29286,N_24619,N_26740);
nor U29287 (N_29287,N_26126,N_24485);
nand U29288 (N_29288,N_24545,N_26501);
xor U29289 (N_29289,N_26340,N_24570);
and U29290 (N_29290,N_26528,N_25500);
and U29291 (N_29291,N_24002,N_24479);
or U29292 (N_29292,N_25310,N_26406);
nor U29293 (N_29293,N_26953,N_24224);
and U29294 (N_29294,N_25309,N_24367);
xor U29295 (N_29295,N_24124,N_24341);
xnor U29296 (N_29296,N_25986,N_25977);
or U29297 (N_29297,N_24763,N_26819);
nor U29298 (N_29298,N_24021,N_26019);
or U29299 (N_29299,N_25165,N_26756);
and U29300 (N_29300,N_24967,N_24603);
nand U29301 (N_29301,N_25896,N_26797);
and U29302 (N_29302,N_25771,N_24480);
xor U29303 (N_29303,N_26634,N_26922);
nor U29304 (N_29304,N_24450,N_25327);
or U29305 (N_29305,N_26975,N_24382);
and U29306 (N_29306,N_24147,N_26308);
and U29307 (N_29307,N_26086,N_25858);
or U29308 (N_29308,N_24352,N_26945);
or U29309 (N_29309,N_24029,N_26937);
and U29310 (N_29310,N_26815,N_24954);
nor U29311 (N_29311,N_25801,N_26633);
nand U29312 (N_29312,N_26900,N_26453);
nand U29313 (N_29313,N_26211,N_25934);
and U29314 (N_29314,N_25056,N_26186);
and U29315 (N_29315,N_24222,N_24719);
nand U29316 (N_29316,N_24095,N_26543);
and U29317 (N_29317,N_25346,N_24141);
and U29318 (N_29318,N_26278,N_25586);
nand U29319 (N_29319,N_25348,N_24777);
and U29320 (N_29320,N_24140,N_25832);
or U29321 (N_29321,N_24272,N_25730);
xnor U29322 (N_29322,N_24284,N_24182);
or U29323 (N_29323,N_25969,N_24429);
nor U29324 (N_29324,N_25609,N_25503);
and U29325 (N_29325,N_25478,N_26467);
nor U29326 (N_29326,N_26875,N_26895);
and U29327 (N_29327,N_25747,N_24990);
nand U29328 (N_29328,N_24489,N_25242);
or U29329 (N_29329,N_25995,N_25629);
and U29330 (N_29330,N_26348,N_26850);
and U29331 (N_29331,N_26101,N_26170);
nand U29332 (N_29332,N_25020,N_25591);
xor U29333 (N_29333,N_24470,N_24123);
nor U29334 (N_29334,N_24822,N_25694);
and U29335 (N_29335,N_25495,N_25546);
nor U29336 (N_29336,N_25787,N_26212);
nand U29337 (N_29337,N_25428,N_24486);
or U29338 (N_29338,N_24811,N_24895);
and U29339 (N_29339,N_24347,N_25817);
nand U29340 (N_29340,N_26944,N_24565);
and U29341 (N_29341,N_26804,N_25418);
xor U29342 (N_29342,N_24150,N_24080);
nor U29343 (N_29343,N_26647,N_26430);
nor U29344 (N_29344,N_24402,N_26453);
nor U29345 (N_29345,N_25575,N_24505);
and U29346 (N_29346,N_24354,N_26653);
nor U29347 (N_29347,N_25396,N_25078);
nor U29348 (N_29348,N_25951,N_26262);
and U29349 (N_29349,N_24981,N_26800);
nand U29350 (N_29350,N_25964,N_24594);
nand U29351 (N_29351,N_25685,N_26651);
or U29352 (N_29352,N_26953,N_26637);
and U29353 (N_29353,N_25153,N_26667);
and U29354 (N_29354,N_24761,N_24342);
xor U29355 (N_29355,N_26590,N_24527);
or U29356 (N_29356,N_24192,N_26023);
or U29357 (N_29357,N_25878,N_25412);
xor U29358 (N_29358,N_24192,N_25808);
or U29359 (N_29359,N_24097,N_24017);
nor U29360 (N_29360,N_26737,N_24423);
nand U29361 (N_29361,N_26433,N_24808);
xor U29362 (N_29362,N_24552,N_25692);
nor U29363 (N_29363,N_25319,N_25229);
or U29364 (N_29364,N_25299,N_26098);
and U29365 (N_29365,N_25580,N_25604);
xor U29366 (N_29366,N_25575,N_24343);
nor U29367 (N_29367,N_24793,N_26849);
nand U29368 (N_29368,N_24763,N_25366);
nand U29369 (N_29369,N_26993,N_25492);
or U29370 (N_29370,N_25245,N_26255);
or U29371 (N_29371,N_25457,N_24191);
and U29372 (N_29372,N_26829,N_25194);
or U29373 (N_29373,N_25542,N_25770);
nand U29374 (N_29374,N_24236,N_26045);
and U29375 (N_29375,N_26712,N_24099);
xor U29376 (N_29376,N_24328,N_25556);
xnor U29377 (N_29377,N_26441,N_26464);
nor U29378 (N_29378,N_26824,N_25659);
xor U29379 (N_29379,N_25544,N_25913);
or U29380 (N_29380,N_24486,N_26247);
nand U29381 (N_29381,N_26829,N_24686);
and U29382 (N_29382,N_26224,N_26642);
nor U29383 (N_29383,N_25414,N_24880);
nand U29384 (N_29384,N_25983,N_25891);
xor U29385 (N_29385,N_26145,N_25100);
or U29386 (N_29386,N_25532,N_25103);
nand U29387 (N_29387,N_25886,N_24668);
or U29388 (N_29388,N_26154,N_24346);
xor U29389 (N_29389,N_26858,N_26298);
xnor U29390 (N_29390,N_26090,N_26424);
xnor U29391 (N_29391,N_26100,N_25948);
nand U29392 (N_29392,N_24326,N_24253);
xnor U29393 (N_29393,N_24487,N_24461);
or U29394 (N_29394,N_26703,N_25250);
or U29395 (N_29395,N_26199,N_25706);
nor U29396 (N_29396,N_26216,N_26289);
or U29397 (N_29397,N_24317,N_25379);
nor U29398 (N_29398,N_24531,N_25234);
xnor U29399 (N_29399,N_26578,N_26959);
or U29400 (N_29400,N_26546,N_25477);
and U29401 (N_29401,N_25244,N_24406);
and U29402 (N_29402,N_25986,N_25466);
or U29403 (N_29403,N_26443,N_26305);
nor U29404 (N_29404,N_26559,N_26311);
nor U29405 (N_29405,N_25662,N_24833);
nand U29406 (N_29406,N_25550,N_24603);
nor U29407 (N_29407,N_26922,N_26185);
nor U29408 (N_29408,N_25795,N_26523);
nor U29409 (N_29409,N_25327,N_24253);
nor U29410 (N_29410,N_24865,N_26479);
xnor U29411 (N_29411,N_26508,N_26057);
or U29412 (N_29412,N_26937,N_26165);
and U29413 (N_29413,N_24770,N_24321);
and U29414 (N_29414,N_26294,N_24509);
xnor U29415 (N_29415,N_25094,N_26169);
and U29416 (N_29416,N_24843,N_25418);
or U29417 (N_29417,N_26476,N_26037);
and U29418 (N_29418,N_26296,N_25219);
nand U29419 (N_29419,N_24424,N_24787);
nor U29420 (N_29420,N_24220,N_24675);
xnor U29421 (N_29421,N_25576,N_26489);
xnor U29422 (N_29422,N_26692,N_26703);
and U29423 (N_29423,N_26149,N_25921);
xnor U29424 (N_29424,N_24460,N_24562);
xnor U29425 (N_29425,N_25949,N_25390);
and U29426 (N_29426,N_24057,N_25333);
and U29427 (N_29427,N_26072,N_24638);
xnor U29428 (N_29428,N_25062,N_24878);
or U29429 (N_29429,N_26730,N_26647);
and U29430 (N_29430,N_26352,N_26724);
nor U29431 (N_29431,N_26517,N_26879);
nand U29432 (N_29432,N_24055,N_25479);
nor U29433 (N_29433,N_25481,N_24005);
nor U29434 (N_29434,N_24319,N_26234);
and U29435 (N_29435,N_26936,N_26459);
xnor U29436 (N_29436,N_26580,N_24250);
and U29437 (N_29437,N_26720,N_26930);
nand U29438 (N_29438,N_24793,N_25277);
nor U29439 (N_29439,N_24995,N_26122);
xnor U29440 (N_29440,N_25799,N_26426);
nor U29441 (N_29441,N_26795,N_26823);
or U29442 (N_29442,N_25681,N_25885);
nor U29443 (N_29443,N_25549,N_25853);
nand U29444 (N_29444,N_26865,N_25089);
or U29445 (N_29445,N_26181,N_26372);
or U29446 (N_29446,N_25743,N_26881);
or U29447 (N_29447,N_24941,N_26085);
and U29448 (N_29448,N_24568,N_26827);
and U29449 (N_29449,N_26396,N_25451);
and U29450 (N_29450,N_26987,N_24041);
or U29451 (N_29451,N_24815,N_25816);
nand U29452 (N_29452,N_25480,N_24139);
nand U29453 (N_29453,N_24724,N_25397);
xor U29454 (N_29454,N_25095,N_26227);
and U29455 (N_29455,N_25081,N_26059);
or U29456 (N_29456,N_25736,N_25320);
xor U29457 (N_29457,N_26377,N_26471);
and U29458 (N_29458,N_25879,N_24248);
nor U29459 (N_29459,N_26575,N_26403);
nand U29460 (N_29460,N_25958,N_24312);
nor U29461 (N_29461,N_24949,N_25909);
xor U29462 (N_29462,N_24819,N_26130);
nor U29463 (N_29463,N_25124,N_26536);
nor U29464 (N_29464,N_25425,N_26063);
nand U29465 (N_29465,N_24585,N_26750);
or U29466 (N_29466,N_25694,N_25074);
nand U29467 (N_29467,N_26811,N_26604);
or U29468 (N_29468,N_24618,N_24010);
nand U29469 (N_29469,N_26733,N_25502);
or U29470 (N_29470,N_25771,N_25634);
or U29471 (N_29471,N_25238,N_24743);
nand U29472 (N_29472,N_26389,N_26222);
nor U29473 (N_29473,N_24985,N_26182);
xnor U29474 (N_29474,N_25965,N_24890);
nor U29475 (N_29475,N_24152,N_25869);
xor U29476 (N_29476,N_26347,N_26686);
or U29477 (N_29477,N_26223,N_24277);
xnor U29478 (N_29478,N_26409,N_24332);
and U29479 (N_29479,N_25322,N_26557);
and U29480 (N_29480,N_25417,N_25084);
nand U29481 (N_29481,N_24587,N_24579);
or U29482 (N_29482,N_26307,N_24365);
nor U29483 (N_29483,N_26339,N_24870);
and U29484 (N_29484,N_25318,N_24923);
nor U29485 (N_29485,N_25062,N_24110);
nor U29486 (N_29486,N_26589,N_24228);
or U29487 (N_29487,N_25790,N_24321);
nor U29488 (N_29488,N_26563,N_26118);
or U29489 (N_29489,N_25521,N_24516);
or U29490 (N_29490,N_25265,N_26768);
and U29491 (N_29491,N_26637,N_24418);
xnor U29492 (N_29492,N_26532,N_26200);
nand U29493 (N_29493,N_25228,N_24209);
nand U29494 (N_29494,N_24579,N_24461);
and U29495 (N_29495,N_25735,N_24314);
xor U29496 (N_29496,N_24324,N_25725);
xnor U29497 (N_29497,N_26628,N_24167);
or U29498 (N_29498,N_24857,N_24017);
nand U29499 (N_29499,N_26197,N_26342);
or U29500 (N_29500,N_26686,N_25886);
or U29501 (N_29501,N_26543,N_25288);
nand U29502 (N_29502,N_26672,N_26236);
and U29503 (N_29503,N_26746,N_26595);
and U29504 (N_29504,N_24036,N_26470);
or U29505 (N_29505,N_26179,N_26787);
xnor U29506 (N_29506,N_25953,N_26840);
nand U29507 (N_29507,N_26614,N_25740);
nand U29508 (N_29508,N_24248,N_26663);
and U29509 (N_29509,N_24363,N_26755);
nor U29510 (N_29510,N_25735,N_26497);
nand U29511 (N_29511,N_25381,N_25264);
and U29512 (N_29512,N_24698,N_26868);
xor U29513 (N_29513,N_26171,N_24635);
or U29514 (N_29514,N_26077,N_25264);
nand U29515 (N_29515,N_24819,N_26828);
nand U29516 (N_29516,N_24085,N_25659);
nand U29517 (N_29517,N_24600,N_25203);
xor U29518 (N_29518,N_26163,N_24571);
and U29519 (N_29519,N_24279,N_25355);
nand U29520 (N_29520,N_26296,N_25701);
nand U29521 (N_29521,N_25476,N_24897);
nor U29522 (N_29522,N_25868,N_24898);
xnor U29523 (N_29523,N_25735,N_24587);
or U29524 (N_29524,N_26392,N_24457);
nand U29525 (N_29525,N_24051,N_24773);
xor U29526 (N_29526,N_24174,N_25824);
nand U29527 (N_29527,N_26507,N_25218);
and U29528 (N_29528,N_24712,N_26556);
or U29529 (N_29529,N_26316,N_26673);
or U29530 (N_29530,N_24409,N_26578);
xor U29531 (N_29531,N_24347,N_24164);
and U29532 (N_29532,N_24608,N_24746);
nor U29533 (N_29533,N_24647,N_25027);
xnor U29534 (N_29534,N_24906,N_25553);
nor U29535 (N_29535,N_24065,N_24724);
xor U29536 (N_29536,N_24181,N_26329);
and U29537 (N_29537,N_25228,N_24992);
xnor U29538 (N_29538,N_24784,N_25684);
or U29539 (N_29539,N_25736,N_26635);
xor U29540 (N_29540,N_25932,N_26618);
or U29541 (N_29541,N_25555,N_25662);
or U29542 (N_29542,N_26945,N_24921);
nand U29543 (N_29543,N_25432,N_26914);
xnor U29544 (N_29544,N_24135,N_25354);
or U29545 (N_29545,N_25742,N_24927);
nor U29546 (N_29546,N_26781,N_25569);
nor U29547 (N_29547,N_26144,N_24297);
xnor U29548 (N_29548,N_24575,N_24840);
and U29549 (N_29549,N_24766,N_24463);
nor U29550 (N_29550,N_26772,N_24405);
nand U29551 (N_29551,N_25113,N_24708);
and U29552 (N_29552,N_25319,N_24611);
xor U29553 (N_29553,N_26742,N_24122);
and U29554 (N_29554,N_26975,N_24955);
nor U29555 (N_29555,N_26789,N_24467);
nand U29556 (N_29556,N_25690,N_25688);
or U29557 (N_29557,N_26848,N_25738);
xor U29558 (N_29558,N_24711,N_25800);
xnor U29559 (N_29559,N_25996,N_26469);
or U29560 (N_29560,N_26425,N_24156);
nand U29561 (N_29561,N_26358,N_26166);
nand U29562 (N_29562,N_25900,N_25348);
and U29563 (N_29563,N_26170,N_25591);
xnor U29564 (N_29564,N_26929,N_26468);
and U29565 (N_29565,N_26403,N_25388);
and U29566 (N_29566,N_25059,N_24136);
nand U29567 (N_29567,N_26503,N_25864);
and U29568 (N_29568,N_24190,N_25769);
or U29569 (N_29569,N_24658,N_24860);
nor U29570 (N_29570,N_26265,N_26664);
and U29571 (N_29571,N_25321,N_26349);
nor U29572 (N_29572,N_24658,N_24938);
nor U29573 (N_29573,N_25045,N_26639);
or U29574 (N_29574,N_24812,N_25635);
xor U29575 (N_29575,N_25331,N_24333);
xor U29576 (N_29576,N_24708,N_24209);
nor U29577 (N_29577,N_24508,N_26473);
or U29578 (N_29578,N_24095,N_26141);
or U29579 (N_29579,N_25921,N_24234);
and U29580 (N_29580,N_24315,N_26338);
nand U29581 (N_29581,N_24131,N_24476);
or U29582 (N_29582,N_26527,N_25807);
nor U29583 (N_29583,N_24376,N_25873);
and U29584 (N_29584,N_25997,N_25198);
nand U29585 (N_29585,N_25356,N_24750);
nor U29586 (N_29586,N_24361,N_26160);
nand U29587 (N_29587,N_26278,N_25141);
nand U29588 (N_29588,N_26927,N_25131);
and U29589 (N_29589,N_24754,N_26741);
and U29590 (N_29590,N_26584,N_26014);
or U29591 (N_29591,N_25317,N_26345);
nand U29592 (N_29592,N_25758,N_24144);
nor U29593 (N_29593,N_25366,N_24735);
xnor U29594 (N_29594,N_25305,N_26094);
nor U29595 (N_29595,N_25719,N_25732);
nor U29596 (N_29596,N_26739,N_26281);
and U29597 (N_29597,N_26515,N_26802);
nor U29598 (N_29598,N_24454,N_25905);
nand U29599 (N_29599,N_25610,N_26371);
xor U29600 (N_29600,N_25619,N_26971);
and U29601 (N_29601,N_26552,N_25281);
and U29602 (N_29602,N_26741,N_24156);
xor U29603 (N_29603,N_25894,N_26575);
and U29604 (N_29604,N_26786,N_26171);
and U29605 (N_29605,N_24458,N_24790);
or U29606 (N_29606,N_26271,N_24939);
xnor U29607 (N_29607,N_26756,N_26177);
and U29608 (N_29608,N_26142,N_25124);
nand U29609 (N_29609,N_25493,N_24401);
nand U29610 (N_29610,N_26810,N_25850);
nand U29611 (N_29611,N_26928,N_24895);
nand U29612 (N_29612,N_26661,N_26574);
and U29613 (N_29613,N_24170,N_25764);
xnor U29614 (N_29614,N_25769,N_25778);
xor U29615 (N_29615,N_25912,N_24929);
and U29616 (N_29616,N_25567,N_25507);
nand U29617 (N_29617,N_24738,N_26497);
nand U29618 (N_29618,N_26166,N_25689);
nor U29619 (N_29619,N_26262,N_25968);
and U29620 (N_29620,N_24549,N_26898);
and U29621 (N_29621,N_25646,N_26794);
xor U29622 (N_29622,N_25764,N_24007);
nand U29623 (N_29623,N_25244,N_26740);
xor U29624 (N_29624,N_24465,N_25530);
and U29625 (N_29625,N_25765,N_24001);
nand U29626 (N_29626,N_24584,N_25745);
xor U29627 (N_29627,N_26501,N_24531);
nand U29628 (N_29628,N_24245,N_24823);
nand U29629 (N_29629,N_24326,N_25797);
nor U29630 (N_29630,N_24955,N_26733);
xor U29631 (N_29631,N_26454,N_26886);
xor U29632 (N_29632,N_26803,N_26032);
and U29633 (N_29633,N_24087,N_24675);
and U29634 (N_29634,N_25693,N_25700);
nand U29635 (N_29635,N_24923,N_24679);
nor U29636 (N_29636,N_26150,N_26998);
and U29637 (N_29637,N_25904,N_25308);
and U29638 (N_29638,N_26270,N_25510);
and U29639 (N_29639,N_24185,N_25828);
or U29640 (N_29640,N_25650,N_26900);
and U29641 (N_29641,N_25096,N_25887);
nor U29642 (N_29642,N_25879,N_26583);
or U29643 (N_29643,N_24983,N_26568);
or U29644 (N_29644,N_26783,N_25646);
xnor U29645 (N_29645,N_26823,N_25449);
nand U29646 (N_29646,N_26720,N_24644);
nor U29647 (N_29647,N_26817,N_25600);
nand U29648 (N_29648,N_25679,N_24120);
nor U29649 (N_29649,N_26990,N_26964);
nand U29650 (N_29650,N_26930,N_26099);
and U29651 (N_29651,N_24900,N_25190);
xor U29652 (N_29652,N_24799,N_24295);
and U29653 (N_29653,N_25924,N_25678);
and U29654 (N_29654,N_25423,N_25116);
nand U29655 (N_29655,N_26896,N_25630);
and U29656 (N_29656,N_24623,N_26984);
and U29657 (N_29657,N_25489,N_26301);
or U29658 (N_29658,N_25778,N_25562);
and U29659 (N_29659,N_26471,N_24783);
nor U29660 (N_29660,N_24847,N_24969);
nor U29661 (N_29661,N_26858,N_25593);
nor U29662 (N_29662,N_26532,N_26090);
nor U29663 (N_29663,N_24305,N_25115);
or U29664 (N_29664,N_24719,N_26643);
xnor U29665 (N_29665,N_24534,N_26593);
nor U29666 (N_29666,N_24485,N_25467);
nor U29667 (N_29667,N_24778,N_24648);
nand U29668 (N_29668,N_26822,N_24261);
and U29669 (N_29669,N_25357,N_26122);
or U29670 (N_29670,N_25244,N_24944);
xnor U29671 (N_29671,N_26168,N_25635);
and U29672 (N_29672,N_24461,N_24092);
nand U29673 (N_29673,N_26663,N_24405);
xor U29674 (N_29674,N_24963,N_26669);
nand U29675 (N_29675,N_25757,N_26371);
nand U29676 (N_29676,N_24976,N_25019);
and U29677 (N_29677,N_25420,N_26897);
nor U29678 (N_29678,N_25856,N_24153);
or U29679 (N_29679,N_25493,N_26075);
nor U29680 (N_29680,N_25705,N_26803);
nor U29681 (N_29681,N_24327,N_26280);
and U29682 (N_29682,N_26209,N_24435);
nand U29683 (N_29683,N_25911,N_25798);
and U29684 (N_29684,N_26263,N_25754);
and U29685 (N_29685,N_24652,N_26369);
and U29686 (N_29686,N_25575,N_26076);
or U29687 (N_29687,N_26882,N_25901);
xnor U29688 (N_29688,N_26717,N_25366);
nand U29689 (N_29689,N_26378,N_25992);
nand U29690 (N_29690,N_26920,N_26666);
nor U29691 (N_29691,N_26735,N_26544);
or U29692 (N_29692,N_26792,N_24063);
nand U29693 (N_29693,N_26186,N_25882);
and U29694 (N_29694,N_24175,N_24731);
or U29695 (N_29695,N_26987,N_25660);
nor U29696 (N_29696,N_26870,N_26066);
or U29697 (N_29697,N_25645,N_25121);
nor U29698 (N_29698,N_24894,N_26691);
and U29699 (N_29699,N_25750,N_26088);
xnor U29700 (N_29700,N_25648,N_25716);
and U29701 (N_29701,N_24999,N_24101);
or U29702 (N_29702,N_26369,N_25874);
xor U29703 (N_29703,N_26708,N_26345);
xnor U29704 (N_29704,N_24726,N_25229);
and U29705 (N_29705,N_26332,N_26983);
and U29706 (N_29706,N_25547,N_24454);
xnor U29707 (N_29707,N_25214,N_25485);
nor U29708 (N_29708,N_24576,N_26024);
xnor U29709 (N_29709,N_24175,N_25452);
and U29710 (N_29710,N_24523,N_24521);
or U29711 (N_29711,N_24645,N_25284);
and U29712 (N_29712,N_25331,N_25094);
nor U29713 (N_29713,N_26820,N_26172);
and U29714 (N_29714,N_25972,N_25859);
nor U29715 (N_29715,N_25062,N_24188);
and U29716 (N_29716,N_26128,N_25503);
xor U29717 (N_29717,N_26020,N_25364);
nand U29718 (N_29718,N_26348,N_26569);
nor U29719 (N_29719,N_24199,N_25141);
and U29720 (N_29720,N_26100,N_24108);
xnor U29721 (N_29721,N_25326,N_24129);
or U29722 (N_29722,N_25712,N_26993);
nand U29723 (N_29723,N_26753,N_24288);
or U29724 (N_29724,N_25432,N_24971);
and U29725 (N_29725,N_26900,N_25969);
xnor U29726 (N_29726,N_25184,N_26362);
nor U29727 (N_29727,N_25916,N_26822);
nand U29728 (N_29728,N_26757,N_25445);
and U29729 (N_29729,N_24894,N_25132);
nor U29730 (N_29730,N_26332,N_26272);
nand U29731 (N_29731,N_24455,N_24460);
or U29732 (N_29732,N_26274,N_24839);
nand U29733 (N_29733,N_25239,N_25217);
and U29734 (N_29734,N_24340,N_25778);
or U29735 (N_29735,N_24610,N_26104);
nand U29736 (N_29736,N_26956,N_24146);
xor U29737 (N_29737,N_26997,N_26237);
or U29738 (N_29738,N_24565,N_24628);
or U29739 (N_29739,N_25344,N_24090);
xor U29740 (N_29740,N_25608,N_25468);
or U29741 (N_29741,N_24656,N_26049);
and U29742 (N_29742,N_24340,N_25680);
or U29743 (N_29743,N_26592,N_25993);
or U29744 (N_29744,N_26919,N_24826);
nand U29745 (N_29745,N_26645,N_25745);
nand U29746 (N_29746,N_26386,N_24879);
and U29747 (N_29747,N_25450,N_24707);
or U29748 (N_29748,N_25280,N_25560);
nor U29749 (N_29749,N_26710,N_25976);
xor U29750 (N_29750,N_26800,N_24767);
or U29751 (N_29751,N_24633,N_25937);
or U29752 (N_29752,N_25691,N_25339);
nand U29753 (N_29753,N_25798,N_26590);
nand U29754 (N_29754,N_26662,N_26840);
nor U29755 (N_29755,N_25772,N_26297);
nor U29756 (N_29756,N_24506,N_25733);
nor U29757 (N_29757,N_26375,N_25996);
nand U29758 (N_29758,N_25862,N_25686);
and U29759 (N_29759,N_26818,N_24923);
nor U29760 (N_29760,N_26361,N_25056);
nor U29761 (N_29761,N_25890,N_25440);
and U29762 (N_29762,N_25801,N_26746);
nor U29763 (N_29763,N_25054,N_26082);
nor U29764 (N_29764,N_26059,N_26931);
and U29765 (N_29765,N_26090,N_26726);
or U29766 (N_29766,N_25395,N_24125);
nand U29767 (N_29767,N_25975,N_25143);
or U29768 (N_29768,N_24051,N_25731);
or U29769 (N_29769,N_24560,N_25049);
and U29770 (N_29770,N_26520,N_26603);
and U29771 (N_29771,N_24288,N_24735);
or U29772 (N_29772,N_25462,N_24431);
or U29773 (N_29773,N_26170,N_25343);
or U29774 (N_29774,N_25557,N_24378);
nand U29775 (N_29775,N_24901,N_26128);
xor U29776 (N_29776,N_26968,N_24466);
and U29777 (N_29777,N_25562,N_25657);
nor U29778 (N_29778,N_24122,N_25162);
nand U29779 (N_29779,N_26774,N_24454);
and U29780 (N_29780,N_24057,N_26537);
xnor U29781 (N_29781,N_25097,N_26633);
xnor U29782 (N_29782,N_24275,N_24321);
and U29783 (N_29783,N_24209,N_26446);
xnor U29784 (N_29784,N_25161,N_26938);
or U29785 (N_29785,N_25025,N_25083);
and U29786 (N_29786,N_26039,N_25167);
xnor U29787 (N_29787,N_24457,N_24288);
xnor U29788 (N_29788,N_25028,N_24559);
xnor U29789 (N_29789,N_26213,N_25865);
xnor U29790 (N_29790,N_24764,N_24859);
nor U29791 (N_29791,N_26040,N_25403);
nand U29792 (N_29792,N_25907,N_24776);
nor U29793 (N_29793,N_25616,N_25154);
nor U29794 (N_29794,N_26471,N_25871);
and U29795 (N_29795,N_26232,N_25330);
nor U29796 (N_29796,N_24383,N_24127);
and U29797 (N_29797,N_24441,N_24380);
nor U29798 (N_29798,N_25106,N_25482);
nand U29799 (N_29799,N_26983,N_25845);
nand U29800 (N_29800,N_26564,N_26843);
xor U29801 (N_29801,N_26473,N_25897);
nand U29802 (N_29802,N_26762,N_26892);
nand U29803 (N_29803,N_24378,N_25799);
nor U29804 (N_29804,N_24421,N_24188);
and U29805 (N_29805,N_26771,N_26615);
and U29806 (N_29806,N_24539,N_26504);
or U29807 (N_29807,N_25122,N_26614);
or U29808 (N_29808,N_26284,N_24720);
xnor U29809 (N_29809,N_24280,N_26901);
nor U29810 (N_29810,N_26533,N_25644);
xnor U29811 (N_29811,N_24246,N_24773);
and U29812 (N_29812,N_24007,N_25902);
nand U29813 (N_29813,N_25392,N_26737);
and U29814 (N_29814,N_24133,N_24801);
nor U29815 (N_29815,N_26658,N_25306);
xnor U29816 (N_29816,N_24086,N_25768);
nand U29817 (N_29817,N_26369,N_25603);
nor U29818 (N_29818,N_26230,N_26888);
and U29819 (N_29819,N_25234,N_24698);
and U29820 (N_29820,N_26316,N_25393);
xnor U29821 (N_29821,N_26286,N_24705);
xor U29822 (N_29822,N_25664,N_24264);
and U29823 (N_29823,N_26653,N_24205);
or U29824 (N_29824,N_26986,N_25660);
nor U29825 (N_29825,N_25691,N_24603);
and U29826 (N_29826,N_26264,N_24793);
nand U29827 (N_29827,N_25244,N_26800);
and U29828 (N_29828,N_26411,N_25997);
or U29829 (N_29829,N_24118,N_25418);
or U29830 (N_29830,N_24746,N_25021);
nor U29831 (N_29831,N_26320,N_25183);
nand U29832 (N_29832,N_24046,N_25326);
nor U29833 (N_29833,N_26238,N_24254);
xor U29834 (N_29834,N_25894,N_26033);
xor U29835 (N_29835,N_26777,N_24248);
nand U29836 (N_29836,N_25688,N_24801);
nor U29837 (N_29837,N_24599,N_24001);
and U29838 (N_29838,N_24270,N_26996);
and U29839 (N_29839,N_26864,N_24729);
xnor U29840 (N_29840,N_25455,N_24850);
and U29841 (N_29841,N_25249,N_26510);
nand U29842 (N_29842,N_26747,N_26175);
nor U29843 (N_29843,N_24598,N_26183);
and U29844 (N_29844,N_25184,N_24816);
nand U29845 (N_29845,N_26737,N_24604);
and U29846 (N_29846,N_24317,N_26006);
nand U29847 (N_29847,N_26318,N_24624);
or U29848 (N_29848,N_24621,N_25818);
nor U29849 (N_29849,N_25660,N_25450);
or U29850 (N_29850,N_24838,N_25113);
or U29851 (N_29851,N_24625,N_26218);
nand U29852 (N_29852,N_25835,N_26451);
or U29853 (N_29853,N_26970,N_26763);
and U29854 (N_29854,N_26473,N_25726);
nand U29855 (N_29855,N_24042,N_26823);
and U29856 (N_29856,N_26762,N_25307);
or U29857 (N_29857,N_26898,N_25773);
xnor U29858 (N_29858,N_25014,N_24344);
nor U29859 (N_29859,N_26873,N_26517);
nor U29860 (N_29860,N_24505,N_26202);
or U29861 (N_29861,N_26956,N_24239);
nand U29862 (N_29862,N_25602,N_26654);
or U29863 (N_29863,N_24370,N_24633);
nor U29864 (N_29864,N_25633,N_26377);
xor U29865 (N_29865,N_25320,N_24412);
nand U29866 (N_29866,N_25649,N_26376);
nor U29867 (N_29867,N_26239,N_25160);
nor U29868 (N_29868,N_24975,N_26728);
or U29869 (N_29869,N_26938,N_24077);
xnor U29870 (N_29870,N_24576,N_25054);
and U29871 (N_29871,N_25447,N_24144);
nor U29872 (N_29872,N_26748,N_26456);
xnor U29873 (N_29873,N_26898,N_25579);
or U29874 (N_29874,N_25602,N_26628);
nand U29875 (N_29875,N_25198,N_25447);
nand U29876 (N_29876,N_24042,N_25719);
nand U29877 (N_29877,N_25006,N_24420);
nand U29878 (N_29878,N_25180,N_26685);
nand U29879 (N_29879,N_26424,N_26392);
nor U29880 (N_29880,N_24170,N_25811);
nand U29881 (N_29881,N_25474,N_25057);
xor U29882 (N_29882,N_26168,N_26477);
xor U29883 (N_29883,N_24666,N_26190);
and U29884 (N_29884,N_26333,N_24394);
nor U29885 (N_29885,N_24664,N_26024);
nor U29886 (N_29886,N_25820,N_24804);
and U29887 (N_29887,N_25810,N_24015);
xor U29888 (N_29888,N_25290,N_24430);
nor U29889 (N_29889,N_26729,N_26949);
or U29890 (N_29890,N_25670,N_26280);
xnor U29891 (N_29891,N_25075,N_26695);
nor U29892 (N_29892,N_25628,N_26456);
nand U29893 (N_29893,N_25715,N_25906);
nor U29894 (N_29894,N_26947,N_25629);
and U29895 (N_29895,N_24172,N_25765);
nand U29896 (N_29896,N_26355,N_26765);
xnor U29897 (N_29897,N_26841,N_24275);
xor U29898 (N_29898,N_25531,N_25150);
and U29899 (N_29899,N_25379,N_24557);
nand U29900 (N_29900,N_25925,N_25508);
nand U29901 (N_29901,N_24139,N_24474);
and U29902 (N_29902,N_24710,N_26956);
nor U29903 (N_29903,N_24359,N_24750);
xor U29904 (N_29904,N_24375,N_25199);
nand U29905 (N_29905,N_26909,N_26413);
and U29906 (N_29906,N_25517,N_26745);
nand U29907 (N_29907,N_26635,N_24658);
xnor U29908 (N_29908,N_24062,N_24105);
nor U29909 (N_29909,N_24751,N_26659);
nand U29910 (N_29910,N_24404,N_25149);
or U29911 (N_29911,N_25196,N_24194);
or U29912 (N_29912,N_25787,N_25094);
or U29913 (N_29913,N_25797,N_26350);
nand U29914 (N_29914,N_26120,N_25476);
nand U29915 (N_29915,N_26273,N_25233);
nand U29916 (N_29916,N_25378,N_24422);
nand U29917 (N_29917,N_26035,N_25559);
and U29918 (N_29918,N_26955,N_24178);
xnor U29919 (N_29919,N_26317,N_24529);
and U29920 (N_29920,N_24339,N_26067);
or U29921 (N_29921,N_26613,N_26859);
or U29922 (N_29922,N_25211,N_25479);
xnor U29923 (N_29923,N_26692,N_26381);
or U29924 (N_29924,N_25202,N_26451);
nor U29925 (N_29925,N_26767,N_24594);
or U29926 (N_29926,N_24258,N_25082);
and U29927 (N_29927,N_25924,N_24793);
or U29928 (N_29928,N_24897,N_24117);
nand U29929 (N_29929,N_25861,N_24455);
or U29930 (N_29930,N_26914,N_26436);
and U29931 (N_29931,N_26508,N_26495);
and U29932 (N_29932,N_26213,N_24421);
xnor U29933 (N_29933,N_24612,N_26865);
nand U29934 (N_29934,N_26830,N_26097);
or U29935 (N_29935,N_25969,N_25767);
nor U29936 (N_29936,N_26934,N_24603);
and U29937 (N_29937,N_26708,N_25728);
nand U29938 (N_29938,N_25798,N_26317);
xnor U29939 (N_29939,N_26274,N_26952);
xnor U29940 (N_29940,N_26071,N_25820);
xor U29941 (N_29941,N_25083,N_24066);
or U29942 (N_29942,N_24099,N_26940);
or U29943 (N_29943,N_25848,N_26811);
xor U29944 (N_29944,N_26190,N_25460);
or U29945 (N_29945,N_25787,N_25006);
nor U29946 (N_29946,N_25966,N_25573);
and U29947 (N_29947,N_26437,N_25681);
and U29948 (N_29948,N_24275,N_25525);
nand U29949 (N_29949,N_24881,N_25056);
xnor U29950 (N_29950,N_26402,N_25035);
and U29951 (N_29951,N_24327,N_25116);
nand U29952 (N_29952,N_24237,N_24926);
nor U29953 (N_29953,N_24072,N_26109);
xor U29954 (N_29954,N_25480,N_25000);
xnor U29955 (N_29955,N_26728,N_24636);
xor U29956 (N_29956,N_26197,N_24826);
nand U29957 (N_29957,N_24098,N_25101);
or U29958 (N_29958,N_24064,N_25251);
and U29959 (N_29959,N_26173,N_26070);
nand U29960 (N_29960,N_24138,N_24075);
nand U29961 (N_29961,N_25948,N_26020);
nor U29962 (N_29962,N_24398,N_24022);
and U29963 (N_29963,N_26193,N_26618);
xor U29964 (N_29964,N_24094,N_24192);
xor U29965 (N_29965,N_24305,N_24243);
nor U29966 (N_29966,N_24462,N_25999);
nor U29967 (N_29967,N_25459,N_25243);
xor U29968 (N_29968,N_26175,N_25015);
nand U29969 (N_29969,N_24351,N_25015);
and U29970 (N_29970,N_26897,N_25314);
and U29971 (N_29971,N_26405,N_25314);
nand U29972 (N_29972,N_24573,N_26143);
xnor U29973 (N_29973,N_26557,N_25684);
and U29974 (N_29974,N_25929,N_25363);
xor U29975 (N_29975,N_26781,N_26114);
and U29976 (N_29976,N_26040,N_24542);
xor U29977 (N_29977,N_26295,N_25280);
xnor U29978 (N_29978,N_26694,N_25940);
nor U29979 (N_29979,N_24555,N_25050);
or U29980 (N_29980,N_26840,N_25310);
and U29981 (N_29981,N_24376,N_24343);
or U29982 (N_29982,N_25256,N_26869);
nand U29983 (N_29983,N_25861,N_25619);
nor U29984 (N_29984,N_24376,N_25409);
or U29985 (N_29985,N_24047,N_25936);
nor U29986 (N_29986,N_25808,N_24052);
or U29987 (N_29987,N_25849,N_25428);
nor U29988 (N_29988,N_25817,N_25867);
and U29989 (N_29989,N_24269,N_26550);
nor U29990 (N_29990,N_24570,N_24545);
nor U29991 (N_29991,N_25391,N_26562);
or U29992 (N_29992,N_24334,N_24079);
or U29993 (N_29993,N_25487,N_25713);
xnor U29994 (N_29994,N_25645,N_24923);
and U29995 (N_29995,N_24517,N_26510);
nand U29996 (N_29996,N_26677,N_26100);
xnor U29997 (N_29997,N_25609,N_26763);
nor U29998 (N_29998,N_25271,N_24437);
nor U29999 (N_29999,N_24113,N_24918);
nand UO_0 (O_0,N_27828,N_27355);
xor UO_1 (O_1,N_28274,N_28466);
nor UO_2 (O_2,N_29915,N_27904);
or UO_3 (O_3,N_29634,N_29792);
or UO_4 (O_4,N_27915,N_27054);
or UO_5 (O_5,N_27771,N_27881);
or UO_6 (O_6,N_27349,N_27795);
nor UO_7 (O_7,N_28362,N_28069);
nor UO_8 (O_8,N_28027,N_29407);
and UO_9 (O_9,N_28773,N_27197);
xnor UO_10 (O_10,N_28646,N_28864);
nand UO_11 (O_11,N_28538,N_29283);
or UO_12 (O_12,N_27065,N_27799);
or UO_13 (O_13,N_28517,N_28312);
or UO_14 (O_14,N_27929,N_28869);
nand UO_15 (O_15,N_27069,N_28028);
nand UO_16 (O_16,N_28917,N_29472);
nand UO_17 (O_17,N_28014,N_28657);
xnor UO_18 (O_18,N_29450,N_27288);
nand UO_19 (O_19,N_29344,N_27954);
and UO_20 (O_20,N_28151,N_28201);
nand UO_21 (O_21,N_27606,N_27284);
and UO_22 (O_22,N_27143,N_29107);
or UO_23 (O_23,N_29695,N_27147);
and UO_24 (O_24,N_28039,N_29958);
nand UO_25 (O_25,N_27180,N_29434);
or UO_26 (O_26,N_29805,N_29370);
nand UO_27 (O_27,N_27531,N_29252);
and UO_28 (O_28,N_29365,N_27549);
or UO_29 (O_29,N_29035,N_28254);
or UO_30 (O_30,N_27872,N_29826);
nand UO_31 (O_31,N_29421,N_29622);
or UO_32 (O_32,N_27047,N_29770);
xor UO_33 (O_33,N_29335,N_27938);
xnor UO_34 (O_34,N_27420,N_27607);
nand UO_35 (O_35,N_27746,N_29813);
nor UO_36 (O_36,N_29464,N_28695);
or UO_37 (O_37,N_27679,N_27485);
nor UO_38 (O_38,N_27983,N_28992);
nor UO_39 (O_39,N_28862,N_29470);
xnor UO_40 (O_40,N_27913,N_29295);
and UO_41 (O_41,N_28412,N_29497);
xnor UO_42 (O_42,N_28086,N_29588);
nor UO_43 (O_43,N_27968,N_28831);
or UO_44 (O_44,N_27684,N_28943);
nand UO_45 (O_45,N_29843,N_29362);
or UO_46 (O_46,N_29153,N_29590);
xnor UO_47 (O_47,N_28623,N_29156);
or UO_48 (O_48,N_27481,N_29898);
nand UO_49 (O_49,N_28873,N_27240);
nand UO_50 (O_50,N_29929,N_28867);
xnor UO_51 (O_51,N_28585,N_28540);
and UO_52 (O_52,N_28394,N_27412);
nand UO_53 (O_53,N_28922,N_28977);
or UO_54 (O_54,N_27472,N_28562);
and UO_55 (O_55,N_29614,N_29419);
and UO_56 (O_56,N_27057,N_27505);
xor UO_57 (O_57,N_28127,N_28124);
xor UO_58 (O_58,N_29998,N_28559);
nor UO_59 (O_59,N_29664,N_27347);
xor UO_60 (O_60,N_29267,N_27437);
xnor UO_61 (O_61,N_28987,N_28146);
and UO_62 (O_62,N_28512,N_28927);
nor UO_63 (O_63,N_28957,N_29908);
or UO_64 (O_64,N_27368,N_29255);
or UO_65 (O_65,N_28181,N_27643);
xnor UO_66 (O_66,N_28104,N_28207);
nor UO_67 (O_67,N_28829,N_27579);
nor UO_68 (O_68,N_27304,N_27011);
nor UO_69 (O_69,N_29055,N_27092);
nor UO_70 (O_70,N_27949,N_29961);
and UO_71 (O_71,N_27491,N_29866);
xor UO_72 (O_72,N_27845,N_27093);
nand UO_73 (O_73,N_27246,N_29340);
or UO_74 (O_74,N_28598,N_28488);
nand UO_75 (O_75,N_27713,N_28091);
and UO_76 (O_76,N_27022,N_29905);
nand UO_77 (O_77,N_27910,N_28492);
nand UO_78 (O_78,N_29538,N_27609);
nor UO_79 (O_79,N_27757,N_27478);
xnor UO_80 (O_80,N_29587,N_28659);
xor UO_81 (O_81,N_29988,N_28705);
xnor UO_82 (O_82,N_28483,N_29900);
xor UO_83 (O_83,N_27149,N_27048);
or UO_84 (O_84,N_28555,N_28527);
and UO_85 (O_85,N_28473,N_29330);
nand UO_86 (O_86,N_29842,N_29973);
xor UO_87 (O_87,N_28843,N_29563);
and UO_88 (O_88,N_28134,N_28637);
and UO_89 (O_89,N_27561,N_29662);
or UO_90 (O_90,N_28071,N_28001);
nand UO_91 (O_91,N_27600,N_29269);
and UO_92 (O_92,N_27411,N_29561);
or UO_93 (O_93,N_29305,N_28257);
nand UO_94 (O_94,N_29226,N_27948);
or UO_95 (O_95,N_28894,N_28851);
nor UO_96 (O_96,N_29606,N_27423);
xor UO_97 (O_97,N_29720,N_28836);
nand UO_98 (O_98,N_29965,N_28696);
nand UO_99 (O_99,N_29122,N_27375);
and UO_100 (O_100,N_29241,N_29240);
and UO_101 (O_101,N_28444,N_27178);
nor UO_102 (O_102,N_28465,N_29747);
nand UO_103 (O_103,N_27840,N_29387);
nor UO_104 (O_104,N_27519,N_29758);
and UO_105 (O_105,N_27348,N_27198);
xor UO_106 (O_106,N_27639,N_28744);
nand UO_107 (O_107,N_29672,N_28842);
or UO_108 (O_108,N_29498,N_27435);
nand UO_109 (O_109,N_27283,N_27729);
or UO_110 (O_110,N_28322,N_29475);
and UO_111 (O_111,N_29086,N_29506);
xnor UO_112 (O_112,N_27131,N_27865);
and UO_113 (O_113,N_29835,N_29056);
nor UO_114 (O_114,N_27596,N_29219);
and UO_115 (O_115,N_28626,N_29490);
nand UO_116 (O_116,N_28248,N_28338);
nand UO_117 (O_117,N_28478,N_29266);
nand UO_118 (O_118,N_29531,N_28010);
or UO_119 (O_119,N_28184,N_29595);
nor UO_120 (O_120,N_27803,N_28948);
xnor UO_121 (O_121,N_27926,N_27170);
and UO_122 (O_122,N_28963,N_27381);
or UO_123 (O_123,N_27253,N_29479);
nand UO_124 (O_124,N_27043,N_27547);
xor UO_125 (O_125,N_27853,N_29336);
and UO_126 (O_126,N_27740,N_27784);
nand UO_127 (O_127,N_29778,N_28431);
nand UO_128 (O_128,N_29856,N_29947);
xnor UO_129 (O_129,N_29142,N_28343);
nand UO_130 (O_130,N_27279,N_28956);
or UO_131 (O_131,N_28183,N_29967);
or UO_132 (O_132,N_28614,N_27203);
or UO_133 (O_133,N_27138,N_29771);
nor UO_134 (O_134,N_28164,N_27275);
nor UO_135 (O_135,N_27085,N_28721);
nor UO_136 (O_136,N_29458,N_28346);
xor UO_137 (O_137,N_27134,N_27861);
or UO_138 (O_138,N_28653,N_29936);
and UO_139 (O_139,N_27651,N_29129);
nor UO_140 (O_140,N_29567,N_29041);
nand UO_141 (O_141,N_28405,N_29050);
or UO_142 (O_142,N_27438,N_27739);
xnor UO_143 (O_143,N_28266,N_28472);
nor UO_144 (O_144,N_27712,N_29933);
nor UO_145 (O_145,N_28803,N_27500);
and UO_146 (O_146,N_28032,N_27220);
or UO_147 (O_147,N_29348,N_29512);
or UO_148 (O_148,N_27779,N_29053);
or UO_149 (O_149,N_27414,N_27082);
nor UO_150 (O_150,N_28938,N_28441);
xnor UO_151 (O_151,N_29198,N_28616);
nor UO_152 (O_152,N_27939,N_29289);
or UO_153 (O_153,N_27802,N_29399);
nand UO_154 (O_154,N_28462,N_29482);
nand UO_155 (O_155,N_27492,N_27666);
xor UO_156 (O_156,N_29070,N_27272);
nor UO_157 (O_157,N_27855,N_29465);
and UO_158 (O_158,N_27695,N_27574);
and UO_159 (O_159,N_29769,N_29124);
and UO_160 (O_160,N_29510,N_29751);
xor UO_161 (O_161,N_27632,N_27690);
and UO_162 (O_162,N_27829,N_29048);
xor UO_163 (O_163,N_28357,N_29701);
nand UO_164 (O_164,N_29331,N_29426);
nor UO_165 (O_165,N_28299,N_29786);
nor UO_166 (O_166,N_29678,N_29794);
nand UO_167 (O_167,N_28844,N_29889);
xnor UO_168 (O_168,N_27526,N_27384);
and UO_169 (O_169,N_29609,N_27979);
nand UO_170 (O_170,N_28752,N_28931);
nand UO_171 (O_171,N_28258,N_27141);
nor UO_172 (O_172,N_28451,N_27852);
nor UO_173 (O_173,N_28973,N_29101);
nor UO_174 (O_174,N_28656,N_29621);
xnor UO_175 (O_175,N_29602,N_29864);
and UO_176 (O_176,N_29183,N_28413);
xnor UO_177 (O_177,N_29140,N_29368);
nor UO_178 (O_178,N_29317,N_28120);
nor UO_179 (O_179,N_27707,N_27517);
nor UO_180 (O_180,N_28751,N_27495);
or UO_181 (O_181,N_28092,N_28447);
nor UO_182 (O_182,N_29447,N_27184);
xor UO_183 (O_183,N_29028,N_29733);
nor UO_184 (O_184,N_28410,N_29617);
xor UO_185 (O_185,N_28971,N_29298);
nand UO_186 (O_186,N_27833,N_28967);
nor UO_187 (O_187,N_29078,N_28731);
nand UO_188 (O_188,N_28255,N_27075);
xor UO_189 (O_189,N_29554,N_28541);
nor UO_190 (O_190,N_27996,N_29005);
nand UO_191 (O_191,N_29626,N_29815);
or UO_192 (O_192,N_28595,N_28321);
or UO_193 (O_193,N_28213,N_29945);
and UO_194 (O_194,N_27940,N_28514);
nand UO_195 (O_195,N_27775,N_27274);
nor UO_196 (O_196,N_27417,N_29741);
and UO_197 (O_197,N_28423,N_28935);
and UO_198 (O_198,N_27094,N_28619);
nor UO_199 (O_199,N_28220,N_27677);
xor UO_200 (O_200,N_29740,N_28966);
or UO_201 (O_201,N_27339,N_29364);
or UO_202 (O_202,N_29023,N_27313);
or UO_203 (O_203,N_28883,N_27837);
or UO_204 (O_204,N_29990,N_28141);
or UO_205 (O_205,N_29062,N_28895);
or UO_206 (O_206,N_28436,N_29222);
and UO_207 (O_207,N_28211,N_29310);
nand UO_208 (O_208,N_27953,N_27107);
xnor UO_209 (O_209,N_28530,N_28769);
and UO_210 (O_210,N_28205,N_27422);
nor UO_211 (O_211,N_29804,N_28772);
nor UO_212 (O_212,N_27498,N_27287);
nand UO_213 (O_213,N_28041,N_29890);
xor UO_214 (O_214,N_29956,N_28763);
and UO_215 (O_215,N_29111,N_28794);
nor UO_216 (O_216,N_28226,N_29011);
and UO_217 (O_217,N_28972,N_29322);
nand UO_218 (O_218,N_28665,N_29233);
xnor UO_219 (O_219,N_28936,N_29109);
and UO_220 (O_220,N_28275,N_27760);
nand UO_221 (O_221,N_28556,N_27682);
or UO_222 (O_222,N_27187,N_27545);
and UO_223 (O_223,N_29359,N_27496);
and UO_224 (O_224,N_28100,N_28951);
nand UO_225 (O_225,N_27937,N_28612);
nor UO_226 (O_226,N_27127,N_28398);
xor UO_227 (O_227,N_29392,N_27614);
nand UO_228 (O_228,N_27504,N_29756);
and UO_229 (O_229,N_27398,N_29524);
nand UO_230 (O_230,N_27997,N_28233);
xor UO_231 (O_231,N_28073,N_29928);
nor UO_232 (O_232,N_27860,N_29635);
nand UO_233 (O_233,N_29025,N_29120);
xnor UO_234 (O_234,N_28040,N_27534);
nand UO_235 (O_235,N_27362,N_27158);
nand UO_236 (O_236,N_29073,N_27925);
or UO_237 (O_237,N_28680,N_27215);
nor UO_238 (O_238,N_28425,N_28250);
or UO_239 (O_239,N_28793,N_27192);
nand UO_240 (O_240,N_28663,N_28349);
nand UO_241 (O_241,N_29227,N_27708);
or UO_242 (O_242,N_27693,N_28900);
and UO_243 (O_243,N_28551,N_29215);
nor UO_244 (O_244,N_27839,N_29301);
nor UO_245 (O_245,N_28459,N_27963);
and UO_246 (O_246,N_29702,N_28600);
nand UO_247 (O_247,N_27645,N_27366);
nand UO_248 (O_248,N_29189,N_29063);
or UO_249 (O_249,N_28745,N_27539);
xnor UO_250 (O_250,N_27722,N_29941);
xor UO_251 (O_251,N_27623,N_29249);
or UO_252 (O_252,N_27697,N_28239);
xor UO_253 (O_253,N_28545,N_27301);
xnor UO_254 (O_254,N_29456,N_28592);
nand UO_255 (O_255,N_29784,N_27255);
or UO_256 (O_256,N_27305,N_28022);
or UO_257 (O_257,N_27919,N_27055);
nand UO_258 (O_258,N_27777,N_29286);
or UO_259 (O_259,N_27165,N_29341);
xor UO_260 (O_260,N_27140,N_29093);
nor UO_261 (O_261,N_27624,N_28984);
nor UO_262 (O_262,N_27151,N_28382);
xor UO_263 (O_263,N_29476,N_27433);
nor UO_264 (O_264,N_29663,N_28417);
xnor UO_265 (O_265,N_29081,N_29568);
and UO_266 (O_266,N_29160,N_28819);
or UO_267 (O_267,N_29721,N_27916);
nand UO_268 (O_268,N_29262,N_29044);
xor UO_269 (O_269,N_28911,N_28456);
nor UO_270 (O_270,N_29151,N_27583);
nor UO_271 (O_271,N_29987,N_29666);
nand UO_272 (O_272,N_27764,N_28361);
nor UO_273 (O_273,N_27238,N_27115);
and UO_274 (O_274,N_27563,N_27298);
xor UO_275 (O_275,N_27258,N_28796);
and UO_276 (O_276,N_29766,N_27052);
nor UO_277 (O_277,N_27335,N_29765);
nand UO_278 (O_278,N_28324,N_27778);
nor UO_279 (O_279,N_28923,N_29155);
and UO_280 (O_280,N_28428,N_27211);
nor UO_281 (O_281,N_27877,N_27183);
xnor UO_282 (O_282,N_29352,N_27792);
and UO_283 (O_283,N_28681,N_29573);
nand UO_284 (O_284,N_28502,N_29003);
xor UO_285 (O_285,N_29952,N_28854);
nand UO_286 (O_286,N_27903,N_28983);
and UO_287 (O_287,N_27006,N_28161);
and UO_288 (O_288,N_27789,N_28610);
or UO_289 (O_289,N_29966,N_27447);
and UO_290 (O_290,N_28045,N_28937);
nor UO_291 (O_291,N_29696,N_29357);
nor UO_292 (O_292,N_27020,N_27307);
xnor UO_293 (O_293,N_28669,N_27262);
or UO_294 (O_294,N_28126,N_29457);
nand UO_295 (O_295,N_27487,N_27823);
and UO_296 (O_296,N_28224,N_28318);
or UO_297 (O_297,N_29681,N_27756);
nor UO_298 (O_298,N_28606,N_27462);
xor UO_299 (O_299,N_29660,N_27945);
or UO_300 (O_300,N_28287,N_28887);
xor UO_301 (O_301,N_27681,N_27377);
nor UO_302 (O_302,N_27074,N_28755);
nor UO_303 (O_303,N_27538,N_27879);
nor UO_304 (O_304,N_28761,N_29557);
xor UO_305 (O_305,N_29895,N_29128);
nor UO_306 (O_306,N_28131,N_29572);
and UO_307 (O_307,N_29452,N_27542);
and UO_308 (O_308,N_29488,N_29213);
xnor UO_309 (O_309,N_27971,N_29934);
and UO_310 (O_310,N_28476,N_28358);
xor UO_311 (O_311,N_28125,N_27315);
xor UO_312 (O_312,N_27742,N_28267);
and UO_313 (O_313,N_27125,N_27400);
nor UO_314 (O_314,N_27914,N_29074);
nand UO_315 (O_315,N_29173,N_28493);
nand UO_316 (O_316,N_29871,N_29578);
xnor UO_317 (O_317,N_28305,N_27465);
nor UO_318 (O_318,N_29367,N_27815);
and UO_319 (O_319,N_28857,N_29867);
nor UO_320 (O_320,N_27647,N_27444);
nor UO_321 (O_321,N_28317,N_28196);
nand UO_322 (O_322,N_28345,N_27120);
nand UO_323 (O_323,N_28415,N_27111);
or UO_324 (O_324,N_27237,N_29833);
xnor UO_325 (O_325,N_29657,N_27232);
nand UO_326 (O_326,N_29019,N_28310);
nor UO_327 (O_327,N_27330,N_29326);
nor UO_328 (O_328,N_28158,N_29661);
or UO_329 (O_329,N_27109,N_28809);
nor UO_330 (O_330,N_29026,N_29200);
xnor UO_331 (O_331,N_27748,N_27148);
or UO_332 (O_332,N_29558,N_28188);
nor UO_333 (O_333,N_27228,N_27933);
or UO_334 (O_334,N_28486,N_27144);
nor UO_335 (O_335,N_28244,N_29260);
nand UO_336 (O_336,N_27387,N_28171);
nand UO_337 (O_337,N_28366,N_29207);
xor UO_338 (O_338,N_27988,N_28750);
xnor UO_339 (O_339,N_29974,N_28391);
nor UO_340 (O_340,N_28364,N_27322);
xnor UO_341 (O_341,N_29604,N_27678);
nand UO_342 (O_342,N_29206,N_27475);
or UO_343 (O_343,N_29135,N_29653);
and UO_344 (O_344,N_28276,N_28206);
nand UO_345 (O_345,N_29519,N_28090);
nand UO_346 (O_346,N_27419,N_27692);
and UO_347 (O_347,N_27293,N_29690);
xor UO_348 (O_348,N_29265,N_28640);
xnor UO_349 (O_349,N_29398,N_28056);
nand UO_350 (O_350,N_27280,N_27331);
and UO_351 (O_351,N_28074,N_29704);
nand UO_352 (O_352,N_27886,N_29292);
or UO_353 (O_353,N_27089,N_28889);
and UO_354 (O_354,N_27123,N_29027);
xor UO_355 (O_355,N_28674,N_29920);
and UO_356 (O_356,N_27430,N_27429);
or UO_357 (O_357,N_28682,N_29203);
nand UO_358 (O_358,N_28990,N_27181);
xor UO_359 (O_359,N_27720,N_29569);
nor UO_360 (O_360,N_27701,N_27595);
or UO_361 (O_361,N_29039,N_27161);
nor UO_362 (O_362,N_28976,N_29248);
xnor UO_363 (O_363,N_29633,N_28609);
nor UO_364 (O_364,N_27832,N_27995);
nor UO_365 (O_365,N_29692,N_29049);
or UO_366 (O_366,N_29738,N_28075);
or UO_367 (O_367,N_27696,N_29954);
nand UO_368 (O_368,N_27811,N_27302);
or UO_369 (O_369,N_28526,N_29247);
nor UO_370 (O_370,N_27233,N_27658);
nor UO_371 (O_371,N_29923,N_28633);
nor UO_372 (O_372,N_27227,N_28715);
nor UO_373 (O_373,N_29860,N_28470);
xnor UO_374 (O_374,N_29553,N_29526);
and UO_375 (O_375,N_29985,N_28295);
and UO_376 (O_376,N_29437,N_28121);
xor UO_377 (O_377,N_29284,N_27025);
nand UO_378 (O_378,N_29984,N_29195);
and UO_379 (O_379,N_29217,N_28841);
and UO_380 (O_380,N_29433,N_27365);
nand UO_381 (O_381,N_28611,N_29791);
xnor UO_382 (O_382,N_28102,N_28438);
xnor UO_383 (O_383,N_27392,N_29268);
and UO_384 (O_384,N_27530,N_29459);
and UO_385 (O_385,N_28252,N_27397);
nand UO_386 (O_386,N_28445,N_28286);
or UO_387 (O_387,N_28563,N_28009);
nor UO_388 (O_388,N_28202,N_28076);
nand UO_389 (O_389,N_29302,N_28198);
nor UO_390 (O_390,N_27918,N_29716);
or UO_391 (O_391,N_29729,N_27359);
or UO_392 (O_392,N_29300,N_28615);
nor UO_393 (O_393,N_28095,N_28876);
nand UO_394 (O_394,N_29391,N_29319);
and UO_395 (O_395,N_28360,N_28639);
or UO_396 (O_396,N_28007,N_29539);
nand UO_397 (O_397,N_29855,N_29992);
or UO_398 (O_398,N_27058,N_28469);
xnor UO_399 (O_399,N_28578,N_28411);
or UO_400 (O_400,N_28550,N_28426);
and UO_401 (O_401,N_28328,N_29601);
nor UO_402 (O_402,N_28520,N_27281);
xor UO_403 (O_403,N_27027,N_28714);
xnor UO_404 (O_404,N_28173,N_28263);
xor UO_405 (O_405,N_29818,N_28498);
xor UO_406 (O_406,N_28241,N_28823);
nand UO_407 (O_407,N_28108,N_27834);
and UO_408 (O_408,N_29354,N_29192);
and UO_409 (O_409,N_29673,N_27501);
nor UO_410 (O_410,N_27866,N_28632);
xnor UO_411 (O_411,N_28182,N_27480);
nand UO_412 (O_412,N_28347,N_28711);
or UO_413 (O_413,N_28297,N_29658);
and UO_414 (O_414,N_29586,N_29718);
and UO_415 (O_415,N_29119,N_27984);
or UO_416 (O_416,N_27617,N_27320);
nor UO_417 (O_417,N_28416,N_28875);
nand UO_418 (O_418,N_29068,N_28970);
and UO_419 (O_419,N_27659,N_29862);
and UO_420 (O_420,N_28246,N_29126);
or UO_421 (O_421,N_29214,N_28720);
nand UO_422 (O_422,N_28993,N_28918);
xnor UO_423 (O_423,N_28060,N_29694);
and UO_424 (O_424,N_29123,N_27602);
or UO_425 (O_425,N_28620,N_29170);
or UO_426 (O_426,N_28392,N_27257);
and UO_427 (O_427,N_27005,N_28115);
nand UO_428 (O_428,N_29706,N_29793);
and UO_429 (O_429,N_29036,N_28320);
and UO_430 (O_430,N_27669,N_27106);
xor UO_431 (O_431,N_27030,N_29040);
nor UO_432 (O_432,N_27277,N_28868);
and UO_433 (O_433,N_29320,N_29401);
and UO_434 (O_434,N_29083,N_27096);
xor UO_435 (O_435,N_29304,N_27518);
nand UO_436 (O_436,N_28306,N_28292);
and UO_437 (O_437,N_28511,N_27978);
xnor UO_438 (O_438,N_28348,N_29735);
and UO_439 (O_439,N_27252,N_29907);
and UO_440 (O_440,N_28515,N_29651);
xor UO_441 (O_441,N_27004,N_28025);
and UO_442 (O_442,N_29989,N_27230);
xor UO_443 (O_443,N_29318,N_28078);
xor UO_444 (O_444,N_29630,N_28838);
and UO_445 (O_445,N_27186,N_27212);
and UO_446 (O_446,N_28830,N_27142);
xor UO_447 (O_447,N_29809,N_28023);
xor UO_448 (O_448,N_29535,N_27226);
xor UO_449 (O_449,N_29500,N_29618);
xnor UO_450 (O_450,N_29356,N_29487);
and UO_451 (O_451,N_28049,N_28934);
nor UO_452 (O_452,N_27256,N_28142);
or UO_453 (O_453,N_29258,N_27993);
nor UO_454 (O_454,N_29009,N_27234);
or UO_455 (O_455,N_28225,N_27615);
or UO_456 (O_456,N_27071,N_27388);
nand UO_457 (O_457,N_28953,N_29976);
nand UO_458 (O_458,N_29594,N_28582);
xnor UO_459 (O_459,N_27683,N_29016);
nand UO_460 (O_460,N_29199,N_28268);
nor UO_461 (O_461,N_27408,N_28892);
nor UO_462 (O_462,N_27482,N_27808);
and UO_463 (O_463,N_28152,N_27273);
and UO_464 (O_464,N_29808,N_29236);
nand UO_465 (O_465,N_27449,N_27163);
nor UO_466 (O_466,N_29520,N_28567);
or UO_467 (O_467,N_28458,N_29275);
nand UO_468 (O_468,N_28636,N_27665);
and UO_469 (O_469,N_28433,N_29225);
nor UO_470 (O_470,N_27841,N_28754);
nand UO_471 (O_471,N_29949,N_29418);
and UO_472 (O_472,N_28708,N_29211);
xor UO_473 (O_473,N_28407,N_28387);
xor UO_474 (O_474,N_29060,N_27849);
or UO_475 (O_475,N_29795,N_28568);
or UO_476 (O_476,N_29816,N_28523);
or UO_477 (O_477,N_27079,N_28003);
nand UO_478 (O_478,N_28723,N_28625);
nor UO_479 (O_479,N_27568,N_27316);
nand UO_480 (O_480,N_28690,N_27452);
nand UO_481 (O_481,N_29968,N_29548);
or UO_482 (O_482,N_29386,N_29655);
nor UO_483 (O_483,N_29722,N_28904);
nor UO_484 (O_484,N_28051,N_29066);
nand UO_485 (O_485,N_27067,N_28678);
and UO_486 (O_486,N_27502,N_29811);
nor UO_487 (O_487,N_29824,N_27575);
and UO_488 (O_488,N_28933,N_28654);
and UO_489 (O_489,N_28879,N_29480);
and UO_490 (O_490,N_27625,N_28208);
and UO_491 (O_491,N_27146,N_28427);
xor UO_492 (O_492,N_29468,N_28733);
xnor UO_493 (O_493,N_29012,N_27461);
nor UO_494 (O_494,N_28140,N_27072);
nor UO_495 (O_495,N_27150,N_29010);
or UO_496 (O_496,N_27987,N_27770);
xor UO_497 (O_497,N_27867,N_28150);
nor UO_498 (O_498,N_27064,N_28914);
xnor UO_499 (O_499,N_27490,N_29518);
nor UO_500 (O_500,N_27208,N_28912);
and UO_501 (O_501,N_29004,N_29684);
nand UO_502 (O_502,N_28719,N_28510);
and UO_503 (O_503,N_29579,N_28155);
or UO_504 (O_504,N_27370,N_28109);
and UO_505 (O_505,N_27489,N_29112);
and UO_506 (O_506,N_28000,N_27664);
xor UO_507 (O_507,N_27294,N_29346);
nand UO_508 (O_508,N_29303,N_28026);
xnor UO_509 (O_509,N_29430,N_28052);
or UO_510 (O_510,N_27941,N_29957);
and UO_511 (O_511,N_28163,N_28638);
or UO_512 (O_512,N_28389,N_29371);
nand UO_513 (O_513,N_27344,N_28650);
nor UO_514 (O_514,N_29537,N_29647);
xnor UO_515 (O_515,N_29592,N_28210);
nand UO_516 (O_516,N_29469,N_29550);
nand UO_517 (O_517,N_28978,N_27050);
or UO_518 (O_518,N_29744,N_29202);
nor UO_519 (O_519,N_28005,N_27725);
xor UO_520 (O_520,N_27382,N_29754);
xnor UO_521 (O_521,N_29282,N_27822);
and UO_522 (O_522,N_28701,N_28813);
nor UO_523 (O_523,N_28490,N_28749);
or UO_524 (O_524,N_27189,N_27734);
and UO_525 (O_525,N_27413,N_29406);
and UO_526 (O_526,N_28500,N_29880);
xnor UO_527 (O_527,N_27373,N_29394);
and UO_528 (O_528,N_28790,N_28375);
nor UO_529 (O_529,N_27890,N_28116);
or UO_530 (O_530,N_29814,N_27548);
xnor UO_531 (O_531,N_29090,N_27900);
and UO_532 (O_532,N_27217,N_28169);
nand UO_533 (O_533,N_27888,N_28645);
nor UO_534 (O_534,N_29201,N_29316);
xor UO_535 (O_535,N_27070,N_28186);
nand UO_536 (O_536,N_29581,N_28635);
and UO_537 (O_537,N_27367,N_29237);
and UO_538 (O_538,N_29259,N_27648);
nor UO_539 (O_539,N_29423,N_27924);
nand UO_540 (O_540,N_27767,N_29067);
and UO_541 (O_541,N_27479,N_28017);
or UO_542 (O_542,N_28542,N_28437);
xor UO_543 (O_543,N_28372,N_28979);
xor UO_544 (O_544,N_28688,N_28756);
xor UO_545 (O_545,N_29245,N_28553);
or UO_546 (O_546,N_27620,N_29625);
and UO_547 (O_547,N_29428,N_28577);
and UO_548 (O_548,N_28291,N_29707);
and UO_549 (O_549,N_29713,N_28495);
nor UO_550 (O_550,N_28399,N_28776);
or UO_551 (O_551,N_27536,N_29100);
xnor UO_552 (O_552,N_29020,N_28177);
and UO_553 (O_553,N_29820,N_28546);
nand UO_554 (O_554,N_29138,N_29847);
nor UO_555 (O_555,N_27966,N_27426);
nor UO_556 (O_556,N_28893,N_29184);
and UO_557 (O_557,N_28218,N_29832);
nand UO_558 (O_558,N_27225,N_27383);
xor UO_559 (O_559,N_27952,N_28068);
and UO_560 (O_560,N_28940,N_29489);
xnor UO_561 (O_561,N_27884,N_28722);
and UO_562 (O_562,N_28528,N_28153);
nand UO_563 (O_563,N_27603,N_27759);
xnor UO_564 (O_564,N_27550,N_29714);
nor UO_565 (O_565,N_28965,N_27577);
xor UO_566 (O_566,N_28353,N_28770);
nand UO_567 (O_567,N_27156,N_29925);
and UO_568 (O_568,N_27622,N_29971);
nand UO_569 (O_569,N_28961,N_27045);
or UO_570 (O_570,N_27406,N_27137);
nand UO_571 (O_571,N_29099,N_27110);
nor UO_572 (O_572,N_27975,N_29393);
nand UO_573 (O_573,N_27464,N_29963);
nor UO_574 (O_574,N_28800,N_28455);
xnor UO_575 (O_575,N_27882,N_27099);
xor UO_576 (O_576,N_28789,N_29853);
or UO_577 (O_577,N_28539,N_28576);
xor UO_578 (O_578,N_29844,N_27875);
nor UO_579 (O_579,N_28402,N_29382);
and UO_580 (O_580,N_28847,N_28084);
or UO_581 (O_581,N_29649,N_29903);
and UO_582 (O_582,N_29297,N_28325);
xnor UO_583 (O_583,N_27844,N_27980);
and UO_584 (O_584,N_28132,N_27193);
xnor UO_585 (O_585,N_27044,N_27241);
or UO_586 (O_586,N_29276,N_27276);
nor UO_587 (O_587,N_28033,N_27040);
and UO_588 (O_588,N_27154,N_29314);
nand UO_589 (O_589,N_29404,N_29763);
nor UO_590 (O_590,N_27629,N_27076);
and UO_591 (O_591,N_29047,N_28053);
or UO_592 (O_592,N_28335,N_29130);
and UO_593 (O_593,N_27646,N_27733);
nand UO_594 (O_594,N_28002,N_28590);
and UO_595 (O_595,N_29461,N_29600);
and UO_596 (O_596,N_27338,N_27512);
xor UO_597 (O_597,N_27891,N_27587);
nand UO_598 (O_598,N_28771,N_29454);
or UO_599 (O_599,N_28762,N_27391);
or UO_600 (O_600,N_29444,N_29451);
nand UO_601 (O_601,N_27719,N_28718);
nor UO_602 (O_602,N_29342,N_29311);
nor UO_603 (O_603,N_27737,N_28525);
nor UO_604 (O_604,N_29910,N_29632);
and UO_605 (O_605,N_29620,N_27905);
nand UO_606 (O_606,N_28439,N_27345);
nand UO_607 (O_607,N_27455,N_27599);
and UO_608 (O_608,N_29891,N_27728);
nor UO_609 (O_609,N_29376,N_29261);
nand UO_610 (O_610,N_29801,N_28031);
and UO_611 (O_611,N_27474,N_29108);
xor UO_612 (O_612,N_28533,N_28985);
or UO_613 (O_613,N_27970,N_29552);
nor UO_614 (O_614,N_28418,N_29521);
and UO_615 (O_615,N_28062,N_28379);
or UO_616 (O_616,N_29612,N_29533);
xor UO_617 (O_617,N_28913,N_29505);
or UO_618 (O_618,N_27732,N_27343);
and UO_619 (O_619,N_27242,N_29611);
nor UO_620 (O_620,N_29736,N_29946);
nor UO_621 (O_621,N_27470,N_27567);
and UO_622 (O_622,N_29589,N_28547);
nand UO_623 (O_623,N_27885,N_27083);
nor UO_624 (O_624,N_28044,N_28580);
and UO_625 (O_625,N_29980,N_29737);
xor UO_626 (O_626,N_28518,N_29442);
nor UO_627 (O_627,N_27899,N_28390);
nor UO_628 (O_628,N_27494,N_28702);
or UO_629 (O_629,N_27515,N_28741);
and UO_630 (O_630,N_28627,N_28117);
nand UO_631 (O_631,N_29624,N_27152);
xnor UO_632 (O_632,N_28315,N_28662);
and UO_633 (O_633,N_29256,N_28370);
nand UO_634 (O_634,N_28624,N_27626);
nand UO_635 (O_635,N_29299,N_28534);
xnor UO_636 (O_636,N_28256,N_29014);
xor UO_637 (O_637,N_27921,N_27731);
xnor UO_638 (O_638,N_27191,N_27102);
xnor UO_639 (O_639,N_27299,N_27655);
nor UO_640 (O_640,N_28753,N_29644);
xor UO_641 (O_641,N_29839,N_29845);
or UO_642 (O_642,N_29415,N_27747);
nand UO_643 (O_643,N_27698,N_29175);
xnor UO_644 (O_644,N_27569,N_27454);
and UO_645 (O_645,N_28907,N_28670);
and UO_646 (O_646,N_27723,N_27738);
nor UO_647 (O_647,N_28189,N_29623);
or UO_648 (O_648,N_29495,N_28660);
or UO_649 (O_649,N_27159,N_27752);
nor UO_650 (O_650,N_28903,N_27222);
and UO_651 (O_651,N_29077,N_28552);
xnor UO_652 (O_652,N_29648,N_27360);
nand UO_653 (O_653,N_28374,N_29975);
and UO_654 (O_654,N_29870,N_29857);
or UO_655 (O_655,N_28958,N_27976);
and UO_656 (O_656,N_28710,N_29850);
xor UO_657 (O_657,N_27540,N_28376);
and UO_658 (O_658,N_28508,N_27585);
or UO_659 (O_659,N_28855,N_29727);
xnor UO_660 (O_660,N_28199,N_28247);
and UO_661 (O_661,N_29582,N_27843);
and UO_662 (O_662,N_27473,N_29379);
and UO_663 (O_663,N_27017,N_28113);
xor UO_664 (O_664,N_27235,N_27428);
nor UO_665 (O_665,N_28807,N_27532);
or UO_666 (O_666,N_28888,N_27847);
nand UO_667 (O_667,N_28180,N_29257);
nand UO_668 (O_668,N_29043,N_28676);
and UO_669 (O_669,N_28947,N_28964);
and UO_670 (O_670,N_28814,N_29054);
or UO_671 (O_671,N_29445,N_28420);
or UO_672 (O_672,N_28833,N_29460);
nand UO_673 (O_673,N_29246,N_29492);
nand UO_674 (O_674,N_27103,N_28898);
or UO_675 (O_675,N_28135,N_29499);
and UO_676 (O_676,N_29037,N_27848);
and UO_677 (O_677,N_27956,N_28006);
and UO_678 (O_678,N_27363,N_28969);
xnor UO_679 (O_679,N_28414,N_27951);
nor UO_680 (O_680,N_28229,N_28093);
and UO_681 (O_681,N_27104,N_28516);
nand UO_682 (O_682,N_29755,N_29105);
and UO_683 (O_683,N_29405,N_27357);
xnor UO_684 (O_684,N_29631,N_29205);
nand UO_685 (O_685,N_29242,N_29429);
nand UO_686 (O_686,N_27950,N_29193);
and UO_687 (O_687,N_29477,N_28760);
nand UO_688 (O_688,N_27817,N_27249);
xnor UO_689 (O_689,N_27959,N_29231);
nand UO_690 (O_690,N_27312,N_27488);
nand UO_691 (O_691,N_27990,N_27907);
xor UO_692 (O_692,N_29551,N_29541);
xor UO_693 (O_693,N_27442,N_28865);
nor UO_694 (O_694,N_27755,N_29576);
nor UO_695 (O_695,N_27018,N_28187);
or UO_696 (O_696,N_28901,N_29191);
or UO_697 (O_697,N_29334,N_29774);
nor UO_698 (O_698,N_28344,N_29777);
or UO_699 (O_699,N_28449,N_29064);
nor UO_700 (O_700,N_29024,N_28137);
nand UO_701 (O_701,N_29313,N_28924);
nand UO_702 (O_702,N_27171,N_27218);
or UO_703 (O_703,N_27593,N_27851);
nor UO_704 (O_704,N_28945,N_28536);
nand UO_705 (O_705,N_27578,N_29486);
and UO_706 (O_706,N_27680,N_28629);
nand UO_707 (O_707,N_28858,N_28269);
nor UO_708 (O_708,N_29216,N_28018);
xnor UO_709 (O_709,N_28782,N_28928);
and UO_710 (O_710,N_28531,N_29899);
nand UO_711 (O_711,N_29608,N_28692);
xor UO_712 (O_712,N_28046,N_28950);
or UO_713 (O_713,N_27935,N_27576);
nand UO_714 (O_714,N_27476,N_29745);
or UO_715 (O_715,N_28087,N_27195);
or UO_716 (O_716,N_27060,N_29096);
nand UO_717 (O_717,N_29530,N_29575);
or UO_718 (O_718,N_27564,N_27441);
nand UO_719 (O_719,N_27898,N_28440);
and UO_720 (O_720,N_29669,N_28837);
nor UO_721 (O_721,N_28064,N_27396);
nor UO_722 (O_722,N_29337,N_28434);
nand UO_723 (O_723,N_27726,N_27836);
or UO_724 (O_724,N_27327,N_29679);
nand UO_725 (O_725,N_27453,N_28726);
or UO_726 (O_726,N_27917,N_29515);
nand UO_727 (O_727,N_28675,N_29938);
or UO_728 (O_728,N_28998,N_29264);
nand UO_729 (O_729,N_27735,N_27619);
nor UO_730 (O_730,N_29159,N_28079);
and UO_731 (O_731,N_27167,N_29157);
xnor UO_732 (O_732,N_29788,N_27418);
and UO_733 (O_733,N_27529,N_27762);
nand UO_734 (O_734,N_28197,N_27466);
nand UO_735 (O_735,N_29502,N_28430);
or UO_736 (O_736,N_27565,N_27998);
nor UO_737 (O_737,N_28260,N_27329);
xor UO_738 (O_738,N_28474,N_29496);
nand UO_739 (O_739,N_28200,N_29483);
nor UO_740 (O_740,N_27706,N_27088);
and UO_741 (O_741,N_27895,N_27221);
xnor UO_742 (O_742,N_27264,N_28505);
nand UO_743 (O_743,N_28191,N_28544);
nor UO_744 (O_744,N_27668,N_27636);
or UO_745 (O_745,N_28856,N_27807);
nand UO_746 (O_746,N_29094,N_27700);
nor UO_747 (O_747,N_27034,N_29463);
xor UO_748 (O_748,N_29332,N_28145);
or UO_749 (O_749,N_29628,N_29865);
or UO_750 (O_750,N_28878,N_29761);
nand UO_751 (O_751,N_28974,N_28565);
or UO_752 (O_752,N_29462,N_28739);
xnor UO_753 (O_753,N_29355,N_27073);
and UO_754 (O_754,N_28067,N_27685);
or UO_755 (O_755,N_28442,N_27551);
nor UO_756 (O_756,N_27023,N_28479);
nor UO_757 (O_757,N_29599,N_29210);
and UO_758 (O_758,N_29559,N_28309);
xnor UO_759 (O_759,N_28812,N_28827);
xnor UO_760 (O_760,N_27977,N_27399);
xnor UO_761 (O_761,N_28094,N_29705);
nor UO_762 (O_762,N_27393,N_28691);
and UO_763 (O_763,N_27704,N_29221);
nor UO_764 (O_764,N_29503,N_28955);
or UO_765 (O_765,N_28925,N_27084);
and UO_766 (O_766,N_27744,N_29671);
nor UO_767 (O_767,N_27483,N_28932);
and UO_768 (O_768,N_27164,N_29161);
xnor UO_769 (O_769,N_28397,N_27982);
nand UO_770 (O_770,N_28897,N_28758);
nand UO_771 (O_771,N_29273,N_29603);
nor UO_772 (O_772,N_28860,N_29642);
nor UO_773 (O_773,N_29711,N_28507);
nand UO_774 (O_774,N_27835,N_29686);
nor UO_775 (O_775,N_27544,N_28778);
nand UO_776 (O_776,N_28329,N_29918);
nor UO_777 (O_777,N_27714,N_27524);
xnor UO_778 (O_778,N_27122,N_27061);
xor UO_779 (O_779,N_27781,N_28422);
xor UO_780 (O_780,N_29345,N_27326);
and UO_781 (O_781,N_27378,N_29144);
xnor UO_782 (O_782,N_27724,N_27663);
or UO_783 (O_783,N_29691,N_27204);
or UO_784 (O_784,N_27831,N_27657);
nand UO_785 (O_785,N_29849,N_27101);
nand UO_786 (O_786,N_27631,N_28825);
and UO_787 (O_787,N_27511,N_28070);
nor UO_788 (O_788,N_28765,N_29015);
and UO_789 (O_789,N_28302,N_27342);
nor UO_790 (O_790,N_29413,N_28713);
or UO_791 (O_791,N_29831,N_28054);
nor UO_792 (O_792,N_27986,N_27003);
nor UO_793 (O_793,N_28902,N_28396);
and UO_794 (O_794,N_29909,N_28363);
xor UO_795 (O_795,N_29396,N_29693);
nor UO_796 (O_796,N_29435,N_27434);
nand UO_797 (O_797,N_28296,N_27821);
nand UO_798 (O_798,N_29646,N_27944);
nand UO_799 (O_799,N_29543,N_29424);
nor UO_800 (O_800,N_29104,N_28941);
and UO_801 (O_801,N_29080,N_27376);
nor UO_802 (O_802,N_29848,N_27033);
xnor UO_803 (O_803,N_29955,N_28111);
xnor UO_804 (O_804,N_29125,N_28285);
and UO_805 (O_805,N_28350,N_28195);
xnor UO_806 (O_806,N_27946,N_28631);
nor UO_807 (O_807,N_27590,N_28698);
nor UO_808 (O_808,N_27594,N_27100);
xor UO_809 (O_809,N_27244,N_27323);
and UO_810 (O_810,N_27194,N_29680);
nor UO_811 (O_811,N_29780,N_29188);
and UO_812 (O_812,N_29484,N_29861);
xor UO_813 (O_813,N_28641,N_29018);
xor UO_814 (O_814,N_27800,N_29285);
nand UO_815 (O_815,N_27661,N_27484);
or UO_816 (O_816,N_27416,N_27379);
xor UO_817 (O_817,N_27369,N_28249);
and UO_818 (O_818,N_29607,N_29353);
and UO_819 (O_819,N_27112,N_27640);
nand UO_820 (O_820,N_28621,N_28846);
xnor UO_821 (O_821,N_29858,N_28340);
or UO_822 (O_822,N_27436,N_27380);
nor UO_823 (O_823,N_28651,N_29250);
nand UO_824 (O_824,N_29038,N_29471);
nor UO_825 (O_825,N_28409,N_27618);
nand UO_826 (O_826,N_28277,N_27037);
and UO_827 (O_827,N_29981,N_28944);
nor UO_828 (O_828,N_27361,N_28828);
xor UO_829 (O_829,N_27958,N_28622);
nand UO_830 (O_830,N_28740,N_29821);
or UO_831 (O_831,N_28687,N_29783);
nand UO_832 (O_832,N_29757,N_28589);
nand UO_833 (O_833,N_27897,N_27533);
or UO_834 (O_834,N_29029,N_29724);
nor UO_835 (O_835,N_27523,N_29501);
nor UO_836 (O_836,N_29750,N_27960);
xnor UO_837 (O_837,N_27458,N_29061);
and UO_838 (O_838,N_29872,N_27743);
and UO_839 (O_839,N_29017,N_28175);
or UO_840 (O_840,N_27927,N_27266);
nand UO_841 (O_841,N_27964,N_29921);
and UO_842 (O_842,N_28106,N_27503);
nor UO_843 (O_843,N_27763,N_29089);
xor UO_844 (O_844,N_27782,N_27902);
nand UO_845 (O_845,N_28880,N_27202);
xor UO_846 (O_846,N_28480,N_28048);
or UO_847 (O_847,N_29698,N_28792);
or UO_848 (O_848,N_27992,N_28916);
and UO_849 (O_849,N_29819,N_28047);
and UO_850 (O_850,N_28596,N_28149);
and UO_851 (O_851,N_28089,N_28118);
or UO_852 (O_852,N_28549,N_28136);
nand UO_853 (O_853,N_27873,N_29940);
nand UO_854 (O_854,N_27260,N_28450);
nor UO_855 (O_855,N_28591,N_29924);
xnor UO_856 (O_856,N_27850,N_29190);
xnor UO_857 (O_857,N_29509,N_28491);
nand UO_858 (O_858,N_29127,N_29516);
nor UO_859 (O_859,N_27901,N_28899);
nand UO_860 (O_860,N_27095,N_28042);
xnor UO_861 (O_861,N_29799,N_29001);
or UO_862 (O_862,N_28929,N_28243);
nor UO_863 (O_863,N_28029,N_27053);
or UO_864 (O_864,N_29562,N_28881);
and UO_865 (O_865,N_29293,N_27633);
nor UO_866 (O_866,N_27967,N_29134);
xor UO_867 (O_867,N_27947,N_27616);
xor UO_868 (O_868,N_27351,N_27440);
nand UO_869 (O_869,N_27401,N_28579);
nor UO_870 (O_870,N_28088,N_29829);
nor UO_871 (O_871,N_27634,N_28694);
nor UO_872 (O_872,N_27974,N_29841);
xor UO_873 (O_873,N_29389,N_29087);
nand UO_874 (O_874,N_28174,N_28734);
xor UO_875 (O_875,N_28160,N_27080);
or UO_876 (O_876,N_29069,N_28801);
or UO_877 (O_877,N_28982,N_28601);
or UO_878 (O_878,N_28786,N_27773);
nor UO_879 (O_879,N_28219,N_27820);
xor UO_880 (O_880,N_29885,N_28824);
nand UO_881 (O_881,N_28791,N_28779);
and UO_882 (O_882,N_28835,N_27871);
nor UO_883 (O_883,N_27691,N_29229);
or UO_884 (O_884,N_29930,N_28463);
or UO_885 (O_885,N_28628,N_29443);
or UO_886 (O_886,N_27932,N_29743);
and UO_887 (O_887,N_29290,N_27179);
or UO_888 (O_888,N_28648,N_28242);
or UO_889 (O_889,N_29223,N_27209);
or UO_890 (O_890,N_27922,N_28891);
nand UO_891 (O_891,N_28535,N_28264);
xnor UO_892 (O_892,N_27838,N_28395);
and UO_893 (O_893,N_27522,N_29627);
nor UO_894 (O_894,N_29212,N_29914);
xor UO_895 (O_895,N_29523,N_28815);
nand UO_896 (O_896,N_29166,N_28724);
xnor UO_897 (O_897,N_27145,N_29278);
nand UO_898 (O_898,N_28316,N_29402);
or UO_899 (O_899,N_28871,N_28727);
nor UO_900 (O_900,N_27627,N_28331);
nor UO_901 (O_901,N_28775,N_29760);
or UO_902 (O_902,N_29375,N_28866);
nor UO_903 (O_903,N_27931,N_29659);
and UO_904 (O_904,N_29165,N_29238);
and UO_905 (O_905,N_29846,N_28351);
xor UO_906 (O_906,N_27300,N_28997);
or UO_907 (O_907,N_28781,N_28144);
xor UO_908 (O_908,N_27019,N_28989);
xor UO_909 (O_909,N_28962,N_28840);
or UO_910 (O_910,N_29639,N_28513);
xor UO_911 (O_911,N_28748,N_27749);
nand UO_912 (O_912,N_28103,N_29360);
nor UO_913 (O_913,N_27468,N_28811);
and UO_914 (O_914,N_29922,N_27541);
nand UO_915 (O_915,N_28419,N_27214);
or UO_916 (O_916,N_27162,N_27601);
and UO_917 (O_917,N_27591,N_28119);
and UO_918 (O_918,N_28464,N_29439);
xnor UO_919 (O_919,N_27309,N_27002);
xor UO_920 (O_920,N_29136,N_29281);
xnor UO_921 (O_921,N_29307,N_29441);
or UO_922 (O_922,N_27589,N_27710);
or UO_923 (O_923,N_29703,N_28919);
and UO_924 (O_924,N_29084,N_28308);
nand UO_925 (O_925,N_27892,N_27271);
nor UO_926 (O_926,N_27333,N_28058);
or UO_927 (O_927,N_29349,N_29997);
xnor UO_928 (O_928,N_27635,N_28300);
and UO_929 (O_929,N_27868,N_28314);
xnor UO_930 (O_930,N_27553,N_28334);
and UO_931 (O_931,N_28798,N_27957);
xnor UO_932 (O_932,N_28884,N_27153);
or UO_933 (O_933,N_29007,N_29467);
xnor UO_934 (O_934,N_28035,N_29508);
nor UO_935 (O_935,N_28170,N_29244);
xor UO_936 (O_936,N_29146,N_29717);
xnor UO_937 (O_937,N_29699,N_29616);
or UO_938 (O_938,N_29580,N_29719);
or UO_939 (O_939,N_29677,N_29593);
nor UO_940 (O_940,N_27906,N_27160);
nand UO_941 (O_941,N_27013,N_28787);
and UO_942 (O_942,N_28475,N_28154);
nor UO_943 (O_943,N_29186,N_27790);
nand UO_944 (O_944,N_29395,N_27086);
nand UO_945 (O_945,N_27356,N_28667);
xnor UO_946 (O_946,N_29605,N_29410);
xor UO_947 (O_947,N_29321,N_27675);
or UO_948 (O_948,N_27705,N_29881);
xnor UO_949 (O_949,N_27190,N_27686);
nor UO_950 (O_950,N_27842,N_27934);
and UO_951 (O_951,N_29710,N_27421);
and UO_952 (O_952,N_28388,N_28354);
or UO_953 (O_953,N_27261,N_29121);
or UO_954 (O_954,N_27289,N_28057);
nor UO_955 (O_955,N_29904,N_28016);
or UO_956 (O_956,N_29139,N_27750);
nand UO_957 (O_957,N_28529,N_29759);
nand UO_958 (O_958,N_29953,N_29772);
or UO_959 (O_959,N_29228,N_27321);
xor UO_960 (O_960,N_29685,N_28460);
and UO_961 (O_961,N_28110,N_29013);
and UO_962 (O_962,N_27894,N_29085);
and UO_963 (O_963,N_27702,N_28991);
or UO_964 (O_964,N_29182,N_29874);
nor UO_965 (O_965,N_27139,N_27509);
nand UO_966 (O_966,N_29978,N_27295);
nor UO_967 (O_967,N_29141,N_27010);
nor UO_968 (O_968,N_28139,N_27346);
nand UO_969 (O_969,N_27819,N_29837);
nor UO_970 (O_970,N_28367,N_28643);
nor UO_971 (O_971,N_27588,N_29892);
nor UO_972 (O_972,N_28613,N_29597);
xnor UO_973 (O_973,N_27943,N_29381);
or UO_974 (O_974,N_27508,N_27097);
xor UO_975 (O_975,N_27546,N_29931);
xor UO_976 (O_976,N_27049,N_29158);
xor UO_977 (O_977,N_27059,N_27056);
or UO_978 (O_978,N_28839,N_29412);
and UO_979 (O_979,N_28587,N_29970);
or UO_980 (O_980,N_29838,N_28634);
and UO_981 (O_981,N_28584,N_29181);
and UO_982 (O_982,N_29294,N_29951);
and UO_983 (O_983,N_28738,N_28383);
nor UO_984 (O_984,N_27662,N_27201);
nor UO_985 (O_985,N_27358,N_27063);
xnor UO_986 (O_986,N_28872,N_29031);
and UO_987 (O_987,N_29366,N_28693);
xor UO_988 (O_988,N_27558,N_29374);
xor UO_989 (O_989,N_28063,N_27039);
nor UO_990 (O_990,N_27911,N_27306);
xor UO_991 (O_991,N_27029,N_27673);
nor UO_992 (O_992,N_28461,N_29185);
or UO_993 (O_993,N_28129,N_29540);
and UO_994 (O_994,N_28747,N_27928);
or UO_995 (O_995,N_28214,N_28393);
nand UO_996 (O_996,N_29079,N_28571);
nand UO_997 (O_997,N_27038,N_28081);
nor UO_998 (O_998,N_27486,N_29178);
or UO_999 (O_999,N_27087,N_27793);
nand UO_1000 (O_1000,N_29274,N_29768);
nand UO_1001 (O_1001,N_29271,N_28034);
xor UO_1002 (O_1002,N_27715,N_28886);
xnor UO_1003 (O_1003,N_29547,N_27169);
or UO_1004 (O_1004,N_29851,N_27912);
nand UO_1005 (O_1005,N_29196,N_29449);
nand UO_1006 (O_1006,N_28554,N_28522);
xor UO_1007 (O_1007,N_29812,N_29071);
nor UO_1008 (O_1008,N_29378,N_27613);
xor UO_1009 (O_1009,N_28290,N_27981);
xor UO_1010 (O_1010,N_28408,N_29876);
nand UO_1011 (O_1011,N_27207,N_27386);
nor UO_1012 (O_1012,N_27098,N_29927);
xnor UO_1013 (O_1013,N_27818,N_27032);
and UO_1014 (O_1014,N_28128,N_28729);
nand UO_1015 (O_1015,N_29566,N_28597);
nor UO_1016 (O_1016,N_28561,N_29674);
nand UO_1017 (O_1017,N_27290,N_28072);
nand UO_1018 (O_1018,N_28960,N_27521);
xor UO_1019 (O_1019,N_29383,N_27296);
nor UO_1020 (O_1020,N_28404,N_29688);
nor UO_1021 (O_1021,N_28503,N_28496);
nand UO_1022 (O_1022,N_27827,N_29328);
nand UO_1023 (O_1023,N_29544,N_29154);
and UO_1024 (O_1024,N_28604,N_27325);
xnor UO_1025 (O_1025,N_28683,N_29033);
or UO_1026 (O_1026,N_29172,N_29095);
or UO_1027 (O_1027,N_27128,N_27825);
xor UO_1028 (O_1028,N_27688,N_28013);
nand UO_1029 (O_1029,N_29528,N_27176);
nor UO_1030 (O_1030,N_27199,N_29131);
nand UO_1031 (O_1031,N_29338,N_28684);
nand UO_1032 (O_1032,N_28238,N_28564);
nand UO_1033 (O_1033,N_29749,N_28672);
nor UO_1034 (O_1034,N_27582,N_27292);
and UO_1035 (O_1035,N_27962,N_29239);
xnor UO_1036 (O_1036,N_29251,N_29879);
xnor UO_1037 (O_1037,N_29715,N_28649);
nand UO_1038 (O_1038,N_27353,N_29742);
nor UO_1039 (O_1039,N_28930,N_27812);
and UO_1040 (O_1040,N_27671,N_27185);
and UO_1041 (O_1041,N_28284,N_28323);
xor UO_1042 (O_1042,N_29823,N_28271);
nor UO_1043 (O_1043,N_27467,N_27035);
xnor UO_1044 (O_1044,N_28281,N_28228);
and UO_1045 (O_1045,N_28548,N_27324);
and UO_1046 (O_1046,N_28737,N_28700);
nor UO_1047 (O_1047,N_28501,N_27991);
nand UO_1048 (O_1048,N_29995,N_29408);
xor UO_1049 (O_1049,N_27826,N_29306);
or UO_1050 (O_1050,N_28304,N_28644);
nor UO_1051 (O_1051,N_28996,N_27188);
or UO_1052 (O_1052,N_28435,N_29800);
xor UO_1053 (O_1053,N_28203,N_27572);
or UO_1054 (O_1054,N_29522,N_29309);
xnor UO_1055 (O_1055,N_29884,N_29863);
nor UO_1056 (O_1056,N_29629,N_27443);
nand UO_1057 (O_1057,N_28607,N_29390);
or UO_1058 (O_1058,N_28259,N_29555);
nor UO_1059 (O_1059,N_29708,N_29962);
nor UO_1060 (O_1060,N_28234,N_28036);
and UO_1061 (O_1061,N_28910,N_29873);
and UO_1062 (O_1062,N_27341,N_27703);
xor UO_1063 (O_1063,N_27994,N_27766);
nor UO_1064 (O_1064,N_27846,N_29779);
and UO_1065 (O_1065,N_27200,N_27471);
xnor UO_1066 (O_1066,N_28293,N_29327);
or UO_1067 (O_1067,N_29911,N_29893);
and UO_1068 (O_1068,N_27205,N_28506);
and UO_1069 (O_1069,N_29944,N_27674);
or UO_1070 (O_1070,N_28519,N_29935);
or UO_1071 (O_1071,N_27783,N_29373);
and UO_1072 (O_1072,N_29532,N_29474);
or UO_1073 (O_1073,N_28099,N_28939);
nand UO_1074 (O_1074,N_27126,N_27042);
or UO_1075 (O_1075,N_28352,N_28332);
nor UO_1076 (O_1076,N_27133,N_27791);
or UO_1077 (O_1077,N_28098,N_27424);
nand UO_1078 (O_1078,N_29400,N_28834);
and UO_1079 (O_1079,N_27445,N_29959);
or UO_1080 (O_1080,N_28949,N_27794);
xnor UO_1081 (O_1081,N_29834,N_28319);
xnor UO_1082 (O_1082,N_29513,N_28138);
xnor UO_1083 (O_1083,N_27554,N_27670);
nor UO_1084 (O_1084,N_27328,N_27896);
nand UO_1085 (O_1085,N_29021,N_28573);
xnor UO_1086 (O_1086,N_28569,N_29312);
nand UO_1087 (O_1087,N_28706,N_27727);
or UO_1088 (O_1088,N_29712,N_27270);
xor UO_1089 (O_1089,N_27758,N_27334);
nor UO_1090 (O_1090,N_27573,N_28330);
or UO_1091 (O_1091,N_27395,N_27608);
nor UO_1092 (O_1092,N_29982,N_29802);
xor UO_1093 (O_1093,N_28504,N_27229);
xor UO_1094 (O_1094,N_28021,N_28467);
and UO_1095 (O_1095,N_28133,N_29380);
or UO_1096 (O_1096,N_28004,N_28652);
xor UO_1097 (O_1097,N_27402,N_28368);
nand UO_1098 (O_1098,N_29143,N_27078);
or UO_1099 (O_1099,N_27862,N_27236);
and UO_1100 (O_1100,N_27730,N_28356);
nand UO_1101 (O_1101,N_29613,N_29385);
xnor UO_1102 (O_1102,N_29052,N_28658);
nor UO_1103 (O_1103,N_28217,N_29939);
nor UO_1104 (O_1104,N_28223,N_29746);
nand UO_1105 (O_1105,N_27114,N_29596);
and UO_1106 (O_1106,N_29168,N_28178);
and UO_1107 (O_1107,N_28712,N_27741);
xor UO_1108 (O_1108,N_27354,N_27637);
and UO_1109 (O_1109,N_27788,N_29325);
and UO_1110 (O_1110,N_29224,N_29287);
or UO_1111 (O_1111,N_29148,N_27389);
nand UO_1112 (O_1112,N_27407,N_27876);
nand UO_1113 (O_1113,N_28566,N_27174);
and UO_1114 (O_1114,N_27566,N_27091);
nand UO_1115 (O_1115,N_28337,N_29534);
xnor UO_1116 (O_1116,N_27062,N_29636);
xor UO_1117 (O_1117,N_28377,N_29504);
nand UO_1118 (O_1118,N_29902,N_29868);
or UO_1119 (O_1119,N_28485,N_27166);
nor UO_1120 (O_1120,N_29972,N_27248);
or UO_1121 (O_1121,N_28313,N_29315);
nor UO_1122 (O_1122,N_28558,N_28832);
xor UO_1123 (O_1123,N_29220,N_28730);
or UO_1124 (O_1124,N_29323,N_28336);
nor UO_1125 (O_1125,N_28605,N_27285);
xnor UO_1126 (O_1126,N_28159,N_29906);
or UO_1127 (O_1127,N_27008,N_27007);
xor UO_1128 (O_1128,N_27041,N_27543);
xor UO_1129 (O_1129,N_29776,N_27776);
and UO_1130 (O_1130,N_29854,N_27001);
xor UO_1131 (O_1131,N_29787,N_29840);
or UO_1132 (O_1132,N_29782,N_29088);
xnor UO_1133 (O_1133,N_28294,N_28717);
and UO_1134 (O_1134,N_27259,N_28097);
nand UO_1135 (O_1135,N_28608,N_27340);
nor UO_1136 (O_1136,N_29358,N_29748);
nand UO_1137 (O_1137,N_27942,N_28471);
nand UO_1138 (O_1138,N_28452,N_29171);
xnor UO_1139 (O_1139,N_29347,N_28759);
xnor UO_1140 (O_1140,N_27278,N_27650);
xor UO_1141 (O_1141,N_29194,N_27562);
nand UO_1142 (O_1142,N_27427,N_27135);
nor UO_1143 (O_1143,N_29006,N_28981);
or UO_1144 (O_1144,N_27597,N_29150);
and UO_1145 (O_1145,N_28185,N_28952);
nand UO_1146 (O_1146,N_29996,N_28699);
or UO_1147 (O_1147,N_29091,N_29767);
or UO_1148 (O_1148,N_27051,N_28327);
or UO_1149 (O_1149,N_29272,N_27870);
xor UO_1150 (O_1150,N_27409,N_28457);
and UO_1151 (O_1151,N_28194,N_29032);
xnor UO_1152 (O_1152,N_27711,N_28403);
and UO_1153 (O_1153,N_27930,N_29277);
xnor UO_1154 (O_1154,N_28572,N_27989);
nor UO_1155 (O_1155,N_29403,N_28066);
and UO_1156 (O_1156,N_27972,N_27116);
xnor UO_1157 (O_1157,N_28221,N_28767);
or UO_1158 (O_1158,N_28167,N_29827);
xnor UO_1159 (O_1159,N_29991,N_29163);
or UO_1160 (O_1160,N_28157,N_27431);
nor UO_1161 (O_1161,N_27889,N_27999);
nor UO_1162 (O_1162,N_29180,N_27310);
or UO_1163 (O_1163,N_28909,N_29167);
xor UO_1164 (O_1164,N_28908,N_29689);
nor UO_1165 (O_1165,N_29059,N_29384);
nor UO_1166 (O_1166,N_27450,N_27439);
or UO_1167 (O_1167,N_28147,N_29773);
nor UO_1168 (O_1168,N_29448,N_27656);
nand UO_1169 (O_1169,N_27570,N_27806);
and UO_1170 (O_1170,N_29082,N_27291);
nor UO_1171 (O_1171,N_27667,N_29810);
nor UO_1172 (O_1172,N_28204,N_27936);
nand UO_1173 (O_1173,N_27015,N_29324);
nand UO_1174 (O_1174,N_27514,N_28020);
nand UO_1175 (O_1175,N_28341,N_29361);
nand UO_1176 (O_1176,N_28038,N_29943);
or UO_1177 (O_1177,N_29571,N_29570);
nand UO_1178 (O_1178,N_29700,N_29583);
nor UO_1179 (O_1179,N_29263,N_27231);
or UO_1180 (O_1180,N_28849,N_28570);
or UO_1181 (O_1181,N_27592,N_29372);
or UO_1182 (O_1182,N_29525,N_29882);
xor UO_1183 (O_1183,N_27250,N_28521);
nand UO_1184 (O_1184,N_27415,N_28774);
nor UO_1185 (O_1185,N_29113,N_27555);
or UO_1186 (O_1186,N_29615,N_28821);
or UO_1187 (O_1187,N_27804,N_29886);
nand UO_1188 (O_1188,N_29728,N_29339);
or UO_1189 (O_1189,N_27499,N_28065);
xnor UO_1190 (O_1190,N_28101,N_27780);
and UO_1191 (O_1191,N_29730,N_27314);
nor UO_1192 (O_1192,N_27009,N_29560);
and UO_1193 (O_1193,N_27269,N_29806);
or UO_1194 (O_1194,N_28386,N_27787);
nor UO_1195 (O_1195,N_27638,N_29425);
nand UO_1196 (O_1196,N_27507,N_29279);
and UO_1197 (O_1197,N_29697,N_29869);
nand UO_1198 (O_1198,N_27653,N_29790);
and UO_1199 (O_1199,N_27874,N_28279);
nand UO_1200 (O_1200,N_29652,N_29897);
and UO_1201 (O_1201,N_28716,N_29042);
xor UO_1202 (O_1202,N_29883,N_28850);
and UO_1203 (O_1203,N_28365,N_28400);
nor UO_1204 (O_1204,N_28877,N_28845);
nand UO_1205 (O_1205,N_28162,N_29176);
or UO_1206 (O_1206,N_27297,N_29796);
or UO_1207 (O_1207,N_28642,N_29350);
nand UO_1208 (O_1208,N_29852,N_28406);
nor UO_1209 (O_1209,N_29545,N_27556);
nor UO_1210 (O_1210,N_29420,N_27493);
nand UO_1211 (O_1211,N_27824,N_28380);
or UO_1212 (O_1212,N_28861,N_29739);
nor UO_1213 (O_1213,N_29709,N_28222);
xor UO_1214 (O_1214,N_29638,N_28655);
nand UO_1215 (O_1215,N_28797,N_28743);
nand UO_1216 (O_1216,N_28764,N_27247);
nand UO_1217 (O_1217,N_29098,N_27172);
nor UO_1218 (O_1218,N_28994,N_27210);
nand UO_1219 (O_1219,N_29643,N_28355);
or UO_1220 (O_1220,N_27028,N_29343);
or UO_1221 (O_1221,N_27560,N_28172);
and UO_1222 (O_1222,N_29333,N_27336);
and UO_1223 (O_1223,N_29208,N_27630);
nand UO_1224 (O_1224,N_27969,N_27785);
nand UO_1225 (O_1225,N_28019,N_28166);
nor UO_1226 (O_1226,N_27857,N_29494);
or UO_1227 (O_1227,N_27457,N_29731);
and UO_1228 (O_1228,N_27130,N_28581);
or UO_1229 (O_1229,N_27604,N_29878);
or UO_1230 (O_1230,N_29654,N_29789);
nor UO_1231 (O_1231,N_28882,N_29797);
nand UO_1232 (O_1232,N_27649,N_29411);
xor UO_1233 (O_1233,N_28668,N_27451);
nand UO_1234 (O_1234,N_28265,N_28805);
and UO_1235 (O_1235,N_28443,N_29896);
nor UO_1236 (O_1236,N_28618,N_28664);
xor UO_1237 (O_1237,N_28123,N_27880);
and UO_1238 (O_1238,N_28647,N_27404);
xnor UO_1239 (O_1239,N_28806,N_27000);
nand UO_1240 (O_1240,N_27119,N_28280);
nand UO_1241 (O_1241,N_28810,N_28012);
xnor UO_1242 (O_1242,N_29174,N_29116);
or UO_1243 (O_1243,N_27245,N_28193);
nand UO_1244 (O_1244,N_27090,N_27036);
nor UO_1245 (O_1245,N_29072,N_28484);
nor UO_1246 (O_1246,N_29363,N_28059);
nand UO_1247 (O_1247,N_28975,N_29912);
nor UO_1248 (O_1248,N_27859,N_27586);
or UO_1249 (O_1249,N_29097,N_29732);
xor UO_1250 (O_1250,N_28209,N_28746);
xor UO_1251 (O_1251,N_28859,N_29485);
nand UO_1252 (O_1252,N_27858,N_27571);
nor UO_1253 (O_1253,N_29817,N_27751);
nand UO_1254 (O_1254,N_27864,N_28245);
nor UO_1255 (O_1255,N_27786,N_28055);
or UO_1256 (O_1256,N_27337,N_27223);
and UO_1257 (O_1257,N_28253,N_27372);
or UO_1258 (O_1258,N_27768,N_27772);
nor UO_1259 (O_1259,N_29574,N_28818);
and UO_1260 (O_1260,N_27612,N_29999);
and UO_1261 (O_1261,N_28920,N_28826);
and UO_1262 (O_1262,N_29556,N_27610);
nor UO_1263 (O_1263,N_29351,N_28083);
nor UO_1264 (O_1264,N_27887,N_27805);
and UO_1265 (O_1265,N_28906,N_28804);
or UO_1266 (O_1266,N_29102,N_28130);
and UO_1267 (O_1267,N_27769,N_28251);
and UO_1268 (O_1268,N_27124,N_29254);
and UO_1269 (O_1269,N_29455,N_28424);
nand UO_1270 (O_1270,N_29065,N_27024);
nand UO_1271 (O_1271,N_28822,N_28870);
and UO_1272 (O_1272,N_28802,N_28942);
and UO_1273 (O_1273,N_27177,N_29132);
or UO_1274 (O_1274,N_28679,N_27317);
and UO_1275 (O_1275,N_27863,N_29288);
or UO_1276 (O_1276,N_28235,N_29187);
nor UO_1277 (O_1277,N_28261,N_29875);
nor UO_1278 (O_1278,N_29585,N_27506);
nand UO_1279 (O_1279,N_27694,N_29948);
nand UO_1280 (O_1280,N_29960,N_28586);
nor UO_1281 (O_1281,N_28817,N_27654);
nor UO_1282 (O_1282,N_28788,N_28768);
xor UO_1283 (O_1283,N_28082,N_28148);
nand UO_1284 (O_1284,N_28487,N_29115);
nor UO_1285 (O_1285,N_29650,N_29409);
xor UO_1286 (O_1286,N_28156,N_29478);
xnor UO_1287 (O_1287,N_28574,N_29994);
or UO_1288 (O_1288,N_27801,N_29149);
nand UO_1289 (O_1289,N_27267,N_29514);
xor UO_1290 (O_1290,N_28494,N_27265);
nor UO_1291 (O_1291,N_27469,N_28369);
or UO_1292 (O_1292,N_29926,N_28429);
nor UO_1293 (O_1293,N_29110,N_27477);
nand UO_1294 (O_1294,N_28968,N_29177);
and UO_1295 (O_1295,N_28661,N_27893);
xor UO_1296 (O_1296,N_29667,N_27520);
or UO_1297 (O_1297,N_27718,N_28272);
nor UO_1298 (O_1298,N_27699,N_29397);
nand UO_1299 (O_1299,N_28593,N_27350);
or UO_1300 (O_1300,N_27753,N_29075);
or UO_1301 (O_1301,N_29045,N_29775);
nor UO_1302 (O_1302,N_28289,N_28342);
nand UO_1303 (O_1303,N_27581,N_28381);
nand UO_1304 (O_1304,N_27813,N_28986);
nand UO_1305 (O_1305,N_29022,N_28921);
and UO_1306 (O_1306,N_28482,N_28557);
and UO_1307 (O_1307,N_28959,N_29416);
xnor UO_1308 (O_1308,N_29964,N_29296);
xor UO_1309 (O_1309,N_27446,N_29002);
or UO_1310 (O_1310,N_27254,N_27066);
xor UO_1311 (O_1311,N_28617,N_27687);
nor UO_1312 (O_1312,N_28697,N_27528);
or UO_1313 (O_1313,N_27774,N_27308);
nand UO_1314 (O_1314,N_28735,N_28278);
or UO_1315 (O_1315,N_29076,N_28671);
and UO_1316 (O_1316,N_28757,N_27213);
nand UO_1317 (O_1317,N_28107,N_29446);
nand UO_1318 (O_1318,N_28043,N_29204);
or UO_1319 (O_1319,N_27077,N_28852);
and UO_1320 (O_1320,N_27809,N_28709);
nand UO_1321 (O_1321,N_28499,N_28780);
or UO_1322 (O_1322,N_28112,N_28560);
and UO_1323 (O_1323,N_29169,N_29822);
xor UO_1324 (O_1324,N_27584,N_27605);
nor UO_1325 (O_1325,N_29517,N_27448);
or UO_1326 (O_1326,N_28707,N_28863);
nor UO_1327 (O_1327,N_27642,N_29836);
or UO_1328 (O_1328,N_29546,N_29901);
nand UO_1329 (O_1329,N_27021,N_28227);
or UO_1330 (O_1330,N_28307,N_28114);
or UO_1331 (O_1331,N_27081,N_29473);
or UO_1332 (O_1332,N_27374,N_27031);
and UO_1333 (O_1333,N_28190,N_27908);
and UO_1334 (O_1334,N_27459,N_28905);
nand UO_1335 (O_1335,N_29046,N_29917);
nor UO_1336 (O_1336,N_27405,N_29234);
nor UO_1337 (O_1337,N_29230,N_28677);
nand UO_1338 (O_1338,N_27432,N_29232);
nor UO_1339 (O_1339,N_27394,N_29000);
xnor UO_1340 (O_1340,N_28303,N_28481);
or UO_1341 (O_1341,N_28236,N_28524);
nand UO_1342 (O_1342,N_28262,N_29466);
or UO_1343 (O_1343,N_29753,N_27157);
or UO_1344 (O_1344,N_28588,N_28240);
nor UO_1345 (O_1345,N_29979,N_29197);
and UO_1346 (O_1346,N_27068,N_28926);
nand UO_1347 (O_1347,N_28015,N_29218);
xnor UO_1348 (O_1348,N_29057,N_27224);
or UO_1349 (O_1349,N_28192,N_28509);
nand UO_1350 (O_1350,N_29564,N_29291);
and UO_1351 (O_1351,N_29417,N_29825);
and UO_1352 (O_1352,N_28725,N_27219);
nand UO_1353 (O_1353,N_28995,N_29536);
and UO_1354 (O_1354,N_28732,N_28096);
nand UO_1355 (O_1355,N_28037,N_28575);
nand UO_1356 (O_1356,N_28212,N_27716);
and UO_1357 (O_1357,N_29676,N_28795);
nor UO_1358 (O_1358,N_28477,N_27765);
nor UO_1359 (O_1359,N_27973,N_27920);
or UO_1360 (O_1360,N_29993,N_27689);
and UO_1361 (O_1361,N_29675,N_29280);
nand UO_1362 (O_1362,N_27961,N_29932);
and UO_1363 (O_1363,N_28785,N_27652);
and UO_1364 (O_1364,N_27016,N_29253);
or UO_1365 (O_1365,N_29133,N_27173);
or UO_1366 (O_1366,N_28497,N_27251);
or UO_1367 (O_1367,N_28602,N_28468);
nor UO_1368 (O_1368,N_27014,N_27463);
and UO_1369 (O_1369,N_29986,N_28421);
nor UO_1370 (O_1370,N_29726,N_29637);
and UO_1371 (O_1371,N_27364,N_29243);
xnor UO_1372 (O_1372,N_29431,N_28848);
xor UO_1373 (O_1373,N_27239,N_28728);
nor UO_1374 (O_1374,N_29785,N_29734);
and UO_1375 (O_1375,N_28543,N_28230);
or UO_1376 (O_1376,N_28373,N_29422);
nor UO_1377 (O_1377,N_27798,N_27132);
nand UO_1378 (O_1378,N_28532,N_29511);
xnor UO_1379 (O_1379,N_28766,N_29645);
nor UO_1380 (O_1380,N_29058,N_28896);
nand UO_1381 (O_1381,N_27318,N_27243);
or UO_1382 (O_1382,N_29610,N_28030);
nand UO_1383 (O_1383,N_27878,N_29308);
and UO_1384 (O_1384,N_28050,N_27644);
xor UO_1385 (O_1385,N_27352,N_28777);
nor UO_1386 (O_1386,N_28105,N_29432);
xnor UO_1387 (O_1387,N_27854,N_29030);
or UO_1388 (O_1388,N_29913,N_29103);
nand UO_1389 (O_1389,N_29807,N_28401);
xnor UO_1390 (O_1390,N_29762,N_27129);
xnor UO_1391 (O_1391,N_29764,N_29549);
or UO_1392 (O_1392,N_29598,N_27319);
and UO_1393 (O_1393,N_27797,N_29114);
nor UO_1394 (O_1394,N_28980,N_27660);
nand UO_1395 (O_1395,N_28216,N_28024);
nor UO_1396 (O_1396,N_28371,N_29950);
nor UO_1397 (O_1397,N_28999,N_27371);
or UO_1398 (O_1398,N_28326,N_29051);
xor UO_1399 (O_1399,N_27385,N_28816);
nor UO_1400 (O_1400,N_27810,N_27985);
or UO_1401 (O_1401,N_29683,N_29665);
and UO_1402 (O_1402,N_27717,N_28176);
or UO_1403 (O_1403,N_27513,N_27175);
nor UO_1404 (O_1404,N_28333,N_28537);
xor UO_1405 (O_1405,N_29164,N_29493);
or UO_1406 (O_1406,N_28885,N_27816);
nand UO_1407 (O_1407,N_28448,N_29427);
nor UO_1408 (O_1408,N_27046,N_27611);
or UO_1409 (O_1409,N_29137,N_27282);
or UO_1410 (O_1410,N_27559,N_29542);
or UO_1411 (O_1411,N_29527,N_28080);
xnor UO_1412 (O_1412,N_27390,N_29162);
nand UO_1413 (O_1413,N_29147,N_28685);
or UO_1414 (O_1414,N_29888,N_27118);
nor UO_1415 (O_1415,N_29781,N_28446);
or UO_1416 (O_1416,N_27286,N_28489);
and UO_1417 (O_1417,N_29440,N_29894);
nor UO_1418 (O_1418,N_27263,N_27403);
nand UO_1419 (O_1419,N_29687,N_29641);
nand UO_1420 (O_1420,N_28061,N_29828);
xor UO_1421 (O_1421,N_27535,N_27856);
and UO_1422 (O_1422,N_27303,N_29916);
nand UO_1423 (O_1423,N_27709,N_29887);
nand UO_1424 (O_1424,N_29529,N_29919);
and UO_1425 (O_1425,N_28378,N_27676);
or UO_1426 (O_1426,N_27268,N_27113);
and UO_1427 (O_1427,N_27580,N_28453);
and UO_1428 (O_1428,N_27552,N_29619);
or UO_1429 (O_1429,N_28311,N_29481);
nand UO_1430 (O_1430,N_28237,N_27955);
nor UO_1431 (O_1431,N_29453,N_28890);
or UO_1432 (O_1432,N_28583,N_28298);
nor UO_1433 (O_1433,N_27761,N_27721);
nor UO_1434 (O_1434,N_29270,N_28630);
nor UO_1435 (O_1435,N_27206,N_29577);
or UO_1436 (O_1436,N_27641,N_28231);
and UO_1437 (O_1437,N_29008,N_29117);
or UO_1438 (O_1438,N_29752,N_29179);
and UO_1439 (O_1439,N_29491,N_29591);
xor UO_1440 (O_1440,N_28820,N_27621);
nor UO_1441 (O_1441,N_29803,N_27456);
nor UO_1442 (O_1442,N_28270,N_28742);
nand UO_1443 (O_1443,N_29723,N_27965);
nor UO_1444 (O_1444,N_28122,N_28165);
or UO_1445 (O_1445,N_28384,N_29034);
nor UO_1446 (O_1446,N_29106,N_29977);
nor UO_1447 (O_1447,N_28454,N_29145);
nand UO_1448 (O_1448,N_29640,N_29798);
nor UO_1449 (O_1449,N_29942,N_29388);
or UO_1450 (O_1450,N_29584,N_27909);
xnor UO_1451 (O_1451,N_27460,N_28008);
or UO_1452 (O_1452,N_27510,N_29656);
nor UO_1453 (O_1453,N_27196,N_27672);
or UO_1454 (O_1454,N_28689,N_29235);
and UO_1455 (O_1455,N_29725,N_27537);
or UO_1456 (O_1456,N_29877,N_28288);
or UO_1457 (O_1457,N_28599,N_27796);
xor UO_1458 (O_1458,N_28359,N_28143);
nand UO_1459 (O_1459,N_27117,N_28666);
nor UO_1460 (O_1460,N_28673,N_28273);
nand UO_1461 (O_1461,N_29209,N_28432);
or UO_1462 (O_1462,N_29118,N_29377);
and UO_1463 (O_1463,N_28704,N_28603);
nand UO_1464 (O_1464,N_27869,N_28077);
nor UO_1465 (O_1465,N_27516,N_27497);
nor UO_1466 (O_1466,N_27026,N_27598);
and UO_1467 (O_1467,N_27155,N_28283);
nor UO_1468 (O_1468,N_27105,N_28853);
nand UO_1469 (O_1469,N_28946,N_29507);
and UO_1470 (O_1470,N_27168,N_27527);
and UO_1471 (O_1471,N_29565,N_27557);
and UO_1472 (O_1472,N_28232,N_27628);
or UO_1473 (O_1473,N_28385,N_27136);
xor UO_1474 (O_1474,N_27216,N_27923);
or UO_1475 (O_1475,N_27121,N_27883);
nor UO_1476 (O_1476,N_29668,N_27830);
xnor UO_1477 (O_1477,N_27425,N_29369);
or UO_1478 (O_1478,N_27745,N_29414);
and UO_1479 (O_1479,N_28301,N_27311);
nand UO_1480 (O_1480,N_29092,N_29436);
xnor UO_1481 (O_1481,N_28954,N_29152);
and UO_1482 (O_1482,N_28736,N_29937);
nor UO_1483 (O_1483,N_28784,N_29438);
or UO_1484 (O_1484,N_28168,N_27182);
nor UO_1485 (O_1485,N_28783,N_29830);
xnor UO_1486 (O_1486,N_28874,N_27754);
xor UO_1487 (O_1487,N_29670,N_27108);
nor UO_1488 (O_1488,N_29682,N_27410);
xnor UO_1489 (O_1489,N_28011,N_28085);
or UO_1490 (O_1490,N_29329,N_29859);
nor UO_1491 (O_1491,N_28339,N_28686);
and UO_1492 (O_1492,N_29969,N_27814);
xor UO_1493 (O_1493,N_27736,N_28282);
xnor UO_1494 (O_1494,N_27012,N_27525);
nor UO_1495 (O_1495,N_28915,N_28703);
or UO_1496 (O_1496,N_28808,N_28988);
xor UO_1497 (O_1497,N_28799,N_28179);
and UO_1498 (O_1498,N_28215,N_28594);
xor UO_1499 (O_1499,N_29983,N_27332);
and UO_1500 (O_1500,N_27112,N_27264);
nor UO_1501 (O_1501,N_29181,N_27451);
nor UO_1502 (O_1502,N_28306,N_28034);
or UO_1503 (O_1503,N_29694,N_29539);
xor UO_1504 (O_1504,N_27329,N_27414);
or UO_1505 (O_1505,N_28667,N_29583);
nor UO_1506 (O_1506,N_28901,N_28687);
or UO_1507 (O_1507,N_27649,N_27335);
and UO_1508 (O_1508,N_27153,N_29742);
and UO_1509 (O_1509,N_28463,N_29777);
and UO_1510 (O_1510,N_28921,N_28513);
and UO_1511 (O_1511,N_28171,N_28459);
and UO_1512 (O_1512,N_28940,N_29009);
nor UO_1513 (O_1513,N_29667,N_27702);
nor UO_1514 (O_1514,N_27827,N_29553);
and UO_1515 (O_1515,N_29584,N_27146);
or UO_1516 (O_1516,N_29636,N_28555);
or UO_1517 (O_1517,N_27919,N_27018);
or UO_1518 (O_1518,N_29467,N_28824);
nor UO_1519 (O_1519,N_28080,N_29403);
xor UO_1520 (O_1520,N_27267,N_28230);
and UO_1521 (O_1521,N_29384,N_29319);
xor UO_1522 (O_1522,N_29028,N_27557);
or UO_1523 (O_1523,N_28962,N_29372);
or UO_1524 (O_1524,N_27052,N_27236);
and UO_1525 (O_1525,N_28507,N_27093);
or UO_1526 (O_1526,N_28097,N_28970);
or UO_1527 (O_1527,N_28711,N_27365);
xnor UO_1528 (O_1528,N_27001,N_27528);
nand UO_1529 (O_1529,N_27624,N_27301);
and UO_1530 (O_1530,N_29471,N_28736);
nand UO_1531 (O_1531,N_28243,N_29867);
or UO_1532 (O_1532,N_28389,N_28266);
nor UO_1533 (O_1533,N_29639,N_29901);
and UO_1534 (O_1534,N_27512,N_27393);
nor UO_1535 (O_1535,N_29744,N_27434);
or UO_1536 (O_1536,N_27781,N_27580);
and UO_1537 (O_1537,N_28751,N_27089);
or UO_1538 (O_1538,N_27340,N_28813);
or UO_1539 (O_1539,N_27057,N_27723);
xnor UO_1540 (O_1540,N_29677,N_27573);
or UO_1541 (O_1541,N_29816,N_28432);
xor UO_1542 (O_1542,N_29131,N_29096);
and UO_1543 (O_1543,N_27551,N_27466);
xnor UO_1544 (O_1544,N_28074,N_28085);
nand UO_1545 (O_1545,N_28531,N_29081);
and UO_1546 (O_1546,N_27211,N_29302);
or UO_1547 (O_1547,N_27137,N_29776);
and UO_1548 (O_1548,N_27473,N_29186);
and UO_1549 (O_1549,N_29882,N_28159);
xor UO_1550 (O_1550,N_29769,N_29529);
or UO_1551 (O_1551,N_28431,N_27786);
xor UO_1552 (O_1552,N_29433,N_29635);
xnor UO_1553 (O_1553,N_28346,N_27674);
and UO_1554 (O_1554,N_29018,N_27705);
nor UO_1555 (O_1555,N_27166,N_27539);
xnor UO_1556 (O_1556,N_29030,N_29641);
nor UO_1557 (O_1557,N_27245,N_29926);
nand UO_1558 (O_1558,N_29412,N_29148);
nand UO_1559 (O_1559,N_28430,N_29778);
nand UO_1560 (O_1560,N_29316,N_29422);
xor UO_1561 (O_1561,N_29305,N_27161);
nand UO_1562 (O_1562,N_29962,N_28186);
and UO_1563 (O_1563,N_29491,N_28964);
xnor UO_1564 (O_1564,N_27630,N_29936);
and UO_1565 (O_1565,N_27208,N_27942);
nand UO_1566 (O_1566,N_27721,N_27207);
xnor UO_1567 (O_1567,N_29536,N_28487);
or UO_1568 (O_1568,N_29280,N_29545);
xor UO_1569 (O_1569,N_28724,N_29885);
nand UO_1570 (O_1570,N_28233,N_28061);
or UO_1571 (O_1571,N_28433,N_27577);
or UO_1572 (O_1572,N_27499,N_27438);
xnor UO_1573 (O_1573,N_27211,N_29286);
or UO_1574 (O_1574,N_28395,N_29451);
nor UO_1575 (O_1575,N_29970,N_27165);
xnor UO_1576 (O_1576,N_29663,N_28835);
or UO_1577 (O_1577,N_28012,N_28453);
xnor UO_1578 (O_1578,N_28765,N_29214);
nand UO_1579 (O_1579,N_28128,N_29805);
or UO_1580 (O_1580,N_29395,N_27570);
nand UO_1581 (O_1581,N_29858,N_28336);
xnor UO_1582 (O_1582,N_29322,N_28852);
nand UO_1583 (O_1583,N_27260,N_28223);
and UO_1584 (O_1584,N_28702,N_29555);
nor UO_1585 (O_1585,N_27628,N_29049);
nor UO_1586 (O_1586,N_27843,N_27157);
and UO_1587 (O_1587,N_29757,N_28423);
nand UO_1588 (O_1588,N_29312,N_27183);
or UO_1589 (O_1589,N_28294,N_29975);
or UO_1590 (O_1590,N_28561,N_29052);
or UO_1591 (O_1591,N_28556,N_27982);
nor UO_1592 (O_1592,N_27743,N_27147);
and UO_1593 (O_1593,N_27990,N_27753);
and UO_1594 (O_1594,N_27565,N_27261);
nand UO_1595 (O_1595,N_29801,N_28594);
nand UO_1596 (O_1596,N_28245,N_27850);
and UO_1597 (O_1597,N_28645,N_29846);
and UO_1598 (O_1598,N_27367,N_29130);
and UO_1599 (O_1599,N_29341,N_27624);
nor UO_1600 (O_1600,N_29676,N_28731);
nand UO_1601 (O_1601,N_27136,N_29060);
or UO_1602 (O_1602,N_29664,N_29003);
or UO_1603 (O_1603,N_28953,N_28714);
or UO_1604 (O_1604,N_28302,N_28757);
nand UO_1605 (O_1605,N_27519,N_27553);
xor UO_1606 (O_1606,N_27307,N_28745);
nand UO_1607 (O_1607,N_27086,N_29007);
xor UO_1608 (O_1608,N_29187,N_27670);
nand UO_1609 (O_1609,N_28004,N_27533);
and UO_1610 (O_1610,N_28726,N_28682);
nand UO_1611 (O_1611,N_29524,N_27370);
and UO_1612 (O_1612,N_27670,N_27643);
nand UO_1613 (O_1613,N_28889,N_27003);
nor UO_1614 (O_1614,N_29736,N_28191);
or UO_1615 (O_1615,N_28234,N_29648);
xnor UO_1616 (O_1616,N_27481,N_27280);
xnor UO_1617 (O_1617,N_27536,N_29337);
nand UO_1618 (O_1618,N_27635,N_29686);
nand UO_1619 (O_1619,N_28796,N_29864);
or UO_1620 (O_1620,N_29777,N_28077);
nand UO_1621 (O_1621,N_27071,N_29591);
or UO_1622 (O_1622,N_28209,N_27646);
or UO_1623 (O_1623,N_28201,N_28962);
nor UO_1624 (O_1624,N_29856,N_27707);
or UO_1625 (O_1625,N_29450,N_29686);
or UO_1626 (O_1626,N_27720,N_28164);
and UO_1627 (O_1627,N_27739,N_29579);
and UO_1628 (O_1628,N_27411,N_29949);
nand UO_1629 (O_1629,N_27767,N_28452);
nand UO_1630 (O_1630,N_27648,N_27778);
xnor UO_1631 (O_1631,N_28796,N_29602);
nor UO_1632 (O_1632,N_29756,N_28942);
nand UO_1633 (O_1633,N_29367,N_27462);
or UO_1634 (O_1634,N_28468,N_28395);
nand UO_1635 (O_1635,N_29935,N_27683);
xor UO_1636 (O_1636,N_29851,N_28395);
nor UO_1637 (O_1637,N_27391,N_29249);
and UO_1638 (O_1638,N_28273,N_28433);
nand UO_1639 (O_1639,N_29351,N_27072);
nor UO_1640 (O_1640,N_29000,N_27778);
nand UO_1641 (O_1641,N_27919,N_27858);
and UO_1642 (O_1642,N_27281,N_28799);
nand UO_1643 (O_1643,N_28576,N_27663);
xnor UO_1644 (O_1644,N_29625,N_27539);
or UO_1645 (O_1645,N_27405,N_28875);
nor UO_1646 (O_1646,N_28944,N_28962);
and UO_1647 (O_1647,N_27456,N_29391);
and UO_1648 (O_1648,N_28638,N_29213);
nand UO_1649 (O_1649,N_27466,N_28576);
and UO_1650 (O_1650,N_29962,N_27363);
nand UO_1651 (O_1651,N_29244,N_28985);
nor UO_1652 (O_1652,N_28684,N_29187);
and UO_1653 (O_1653,N_28646,N_28090);
nand UO_1654 (O_1654,N_27543,N_27253);
and UO_1655 (O_1655,N_28286,N_27001);
nor UO_1656 (O_1656,N_27360,N_28400);
nor UO_1657 (O_1657,N_29384,N_29009);
nor UO_1658 (O_1658,N_27995,N_29812);
and UO_1659 (O_1659,N_29668,N_27666);
nand UO_1660 (O_1660,N_27463,N_28144);
nand UO_1661 (O_1661,N_27279,N_28067);
nand UO_1662 (O_1662,N_28693,N_28832);
and UO_1663 (O_1663,N_28130,N_28488);
or UO_1664 (O_1664,N_27087,N_27721);
nor UO_1665 (O_1665,N_28746,N_28634);
nand UO_1666 (O_1666,N_29502,N_27488);
nand UO_1667 (O_1667,N_29874,N_28897);
xor UO_1668 (O_1668,N_28243,N_27251);
or UO_1669 (O_1669,N_28566,N_29158);
or UO_1670 (O_1670,N_29214,N_27853);
or UO_1671 (O_1671,N_29732,N_27771);
or UO_1672 (O_1672,N_27883,N_28569);
and UO_1673 (O_1673,N_28970,N_27745);
xnor UO_1674 (O_1674,N_29835,N_28945);
or UO_1675 (O_1675,N_28056,N_28126);
or UO_1676 (O_1676,N_29446,N_28148);
xor UO_1677 (O_1677,N_28222,N_27734);
nor UO_1678 (O_1678,N_28986,N_27309);
or UO_1679 (O_1679,N_29260,N_27028);
nor UO_1680 (O_1680,N_29908,N_28191);
nor UO_1681 (O_1681,N_29260,N_28625);
or UO_1682 (O_1682,N_29865,N_29755);
nand UO_1683 (O_1683,N_29323,N_27918);
xnor UO_1684 (O_1684,N_28960,N_28041);
or UO_1685 (O_1685,N_27223,N_28837);
nand UO_1686 (O_1686,N_27809,N_29222);
and UO_1687 (O_1687,N_28930,N_27950);
xor UO_1688 (O_1688,N_29409,N_27294);
nor UO_1689 (O_1689,N_28659,N_27836);
or UO_1690 (O_1690,N_29453,N_28225);
xnor UO_1691 (O_1691,N_28718,N_27317);
or UO_1692 (O_1692,N_28659,N_29960);
or UO_1693 (O_1693,N_28635,N_27894);
xor UO_1694 (O_1694,N_29390,N_27675);
nor UO_1695 (O_1695,N_29080,N_27480);
or UO_1696 (O_1696,N_27948,N_27928);
nand UO_1697 (O_1697,N_29192,N_28376);
and UO_1698 (O_1698,N_27612,N_28485);
nor UO_1699 (O_1699,N_27361,N_28339);
xor UO_1700 (O_1700,N_27686,N_28407);
nor UO_1701 (O_1701,N_28303,N_28392);
nor UO_1702 (O_1702,N_29145,N_27821);
nor UO_1703 (O_1703,N_28732,N_27514);
nand UO_1704 (O_1704,N_29370,N_27031);
nor UO_1705 (O_1705,N_28616,N_29556);
nor UO_1706 (O_1706,N_28928,N_29516);
or UO_1707 (O_1707,N_28543,N_27800);
nand UO_1708 (O_1708,N_29515,N_28522);
xnor UO_1709 (O_1709,N_27049,N_28346);
nand UO_1710 (O_1710,N_28346,N_28583);
nor UO_1711 (O_1711,N_27900,N_29012);
xnor UO_1712 (O_1712,N_28293,N_29512);
nor UO_1713 (O_1713,N_27845,N_27388);
or UO_1714 (O_1714,N_28516,N_29834);
nand UO_1715 (O_1715,N_29316,N_27701);
or UO_1716 (O_1716,N_27761,N_29891);
xor UO_1717 (O_1717,N_29873,N_27291);
nor UO_1718 (O_1718,N_27313,N_29602);
xnor UO_1719 (O_1719,N_28646,N_29363);
nand UO_1720 (O_1720,N_28711,N_27448);
nand UO_1721 (O_1721,N_28736,N_28932);
xor UO_1722 (O_1722,N_29501,N_28694);
nor UO_1723 (O_1723,N_27333,N_27658);
and UO_1724 (O_1724,N_29047,N_28665);
nand UO_1725 (O_1725,N_28082,N_28077);
or UO_1726 (O_1726,N_29606,N_29035);
and UO_1727 (O_1727,N_29620,N_28258);
xnor UO_1728 (O_1728,N_27788,N_29872);
and UO_1729 (O_1729,N_29443,N_29894);
nor UO_1730 (O_1730,N_27536,N_27008);
nor UO_1731 (O_1731,N_29965,N_27841);
nor UO_1732 (O_1732,N_28756,N_27071);
or UO_1733 (O_1733,N_29528,N_28271);
nor UO_1734 (O_1734,N_28982,N_28156);
and UO_1735 (O_1735,N_28297,N_28536);
nor UO_1736 (O_1736,N_28985,N_29627);
nand UO_1737 (O_1737,N_28273,N_27761);
xnor UO_1738 (O_1738,N_29129,N_28244);
nand UO_1739 (O_1739,N_28234,N_28162);
nor UO_1740 (O_1740,N_27648,N_27605);
or UO_1741 (O_1741,N_28747,N_29197);
or UO_1742 (O_1742,N_27757,N_28228);
nor UO_1743 (O_1743,N_29624,N_29162);
nand UO_1744 (O_1744,N_27086,N_28956);
xor UO_1745 (O_1745,N_27519,N_27201);
and UO_1746 (O_1746,N_29613,N_28418);
nand UO_1747 (O_1747,N_27403,N_28960);
nand UO_1748 (O_1748,N_28207,N_29202);
xnor UO_1749 (O_1749,N_29411,N_28121);
or UO_1750 (O_1750,N_29720,N_29041);
nor UO_1751 (O_1751,N_27071,N_28156);
nand UO_1752 (O_1752,N_27592,N_28527);
nand UO_1753 (O_1753,N_28516,N_29115);
nand UO_1754 (O_1754,N_27312,N_27969);
or UO_1755 (O_1755,N_27897,N_29046);
or UO_1756 (O_1756,N_29647,N_28492);
nor UO_1757 (O_1757,N_28443,N_29408);
nor UO_1758 (O_1758,N_27454,N_28469);
or UO_1759 (O_1759,N_27889,N_28903);
or UO_1760 (O_1760,N_29998,N_28387);
nand UO_1761 (O_1761,N_27684,N_28222);
or UO_1762 (O_1762,N_28120,N_27932);
nor UO_1763 (O_1763,N_28018,N_27048);
or UO_1764 (O_1764,N_29516,N_29883);
nor UO_1765 (O_1765,N_27563,N_28318);
xor UO_1766 (O_1766,N_29947,N_28991);
nor UO_1767 (O_1767,N_29494,N_28396);
nor UO_1768 (O_1768,N_28148,N_29912);
xor UO_1769 (O_1769,N_27114,N_29346);
nand UO_1770 (O_1770,N_29001,N_28445);
xnor UO_1771 (O_1771,N_29363,N_28861);
xnor UO_1772 (O_1772,N_27974,N_29285);
or UO_1773 (O_1773,N_28842,N_27826);
xnor UO_1774 (O_1774,N_27755,N_27319);
xnor UO_1775 (O_1775,N_27351,N_28686);
nand UO_1776 (O_1776,N_28555,N_28887);
and UO_1777 (O_1777,N_28773,N_29204);
and UO_1778 (O_1778,N_29266,N_27250);
or UO_1779 (O_1779,N_28086,N_28823);
or UO_1780 (O_1780,N_27835,N_29528);
or UO_1781 (O_1781,N_29312,N_29343);
xor UO_1782 (O_1782,N_28486,N_29174);
nor UO_1783 (O_1783,N_27919,N_28291);
and UO_1784 (O_1784,N_28414,N_28861);
nand UO_1785 (O_1785,N_28366,N_28081);
and UO_1786 (O_1786,N_28258,N_28325);
nand UO_1787 (O_1787,N_27154,N_28967);
nand UO_1788 (O_1788,N_27751,N_27666);
nand UO_1789 (O_1789,N_29085,N_29981);
or UO_1790 (O_1790,N_27433,N_28119);
nor UO_1791 (O_1791,N_29054,N_27094);
nor UO_1792 (O_1792,N_27616,N_27372);
nand UO_1793 (O_1793,N_28696,N_29882);
nor UO_1794 (O_1794,N_29567,N_27264);
nand UO_1795 (O_1795,N_29405,N_28384);
and UO_1796 (O_1796,N_27830,N_28904);
nor UO_1797 (O_1797,N_28441,N_28535);
nand UO_1798 (O_1798,N_28698,N_28908);
nor UO_1799 (O_1799,N_27225,N_27093);
xnor UO_1800 (O_1800,N_29241,N_29707);
xor UO_1801 (O_1801,N_27744,N_29881);
or UO_1802 (O_1802,N_28867,N_29503);
nor UO_1803 (O_1803,N_28940,N_28441);
nor UO_1804 (O_1804,N_27880,N_28513);
and UO_1805 (O_1805,N_27154,N_27993);
xnor UO_1806 (O_1806,N_29190,N_29665);
or UO_1807 (O_1807,N_28668,N_28062);
or UO_1808 (O_1808,N_28285,N_28089);
xor UO_1809 (O_1809,N_27789,N_27710);
nand UO_1810 (O_1810,N_28015,N_28741);
nand UO_1811 (O_1811,N_29724,N_29570);
or UO_1812 (O_1812,N_29171,N_29982);
xnor UO_1813 (O_1813,N_29400,N_29680);
nand UO_1814 (O_1814,N_27004,N_28516);
or UO_1815 (O_1815,N_29922,N_28617);
and UO_1816 (O_1816,N_27973,N_29656);
and UO_1817 (O_1817,N_29273,N_29772);
xor UO_1818 (O_1818,N_27368,N_29918);
xor UO_1819 (O_1819,N_28837,N_29303);
and UO_1820 (O_1820,N_27027,N_29973);
and UO_1821 (O_1821,N_27129,N_28496);
nand UO_1822 (O_1822,N_27127,N_28742);
nor UO_1823 (O_1823,N_29111,N_29243);
xnor UO_1824 (O_1824,N_28592,N_29215);
nor UO_1825 (O_1825,N_29784,N_28481);
or UO_1826 (O_1826,N_28503,N_27715);
nand UO_1827 (O_1827,N_27494,N_28152);
and UO_1828 (O_1828,N_27387,N_29408);
nor UO_1829 (O_1829,N_27581,N_29389);
or UO_1830 (O_1830,N_28108,N_29123);
and UO_1831 (O_1831,N_29248,N_29215);
nor UO_1832 (O_1832,N_28917,N_29052);
xnor UO_1833 (O_1833,N_29731,N_29340);
xor UO_1834 (O_1834,N_29011,N_28420);
and UO_1835 (O_1835,N_28213,N_27531);
and UO_1836 (O_1836,N_28763,N_27765);
xor UO_1837 (O_1837,N_27621,N_27628);
and UO_1838 (O_1838,N_28082,N_29846);
and UO_1839 (O_1839,N_29887,N_28333);
nor UO_1840 (O_1840,N_28729,N_29891);
or UO_1841 (O_1841,N_28020,N_28886);
xnor UO_1842 (O_1842,N_28559,N_28811);
and UO_1843 (O_1843,N_29214,N_27589);
or UO_1844 (O_1844,N_29092,N_29822);
and UO_1845 (O_1845,N_27398,N_28503);
nor UO_1846 (O_1846,N_28656,N_27555);
xor UO_1847 (O_1847,N_27214,N_29123);
or UO_1848 (O_1848,N_29665,N_29881);
xor UO_1849 (O_1849,N_27873,N_27061);
and UO_1850 (O_1850,N_27077,N_29766);
or UO_1851 (O_1851,N_27909,N_28595);
nor UO_1852 (O_1852,N_29423,N_27886);
and UO_1853 (O_1853,N_28922,N_28864);
nor UO_1854 (O_1854,N_29797,N_29661);
xnor UO_1855 (O_1855,N_29418,N_27024);
xnor UO_1856 (O_1856,N_27397,N_29976);
nand UO_1857 (O_1857,N_28740,N_28535);
or UO_1858 (O_1858,N_27161,N_27271);
xnor UO_1859 (O_1859,N_28666,N_28280);
nand UO_1860 (O_1860,N_27963,N_29954);
or UO_1861 (O_1861,N_28633,N_29197);
nand UO_1862 (O_1862,N_29565,N_28792);
nor UO_1863 (O_1863,N_29152,N_27677);
xor UO_1864 (O_1864,N_29206,N_28109);
and UO_1865 (O_1865,N_29435,N_27212);
nand UO_1866 (O_1866,N_27750,N_28482);
or UO_1867 (O_1867,N_27800,N_27517);
nand UO_1868 (O_1868,N_28692,N_27493);
and UO_1869 (O_1869,N_29980,N_29066);
nand UO_1870 (O_1870,N_29692,N_28075);
or UO_1871 (O_1871,N_27450,N_29874);
or UO_1872 (O_1872,N_29529,N_27258);
or UO_1873 (O_1873,N_27937,N_27358);
and UO_1874 (O_1874,N_27492,N_29399);
or UO_1875 (O_1875,N_27621,N_29461);
xnor UO_1876 (O_1876,N_27624,N_28372);
and UO_1877 (O_1877,N_29518,N_27713);
nand UO_1878 (O_1878,N_29851,N_27014);
or UO_1879 (O_1879,N_29484,N_27774);
xor UO_1880 (O_1880,N_28452,N_28899);
and UO_1881 (O_1881,N_27110,N_27709);
xor UO_1882 (O_1882,N_27395,N_29897);
or UO_1883 (O_1883,N_28809,N_27118);
or UO_1884 (O_1884,N_27164,N_28358);
and UO_1885 (O_1885,N_28442,N_29406);
xnor UO_1886 (O_1886,N_27895,N_27423);
xnor UO_1887 (O_1887,N_29132,N_29130);
and UO_1888 (O_1888,N_27825,N_29549);
or UO_1889 (O_1889,N_28062,N_29794);
or UO_1890 (O_1890,N_28810,N_28630);
xnor UO_1891 (O_1891,N_27356,N_27428);
and UO_1892 (O_1892,N_27512,N_27636);
xor UO_1893 (O_1893,N_29823,N_29333);
and UO_1894 (O_1894,N_29585,N_27776);
nand UO_1895 (O_1895,N_27214,N_28323);
and UO_1896 (O_1896,N_28930,N_28441);
nor UO_1897 (O_1897,N_28307,N_29541);
xor UO_1898 (O_1898,N_28548,N_28456);
nor UO_1899 (O_1899,N_29479,N_29520);
nand UO_1900 (O_1900,N_29723,N_27236);
nand UO_1901 (O_1901,N_29303,N_27775);
or UO_1902 (O_1902,N_29708,N_29225);
nor UO_1903 (O_1903,N_28405,N_27795);
nor UO_1904 (O_1904,N_29083,N_28388);
nand UO_1905 (O_1905,N_27605,N_29506);
or UO_1906 (O_1906,N_28159,N_28955);
or UO_1907 (O_1907,N_29728,N_28783);
and UO_1908 (O_1908,N_28861,N_27049);
xnor UO_1909 (O_1909,N_27457,N_27353);
and UO_1910 (O_1910,N_27709,N_28346);
and UO_1911 (O_1911,N_28248,N_28585);
nor UO_1912 (O_1912,N_28753,N_28722);
nand UO_1913 (O_1913,N_27767,N_29713);
xnor UO_1914 (O_1914,N_29345,N_28067);
and UO_1915 (O_1915,N_27680,N_29480);
nand UO_1916 (O_1916,N_29776,N_28389);
or UO_1917 (O_1917,N_27389,N_29124);
nand UO_1918 (O_1918,N_28842,N_27600);
nor UO_1919 (O_1919,N_29157,N_27980);
and UO_1920 (O_1920,N_27201,N_29935);
nor UO_1921 (O_1921,N_27058,N_28187);
xnor UO_1922 (O_1922,N_27589,N_28508);
nor UO_1923 (O_1923,N_28026,N_27404);
nand UO_1924 (O_1924,N_29817,N_29561);
nand UO_1925 (O_1925,N_28310,N_28693);
xor UO_1926 (O_1926,N_29663,N_27834);
or UO_1927 (O_1927,N_27945,N_27145);
or UO_1928 (O_1928,N_29765,N_27991);
nor UO_1929 (O_1929,N_29677,N_28853);
nand UO_1930 (O_1930,N_29494,N_27055);
and UO_1931 (O_1931,N_28251,N_29499);
xor UO_1932 (O_1932,N_29585,N_27520);
or UO_1933 (O_1933,N_29767,N_28242);
and UO_1934 (O_1934,N_28060,N_29774);
nand UO_1935 (O_1935,N_29389,N_27039);
and UO_1936 (O_1936,N_29593,N_27977);
or UO_1937 (O_1937,N_27946,N_28270);
nor UO_1938 (O_1938,N_28219,N_27049);
nand UO_1939 (O_1939,N_29063,N_29087);
and UO_1940 (O_1940,N_28011,N_29493);
nor UO_1941 (O_1941,N_28964,N_28506);
nand UO_1942 (O_1942,N_29333,N_28602);
or UO_1943 (O_1943,N_29737,N_29846);
or UO_1944 (O_1944,N_27365,N_28008);
nand UO_1945 (O_1945,N_29664,N_27445);
nor UO_1946 (O_1946,N_29679,N_28688);
or UO_1947 (O_1947,N_29349,N_28955);
nand UO_1948 (O_1948,N_28766,N_28006);
nand UO_1949 (O_1949,N_28765,N_29498);
xor UO_1950 (O_1950,N_28955,N_29362);
nor UO_1951 (O_1951,N_27451,N_27394);
or UO_1952 (O_1952,N_28399,N_29191);
or UO_1953 (O_1953,N_28054,N_29242);
nor UO_1954 (O_1954,N_28326,N_27747);
nor UO_1955 (O_1955,N_29337,N_29334);
and UO_1956 (O_1956,N_27958,N_28057);
nor UO_1957 (O_1957,N_27898,N_29709);
or UO_1958 (O_1958,N_28478,N_29718);
xnor UO_1959 (O_1959,N_27698,N_29385);
or UO_1960 (O_1960,N_28269,N_28380);
nand UO_1961 (O_1961,N_27392,N_28256);
nand UO_1962 (O_1962,N_29263,N_27283);
nor UO_1963 (O_1963,N_28796,N_29764);
or UO_1964 (O_1964,N_28856,N_27679);
nand UO_1965 (O_1965,N_27981,N_28783);
nor UO_1966 (O_1966,N_29069,N_27087);
and UO_1967 (O_1967,N_29423,N_28885);
xor UO_1968 (O_1968,N_29728,N_29990);
nor UO_1969 (O_1969,N_29647,N_27691);
and UO_1970 (O_1970,N_29989,N_29938);
or UO_1971 (O_1971,N_29287,N_28875);
xor UO_1972 (O_1972,N_28784,N_27059);
or UO_1973 (O_1973,N_27079,N_28513);
and UO_1974 (O_1974,N_29093,N_29830);
xor UO_1975 (O_1975,N_28338,N_29735);
xor UO_1976 (O_1976,N_27882,N_29425);
or UO_1977 (O_1977,N_28741,N_29750);
xnor UO_1978 (O_1978,N_27941,N_29307);
and UO_1979 (O_1979,N_29370,N_28618);
xor UO_1980 (O_1980,N_28412,N_28938);
nor UO_1981 (O_1981,N_28902,N_28670);
and UO_1982 (O_1982,N_27338,N_28276);
nor UO_1983 (O_1983,N_27101,N_29584);
or UO_1984 (O_1984,N_29471,N_27802);
and UO_1985 (O_1985,N_28003,N_29240);
or UO_1986 (O_1986,N_27728,N_27832);
and UO_1987 (O_1987,N_28608,N_27858);
nor UO_1988 (O_1988,N_29750,N_27721);
and UO_1989 (O_1989,N_28283,N_28121);
or UO_1990 (O_1990,N_28000,N_27558);
and UO_1991 (O_1991,N_28582,N_28527);
nand UO_1992 (O_1992,N_28731,N_28514);
nand UO_1993 (O_1993,N_29383,N_29167);
nand UO_1994 (O_1994,N_28858,N_27817);
xnor UO_1995 (O_1995,N_29454,N_29697);
nor UO_1996 (O_1996,N_29656,N_27439);
xor UO_1997 (O_1997,N_28027,N_27671);
or UO_1998 (O_1998,N_28735,N_27062);
and UO_1999 (O_1999,N_28473,N_29687);
nand UO_2000 (O_2000,N_28042,N_27800);
or UO_2001 (O_2001,N_28879,N_27350);
xnor UO_2002 (O_2002,N_28581,N_27115);
nor UO_2003 (O_2003,N_28865,N_29169);
nand UO_2004 (O_2004,N_29727,N_27416);
and UO_2005 (O_2005,N_29936,N_28456);
or UO_2006 (O_2006,N_28331,N_29611);
nor UO_2007 (O_2007,N_28318,N_29233);
xnor UO_2008 (O_2008,N_28485,N_27362);
or UO_2009 (O_2009,N_28816,N_27904);
and UO_2010 (O_2010,N_27793,N_28919);
nand UO_2011 (O_2011,N_27473,N_28584);
nor UO_2012 (O_2012,N_29617,N_28314);
xnor UO_2013 (O_2013,N_28678,N_29598);
xnor UO_2014 (O_2014,N_27799,N_27371);
xnor UO_2015 (O_2015,N_28493,N_29694);
nand UO_2016 (O_2016,N_28643,N_27441);
nand UO_2017 (O_2017,N_28630,N_28114);
nor UO_2018 (O_2018,N_29337,N_29766);
or UO_2019 (O_2019,N_28156,N_28974);
xnor UO_2020 (O_2020,N_27155,N_29062);
or UO_2021 (O_2021,N_28813,N_28952);
xnor UO_2022 (O_2022,N_29151,N_28505);
nor UO_2023 (O_2023,N_27890,N_27744);
and UO_2024 (O_2024,N_28572,N_27084);
xnor UO_2025 (O_2025,N_27460,N_27974);
nor UO_2026 (O_2026,N_27881,N_27361);
and UO_2027 (O_2027,N_28272,N_29531);
nand UO_2028 (O_2028,N_29759,N_27656);
and UO_2029 (O_2029,N_27211,N_29928);
xnor UO_2030 (O_2030,N_28843,N_29172);
nor UO_2031 (O_2031,N_27418,N_27235);
xnor UO_2032 (O_2032,N_28435,N_29044);
nand UO_2033 (O_2033,N_27269,N_27550);
xor UO_2034 (O_2034,N_29945,N_28837);
nor UO_2035 (O_2035,N_27253,N_27463);
nor UO_2036 (O_2036,N_28094,N_28547);
and UO_2037 (O_2037,N_27921,N_27367);
or UO_2038 (O_2038,N_27633,N_27802);
and UO_2039 (O_2039,N_29175,N_27989);
and UO_2040 (O_2040,N_28742,N_29075);
and UO_2041 (O_2041,N_28396,N_28750);
nor UO_2042 (O_2042,N_27760,N_29032);
nand UO_2043 (O_2043,N_27813,N_27439);
nor UO_2044 (O_2044,N_27186,N_28178);
nor UO_2045 (O_2045,N_27558,N_27552);
nand UO_2046 (O_2046,N_28324,N_28517);
or UO_2047 (O_2047,N_29380,N_29884);
xnor UO_2048 (O_2048,N_29916,N_29867);
nand UO_2049 (O_2049,N_27856,N_29158);
or UO_2050 (O_2050,N_29258,N_28182);
or UO_2051 (O_2051,N_28882,N_29627);
xor UO_2052 (O_2052,N_28340,N_29109);
and UO_2053 (O_2053,N_28012,N_29261);
and UO_2054 (O_2054,N_29245,N_28980);
or UO_2055 (O_2055,N_27025,N_27825);
xor UO_2056 (O_2056,N_29266,N_29440);
and UO_2057 (O_2057,N_29142,N_27691);
xnor UO_2058 (O_2058,N_28922,N_28516);
and UO_2059 (O_2059,N_27665,N_28097);
and UO_2060 (O_2060,N_27095,N_27374);
nand UO_2061 (O_2061,N_27250,N_28714);
nor UO_2062 (O_2062,N_27958,N_27343);
xnor UO_2063 (O_2063,N_27709,N_27200);
nor UO_2064 (O_2064,N_28818,N_27106);
xor UO_2065 (O_2065,N_29746,N_28642);
or UO_2066 (O_2066,N_29491,N_27335);
nand UO_2067 (O_2067,N_27622,N_29124);
nand UO_2068 (O_2068,N_27911,N_28615);
or UO_2069 (O_2069,N_27605,N_28346);
nand UO_2070 (O_2070,N_27122,N_28569);
or UO_2071 (O_2071,N_29350,N_27460);
xnor UO_2072 (O_2072,N_27702,N_27073);
nor UO_2073 (O_2073,N_29061,N_28898);
or UO_2074 (O_2074,N_28237,N_27920);
or UO_2075 (O_2075,N_29969,N_27827);
or UO_2076 (O_2076,N_29885,N_28067);
nand UO_2077 (O_2077,N_29693,N_28854);
or UO_2078 (O_2078,N_27972,N_27047);
and UO_2079 (O_2079,N_27519,N_27748);
and UO_2080 (O_2080,N_27003,N_28042);
xnor UO_2081 (O_2081,N_29158,N_29391);
nand UO_2082 (O_2082,N_28827,N_28336);
nor UO_2083 (O_2083,N_29324,N_27496);
xor UO_2084 (O_2084,N_28353,N_27221);
and UO_2085 (O_2085,N_27846,N_29011);
or UO_2086 (O_2086,N_28685,N_29367);
or UO_2087 (O_2087,N_27539,N_27496);
nor UO_2088 (O_2088,N_28846,N_29077);
xnor UO_2089 (O_2089,N_29930,N_28150);
or UO_2090 (O_2090,N_29523,N_27472);
and UO_2091 (O_2091,N_29865,N_27359);
xnor UO_2092 (O_2092,N_27262,N_27665);
or UO_2093 (O_2093,N_29817,N_29648);
nor UO_2094 (O_2094,N_27535,N_27264);
and UO_2095 (O_2095,N_28079,N_28288);
nor UO_2096 (O_2096,N_29684,N_27611);
nand UO_2097 (O_2097,N_29790,N_29760);
and UO_2098 (O_2098,N_29123,N_29188);
and UO_2099 (O_2099,N_27157,N_28231);
or UO_2100 (O_2100,N_28943,N_29249);
and UO_2101 (O_2101,N_27234,N_28999);
or UO_2102 (O_2102,N_28944,N_28945);
nor UO_2103 (O_2103,N_27920,N_28639);
and UO_2104 (O_2104,N_27373,N_29148);
and UO_2105 (O_2105,N_28723,N_27605);
nand UO_2106 (O_2106,N_27478,N_28102);
and UO_2107 (O_2107,N_29789,N_29017);
or UO_2108 (O_2108,N_29329,N_27969);
xnor UO_2109 (O_2109,N_27499,N_28353);
or UO_2110 (O_2110,N_28266,N_28141);
xor UO_2111 (O_2111,N_28838,N_27819);
nor UO_2112 (O_2112,N_28048,N_29861);
xnor UO_2113 (O_2113,N_28411,N_27875);
and UO_2114 (O_2114,N_27757,N_27901);
or UO_2115 (O_2115,N_28181,N_28236);
and UO_2116 (O_2116,N_27081,N_28873);
xor UO_2117 (O_2117,N_29378,N_29420);
and UO_2118 (O_2118,N_29129,N_28915);
or UO_2119 (O_2119,N_29481,N_28933);
and UO_2120 (O_2120,N_28594,N_28276);
nor UO_2121 (O_2121,N_29572,N_27935);
or UO_2122 (O_2122,N_29693,N_27925);
or UO_2123 (O_2123,N_29180,N_27828);
and UO_2124 (O_2124,N_28276,N_29071);
and UO_2125 (O_2125,N_28095,N_27716);
nor UO_2126 (O_2126,N_28706,N_27310);
nor UO_2127 (O_2127,N_29689,N_27024);
nand UO_2128 (O_2128,N_28035,N_29669);
or UO_2129 (O_2129,N_28345,N_27687);
xor UO_2130 (O_2130,N_29248,N_27715);
nor UO_2131 (O_2131,N_28417,N_29038);
nand UO_2132 (O_2132,N_27999,N_28313);
nor UO_2133 (O_2133,N_28439,N_27883);
nor UO_2134 (O_2134,N_27940,N_27785);
nor UO_2135 (O_2135,N_27242,N_27915);
xnor UO_2136 (O_2136,N_29417,N_28921);
xor UO_2137 (O_2137,N_28565,N_29030);
nand UO_2138 (O_2138,N_27159,N_28515);
or UO_2139 (O_2139,N_28276,N_29947);
xnor UO_2140 (O_2140,N_28329,N_28266);
nor UO_2141 (O_2141,N_28739,N_28135);
nand UO_2142 (O_2142,N_27956,N_28261);
xnor UO_2143 (O_2143,N_28186,N_29483);
nand UO_2144 (O_2144,N_29151,N_27173);
or UO_2145 (O_2145,N_27395,N_28995);
nor UO_2146 (O_2146,N_28135,N_27454);
nor UO_2147 (O_2147,N_28884,N_27769);
and UO_2148 (O_2148,N_29561,N_29528);
xnor UO_2149 (O_2149,N_29022,N_27571);
xor UO_2150 (O_2150,N_28754,N_28889);
nor UO_2151 (O_2151,N_29045,N_28063);
xnor UO_2152 (O_2152,N_29413,N_29723);
xor UO_2153 (O_2153,N_28837,N_27605);
nor UO_2154 (O_2154,N_27508,N_28461);
nor UO_2155 (O_2155,N_29007,N_28338);
or UO_2156 (O_2156,N_27432,N_27817);
and UO_2157 (O_2157,N_29491,N_29438);
xor UO_2158 (O_2158,N_29487,N_28263);
and UO_2159 (O_2159,N_28229,N_28546);
and UO_2160 (O_2160,N_28349,N_28550);
nor UO_2161 (O_2161,N_28050,N_28488);
nor UO_2162 (O_2162,N_29646,N_27867);
nor UO_2163 (O_2163,N_29128,N_27118);
or UO_2164 (O_2164,N_27346,N_29216);
and UO_2165 (O_2165,N_28825,N_29982);
or UO_2166 (O_2166,N_27489,N_28515);
and UO_2167 (O_2167,N_27648,N_27725);
nand UO_2168 (O_2168,N_28719,N_28502);
xor UO_2169 (O_2169,N_27352,N_29919);
nor UO_2170 (O_2170,N_29890,N_27883);
xnor UO_2171 (O_2171,N_29028,N_29139);
nor UO_2172 (O_2172,N_29880,N_29481);
nor UO_2173 (O_2173,N_27959,N_28433);
nand UO_2174 (O_2174,N_27335,N_28216);
xor UO_2175 (O_2175,N_28882,N_29262);
and UO_2176 (O_2176,N_27702,N_27215);
nand UO_2177 (O_2177,N_29901,N_27433);
xor UO_2178 (O_2178,N_28064,N_27125);
nand UO_2179 (O_2179,N_27827,N_27020);
and UO_2180 (O_2180,N_27487,N_29363);
or UO_2181 (O_2181,N_29228,N_29762);
and UO_2182 (O_2182,N_27365,N_27512);
or UO_2183 (O_2183,N_27087,N_28361);
and UO_2184 (O_2184,N_29882,N_29788);
nand UO_2185 (O_2185,N_27266,N_29988);
nand UO_2186 (O_2186,N_28840,N_29806);
nand UO_2187 (O_2187,N_27019,N_28215);
xor UO_2188 (O_2188,N_27759,N_28068);
and UO_2189 (O_2189,N_27341,N_27859);
and UO_2190 (O_2190,N_27588,N_29891);
nand UO_2191 (O_2191,N_27612,N_27004);
nor UO_2192 (O_2192,N_27330,N_29038);
or UO_2193 (O_2193,N_28759,N_27180);
xnor UO_2194 (O_2194,N_28840,N_29654);
and UO_2195 (O_2195,N_28666,N_28776);
xor UO_2196 (O_2196,N_29755,N_27458);
and UO_2197 (O_2197,N_27250,N_27728);
nor UO_2198 (O_2198,N_29178,N_29285);
nor UO_2199 (O_2199,N_27066,N_29176);
and UO_2200 (O_2200,N_29998,N_27983);
xnor UO_2201 (O_2201,N_29106,N_29889);
nand UO_2202 (O_2202,N_28180,N_27424);
xnor UO_2203 (O_2203,N_27142,N_27865);
or UO_2204 (O_2204,N_27581,N_29338);
nor UO_2205 (O_2205,N_29231,N_27324);
and UO_2206 (O_2206,N_27369,N_28254);
and UO_2207 (O_2207,N_28863,N_29081);
and UO_2208 (O_2208,N_27890,N_28801);
nor UO_2209 (O_2209,N_28382,N_27406);
nor UO_2210 (O_2210,N_28566,N_27885);
nand UO_2211 (O_2211,N_27470,N_27266);
nand UO_2212 (O_2212,N_29492,N_27846);
or UO_2213 (O_2213,N_29175,N_28835);
nor UO_2214 (O_2214,N_29174,N_27399);
nor UO_2215 (O_2215,N_29971,N_28232);
xor UO_2216 (O_2216,N_27816,N_28764);
nand UO_2217 (O_2217,N_29128,N_29075);
or UO_2218 (O_2218,N_28410,N_27809);
or UO_2219 (O_2219,N_29263,N_28589);
xnor UO_2220 (O_2220,N_28881,N_27419);
nor UO_2221 (O_2221,N_28352,N_29646);
nor UO_2222 (O_2222,N_29656,N_29198);
and UO_2223 (O_2223,N_27227,N_28452);
nor UO_2224 (O_2224,N_29682,N_28478);
nor UO_2225 (O_2225,N_29820,N_28041);
nor UO_2226 (O_2226,N_27673,N_27166);
xnor UO_2227 (O_2227,N_28538,N_29388);
xnor UO_2228 (O_2228,N_27937,N_29897);
nand UO_2229 (O_2229,N_29583,N_28250);
xnor UO_2230 (O_2230,N_28924,N_28788);
nand UO_2231 (O_2231,N_27908,N_28480);
nand UO_2232 (O_2232,N_27758,N_27326);
and UO_2233 (O_2233,N_27147,N_29792);
nor UO_2234 (O_2234,N_28824,N_27130);
xnor UO_2235 (O_2235,N_27972,N_28045);
xnor UO_2236 (O_2236,N_29784,N_29780);
or UO_2237 (O_2237,N_28505,N_29316);
nand UO_2238 (O_2238,N_27540,N_27212);
and UO_2239 (O_2239,N_27890,N_28689);
nor UO_2240 (O_2240,N_27179,N_28463);
or UO_2241 (O_2241,N_29789,N_28368);
or UO_2242 (O_2242,N_27730,N_27183);
xor UO_2243 (O_2243,N_27849,N_29784);
xnor UO_2244 (O_2244,N_29760,N_27151);
xnor UO_2245 (O_2245,N_27888,N_28222);
and UO_2246 (O_2246,N_27229,N_27758);
xnor UO_2247 (O_2247,N_27869,N_27414);
nor UO_2248 (O_2248,N_27500,N_28947);
and UO_2249 (O_2249,N_29001,N_28224);
and UO_2250 (O_2250,N_27972,N_27823);
nand UO_2251 (O_2251,N_27940,N_27612);
or UO_2252 (O_2252,N_28020,N_28519);
nor UO_2253 (O_2253,N_28248,N_27160);
xnor UO_2254 (O_2254,N_28697,N_27904);
and UO_2255 (O_2255,N_29358,N_28436);
nor UO_2256 (O_2256,N_28707,N_29911);
xnor UO_2257 (O_2257,N_28336,N_29437);
and UO_2258 (O_2258,N_29190,N_28546);
xor UO_2259 (O_2259,N_27617,N_28677);
nand UO_2260 (O_2260,N_27480,N_28848);
nor UO_2261 (O_2261,N_28032,N_28400);
xor UO_2262 (O_2262,N_29539,N_27731);
and UO_2263 (O_2263,N_27794,N_27051);
nand UO_2264 (O_2264,N_29381,N_28651);
xor UO_2265 (O_2265,N_27576,N_29862);
or UO_2266 (O_2266,N_27642,N_27462);
and UO_2267 (O_2267,N_27961,N_27412);
or UO_2268 (O_2268,N_27481,N_29388);
xnor UO_2269 (O_2269,N_29394,N_29990);
or UO_2270 (O_2270,N_28559,N_28259);
xnor UO_2271 (O_2271,N_27331,N_29195);
nand UO_2272 (O_2272,N_27065,N_27310);
xnor UO_2273 (O_2273,N_27346,N_29723);
xnor UO_2274 (O_2274,N_28172,N_28882);
or UO_2275 (O_2275,N_27639,N_27916);
xor UO_2276 (O_2276,N_29291,N_27602);
xnor UO_2277 (O_2277,N_29130,N_29165);
and UO_2278 (O_2278,N_27179,N_27583);
nand UO_2279 (O_2279,N_27508,N_28963);
or UO_2280 (O_2280,N_28749,N_28026);
nand UO_2281 (O_2281,N_28019,N_29861);
or UO_2282 (O_2282,N_29782,N_27247);
nor UO_2283 (O_2283,N_28403,N_27377);
and UO_2284 (O_2284,N_27087,N_27622);
xor UO_2285 (O_2285,N_29191,N_28372);
nor UO_2286 (O_2286,N_28170,N_28887);
xor UO_2287 (O_2287,N_29026,N_29791);
or UO_2288 (O_2288,N_29570,N_27148);
and UO_2289 (O_2289,N_28351,N_28957);
nor UO_2290 (O_2290,N_27140,N_28279);
and UO_2291 (O_2291,N_27311,N_29165);
nor UO_2292 (O_2292,N_27273,N_29266);
nand UO_2293 (O_2293,N_27371,N_28634);
nand UO_2294 (O_2294,N_29629,N_28697);
nor UO_2295 (O_2295,N_27703,N_29425);
and UO_2296 (O_2296,N_29493,N_28230);
xor UO_2297 (O_2297,N_29513,N_27829);
nand UO_2298 (O_2298,N_29636,N_28091);
nor UO_2299 (O_2299,N_27492,N_29707);
nand UO_2300 (O_2300,N_27442,N_29857);
or UO_2301 (O_2301,N_27572,N_28273);
and UO_2302 (O_2302,N_27928,N_28449);
nand UO_2303 (O_2303,N_29076,N_29174);
xnor UO_2304 (O_2304,N_29352,N_29014);
nand UO_2305 (O_2305,N_29734,N_28737);
nor UO_2306 (O_2306,N_27320,N_27301);
and UO_2307 (O_2307,N_28204,N_27839);
xor UO_2308 (O_2308,N_28624,N_29769);
xnor UO_2309 (O_2309,N_28916,N_29339);
and UO_2310 (O_2310,N_28826,N_29576);
nor UO_2311 (O_2311,N_27557,N_27600);
xor UO_2312 (O_2312,N_28777,N_29576);
nor UO_2313 (O_2313,N_27364,N_29993);
nor UO_2314 (O_2314,N_28624,N_29522);
or UO_2315 (O_2315,N_29764,N_27910);
and UO_2316 (O_2316,N_28655,N_27192);
nand UO_2317 (O_2317,N_29817,N_29620);
nor UO_2318 (O_2318,N_29957,N_28981);
xnor UO_2319 (O_2319,N_27421,N_28133);
and UO_2320 (O_2320,N_27558,N_28712);
xor UO_2321 (O_2321,N_27618,N_28496);
nor UO_2322 (O_2322,N_28999,N_29745);
nand UO_2323 (O_2323,N_29192,N_28823);
nor UO_2324 (O_2324,N_27431,N_27470);
and UO_2325 (O_2325,N_27003,N_27467);
xor UO_2326 (O_2326,N_29271,N_27581);
xor UO_2327 (O_2327,N_29371,N_28453);
nand UO_2328 (O_2328,N_27489,N_27152);
or UO_2329 (O_2329,N_27017,N_27717);
nand UO_2330 (O_2330,N_29884,N_27005);
nor UO_2331 (O_2331,N_28672,N_28114);
xor UO_2332 (O_2332,N_28144,N_28143);
nor UO_2333 (O_2333,N_27109,N_29880);
nor UO_2334 (O_2334,N_28418,N_28375);
or UO_2335 (O_2335,N_27157,N_27112);
xnor UO_2336 (O_2336,N_27004,N_28086);
nand UO_2337 (O_2337,N_28678,N_27064);
xor UO_2338 (O_2338,N_29012,N_28774);
and UO_2339 (O_2339,N_27484,N_29153);
nand UO_2340 (O_2340,N_29555,N_27044);
nand UO_2341 (O_2341,N_28992,N_28329);
or UO_2342 (O_2342,N_27557,N_29519);
or UO_2343 (O_2343,N_28774,N_28736);
or UO_2344 (O_2344,N_29818,N_28296);
xor UO_2345 (O_2345,N_28760,N_28200);
and UO_2346 (O_2346,N_27511,N_27340);
or UO_2347 (O_2347,N_28405,N_27434);
or UO_2348 (O_2348,N_29787,N_29972);
nand UO_2349 (O_2349,N_27833,N_28333);
nand UO_2350 (O_2350,N_28073,N_28723);
nand UO_2351 (O_2351,N_28143,N_29014);
nor UO_2352 (O_2352,N_27187,N_29380);
and UO_2353 (O_2353,N_27692,N_29814);
or UO_2354 (O_2354,N_29879,N_29308);
or UO_2355 (O_2355,N_28653,N_27680);
and UO_2356 (O_2356,N_29470,N_28621);
or UO_2357 (O_2357,N_28607,N_28713);
and UO_2358 (O_2358,N_28087,N_28343);
or UO_2359 (O_2359,N_28629,N_27501);
nor UO_2360 (O_2360,N_27767,N_28952);
xnor UO_2361 (O_2361,N_29288,N_28192);
nor UO_2362 (O_2362,N_27179,N_29843);
or UO_2363 (O_2363,N_28181,N_28933);
or UO_2364 (O_2364,N_27630,N_29521);
nand UO_2365 (O_2365,N_29407,N_27183);
xor UO_2366 (O_2366,N_27321,N_28043);
nand UO_2367 (O_2367,N_27129,N_29198);
xor UO_2368 (O_2368,N_28466,N_29942);
nor UO_2369 (O_2369,N_27927,N_27229);
nand UO_2370 (O_2370,N_28708,N_29206);
or UO_2371 (O_2371,N_29018,N_28923);
nand UO_2372 (O_2372,N_27377,N_28633);
or UO_2373 (O_2373,N_29635,N_27212);
nand UO_2374 (O_2374,N_28402,N_28472);
and UO_2375 (O_2375,N_28958,N_29064);
nand UO_2376 (O_2376,N_29068,N_27451);
xnor UO_2377 (O_2377,N_27829,N_29785);
nand UO_2378 (O_2378,N_28747,N_27604);
nand UO_2379 (O_2379,N_27186,N_29251);
nand UO_2380 (O_2380,N_27368,N_29010);
xnor UO_2381 (O_2381,N_29558,N_28752);
nand UO_2382 (O_2382,N_28464,N_29316);
nor UO_2383 (O_2383,N_27767,N_27300);
and UO_2384 (O_2384,N_28668,N_28184);
nor UO_2385 (O_2385,N_27589,N_28939);
or UO_2386 (O_2386,N_28041,N_28930);
or UO_2387 (O_2387,N_27891,N_28825);
xor UO_2388 (O_2388,N_29028,N_29600);
and UO_2389 (O_2389,N_28861,N_29454);
nand UO_2390 (O_2390,N_28478,N_27416);
nand UO_2391 (O_2391,N_29552,N_28426);
and UO_2392 (O_2392,N_27039,N_27085);
nor UO_2393 (O_2393,N_27925,N_28395);
xor UO_2394 (O_2394,N_28949,N_27430);
nor UO_2395 (O_2395,N_29467,N_28597);
xor UO_2396 (O_2396,N_27831,N_27687);
or UO_2397 (O_2397,N_29443,N_27852);
nand UO_2398 (O_2398,N_28251,N_28553);
or UO_2399 (O_2399,N_28758,N_28551);
and UO_2400 (O_2400,N_28286,N_27776);
or UO_2401 (O_2401,N_29939,N_28667);
or UO_2402 (O_2402,N_28794,N_27963);
xnor UO_2403 (O_2403,N_29721,N_28816);
or UO_2404 (O_2404,N_28767,N_29014);
and UO_2405 (O_2405,N_28204,N_29702);
and UO_2406 (O_2406,N_27626,N_29697);
and UO_2407 (O_2407,N_29359,N_27903);
or UO_2408 (O_2408,N_27781,N_29672);
nand UO_2409 (O_2409,N_27729,N_27255);
and UO_2410 (O_2410,N_27491,N_28590);
xnor UO_2411 (O_2411,N_29200,N_29684);
xor UO_2412 (O_2412,N_29985,N_28905);
and UO_2413 (O_2413,N_27240,N_28278);
and UO_2414 (O_2414,N_27914,N_28261);
nand UO_2415 (O_2415,N_28477,N_28491);
xor UO_2416 (O_2416,N_28449,N_29166);
or UO_2417 (O_2417,N_29695,N_28420);
nor UO_2418 (O_2418,N_27042,N_29996);
nand UO_2419 (O_2419,N_28012,N_28876);
xnor UO_2420 (O_2420,N_28118,N_27196);
or UO_2421 (O_2421,N_29469,N_29637);
and UO_2422 (O_2422,N_28584,N_28151);
xnor UO_2423 (O_2423,N_29930,N_29886);
or UO_2424 (O_2424,N_27399,N_28821);
xnor UO_2425 (O_2425,N_29039,N_27532);
and UO_2426 (O_2426,N_28667,N_29648);
xnor UO_2427 (O_2427,N_27745,N_28798);
xnor UO_2428 (O_2428,N_28504,N_28816);
nand UO_2429 (O_2429,N_27841,N_29666);
nor UO_2430 (O_2430,N_27582,N_28143);
and UO_2431 (O_2431,N_29762,N_29783);
xor UO_2432 (O_2432,N_28497,N_27368);
nor UO_2433 (O_2433,N_27321,N_28842);
nand UO_2434 (O_2434,N_28294,N_27421);
xor UO_2435 (O_2435,N_29506,N_29248);
nor UO_2436 (O_2436,N_28923,N_27800);
or UO_2437 (O_2437,N_29192,N_29632);
nand UO_2438 (O_2438,N_29807,N_28086);
nand UO_2439 (O_2439,N_29756,N_28690);
or UO_2440 (O_2440,N_27438,N_27845);
nor UO_2441 (O_2441,N_27705,N_29294);
or UO_2442 (O_2442,N_29885,N_27627);
nor UO_2443 (O_2443,N_27876,N_29923);
xor UO_2444 (O_2444,N_27045,N_28540);
xor UO_2445 (O_2445,N_27584,N_27013);
and UO_2446 (O_2446,N_29109,N_28378);
nand UO_2447 (O_2447,N_28187,N_28795);
or UO_2448 (O_2448,N_29522,N_28498);
or UO_2449 (O_2449,N_28515,N_29103);
or UO_2450 (O_2450,N_27749,N_27643);
nand UO_2451 (O_2451,N_29049,N_28684);
or UO_2452 (O_2452,N_27339,N_27758);
and UO_2453 (O_2453,N_28991,N_29225);
nor UO_2454 (O_2454,N_28296,N_29088);
nand UO_2455 (O_2455,N_28841,N_29729);
nand UO_2456 (O_2456,N_27468,N_28627);
and UO_2457 (O_2457,N_27556,N_28162);
xor UO_2458 (O_2458,N_27365,N_28155);
nor UO_2459 (O_2459,N_27898,N_29085);
or UO_2460 (O_2460,N_28402,N_28689);
xor UO_2461 (O_2461,N_27554,N_28790);
nand UO_2462 (O_2462,N_29612,N_29952);
nor UO_2463 (O_2463,N_27157,N_27410);
and UO_2464 (O_2464,N_27161,N_27718);
xnor UO_2465 (O_2465,N_28148,N_29864);
nand UO_2466 (O_2466,N_28402,N_27780);
nor UO_2467 (O_2467,N_27895,N_27593);
xor UO_2468 (O_2468,N_28974,N_29799);
xnor UO_2469 (O_2469,N_27456,N_29976);
nor UO_2470 (O_2470,N_27332,N_29560);
xor UO_2471 (O_2471,N_29121,N_28834);
and UO_2472 (O_2472,N_29759,N_28173);
or UO_2473 (O_2473,N_28489,N_27520);
xnor UO_2474 (O_2474,N_27448,N_27731);
nor UO_2475 (O_2475,N_28241,N_29947);
xnor UO_2476 (O_2476,N_27999,N_27070);
xnor UO_2477 (O_2477,N_27891,N_28520);
xor UO_2478 (O_2478,N_29199,N_28568);
or UO_2479 (O_2479,N_27334,N_28424);
and UO_2480 (O_2480,N_27600,N_28736);
nand UO_2481 (O_2481,N_29291,N_28604);
nor UO_2482 (O_2482,N_27319,N_28928);
nor UO_2483 (O_2483,N_27306,N_28214);
nor UO_2484 (O_2484,N_29793,N_29099);
nand UO_2485 (O_2485,N_27687,N_28733);
or UO_2486 (O_2486,N_29117,N_28779);
nand UO_2487 (O_2487,N_27177,N_27381);
and UO_2488 (O_2488,N_28083,N_28125);
nand UO_2489 (O_2489,N_28911,N_27649);
or UO_2490 (O_2490,N_27288,N_28107);
or UO_2491 (O_2491,N_27432,N_27178);
nand UO_2492 (O_2492,N_28722,N_29068);
and UO_2493 (O_2493,N_27667,N_29479);
or UO_2494 (O_2494,N_28400,N_29654);
and UO_2495 (O_2495,N_29489,N_27398);
or UO_2496 (O_2496,N_29073,N_29618);
and UO_2497 (O_2497,N_27620,N_29105);
and UO_2498 (O_2498,N_29342,N_28934);
or UO_2499 (O_2499,N_28068,N_27102);
or UO_2500 (O_2500,N_27786,N_28745);
nand UO_2501 (O_2501,N_29884,N_28671);
nor UO_2502 (O_2502,N_28443,N_29428);
or UO_2503 (O_2503,N_28099,N_27093);
and UO_2504 (O_2504,N_29742,N_28227);
and UO_2505 (O_2505,N_29673,N_27295);
or UO_2506 (O_2506,N_28249,N_27514);
nor UO_2507 (O_2507,N_29646,N_28213);
or UO_2508 (O_2508,N_29762,N_29332);
xor UO_2509 (O_2509,N_28801,N_29834);
nand UO_2510 (O_2510,N_29942,N_28569);
nand UO_2511 (O_2511,N_29067,N_29232);
or UO_2512 (O_2512,N_28394,N_29997);
xnor UO_2513 (O_2513,N_28126,N_29538);
xnor UO_2514 (O_2514,N_28389,N_27011);
nand UO_2515 (O_2515,N_28518,N_27612);
nand UO_2516 (O_2516,N_29760,N_27333);
nor UO_2517 (O_2517,N_28509,N_27450);
nand UO_2518 (O_2518,N_28503,N_29198);
nor UO_2519 (O_2519,N_28302,N_29352);
or UO_2520 (O_2520,N_28193,N_28859);
nor UO_2521 (O_2521,N_27070,N_27750);
nand UO_2522 (O_2522,N_29512,N_27872);
xnor UO_2523 (O_2523,N_27002,N_28828);
or UO_2524 (O_2524,N_27901,N_27972);
and UO_2525 (O_2525,N_28157,N_28566);
and UO_2526 (O_2526,N_27945,N_27382);
nand UO_2527 (O_2527,N_29001,N_28844);
and UO_2528 (O_2528,N_28690,N_29436);
xnor UO_2529 (O_2529,N_29439,N_27237);
or UO_2530 (O_2530,N_27062,N_29747);
nor UO_2531 (O_2531,N_29860,N_27641);
or UO_2532 (O_2532,N_29447,N_28387);
and UO_2533 (O_2533,N_29410,N_29612);
and UO_2534 (O_2534,N_27408,N_28535);
xnor UO_2535 (O_2535,N_27693,N_27510);
nor UO_2536 (O_2536,N_29902,N_28954);
nor UO_2537 (O_2537,N_28952,N_29197);
nand UO_2538 (O_2538,N_28600,N_28930);
nand UO_2539 (O_2539,N_28926,N_28520);
or UO_2540 (O_2540,N_29314,N_27727);
or UO_2541 (O_2541,N_28343,N_29227);
nor UO_2542 (O_2542,N_27864,N_28683);
and UO_2543 (O_2543,N_28628,N_29681);
and UO_2544 (O_2544,N_27189,N_28809);
nor UO_2545 (O_2545,N_27656,N_27259);
xnor UO_2546 (O_2546,N_29273,N_28306);
nor UO_2547 (O_2547,N_28810,N_27367);
xor UO_2548 (O_2548,N_27636,N_28404);
and UO_2549 (O_2549,N_29936,N_27449);
xor UO_2550 (O_2550,N_29956,N_28773);
and UO_2551 (O_2551,N_29562,N_28852);
nand UO_2552 (O_2552,N_27176,N_27413);
or UO_2553 (O_2553,N_29557,N_29301);
nand UO_2554 (O_2554,N_27513,N_28269);
xor UO_2555 (O_2555,N_29047,N_28858);
nand UO_2556 (O_2556,N_28490,N_28449);
or UO_2557 (O_2557,N_29982,N_29678);
and UO_2558 (O_2558,N_29573,N_27831);
nor UO_2559 (O_2559,N_27269,N_29104);
nor UO_2560 (O_2560,N_29414,N_29818);
and UO_2561 (O_2561,N_29573,N_29442);
nor UO_2562 (O_2562,N_28477,N_28825);
nand UO_2563 (O_2563,N_28180,N_28679);
nor UO_2564 (O_2564,N_29452,N_27140);
and UO_2565 (O_2565,N_29128,N_27109);
and UO_2566 (O_2566,N_29016,N_28131);
xnor UO_2567 (O_2567,N_29763,N_27601);
or UO_2568 (O_2568,N_29098,N_27564);
and UO_2569 (O_2569,N_29365,N_28591);
nand UO_2570 (O_2570,N_28189,N_27728);
or UO_2571 (O_2571,N_27520,N_27562);
nand UO_2572 (O_2572,N_29294,N_28583);
xor UO_2573 (O_2573,N_28627,N_29268);
or UO_2574 (O_2574,N_27977,N_28832);
xnor UO_2575 (O_2575,N_29043,N_28602);
or UO_2576 (O_2576,N_27657,N_29679);
nand UO_2577 (O_2577,N_27852,N_29021);
nand UO_2578 (O_2578,N_29486,N_28286);
nor UO_2579 (O_2579,N_28377,N_28281);
xnor UO_2580 (O_2580,N_28131,N_27783);
xnor UO_2581 (O_2581,N_27845,N_28743);
xnor UO_2582 (O_2582,N_28425,N_28440);
or UO_2583 (O_2583,N_29021,N_29201);
or UO_2584 (O_2584,N_27741,N_29436);
or UO_2585 (O_2585,N_29006,N_29013);
nor UO_2586 (O_2586,N_29147,N_28548);
or UO_2587 (O_2587,N_27484,N_29510);
nand UO_2588 (O_2588,N_29030,N_27363);
or UO_2589 (O_2589,N_27499,N_29757);
or UO_2590 (O_2590,N_29500,N_27486);
nor UO_2591 (O_2591,N_28367,N_29101);
nand UO_2592 (O_2592,N_29855,N_28042);
and UO_2593 (O_2593,N_27486,N_28736);
and UO_2594 (O_2594,N_29493,N_29938);
nand UO_2595 (O_2595,N_27351,N_27429);
xnor UO_2596 (O_2596,N_29071,N_29181);
or UO_2597 (O_2597,N_29523,N_28879);
nand UO_2598 (O_2598,N_29356,N_28072);
xnor UO_2599 (O_2599,N_28217,N_27521);
and UO_2600 (O_2600,N_29993,N_28376);
or UO_2601 (O_2601,N_28730,N_28687);
or UO_2602 (O_2602,N_27695,N_27134);
or UO_2603 (O_2603,N_27202,N_29245);
xnor UO_2604 (O_2604,N_29803,N_28434);
and UO_2605 (O_2605,N_27599,N_29372);
nand UO_2606 (O_2606,N_29296,N_28252);
nand UO_2607 (O_2607,N_27606,N_28699);
nand UO_2608 (O_2608,N_28088,N_28507);
nand UO_2609 (O_2609,N_27807,N_27182);
xnor UO_2610 (O_2610,N_29280,N_27769);
and UO_2611 (O_2611,N_29915,N_28800);
nor UO_2612 (O_2612,N_27888,N_29824);
or UO_2613 (O_2613,N_27320,N_27498);
nor UO_2614 (O_2614,N_28068,N_28859);
nand UO_2615 (O_2615,N_29899,N_28389);
or UO_2616 (O_2616,N_27841,N_28434);
or UO_2617 (O_2617,N_28146,N_28131);
nor UO_2618 (O_2618,N_28008,N_27609);
xor UO_2619 (O_2619,N_28941,N_29003);
nand UO_2620 (O_2620,N_27228,N_27101);
nor UO_2621 (O_2621,N_27591,N_29891);
or UO_2622 (O_2622,N_27594,N_29520);
xnor UO_2623 (O_2623,N_28826,N_28240);
and UO_2624 (O_2624,N_28382,N_27259);
or UO_2625 (O_2625,N_29495,N_28845);
nand UO_2626 (O_2626,N_28307,N_28503);
nor UO_2627 (O_2627,N_28943,N_27894);
nand UO_2628 (O_2628,N_28604,N_28774);
and UO_2629 (O_2629,N_28304,N_27867);
nor UO_2630 (O_2630,N_27732,N_28657);
xor UO_2631 (O_2631,N_29437,N_29959);
and UO_2632 (O_2632,N_28917,N_29772);
xor UO_2633 (O_2633,N_28306,N_27332);
and UO_2634 (O_2634,N_29721,N_28311);
nor UO_2635 (O_2635,N_27961,N_28868);
nor UO_2636 (O_2636,N_28708,N_29938);
nor UO_2637 (O_2637,N_29828,N_29953);
xor UO_2638 (O_2638,N_28094,N_29438);
xor UO_2639 (O_2639,N_27944,N_27841);
xnor UO_2640 (O_2640,N_28152,N_29105);
nor UO_2641 (O_2641,N_27752,N_29954);
or UO_2642 (O_2642,N_28500,N_27601);
xor UO_2643 (O_2643,N_29432,N_29753);
xor UO_2644 (O_2644,N_27065,N_27222);
xor UO_2645 (O_2645,N_27917,N_28120);
or UO_2646 (O_2646,N_27286,N_28871);
nor UO_2647 (O_2647,N_28209,N_28467);
nand UO_2648 (O_2648,N_27117,N_29715);
xnor UO_2649 (O_2649,N_27125,N_29818);
xnor UO_2650 (O_2650,N_28862,N_27734);
xnor UO_2651 (O_2651,N_28365,N_29433);
nor UO_2652 (O_2652,N_27660,N_29805);
xor UO_2653 (O_2653,N_29679,N_28012);
and UO_2654 (O_2654,N_29057,N_28194);
nor UO_2655 (O_2655,N_27561,N_28111);
nor UO_2656 (O_2656,N_29703,N_29930);
nor UO_2657 (O_2657,N_27566,N_29216);
nor UO_2658 (O_2658,N_29855,N_27570);
nand UO_2659 (O_2659,N_27304,N_29690);
and UO_2660 (O_2660,N_27777,N_29543);
or UO_2661 (O_2661,N_28327,N_28029);
nand UO_2662 (O_2662,N_27175,N_29645);
and UO_2663 (O_2663,N_27183,N_29817);
nand UO_2664 (O_2664,N_28687,N_27330);
nor UO_2665 (O_2665,N_29358,N_28757);
or UO_2666 (O_2666,N_29775,N_27538);
xor UO_2667 (O_2667,N_27989,N_27416);
or UO_2668 (O_2668,N_29249,N_28625);
nor UO_2669 (O_2669,N_28726,N_29646);
xor UO_2670 (O_2670,N_29952,N_28739);
nor UO_2671 (O_2671,N_28246,N_28151);
and UO_2672 (O_2672,N_29074,N_27396);
or UO_2673 (O_2673,N_29954,N_29265);
or UO_2674 (O_2674,N_27314,N_29898);
nor UO_2675 (O_2675,N_27001,N_29586);
nand UO_2676 (O_2676,N_27211,N_29656);
and UO_2677 (O_2677,N_29719,N_28237);
nand UO_2678 (O_2678,N_27614,N_29035);
or UO_2679 (O_2679,N_29095,N_28116);
nor UO_2680 (O_2680,N_28025,N_28442);
nand UO_2681 (O_2681,N_28061,N_29829);
or UO_2682 (O_2682,N_27978,N_29708);
nand UO_2683 (O_2683,N_28469,N_27185);
and UO_2684 (O_2684,N_29853,N_28871);
or UO_2685 (O_2685,N_28294,N_27462);
and UO_2686 (O_2686,N_27827,N_28415);
nor UO_2687 (O_2687,N_29486,N_28039);
xnor UO_2688 (O_2688,N_28520,N_27326);
or UO_2689 (O_2689,N_29702,N_27444);
and UO_2690 (O_2690,N_28818,N_29616);
xnor UO_2691 (O_2691,N_28423,N_28632);
nor UO_2692 (O_2692,N_28071,N_29706);
or UO_2693 (O_2693,N_27382,N_28080);
and UO_2694 (O_2694,N_27982,N_28035);
and UO_2695 (O_2695,N_27235,N_27920);
or UO_2696 (O_2696,N_29252,N_27092);
nand UO_2697 (O_2697,N_29300,N_29357);
nor UO_2698 (O_2698,N_27416,N_28437);
and UO_2699 (O_2699,N_29659,N_28078);
xnor UO_2700 (O_2700,N_27831,N_29983);
xor UO_2701 (O_2701,N_29781,N_28068);
xnor UO_2702 (O_2702,N_28391,N_28241);
and UO_2703 (O_2703,N_27592,N_29631);
xor UO_2704 (O_2704,N_28422,N_27435);
xor UO_2705 (O_2705,N_28531,N_28082);
nor UO_2706 (O_2706,N_27369,N_27317);
xor UO_2707 (O_2707,N_27816,N_28541);
xor UO_2708 (O_2708,N_27104,N_27480);
nand UO_2709 (O_2709,N_27841,N_29308);
xor UO_2710 (O_2710,N_28201,N_28949);
nor UO_2711 (O_2711,N_27604,N_27591);
nand UO_2712 (O_2712,N_27021,N_27891);
or UO_2713 (O_2713,N_27674,N_27454);
nand UO_2714 (O_2714,N_28086,N_29393);
xor UO_2715 (O_2715,N_28904,N_29684);
and UO_2716 (O_2716,N_29947,N_27599);
nand UO_2717 (O_2717,N_29975,N_28187);
xor UO_2718 (O_2718,N_29099,N_28679);
and UO_2719 (O_2719,N_28233,N_28562);
xor UO_2720 (O_2720,N_27075,N_29746);
and UO_2721 (O_2721,N_27135,N_29081);
nor UO_2722 (O_2722,N_28654,N_27402);
nor UO_2723 (O_2723,N_28436,N_29077);
nand UO_2724 (O_2724,N_27090,N_27550);
and UO_2725 (O_2725,N_29188,N_28157);
nor UO_2726 (O_2726,N_28194,N_29253);
and UO_2727 (O_2727,N_29132,N_28719);
nor UO_2728 (O_2728,N_28171,N_29958);
and UO_2729 (O_2729,N_27792,N_27605);
xnor UO_2730 (O_2730,N_28284,N_29379);
or UO_2731 (O_2731,N_27934,N_27222);
or UO_2732 (O_2732,N_27710,N_27003);
and UO_2733 (O_2733,N_29496,N_29644);
nand UO_2734 (O_2734,N_27612,N_28949);
or UO_2735 (O_2735,N_27634,N_28468);
xnor UO_2736 (O_2736,N_29008,N_27347);
and UO_2737 (O_2737,N_27372,N_28125);
or UO_2738 (O_2738,N_29396,N_29863);
or UO_2739 (O_2739,N_29469,N_28573);
and UO_2740 (O_2740,N_28776,N_28862);
xor UO_2741 (O_2741,N_29106,N_27763);
and UO_2742 (O_2742,N_28787,N_28710);
or UO_2743 (O_2743,N_28658,N_29486);
or UO_2744 (O_2744,N_29055,N_28667);
xor UO_2745 (O_2745,N_28623,N_28944);
nand UO_2746 (O_2746,N_28363,N_27817);
nand UO_2747 (O_2747,N_27446,N_29378);
nor UO_2748 (O_2748,N_28026,N_29931);
xnor UO_2749 (O_2749,N_29788,N_28186);
nor UO_2750 (O_2750,N_28056,N_29567);
or UO_2751 (O_2751,N_29530,N_29272);
nor UO_2752 (O_2752,N_29664,N_27041);
or UO_2753 (O_2753,N_27746,N_27677);
and UO_2754 (O_2754,N_27753,N_28333);
xor UO_2755 (O_2755,N_28073,N_29340);
or UO_2756 (O_2756,N_28030,N_29390);
or UO_2757 (O_2757,N_29237,N_28266);
or UO_2758 (O_2758,N_28538,N_27935);
and UO_2759 (O_2759,N_27384,N_28436);
xor UO_2760 (O_2760,N_29231,N_29156);
nor UO_2761 (O_2761,N_29580,N_28892);
or UO_2762 (O_2762,N_28493,N_28952);
and UO_2763 (O_2763,N_29594,N_28899);
xnor UO_2764 (O_2764,N_28916,N_27254);
xnor UO_2765 (O_2765,N_28393,N_29811);
nand UO_2766 (O_2766,N_29648,N_27578);
and UO_2767 (O_2767,N_29109,N_27133);
or UO_2768 (O_2768,N_27456,N_29472);
nand UO_2769 (O_2769,N_28624,N_27143);
xor UO_2770 (O_2770,N_28708,N_27977);
or UO_2771 (O_2771,N_28338,N_27829);
xnor UO_2772 (O_2772,N_28874,N_29973);
nand UO_2773 (O_2773,N_28815,N_28962);
xnor UO_2774 (O_2774,N_29305,N_29044);
or UO_2775 (O_2775,N_29066,N_27080);
or UO_2776 (O_2776,N_27034,N_29025);
or UO_2777 (O_2777,N_27930,N_29035);
nand UO_2778 (O_2778,N_29651,N_27604);
or UO_2779 (O_2779,N_27371,N_27325);
or UO_2780 (O_2780,N_28485,N_27295);
and UO_2781 (O_2781,N_27836,N_28924);
and UO_2782 (O_2782,N_27531,N_27284);
nand UO_2783 (O_2783,N_28726,N_29438);
nor UO_2784 (O_2784,N_28516,N_28683);
nor UO_2785 (O_2785,N_28713,N_27870);
nand UO_2786 (O_2786,N_28268,N_29170);
nor UO_2787 (O_2787,N_27202,N_29855);
and UO_2788 (O_2788,N_28159,N_28106);
xor UO_2789 (O_2789,N_29981,N_29856);
nand UO_2790 (O_2790,N_29554,N_27327);
nor UO_2791 (O_2791,N_28000,N_29003);
nor UO_2792 (O_2792,N_29434,N_27086);
nor UO_2793 (O_2793,N_28396,N_28270);
nor UO_2794 (O_2794,N_29048,N_28617);
nand UO_2795 (O_2795,N_27530,N_27360);
or UO_2796 (O_2796,N_27976,N_27708);
nand UO_2797 (O_2797,N_29824,N_28798);
nand UO_2798 (O_2798,N_27428,N_28291);
xnor UO_2799 (O_2799,N_27193,N_27693);
or UO_2800 (O_2800,N_29080,N_27234);
or UO_2801 (O_2801,N_27778,N_27713);
xor UO_2802 (O_2802,N_27228,N_28368);
and UO_2803 (O_2803,N_28634,N_27098);
and UO_2804 (O_2804,N_28526,N_28539);
or UO_2805 (O_2805,N_29207,N_27525);
nand UO_2806 (O_2806,N_28131,N_29403);
nor UO_2807 (O_2807,N_27629,N_27365);
or UO_2808 (O_2808,N_29328,N_28589);
nor UO_2809 (O_2809,N_28879,N_27364);
and UO_2810 (O_2810,N_29929,N_29147);
or UO_2811 (O_2811,N_28391,N_27885);
or UO_2812 (O_2812,N_29557,N_29782);
xor UO_2813 (O_2813,N_27132,N_28151);
or UO_2814 (O_2814,N_27787,N_28088);
and UO_2815 (O_2815,N_29016,N_27742);
xnor UO_2816 (O_2816,N_29481,N_27654);
nand UO_2817 (O_2817,N_27098,N_27796);
nand UO_2818 (O_2818,N_27446,N_28051);
or UO_2819 (O_2819,N_29654,N_29479);
nor UO_2820 (O_2820,N_28739,N_29610);
nand UO_2821 (O_2821,N_27767,N_28955);
nor UO_2822 (O_2822,N_28879,N_29682);
nor UO_2823 (O_2823,N_27314,N_28922);
or UO_2824 (O_2824,N_28114,N_27347);
xnor UO_2825 (O_2825,N_27206,N_27239);
nor UO_2826 (O_2826,N_27613,N_29176);
nor UO_2827 (O_2827,N_29649,N_27001);
nand UO_2828 (O_2828,N_29747,N_28529);
and UO_2829 (O_2829,N_27319,N_29008);
and UO_2830 (O_2830,N_28498,N_27047);
and UO_2831 (O_2831,N_29969,N_29427);
xor UO_2832 (O_2832,N_27392,N_29347);
nor UO_2833 (O_2833,N_27620,N_28356);
nand UO_2834 (O_2834,N_28800,N_27514);
nand UO_2835 (O_2835,N_29031,N_27083);
xnor UO_2836 (O_2836,N_28879,N_27008);
and UO_2837 (O_2837,N_29902,N_28162);
nor UO_2838 (O_2838,N_29930,N_27180);
and UO_2839 (O_2839,N_29795,N_28392);
nand UO_2840 (O_2840,N_28236,N_29369);
nand UO_2841 (O_2841,N_27129,N_29531);
xor UO_2842 (O_2842,N_29190,N_28556);
xnor UO_2843 (O_2843,N_28703,N_27569);
xnor UO_2844 (O_2844,N_29065,N_28207);
and UO_2845 (O_2845,N_27007,N_27346);
and UO_2846 (O_2846,N_27573,N_29285);
nor UO_2847 (O_2847,N_28161,N_27273);
nor UO_2848 (O_2848,N_29688,N_29436);
nor UO_2849 (O_2849,N_27270,N_27393);
and UO_2850 (O_2850,N_27478,N_28654);
xor UO_2851 (O_2851,N_27421,N_27941);
or UO_2852 (O_2852,N_29288,N_29119);
or UO_2853 (O_2853,N_27898,N_29938);
nor UO_2854 (O_2854,N_28039,N_29030);
nor UO_2855 (O_2855,N_28577,N_29154);
and UO_2856 (O_2856,N_28906,N_27554);
xnor UO_2857 (O_2857,N_28703,N_28363);
or UO_2858 (O_2858,N_29811,N_29225);
and UO_2859 (O_2859,N_29500,N_27733);
nand UO_2860 (O_2860,N_27299,N_27510);
nand UO_2861 (O_2861,N_27771,N_28970);
and UO_2862 (O_2862,N_27431,N_28510);
nand UO_2863 (O_2863,N_27637,N_28584);
nand UO_2864 (O_2864,N_28326,N_28120);
nor UO_2865 (O_2865,N_28525,N_28196);
xnor UO_2866 (O_2866,N_29374,N_28275);
nor UO_2867 (O_2867,N_29053,N_27950);
xnor UO_2868 (O_2868,N_28482,N_28414);
xnor UO_2869 (O_2869,N_28185,N_28536);
xnor UO_2870 (O_2870,N_28985,N_28001);
or UO_2871 (O_2871,N_27920,N_29707);
nor UO_2872 (O_2872,N_27861,N_28548);
xnor UO_2873 (O_2873,N_28086,N_29254);
or UO_2874 (O_2874,N_28624,N_28482);
or UO_2875 (O_2875,N_27044,N_28098);
or UO_2876 (O_2876,N_28232,N_29854);
nor UO_2877 (O_2877,N_29876,N_29304);
xnor UO_2878 (O_2878,N_28960,N_28248);
xor UO_2879 (O_2879,N_28865,N_27941);
and UO_2880 (O_2880,N_27309,N_28156);
or UO_2881 (O_2881,N_29007,N_27834);
nor UO_2882 (O_2882,N_28126,N_27045);
or UO_2883 (O_2883,N_29678,N_29148);
nor UO_2884 (O_2884,N_29501,N_29157);
and UO_2885 (O_2885,N_29483,N_28102);
nand UO_2886 (O_2886,N_27626,N_28259);
nor UO_2887 (O_2887,N_28373,N_29853);
and UO_2888 (O_2888,N_27866,N_28458);
nor UO_2889 (O_2889,N_28277,N_27691);
and UO_2890 (O_2890,N_29075,N_28411);
and UO_2891 (O_2891,N_27566,N_29787);
nor UO_2892 (O_2892,N_28432,N_29686);
and UO_2893 (O_2893,N_29335,N_28957);
and UO_2894 (O_2894,N_27165,N_27414);
or UO_2895 (O_2895,N_29923,N_27005);
or UO_2896 (O_2896,N_27468,N_27002);
or UO_2897 (O_2897,N_29492,N_29235);
and UO_2898 (O_2898,N_28980,N_27133);
nor UO_2899 (O_2899,N_27114,N_29684);
xnor UO_2900 (O_2900,N_27862,N_28218);
xor UO_2901 (O_2901,N_27447,N_28891);
xor UO_2902 (O_2902,N_27304,N_28154);
and UO_2903 (O_2903,N_29036,N_29631);
or UO_2904 (O_2904,N_28365,N_29837);
nor UO_2905 (O_2905,N_29152,N_29653);
xor UO_2906 (O_2906,N_28717,N_28062);
nor UO_2907 (O_2907,N_27957,N_29249);
nand UO_2908 (O_2908,N_27046,N_28001);
xnor UO_2909 (O_2909,N_27609,N_29704);
and UO_2910 (O_2910,N_28288,N_29966);
nor UO_2911 (O_2911,N_28220,N_29879);
nand UO_2912 (O_2912,N_27663,N_28360);
xor UO_2913 (O_2913,N_29289,N_27043);
or UO_2914 (O_2914,N_28012,N_28132);
or UO_2915 (O_2915,N_29709,N_29771);
xnor UO_2916 (O_2916,N_27414,N_29757);
or UO_2917 (O_2917,N_27506,N_28278);
xor UO_2918 (O_2918,N_28170,N_28870);
or UO_2919 (O_2919,N_29839,N_28555);
nand UO_2920 (O_2920,N_28588,N_27032);
xnor UO_2921 (O_2921,N_27422,N_28710);
or UO_2922 (O_2922,N_27625,N_28374);
xnor UO_2923 (O_2923,N_28069,N_28361);
xor UO_2924 (O_2924,N_27907,N_29421);
and UO_2925 (O_2925,N_28161,N_28361);
and UO_2926 (O_2926,N_29662,N_29448);
and UO_2927 (O_2927,N_28038,N_28764);
nor UO_2928 (O_2928,N_29959,N_27696);
or UO_2929 (O_2929,N_29738,N_28585);
nand UO_2930 (O_2930,N_29654,N_29701);
or UO_2931 (O_2931,N_28897,N_29698);
nand UO_2932 (O_2932,N_27849,N_28136);
nor UO_2933 (O_2933,N_27315,N_28751);
nor UO_2934 (O_2934,N_28942,N_28873);
nand UO_2935 (O_2935,N_28912,N_28916);
or UO_2936 (O_2936,N_27269,N_29921);
nor UO_2937 (O_2937,N_27287,N_27726);
and UO_2938 (O_2938,N_29913,N_29797);
or UO_2939 (O_2939,N_27846,N_27687);
nand UO_2940 (O_2940,N_28397,N_29893);
nand UO_2941 (O_2941,N_29874,N_28075);
nor UO_2942 (O_2942,N_27039,N_27089);
and UO_2943 (O_2943,N_28972,N_27165);
nand UO_2944 (O_2944,N_28724,N_27719);
and UO_2945 (O_2945,N_28664,N_28109);
and UO_2946 (O_2946,N_28970,N_27609);
and UO_2947 (O_2947,N_29771,N_27041);
or UO_2948 (O_2948,N_27541,N_29457);
nor UO_2949 (O_2949,N_28850,N_29753);
and UO_2950 (O_2950,N_29411,N_29570);
and UO_2951 (O_2951,N_27377,N_27994);
or UO_2952 (O_2952,N_27026,N_29497);
and UO_2953 (O_2953,N_28008,N_27328);
nor UO_2954 (O_2954,N_28552,N_28785);
or UO_2955 (O_2955,N_28291,N_28165);
nor UO_2956 (O_2956,N_28189,N_29017);
nor UO_2957 (O_2957,N_27169,N_27743);
or UO_2958 (O_2958,N_27451,N_29815);
and UO_2959 (O_2959,N_27673,N_29108);
nand UO_2960 (O_2960,N_27477,N_29092);
or UO_2961 (O_2961,N_29089,N_29735);
and UO_2962 (O_2962,N_29480,N_28458);
and UO_2963 (O_2963,N_29765,N_27083);
xor UO_2964 (O_2964,N_29732,N_29570);
nor UO_2965 (O_2965,N_28640,N_27405);
or UO_2966 (O_2966,N_28909,N_29164);
and UO_2967 (O_2967,N_27547,N_28253);
or UO_2968 (O_2968,N_29809,N_28609);
and UO_2969 (O_2969,N_28041,N_28462);
nand UO_2970 (O_2970,N_28882,N_29381);
xor UO_2971 (O_2971,N_29967,N_28377);
nor UO_2972 (O_2972,N_28799,N_28746);
or UO_2973 (O_2973,N_27866,N_29181);
and UO_2974 (O_2974,N_29101,N_28472);
nand UO_2975 (O_2975,N_28108,N_29088);
nand UO_2976 (O_2976,N_27355,N_29529);
nor UO_2977 (O_2977,N_29302,N_27584);
or UO_2978 (O_2978,N_28522,N_28614);
and UO_2979 (O_2979,N_27965,N_29341);
or UO_2980 (O_2980,N_28334,N_29877);
nor UO_2981 (O_2981,N_28861,N_28982);
and UO_2982 (O_2982,N_28728,N_28842);
nor UO_2983 (O_2983,N_28730,N_27022);
and UO_2984 (O_2984,N_29380,N_27274);
xor UO_2985 (O_2985,N_27365,N_27763);
nor UO_2986 (O_2986,N_29462,N_28303);
nor UO_2987 (O_2987,N_27428,N_27997);
xor UO_2988 (O_2988,N_29527,N_27907);
xnor UO_2989 (O_2989,N_29363,N_28774);
and UO_2990 (O_2990,N_27423,N_29266);
xnor UO_2991 (O_2991,N_28717,N_28631);
nand UO_2992 (O_2992,N_27162,N_29257);
or UO_2993 (O_2993,N_27070,N_29726);
and UO_2994 (O_2994,N_27971,N_27519);
or UO_2995 (O_2995,N_28921,N_28033);
nand UO_2996 (O_2996,N_28175,N_29770);
nand UO_2997 (O_2997,N_29372,N_28985);
nor UO_2998 (O_2998,N_28605,N_27915);
nand UO_2999 (O_2999,N_27445,N_29425);
nand UO_3000 (O_3000,N_28340,N_27742);
nand UO_3001 (O_3001,N_28269,N_29112);
nand UO_3002 (O_3002,N_27949,N_27164);
xnor UO_3003 (O_3003,N_28367,N_28888);
xor UO_3004 (O_3004,N_29989,N_28365);
or UO_3005 (O_3005,N_28409,N_28671);
nand UO_3006 (O_3006,N_27844,N_29494);
and UO_3007 (O_3007,N_27237,N_28162);
nand UO_3008 (O_3008,N_28902,N_28176);
and UO_3009 (O_3009,N_27228,N_28380);
and UO_3010 (O_3010,N_28627,N_29441);
and UO_3011 (O_3011,N_29696,N_29783);
and UO_3012 (O_3012,N_29051,N_27688);
nor UO_3013 (O_3013,N_29283,N_29382);
or UO_3014 (O_3014,N_27490,N_29699);
or UO_3015 (O_3015,N_27053,N_29183);
and UO_3016 (O_3016,N_28901,N_29334);
or UO_3017 (O_3017,N_29221,N_28682);
or UO_3018 (O_3018,N_29012,N_28077);
nor UO_3019 (O_3019,N_27993,N_29224);
nand UO_3020 (O_3020,N_29259,N_27066);
or UO_3021 (O_3021,N_29682,N_28193);
nand UO_3022 (O_3022,N_29851,N_28455);
nand UO_3023 (O_3023,N_28435,N_28650);
nand UO_3024 (O_3024,N_28927,N_27253);
and UO_3025 (O_3025,N_27188,N_28575);
nand UO_3026 (O_3026,N_28271,N_27538);
xor UO_3027 (O_3027,N_28140,N_29795);
nand UO_3028 (O_3028,N_28454,N_27371);
nand UO_3029 (O_3029,N_28097,N_29967);
nand UO_3030 (O_3030,N_28430,N_28856);
and UO_3031 (O_3031,N_28600,N_29473);
or UO_3032 (O_3032,N_29571,N_28941);
and UO_3033 (O_3033,N_28177,N_28728);
xor UO_3034 (O_3034,N_29360,N_28734);
or UO_3035 (O_3035,N_29906,N_28427);
xnor UO_3036 (O_3036,N_27864,N_29027);
nor UO_3037 (O_3037,N_28079,N_27568);
xnor UO_3038 (O_3038,N_29709,N_28214);
nor UO_3039 (O_3039,N_29130,N_28472);
and UO_3040 (O_3040,N_27970,N_28106);
and UO_3041 (O_3041,N_28330,N_27999);
nand UO_3042 (O_3042,N_27988,N_28922);
nand UO_3043 (O_3043,N_27566,N_27027);
nand UO_3044 (O_3044,N_28690,N_28248);
nor UO_3045 (O_3045,N_27543,N_29129);
nor UO_3046 (O_3046,N_27961,N_28382);
nor UO_3047 (O_3047,N_27855,N_29212);
xor UO_3048 (O_3048,N_27756,N_29042);
nand UO_3049 (O_3049,N_28701,N_27260);
nor UO_3050 (O_3050,N_27954,N_27721);
xor UO_3051 (O_3051,N_27417,N_28108);
or UO_3052 (O_3052,N_28173,N_29627);
nor UO_3053 (O_3053,N_27359,N_29175);
and UO_3054 (O_3054,N_27646,N_27467);
xor UO_3055 (O_3055,N_27690,N_29061);
xor UO_3056 (O_3056,N_29322,N_29578);
or UO_3057 (O_3057,N_28486,N_29390);
nand UO_3058 (O_3058,N_29951,N_27878);
nand UO_3059 (O_3059,N_29115,N_27936);
nor UO_3060 (O_3060,N_29211,N_28227);
and UO_3061 (O_3061,N_28330,N_29137);
nand UO_3062 (O_3062,N_28060,N_28953);
and UO_3063 (O_3063,N_29805,N_29397);
nor UO_3064 (O_3064,N_28660,N_28411);
xor UO_3065 (O_3065,N_29820,N_29990);
and UO_3066 (O_3066,N_29976,N_28015);
or UO_3067 (O_3067,N_29649,N_29713);
nor UO_3068 (O_3068,N_27137,N_27394);
xor UO_3069 (O_3069,N_27914,N_27337);
nand UO_3070 (O_3070,N_27293,N_27064);
xor UO_3071 (O_3071,N_29534,N_27159);
nor UO_3072 (O_3072,N_28834,N_28578);
and UO_3073 (O_3073,N_28841,N_29028);
and UO_3074 (O_3074,N_27739,N_27102);
or UO_3075 (O_3075,N_29153,N_27735);
nor UO_3076 (O_3076,N_27749,N_28230);
nand UO_3077 (O_3077,N_29782,N_27547);
xor UO_3078 (O_3078,N_29166,N_27261);
and UO_3079 (O_3079,N_27617,N_28371);
nand UO_3080 (O_3080,N_28005,N_28649);
xor UO_3081 (O_3081,N_28242,N_28272);
xor UO_3082 (O_3082,N_28714,N_28096);
nor UO_3083 (O_3083,N_29168,N_28055);
nand UO_3084 (O_3084,N_27442,N_27292);
and UO_3085 (O_3085,N_28677,N_28767);
or UO_3086 (O_3086,N_27934,N_29612);
nand UO_3087 (O_3087,N_27541,N_28021);
nor UO_3088 (O_3088,N_28201,N_28283);
or UO_3089 (O_3089,N_28763,N_29408);
and UO_3090 (O_3090,N_27856,N_28960);
and UO_3091 (O_3091,N_28967,N_29540);
nor UO_3092 (O_3092,N_28758,N_28419);
or UO_3093 (O_3093,N_28414,N_28425);
nor UO_3094 (O_3094,N_28749,N_29468);
nor UO_3095 (O_3095,N_28404,N_28303);
nand UO_3096 (O_3096,N_27313,N_28375);
nor UO_3097 (O_3097,N_27333,N_29771);
or UO_3098 (O_3098,N_27519,N_29431);
xnor UO_3099 (O_3099,N_28362,N_29920);
nor UO_3100 (O_3100,N_29378,N_29430);
xnor UO_3101 (O_3101,N_27447,N_29566);
or UO_3102 (O_3102,N_29323,N_29069);
nand UO_3103 (O_3103,N_29110,N_29957);
or UO_3104 (O_3104,N_27750,N_28121);
xor UO_3105 (O_3105,N_29505,N_27098);
nand UO_3106 (O_3106,N_29090,N_28809);
nand UO_3107 (O_3107,N_29939,N_27490);
and UO_3108 (O_3108,N_28945,N_28148);
xor UO_3109 (O_3109,N_29860,N_27185);
nand UO_3110 (O_3110,N_29636,N_29148);
nand UO_3111 (O_3111,N_29028,N_28954);
or UO_3112 (O_3112,N_29567,N_28060);
and UO_3113 (O_3113,N_27130,N_27669);
xor UO_3114 (O_3114,N_27167,N_28906);
and UO_3115 (O_3115,N_28758,N_28225);
nor UO_3116 (O_3116,N_28599,N_28024);
or UO_3117 (O_3117,N_28386,N_29770);
nand UO_3118 (O_3118,N_28928,N_27535);
xor UO_3119 (O_3119,N_28592,N_28951);
or UO_3120 (O_3120,N_29530,N_29135);
nand UO_3121 (O_3121,N_27756,N_29357);
or UO_3122 (O_3122,N_29396,N_29269);
or UO_3123 (O_3123,N_29146,N_27304);
and UO_3124 (O_3124,N_28817,N_28966);
nand UO_3125 (O_3125,N_28908,N_29090);
or UO_3126 (O_3126,N_29620,N_29147);
nand UO_3127 (O_3127,N_29718,N_28226);
nand UO_3128 (O_3128,N_27192,N_28422);
nor UO_3129 (O_3129,N_27493,N_27813);
nand UO_3130 (O_3130,N_29914,N_29975);
xor UO_3131 (O_3131,N_29128,N_28259);
or UO_3132 (O_3132,N_28805,N_28219);
xor UO_3133 (O_3133,N_28339,N_27149);
and UO_3134 (O_3134,N_29814,N_27394);
or UO_3135 (O_3135,N_28767,N_27765);
and UO_3136 (O_3136,N_27689,N_29939);
nand UO_3137 (O_3137,N_29955,N_29957);
or UO_3138 (O_3138,N_27216,N_29248);
xnor UO_3139 (O_3139,N_27951,N_29187);
nor UO_3140 (O_3140,N_29783,N_29303);
and UO_3141 (O_3141,N_29035,N_27390);
and UO_3142 (O_3142,N_27226,N_28241);
nand UO_3143 (O_3143,N_29292,N_29152);
or UO_3144 (O_3144,N_28013,N_29055);
nand UO_3145 (O_3145,N_27341,N_29197);
nor UO_3146 (O_3146,N_29437,N_28413);
nor UO_3147 (O_3147,N_28556,N_29545);
nand UO_3148 (O_3148,N_29531,N_29652);
nand UO_3149 (O_3149,N_27125,N_27182);
and UO_3150 (O_3150,N_29008,N_27044);
xnor UO_3151 (O_3151,N_29149,N_29009);
or UO_3152 (O_3152,N_27561,N_27628);
and UO_3153 (O_3153,N_28700,N_29214);
nor UO_3154 (O_3154,N_29383,N_29458);
xor UO_3155 (O_3155,N_28725,N_28334);
nor UO_3156 (O_3156,N_29097,N_28514);
nand UO_3157 (O_3157,N_27846,N_27798);
and UO_3158 (O_3158,N_28412,N_29821);
nor UO_3159 (O_3159,N_29363,N_28475);
nand UO_3160 (O_3160,N_28532,N_27129);
xnor UO_3161 (O_3161,N_29908,N_28512);
or UO_3162 (O_3162,N_29252,N_28135);
nor UO_3163 (O_3163,N_28706,N_27300);
nand UO_3164 (O_3164,N_27278,N_28165);
or UO_3165 (O_3165,N_29588,N_27538);
xor UO_3166 (O_3166,N_27418,N_28215);
nor UO_3167 (O_3167,N_28417,N_29972);
or UO_3168 (O_3168,N_28924,N_27042);
or UO_3169 (O_3169,N_28324,N_28419);
and UO_3170 (O_3170,N_28233,N_28250);
or UO_3171 (O_3171,N_28149,N_27903);
xor UO_3172 (O_3172,N_29552,N_28751);
or UO_3173 (O_3173,N_28614,N_28271);
xnor UO_3174 (O_3174,N_27816,N_29830);
nor UO_3175 (O_3175,N_27495,N_28016);
nor UO_3176 (O_3176,N_28773,N_27701);
nand UO_3177 (O_3177,N_27320,N_28496);
nand UO_3178 (O_3178,N_27674,N_29038);
and UO_3179 (O_3179,N_28451,N_28623);
or UO_3180 (O_3180,N_28129,N_28964);
or UO_3181 (O_3181,N_28071,N_27788);
nand UO_3182 (O_3182,N_29996,N_28347);
nand UO_3183 (O_3183,N_29578,N_27748);
or UO_3184 (O_3184,N_29297,N_29543);
xnor UO_3185 (O_3185,N_27678,N_29352);
or UO_3186 (O_3186,N_27635,N_29526);
or UO_3187 (O_3187,N_27448,N_28206);
or UO_3188 (O_3188,N_29609,N_28837);
and UO_3189 (O_3189,N_28664,N_28175);
or UO_3190 (O_3190,N_29225,N_28909);
nand UO_3191 (O_3191,N_29998,N_29310);
or UO_3192 (O_3192,N_29396,N_29059);
and UO_3193 (O_3193,N_28541,N_27132);
nor UO_3194 (O_3194,N_28513,N_27995);
and UO_3195 (O_3195,N_28130,N_28511);
xnor UO_3196 (O_3196,N_29648,N_28779);
and UO_3197 (O_3197,N_29343,N_27301);
nand UO_3198 (O_3198,N_28782,N_27959);
and UO_3199 (O_3199,N_27948,N_29073);
xnor UO_3200 (O_3200,N_29600,N_28302);
or UO_3201 (O_3201,N_29139,N_27551);
nand UO_3202 (O_3202,N_28197,N_28777);
xor UO_3203 (O_3203,N_27786,N_28998);
nor UO_3204 (O_3204,N_27487,N_29883);
or UO_3205 (O_3205,N_28733,N_27980);
and UO_3206 (O_3206,N_29113,N_28204);
nor UO_3207 (O_3207,N_29512,N_28414);
nor UO_3208 (O_3208,N_29779,N_29331);
or UO_3209 (O_3209,N_29222,N_29399);
nor UO_3210 (O_3210,N_27296,N_29908);
and UO_3211 (O_3211,N_27466,N_29789);
nor UO_3212 (O_3212,N_27343,N_27196);
and UO_3213 (O_3213,N_29077,N_29898);
xnor UO_3214 (O_3214,N_29699,N_28375);
nor UO_3215 (O_3215,N_28444,N_28463);
nor UO_3216 (O_3216,N_28337,N_27957);
nor UO_3217 (O_3217,N_27304,N_29845);
xnor UO_3218 (O_3218,N_28892,N_27639);
or UO_3219 (O_3219,N_27701,N_28111);
xor UO_3220 (O_3220,N_29934,N_28728);
and UO_3221 (O_3221,N_28324,N_28958);
nand UO_3222 (O_3222,N_29404,N_29455);
xnor UO_3223 (O_3223,N_27497,N_28348);
or UO_3224 (O_3224,N_28393,N_29743);
xnor UO_3225 (O_3225,N_29635,N_29886);
xor UO_3226 (O_3226,N_29366,N_27466);
nand UO_3227 (O_3227,N_27366,N_28279);
and UO_3228 (O_3228,N_29878,N_29539);
or UO_3229 (O_3229,N_28766,N_28462);
nor UO_3230 (O_3230,N_29326,N_27443);
nand UO_3231 (O_3231,N_28550,N_28222);
nand UO_3232 (O_3232,N_28191,N_28383);
nand UO_3233 (O_3233,N_28389,N_29599);
xnor UO_3234 (O_3234,N_27364,N_28026);
nand UO_3235 (O_3235,N_28564,N_29209);
nand UO_3236 (O_3236,N_28934,N_27665);
xnor UO_3237 (O_3237,N_29233,N_29821);
or UO_3238 (O_3238,N_28681,N_29603);
and UO_3239 (O_3239,N_27262,N_28779);
xnor UO_3240 (O_3240,N_27485,N_27620);
nor UO_3241 (O_3241,N_27212,N_28682);
xnor UO_3242 (O_3242,N_27120,N_27293);
and UO_3243 (O_3243,N_29809,N_29881);
and UO_3244 (O_3244,N_27315,N_28124);
and UO_3245 (O_3245,N_27606,N_27656);
and UO_3246 (O_3246,N_29253,N_28969);
nand UO_3247 (O_3247,N_29471,N_27736);
nor UO_3248 (O_3248,N_29742,N_29958);
nor UO_3249 (O_3249,N_29302,N_28202);
xor UO_3250 (O_3250,N_28452,N_29452);
or UO_3251 (O_3251,N_28176,N_28762);
xor UO_3252 (O_3252,N_27755,N_27968);
nor UO_3253 (O_3253,N_28208,N_27765);
nor UO_3254 (O_3254,N_27627,N_27049);
or UO_3255 (O_3255,N_29408,N_29430);
nor UO_3256 (O_3256,N_29364,N_27974);
or UO_3257 (O_3257,N_29110,N_28716);
xnor UO_3258 (O_3258,N_29569,N_28368);
and UO_3259 (O_3259,N_28781,N_29159);
nand UO_3260 (O_3260,N_27732,N_27545);
or UO_3261 (O_3261,N_29928,N_27321);
nor UO_3262 (O_3262,N_28375,N_28469);
nor UO_3263 (O_3263,N_28762,N_28484);
nor UO_3264 (O_3264,N_27153,N_27623);
nor UO_3265 (O_3265,N_28746,N_29753);
or UO_3266 (O_3266,N_27019,N_29822);
nor UO_3267 (O_3267,N_29373,N_28566);
nand UO_3268 (O_3268,N_28699,N_29134);
or UO_3269 (O_3269,N_28967,N_29593);
nand UO_3270 (O_3270,N_29630,N_28178);
nand UO_3271 (O_3271,N_29776,N_28690);
nor UO_3272 (O_3272,N_29691,N_27993);
nand UO_3273 (O_3273,N_28489,N_27974);
and UO_3274 (O_3274,N_28533,N_29544);
or UO_3275 (O_3275,N_29452,N_27332);
nor UO_3276 (O_3276,N_27410,N_29568);
and UO_3277 (O_3277,N_28316,N_27044);
nand UO_3278 (O_3278,N_27797,N_28628);
xnor UO_3279 (O_3279,N_27808,N_29107);
nand UO_3280 (O_3280,N_29598,N_29704);
nor UO_3281 (O_3281,N_28268,N_27974);
nor UO_3282 (O_3282,N_28418,N_29572);
and UO_3283 (O_3283,N_28911,N_29733);
nand UO_3284 (O_3284,N_29350,N_28867);
xnor UO_3285 (O_3285,N_27231,N_27166);
xnor UO_3286 (O_3286,N_29710,N_29532);
or UO_3287 (O_3287,N_27189,N_28330);
and UO_3288 (O_3288,N_27450,N_29494);
nor UO_3289 (O_3289,N_29892,N_29156);
nor UO_3290 (O_3290,N_29584,N_28357);
nor UO_3291 (O_3291,N_28510,N_27587);
nand UO_3292 (O_3292,N_28545,N_29914);
nor UO_3293 (O_3293,N_29901,N_28461);
nand UO_3294 (O_3294,N_29891,N_27758);
xor UO_3295 (O_3295,N_28970,N_27456);
or UO_3296 (O_3296,N_29011,N_28592);
or UO_3297 (O_3297,N_28087,N_29092);
xnor UO_3298 (O_3298,N_28016,N_29976);
xnor UO_3299 (O_3299,N_29286,N_29624);
nand UO_3300 (O_3300,N_28318,N_27600);
or UO_3301 (O_3301,N_27488,N_29390);
nor UO_3302 (O_3302,N_28139,N_27362);
nand UO_3303 (O_3303,N_27850,N_27526);
xor UO_3304 (O_3304,N_27583,N_29038);
nor UO_3305 (O_3305,N_28278,N_27946);
and UO_3306 (O_3306,N_28196,N_27766);
nor UO_3307 (O_3307,N_28691,N_27549);
nor UO_3308 (O_3308,N_29624,N_28877);
and UO_3309 (O_3309,N_27078,N_29416);
and UO_3310 (O_3310,N_27768,N_27369);
nor UO_3311 (O_3311,N_28166,N_29751);
or UO_3312 (O_3312,N_27375,N_27746);
nor UO_3313 (O_3313,N_29043,N_28297);
xnor UO_3314 (O_3314,N_27445,N_27123);
nor UO_3315 (O_3315,N_27196,N_28181);
and UO_3316 (O_3316,N_27163,N_28104);
and UO_3317 (O_3317,N_28180,N_27435);
and UO_3318 (O_3318,N_28052,N_29529);
and UO_3319 (O_3319,N_29715,N_29527);
nand UO_3320 (O_3320,N_29124,N_29734);
nor UO_3321 (O_3321,N_27596,N_28933);
and UO_3322 (O_3322,N_28981,N_27116);
or UO_3323 (O_3323,N_27626,N_29984);
or UO_3324 (O_3324,N_29590,N_29555);
nor UO_3325 (O_3325,N_27888,N_27128);
nor UO_3326 (O_3326,N_27445,N_29312);
and UO_3327 (O_3327,N_27952,N_27174);
nand UO_3328 (O_3328,N_28629,N_28881);
nor UO_3329 (O_3329,N_27194,N_27763);
nand UO_3330 (O_3330,N_29076,N_27318);
and UO_3331 (O_3331,N_29931,N_28166);
or UO_3332 (O_3332,N_28013,N_27125);
and UO_3333 (O_3333,N_29220,N_29477);
nor UO_3334 (O_3334,N_29331,N_29873);
or UO_3335 (O_3335,N_27426,N_28624);
nor UO_3336 (O_3336,N_28959,N_27643);
nand UO_3337 (O_3337,N_27150,N_28187);
nor UO_3338 (O_3338,N_28236,N_28034);
and UO_3339 (O_3339,N_29685,N_28471);
nor UO_3340 (O_3340,N_27949,N_29607);
xor UO_3341 (O_3341,N_28274,N_27929);
and UO_3342 (O_3342,N_29142,N_29233);
and UO_3343 (O_3343,N_29777,N_28467);
nand UO_3344 (O_3344,N_29217,N_27815);
nor UO_3345 (O_3345,N_27768,N_28858);
xnor UO_3346 (O_3346,N_29523,N_28605);
and UO_3347 (O_3347,N_27551,N_27888);
or UO_3348 (O_3348,N_27007,N_27180);
and UO_3349 (O_3349,N_29393,N_28296);
nand UO_3350 (O_3350,N_28500,N_29559);
nor UO_3351 (O_3351,N_27512,N_29861);
or UO_3352 (O_3352,N_28260,N_29000);
or UO_3353 (O_3353,N_27921,N_29432);
xnor UO_3354 (O_3354,N_28676,N_29847);
nand UO_3355 (O_3355,N_27171,N_27703);
nand UO_3356 (O_3356,N_29871,N_27322);
nand UO_3357 (O_3357,N_28777,N_28367);
xnor UO_3358 (O_3358,N_29361,N_27661);
xor UO_3359 (O_3359,N_29110,N_28116);
and UO_3360 (O_3360,N_28567,N_29459);
nor UO_3361 (O_3361,N_29031,N_29687);
xnor UO_3362 (O_3362,N_29678,N_28064);
or UO_3363 (O_3363,N_28587,N_27756);
or UO_3364 (O_3364,N_28784,N_28439);
or UO_3365 (O_3365,N_28905,N_28791);
or UO_3366 (O_3366,N_28208,N_29779);
xor UO_3367 (O_3367,N_28926,N_27328);
nor UO_3368 (O_3368,N_27190,N_28823);
and UO_3369 (O_3369,N_29803,N_27602);
nand UO_3370 (O_3370,N_28603,N_27244);
nand UO_3371 (O_3371,N_29494,N_29235);
and UO_3372 (O_3372,N_27725,N_27979);
xnor UO_3373 (O_3373,N_28021,N_28015);
nand UO_3374 (O_3374,N_29299,N_29262);
nand UO_3375 (O_3375,N_27698,N_27349);
xnor UO_3376 (O_3376,N_28615,N_28701);
nand UO_3377 (O_3377,N_28573,N_28638);
nor UO_3378 (O_3378,N_27877,N_27632);
nand UO_3379 (O_3379,N_27808,N_29756);
nor UO_3380 (O_3380,N_27874,N_29897);
nand UO_3381 (O_3381,N_29502,N_29944);
nor UO_3382 (O_3382,N_29544,N_29658);
xor UO_3383 (O_3383,N_29651,N_27233);
or UO_3384 (O_3384,N_27079,N_27220);
xor UO_3385 (O_3385,N_28873,N_29645);
nor UO_3386 (O_3386,N_29823,N_29453);
nor UO_3387 (O_3387,N_28754,N_28804);
or UO_3388 (O_3388,N_29309,N_27216);
or UO_3389 (O_3389,N_27463,N_29072);
xnor UO_3390 (O_3390,N_28255,N_29639);
xnor UO_3391 (O_3391,N_27566,N_27986);
or UO_3392 (O_3392,N_28240,N_29983);
nand UO_3393 (O_3393,N_28807,N_29922);
or UO_3394 (O_3394,N_27277,N_29200);
or UO_3395 (O_3395,N_28132,N_27762);
nand UO_3396 (O_3396,N_27700,N_27687);
nand UO_3397 (O_3397,N_28925,N_28145);
nand UO_3398 (O_3398,N_28620,N_28808);
and UO_3399 (O_3399,N_29850,N_29758);
or UO_3400 (O_3400,N_28555,N_27099);
nor UO_3401 (O_3401,N_29833,N_27695);
xor UO_3402 (O_3402,N_27950,N_28387);
xnor UO_3403 (O_3403,N_29575,N_28331);
nand UO_3404 (O_3404,N_27516,N_27136);
nor UO_3405 (O_3405,N_27219,N_29140);
xnor UO_3406 (O_3406,N_27855,N_27679);
nor UO_3407 (O_3407,N_29476,N_27238);
nand UO_3408 (O_3408,N_29121,N_28600);
nand UO_3409 (O_3409,N_29737,N_27319);
xor UO_3410 (O_3410,N_28768,N_27931);
nor UO_3411 (O_3411,N_28540,N_27338);
nand UO_3412 (O_3412,N_29160,N_28541);
or UO_3413 (O_3413,N_27618,N_29803);
xnor UO_3414 (O_3414,N_29865,N_27709);
nand UO_3415 (O_3415,N_29188,N_29946);
and UO_3416 (O_3416,N_29254,N_29701);
xnor UO_3417 (O_3417,N_27450,N_28989);
nand UO_3418 (O_3418,N_27528,N_29526);
nand UO_3419 (O_3419,N_27269,N_29755);
nor UO_3420 (O_3420,N_29188,N_29903);
or UO_3421 (O_3421,N_28624,N_27367);
nor UO_3422 (O_3422,N_27375,N_29874);
nand UO_3423 (O_3423,N_28645,N_29739);
xnor UO_3424 (O_3424,N_29102,N_27958);
nor UO_3425 (O_3425,N_29547,N_28682);
or UO_3426 (O_3426,N_29618,N_28126);
nor UO_3427 (O_3427,N_29334,N_28924);
nor UO_3428 (O_3428,N_29078,N_29066);
nor UO_3429 (O_3429,N_27835,N_27433);
xnor UO_3430 (O_3430,N_28525,N_29065);
and UO_3431 (O_3431,N_27182,N_27679);
or UO_3432 (O_3432,N_29732,N_27768);
xor UO_3433 (O_3433,N_27144,N_29227);
nand UO_3434 (O_3434,N_28287,N_28955);
xor UO_3435 (O_3435,N_29959,N_28500);
or UO_3436 (O_3436,N_29417,N_29792);
and UO_3437 (O_3437,N_29793,N_27645);
xnor UO_3438 (O_3438,N_29224,N_29251);
nor UO_3439 (O_3439,N_28968,N_28573);
and UO_3440 (O_3440,N_27000,N_29395);
nor UO_3441 (O_3441,N_29402,N_27977);
and UO_3442 (O_3442,N_29279,N_28057);
or UO_3443 (O_3443,N_27713,N_27501);
xor UO_3444 (O_3444,N_28655,N_28114);
or UO_3445 (O_3445,N_27391,N_27823);
nor UO_3446 (O_3446,N_27308,N_29551);
nor UO_3447 (O_3447,N_28079,N_28303);
or UO_3448 (O_3448,N_29117,N_27152);
or UO_3449 (O_3449,N_28089,N_27093);
nor UO_3450 (O_3450,N_29418,N_27460);
nor UO_3451 (O_3451,N_28832,N_27661);
nor UO_3452 (O_3452,N_27383,N_29342);
nand UO_3453 (O_3453,N_27108,N_28908);
nand UO_3454 (O_3454,N_28759,N_29311);
and UO_3455 (O_3455,N_29504,N_28093);
nor UO_3456 (O_3456,N_29891,N_29630);
nand UO_3457 (O_3457,N_28308,N_27971);
and UO_3458 (O_3458,N_28772,N_29246);
xor UO_3459 (O_3459,N_27921,N_29352);
xor UO_3460 (O_3460,N_28655,N_27300);
nand UO_3461 (O_3461,N_28917,N_27761);
nor UO_3462 (O_3462,N_28363,N_29392);
and UO_3463 (O_3463,N_29807,N_27664);
xor UO_3464 (O_3464,N_29671,N_27189);
nand UO_3465 (O_3465,N_28573,N_27395);
nand UO_3466 (O_3466,N_27113,N_28512);
and UO_3467 (O_3467,N_27301,N_29040);
or UO_3468 (O_3468,N_29765,N_28656);
xor UO_3469 (O_3469,N_28268,N_27313);
and UO_3470 (O_3470,N_27834,N_27593);
nand UO_3471 (O_3471,N_29387,N_28976);
and UO_3472 (O_3472,N_28221,N_29289);
or UO_3473 (O_3473,N_27465,N_28686);
nand UO_3474 (O_3474,N_27384,N_29311);
nand UO_3475 (O_3475,N_28642,N_29777);
nand UO_3476 (O_3476,N_27755,N_27962);
xor UO_3477 (O_3477,N_28556,N_28364);
nor UO_3478 (O_3478,N_29122,N_29902);
xnor UO_3479 (O_3479,N_28908,N_29713);
and UO_3480 (O_3480,N_29475,N_28653);
nand UO_3481 (O_3481,N_29563,N_28819);
nand UO_3482 (O_3482,N_27564,N_29961);
nor UO_3483 (O_3483,N_28232,N_28635);
and UO_3484 (O_3484,N_29081,N_27531);
xnor UO_3485 (O_3485,N_27075,N_29441);
xor UO_3486 (O_3486,N_27860,N_28543);
nor UO_3487 (O_3487,N_27657,N_29546);
xor UO_3488 (O_3488,N_29452,N_29190);
or UO_3489 (O_3489,N_29741,N_28191);
and UO_3490 (O_3490,N_28714,N_29707);
or UO_3491 (O_3491,N_29386,N_27100);
nor UO_3492 (O_3492,N_29547,N_27102);
nand UO_3493 (O_3493,N_29939,N_28935);
nor UO_3494 (O_3494,N_29244,N_29704);
nand UO_3495 (O_3495,N_28535,N_27854);
or UO_3496 (O_3496,N_29864,N_28037);
nand UO_3497 (O_3497,N_28022,N_27472);
nor UO_3498 (O_3498,N_29276,N_28820);
nor UO_3499 (O_3499,N_29204,N_27184);
endmodule