module basic_500_3000_500_15_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_416,In_452);
nor U1 (N_1,In_151,In_178);
nor U2 (N_2,In_67,In_74);
or U3 (N_3,In_302,In_454);
nor U4 (N_4,In_110,In_356);
nor U5 (N_5,In_13,In_282);
and U6 (N_6,In_426,In_180);
and U7 (N_7,In_372,In_8);
or U8 (N_8,In_158,In_487);
or U9 (N_9,In_106,In_171);
and U10 (N_10,In_463,In_131);
and U11 (N_11,In_207,In_437);
and U12 (N_12,In_232,In_137);
nor U13 (N_13,In_192,In_223);
and U14 (N_14,In_349,In_436);
nor U15 (N_15,In_287,In_371);
nor U16 (N_16,In_98,In_147);
nor U17 (N_17,In_145,In_239);
and U18 (N_18,In_225,In_400);
or U19 (N_19,In_319,In_99);
xor U20 (N_20,In_182,In_275);
nor U21 (N_21,In_26,In_217);
nand U22 (N_22,In_176,In_21);
nand U23 (N_23,In_413,In_261);
and U24 (N_24,In_230,In_353);
nor U25 (N_25,In_332,In_189);
or U26 (N_26,In_85,In_414);
and U27 (N_27,In_455,In_245);
nor U28 (N_28,In_377,In_354);
nor U29 (N_29,In_72,In_485);
and U30 (N_30,In_351,In_36);
nor U31 (N_31,In_34,In_61);
nand U32 (N_32,In_347,In_394);
and U33 (N_33,In_248,In_361);
nand U34 (N_34,In_267,In_272);
xor U35 (N_35,In_247,In_144);
nand U36 (N_36,In_474,In_270);
nand U37 (N_37,In_493,In_460);
nor U38 (N_38,In_136,In_105);
and U39 (N_39,In_308,In_316);
nand U40 (N_40,In_38,In_3);
or U41 (N_41,In_459,In_229);
nand U42 (N_42,In_100,In_449);
and U43 (N_43,In_325,In_305);
and U44 (N_44,In_9,In_32);
nand U45 (N_45,In_54,In_381);
or U46 (N_46,In_346,In_139);
and U47 (N_47,In_355,In_240);
nor U48 (N_48,In_7,In_0);
or U49 (N_49,In_333,In_309);
nor U50 (N_50,In_458,In_200);
nand U51 (N_51,In_42,In_24);
and U52 (N_52,In_29,In_442);
or U53 (N_53,In_484,In_107);
nor U54 (N_54,In_15,In_256);
nor U55 (N_55,In_89,In_111);
and U56 (N_56,In_411,In_167);
and U57 (N_57,In_191,In_380);
nor U58 (N_58,In_255,In_64);
nand U59 (N_59,In_90,In_314);
and U60 (N_60,In_165,In_370);
and U61 (N_61,In_258,In_159);
nand U62 (N_62,In_253,In_296);
nor U63 (N_63,In_284,In_448);
and U64 (N_64,In_271,In_367);
or U65 (N_65,In_249,In_444);
nand U66 (N_66,In_430,In_334);
nand U67 (N_67,In_93,In_423);
or U68 (N_68,In_175,In_348);
xor U69 (N_69,In_149,In_386);
and U70 (N_70,In_121,In_198);
nor U71 (N_71,In_290,In_483);
nor U72 (N_72,In_438,In_273);
or U73 (N_73,In_83,In_395);
or U74 (N_74,In_1,In_286);
or U75 (N_75,In_146,In_174);
nor U76 (N_76,In_57,In_405);
and U77 (N_77,In_119,In_257);
and U78 (N_78,In_313,In_221);
nor U79 (N_79,In_6,In_476);
nor U80 (N_80,In_404,In_213);
or U81 (N_81,In_350,In_120);
and U82 (N_82,In_109,In_373);
or U83 (N_83,In_441,In_219);
and U84 (N_84,In_73,In_445);
xor U85 (N_85,In_301,In_335);
xor U86 (N_86,In_478,In_48);
and U87 (N_87,In_37,In_86);
and U88 (N_88,In_201,In_469);
or U89 (N_89,In_447,In_51);
nand U90 (N_90,In_244,In_234);
or U91 (N_91,In_135,In_456);
and U92 (N_92,In_71,In_79);
nor U93 (N_93,In_376,In_419);
nand U94 (N_94,In_362,In_88);
and U95 (N_95,In_443,In_410);
or U96 (N_96,In_62,In_418);
nor U97 (N_97,In_22,In_33);
or U98 (N_98,In_125,In_196);
nor U99 (N_99,In_66,In_124);
nor U100 (N_100,In_431,In_337);
and U101 (N_101,In_17,In_291);
and U102 (N_102,In_277,In_278);
nand U103 (N_103,In_123,In_492);
or U104 (N_104,In_81,In_231);
or U105 (N_105,In_163,In_220);
nor U106 (N_106,In_162,In_461);
nor U107 (N_107,In_96,In_269);
nor U108 (N_108,In_28,In_297);
nor U109 (N_109,In_409,In_358);
nor U110 (N_110,In_339,In_439);
and U111 (N_111,In_303,In_10);
or U112 (N_112,In_133,In_237);
nor U113 (N_113,In_104,In_364);
and U114 (N_114,In_14,In_154);
or U115 (N_115,In_369,In_477);
nand U116 (N_116,In_389,In_491);
nand U117 (N_117,In_170,In_417);
nand U118 (N_118,In_482,In_31);
or U119 (N_119,In_429,In_49);
nor U120 (N_120,In_343,In_388);
nor U121 (N_121,In_4,In_479);
nor U122 (N_122,In_473,In_412);
nor U123 (N_123,In_243,In_58);
and U124 (N_124,In_65,In_307);
and U125 (N_125,In_481,In_315);
nand U126 (N_126,In_166,In_11);
or U127 (N_127,In_20,In_428);
nand U128 (N_128,In_462,In_311);
or U129 (N_129,In_306,In_70);
nand U130 (N_130,In_424,In_490);
or U131 (N_131,In_30,In_132);
or U132 (N_132,In_108,In_103);
nand U133 (N_133,In_366,In_496);
or U134 (N_134,In_262,In_345);
nor U135 (N_135,In_294,In_330);
and U136 (N_136,In_384,In_45);
or U137 (N_137,In_401,In_352);
or U138 (N_138,In_266,In_187);
and U139 (N_139,In_450,In_489);
nor U140 (N_140,In_84,In_78);
or U141 (N_141,In_202,In_128);
or U142 (N_142,In_295,In_112);
nor U143 (N_143,In_16,In_322);
and U144 (N_144,In_194,In_224);
or U145 (N_145,In_457,In_293);
nand U146 (N_146,In_265,In_357);
nand U147 (N_147,In_238,In_263);
or U148 (N_148,In_396,In_391);
or U149 (N_149,In_47,In_276);
nand U150 (N_150,In_177,In_172);
nor U151 (N_151,In_344,In_129);
nand U152 (N_152,In_91,In_43);
nor U153 (N_153,In_206,In_304);
or U154 (N_154,In_211,In_18);
nor U155 (N_155,In_77,In_402);
and U156 (N_156,In_365,In_102);
and U157 (N_157,In_101,In_499);
nor U158 (N_158,In_233,In_209);
nor U159 (N_159,In_113,In_408);
and U160 (N_160,In_63,In_27);
and U161 (N_161,In_134,In_292);
and U162 (N_162,In_497,In_299);
and U163 (N_163,In_130,In_374);
nor U164 (N_164,In_59,In_385);
or U165 (N_165,In_155,In_216);
or U166 (N_166,In_480,In_420);
or U167 (N_167,In_368,In_185);
nand U168 (N_168,In_279,In_117);
or U169 (N_169,In_427,In_390);
nor U170 (N_170,In_251,In_387);
or U171 (N_171,In_212,In_310);
and U172 (N_172,In_2,In_226);
nand U173 (N_173,In_241,In_56);
and U174 (N_174,In_183,In_186);
or U175 (N_175,In_324,In_252);
nor U176 (N_176,In_23,In_235);
nand U177 (N_177,In_157,In_403);
and U178 (N_178,In_60,In_264);
nor U179 (N_179,In_398,In_35);
nor U180 (N_180,In_433,In_25);
or U181 (N_181,In_465,In_421);
or U182 (N_182,In_242,In_190);
nand U183 (N_183,In_44,In_495);
and U184 (N_184,In_40,In_331);
nand U185 (N_185,In_228,In_141);
and U186 (N_186,In_168,In_471);
and U187 (N_187,In_259,In_488);
or U188 (N_188,In_283,In_326);
or U189 (N_189,In_340,In_472);
or U190 (N_190,In_312,In_432);
or U191 (N_191,In_95,In_204);
nor U192 (N_192,In_466,In_328);
and U193 (N_193,In_195,In_289);
nand U194 (N_194,In_298,In_50);
and U195 (N_195,In_281,In_321);
or U196 (N_196,In_161,In_214);
and U197 (N_197,In_378,In_486);
or U198 (N_198,In_375,In_222);
or U199 (N_199,In_288,In_467);
nor U200 (N_200,N_122,In_203);
nand U201 (N_201,In_323,N_135);
nand U202 (N_202,N_0,N_186);
nor U203 (N_203,N_116,In_338);
nand U204 (N_204,N_86,N_156);
nand U205 (N_205,In_254,N_87);
nand U206 (N_206,N_74,In_75);
nor U207 (N_207,N_124,In_280);
or U208 (N_208,N_166,N_157);
and U209 (N_209,N_53,N_27);
and U210 (N_210,N_104,In_122);
and U211 (N_211,N_154,In_152);
and U212 (N_212,N_39,N_136);
nor U213 (N_213,In_173,N_181);
or U214 (N_214,N_89,N_118);
and U215 (N_215,N_127,N_20);
nand U216 (N_216,N_80,N_177);
and U217 (N_217,In_46,In_205);
nor U218 (N_218,N_131,N_54);
xnor U219 (N_219,N_32,In_327);
and U220 (N_220,In_118,In_12);
nor U221 (N_221,N_2,N_187);
or U222 (N_222,N_173,N_119);
and U223 (N_223,In_451,N_183);
and U224 (N_224,N_111,N_129);
nand U225 (N_225,In_184,In_142);
or U226 (N_226,In_197,N_160);
nor U227 (N_227,N_158,N_7);
and U228 (N_228,N_83,N_71);
nor U229 (N_229,In_407,N_78);
nand U230 (N_230,In_425,N_149);
and U231 (N_231,N_22,N_30);
nand U232 (N_232,N_42,N_29);
nand U233 (N_233,In_446,In_329);
nand U234 (N_234,N_151,In_320);
and U235 (N_235,N_199,N_60);
and U236 (N_236,In_215,N_196);
or U237 (N_237,In_336,N_81);
and U238 (N_238,N_55,N_28);
nor U239 (N_239,In_114,N_18);
or U240 (N_240,N_170,In_246);
or U241 (N_241,N_94,N_59);
or U242 (N_242,N_107,N_12);
and U243 (N_243,In_143,N_4);
nand U244 (N_244,N_178,N_148);
nand U245 (N_245,N_134,N_40);
and U246 (N_246,N_140,N_152);
xor U247 (N_247,In_138,N_95);
nand U248 (N_248,N_34,In_97);
nand U249 (N_249,N_146,In_41);
nand U250 (N_250,N_25,In_68);
nor U251 (N_251,N_26,N_184);
nor U252 (N_252,N_162,N_79);
or U253 (N_253,In_285,N_153);
or U254 (N_254,N_37,N_191);
and U255 (N_255,In_250,In_397);
nor U256 (N_256,N_75,In_87);
or U257 (N_257,N_137,N_68);
or U258 (N_258,N_142,N_144);
nor U259 (N_259,N_176,N_123);
nand U260 (N_260,In_69,N_96);
and U261 (N_261,In_53,In_148);
nor U262 (N_262,N_101,In_434);
or U263 (N_263,In_342,N_90);
xor U264 (N_264,In_156,In_498);
nand U265 (N_265,In_169,N_128);
xnor U266 (N_266,N_10,In_360);
nor U267 (N_267,N_47,In_363);
and U268 (N_268,In_260,N_24);
nor U269 (N_269,In_76,N_132);
or U270 (N_270,In_468,N_182);
nand U271 (N_271,In_52,N_161);
nand U272 (N_272,In_494,N_195);
nor U273 (N_273,N_38,N_169);
nor U274 (N_274,N_193,N_82);
nor U275 (N_275,N_159,In_383);
nand U276 (N_276,N_155,N_1);
or U277 (N_277,N_88,N_58);
nand U278 (N_278,N_6,In_164);
nand U279 (N_279,N_63,N_167);
nand U280 (N_280,N_130,In_199);
and U281 (N_281,N_50,N_125);
and U282 (N_282,N_197,In_393);
and U283 (N_283,N_106,N_175);
or U284 (N_284,N_57,N_150);
nand U285 (N_285,In_440,N_33);
or U286 (N_286,In_453,In_127);
nor U287 (N_287,N_121,In_470);
and U288 (N_288,N_43,N_51);
nor U289 (N_289,N_61,N_133);
nand U290 (N_290,N_102,In_406);
nor U291 (N_291,In_140,In_268);
and U292 (N_292,N_190,In_188);
nand U293 (N_293,In_160,In_422);
or U294 (N_294,In_208,In_464);
and U295 (N_295,In_150,N_91);
or U296 (N_296,N_41,N_49);
or U297 (N_297,N_147,N_15);
or U298 (N_298,N_76,N_143);
xor U299 (N_299,N_165,N_103);
nor U300 (N_300,N_114,N_21);
nand U301 (N_301,N_99,In_300);
nor U302 (N_302,N_84,In_415);
and U303 (N_303,N_31,N_110);
nand U304 (N_304,N_141,N_3);
and U305 (N_305,N_19,In_94);
nand U306 (N_306,In_236,N_16);
nor U307 (N_307,In_80,In_193);
or U308 (N_308,N_189,N_174);
xor U309 (N_309,N_70,N_9);
nor U310 (N_310,N_171,N_52);
and U311 (N_311,In_359,In_392);
nor U312 (N_312,In_382,In_435);
nor U313 (N_313,N_44,N_194);
or U314 (N_314,In_39,N_145);
nor U315 (N_315,N_72,In_317);
or U316 (N_316,N_85,N_69);
or U317 (N_317,N_93,In_475);
or U318 (N_318,N_168,N_100);
or U319 (N_319,N_179,N_115);
and U320 (N_320,In_116,N_164);
nor U321 (N_321,N_98,N_65);
and U322 (N_322,N_23,N_139);
nor U323 (N_323,In_153,In_115);
nor U324 (N_324,N_105,N_126);
nand U325 (N_325,N_180,N_109);
nor U326 (N_326,In_19,N_188);
or U327 (N_327,In_318,In_218);
nand U328 (N_328,In_379,N_113);
nand U329 (N_329,N_192,N_120);
nand U330 (N_330,In_274,In_399);
xor U331 (N_331,N_48,N_35);
or U332 (N_332,N_66,N_36);
nand U333 (N_333,In_341,N_62);
nor U334 (N_334,In_179,N_92);
or U335 (N_335,N_112,N_163);
or U336 (N_336,N_77,N_67);
nor U337 (N_337,N_73,N_108);
or U338 (N_338,N_8,N_172);
or U339 (N_339,In_55,N_56);
nor U340 (N_340,In_227,N_14);
nand U341 (N_341,N_117,N_138);
nand U342 (N_342,N_17,In_210);
and U343 (N_343,N_64,In_82);
nor U344 (N_344,N_198,N_46);
and U345 (N_345,In_181,In_5);
and U346 (N_346,N_5,N_185);
nor U347 (N_347,N_45,In_92);
nor U348 (N_348,N_13,N_11);
xnor U349 (N_349,N_97,In_126);
nor U350 (N_350,N_170,N_101);
nor U351 (N_351,N_40,In_82);
or U352 (N_352,N_152,N_26);
nor U353 (N_353,N_46,N_166);
and U354 (N_354,In_179,In_464);
or U355 (N_355,In_379,In_152);
nor U356 (N_356,In_434,In_116);
and U357 (N_357,In_393,N_93);
nand U358 (N_358,N_15,N_156);
nor U359 (N_359,In_246,N_42);
or U360 (N_360,N_199,N_104);
nand U361 (N_361,In_393,In_94);
and U362 (N_362,N_189,N_73);
and U363 (N_363,N_16,N_61);
nor U364 (N_364,In_150,N_40);
nand U365 (N_365,N_197,N_54);
or U366 (N_366,In_80,In_164);
nor U367 (N_367,N_159,N_151);
nand U368 (N_368,In_140,N_184);
and U369 (N_369,In_142,In_360);
and U370 (N_370,N_89,In_260);
nor U371 (N_371,N_55,In_327);
nor U372 (N_372,In_197,In_53);
nand U373 (N_373,In_199,N_117);
or U374 (N_374,N_92,In_336);
nor U375 (N_375,In_285,N_178);
nor U376 (N_376,N_197,N_93);
and U377 (N_377,N_43,N_155);
and U378 (N_378,N_168,N_88);
or U379 (N_379,N_62,N_153);
nand U380 (N_380,N_98,N_62);
nor U381 (N_381,N_94,N_196);
or U382 (N_382,N_22,N_128);
or U383 (N_383,N_11,In_140);
and U384 (N_384,N_36,N_126);
nor U385 (N_385,N_194,N_93);
and U386 (N_386,In_393,N_189);
or U387 (N_387,In_138,In_494);
nand U388 (N_388,N_51,N_1);
or U389 (N_389,N_174,In_68);
or U390 (N_390,N_0,In_494);
or U391 (N_391,N_57,N_172);
or U392 (N_392,N_79,N_193);
nor U393 (N_393,N_143,In_415);
nand U394 (N_394,N_55,N_64);
and U395 (N_395,N_35,In_300);
nand U396 (N_396,N_101,In_446);
or U397 (N_397,In_184,N_24);
or U398 (N_398,In_193,N_27);
or U399 (N_399,N_179,N_96);
and U400 (N_400,N_301,N_319);
or U401 (N_401,N_381,N_386);
nor U402 (N_402,N_318,N_244);
nand U403 (N_403,N_314,N_382);
nand U404 (N_404,N_368,N_294);
nor U405 (N_405,N_284,N_369);
or U406 (N_406,N_327,N_363);
or U407 (N_407,N_234,N_357);
or U408 (N_408,N_384,N_210);
or U409 (N_409,N_277,N_296);
and U410 (N_410,N_252,N_317);
and U411 (N_411,N_356,N_397);
or U412 (N_412,N_205,N_345);
and U413 (N_413,N_392,N_214);
or U414 (N_414,N_344,N_394);
or U415 (N_415,N_324,N_349);
xor U416 (N_416,N_312,N_337);
nor U417 (N_417,N_261,N_389);
and U418 (N_418,N_316,N_200);
nor U419 (N_419,N_377,N_219);
nand U420 (N_420,N_213,N_388);
and U421 (N_421,N_278,N_385);
nand U422 (N_422,N_379,N_291);
nand U423 (N_423,N_226,N_313);
nor U424 (N_424,N_343,N_355);
or U425 (N_425,N_209,N_242);
or U426 (N_426,N_342,N_285);
nand U427 (N_427,N_358,N_235);
nand U428 (N_428,N_274,N_309);
or U429 (N_429,N_231,N_326);
nand U430 (N_430,N_230,N_323);
nor U431 (N_431,N_256,N_346);
nand U432 (N_432,N_399,N_347);
or U433 (N_433,N_216,N_297);
and U434 (N_434,N_300,N_222);
nand U435 (N_435,N_262,N_287);
and U436 (N_436,N_330,N_283);
and U437 (N_437,N_246,N_359);
nand U438 (N_438,N_237,N_239);
nand U439 (N_439,N_281,N_221);
and U440 (N_440,N_223,N_304);
nand U441 (N_441,N_361,N_376);
and U442 (N_442,N_218,N_365);
or U443 (N_443,N_282,N_275);
or U444 (N_444,N_279,N_380);
nand U445 (N_445,N_383,N_206);
and U446 (N_446,N_259,N_390);
or U447 (N_447,N_302,N_398);
nor U448 (N_448,N_232,N_238);
or U449 (N_449,N_350,N_375);
nand U450 (N_450,N_354,N_241);
and U451 (N_451,N_311,N_236);
or U452 (N_452,N_243,N_331);
nand U453 (N_453,N_374,N_351);
nor U454 (N_454,N_270,N_321);
or U455 (N_455,N_245,N_362);
nand U456 (N_456,N_315,N_264);
nand U457 (N_457,N_307,N_254);
or U458 (N_458,N_322,N_266);
or U459 (N_459,N_233,N_260);
and U460 (N_460,N_208,N_265);
nand U461 (N_461,N_305,N_336);
or U462 (N_462,N_371,N_217);
nor U463 (N_463,N_303,N_255);
nor U464 (N_464,N_293,N_258);
and U465 (N_465,N_224,N_370);
nor U466 (N_466,N_396,N_373);
or U467 (N_467,N_268,N_250);
nand U468 (N_468,N_295,N_269);
or U469 (N_469,N_366,N_310);
nand U470 (N_470,N_338,N_247);
and U471 (N_471,N_202,N_360);
nand U472 (N_472,N_348,N_299);
nand U473 (N_473,N_267,N_280);
and U474 (N_474,N_378,N_335);
nor U475 (N_475,N_341,N_329);
and U476 (N_476,N_229,N_288);
nor U477 (N_477,N_340,N_290);
and U478 (N_478,N_228,N_271);
nand U479 (N_479,N_339,N_395);
nor U480 (N_480,N_325,N_276);
nand U481 (N_481,N_215,N_220);
nand U482 (N_482,N_328,N_263);
nand U483 (N_483,N_203,N_367);
nor U484 (N_484,N_251,N_306);
xor U485 (N_485,N_308,N_364);
or U486 (N_486,N_201,N_253);
nand U487 (N_487,N_353,N_249);
or U488 (N_488,N_289,N_204);
or U489 (N_489,N_248,N_372);
nand U490 (N_490,N_225,N_298);
nand U491 (N_491,N_240,N_393);
nand U492 (N_492,N_333,N_227);
nand U493 (N_493,N_211,N_391);
or U494 (N_494,N_286,N_212);
nand U495 (N_495,N_257,N_387);
or U496 (N_496,N_320,N_207);
or U497 (N_497,N_272,N_273);
or U498 (N_498,N_332,N_334);
nand U499 (N_499,N_292,N_352);
or U500 (N_500,N_239,N_258);
xor U501 (N_501,N_314,N_396);
nand U502 (N_502,N_340,N_394);
or U503 (N_503,N_391,N_282);
nand U504 (N_504,N_316,N_250);
or U505 (N_505,N_355,N_231);
and U506 (N_506,N_256,N_326);
nand U507 (N_507,N_388,N_225);
nand U508 (N_508,N_223,N_387);
or U509 (N_509,N_205,N_236);
nor U510 (N_510,N_356,N_296);
nor U511 (N_511,N_268,N_302);
or U512 (N_512,N_333,N_275);
nor U513 (N_513,N_352,N_394);
xor U514 (N_514,N_256,N_324);
nor U515 (N_515,N_332,N_276);
nand U516 (N_516,N_393,N_301);
nand U517 (N_517,N_321,N_311);
or U518 (N_518,N_231,N_255);
or U519 (N_519,N_221,N_291);
or U520 (N_520,N_366,N_200);
nand U521 (N_521,N_249,N_316);
and U522 (N_522,N_332,N_379);
or U523 (N_523,N_219,N_330);
or U524 (N_524,N_204,N_221);
nor U525 (N_525,N_387,N_275);
nor U526 (N_526,N_293,N_251);
nor U527 (N_527,N_222,N_281);
and U528 (N_528,N_372,N_357);
or U529 (N_529,N_259,N_269);
nand U530 (N_530,N_337,N_206);
nand U531 (N_531,N_358,N_203);
nand U532 (N_532,N_230,N_390);
or U533 (N_533,N_365,N_363);
or U534 (N_534,N_318,N_261);
or U535 (N_535,N_258,N_226);
or U536 (N_536,N_251,N_207);
and U537 (N_537,N_340,N_254);
nor U538 (N_538,N_208,N_219);
nor U539 (N_539,N_337,N_285);
and U540 (N_540,N_368,N_388);
and U541 (N_541,N_215,N_290);
nand U542 (N_542,N_274,N_292);
nor U543 (N_543,N_214,N_210);
or U544 (N_544,N_220,N_232);
nor U545 (N_545,N_289,N_365);
and U546 (N_546,N_324,N_370);
and U547 (N_547,N_334,N_267);
or U548 (N_548,N_339,N_347);
or U549 (N_549,N_282,N_263);
nor U550 (N_550,N_293,N_245);
and U551 (N_551,N_386,N_320);
nor U552 (N_552,N_346,N_259);
and U553 (N_553,N_371,N_385);
nor U554 (N_554,N_382,N_217);
or U555 (N_555,N_215,N_249);
xor U556 (N_556,N_212,N_377);
nor U557 (N_557,N_240,N_249);
xor U558 (N_558,N_293,N_377);
nor U559 (N_559,N_269,N_227);
nor U560 (N_560,N_317,N_209);
nand U561 (N_561,N_378,N_374);
nand U562 (N_562,N_225,N_268);
and U563 (N_563,N_201,N_374);
nor U564 (N_564,N_211,N_326);
and U565 (N_565,N_280,N_349);
or U566 (N_566,N_224,N_317);
nor U567 (N_567,N_215,N_361);
nor U568 (N_568,N_217,N_337);
nand U569 (N_569,N_399,N_238);
or U570 (N_570,N_346,N_348);
or U571 (N_571,N_223,N_294);
nand U572 (N_572,N_226,N_377);
or U573 (N_573,N_289,N_239);
nand U574 (N_574,N_273,N_245);
and U575 (N_575,N_208,N_325);
nand U576 (N_576,N_252,N_388);
nor U577 (N_577,N_337,N_341);
nor U578 (N_578,N_247,N_342);
or U579 (N_579,N_313,N_336);
nand U580 (N_580,N_388,N_245);
or U581 (N_581,N_377,N_274);
nor U582 (N_582,N_203,N_218);
or U583 (N_583,N_318,N_344);
or U584 (N_584,N_379,N_344);
nor U585 (N_585,N_391,N_265);
or U586 (N_586,N_384,N_322);
or U587 (N_587,N_346,N_293);
nand U588 (N_588,N_256,N_341);
and U589 (N_589,N_332,N_394);
nor U590 (N_590,N_356,N_232);
nand U591 (N_591,N_233,N_232);
or U592 (N_592,N_384,N_208);
and U593 (N_593,N_301,N_360);
nor U594 (N_594,N_291,N_372);
or U595 (N_595,N_282,N_336);
and U596 (N_596,N_318,N_222);
and U597 (N_597,N_221,N_283);
and U598 (N_598,N_311,N_271);
xor U599 (N_599,N_227,N_397);
nor U600 (N_600,N_423,N_566);
and U601 (N_601,N_574,N_426);
or U602 (N_602,N_444,N_494);
or U603 (N_603,N_583,N_416);
or U604 (N_604,N_593,N_596);
or U605 (N_605,N_403,N_565);
and U606 (N_606,N_471,N_517);
and U607 (N_607,N_487,N_475);
or U608 (N_608,N_548,N_409);
nand U609 (N_609,N_564,N_537);
nand U610 (N_610,N_479,N_459);
xor U611 (N_611,N_567,N_415);
xor U612 (N_612,N_577,N_482);
and U613 (N_613,N_441,N_552);
nor U614 (N_614,N_425,N_506);
and U615 (N_615,N_420,N_525);
or U616 (N_616,N_570,N_547);
nor U617 (N_617,N_568,N_429);
nand U618 (N_618,N_513,N_447);
or U619 (N_619,N_455,N_422);
and U620 (N_620,N_520,N_402);
nand U621 (N_621,N_435,N_448);
nand U622 (N_622,N_551,N_500);
nor U623 (N_623,N_523,N_438);
and U624 (N_624,N_432,N_401);
and U625 (N_625,N_497,N_539);
and U626 (N_626,N_554,N_524);
or U627 (N_627,N_427,N_412);
or U628 (N_628,N_549,N_417);
nor U629 (N_629,N_527,N_458);
nand U630 (N_630,N_421,N_498);
nand U631 (N_631,N_507,N_542);
or U632 (N_632,N_464,N_530);
or U633 (N_633,N_483,N_585);
nand U634 (N_634,N_499,N_405);
nand U635 (N_635,N_460,N_454);
or U636 (N_636,N_519,N_414);
and U637 (N_637,N_514,N_442);
and U638 (N_638,N_571,N_468);
or U639 (N_639,N_474,N_491);
nand U640 (N_640,N_408,N_543);
nor U641 (N_641,N_598,N_510);
or U642 (N_642,N_558,N_461);
nor U643 (N_643,N_451,N_436);
or U644 (N_644,N_440,N_489);
and U645 (N_645,N_594,N_550);
or U646 (N_646,N_439,N_457);
and U647 (N_647,N_450,N_452);
or U648 (N_648,N_545,N_467);
and U649 (N_649,N_518,N_469);
nand U650 (N_650,N_526,N_477);
nor U651 (N_651,N_555,N_553);
and U652 (N_652,N_472,N_466);
nand U653 (N_653,N_485,N_470);
or U654 (N_654,N_516,N_410);
nor U655 (N_655,N_509,N_540);
and U656 (N_656,N_488,N_493);
nor U657 (N_657,N_404,N_559);
nand U658 (N_658,N_434,N_572);
and U659 (N_659,N_591,N_541);
nand U660 (N_660,N_508,N_486);
nand U661 (N_661,N_465,N_587);
nand U662 (N_662,N_556,N_419);
or U663 (N_663,N_446,N_481);
and U664 (N_664,N_560,N_579);
nor U665 (N_665,N_411,N_580);
and U666 (N_666,N_430,N_531);
and U667 (N_667,N_589,N_437);
nand U668 (N_668,N_535,N_534);
and U669 (N_669,N_582,N_490);
or U670 (N_670,N_463,N_406);
or U671 (N_671,N_495,N_502);
nand U672 (N_672,N_561,N_590);
nand U673 (N_673,N_536,N_586);
or U674 (N_674,N_515,N_592);
and U675 (N_675,N_496,N_431);
nor U676 (N_676,N_599,N_473);
or U677 (N_677,N_588,N_400);
nor U678 (N_678,N_597,N_413);
and U679 (N_679,N_462,N_511);
or U680 (N_680,N_562,N_505);
and U681 (N_681,N_573,N_480);
nor U682 (N_682,N_428,N_546);
or U683 (N_683,N_522,N_501);
nor U684 (N_684,N_532,N_576);
nand U685 (N_685,N_484,N_504);
nand U686 (N_686,N_476,N_538);
nand U687 (N_687,N_529,N_544);
and U688 (N_688,N_563,N_528);
nor U689 (N_689,N_575,N_418);
nand U690 (N_690,N_424,N_581);
and U691 (N_691,N_584,N_456);
or U692 (N_692,N_503,N_512);
xnor U693 (N_693,N_445,N_407);
or U694 (N_694,N_533,N_443);
nand U695 (N_695,N_492,N_449);
nor U696 (N_696,N_578,N_521);
or U697 (N_697,N_569,N_453);
or U698 (N_698,N_433,N_478);
nor U699 (N_699,N_557,N_595);
nor U700 (N_700,N_515,N_434);
nand U701 (N_701,N_565,N_463);
and U702 (N_702,N_455,N_551);
nor U703 (N_703,N_598,N_533);
or U704 (N_704,N_540,N_557);
xor U705 (N_705,N_560,N_588);
nor U706 (N_706,N_599,N_565);
nand U707 (N_707,N_531,N_513);
and U708 (N_708,N_434,N_456);
nor U709 (N_709,N_597,N_451);
and U710 (N_710,N_489,N_505);
nor U711 (N_711,N_599,N_491);
or U712 (N_712,N_413,N_491);
or U713 (N_713,N_563,N_538);
or U714 (N_714,N_513,N_408);
nand U715 (N_715,N_531,N_479);
nand U716 (N_716,N_543,N_538);
or U717 (N_717,N_447,N_566);
xor U718 (N_718,N_438,N_472);
nor U719 (N_719,N_586,N_457);
and U720 (N_720,N_451,N_412);
and U721 (N_721,N_577,N_541);
nor U722 (N_722,N_570,N_443);
or U723 (N_723,N_580,N_532);
and U724 (N_724,N_444,N_411);
or U725 (N_725,N_554,N_455);
nor U726 (N_726,N_503,N_447);
nand U727 (N_727,N_529,N_582);
and U728 (N_728,N_447,N_451);
xnor U729 (N_729,N_515,N_425);
nor U730 (N_730,N_401,N_530);
or U731 (N_731,N_563,N_527);
and U732 (N_732,N_546,N_416);
or U733 (N_733,N_595,N_456);
and U734 (N_734,N_470,N_529);
nand U735 (N_735,N_486,N_401);
and U736 (N_736,N_435,N_577);
and U737 (N_737,N_407,N_521);
xor U738 (N_738,N_532,N_575);
nand U739 (N_739,N_592,N_496);
or U740 (N_740,N_449,N_537);
nand U741 (N_741,N_520,N_575);
xor U742 (N_742,N_598,N_438);
or U743 (N_743,N_449,N_559);
nor U744 (N_744,N_502,N_546);
nand U745 (N_745,N_425,N_568);
nand U746 (N_746,N_403,N_471);
nor U747 (N_747,N_525,N_475);
nor U748 (N_748,N_594,N_433);
and U749 (N_749,N_528,N_403);
or U750 (N_750,N_550,N_575);
nor U751 (N_751,N_415,N_581);
nor U752 (N_752,N_416,N_451);
and U753 (N_753,N_582,N_522);
or U754 (N_754,N_431,N_419);
or U755 (N_755,N_532,N_595);
and U756 (N_756,N_474,N_486);
and U757 (N_757,N_411,N_433);
nand U758 (N_758,N_532,N_452);
nor U759 (N_759,N_505,N_581);
nand U760 (N_760,N_530,N_433);
nand U761 (N_761,N_554,N_553);
nand U762 (N_762,N_401,N_543);
or U763 (N_763,N_494,N_504);
nand U764 (N_764,N_532,N_485);
and U765 (N_765,N_483,N_501);
nor U766 (N_766,N_490,N_554);
and U767 (N_767,N_590,N_433);
or U768 (N_768,N_511,N_492);
or U769 (N_769,N_473,N_524);
or U770 (N_770,N_589,N_517);
and U771 (N_771,N_588,N_415);
nor U772 (N_772,N_595,N_517);
nor U773 (N_773,N_568,N_574);
and U774 (N_774,N_547,N_529);
and U775 (N_775,N_400,N_563);
and U776 (N_776,N_527,N_474);
nor U777 (N_777,N_532,N_436);
nand U778 (N_778,N_436,N_519);
and U779 (N_779,N_442,N_438);
and U780 (N_780,N_411,N_565);
nand U781 (N_781,N_573,N_533);
or U782 (N_782,N_577,N_507);
and U783 (N_783,N_541,N_472);
and U784 (N_784,N_529,N_591);
nand U785 (N_785,N_449,N_574);
nand U786 (N_786,N_557,N_524);
and U787 (N_787,N_497,N_412);
nor U788 (N_788,N_457,N_469);
and U789 (N_789,N_485,N_428);
and U790 (N_790,N_485,N_446);
or U791 (N_791,N_510,N_434);
nand U792 (N_792,N_504,N_562);
nor U793 (N_793,N_468,N_561);
nor U794 (N_794,N_539,N_512);
xnor U795 (N_795,N_464,N_501);
and U796 (N_796,N_509,N_446);
and U797 (N_797,N_477,N_537);
nor U798 (N_798,N_537,N_515);
and U799 (N_799,N_502,N_444);
and U800 (N_800,N_636,N_704);
and U801 (N_801,N_608,N_770);
and U802 (N_802,N_671,N_615);
or U803 (N_803,N_769,N_668);
and U804 (N_804,N_765,N_652);
nor U805 (N_805,N_749,N_600);
and U806 (N_806,N_681,N_620);
xor U807 (N_807,N_662,N_670);
or U808 (N_808,N_734,N_754);
nand U809 (N_809,N_611,N_758);
xnor U810 (N_810,N_763,N_747);
and U811 (N_811,N_742,N_716);
and U812 (N_812,N_773,N_762);
nand U813 (N_813,N_721,N_759);
nand U814 (N_814,N_774,N_691);
or U815 (N_815,N_743,N_703);
nor U816 (N_816,N_603,N_637);
and U817 (N_817,N_630,N_635);
and U818 (N_818,N_722,N_659);
nand U819 (N_819,N_641,N_776);
xnor U820 (N_820,N_651,N_669);
or U821 (N_821,N_791,N_673);
nor U822 (N_822,N_656,N_667);
or U823 (N_823,N_727,N_702);
nor U824 (N_824,N_610,N_753);
and U825 (N_825,N_755,N_751);
nand U826 (N_826,N_606,N_725);
nand U827 (N_827,N_764,N_729);
nand U828 (N_828,N_746,N_686);
and U829 (N_829,N_674,N_728);
nand U830 (N_830,N_665,N_739);
nor U831 (N_831,N_797,N_694);
nor U832 (N_832,N_622,N_616);
and U833 (N_833,N_719,N_609);
nand U834 (N_834,N_771,N_666);
nor U835 (N_835,N_617,N_766);
nor U836 (N_836,N_643,N_650);
or U837 (N_837,N_798,N_661);
or U838 (N_838,N_654,N_752);
xnor U839 (N_839,N_607,N_711);
or U840 (N_840,N_738,N_647);
nor U841 (N_841,N_736,N_642);
nand U842 (N_842,N_788,N_660);
nand U843 (N_843,N_783,N_612);
or U844 (N_844,N_779,N_624);
nand U845 (N_845,N_602,N_680);
or U846 (N_846,N_757,N_794);
and U847 (N_847,N_677,N_623);
or U848 (N_848,N_784,N_732);
nor U849 (N_849,N_740,N_750);
nor U850 (N_850,N_799,N_693);
nor U851 (N_851,N_699,N_678);
and U852 (N_852,N_741,N_782);
nand U853 (N_853,N_731,N_634);
xor U854 (N_854,N_787,N_767);
nor U855 (N_855,N_785,N_649);
and U856 (N_856,N_655,N_723);
or U857 (N_857,N_631,N_772);
nor U858 (N_858,N_724,N_684);
nor U859 (N_859,N_789,N_717);
nand U860 (N_860,N_627,N_688);
nand U861 (N_861,N_628,N_715);
nand U862 (N_862,N_676,N_626);
and U863 (N_863,N_712,N_683);
nand U864 (N_864,N_735,N_679);
and U865 (N_865,N_639,N_605);
nand U866 (N_866,N_710,N_658);
nand U867 (N_867,N_707,N_705);
nand U868 (N_868,N_760,N_685);
and U869 (N_869,N_644,N_761);
nor U870 (N_870,N_768,N_672);
or U871 (N_871,N_730,N_720);
nand U872 (N_872,N_718,N_653);
nor U873 (N_873,N_698,N_675);
nand U874 (N_874,N_621,N_786);
nand U875 (N_875,N_795,N_638);
nand U876 (N_876,N_695,N_777);
nor U877 (N_877,N_682,N_790);
nor U878 (N_878,N_687,N_633);
and U879 (N_879,N_714,N_706);
or U880 (N_880,N_756,N_780);
or U881 (N_881,N_778,N_733);
or U882 (N_882,N_657,N_796);
nand U883 (N_883,N_744,N_726);
or U884 (N_884,N_793,N_745);
nor U885 (N_885,N_625,N_775);
and U886 (N_886,N_646,N_664);
and U887 (N_887,N_748,N_700);
or U888 (N_888,N_697,N_708);
nand U889 (N_889,N_696,N_601);
and U890 (N_890,N_640,N_701);
and U891 (N_891,N_781,N_648);
nor U892 (N_892,N_629,N_692);
and U893 (N_893,N_614,N_604);
and U894 (N_894,N_713,N_619);
and U895 (N_895,N_613,N_689);
or U896 (N_896,N_709,N_663);
nor U897 (N_897,N_632,N_737);
or U898 (N_898,N_645,N_792);
nor U899 (N_899,N_690,N_618);
or U900 (N_900,N_684,N_600);
or U901 (N_901,N_769,N_611);
and U902 (N_902,N_602,N_638);
or U903 (N_903,N_687,N_694);
nor U904 (N_904,N_698,N_641);
and U905 (N_905,N_667,N_668);
and U906 (N_906,N_736,N_718);
nand U907 (N_907,N_621,N_758);
nand U908 (N_908,N_708,N_695);
or U909 (N_909,N_792,N_753);
nor U910 (N_910,N_765,N_711);
nand U911 (N_911,N_612,N_785);
nor U912 (N_912,N_774,N_603);
and U913 (N_913,N_756,N_644);
xor U914 (N_914,N_690,N_700);
nor U915 (N_915,N_715,N_799);
nor U916 (N_916,N_733,N_609);
nand U917 (N_917,N_743,N_759);
nor U918 (N_918,N_697,N_670);
nor U919 (N_919,N_789,N_655);
or U920 (N_920,N_694,N_715);
and U921 (N_921,N_792,N_658);
nand U922 (N_922,N_683,N_659);
nand U923 (N_923,N_683,N_684);
or U924 (N_924,N_766,N_753);
and U925 (N_925,N_706,N_690);
nor U926 (N_926,N_697,N_620);
nor U927 (N_927,N_630,N_790);
or U928 (N_928,N_646,N_794);
or U929 (N_929,N_796,N_778);
and U930 (N_930,N_678,N_666);
or U931 (N_931,N_744,N_735);
nor U932 (N_932,N_794,N_612);
nand U933 (N_933,N_606,N_774);
nor U934 (N_934,N_788,N_696);
and U935 (N_935,N_747,N_694);
and U936 (N_936,N_669,N_785);
or U937 (N_937,N_625,N_751);
or U938 (N_938,N_745,N_640);
nor U939 (N_939,N_640,N_686);
nor U940 (N_940,N_791,N_665);
or U941 (N_941,N_647,N_792);
nand U942 (N_942,N_604,N_685);
nand U943 (N_943,N_619,N_641);
and U944 (N_944,N_618,N_702);
nor U945 (N_945,N_635,N_601);
nand U946 (N_946,N_792,N_643);
and U947 (N_947,N_645,N_674);
and U948 (N_948,N_718,N_707);
and U949 (N_949,N_794,N_728);
nor U950 (N_950,N_734,N_622);
or U951 (N_951,N_600,N_746);
or U952 (N_952,N_709,N_700);
and U953 (N_953,N_740,N_658);
or U954 (N_954,N_706,N_735);
and U955 (N_955,N_785,N_747);
or U956 (N_956,N_790,N_783);
or U957 (N_957,N_772,N_798);
nand U958 (N_958,N_793,N_621);
nor U959 (N_959,N_726,N_762);
nor U960 (N_960,N_711,N_696);
nor U961 (N_961,N_793,N_789);
and U962 (N_962,N_612,N_755);
or U963 (N_963,N_607,N_625);
or U964 (N_964,N_799,N_636);
nor U965 (N_965,N_790,N_672);
xor U966 (N_966,N_639,N_738);
or U967 (N_967,N_710,N_793);
and U968 (N_968,N_669,N_653);
or U969 (N_969,N_718,N_791);
and U970 (N_970,N_781,N_763);
nand U971 (N_971,N_691,N_720);
nand U972 (N_972,N_776,N_655);
and U973 (N_973,N_775,N_688);
and U974 (N_974,N_721,N_772);
or U975 (N_975,N_640,N_622);
nand U976 (N_976,N_687,N_624);
or U977 (N_977,N_771,N_685);
nor U978 (N_978,N_617,N_792);
and U979 (N_979,N_625,N_628);
and U980 (N_980,N_719,N_657);
nor U981 (N_981,N_622,N_672);
or U982 (N_982,N_742,N_799);
nand U983 (N_983,N_680,N_702);
or U984 (N_984,N_753,N_623);
nor U985 (N_985,N_633,N_762);
or U986 (N_986,N_614,N_709);
nand U987 (N_987,N_691,N_613);
and U988 (N_988,N_664,N_654);
or U989 (N_989,N_762,N_614);
and U990 (N_990,N_694,N_643);
nor U991 (N_991,N_689,N_701);
nand U992 (N_992,N_602,N_716);
nor U993 (N_993,N_663,N_698);
and U994 (N_994,N_773,N_724);
nand U995 (N_995,N_751,N_785);
nand U996 (N_996,N_737,N_788);
nand U997 (N_997,N_704,N_624);
nand U998 (N_998,N_627,N_764);
nand U999 (N_999,N_764,N_780);
or U1000 (N_1000,N_897,N_823);
nor U1001 (N_1001,N_955,N_814);
and U1002 (N_1002,N_883,N_925);
nor U1003 (N_1003,N_998,N_937);
and U1004 (N_1004,N_900,N_870);
nand U1005 (N_1005,N_833,N_856);
nand U1006 (N_1006,N_996,N_887);
nor U1007 (N_1007,N_827,N_974);
nor U1008 (N_1008,N_958,N_946);
nand U1009 (N_1009,N_986,N_939);
nor U1010 (N_1010,N_993,N_934);
nand U1011 (N_1011,N_959,N_818);
nor U1012 (N_1012,N_926,N_964);
or U1013 (N_1013,N_953,N_961);
nand U1014 (N_1014,N_947,N_901);
or U1015 (N_1015,N_973,N_891);
or U1016 (N_1016,N_991,N_999);
nor U1017 (N_1017,N_917,N_932);
nor U1018 (N_1018,N_997,N_889);
or U1019 (N_1019,N_976,N_944);
nand U1020 (N_1020,N_984,N_878);
or U1021 (N_1021,N_832,N_863);
and U1022 (N_1022,N_988,N_815);
nor U1023 (N_1023,N_972,N_910);
or U1024 (N_1024,N_916,N_924);
nor U1025 (N_1025,N_969,N_855);
and U1026 (N_1026,N_884,N_864);
nor U1027 (N_1027,N_828,N_850);
nand U1028 (N_1028,N_963,N_957);
or U1029 (N_1029,N_888,N_948);
nor U1030 (N_1030,N_979,N_949);
and U1031 (N_1031,N_848,N_844);
nand U1032 (N_1032,N_985,N_980);
nand U1033 (N_1033,N_825,N_820);
nor U1034 (N_1034,N_904,N_920);
xor U1035 (N_1035,N_954,N_835);
nor U1036 (N_1036,N_995,N_822);
and U1037 (N_1037,N_908,N_803);
or U1038 (N_1038,N_852,N_970);
nor U1039 (N_1039,N_853,N_837);
nor U1040 (N_1040,N_893,N_866);
and U1041 (N_1041,N_869,N_951);
and U1042 (N_1042,N_895,N_811);
and U1043 (N_1043,N_965,N_862);
xnor U1044 (N_1044,N_872,N_927);
and U1045 (N_1045,N_914,N_840);
xor U1046 (N_1046,N_978,N_923);
nor U1047 (N_1047,N_843,N_868);
nor U1048 (N_1048,N_831,N_921);
and U1049 (N_1049,N_817,N_890);
and U1050 (N_1050,N_807,N_865);
nand U1051 (N_1051,N_860,N_896);
or U1052 (N_1052,N_819,N_829);
nand U1053 (N_1053,N_956,N_968);
nand U1054 (N_1054,N_892,N_847);
and U1055 (N_1055,N_874,N_804);
and U1056 (N_1056,N_805,N_810);
nor U1057 (N_1057,N_881,N_812);
or U1058 (N_1058,N_922,N_845);
and U1059 (N_1059,N_919,N_909);
nand U1060 (N_1060,N_824,N_857);
xnor U1061 (N_1061,N_928,N_800);
or U1062 (N_1062,N_841,N_912);
nand U1063 (N_1063,N_861,N_858);
or U1064 (N_1064,N_834,N_894);
or U1065 (N_1065,N_816,N_941);
and U1066 (N_1066,N_898,N_838);
and U1067 (N_1067,N_938,N_880);
nand U1068 (N_1068,N_885,N_981);
nand U1069 (N_1069,N_802,N_966);
or U1070 (N_1070,N_907,N_940);
xnor U1071 (N_1071,N_906,N_992);
nand U1072 (N_1072,N_877,N_905);
and U1073 (N_1073,N_902,N_915);
and U1074 (N_1074,N_911,N_846);
nor U1075 (N_1075,N_886,N_839);
nor U1076 (N_1076,N_950,N_967);
and U1077 (N_1077,N_930,N_842);
and U1078 (N_1078,N_962,N_935);
or U1079 (N_1079,N_806,N_867);
nor U1080 (N_1080,N_903,N_849);
and U1081 (N_1081,N_994,N_808);
nor U1082 (N_1082,N_990,N_971);
nand U1083 (N_1083,N_977,N_813);
and U1084 (N_1084,N_960,N_826);
nand U1085 (N_1085,N_918,N_821);
xor U1086 (N_1086,N_879,N_836);
nand U1087 (N_1087,N_871,N_929);
nor U1088 (N_1088,N_943,N_933);
and U1089 (N_1089,N_876,N_952);
xnor U1090 (N_1090,N_851,N_854);
xnor U1091 (N_1091,N_899,N_945);
nand U1092 (N_1092,N_830,N_875);
nor U1093 (N_1093,N_913,N_982);
nor U1094 (N_1094,N_989,N_859);
and U1095 (N_1095,N_873,N_987);
and U1096 (N_1096,N_983,N_882);
nand U1097 (N_1097,N_801,N_931);
nor U1098 (N_1098,N_942,N_936);
nor U1099 (N_1099,N_975,N_809);
nand U1100 (N_1100,N_917,N_955);
and U1101 (N_1101,N_976,N_954);
nor U1102 (N_1102,N_823,N_806);
nand U1103 (N_1103,N_932,N_888);
or U1104 (N_1104,N_997,N_818);
and U1105 (N_1105,N_869,N_825);
nor U1106 (N_1106,N_930,N_952);
and U1107 (N_1107,N_969,N_902);
nand U1108 (N_1108,N_986,N_979);
nand U1109 (N_1109,N_893,N_947);
nor U1110 (N_1110,N_954,N_881);
or U1111 (N_1111,N_823,N_876);
nor U1112 (N_1112,N_834,N_807);
and U1113 (N_1113,N_973,N_919);
nor U1114 (N_1114,N_836,N_859);
nand U1115 (N_1115,N_844,N_896);
and U1116 (N_1116,N_999,N_917);
nor U1117 (N_1117,N_924,N_951);
nand U1118 (N_1118,N_896,N_980);
nand U1119 (N_1119,N_804,N_826);
nand U1120 (N_1120,N_954,N_879);
nor U1121 (N_1121,N_863,N_857);
and U1122 (N_1122,N_977,N_825);
or U1123 (N_1123,N_897,N_810);
or U1124 (N_1124,N_818,N_897);
or U1125 (N_1125,N_995,N_852);
and U1126 (N_1126,N_943,N_903);
nor U1127 (N_1127,N_902,N_884);
nor U1128 (N_1128,N_938,N_883);
nand U1129 (N_1129,N_817,N_880);
or U1130 (N_1130,N_936,N_976);
nor U1131 (N_1131,N_839,N_882);
nor U1132 (N_1132,N_880,N_892);
nor U1133 (N_1133,N_940,N_830);
nand U1134 (N_1134,N_823,N_830);
and U1135 (N_1135,N_950,N_915);
and U1136 (N_1136,N_873,N_942);
and U1137 (N_1137,N_917,N_830);
nand U1138 (N_1138,N_944,N_942);
nor U1139 (N_1139,N_894,N_985);
nand U1140 (N_1140,N_953,N_972);
nand U1141 (N_1141,N_965,N_988);
and U1142 (N_1142,N_822,N_936);
nor U1143 (N_1143,N_921,N_987);
nor U1144 (N_1144,N_887,N_874);
nor U1145 (N_1145,N_819,N_814);
or U1146 (N_1146,N_833,N_887);
nand U1147 (N_1147,N_961,N_985);
or U1148 (N_1148,N_950,N_988);
and U1149 (N_1149,N_814,N_826);
nor U1150 (N_1150,N_888,N_937);
and U1151 (N_1151,N_945,N_966);
and U1152 (N_1152,N_930,N_826);
or U1153 (N_1153,N_809,N_816);
nor U1154 (N_1154,N_824,N_921);
nand U1155 (N_1155,N_956,N_835);
or U1156 (N_1156,N_891,N_981);
and U1157 (N_1157,N_819,N_928);
or U1158 (N_1158,N_854,N_852);
and U1159 (N_1159,N_804,N_967);
or U1160 (N_1160,N_813,N_810);
or U1161 (N_1161,N_919,N_888);
nand U1162 (N_1162,N_847,N_968);
or U1163 (N_1163,N_878,N_945);
or U1164 (N_1164,N_833,N_847);
or U1165 (N_1165,N_868,N_947);
or U1166 (N_1166,N_984,N_859);
xor U1167 (N_1167,N_924,N_913);
xor U1168 (N_1168,N_876,N_973);
nand U1169 (N_1169,N_820,N_902);
nor U1170 (N_1170,N_854,N_972);
nand U1171 (N_1171,N_874,N_997);
nor U1172 (N_1172,N_847,N_922);
and U1173 (N_1173,N_878,N_851);
and U1174 (N_1174,N_923,N_908);
and U1175 (N_1175,N_864,N_942);
and U1176 (N_1176,N_833,N_843);
nor U1177 (N_1177,N_974,N_828);
nand U1178 (N_1178,N_817,N_911);
nand U1179 (N_1179,N_820,N_812);
or U1180 (N_1180,N_931,N_840);
or U1181 (N_1181,N_885,N_989);
and U1182 (N_1182,N_992,N_937);
nor U1183 (N_1183,N_897,N_841);
nand U1184 (N_1184,N_925,N_975);
or U1185 (N_1185,N_970,N_883);
nand U1186 (N_1186,N_966,N_990);
or U1187 (N_1187,N_858,N_854);
nand U1188 (N_1188,N_943,N_845);
and U1189 (N_1189,N_855,N_925);
nand U1190 (N_1190,N_802,N_821);
nand U1191 (N_1191,N_819,N_890);
nor U1192 (N_1192,N_884,N_847);
nor U1193 (N_1193,N_879,N_887);
nand U1194 (N_1194,N_962,N_837);
or U1195 (N_1195,N_941,N_994);
nor U1196 (N_1196,N_908,N_828);
or U1197 (N_1197,N_980,N_874);
and U1198 (N_1198,N_877,N_894);
nand U1199 (N_1199,N_978,N_828);
nand U1200 (N_1200,N_1013,N_1104);
or U1201 (N_1201,N_1139,N_1182);
nand U1202 (N_1202,N_1006,N_1144);
and U1203 (N_1203,N_1045,N_1059);
or U1204 (N_1204,N_1030,N_1170);
or U1205 (N_1205,N_1143,N_1153);
nor U1206 (N_1206,N_1075,N_1055);
nand U1207 (N_1207,N_1057,N_1109);
nand U1208 (N_1208,N_1178,N_1088);
nand U1209 (N_1209,N_1014,N_1051);
nor U1210 (N_1210,N_1085,N_1167);
and U1211 (N_1211,N_1081,N_1184);
nand U1212 (N_1212,N_1133,N_1046);
nor U1213 (N_1213,N_1192,N_1146);
or U1214 (N_1214,N_1107,N_1117);
or U1215 (N_1215,N_1127,N_1084);
nand U1216 (N_1216,N_1163,N_1063);
and U1217 (N_1217,N_1062,N_1187);
and U1218 (N_1218,N_1004,N_1173);
nor U1219 (N_1219,N_1154,N_1066);
or U1220 (N_1220,N_1042,N_1124);
nor U1221 (N_1221,N_1003,N_1070);
nor U1222 (N_1222,N_1102,N_1140);
and U1223 (N_1223,N_1198,N_1002);
xor U1224 (N_1224,N_1098,N_1017);
or U1225 (N_1225,N_1005,N_1018);
nor U1226 (N_1226,N_1141,N_1190);
or U1227 (N_1227,N_1068,N_1039);
and U1228 (N_1228,N_1194,N_1118);
nor U1229 (N_1229,N_1099,N_1001);
or U1230 (N_1230,N_1089,N_1067);
or U1231 (N_1231,N_1058,N_1023);
nand U1232 (N_1232,N_1056,N_1082);
nand U1233 (N_1233,N_1080,N_1019);
nand U1234 (N_1234,N_1155,N_1032);
nand U1235 (N_1235,N_1129,N_1158);
nand U1236 (N_1236,N_1061,N_1120);
nand U1237 (N_1237,N_1071,N_1083);
and U1238 (N_1238,N_1064,N_1165);
or U1239 (N_1239,N_1161,N_1175);
xor U1240 (N_1240,N_1103,N_1016);
nor U1241 (N_1241,N_1091,N_1131);
nand U1242 (N_1242,N_1149,N_1072);
nand U1243 (N_1243,N_1180,N_1028);
and U1244 (N_1244,N_1162,N_1021);
or U1245 (N_1245,N_1087,N_1150);
and U1246 (N_1246,N_1047,N_1108);
nor U1247 (N_1247,N_1199,N_1112);
nor U1248 (N_1248,N_1037,N_1186);
or U1249 (N_1249,N_1196,N_1106);
or U1250 (N_1250,N_1034,N_1052);
or U1251 (N_1251,N_1024,N_1137);
or U1252 (N_1252,N_1145,N_1012);
nor U1253 (N_1253,N_1113,N_1027);
and U1254 (N_1254,N_1132,N_1025);
or U1255 (N_1255,N_1044,N_1147);
nand U1256 (N_1256,N_1151,N_1176);
and U1257 (N_1257,N_1060,N_1130);
or U1258 (N_1258,N_1135,N_1086);
or U1259 (N_1259,N_1166,N_1040);
or U1260 (N_1260,N_1188,N_1156);
nor U1261 (N_1261,N_1122,N_1048);
nand U1262 (N_1262,N_1093,N_1090);
nor U1263 (N_1263,N_1185,N_1134);
or U1264 (N_1264,N_1008,N_1157);
nand U1265 (N_1265,N_1035,N_1121);
nor U1266 (N_1266,N_1193,N_1010);
nor U1267 (N_1267,N_1111,N_1043);
and U1268 (N_1268,N_1073,N_1177);
or U1269 (N_1269,N_1011,N_1142);
nand U1270 (N_1270,N_1100,N_1119);
nand U1271 (N_1271,N_1179,N_1096);
nor U1272 (N_1272,N_1065,N_1054);
xor U1273 (N_1273,N_1022,N_1172);
and U1274 (N_1274,N_1123,N_1097);
nand U1275 (N_1275,N_1015,N_1164);
and U1276 (N_1276,N_1049,N_1069);
or U1277 (N_1277,N_1079,N_1115);
or U1278 (N_1278,N_1041,N_1191);
nor U1279 (N_1279,N_1076,N_1078);
and U1280 (N_1280,N_1136,N_1077);
nor U1281 (N_1281,N_1092,N_1053);
or U1282 (N_1282,N_1171,N_1029);
and U1283 (N_1283,N_1095,N_1101);
and U1284 (N_1284,N_1009,N_1183);
or U1285 (N_1285,N_1195,N_1125);
nand U1286 (N_1286,N_1074,N_1110);
nand U1287 (N_1287,N_1174,N_1038);
nor U1288 (N_1288,N_1007,N_1189);
nor U1289 (N_1289,N_1128,N_1159);
and U1290 (N_1290,N_1105,N_1169);
nand U1291 (N_1291,N_1116,N_1148);
nor U1292 (N_1292,N_1152,N_1138);
nor U1293 (N_1293,N_1197,N_1000);
and U1294 (N_1294,N_1026,N_1094);
and U1295 (N_1295,N_1031,N_1126);
nor U1296 (N_1296,N_1114,N_1036);
xnor U1297 (N_1297,N_1181,N_1020);
or U1298 (N_1298,N_1168,N_1033);
nand U1299 (N_1299,N_1160,N_1050);
and U1300 (N_1300,N_1121,N_1137);
and U1301 (N_1301,N_1100,N_1147);
xnor U1302 (N_1302,N_1055,N_1116);
xnor U1303 (N_1303,N_1044,N_1133);
nor U1304 (N_1304,N_1024,N_1119);
nor U1305 (N_1305,N_1008,N_1089);
or U1306 (N_1306,N_1186,N_1038);
nor U1307 (N_1307,N_1057,N_1105);
and U1308 (N_1308,N_1041,N_1049);
and U1309 (N_1309,N_1029,N_1176);
nor U1310 (N_1310,N_1105,N_1076);
nand U1311 (N_1311,N_1018,N_1045);
or U1312 (N_1312,N_1130,N_1099);
and U1313 (N_1313,N_1107,N_1110);
nor U1314 (N_1314,N_1195,N_1189);
nor U1315 (N_1315,N_1093,N_1188);
nand U1316 (N_1316,N_1086,N_1133);
nor U1317 (N_1317,N_1165,N_1060);
or U1318 (N_1318,N_1108,N_1130);
and U1319 (N_1319,N_1152,N_1035);
or U1320 (N_1320,N_1118,N_1137);
nand U1321 (N_1321,N_1001,N_1115);
xor U1322 (N_1322,N_1126,N_1102);
and U1323 (N_1323,N_1007,N_1191);
nand U1324 (N_1324,N_1075,N_1043);
and U1325 (N_1325,N_1071,N_1027);
or U1326 (N_1326,N_1059,N_1077);
or U1327 (N_1327,N_1113,N_1065);
or U1328 (N_1328,N_1042,N_1062);
and U1329 (N_1329,N_1073,N_1149);
and U1330 (N_1330,N_1199,N_1000);
nor U1331 (N_1331,N_1132,N_1092);
nor U1332 (N_1332,N_1134,N_1199);
nand U1333 (N_1333,N_1064,N_1193);
and U1334 (N_1334,N_1005,N_1078);
nand U1335 (N_1335,N_1127,N_1131);
nor U1336 (N_1336,N_1166,N_1030);
or U1337 (N_1337,N_1068,N_1143);
or U1338 (N_1338,N_1174,N_1031);
nand U1339 (N_1339,N_1140,N_1054);
or U1340 (N_1340,N_1159,N_1108);
and U1341 (N_1341,N_1159,N_1019);
or U1342 (N_1342,N_1085,N_1130);
nor U1343 (N_1343,N_1158,N_1143);
nor U1344 (N_1344,N_1105,N_1107);
nand U1345 (N_1345,N_1158,N_1002);
and U1346 (N_1346,N_1005,N_1115);
and U1347 (N_1347,N_1075,N_1184);
and U1348 (N_1348,N_1170,N_1049);
nor U1349 (N_1349,N_1071,N_1161);
nand U1350 (N_1350,N_1073,N_1170);
nor U1351 (N_1351,N_1172,N_1167);
nor U1352 (N_1352,N_1176,N_1025);
or U1353 (N_1353,N_1176,N_1079);
nor U1354 (N_1354,N_1066,N_1006);
and U1355 (N_1355,N_1153,N_1116);
and U1356 (N_1356,N_1071,N_1157);
nor U1357 (N_1357,N_1058,N_1042);
xnor U1358 (N_1358,N_1095,N_1020);
nand U1359 (N_1359,N_1001,N_1018);
or U1360 (N_1360,N_1035,N_1180);
or U1361 (N_1361,N_1106,N_1195);
nor U1362 (N_1362,N_1057,N_1072);
nor U1363 (N_1363,N_1096,N_1065);
nand U1364 (N_1364,N_1013,N_1158);
and U1365 (N_1365,N_1038,N_1049);
nand U1366 (N_1366,N_1193,N_1030);
and U1367 (N_1367,N_1113,N_1104);
or U1368 (N_1368,N_1187,N_1126);
nand U1369 (N_1369,N_1175,N_1087);
and U1370 (N_1370,N_1189,N_1056);
nand U1371 (N_1371,N_1039,N_1124);
nor U1372 (N_1372,N_1097,N_1048);
or U1373 (N_1373,N_1108,N_1001);
and U1374 (N_1374,N_1086,N_1180);
or U1375 (N_1375,N_1078,N_1108);
or U1376 (N_1376,N_1184,N_1069);
and U1377 (N_1377,N_1172,N_1139);
and U1378 (N_1378,N_1135,N_1072);
or U1379 (N_1379,N_1095,N_1047);
or U1380 (N_1380,N_1028,N_1085);
nor U1381 (N_1381,N_1042,N_1057);
xor U1382 (N_1382,N_1072,N_1171);
nor U1383 (N_1383,N_1015,N_1090);
nand U1384 (N_1384,N_1034,N_1153);
or U1385 (N_1385,N_1099,N_1169);
or U1386 (N_1386,N_1083,N_1084);
or U1387 (N_1387,N_1135,N_1112);
nand U1388 (N_1388,N_1094,N_1056);
nand U1389 (N_1389,N_1152,N_1124);
nor U1390 (N_1390,N_1179,N_1083);
and U1391 (N_1391,N_1018,N_1042);
nor U1392 (N_1392,N_1089,N_1050);
or U1393 (N_1393,N_1140,N_1174);
xor U1394 (N_1394,N_1113,N_1068);
nand U1395 (N_1395,N_1186,N_1051);
and U1396 (N_1396,N_1075,N_1171);
or U1397 (N_1397,N_1024,N_1057);
nand U1398 (N_1398,N_1016,N_1083);
or U1399 (N_1399,N_1034,N_1169);
and U1400 (N_1400,N_1323,N_1262);
nor U1401 (N_1401,N_1398,N_1349);
and U1402 (N_1402,N_1280,N_1229);
nand U1403 (N_1403,N_1240,N_1288);
or U1404 (N_1404,N_1378,N_1319);
nor U1405 (N_1405,N_1223,N_1308);
and U1406 (N_1406,N_1351,N_1382);
and U1407 (N_1407,N_1213,N_1375);
and U1408 (N_1408,N_1331,N_1325);
or U1409 (N_1409,N_1304,N_1295);
nor U1410 (N_1410,N_1348,N_1285);
or U1411 (N_1411,N_1362,N_1340);
and U1412 (N_1412,N_1318,N_1283);
or U1413 (N_1413,N_1356,N_1233);
or U1414 (N_1414,N_1289,N_1200);
and U1415 (N_1415,N_1307,N_1207);
nand U1416 (N_1416,N_1274,N_1330);
or U1417 (N_1417,N_1371,N_1236);
and U1418 (N_1418,N_1328,N_1224);
and U1419 (N_1419,N_1374,N_1296);
nor U1420 (N_1420,N_1366,N_1367);
nor U1421 (N_1421,N_1248,N_1395);
nand U1422 (N_1422,N_1202,N_1214);
nand U1423 (N_1423,N_1335,N_1352);
and U1424 (N_1424,N_1279,N_1257);
or U1425 (N_1425,N_1327,N_1263);
nand U1426 (N_1426,N_1373,N_1222);
nor U1427 (N_1427,N_1282,N_1346);
nand U1428 (N_1428,N_1254,N_1302);
nor U1429 (N_1429,N_1394,N_1210);
or U1430 (N_1430,N_1251,N_1357);
nand U1431 (N_1431,N_1358,N_1321);
nor U1432 (N_1432,N_1238,N_1270);
and U1433 (N_1433,N_1332,N_1324);
xnor U1434 (N_1434,N_1291,N_1388);
or U1435 (N_1435,N_1230,N_1384);
nand U1436 (N_1436,N_1312,N_1347);
or U1437 (N_1437,N_1292,N_1255);
xor U1438 (N_1438,N_1290,N_1294);
or U1439 (N_1439,N_1343,N_1284);
and U1440 (N_1440,N_1281,N_1381);
and U1441 (N_1441,N_1370,N_1249);
or U1442 (N_1442,N_1361,N_1309);
and U1443 (N_1443,N_1221,N_1297);
nand U1444 (N_1444,N_1228,N_1344);
nor U1445 (N_1445,N_1271,N_1300);
and U1446 (N_1446,N_1258,N_1306);
and U1447 (N_1447,N_1365,N_1326);
nor U1448 (N_1448,N_1242,N_1208);
xor U1449 (N_1449,N_1341,N_1286);
or U1450 (N_1450,N_1231,N_1239);
and U1451 (N_1451,N_1252,N_1314);
and U1452 (N_1452,N_1215,N_1369);
or U1453 (N_1453,N_1276,N_1303);
xnor U1454 (N_1454,N_1336,N_1393);
or U1455 (N_1455,N_1338,N_1260);
nor U1456 (N_1456,N_1206,N_1219);
nand U1457 (N_1457,N_1265,N_1354);
nand U1458 (N_1458,N_1261,N_1277);
nor U1459 (N_1459,N_1272,N_1397);
nand U1460 (N_1460,N_1387,N_1390);
or U1461 (N_1461,N_1316,N_1235);
nor U1462 (N_1462,N_1256,N_1216);
and U1463 (N_1463,N_1350,N_1359);
nor U1464 (N_1464,N_1278,N_1264);
nand U1465 (N_1465,N_1315,N_1287);
and U1466 (N_1466,N_1396,N_1339);
and U1467 (N_1467,N_1203,N_1368);
nor U1468 (N_1468,N_1329,N_1201);
and U1469 (N_1469,N_1333,N_1334);
nor U1470 (N_1470,N_1268,N_1266);
or U1471 (N_1471,N_1386,N_1363);
and U1472 (N_1472,N_1345,N_1311);
or U1473 (N_1473,N_1391,N_1275);
xor U1474 (N_1474,N_1389,N_1246);
nand U1475 (N_1475,N_1205,N_1227);
nor U1476 (N_1476,N_1241,N_1320);
nor U1477 (N_1477,N_1392,N_1298);
and U1478 (N_1478,N_1209,N_1226);
nor U1479 (N_1479,N_1353,N_1372);
nor U1480 (N_1480,N_1220,N_1399);
and U1481 (N_1481,N_1310,N_1234);
and U1482 (N_1482,N_1376,N_1379);
and U1483 (N_1483,N_1243,N_1212);
xnor U1484 (N_1484,N_1247,N_1244);
nor U1485 (N_1485,N_1301,N_1322);
nor U1486 (N_1486,N_1313,N_1317);
or U1487 (N_1487,N_1232,N_1259);
nor U1488 (N_1488,N_1217,N_1299);
nand U1489 (N_1489,N_1253,N_1305);
nand U1490 (N_1490,N_1237,N_1385);
and U1491 (N_1491,N_1337,N_1364);
and U1492 (N_1492,N_1383,N_1211);
or U1493 (N_1493,N_1273,N_1377);
or U1494 (N_1494,N_1293,N_1250);
nor U1495 (N_1495,N_1225,N_1380);
and U1496 (N_1496,N_1342,N_1245);
and U1497 (N_1497,N_1269,N_1360);
and U1498 (N_1498,N_1204,N_1355);
or U1499 (N_1499,N_1267,N_1218);
and U1500 (N_1500,N_1294,N_1323);
or U1501 (N_1501,N_1241,N_1202);
nand U1502 (N_1502,N_1348,N_1263);
nand U1503 (N_1503,N_1324,N_1242);
nor U1504 (N_1504,N_1312,N_1284);
and U1505 (N_1505,N_1242,N_1307);
nand U1506 (N_1506,N_1305,N_1354);
nor U1507 (N_1507,N_1368,N_1261);
and U1508 (N_1508,N_1369,N_1301);
nor U1509 (N_1509,N_1378,N_1227);
or U1510 (N_1510,N_1210,N_1335);
and U1511 (N_1511,N_1311,N_1265);
or U1512 (N_1512,N_1222,N_1335);
nand U1513 (N_1513,N_1242,N_1272);
or U1514 (N_1514,N_1212,N_1371);
nor U1515 (N_1515,N_1341,N_1240);
or U1516 (N_1516,N_1304,N_1310);
nor U1517 (N_1517,N_1281,N_1330);
xor U1518 (N_1518,N_1330,N_1360);
or U1519 (N_1519,N_1217,N_1301);
nor U1520 (N_1520,N_1275,N_1272);
or U1521 (N_1521,N_1229,N_1396);
nor U1522 (N_1522,N_1266,N_1299);
nor U1523 (N_1523,N_1201,N_1350);
nand U1524 (N_1524,N_1328,N_1250);
and U1525 (N_1525,N_1339,N_1280);
nor U1526 (N_1526,N_1252,N_1229);
and U1527 (N_1527,N_1262,N_1395);
or U1528 (N_1528,N_1268,N_1257);
nor U1529 (N_1529,N_1364,N_1386);
and U1530 (N_1530,N_1275,N_1225);
nand U1531 (N_1531,N_1218,N_1279);
and U1532 (N_1532,N_1394,N_1354);
or U1533 (N_1533,N_1280,N_1271);
or U1534 (N_1534,N_1250,N_1225);
and U1535 (N_1535,N_1333,N_1291);
nand U1536 (N_1536,N_1262,N_1211);
xor U1537 (N_1537,N_1273,N_1379);
nand U1538 (N_1538,N_1206,N_1372);
or U1539 (N_1539,N_1349,N_1324);
nor U1540 (N_1540,N_1229,N_1379);
nor U1541 (N_1541,N_1343,N_1330);
nand U1542 (N_1542,N_1345,N_1330);
nor U1543 (N_1543,N_1302,N_1292);
and U1544 (N_1544,N_1272,N_1220);
nor U1545 (N_1545,N_1279,N_1369);
and U1546 (N_1546,N_1382,N_1313);
nand U1547 (N_1547,N_1376,N_1267);
xnor U1548 (N_1548,N_1287,N_1248);
or U1549 (N_1549,N_1334,N_1287);
nand U1550 (N_1550,N_1381,N_1376);
nor U1551 (N_1551,N_1222,N_1280);
or U1552 (N_1552,N_1352,N_1333);
nand U1553 (N_1553,N_1202,N_1385);
or U1554 (N_1554,N_1204,N_1363);
nand U1555 (N_1555,N_1208,N_1323);
nor U1556 (N_1556,N_1342,N_1252);
nor U1557 (N_1557,N_1371,N_1219);
or U1558 (N_1558,N_1290,N_1349);
or U1559 (N_1559,N_1293,N_1370);
and U1560 (N_1560,N_1263,N_1242);
or U1561 (N_1561,N_1237,N_1314);
nor U1562 (N_1562,N_1289,N_1204);
or U1563 (N_1563,N_1304,N_1207);
nand U1564 (N_1564,N_1278,N_1327);
and U1565 (N_1565,N_1296,N_1307);
and U1566 (N_1566,N_1378,N_1271);
nor U1567 (N_1567,N_1349,N_1213);
or U1568 (N_1568,N_1299,N_1287);
or U1569 (N_1569,N_1307,N_1259);
and U1570 (N_1570,N_1319,N_1365);
nand U1571 (N_1571,N_1343,N_1218);
nand U1572 (N_1572,N_1354,N_1350);
or U1573 (N_1573,N_1234,N_1228);
nor U1574 (N_1574,N_1204,N_1380);
nand U1575 (N_1575,N_1341,N_1359);
or U1576 (N_1576,N_1334,N_1392);
nor U1577 (N_1577,N_1225,N_1328);
and U1578 (N_1578,N_1315,N_1391);
or U1579 (N_1579,N_1214,N_1273);
or U1580 (N_1580,N_1272,N_1268);
nor U1581 (N_1581,N_1230,N_1289);
nor U1582 (N_1582,N_1247,N_1266);
nor U1583 (N_1583,N_1281,N_1329);
nand U1584 (N_1584,N_1319,N_1202);
or U1585 (N_1585,N_1361,N_1240);
or U1586 (N_1586,N_1226,N_1319);
or U1587 (N_1587,N_1279,N_1248);
and U1588 (N_1588,N_1204,N_1290);
xnor U1589 (N_1589,N_1272,N_1239);
nand U1590 (N_1590,N_1246,N_1227);
nor U1591 (N_1591,N_1297,N_1238);
and U1592 (N_1592,N_1391,N_1385);
nand U1593 (N_1593,N_1245,N_1387);
xor U1594 (N_1594,N_1268,N_1347);
or U1595 (N_1595,N_1334,N_1281);
nand U1596 (N_1596,N_1342,N_1343);
nor U1597 (N_1597,N_1244,N_1313);
and U1598 (N_1598,N_1394,N_1299);
nand U1599 (N_1599,N_1387,N_1343);
and U1600 (N_1600,N_1538,N_1473);
or U1601 (N_1601,N_1438,N_1520);
nand U1602 (N_1602,N_1483,N_1418);
nor U1603 (N_1603,N_1401,N_1581);
nor U1604 (N_1604,N_1505,N_1465);
nand U1605 (N_1605,N_1569,N_1543);
or U1606 (N_1606,N_1459,N_1453);
xor U1607 (N_1607,N_1468,N_1457);
and U1608 (N_1608,N_1576,N_1404);
nor U1609 (N_1609,N_1405,N_1494);
nor U1610 (N_1610,N_1416,N_1501);
nand U1611 (N_1611,N_1429,N_1564);
nand U1612 (N_1612,N_1574,N_1474);
nand U1613 (N_1613,N_1550,N_1560);
nor U1614 (N_1614,N_1544,N_1534);
nand U1615 (N_1615,N_1570,N_1517);
nand U1616 (N_1616,N_1578,N_1491);
nand U1617 (N_1617,N_1589,N_1565);
or U1618 (N_1618,N_1488,N_1524);
nor U1619 (N_1619,N_1558,N_1500);
nor U1620 (N_1620,N_1423,N_1561);
or U1621 (N_1621,N_1425,N_1419);
nor U1622 (N_1622,N_1499,N_1514);
nand U1623 (N_1623,N_1434,N_1469);
nor U1624 (N_1624,N_1413,N_1446);
or U1625 (N_1625,N_1445,N_1493);
and U1626 (N_1626,N_1542,N_1503);
and U1627 (N_1627,N_1531,N_1489);
or U1628 (N_1628,N_1443,N_1484);
and U1629 (N_1629,N_1479,N_1519);
nand U1630 (N_1630,N_1566,N_1512);
and U1631 (N_1631,N_1596,N_1462);
nor U1632 (N_1632,N_1539,N_1417);
nor U1633 (N_1633,N_1487,N_1593);
nand U1634 (N_1634,N_1412,N_1437);
nand U1635 (N_1635,N_1571,N_1521);
or U1636 (N_1636,N_1495,N_1458);
nor U1637 (N_1637,N_1518,N_1466);
nand U1638 (N_1638,N_1477,N_1448);
nand U1639 (N_1639,N_1553,N_1584);
and U1640 (N_1640,N_1575,N_1470);
or U1641 (N_1641,N_1486,N_1563);
nor U1642 (N_1642,N_1433,N_1400);
nand U1643 (N_1643,N_1594,N_1568);
xor U1644 (N_1644,N_1585,N_1508);
and U1645 (N_1645,N_1573,N_1579);
nor U1646 (N_1646,N_1450,N_1535);
and U1647 (N_1647,N_1454,N_1409);
and U1648 (N_1648,N_1480,N_1440);
and U1649 (N_1649,N_1427,N_1536);
nor U1650 (N_1650,N_1513,N_1464);
nor U1651 (N_1651,N_1452,N_1592);
or U1652 (N_1652,N_1481,N_1410);
nand U1653 (N_1653,N_1547,N_1522);
nor U1654 (N_1654,N_1455,N_1475);
nor U1655 (N_1655,N_1548,N_1421);
and U1656 (N_1656,N_1554,N_1406);
nand U1657 (N_1657,N_1502,N_1567);
and U1658 (N_1658,N_1467,N_1533);
or U1659 (N_1659,N_1580,N_1528);
nand U1660 (N_1660,N_1557,N_1408);
and U1661 (N_1661,N_1583,N_1476);
or U1662 (N_1662,N_1456,N_1598);
nand U1663 (N_1663,N_1595,N_1439);
nand U1664 (N_1664,N_1428,N_1432);
nand U1665 (N_1665,N_1422,N_1478);
nor U1666 (N_1666,N_1496,N_1435);
and U1667 (N_1667,N_1591,N_1451);
nor U1668 (N_1668,N_1444,N_1407);
nor U1669 (N_1669,N_1582,N_1402);
or U1670 (N_1670,N_1590,N_1526);
or U1671 (N_1671,N_1597,N_1449);
nand U1672 (N_1672,N_1507,N_1532);
or U1673 (N_1673,N_1424,N_1463);
nand U1674 (N_1674,N_1461,N_1546);
or U1675 (N_1675,N_1586,N_1414);
and U1676 (N_1676,N_1411,N_1485);
and U1677 (N_1677,N_1497,N_1577);
nand U1678 (N_1678,N_1525,N_1431);
nor U1679 (N_1679,N_1559,N_1552);
nor U1680 (N_1680,N_1545,N_1530);
nand U1681 (N_1681,N_1420,N_1509);
or U1682 (N_1682,N_1556,N_1537);
nand U1683 (N_1683,N_1541,N_1527);
and U1684 (N_1684,N_1540,N_1506);
nor U1685 (N_1685,N_1587,N_1510);
nand U1686 (N_1686,N_1472,N_1482);
and U1687 (N_1687,N_1442,N_1498);
and U1688 (N_1688,N_1430,N_1460);
nand U1689 (N_1689,N_1572,N_1588);
and U1690 (N_1690,N_1504,N_1426);
nand U1691 (N_1691,N_1471,N_1436);
nand U1692 (N_1692,N_1551,N_1529);
and U1693 (N_1693,N_1523,N_1562);
nor U1694 (N_1694,N_1516,N_1549);
or U1695 (N_1695,N_1599,N_1415);
nand U1696 (N_1696,N_1555,N_1490);
nand U1697 (N_1697,N_1492,N_1515);
nor U1698 (N_1698,N_1441,N_1511);
nor U1699 (N_1699,N_1447,N_1403);
and U1700 (N_1700,N_1579,N_1501);
or U1701 (N_1701,N_1436,N_1442);
nor U1702 (N_1702,N_1529,N_1489);
and U1703 (N_1703,N_1521,N_1566);
nor U1704 (N_1704,N_1530,N_1581);
or U1705 (N_1705,N_1538,N_1499);
nand U1706 (N_1706,N_1418,N_1513);
or U1707 (N_1707,N_1468,N_1547);
nand U1708 (N_1708,N_1575,N_1461);
and U1709 (N_1709,N_1487,N_1579);
and U1710 (N_1710,N_1441,N_1422);
nor U1711 (N_1711,N_1581,N_1422);
and U1712 (N_1712,N_1465,N_1452);
nor U1713 (N_1713,N_1567,N_1456);
nand U1714 (N_1714,N_1433,N_1572);
nor U1715 (N_1715,N_1482,N_1521);
nor U1716 (N_1716,N_1456,N_1405);
and U1717 (N_1717,N_1536,N_1584);
and U1718 (N_1718,N_1523,N_1511);
nor U1719 (N_1719,N_1573,N_1429);
and U1720 (N_1720,N_1527,N_1463);
nor U1721 (N_1721,N_1442,N_1486);
and U1722 (N_1722,N_1549,N_1512);
nor U1723 (N_1723,N_1444,N_1502);
or U1724 (N_1724,N_1534,N_1451);
nor U1725 (N_1725,N_1552,N_1537);
nor U1726 (N_1726,N_1413,N_1591);
and U1727 (N_1727,N_1419,N_1529);
and U1728 (N_1728,N_1529,N_1570);
nor U1729 (N_1729,N_1430,N_1585);
or U1730 (N_1730,N_1510,N_1549);
or U1731 (N_1731,N_1541,N_1584);
or U1732 (N_1732,N_1433,N_1509);
nand U1733 (N_1733,N_1462,N_1423);
nand U1734 (N_1734,N_1487,N_1439);
or U1735 (N_1735,N_1428,N_1590);
nand U1736 (N_1736,N_1447,N_1596);
and U1737 (N_1737,N_1560,N_1450);
or U1738 (N_1738,N_1545,N_1415);
nor U1739 (N_1739,N_1482,N_1489);
and U1740 (N_1740,N_1422,N_1540);
and U1741 (N_1741,N_1593,N_1462);
or U1742 (N_1742,N_1408,N_1409);
and U1743 (N_1743,N_1426,N_1571);
or U1744 (N_1744,N_1508,N_1567);
or U1745 (N_1745,N_1478,N_1402);
or U1746 (N_1746,N_1419,N_1554);
nor U1747 (N_1747,N_1485,N_1434);
and U1748 (N_1748,N_1552,N_1589);
nand U1749 (N_1749,N_1564,N_1509);
nand U1750 (N_1750,N_1408,N_1590);
nand U1751 (N_1751,N_1429,N_1532);
nor U1752 (N_1752,N_1554,N_1510);
nand U1753 (N_1753,N_1494,N_1417);
and U1754 (N_1754,N_1599,N_1455);
nor U1755 (N_1755,N_1567,N_1441);
nor U1756 (N_1756,N_1448,N_1483);
nor U1757 (N_1757,N_1450,N_1423);
or U1758 (N_1758,N_1578,N_1544);
nand U1759 (N_1759,N_1556,N_1571);
nor U1760 (N_1760,N_1408,N_1514);
or U1761 (N_1761,N_1554,N_1579);
nand U1762 (N_1762,N_1513,N_1436);
nand U1763 (N_1763,N_1456,N_1510);
or U1764 (N_1764,N_1551,N_1420);
nor U1765 (N_1765,N_1432,N_1473);
and U1766 (N_1766,N_1535,N_1405);
nand U1767 (N_1767,N_1411,N_1573);
or U1768 (N_1768,N_1494,N_1444);
nor U1769 (N_1769,N_1521,N_1593);
or U1770 (N_1770,N_1454,N_1507);
nor U1771 (N_1771,N_1520,N_1404);
or U1772 (N_1772,N_1530,N_1436);
nand U1773 (N_1773,N_1496,N_1409);
nand U1774 (N_1774,N_1454,N_1557);
or U1775 (N_1775,N_1443,N_1578);
nand U1776 (N_1776,N_1559,N_1547);
nand U1777 (N_1777,N_1573,N_1542);
nor U1778 (N_1778,N_1430,N_1421);
nand U1779 (N_1779,N_1544,N_1511);
and U1780 (N_1780,N_1596,N_1537);
nor U1781 (N_1781,N_1578,N_1535);
nand U1782 (N_1782,N_1545,N_1511);
and U1783 (N_1783,N_1545,N_1566);
nand U1784 (N_1784,N_1591,N_1521);
and U1785 (N_1785,N_1540,N_1481);
or U1786 (N_1786,N_1568,N_1468);
and U1787 (N_1787,N_1451,N_1566);
or U1788 (N_1788,N_1570,N_1422);
nor U1789 (N_1789,N_1414,N_1528);
nand U1790 (N_1790,N_1445,N_1581);
nand U1791 (N_1791,N_1496,N_1451);
and U1792 (N_1792,N_1584,N_1498);
nor U1793 (N_1793,N_1594,N_1416);
or U1794 (N_1794,N_1432,N_1516);
nand U1795 (N_1795,N_1435,N_1405);
or U1796 (N_1796,N_1433,N_1546);
or U1797 (N_1797,N_1412,N_1401);
and U1798 (N_1798,N_1591,N_1530);
or U1799 (N_1799,N_1591,N_1487);
or U1800 (N_1800,N_1779,N_1638);
nor U1801 (N_1801,N_1601,N_1753);
or U1802 (N_1802,N_1796,N_1630);
nor U1803 (N_1803,N_1651,N_1609);
or U1804 (N_1804,N_1770,N_1735);
nand U1805 (N_1805,N_1680,N_1765);
or U1806 (N_1806,N_1727,N_1722);
and U1807 (N_1807,N_1681,N_1768);
nor U1808 (N_1808,N_1625,N_1730);
and U1809 (N_1809,N_1613,N_1662);
and U1810 (N_1810,N_1612,N_1707);
or U1811 (N_1811,N_1710,N_1665);
and U1812 (N_1812,N_1658,N_1604);
and U1813 (N_1813,N_1701,N_1628);
nand U1814 (N_1814,N_1700,N_1656);
and U1815 (N_1815,N_1754,N_1783);
nor U1816 (N_1816,N_1782,N_1657);
xnor U1817 (N_1817,N_1745,N_1675);
and U1818 (N_1818,N_1706,N_1702);
and U1819 (N_1819,N_1704,N_1729);
nor U1820 (N_1820,N_1763,N_1611);
nor U1821 (N_1821,N_1679,N_1758);
nor U1822 (N_1822,N_1624,N_1705);
nor U1823 (N_1823,N_1654,N_1622);
or U1824 (N_1824,N_1762,N_1644);
nor U1825 (N_1825,N_1775,N_1797);
or U1826 (N_1826,N_1648,N_1637);
nand U1827 (N_1827,N_1798,N_1607);
and U1828 (N_1828,N_1723,N_1732);
or U1829 (N_1829,N_1635,N_1694);
or U1830 (N_1830,N_1776,N_1653);
nand U1831 (N_1831,N_1716,N_1719);
and U1832 (N_1832,N_1640,N_1688);
or U1833 (N_1833,N_1699,N_1642);
nand U1834 (N_1834,N_1743,N_1731);
or U1835 (N_1835,N_1695,N_1605);
and U1836 (N_1836,N_1767,N_1650);
and U1837 (N_1837,N_1717,N_1713);
xor U1838 (N_1838,N_1616,N_1621);
nand U1839 (N_1839,N_1690,N_1771);
nand U1840 (N_1840,N_1632,N_1666);
and U1841 (N_1841,N_1721,N_1618);
or U1842 (N_1842,N_1684,N_1734);
nand U1843 (N_1843,N_1639,N_1649);
nand U1844 (N_1844,N_1795,N_1691);
nand U1845 (N_1845,N_1655,N_1672);
nor U1846 (N_1846,N_1766,N_1693);
nand U1847 (N_1847,N_1714,N_1617);
and U1848 (N_1848,N_1772,N_1641);
or U1849 (N_1849,N_1606,N_1749);
and U1850 (N_1850,N_1787,N_1646);
and U1851 (N_1851,N_1778,N_1711);
and U1852 (N_1852,N_1603,N_1724);
xor U1853 (N_1853,N_1676,N_1741);
nor U1854 (N_1854,N_1652,N_1739);
nand U1855 (N_1855,N_1687,N_1602);
and U1856 (N_1856,N_1686,N_1627);
nand U1857 (N_1857,N_1788,N_1709);
or U1858 (N_1858,N_1760,N_1789);
nand U1859 (N_1859,N_1769,N_1720);
nand U1860 (N_1860,N_1660,N_1633);
nor U1861 (N_1861,N_1683,N_1751);
nand U1862 (N_1862,N_1623,N_1670);
or U1863 (N_1863,N_1661,N_1764);
nor U1864 (N_1864,N_1696,N_1752);
nand U1865 (N_1865,N_1793,N_1647);
nor U1866 (N_1866,N_1738,N_1733);
or U1867 (N_1867,N_1750,N_1689);
and U1868 (N_1868,N_1792,N_1740);
nand U1869 (N_1869,N_1600,N_1703);
nand U1870 (N_1870,N_1669,N_1664);
nand U1871 (N_1871,N_1742,N_1698);
and U1872 (N_1872,N_1748,N_1626);
and U1873 (N_1873,N_1791,N_1799);
or U1874 (N_1874,N_1744,N_1610);
and U1875 (N_1875,N_1794,N_1774);
nor U1876 (N_1876,N_1608,N_1667);
and U1877 (N_1877,N_1645,N_1682);
or U1878 (N_1878,N_1777,N_1692);
nor U1879 (N_1879,N_1784,N_1629);
xnor U1880 (N_1880,N_1755,N_1790);
nand U1881 (N_1881,N_1785,N_1747);
nand U1882 (N_1882,N_1757,N_1614);
nand U1883 (N_1883,N_1786,N_1718);
xor U1884 (N_1884,N_1697,N_1615);
and U1885 (N_1885,N_1773,N_1659);
and U1886 (N_1886,N_1671,N_1678);
nor U1887 (N_1887,N_1736,N_1715);
or U1888 (N_1888,N_1620,N_1726);
or U1889 (N_1889,N_1728,N_1674);
nor U1890 (N_1890,N_1756,N_1643);
and U1891 (N_1891,N_1668,N_1619);
or U1892 (N_1892,N_1677,N_1737);
or U1893 (N_1893,N_1780,N_1634);
or U1894 (N_1894,N_1636,N_1708);
nor U1895 (N_1895,N_1712,N_1631);
nand U1896 (N_1896,N_1761,N_1759);
nor U1897 (N_1897,N_1781,N_1673);
or U1898 (N_1898,N_1663,N_1746);
nand U1899 (N_1899,N_1725,N_1685);
or U1900 (N_1900,N_1644,N_1707);
nor U1901 (N_1901,N_1789,N_1727);
nor U1902 (N_1902,N_1726,N_1782);
nor U1903 (N_1903,N_1796,N_1658);
xnor U1904 (N_1904,N_1752,N_1656);
nand U1905 (N_1905,N_1638,N_1654);
and U1906 (N_1906,N_1771,N_1698);
and U1907 (N_1907,N_1627,N_1668);
nand U1908 (N_1908,N_1628,N_1699);
or U1909 (N_1909,N_1759,N_1638);
and U1910 (N_1910,N_1610,N_1657);
and U1911 (N_1911,N_1713,N_1687);
and U1912 (N_1912,N_1642,N_1738);
nand U1913 (N_1913,N_1600,N_1677);
and U1914 (N_1914,N_1762,N_1706);
or U1915 (N_1915,N_1601,N_1676);
nor U1916 (N_1916,N_1706,N_1666);
nand U1917 (N_1917,N_1733,N_1647);
nor U1918 (N_1918,N_1618,N_1725);
nor U1919 (N_1919,N_1760,N_1751);
nor U1920 (N_1920,N_1788,N_1675);
and U1921 (N_1921,N_1762,N_1607);
nor U1922 (N_1922,N_1733,N_1610);
or U1923 (N_1923,N_1734,N_1794);
or U1924 (N_1924,N_1792,N_1619);
or U1925 (N_1925,N_1645,N_1611);
nor U1926 (N_1926,N_1758,N_1792);
or U1927 (N_1927,N_1632,N_1692);
nor U1928 (N_1928,N_1658,N_1776);
nand U1929 (N_1929,N_1661,N_1762);
nor U1930 (N_1930,N_1762,N_1754);
or U1931 (N_1931,N_1765,N_1651);
nand U1932 (N_1932,N_1628,N_1795);
nand U1933 (N_1933,N_1643,N_1755);
nor U1934 (N_1934,N_1765,N_1623);
nand U1935 (N_1935,N_1635,N_1639);
nand U1936 (N_1936,N_1654,N_1694);
nand U1937 (N_1937,N_1610,N_1782);
xnor U1938 (N_1938,N_1730,N_1637);
or U1939 (N_1939,N_1680,N_1700);
or U1940 (N_1940,N_1698,N_1769);
nand U1941 (N_1941,N_1777,N_1619);
nand U1942 (N_1942,N_1781,N_1639);
nand U1943 (N_1943,N_1701,N_1600);
or U1944 (N_1944,N_1665,N_1645);
or U1945 (N_1945,N_1713,N_1737);
or U1946 (N_1946,N_1678,N_1700);
or U1947 (N_1947,N_1606,N_1667);
nand U1948 (N_1948,N_1703,N_1769);
nand U1949 (N_1949,N_1605,N_1748);
nand U1950 (N_1950,N_1680,N_1745);
nor U1951 (N_1951,N_1766,N_1673);
nor U1952 (N_1952,N_1779,N_1756);
nand U1953 (N_1953,N_1761,N_1654);
nor U1954 (N_1954,N_1632,N_1678);
nand U1955 (N_1955,N_1795,N_1799);
nand U1956 (N_1956,N_1710,N_1768);
nand U1957 (N_1957,N_1619,N_1602);
or U1958 (N_1958,N_1779,N_1723);
nand U1959 (N_1959,N_1686,N_1689);
nor U1960 (N_1960,N_1792,N_1683);
nand U1961 (N_1961,N_1654,N_1679);
and U1962 (N_1962,N_1627,N_1754);
and U1963 (N_1963,N_1679,N_1717);
and U1964 (N_1964,N_1768,N_1668);
nor U1965 (N_1965,N_1747,N_1707);
or U1966 (N_1966,N_1709,N_1730);
nand U1967 (N_1967,N_1612,N_1724);
nor U1968 (N_1968,N_1675,N_1692);
nand U1969 (N_1969,N_1601,N_1785);
nand U1970 (N_1970,N_1764,N_1759);
nand U1971 (N_1971,N_1636,N_1797);
and U1972 (N_1972,N_1662,N_1758);
nand U1973 (N_1973,N_1733,N_1651);
and U1974 (N_1974,N_1613,N_1687);
nand U1975 (N_1975,N_1771,N_1604);
and U1976 (N_1976,N_1701,N_1789);
and U1977 (N_1977,N_1719,N_1796);
nor U1978 (N_1978,N_1697,N_1797);
and U1979 (N_1979,N_1708,N_1731);
nand U1980 (N_1980,N_1670,N_1681);
and U1981 (N_1981,N_1771,N_1761);
nor U1982 (N_1982,N_1634,N_1755);
nor U1983 (N_1983,N_1782,N_1744);
and U1984 (N_1984,N_1628,N_1767);
or U1985 (N_1985,N_1645,N_1614);
and U1986 (N_1986,N_1605,N_1636);
and U1987 (N_1987,N_1706,N_1653);
nand U1988 (N_1988,N_1600,N_1798);
nand U1989 (N_1989,N_1789,N_1649);
nor U1990 (N_1990,N_1698,N_1692);
and U1991 (N_1991,N_1695,N_1725);
xnor U1992 (N_1992,N_1637,N_1676);
nor U1993 (N_1993,N_1776,N_1623);
nand U1994 (N_1994,N_1768,N_1720);
and U1995 (N_1995,N_1788,N_1605);
nand U1996 (N_1996,N_1623,N_1671);
nand U1997 (N_1997,N_1677,N_1667);
nand U1998 (N_1998,N_1600,N_1761);
or U1999 (N_1999,N_1704,N_1754);
or U2000 (N_2000,N_1982,N_1836);
nor U2001 (N_2001,N_1975,N_1979);
nor U2002 (N_2002,N_1977,N_1919);
or U2003 (N_2003,N_1968,N_1832);
nor U2004 (N_2004,N_1992,N_1825);
and U2005 (N_2005,N_1960,N_1953);
or U2006 (N_2006,N_1964,N_1959);
nand U2007 (N_2007,N_1942,N_1864);
nor U2008 (N_2008,N_1904,N_1830);
nand U2009 (N_2009,N_1926,N_1909);
xnor U2010 (N_2010,N_1954,N_1823);
nor U2011 (N_2011,N_1886,N_1974);
and U2012 (N_2012,N_1885,N_1848);
and U2013 (N_2013,N_1843,N_1944);
or U2014 (N_2014,N_1872,N_1901);
nand U2015 (N_2015,N_1898,N_1950);
nand U2016 (N_2016,N_1859,N_1805);
nor U2017 (N_2017,N_1895,N_1856);
nand U2018 (N_2018,N_1849,N_1932);
and U2019 (N_2019,N_1930,N_1994);
nand U2020 (N_2020,N_1854,N_1833);
nor U2021 (N_2021,N_1837,N_1870);
and U2022 (N_2022,N_1902,N_1815);
or U2023 (N_2023,N_1998,N_1827);
nor U2024 (N_2024,N_1809,N_1946);
and U2025 (N_2025,N_1985,N_1967);
nand U2026 (N_2026,N_1922,N_1881);
or U2027 (N_2027,N_1911,N_1811);
or U2028 (N_2028,N_1966,N_1822);
and U2029 (N_2029,N_1812,N_1853);
nor U2030 (N_2030,N_1842,N_1996);
nor U2031 (N_2031,N_1949,N_1986);
nor U2032 (N_2032,N_1965,N_1973);
nor U2033 (N_2033,N_1857,N_1971);
nor U2034 (N_2034,N_1889,N_1955);
nand U2035 (N_2035,N_1925,N_1816);
or U2036 (N_2036,N_1906,N_1903);
and U2037 (N_2037,N_1999,N_1858);
nor U2038 (N_2038,N_1908,N_1867);
and U2039 (N_2039,N_1957,N_1927);
nor U2040 (N_2040,N_1851,N_1892);
nand U2041 (N_2041,N_1874,N_1875);
and U2042 (N_2042,N_1810,N_1880);
xnor U2043 (N_2043,N_1924,N_1915);
or U2044 (N_2044,N_1988,N_1945);
or U2045 (N_2045,N_1993,N_1984);
or U2046 (N_2046,N_1838,N_1804);
nor U2047 (N_2047,N_1876,N_1987);
or U2048 (N_2048,N_1914,N_1862);
nand U2049 (N_2049,N_1929,N_1978);
or U2050 (N_2050,N_1920,N_1869);
and U2051 (N_2051,N_1890,N_1882);
and U2052 (N_2052,N_1948,N_1800);
and U2053 (N_2053,N_1983,N_1940);
nor U2054 (N_2054,N_1819,N_1845);
nor U2055 (N_2055,N_1861,N_1961);
nand U2056 (N_2056,N_1818,N_1918);
and U2057 (N_2057,N_1888,N_1826);
nor U2058 (N_2058,N_1820,N_1936);
and U2059 (N_2059,N_1990,N_1943);
nand U2060 (N_2060,N_1947,N_1928);
nor U2061 (N_2061,N_1912,N_1962);
and U2062 (N_2062,N_1891,N_1871);
nand U2063 (N_2063,N_1831,N_1807);
and U2064 (N_2064,N_1899,N_1850);
nand U2065 (N_2065,N_1824,N_1860);
or U2066 (N_2066,N_1934,N_1941);
or U2067 (N_2067,N_1879,N_1887);
or U2068 (N_2068,N_1863,N_1835);
nor U2069 (N_2069,N_1802,N_1840);
nor U2070 (N_2070,N_1956,N_1834);
nor U2071 (N_2071,N_1855,N_1923);
nand U2072 (N_2072,N_1893,N_1910);
or U2073 (N_2073,N_1829,N_1817);
nor U2074 (N_2074,N_1896,N_1801);
nor U2075 (N_2075,N_1907,N_1821);
or U2076 (N_2076,N_1852,N_1866);
nand U2077 (N_2077,N_1803,N_1933);
or U2078 (N_2078,N_1917,N_1916);
and U2079 (N_2079,N_1931,N_1958);
nand U2080 (N_2080,N_1813,N_1839);
or U2081 (N_2081,N_1897,N_1970);
nor U2082 (N_2082,N_1841,N_1976);
and U2083 (N_2083,N_1877,N_1963);
and U2084 (N_2084,N_1935,N_1952);
or U2085 (N_2085,N_1913,N_1883);
and U2086 (N_2086,N_1938,N_1969);
or U2087 (N_2087,N_1844,N_1847);
nand U2088 (N_2088,N_1981,N_1980);
or U2089 (N_2089,N_1814,N_1878);
nand U2090 (N_2090,N_1937,N_1991);
and U2091 (N_2091,N_1808,N_1951);
and U2092 (N_2092,N_1865,N_1921);
or U2093 (N_2093,N_1884,N_1828);
nand U2094 (N_2094,N_1995,N_1846);
nand U2095 (N_2095,N_1873,N_1900);
and U2096 (N_2096,N_1894,N_1989);
and U2097 (N_2097,N_1972,N_1939);
and U2098 (N_2098,N_1806,N_1997);
or U2099 (N_2099,N_1868,N_1905);
or U2100 (N_2100,N_1991,N_1824);
or U2101 (N_2101,N_1916,N_1928);
or U2102 (N_2102,N_1944,N_1948);
nand U2103 (N_2103,N_1940,N_1828);
and U2104 (N_2104,N_1927,N_1819);
or U2105 (N_2105,N_1856,N_1924);
and U2106 (N_2106,N_1872,N_1892);
nor U2107 (N_2107,N_1887,N_1827);
or U2108 (N_2108,N_1924,N_1976);
and U2109 (N_2109,N_1881,N_1981);
nor U2110 (N_2110,N_1953,N_1999);
nand U2111 (N_2111,N_1885,N_1842);
nor U2112 (N_2112,N_1821,N_1830);
nor U2113 (N_2113,N_1897,N_1840);
or U2114 (N_2114,N_1952,N_1836);
nor U2115 (N_2115,N_1864,N_1881);
nor U2116 (N_2116,N_1907,N_1888);
nand U2117 (N_2117,N_1879,N_1816);
nor U2118 (N_2118,N_1823,N_1965);
or U2119 (N_2119,N_1804,N_1933);
and U2120 (N_2120,N_1855,N_1858);
or U2121 (N_2121,N_1964,N_1961);
nand U2122 (N_2122,N_1942,N_1862);
and U2123 (N_2123,N_1888,N_1932);
nor U2124 (N_2124,N_1946,N_1838);
or U2125 (N_2125,N_1952,N_1943);
and U2126 (N_2126,N_1937,N_1867);
nand U2127 (N_2127,N_1929,N_1899);
or U2128 (N_2128,N_1878,N_1924);
or U2129 (N_2129,N_1910,N_1903);
and U2130 (N_2130,N_1845,N_1963);
nand U2131 (N_2131,N_1845,N_1940);
nor U2132 (N_2132,N_1884,N_1962);
and U2133 (N_2133,N_1943,N_1941);
or U2134 (N_2134,N_1877,N_1978);
or U2135 (N_2135,N_1801,N_1868);
nand U2136 (N_2136,N_1864,N_1986);
nor U2137 (N_2137,N_1878,N_1916);
or U2138 (N_2138,N_1919,N_1976);
or U2139 (N_2139,N_1926,N_1998);
and U2140 (N_2140,N_1822,N_1905);
or U2141 (N_2141,N_1869,N_1959);
nand U2142 (N_2142,N_1828,N_1955);
nand U2143 (N_2143,N_1838,N_1925);
xnor U2144 (N_2144,N_1801,N_1928);
and U2145 (N_2145,N_1981,N_1859);
nand U2146 (N_2146,N_1933,N_1929);
nor U2147 (N_2147,N_1919,N_1908);
nor U2148 (N_2148,N_1839,N_1832);
or U2149 (N_2149,N_1842,N_1874);
and U2150 (N_2150,N_1928,N_1997);
nand U2151 (N_2151,N_1884,N_1889);
nand U2152 (N_2152,N_1876,N_1804);
or U2153 (N_2153,N_1888,N_1961);
nand U2154 (N_2154,N_1967,N_1986);
or U2155 (N_2155,N_1821,N_1815);
nand U2156 (N_2156,N_1990,N_1880);
or U2157 (N_2157,N_1857,N_1845);
nor U2158 (N_2158,N_1810,N_1914);
nand U2159 (N_2159,N_1849,N_1923);
nand U2160 (N_2160,N_1927,N_1843);
nand U2161 (N_2161,N_1920,N_1808);
nor U2162 (N_2162,N_1965,N_1857);
nor U2163 (N_2163,N_1952,N_1909);
and U2164 (N_2164,N_1803,N_1843);
or U2165 (N_2165,N_1821,N_1810);
nor U2166 (N_2166,N_1940,N_1811);
or U2167 (N_2167,N_1884,N_1987);
nor U2168 (N_2168,N_1901,N_1965);
and U2169 (N_2169,N_1817,N_1803);
nor U2170 (N_2170,N_1882,N_1836);
nor U2171 (N_2171,N_1823,N_1980);
nor U2172 (N_2172,N_1977,N_1900);
nor U2173 (N_2173,N_1827,N_1897);
or U2174 (N_2174,N_1891,N_1835);
and U2175 (N_2175,N_1924,N_1812);
and U2176 (N_2176,N_1857,N_1893);
or U2177 (N_2177,N_1830,N_1892);
and U2178 (N_2178,N_1903,N_1969);
nor U2179 (N_2179,N_1922,N_1877);
xnor U2180 (N_2180,N_1932,N_1812);
or U2181 (N_2181,N_1851,N_1866);
or U2182 (N_2182,N_1964,N_1940);
nand U2183 (N_2183,N_1804,N_1909);
or U2184 (N_2184,N_1898,N_1993);
or U2185 (N_2185,N_1962,N_1844);
or U2186 (N_2186,N_1806,N_1983);
nand U2187 (N_2187,N_1975,N_1876);
nand U2188 (N_2188,N_1924,N_1948);
or U2189 (N_2189,N_1933,N_1957);
nor U2190 (N_2190,N_1880,N_1838);
nand U2191 (N_2191,N_1977,N_1880);
nor U2192 (N_2192,N_1932,N_1802);
nor U2193 (N_2193,N_1992,N_1885);
nand U2194 (N_2194,N_1810,N_1808);
nor U2195 (N_2195,N_1910,N_1868);
and U2196 (N_2196,N_1967,N_1931);
nand U2197 (N_2197,N_1862,N_1868);
nand U2198 (N_2198,N_1944,N_1867);
or U2199 (N_2199,N_1943,N_1914);
nand U2200 (N_2200,N_2086,N_2083);
and U2201 (N_2201,N_2134,N_2131);
nor U2202 (N_2202,N_2140,N_2172);
or U2203 (N_2203,N_2125,N_2181);
and U2204 (N_2204,N_2193,N_2057);
and U2205 (N_2205,N_2069,N_2046);
or U2206 (N_2206,N_2144,N_2042);
nand U2207 (N_2207,N_2010,N_2038);
and U2208 (N_2208,N_2080,N_2154);
nor U2209 (N_2209,N_2074,N_2106);
nand U2210 (N_2210,N_2148,N_2076);
and U2211 (N_2211,N_2009,N_2008);
nor U2212 (N_2212,N_2102,N_2070);
nor U2213 (N_2213,N_2097,N_2081);
nor U2214 (N_2214,N_2177,N_2019);
nand U2215 (N_2215,N_2068,N_2091);
or U2216 (N_2216,N_2045,N_2136);
nor U2217 (N_2217,N_2088,N_2151);
nor U2218 (N_2218,N_2037,N_2049);
nor U2219 (N_2219,N_2174,N_2165);
and U2220 (N_2220,N_2107,N_2061);
nand U2221 (N_2221,N_2022,N_2066);
or U2222 (N_2222,N_2028,N_2122);
nor U2223 (N_2223,N_2043,N_2155);
nand U2224 (N_2224,N_2002,N_2075);
or U2225 (N_2225,N_2011,N_2173);
nor U2226 (N_2226,N_2127,N_2183);
nor U2227 (N_2227,N_2157,N_2179);
and U2228 (N_2228,N_2176,N_2040);
or U2229 (N_2229,N_2044,N_2099);
and U2230 (N_2230,N_2032,N_2185);
and U2231 (N_2231,N_2164,N_2034);
or U2232 (N_2232,N_2138,N_2166);
and U2233 (N_2233,N_2167,N_2189);
and U2234 (N_2234,N_2023,N_2146);
or U2235 (N_2235,N_2039,N_2014);
and U2236 (N_2236,N_2192,N_2145);
nor U2237 (N_2237,N_2143,N_2110);
nor U2238 (N_2238,N_2000,N_2051);
or U2239 (N_2239,N_2082,N_2047);
and U2240 (N_2240,N_2089,N_2194);
and U2241 (N_2241,N_2058,N_2115);
xor U2242 (N_2242,N_2162,N_2120);
nand U2243 (N_2243,N_2033,N_2123);
or U2244 (N_2244,N_2108,N_2053);
nand U2245 (N_2245,N_2130,N_2132);
or U2246 (N_2246,N_2142,N_2161);
or U2247 (N_2247,N_2030,N_2105);
nand U2248 (N_2248,N_2175,N_2078);
nor U2249 (N_2249,N_2139,N_2031);
or U2250 (N_2250,N_2013,N_2095);
or U2251 (N_2251,N_2187,N_2169);
and U2252 (N_2252,N_2050,N_2090);
nor U2253 (N_2253,N_2114,N_2054);
nor U2254 (N_2254,N_2060,N_2178);
nand U2255 (N_2255,N_2059,N_2133);
or U2256 (N_2256,N_2188,N_2035);
or U2257 (N_2257,N_2168,N_2190);
and U2258 (N_2258,N_2048,N_2092);
or U2259 (N_2259,N_2196,N_2093);
nand U2260 (N_2260,N_2073,N_2111);
nor U2261 (N_2261,N_2119,N_2063);
and U2262 (N_2262,N_2158,N_2087);
nor U2263 (N_2263,N_2096,N_2170);
or U2264 (N_2264,N_2017,N_2026);
and U2265 (N_2265,N_2016,N_2056);
nand U2266 (N_2266,N_2129,N_2141);
nor U2267 (N_2267,N_2184,N_2067);
nor U2268 (N_2268,N_2098,N_2171);
and U2269 (N_2269,N_2199,N_2128);
or U2270 (N_2270,N_2003,N_2197);
nand U2271 (N_2271,N_2159,N_2104);
nand U2272 (N_2272,N_2149,N_2121);
nor U2273 (N_2273,N_2079,N_2156);
or U2274 (N_2274,N_2005,N_2135);
nand U2275 (N_2275,N_2018,N_2021);
nand U2276 (N_2276,N_2094,N_2100);
and U2277 (N_2277,N_2072,N_2182);
nor U2278 (N_2278,N_2077,N_2085);
nand U2279 (N_2279,N_2065,N_2006);
or U2280 (N_2280,N_2126,N_2195);
nand U2281 (N_2281,N_2191,N_2137);
nand U2282 (N_2282,N_2198,N_2012);
nor U2283 (N_2283,N_2025,N_2180);
or U2284 (N_2284,N_2103,N_2101);
nand U2285 (N_2285,N_2150,N_2020);
or U2286 (N_2286,N_2186,N_2001);
nand U2287 (N_2287,N_2064,N_2153);
and U2288 (N_2288,N_2116,N_2027);
nand U2289 (N_2289,N_2052,N_2117);
nor U2290 (N_2290,N_2147,N_2084);
nor U2291 (N_2291,N_2124,N_2024);
nor U2292 (N_2292,N_2113,N_2163);
and U2293 (N_2293,N_2160,N_2109);
or U2294 (N_2294,N_2036,N_2007);
nor U2295 (N_2295,N_2029,N_2152);
nor U2296 (N_2296,N_2004,N_2062);
nor U2297 (N_2297,N_2112,N_2015);
nand U2298 (N_2298,N_2055,N_2041);
and U2299 (N_2299,N_2071,N_2118);
nor U2300 (N_2300,N_2084,N_2012);
nand U2301 (N_2301,N_2032,N_2000);
nor U2302 (N_2302,N_2137,N_2022);
or U2303 (N_2303,N_2030,N_2143);
nor U2304 (N_2304,N_2101,N_2172);
and U2305 (N_2305,N_2041,N_2093);
or U2306 (N_2306,N_2111,N_2054);
nor U2307 (N_2307,N_2006,N_2075);
nand U2308 (N_2308,N_2056,N_2148);
or U2309 (N_2309,N_2163,N_2107);
or U2310 (N_2310,N_2079,N_2017);
nand U2311 (N_2311,N_2192,N_2137);
or U2312 (N_2312,N_2075,N_2078);
or U2313 (N_2313,N_2035,N_2009);
or U2314 (N_2314,N_2183,N_2150);
nor U2315 (N_2315,N_2134,N_2037);
or U2316 (N_2316,N_2080,N_2081);
nand U2317 (N_2317,N_2002,N_2136);
or U2318 (N_2318,N_2094,N_2179);
and U2319 (N_2319,N_2190,N_2066);
nand U2320 (N_2320,N_2168,N_2098);
nor U2321 (N_2321,N_2007,N_2191);
and U2322 (N_2322,N_2139,N_2163);
or U2323 (N_2323,N_2099,N_2042);
nor U2324 (N_2324,N_2160,N_2133);
nor U2325 (N_2325,N_2008,N_2125);
xor U2326 (N_2326,N_2023,N_2074);
or U2327 (N_2327,N_2098,N_2189);
and U2328 (N_2328,N_2015,N_2163);
nand U2329 (N_2329,N_2002,N_2191);
nor U2330 (N_2330,N_2135,N_2074);
nand U2331 (N_2331,N_2084,N_2179);
and U2332 (N_2332,N_2068,N_2034);
nand U2333 (N_2333,N_2188,N_2159);
nor U2334 (N_2334,N_2040,N_2053);
and U2335 (N_2335,N_2082,N_2083);
nand U2336 (N_2336,N_2077,N_2117);
or U2337 (N_2337,N_2145,N_2098);
nor U2338 (N_2338,N_2150,N_2050);
or U2339 (N_2339,N_2141,N_2008);
nand U2340 (N_2340,N_2096,N_2033);
and U2341 (N_2341,N_2097,N_2160);
and U2342 (N_2342,N_2154,N_2133);
and U2343 (N_2343,N_2062,N_2045);
or U2344 (N_2344,N_2181,N_2104);
nor U2345 (N_2345,N_2073,N_2099);
and U2346 (N_2346,N_2012,N_2123);
or U2347 (N_2347,N_2040,N_2035);
and U2348 (N_2348,N_2023,N_2160);
or U2349 (N_2349,N_2113,N_2155);
or U2350 (N_2350,N_2108,N_2165);
and U2351 (N_2351,N_2081,N_2070);
nand U2352 (N_2352,N_2139,N_2141);
or U2353 (N_2353,N_2123,N_2114);
or U2354 (N_2354,N_2003,N_2166);
and U2355 (N_2355,N_2110,N_2194);
or U2356 (N_2356,N_2187,N_2197);
nor U2357 (N_2357,N_2191,N_2101);
nand U2358 (N_2358,N_2098,N_2116);
nor U2359 (N_2359,N_2179,N_2052);
nor U2360 (N_2360,N_2125,N_2119);
nor U2361 (N_2361,N_2134,N_2117);
or U2362 (N_2362,N_2070,N_2099);
and U2363 (N_2363,N_2191,N_2160);
nor U2364 (N_2364,N_2018,N_2145);
or U2365 (N_2365,N_2122,N_2188);
nand U2366 (N_2366,N_2077,N_2014);
nor U2367 (N_2367,N_2109,N_2106);
nand U2368 (N_2368,N_2044,N_2162);
nand U2369 (N_2369,N_2089,N_2127);
or U2370 (N_2370,N_2078,N_2033);
xor U2371 (N_2371,N_2125,N_2130);
nor U2372 (N_2372,N_2195,N_2163);
nor U2373 (N_2373,N_2072,N_2094);
or U2374 (N_2374,N_2098,N_2007);
and U2375 (N_2375,N_2068,N_2106);
and U2376 (N_2376,N_2003,N_2020);
and U2377 (N_2377,N_2094,N_2095);
and U2378 (N_2378,N_2094,N_2113);
and U2379 (N_2379,N_2069,N_2107);
xnor U2380 (N_2380,N_2077,N_2199);
nand U2381 (N_2381,N_2137,N_2104);
or U2382 (N_2382,N_2193,N_2145);
or U2383 (N_2383,N_2004,N_2161);
and U2384 (N_2384,N_2031,N_2161);
xnor U2385 (N_2385,N_2052,N_2132);
nor U2386 (N_2386,N_2144,N_2028);
nand U2387 (N_2387,N_2011,N_2139);
nand U2388 (N_2388,N_2085,N_2108);
xnor U2389 (N_2389,N_2117,N_2164);
nand U2390 (N_2390,N_2181,N_2110);
or U2391 (N_2391,N_2190,N_2092);
and U2392 (N_2392,N_2081,N_2157);
xor U2393 (N_2393,N_2154,N_2058);
and U2394 (N_2394,N_2021,N_2117);
and U2395 (N_2395,N_2141,N_2046);
and U2396 (N_2396,N_2194,N_2004);
nand U2397 (N_2397,N_2002,N_2127);
or U2398 (N_2398,N_2055,N_2105);
or U2399 (N_2399,N_2186,N_2170);
nor U2400 (N_2400,N_2368,N_2220);
or U2401 (N_2401,N_2363,N_2315);
nor U2402 (N_2402,N_2318,N_2258);
or U2403 (N_2403,N_2272,N_2237);
or U2404 (N_2404,N_2348,N_2388);
or U2405 (N_2405,N_2278,N_2213);
or U2406 (N_2406,N_2223,N_2352);
nand U2407 (N_2407,N_2224,N_2389);
or U2408 (N_2408,N_2302,N_2338);
nand U2409 (N_2409,N_2308,N_2303);
nand U2410 (N_2410,N_2334,N_2330);
nor U2411 (N_2411,N_2229,N_2286);
nand U2412 (N_2412,N_2214,N_2244);
nor U2413 (N_2413,N_2300,N_2319);
nor U2414 (N_2414,N_2362,N_2274);
nor U2415 (N_2415,N_2385,N_2390);
or U2416 (N_2416,N_2292,N_2290);
or U2417 (N_2417,N_2397,N_2365);
and U2418 (N_2418,N_2230,N_2251);
and U2419 (N_2419,N_2332,N_2234);
and U2420 (N_2420,N_2345,N_2297);
nor U2421 (N_2421,N_2261,N_2395);
nand U2422 (N_2422,N_2280,N_2344);
nor U2423 (N_2423,N_2283,N_2281);
nor U2424 (N_2424,N_2366,N_2265);
nand U2425 (N_2425,N_2225,N_2211);
or U2426 (N_2426,N_2341,N_2243);
nor U2427 (N_2427,N_2347,N_2396);
and U2428 (N_2428,N_2309,N_2255);
and U2429 (N_2429,N_2242,N_2228);
nand U2430 (N_2430,N_2357,N_2305);
nor U2431 (N_2431,N_2252,N_2339);
and U2432 (N_2432,N_2311,N_2316);
and U2433 (N_2433,N_2217,N_2364);
nor U2434 (N_2434,N_2267,N_2253);
nand U2435 (N_2435,N_2378,N_2288);
nor U2436 (N_2436,N_2227,N_2260);
or U2437 (N_2437,N_2247,N_2264);
nand U2438 (N_2438,N_2215,N_2371);
nand U2439 (N_2439,N_2210,N_2293);
and U2440 (N_2440,N_2329,N_2323);
nor U2441 (N_2441,N_2259,N_2337);
nor U2442 (N_2442,N_2373,N_2203);
nand U2443 (N_2443,N_2304,N_2289);
or U2444 (N_2444,N_2239,N_2209);
or U2445 (N_2445,N_2206,N_2350);
nand U2446 (N_2446,N_2353,N_2271);
nor U2447 (N_2447,N_2269,N_2296);
or U2448 (N_2448,N_2369,N_2374);
or U2449 (N_2449,N_2384,N_2355);
nand U2450 (N_2450,N_2248,N_2349);
and U2451 (N_2451,N_2226,N_2383);
xnor U2452 (N_2452,N_2273,N_2276);
nand U2453 (N_2453,N_2375,N_2301);
and U2454 (N_2454,N_2201,N_2351);
or U2455 (N_2455,N_2358,N_2336);
nor U2456 (N_2456,N_2232,N_2287);
or U2457 (N_2457,N_2222,N_2235);
or U2458 (N_2458,N_2333,N_2317);
and U2459 (N_2459,N_2246,N_2256);
nor U2460 (N_2460,N_2221,N_2327);
and U2461 (N_2461,N_2354,N_2393);
or U2462 (N_2462,N_2250,N_2331);
and U2463 (N_2463,N_2284,N_2372);
nand U2464 (N_2464,N_2240,N_2367);
and U2465 (N_2465,N_2322,N_2346);
nand U2466 (N_2466,N_2386,N_2376);
nand U2467 (N_2467,N_2277,N_2335);
or U2468 (N_2468,N_2391,N_2238);
xor U2469 (N_2469,N_2218,N_2200);
and U2470 (N_2470,N_2392,N_2266);
or U2471 (N_2471,N_2370,N_2207);
nor U2472 (N_2472,N_2325,N_2208);
nand U2473 (N_2473,N_2212,N_2342);
nor U2474 (N_2474,N_2340,N_2231);
and U2475 (N_2475,N_2306,N_2257);
or U2476 (N_2476,N_2263,N_2380);
and U2477 (N_2477,N_2328,N_2307);
or U2478 (N_2478,N_2279,N_2382);
nand U2479 (N_2479,N_2249,N_2314);
nand U2480 (N_2480,N_2275,N_2285);
and U2481 (N_2481,N_2236,N_2398);
nand U2482 (N_2482,N_2356,N_2298);
nor U2483 (N_2483,N_2262,N_2282);
xor U2484 (N_2484,N_2291,N_2294);
and U2485 (N_2485,N_2254,N_2205);
nand U2486 (N_2486,N_2359,N_2312);
or U2487 (N_2487,N_2324,N_2233);
or U2488 (N_2488,N_2202,N_2320);
or U2489 (N_2489,N_2216,N_2377);
nand U2490 (N_2490,N_2343,N_2268);
nor U2491 (N_2491,N_2360,N_2299);
nand U2492 (N_2492,N_2321,N_2310);
xor U2493 (N_2493,N_2295,N_2270);
or U2494 (N_2494,N_2313,N_2219);
and U2495 (N_2495,N_2399,N_2379);
and U2496 (N_2496,N_2204,N_2381);
and U2497 (N_2497,N_2245,N_2361);
xor U2498 (N_2498,N_2241,N_2394);
nand U2499 (N_2499,N_2326,N_2387);
nor U2500 (N_2500,N_2318,N_2332);
or U2501 (N_2501,N_2270,N_2245);
or U2502 (N_2502,N_2334,N_2388);
and U2503 (N_2503,N_2235,N_2345);
or U2504 (N_2504,N_2300,N_2236);
or U2505 (N_2505,N_2213,N_2237);
and U2506 (N_2506,N_2286,N_2396);
or U2507 (N_2507,N_2388,N_2368);
and U2508 (N_2508,N_2372,N_2233);
and U2509 (N_2509,N_2213,N_2279);
nand U2510 (N_2510,N_2335,N_2295);
and U2511 (N_2511,N_2220,N_2345);
xnor U2512 (N_2512,N_2274,N_2259);
or U2513 (N_2513,N_2315,N_2397);
nor U2514 (N_2514,N_2268,N_2250);
or U2515 (N_2515,N_2360,N_2323);
or U2516 (N_2516,N_2278,N_2261);
nor U2517 (N_2517,N_2225,N_2380);
nand U2518 (N_2518,N_2320,N_2375);
nor U2519 (N_2519,N_2252,N_2389);
or U2520 (N_2520,N_2281,N_2323);
or U2521 (N_2521,N_2277,N_2387);
and U2522 (N_2522,N_2250,N_2360);
nor U2523 (N_2523,N_2366,N_2332);
nand U2524 (N_2524,N_2353,N_2204);
nor U2525 (N_2525,N_2298,N_2352);
nor U2526 (N_2526,N_2213,N_2249);
or U2527 (N_2527,N_2271,N_2213);
nand U2528 (N_2528,N_2381,N_2319);
and U2529 (N_2529,N_2397,N_2374);
xnor U2530 (N_2530,N_2200,N_2287);
or U2531 (N_2531,N_2253,N_2204);
nand U2532 (N_2532,N_2280,N_2204);
nand U2533 (N_2533,N_2201,N_2230);
xor U2534 (N_2534,N_2399,N_2319);
nand U2535 (N_2535,N_2366,N_2267);
or U2536 (N_2536,N_2276,N_2357);
or U2537 (N_2537,N_2364,N_2368);
and U2538 (N_2538,N_2256,N_2346);
or U2539 (N_2539,N_2325,N_2206);
nand U2540 (N_2540,N_2267,N_2355);
or U2541 (N_2541,N_2230,N_2200);
and U2542 (N_2542,N_2231,N_2240);
and U2543 (N_2543,N_2387,N_2312);
nand U2544 (N_2544,N_2233,N_2371);
xor U2545 (N_2545,N_2336,N_2376);
nand U2546 (N_2546,N_2215,N_2335);
or U2547 (N_2547,N_2313,N_2288);
nor U2548 (N_2548,N_2295,N_2264);
and U2549 (N_2549,N_2379,N_2382);
or U2550 (N_2550,N_2251,N_2280);
xor U2551 (N_2551,N_2333,N_2295);
and U2552 (N_2552,N_2276,N_2230);
nand U2553 (N_2553,N_2206,N_2287);
nand U2554 (N_2554,N_2239,N_2235);
nand U2555 (N_2555,N_2305,N_2252);
xor U2556 (N_2556,N_2330,N_2272);
or U2557 (N_2557,N_2238,N_2399);
nor U2558 (N_2558,N_2238,N_2209);
or U2559 (N_2559,N_2263,N_2225);
and U2560 (N_2560,N_2382,N_2384);
or U2561 (N_2561,N_2300,N_2228);
nor U2562 (N_2562,N_2308,N_2301);
and U2563 (N_2563,N_2280,N_2356);
nand U2564 (N_2564,N_2368,N_2308);
nor U2565 (N_2565,N_2365,N_2312);
and U2566 (N_2566,N_2374,N_2389);
or U2567 (N_2567,N_2337,N_2275);
or U2568 (N_2568,N_2211,N_2298);
or U2569 (N_2569,N_2283,N_2201);
nor U2570 (N_2570,N_2277,N_2333);
or U2571 (N_2571,N_2294,N_2317);
nor U2572 (N_2572,N_2253,N_2201);
or U2573 (N_2573,N_2271,N_2398);
nor U2574 (N_2574,N_2324,N_2202);
nor U2575 (N_2575,N_2224,N_2259);
nand U2576 (N_2576,N_2219,N_2204);
nand U2577 (N_2577,N_2240,N_2343);
and U2578 (N_2578,N_2330,N_2302);
nand U2579 (N_2579,N_2243,N_2262);
nand U2580 (N_2580,N_2293,N_2332);
nor U2581 (N_2581,N_2220,N_2282);
nand U2582 (N_2582,N_2376,N_2276);
xnor U2583 (N_2583,N_2316,N_2227);
or U2584 (N_2584,N_2221,N_2219);
or U2585 (N_2585,N_2312,N_2297);
nand U2586 (N_2586,N_2343,N_2220);
nand U2587 (N_2587,N_2205,N_2299);
or U2588 (N_2588,N_2235,N_2292);
or U2589 (N_2589,N_2225,N_2231);
nor U2590 (N_2590,N_2300,N_2370);
or U2591 (N_2591,N_2345,N_2298);
and U2592 (N_2592,N_2345,N_2365);
nor U2593 (N_2593,N_2233,N_2218);
nor U2594 (N_2594,N_2356,N_2277);
nand U2595 (N_2595,N_2348,N_2332);
or U2596 (N_2596,N_2222,N_2281);
nand U2597 (N_2597,N_2240,N_2317);
and U2598 (N_2598,N_2276,N_2301);
nor U2599 (N_2599,N_2287,N_2379);
nor U2600 (N_2600,N_2525,N_2426);
or U2601 (N_2601,N_2541,N_2454);
nand U2602 (N_2602,N_2491,N_2466);
or U2603 (N_2603,N_2400,N_2515);
or U2604 (N_2604,N_2436,N_2508);
or U2605 (N_2605,N_2566,N_2536);
nand U2606 (N_2606,N_2597,N_2568);
and U2607 (N_2607,N_2527,N_2470);
and U2608 (N_2608,N_2529,N_2472);
xor U2609 (N_2609,N_2496,N_2449);
and U2610 (N_2610,N_2401,N_2517);
nand U2611 (N_2611,N_2430,N_2483);
or U2612 (N_2612,N_2547,N_2585);
and U2613 (N_2613,N_2567,N_2542);
nand U2614 (N_2614,N_2498,N_2512);
and U2615 (N_2615,N_2446,N_2482);
and U2616 (N_2616,N_2422,N_2591);
or U2617 (N_2617,N_2414,N_2576);
and U2618 (N_2618,N_2518,N_2433);
nor U2619 (N_2619,N_2501,N_2461);
nand U2620 (N_2620,N_2502,N_2505);
or U2621 (N_2621,N_2467,N_2440);
and U2622 (N_2622,N_2580,N_2459);
or U2623 (N_2623,N_2458,N_2494);
xnor U2624 (N_2624,N_2545,N_2551);
xor U2625 (N_2625,N_2549,N_2504);
nor U2626 (N_2626,N_2425,N_2444);
nand U2627 (N_2627,N_2456,N_2493);
nor U2628 (N_2628,N_2499,N_2485);
nor U2629 (N_2629,N_2521,N_2593);
nand U2630 (N_2630,N_2537,N_2445);
and U2631 (N_2631,N_2435,N_2556);
or U2632 (N_2632,N_2408,N_2579);
nand U2633 (N_2633,N_2575,N_2540);
or U2634 (N_2634,N_2477,N_2420);
nor U2635 (N_2635,N_2530,N_2571);
and U2636 (N_2636,N_2557,N_2590);
or U2637 (N_2637,N_2594,N_2492);
or U2638 (N_2638,N_2586,N_2524);
xnor U2639 (N_2639,N_2432,N_2592);
or U2640 (N_2640,N_2452,N_2487);
nor U2641 (N_2641,N_2562,N_2559);
and U2642 (N_2642,N_2506,N_2538);
nor U2643 (N_2643,N_2555,N_2564);
and U2644 (N_2644,N_2455,N_2434);
and U2645 (N_2645,N_2453,N_2463);
nor U2646 (N_2646,N_2417,N_2488);
or U2647 (N_2647,N_2429,N_2572);
nor U2648 (N_2648,N_2539,N_2413);
nand U2649 (N_2649,N_2535,N_2596);
xor U2650 (N_2650,N_2569,N_2465);
nor U2651 (N_2651,N_2489,N_2533);
or U2652 (N_2652,N_2418,N_2404);
and U2653 (N_2653,N_2577,N_2478);
and U2654 (N_2654,N_2451,N_2416);
nor U2655 (N_2655,N_2543,N_2411);
or U2656 (N_2656,N_2450,N_2469);
and U2657 (N_2657,N_2419,N_2582);
and U2658 (N_2658,N_2552,N_2481);
and U2659 (N_2659,N_2480,N_2510);
or U2660 (N_2660,N_2473,N_2513);
nor U2661 (N_2661,N_2548,N_2519);
and U2662 (N_2662,N_2428,N_2421);
nor U2663 (N_2663,N_2460,N_2439);
nand U2664 (N_2664,N_2475,N_2405);
nor U2665 (N_2665,N_2507,N_2516);
nor U2666 (N_2666,N_2442,N_2531);
nand U2667 (N_2667,N_2522,N_2570);
nand U2668 (N_2668,N_2523,N_2495);
nor U2669 (N_2669,N_2514,N_2402);
nor U2670 (N_2670,N_2500,N_2471);
or U2671 (N_2671,N_2588,N_2595);
or U2672 (N_2672,N_2520,N_2581);
or U2673 (N_2673,N_2443,N_2412);
nand U2674 (N_2674,N_2528,N_2403);
nor U2675 (N_2675,N_2550,N_2553);
nor U2676 (N_2676,N_2476,N_2589);
nand U2677 (N_2677,N_2474,N_2565);
and U2678 (N_2678,N_2438,N_2497);
and U2679 (N_2679,N_2490,N_2437);
nor U2680 (N_2680,N_2457,N_2583);
or U2681 (N_2681,N_2427,N_2598);
nand U2682 (N_2682,N_2546,N_2431);
and U2683 (N_2683,N_2486,N_2574);
or U2684 (N_2684,N_2468,N_2534);
nand U2685 (N_2685,N_2554,N_2511);
and U2686 (N_2686,N_2532,N_2558);
or U2687 (N_2687,N_2447,N_2424);
and U2688 (N_2688,N_2587,N_2406);
and U2689 (N_2689,N_2410,N_2509);
nand U2690 (N_2690,N_2423,N_2409);
or U2691 (N_2691,N_2448,N_2526);
xor U2692 (N_2692,N_2599,N_2407);
nor U2693 (N_2693,N_2462,N_2561);
and U2694 (N_2694,N_2584,N_2484);
nand U2695 (N_2695,N_2544,N_2503);
and U2696 (N_2696,N_2441,N_2415);
and U2697 (N_2697,N_2479,N_2573);
nand U2698 (N_2698,N_2578,N_2464);
and U2699 (N_2699,N_2563,N_2560);
or U2700 (N_2700,N_2591,N_2403);
nor U2701 (N_2701,N_2548,N_2420);
nor U2702 (N_2702,N_2478,N_2534);
and U2703 (N_2703,N_2515,N_2465);
nor U2704 (N_2704,N_2434,N_2462);
or U2705 (N_2705,N_2519,N_2485);
and U2706 (N_2706,N_2531,N_2599);
and U2707 (N_2707,N_2453,N_2461);
nand U2708 (N_2708,N_2483,N_2459);
nor U2709 (N_2709,N_2451,N_2423);
or U2710 (N_2710,N_2516,N_2557);
nor U2711 (N_2711,N_2586,N_2528);
nor U2712 (N_2712,N_2586,N_2440);
and U2713 (N_2713,N_2566,N_2530);
nand U2714 (N_2714,N_2583,N_2406);
nor U2715 (N_2715,N_2562,N_2548);
nand U2716 (N_2716,N_2563,N_2577);
nand U2717 (N_2717,N_2527,N_2462);
nand U2718 (N_2718,N_2405,N_2402);
or U2719 (N_2719,N_2450,N_2408);
nand U2720 (N_2720,N_2481,N_2569);
xor U2721 (N_2721,N_2531,N_2557);
and U2722 (N_2722,N_2482,N_2577);
nor U2723 (N_2723,N_2447,N_2545);
nand U2724 (N_2724,N_2536,N_2420);
and U2725 (N_2725,N_2535,N_2584);
or U2726 (N_2726,N_2476,N_2420);
and U2727 (N_2727,N_2481,N_2538);
or U2728 (N_2728,N_2573,N_2579);
or U2729 (N_2729,N_2506,N_2599);
nor U2730 (N_2730,N_2429,N_2450);
xnor U2731 (N_2731,N_2474,N_2575);
nor U2732 (N_2732,N_2451,N_2490);
nand U2733 (N_2733,N_2453,N_2412);
nor U2734 (N_2734,N_2476,N_2515);
or U2735 (N_2735,N_2429,N_2494);
and U2736 (N_2736,N_2407,N_2515);
or U2737 (N_2737,N_2477,N_2543);
and U2738 (N_2738,N_2553,N_2479);
or U2739 (N_2739,N_2500,N_2443);
nand U2740 (N_2740,N_2501,N_2420);
nand U2741 (N_2741,N_2490,N_2457);
and U2742 (N_2742,N_2506,N_2593);
or U2743 (N_2743,N_2514,N_2454);
or U2744 (N_2744,N_2526,N_2487);
nand U2745 (N_2745,N_2430,N_2582);
or U2746 (N_2746,N_2585,N_2463);
or U2747 (N_2747,N_2579,N_2562);
nor U2748 (N_2748,N_2442,N_2566);
nor U2749 (N_2749,N_2596,N_2456);
or U2750 (N_2750,N_2484,N_2477);
nand U2751 (N_2751,N_2515,N_2519);
xor U2752 (N_2752,N_2502,N_2529);
nand U2753 (N_2753,N_2452,N_2453);
and U2754 (N_2754,N_2557,N_2404);
or U2755 (N_2755,N_2565,N_2553);
and U2756 (N_2756,N_2498,N_2400);
or U2757 (N_2757,N_2521,N_2499);
and U2758 (N_2758,N_2441,N_2411);
and U2759 (N_2759,N_2415,N_2403);
nand U2760 (N_2760,N_2498,N_2524);
nor U2761 (N_2761,N_2500,N_2562);
and U2762 (N_2762,N_2476,N_2520);
or U2763 (N_2763,N_2546,N_2497);
or U2764 (N_2764,N_2464,N_2543);
or U2765 (N_2765,N_2553,N_2476);
nand U2766 (N_2766,N_2401,N_2423);
or U2767 (N_2767,N_2448,N_2573);
or U2768 (N_2768,N_2558,N_2464);
nor U2769 (N_2769,N_2477,N_2534);
or U2770 (N_2770,N_2479,N_2533);
and U2771 (N_2771,N_2583,N_2582);
or U2772 (N_2772,N_2545,N_2425);
and U2773 (N_2773,N_2598,N_2564);
xnor U2774 (N_2774,N_2553,N_2404);
and U2775 (N_2775,N_2481,N_2471);
nand U2776 (N_2776,N_2572,N_2550);
or U2777 (N_2777,N_2459,N_2529);
nor U2778 (N_2778,N_2460,N_2526);
or U2779 (N_2779,N_2584,N_2577);
xor U2780 (N_2780,N_2536,N_2436);
or U2781 (N_2781,N_2503,N_2520);
or U2782 (N_2782,N_2480,N_2454);
and U2783 (N_2783,N_2548,N_2482);
xnor U2784 (N_2784,N_2548,N_2583);
nor U2785 (N_2785,N_2411,N_2513);
nor U2786 (N_2786,N_2580,N_2591);
or U2787 (N_2787,N_2536,N_2520);
or U2788 (N_2788,N_2572,N_2546);
nor U2789 (N_2789,N_2445,N_2400);
and U2790 (N_2790,N_2586,N_2430);
or U2791 (N_2791,N_2566,N_2570);
nand U2792 (N_2792,N_2431,N_2470);
and U2793 (N_2793,N_2594,N_2588);
nor U2794 (N_2794,N_2586,N_2471);
or U2795 (N_2795,N_2587,N_2522);
or U2796 (N_2796,N_2490,N_2550);
and U2797 (N_2797,N_2592,N_2459);
nand U2798 (N_2798,N_2566,N_2403);
nor U2799 (N_2799,N_2544,N_2535);
or U2800 (N_2800,N_2718,N_2796);
nor U2801 (N_2801,N_2763,N_2742);
nor U2802 (N_2802,N_2703,N_2780);
or U2803 (N_2803,N_2707,N_2783);
or U2804 (N_2804,N_2669,N_2688);
or U2805 (N_2805,N_2690,N_2773);
nor U2806 (N_2806,N_2634,N_2680);
and U2807 (N_2807,N_2650,N_2652);
nand U2808 (N_2808,N_2691,N_2725);
nor U2809 (N_2809,N_2753,N_2750);
nor U2810 (N_2810,N_2785,N_2752);
nand U2811 (N_2811,N_2751,N_2658);
nand U2812 (N_2812,N_2789,N_2629);
nor U2813 (N_2813,N_2655,N_2611);
and U2814 (N_2814,N_2695,N_2618);
nand U2815 (N_2815,N_2661,N_2767);
nand U2816 (N_2816,N_2639,N_2673);
nor U2817 (N_2817,N_2668,N_2626);
nor U2818 (N_2818,N_2798,N_2721);
nor U2819 (N_2819,N_2744,N_2649);
nor U2820 (N_2820,N_2712,N_2714);
or U2821 (N_2821,N_2648,N_2716);
nor U2822 (N_2822,N_2698,N_2689);
nor U2823 (N_2823,N_2743,N_2719);
or U2824 (N_2824,N_2731,N_2622);
and U2825 (N_2825,N_2635,N_2694);
nor U2826 (N_2826,N_2737,N_2747);
or U2827 (N_2827,N_2665,N_2784);
and U2828 (N_2828,N_2709,N_2760);
nor U2829 (N_2829,N_2790,N_2693);
or U2830 (N_2830,N_2758,N_2617);
and U2831 (N_2831,N_2619,N_2630);
xor U2832 (N_2832,N_2706,N_2735);
xor U2833 (N_2833,N_2627,N_2779);
nor U2834 (N_2834,N_2729,N_2638);
nand U2835 (N_2835,N_2621,N_2675);
nor U2836 (N_2836,N_2614,N_2795);
xor U2837 (N_2837,N_2602,N_2624);
or U2838 (N_2838,N_2623,N_2782);
and U2839 (N_2839,N_2741,N_2781);
nand U2840 (N_2840,N_2702,N_2701);
nand U2841 (N_2841,N_2727,N_2775);
nor U2842 (N_2842,N_2757,N_2740);
or U2843 (N_2843,N_2670,N_2605);
nor U2844 (N_2844,N_2769,N_2657);
nor U2845 (N_2845,N_2771,N_2787);
or U2846 (N_2846,N_2754,N_2664);
or U2847 (N_2847,N_2733,N_2726);
nand U2848 (N_2848,N_2604,N_2765);
nand U2849 (N_2849,N_2766,N_2678);
or U2850 (N_2850,N_2609,N_2791);
nor U2851 (N_2851,N_2600,N_2660);
nor U2852 (N_2852,N_2777,N_2632);
nand U2853 (N_2853,N_2667,N_2666);
nand U2854 (N_2854,N_2794,N_2797);
or U2855 (N_2855,N_2641,N_2603);
or U2856 (N_2856,N_2713,N_2730);
nand U2857 (N_2857,N_2762,N_2736);
nand U2858 (N_2858,N_2671,N_2672);
nand U2859 (N_2859,N_2756,N_2644);
nand U2860 (N_2860,N_2633,N_2717);
nor U2861 (N_2861,N_2654,N_2749);
nand U2862 (N_2862,N_2705,N_2683);
or U2863 (N_2863,N_2734,N_2628);
nand U2864 (N_2864,N_2768,N_2776);
or U2865 (N_2865,N_2615,N_2616);
nor U2866 (N_2866,N_2636,N_2620);
or U2867 (N_2867,N_2793,N_2732);
nor U2868 (N_2868,N_2696,N_2631);
and U2869 (N_2869,N_2728,N_2662);
nand U2870 (N_2870,N_2676,N_2715);
and U2871 (N_2871,N_2608,N_2606);
or U2872 (N_2872,N_2651,N_2792);
or U2873 (N_2873,N_2612,N_2704);
nor U2874 (N_2874,N_2799,N_2748);
or U2875 (N_2875,N_2778,N_2692);
nor U2876 (N_2876,N_2640,N_2601);
xnor U2877 (N_2877,N_2761,N_2686);
nor U2878 (N_2878,N_2653,N_2674);
nand U2879 (N_2879,N_2724,N_2759);
nand U2880 (N_2880,N_2687,N_2656);
and U2881 (N_2881,N_2786,N_2625);
nand U2882 (N_2882,N_2708,N_2700);
nor U2883 (N_2883,N_2764,N_2642);
and U2884 (N_2884,N_2637,N_2723);
nor U2885 (N_2885,N_2739,N_2643);
nand U2886 (N_2886,N_2663,N_2681);
nand U2887 (N_2887,N_2699,N_2685);
nor U2888 (N_2888,N_2607,N_2745);
and U2889 (N_2889,N_2710,N_2610);
nor U2890 (N_2890,N_2697,N_2788);
and U2891 (N_2891,N_2645,N_2774);
and U2892 (N_2892,N_2646,N_2613);
nand U2893 (N_2893,N_2682,N_2711);
and U2894 (N_2894,N_2738,N_2647);
and U2895 (N_2895,N_2722,N_2770);
or U2896 (N_2896,N_2746,N_2772);
nor U2897 (N_2897,N_2720,N_2659);
nand U2898 (N_2898,N_2679,N_2684);
or U2899 (N_2899,N_2677,N_2755);
nor U2900 (N_2900,N_2734,N_2620);
nand U2901 (N_2901,N_2629,N_2632);
or U2902 (N_2902,N_2776,N_2787);
and U2903 (N_2903,N_2793,N_2674);
and U2904 (N_2904,N_2606,N_2680);
or U2905 (N_2905,N_2795,N_2714);
or U2906 (N_2906,N_2663,N_2660);
nand U2907 (N_2907,N_2732,N_2741);
and U2908 (N_2908,N_2686,N_2706);
or U2909 (N_2909,N_2681,N_2713);
and U2910 (N_2910,N_2750,N_2703);
or U2911 (N_2911,N_2716,N_2774);
nand U2912 (N_2912,N_2716,N_2714);
or U2913 (N_2913,N_2728,N_2616);
nand U2914 (N_2914,N_2600,N_2667);
and U2915 (N_2915,N_2780,N_2616);
nand U2916 (N_2916,N_2691,N_2675);
nor U2917 (N_2917,N_2702,N_2782);
or U2918 (N_2918,N_2750,N_2726);
nand U2919 (N_2919,N_2687,N_2728);
and U2920 (N_2920,N_2741,N_2690);
nor U2921 (N_2921,N_2775,N_2645);
nand U2922 (N_2922,N_2783,N_2656);
nor U2923 (N_2923,N_2617,N_2715);
nand U2924 (N_2924,N_2637,N_2743);
or U2925 (N_2925,N_2703,N_2742);
nor U2926 (N_2926,N_2729,N_2652);
nor U2927 (N_2927,N_2687,N_2665);
nand U2928 (N_2928,N_2656,N_2742);
or U2929 (N_2929,N_2759,N_2783);
or U2930 (N_2930,N_2783,N_2633);
and U2931 (N_2931,N_2715,N_2770);
xnor U2932 (N_2932,N_2683,N_2708);
nand U2933 (N_2933,N_2793,N_2788);
and U2934 (N_2934,N_2616,N_2741);
and U2935 (N_2935,N_2648,N_2737);
and U2936 (N_2936,N_2773,N_2776);
nand U2937 (N_2937,N_2619,N_2723);
and U2938 (N_2938,N_2725,N_2732);
nand U2939 (N_2939,N_2682,N_2736);
nand U2940 (N_2940,N_2735,N_2763);
nand U2941 (N_2941,N_2741,N_2618);
and U2942 (N_2942,N_2660,N_2673);
or U2943 (N_2943,N_2732,N_2606);
nor U2944 (N_2944,N_2730,N_2790);
or U2945 (N_2945,N_2606,N_2726);
and U2946 (N_2946,N_2648,N_2790);
or U2947 (N_2947,N_2712,N_2759);
or U2948 (N_2948,N_2671,N_2741);
nor U2949 (N_2949,N_2634,N_2742);
nor U2950 (N_2950,N_2654,N_2646);
and U2951 (N_2951,N_2608,N_2760);
nand U2952 (N_2952,N_2712,N_2760);
nand U2953 (N_2953,N_2787,N_2765);
nand U2954 (N_2954,N_2754,N_2744);
and U2955 (N_2955,N_2795,N_2708);
nand U2956 (N_2956,N_2652,N_2665);
nor U2957 (N_2957,N_2721,N_2620);
and U2958 (N_2958,N_2670,N_2797);
nand U2959 (N_2959,N_2710,N_2624);
nor U2960 (N_2960,N_2691,N_2667);
or U2961 (N_2961,N_2717,N_2756);
nand U2962 (N_2962,N_2699,N_2698);
nor U2963 (N_2963,N_2705,N_2623);
or U2964 (N_2964,N_2693,N_2703);
nor U2965 (N_2965,N_2632,N_2771);
nor U2966 (N_2966,N_2696,N_2742);
or U2967 (N_2967,N_2788,N_2641);
nand U2968 (N_2968,N_2693,N_2674);
or U2969 (N_2969,N_2766,N_2629);
nand U2970 (N_2970,N_2647,N_2734);
and U2971 (N_2971,N_2639,N_2620);
or U2972 (N_2972,N_2795,N_2673);
nand U2973 (N_2973,N_2669,N_2639);
nor U2974 (N_2974,N_2698,N_2748);
nor U2975 (N_2975,N_2717,N_2649);
or U2976 (N_2976,N_2642,N_2602);
and U2977 (N_2977,N_2781,N_2660);
nor U2978 (N_2978,N_2712,N_2669);
or U2979 (N_2979,N_2760,N_2742);
nor U2980 (N_2980,N_2600,N_2714);
nor U2981 (N_2981,N_2742,N_2714);
or U2982 (N_2982,N_2708,N_2735);
or U2983 (N_2983,N_2615,N_2665);
and U2984 (N_2984,N_2702,N_2751);
and U2985 (N_2985,N_2618,N_2651);
or U2986 (N_2986,N_2653,N_2737);
and U2987 (N_2987,N_2726,N_2798);
and U2988 (N_2988,N_2726,N_2609);
nand U2989 (N_2989,N_2657,N_2722);
or U2990 (N_2990,N_2791,N_2697);
nor U2991 (N_2991,N_2665,N_2656);
and U2992 (N_2992,N_2674,N_2767);
nor U2993 (N_2993,N_2704,N_2788);
nor U2994 (N_2994,N_2685,N_2793);
or U2995 (N_2995,N_2636,N_2632);
nor U2996 (N_2996,N_2616,N_2632);
and U2997 (N_2997,N_2631,N_2774);
and U2998 (N_2998,N_2763,N_2604);
nor U2999 (N_2999,N_2660,N_2785);
and UO_0 (O_0,N_2838,N_2834);
and UO_1 (O_1,N_2869,N_2857);
or UO_2 (O_2,N_2927,N_2910);
or UO_3 (O_3,N_2823,N_2862);
or UO_4 (O_4,N_2971,N_2893);
or UO_5 (O_5,N_2803,N_2955);
or UO_6 (O_6,N_2957,N_2977);
nand UO_7 (O_7,N_2839,N_2904);
nor UO_8 (O_8,N_2888,N_2921);
nand UO_9 (O_9,N_2938,N_2861);
and UO_10 (O_10,N_2917,N_2885);
or UO_11 (O_11,N_2851,N_2892);
and UO_12 (O_12,N_2867,N_2894);
or UO_13 (O_13,N_2899,N_2986);
xor UO_14 (O_14,N_2874,N_2998);
nand UO_15 (O_15,N_2972,N_2852);
nor UO_16 (O_16,N_2944,N_2808);
nand UO_17 (O_17,N_2868,N_2860);
nor UO_18 (O_18,N_2942,N_2923);
or UO_19 (O_19,N_2877,N_2984);
and UO_20 (O_20,N_2964,N_2922);
or UO_21 (O_21,N_2890,N_2876);
and UO_22 (O_22,N_2990,N_2818);
nor UO_23 (O_23,N_2928,N_2863);
and UO_24 (O_24,N_2858,N_2806);
nor UO_25 (O_25,N_2965,N_2883);
nor UO_26 (O_26,N_2833,N_2901);
nor UO_27 (O_27,N_2967,N_2845);
or UO_28 (O_28,N_2952,N_2933);
nor UO_29 (O_29,N_2994,N_2841);
and UO_30 (O_30,N_2811,N_2884);
nand UO_31 (O_31,N_2958,N_2800);
and UO_32 (O_32,N_2924,N_2988);
and UO_33 (O_33,N_2847,N_2886);
and UO_34 (O_34,N_2887,N_2875);
or UO_35 (O_35,N_2940,N_2880);
nand UO_36 (O_36,N_2912,N_2829);
nand UO_37 (O_37,N_2830,N_2827);
nand UO_38 (O_38,N_2819,N_2945);
or UO_39 (O_39,N_2956,N_2913);
nand UO_40 (O_40,N_2866,N_2812);
or UO_41 (O_41,N_2907,N_2854);
nor UO_42 (O_42,N_2960,N_2962);
nor UO_43 (O_43,N_2911,N_2934);
or UO_44 (O_44,N_2878,N_2985);
and UO_45 (O_45,N_2836,N_2936);
or UO_46 (O_46,N_2896,N_2996);
or UO_47 (O_47,N_2846,N_2973);
nor UO_48 (O_48,N_2840,N_2895);
or UO_49 (O_49,N_2932,N_2983);
nor UO_50 (O_50,N_2939,N_2935);
or UO_51 (O_51,N_2891,N_2864);
or UO_52 (O_52,N_2950,N_2816);
nand UO_53 (O_53,N_2903,N_2961);
nand UO_54 (O_54,N_2814,N_2968);
and UO_55 (O_55,N_2835,N_2954);
nor UO_56 (O_56,N_2930,N_2872);
and UO_57 (O_57,N_2809,N_2915);
or UO_58 (O_58,N_2979,N_2941);
or UO_59 (O_59,N_2970,N_2931);
or UO_60 (O_60,N_2953,N_2881);
or UO_61 (O_61,N_2995,N_2844);
nor UO_62 (O_62,N_2981,N_2825);
and UO_63 (O_63,N_2989,N_2802);
nor UO_64 (O_64,N_2870,N_2929);
nor UO_65 (O_65,N_2848,N_2871);
nor UO_66 (O_66,N_2926,N_2817);
or UO_67 (O_67,N_2991,N_2804);
nand UO_68 (O_68,N_2865,N_2916);
or UO_69 (O_69,N_2906,N_2815);
nand UO_70 (O_70,N_2855,N_2974);
and UO_71 (O_71,N_2850,N_2889);
and UO_72 (O_72,N_2997,N_2943);
nand UO_73 (O_73,N_2897,N_2807);
or UO_74 (O_74,N_2959,N_2837);
nor UO_75 (O_75,N_2882,N_2992);
and UO_76 (O_76,N_2900,N_2978);
nand UO_77 (O_77,N_2925,N_2987);
nand UO_78 (O_78,N_2937,N_2849);
nor UO_79 (O_79,N_2853,N_2976);
nand UO_80 (O_80,N_2879,N_2918);
xor UO_81 (O_81,N_2832,N_2982);
or UO_82 (O_82,N_2902,N_2905);
nor UO_83 (O_83,N_2856,N_2821);
nor UO_84 (O_84,N_2810,N_2801);
nand UO_85 (O_85,N_2909,N_2949);
or UO_86 (O_86,N_2805,N_2908);
nand UO_87 (O_87,N_2842,N_2993);
and UO_88 (O_88,N_2919,N_2914);
nand UO_89 (O_89,N_2820,N_2980);
nand UO_90 (O_90,N_2975,N_2920);
or UO_91 (O_91,N_2843,N_2859);
or UO_92 (O_92,N_2999,N_2951);
nand UO_93 (O_93,N_2898,N_2963);
nand UO_94 (O_94,N_2822,N_2831);
nor UO_95 (O_95,N_2828,N_2969);
nor UO_96 (O_96,N_2873,N_2826);
xor UO_97 (O_97,N_2813,N_2947);
or UO_98 (O_98,N_2946,N_2824);
nor UO_99 (O_99,N_2948,N_2966);
and UO_100 (O_100,N_2865,N_2803);
nand UO_101 (O_101,N_2939,N_2946);
and UO_102 (O_102,N_2935,N_2964);
nand UO_103 (O_103,N_2986,N_2941);
nor UO_104 (O_104,N_2895,N_2936);
nor UO_105 (O_105,N_2842,N_2922);
nand UO_106 (O_106,N_2836,N_2918);
nand UO_107 (O_107,N_2904,N_2975);
or UO_108 (O_108,N_2823,N_2818);
or UO_109 (O_109,N_2825,N_2912);
and UO_110 (O_110,N_2870,N_2845);
and UO_111 (O_111,N_2821,N_2975);
nor UO_112 (O_112,N_2947,N_2982);
and UO_113 (O_113,N_2823,N_2811);
nand UO_114 (O_114,N_2948,N_2864);
and UO_115 (O_115,N_2835,N_2813);
or UO_116 (O_116,N_2803,N_2893);
nor UO_117 (O_117,N_2981,N_2846);
and UO_118 (O_118,N_2875,N_2817);
nor UO_119 (O_119,N_2990,N_2919);
nand UO_120 (O_120,N_2928,N_2895);
or UO_121 (O_121,N_2956,N_2891);
nand UO_122 (O_122,N_2856,N_2888);
and UO_123 (O_123,N_2886,N_2881);
and UO_124 (O_124,N_2981,N_2805);
nand UO_125 (O_125,N_2842,N_2854);
or UO_126 (O_126,N_2954,N_2853);
nand UO_127 (O_127,N_2975,N_2868);
or UO_128 (O_128,N_2920,N_2832);
nor UO_129 (O_129,N_2978,N_2833);
and UO_130 (O_130,N_2916,N_2844);
and UO_131 (O_131,N_2942,N_2901);
and UO_132 (O_132,N_2996,N_2928);
or UO_133 (O_133,N_2876,N_2819);
and UO_134 (O_134,N_2820,N_2808);
nor UO_135 (O_135,N_2881,N_2818);
and UO_136 (O_136,N_2915,N_2892);
nand UO_137 (O_137,N_2807,N_2852);
and UO_138 (O_138,N_2951,N_2911);
nor UO_139 (O_139,N_2883,N_2819);
xor UO_140 (O_140,N_2921,N_2814);
nand UO_141 (O_141,N_2886,N_2971);
nand UO_142 (O_142,N_2857,N_2849);
nand UO_143 (O_143,N_2952,N_2847);
xor UO_144 (O_144,N_2808,N_2954);
and UO_145 (O_145,N_2897,N_2944);
and UO_146 (O_146,N_2847,N_2995);
and UO_147 (O_147,N_2826,N_2832);
or UO_148 (O_148,N_2973,N_2883);
nor UO_149 (O_149,N_2978,N_2975);
nand UO_150 (O_150,N_2818,N_2972);
or UO_151 (O_151,N_2990,N_2842);
or UO_152 (O_152,N_2852,N_2940);
and UO_153 (O_153,N_2804,N_2824);
nor UO_154 (O_154,N_2865,N_2907);
or UO_155 (O_155,N_2944,N_2998);
nor UO_156 (O_156,N_2880,N_2848);
nand UO_157 (O_157,N_2914,N_2873);
xnor UO_158 (O_158,N_2831,N_2904);
nor UO_159 (O_159,N_2918,N_2905);
nor UO_160 (O_160,N_2938,N_2929);
or UO_161 (O_161,N_2812,N_2822);
or UO_162 (O_162,N_2896,N_2862);
or UO_163 (O_163,N_2801,N_2976);
nor UO_164 (O_164,N_2982,N_2977);
nor UO_165 (O_165,N_2855,N_2913);
or UO_166 (O_166,N_2946,N_2985);
or UO_167 (O_167,N_2987,N_2849);
nand UO_168 (O_168,N_2895,N_2847);
nand UO_169 (O_169,N_2970,N_2932);
and UO_170 (O_170,N_2940,N_2887);
or UO_171 (O_171,N_2912,N_2837);
and UO_172 (O_172,N_2932,N_2927);
or UO_173 (O_173,N_2908,N_2950);
nand UO_174 (O_174,N_2813,N_2858);
or UO_175 (O_175,N_2980,N_2817);
and UO_176 (O_176,N_2968,N_2934);
nor UO_177 (O_177,N_2919,N_2833);
nand UO_178 (O_178,N_2803,N_2853);
nor UO_179 (O_179,N_2855,N_2892);
and UO_180 (O_180,N_2988,N_2818);
nor UO_181 (O_181,N_2933,N_2884);
and UO_182 (O_182,N_2938,N_2872);
nor UO_183 (O_183,N_2915,N_2985);
nand UO_184 (O_184,N_2995,N_2922);
nand UO_185 (O_185,N_2916,N_2850);
and UO_186 (O_186,N_2936,N_2832);
nand UO_187 (O_187,N_2891,N_2878);
nand UO_188 (O_188,N_2994,N_2903);
nand UO_189 (O_189,N_2941,N_2897);
or UO_190 (O_190,N_2935,N_2858);
and UO_191 (O_191,N_2924,N_2925);
nand UO_192 (O_192,N_2893,N_2953);
xnor UO_193 (O_193,N_2810,N_2933);
nand UO_194 (O_194,N_2928,N_2953);
and UO_195 (O_195,N_2819,N_2943);
or UO_196 (O_196,N_2971,N_2824);
nand UO_197 (O_197,N_2950,N_2995);
and UO_198 (O_198,N_2817,N_2979);
or UO_199 (O_199,N_2982,N_2939);
nor UO_200 (O_200,N_2845,N_2946);
nand UO_201 (O_201,N_2987,N_2901);
nand UO_202 (O_202,N_2921,N_2943);
nand UO_203 (O_203,N_2969,N_2985);
or UO_204 (O_204,N_2980,N_2964);
or UO_205 (O_205,N_2833,N_2909);
and UO_206 (O_206,N_2904,N_2902);
nand UO_207 (O_207,N_2821,N_2964);
nor UO_208 (O_208,N_2826,N_2992);
and UO_209 (O_209,N_2948,N_2958);
or UO_210 (O_210,N_2929,N_2944);
nand UO_211 (O_211,N_2890,N_2807);
nand UO_212 (O_212,N_2851,N_2994);
and UO_213 (O_213,N_2819,N_2916);
or UO_214 (O_214,N_2918,N_2832);
or UO_215 (O_215,N_2869,N_2986);
or UO_216 (O_216,N_2980,N_2909);
nand UO_217 (O_217,N_2828,N_2991);
nand UO_218 (O_218,N_2803,N_2936);
nand UO_219 (O_219,N_2977,N_2926);
and UO_220 (O_220,N_2865,N_2960);
nor UO_221 (O_221,N_2861,N_2983);
nand UO_222 (O_222,N_2840,N_2989);
or UO_223 (O_223,N_2961,N_2934);
nand UO_224 (O_224,N_2854,N_2945);
or UO_225 (O_225,N_2928,N_2830);
or UO_226 (O_226,N_2831,N_2856);
and UO_227 (O_227,N_2935,N_2848);
nand UO_228 (O_228,N_2905,N_2947);
nor UO_229 (O_229,N_2871,N_2897);
and UO_230 (O_230,N_2875,N_2908);
and UO_231 (O_231,N_2948,N_2930);
nand UO_232 (O_232,N_2942,N_2807);
or UO_233 (O_233,N_2819,N_2927);
or UO_234 (O_234,N_2971,N_2970);
and UO_235 (O_235,N_2983,N_2902);
nand UO_236 (O_236,N_2948,N_2984);
and UO_237 (O_237,N_2976,N_2809);
and UO_238 (O_238,N_2890,N_2809);
and UO_239 (O_239,N_2882,N_2844);
and UO_240 (O_240,N_2914,N_2855);
nor UO_241 (O_241,N_2830,N_2954);
and UO_242 (O_242,N_2993,N_2983);
or UO_243 (O_243,N_2856,N_2903);
nand UO_244 (O_244,N_2998,N_2827);
nand UO_245 (O_245,N_2823,N_2832);
nor UO_246 (O_246,N_2956,N_2919);
nor UO_247 (O_247,N_2865,N_2956);
nor UO_248 (O_248,N_2836,N_2869);
nand UO_249 (O_249,N_2924,N_2868);
and UO_250 (O_250,N_2924,N_2820);
and UO_251 (O_251,N_2851,N_2806);
and UO_252 (O_252,N_2919,N_2841);
and UO_253 (O_253,N_2909,N_2863);
nor UO_254 (O_254,N_2976,N_2826);
nand UO_255 (O_255,N_2925,N_2878);
or UO_256 (O_256,N_2916,N_2894);
nor UO_257 (O_257,N_2800,N_2827);
or UO_258 (O_258,N_2814,N_2903);
xor UO_259 (O_259,N_2803,N_2929);
nor UO_260 (O_260,N_2860,N_2955);
nor UO_261 (O_261,N_2882,N_2862);
nor UO_262 (O_262,N_2918,N_2842);
or UO_263 (O_263,N_2876,N_2888);
and UO_264 (O_264,N_2979,N_2800);
and UO_265 (O_265,N_2855,N_2889);
and UO_266 (O_266,N_2975,N_2993);
or UO_267 (O_267,N_2839,N_2874);
xor UO_268 (O_268,N_2955,N_2901);
and UO_269 (O_269,N_2935,N_2950);
nand UO_270 (O_270,N_2835,N_2883);
or UO_271 (O_271,N_2948,N_2942);
and UO_272 (O_272,N_2851,N_2893);
and UO_273 (O_273,N_2942,N_2861);
or UO_274 (O_274,N_2879,N_2941);
nor UO_275 (O_275,N_2932,N_2925);
or UO_276 (O_276,N_2851,N_2946);
nand UO_277 (O_277,N_2934,N_2953);
or UO_278 (O_278,N_2885,N_2866);
nor UO_279 (O_279,N_2807,N_2952);
or UO_280 (O_280,N_2922,N_2950);
nand UO_281 (O_281,N_2847,N_2902);
nand UO_282 (O_282,N_2924,N_2800);
or UO_283 (O_283,N_2825,N_2859);
nor UO_284 (O_284,N_2898,N_2852);
nor UO_285 (O_285,N_2952,N_2946);
nand UO_286 (O_286,N_2810,N_2846);
and UO_287 (O_287,N_2943,N_2949);
nand UO_288 (O_288,N_2870,N_2882);
nand UO_289 (O_289,N_2849,N_2905);
or UO_290 (O_290,N_2966,N_2927);
and UO_291 (O_291,N_2985,N_2801);
nor UO_292 (O_292,N_2916,N_2883);
nor UO_293 (O_293,N_2831,N_2957);
nor UO_294 (O_294,N_2813,N_2847);
nor UO_295 (O_295,N_2903,N_2900);
nand UO_296 (O_296,N_2872,N_2947);
and UO_297 (O_297,N_2962,N_2891);
and UO_298 (O_298,N_2912,N_2946);
nor UO_299 (O_299,N_2800,N_2899);
or UO_300 (O_300,N_2956,N_2813);
and UO_301 (O_301,N_2848,N_2868);
and UO_302 (O_302,N_2973,N_2993);
nor UO_303 (O_303,N_2914,N_2955);
and UO_304 (O_304,N_2955,N_2926);
or UO_305 (O_305,N_2967,N_2829);
and UO_306 (O_306,N_2910,N_2919);
and UO_307 (O_307,N_2940,N_2855);
nand UO_308 (O_308,N_2808,N_2873);
or UO_309 (O_309,N_2857,N_2883);
nand UO_310 (O_310,N_2926,N_2982);
nand UO_311 (O_311,N_2837,N_2871);
nor UO_312 (O_312,N_2891,N_2958);
nand UO_313 (O_313,N_2971,N_2968);
nand UO_314 (O_314,N_2817,N_2883);
nor UO_315 (O_315,N_2858,N_2851);
or UO_316 (O_316,N_2822,N_2982);
or UO_317 (O_317,N_2815,N_2818);
or UO_318 (O_318,N_2896,N_2820);
or UO_319 (O_319,N_2837,N_2993);
nand UO_320 (O_320,N_2857,N_2964);
xnor UO_321 (O_321,N_2975,N_2944);
nor UO_322 (O_322,N_2983,N_2837);
nor UO_323 (O_323,N_2922,N_2858);
or UO_324 (O_324,N_2982,N_2834);
and UO_325 (O_325,N_2807,N_2822);
nor UO_326 (O_326,N_2859,N_2910);
nand UO_327 (O_327,N_2926,N_2936);
and UO_328 (O_328,N_2972,N_2831);
and UO_329 (O_329,N_2936,N_2912);
xnor UO_330 (O_330,N_2817,N_2881);
or UO_331 (O_331,N_2964,N_2838);
or UO_332 (O_332,N_2958,N_2915);
nor UO_333 (O_333,N_2888,N_2964);
nand UO_334 (O_334,N_2810,N_2906);
nor UO_335 (O_335,N_2821,N_2929);
and UO_336 (O_336,N_2989,N_2873);
and UO_337 (O_337,N_2920,N_2817);
nor UO_338 (O_338,N_2867,N_2986);
or UO_339 (O_339,N_2906,N_2807);
nor UO_340 (O_340,N_2978,N_2822);
or UO_341 (O_341,N_2946,N_2831);
and UO_342 (O_342,N_2898,N_2967);
xnor UO_343 (O_343,N_2984,N_2972);
or UO_344 (O_344,N_2972,N_2993);
or UO_345 (O_345,N_2824,N_2868);
or UO_346 (O_346,N_2919,N_2967);
and UO_347 (O_347,N_2892,N_2968);
xor UO_348 (O_348,N_2926,N_2898);
nand UO_349 (O_349,N_2909,N_2914);
nand UO_350 (O_350,N_2848,N_2819);
nand UO_351 (O_351,N_2913,N_2914);
nand UO_352 (O_352,N_2846,N_2844);
and UO_353 (O_353,N_2844,N_2953);
nand UO_354 (O_354,N_2992,N_2827);
nand UO_355 (O_355,N_2947,N_2943);
or UO_356 (O_356,N_2853,N_2870);
nand UO_357 (O_357,N_2826,N_2821);
nor UO_358 (O_358,N_2995,N_2872);
nor UO_359 (O_359,N_2992,N_2808);
or UO_360 (O_360,N_2938,N_2804);
or UO_361 (O_361,N_2920,N_2851);
and UO_362 (O_362,N_2915,N_2859);
or UO_363 (O_363,N_2846,N_2820);
and UO_364 (O_364,N_2988,N_2917);
nand UO_365 (O_365,N_2981,N_2868);
nand UO_366 (O_366,N_2862,N_2924);
or UO_367 (O_367,N_2813,N_2988);
and UO_368 (O_368,N_2828,N_2819);
or UO_369 (O_369,N_2910,N_2825);
nor UO_370 (O_370,N_2945,N_2823);
nand UO_371 (O_371,N_2864,N_2913);
nor UO_372 (O_372,N_2864,N_2854);
nand UO_373 (O_373,N_2868,N_2810);
nor UO_374 (O_374,N_2878,N_2971);
nor UO_375 (O_375,N_2815,N_2806);
nand UO_376 (O_376,N_2920,N_2910);
or UO_377 (O_377,N_2885,N_2995);
and UO_378 (O_378,N_2860,N_2972);
or UO_379 (O_379,N_2815,N_2880);
and UO_380 (O_380,N_2806,N_2861);
nand UO_381 (O_381,N_2824,N_2877);
nand UO_382 (O_382,N_2898,N_2909);
and UO_383 (O_383,N_2992,N_2923);
and UO_384 (O_384,N_2872,N_2946);
and UO_385 (O_385,N_2984,N_2801);
nor UO_386 (O_386,N_2813,N_2974);
nor UO_387 (O_387,N_2951,N_2865);
and UO_388 (O_388,N_2996,N_2951);
or UO_389 (O_389,N_2965,N_2874);
and UO_390 (O_390,N_2881,N_2875);
nor UO_391 (O_391,N_2908,N_2853);
nor UO_392 (O_392,N_2938,N_2900);
nor UO_393 (O_393,N_2912,N_2853);
or UO_394 (O_394,N_2884,N_2891);
nor UO_395 (O_395,N_2880,N_2876);
nor UO_396 (O_396,N_2921,N_2911);
or UO_397 (O_397,N_2901,N_2906);
nand UO_398 (O_398,N_2825,N_2811);
nand UO_399 (O_399,N_2918,N_2847);
and UO_400 (O_400,N_2981,N_2953);
nor UO_401 (O_401,N_2849,N_2822);
and UO_402 (O_402,N_2975,N_2952);
and UO_403 (O_403,N_2961,N_2895);
nor UO_404 (O_404,N_2884,N_2934);
nor UO_405 (O_405,N_2917,N_2949);
or UO_406 (O_406,N_2815,N_2854);
nand UO_407 (O_407,N_2932,N_2948);
or UO_408 (O_408,N_2967,N_2861);
nand UO_409 (O_409,N_2944,N_2938);
nor UO_410 (O_410,N_2820,N_2957);
or UO_411 (O_411,N_2902,N_2883);
nand UO_412 (O_412,N_2880,N_2886);
and UO_413 (O_413,N_2906,N_2927);
nand UO_414 (O_414,N_2927,N_2823);
and UO_415 (O_415,N_2982,N_2921);
nand UO_416 (O_416,N_2866,N_2939);
and UO_417 (O_417,N_2931,N_2893);
nand UO_418 (O_418,N_2805,N_2959);
nor UO_419 (O_419,N_2926,N_2953);
and UO_420 (O_420,N_2894,N_2812);
and UO_421 (O_421,N_2804,N_2815);
nor UO_422 (O_422,N_2909,N_2939);
or UO_423 (O_423,N_2917,N_2938);
nor UO_424 (O_424,N_2982,N_2873);
nand UO_425 (O_425,N_2904,N_2915);
and UO_426 (O_426,N_2862,N_2907);
nand UO_427 (O_427,N_2805,N_2955);
xnor UO_428 (O_428,N_2800,N_2843);
or UO_429 (O_429,N_2990,N_2917);
nor UO_430 (O_430,N_2944,N_2875);
nand UO_431 (O_431,N_2812,N_2859);
nor UO_432 (O_432,N_2981,N_2923);
or UO_433 (O_433,N_2819,N_2821);
or UO_434 (O_434,N_2969,N_2805);
nand UO_435 (O_435,N_2991,N_2940);
nor UO_436 (O_436,N_2841,N_2881);
or UO_437 (O_437,N_2917,N_2891);
or UO_438 (O_438,N_2889,N_2975);
or UO_439 (O_439,N_2812,N_2961);
xnor UO_440 (O_440,N_2892,N_2909);
and UO_441 (O_441,N_2956,N_2911);
and UO_442 (O_442,N_2836,N_2887);
nand UO_443 (O_443,N_2921,N_2974);
nand UO_444 (O_444,N_2866,N_2877);
and UO_445 (O_445,N_2931,N_2942);
and UO_446 (O_446,N_2934,N_2935);
or UO_447 (O_447,N_2962,N_2827);
nor UO_448 (O_448,N_2981,N_2971);
nor UO_449 (O_449,N_2898,N_2845);
nor UO_450 (O_450,N_2987,N_2827);
or UO_451 (O_451,N_2903,N_2998);
and UO_452 (O_452,N_2850,N_2857);
or UO_453 (O_453,N_2938,N_2867);
or UO_454 (O_454,N_2810,N_2941);
or UO_455 (O_455,N_2898,N_2808);
and UO_456 (O_456,N_2842,N_2949);
and UO_457 (O_457,N_2868,N_2985);
or UO_458 (O_458,N_2988,N_2829);
or UO_459 (O_459,N_2818,N_2822);
nor UO_460 (O_460,N_2881,N_2876);
and UO_461 (O_461,N_2970,N_2818);
nand UO_462 (O_462,N_2827,N_2976);
or UO_463 (O_463,N_2935,N_2802);
or UO_464 (O_464,N_2830,N_2904);
nand UO_465 (O_465,N_2917,N_2819);
nand UO_466 (O_466,N_2807,N_2808);
xor UO_467 (O_467,N_2816,N_2969);
nand UO_468 (O_468,N_2898,N_2950);
nand UO_469 (O_469,N_2832,N_2994);
nand UO_470 (O_470,N_2927,N_2829);
nand UO_471 (O_471,N_2951,N_2929);
nand UO_472 (O_472,N_2829,N_2833);
nor UO_473 (O_473,N_2905,N_2807);
nand UO_474 (O_474,N_2831,N_2875);
and UO_475 (O_475,N_2804,N_2870);
or UO_476 (O_476,N_2941,N_2841);
nand UO_477 (O_477,N_2808,N_2825);
or UO_478 (O_478,N_2976,N_2964);
nor UO_479 (O_479,N_2975,N_2915);
nor UO_480 (O_480,N_2927,N_2937);
or UO_481 (O_481,N_2863,N_2830);
nand UO_482 (O_482,N_2932,N_2837);
and UO_483 (O_483,N_2883,N_2928);
nor UO_484 (O_484,N_2959,N_2822);
nand UO_485 (O_485,N_2806,N_2856);
or UO_486 (O_486,N_2905,N_2886);
nor UO_487 (O_487,N_2859,N_2849);
and UO_488 (O_488,N_2972,N_2813);
nand UO_489 (O_489,N_2830,N_2955);
or UO_490 (O_490,N_2955,N_2903);
nand UO_491 (O_491,N_2889,N_2800);
nor UO_492 (O_492,N_2879,N_2974);
nor UO_493 (O_493,N_2982,N_2891);
nor UO_494 (O_494,N_2866,N_2983);
xor UO_495 (O_495,N_2995,N_2835);
nand UO_496 (O_496,N_2861,N_2880);
and UO_497 (O_497,N_2819,N_2860);
and UO_498 (O_498,N_2935,N_2931);
nand UO_499 (O_499,N_2895,N_2963);
endmodule