module basic_1500_15000_2000_5_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_120,In_1174);
and U1 (N_1,In_450,In_186);
nor U2 (N_2,In_779,In_271);
nor U3 (N_3,In_1391,In_1494);
nand U4 (N_4,In_1088,In_453);
nor U5 (N_5,In_1352,In_1355);
nand U6 (N_6,In_660,In_138);
or U7 (N_7,In_1225,In_949);
nand U8 (N_8,In_1333,In_43);
and U9 (N_9,In_195,In_19);
nor U10 (N_10,In_1415,In_1222);
or U11 (N_11,In_723,In_768);
or U12 (N_12,In_284,In_1047);
nand U13 (N_13,In_833,In_164);
nand U14 (N_14,In_359,In_945);
and U15 (N_15,In_1119,In_1039);
nor U16 (N_16,In_1294,In_1090);
and U17 (N_17,In_534,In_1250);
and U18 (N_18,In_1343,In_572);
or U19 (N_19,In_648,In_889);
nand U20 (N_20,In_1334,In_313);
and U21 (N_21,In_22,In_1271);
nor U22 (N_22,In_474,In_141);
nand U23 (N_23,In_1115,In_12);
and U24 (N_24,In_375,In_1053);
or U25 (N_25,In_1441,In_123);
nand U26 (N_26,In_950,In_806);
nor U27 (N_27,In_79,In_1393);
and U28 (N_28,In_1014,In_306);
and U29 (N_29,In_214,In_1479);
nand U30 (N_30,In_300,In_1094);
or U31 (N_31,In_220,In_161);
nand U32 (N_32,In_155,In_1027);
nor U33 (N_33,In_1487,In_97);
nor U34 (N_34,In_964,In_1073);
and U35 (N_35,In_1298,In_1340);
nor U36 (N_36,In_860,In_574);
nor U37 (N_37,In_912,In_939);
nand U38 (N_38,In_63,In_1011);
nand U39 (N_39,In_490,In_1448);
and U40 (N_40,In_662,In_546);
nand U41 (N_41,In_1336,In_380);
nand U42 (N_42,In_946,In_631);
nor U43 (N_43,In_159,In_83);
nor U44 (N_44,In_1281,In_755);
and U45 (N_45,In_1378,In_551);
nand U46 (N_46,In_738,In_848);
nor U47 (N_47,In_377,In_492);
nor U48 (N_48,In_1165,In_421);
and U49 (N_49,In_248,In_625);
and U50 (N_50,In_1229,In_9);
nor U51 (N_51,In_1499,In_100);
nor U52 (N_52,In_326,In_41);
nand U53 (N_53,In_1432,In_230);
nor U54 (N_54,In_759,In_1316);
or U55 (N_55,In_1282,In_1235);
nor U56 (N_56,In_548,In_1467);
or U57 (N_57,In_980,In_854);
nor U58 (N_58,In_556,In_762);
nand U59 (N_59,In_418,In_263);
or U60 (N_60,In_711,In_91);
or U61 (N_61,In_1248,In_1244);
or U62 (N_62,In_345,In_862);
and U63 (N_63,In_700,In_480);
or U64 (N_64,In_240,In_765);
nand U65 (N_65,In_665,In_521);
or U66 (N_66,In_346,In_330);
and U67 (N_67,In_31,In_211);
nor U68 (N_68,In_259,In_325);
nand U69 (N_69,In_933,In_1347);
nor U70 (N_70,In_443,In_1029);
xnor U71 (N_71,In_301,In_1496);
or U72 (N_72,In_781,In_928);
or U73 (N_73,In_994,In_287);
and U74 (N_74,In_1255,In_72);
nor U75 (N_75,In_793,In_1149);
and U76 (N_76,In_1163,In_469);
nand U77 (N_77,In_517,In_476);
nor U78 (N_78,In_1079,In_1230);
and U79 (N_79,In_1136,In_852);
nand U80 (N_80,In_1327,In_1262);
or U81 (N_81,In_1202,In_639);
nand U82 (N_82,In_504,In_428);
or U83 (N_83,In_1251,In_890);
and U84 (N_84,In_472,In_18);
or U85 (N_85,In_677,In_174);
nand U86 (N_86,In_1193,In_670);
and U87 (N_87,In_1356,In_508);
or U88 (N_88,In_659,In_570);
nand U89 (N_89,In_209,In_686);
nand U90 (N_90,In_1362,In_1042);
nand U91 (N_91,In_6,In_1363);
nand U92 (N_92,In_1371,In_1154);
and U93 (N_93,In_875,In_400);
and U94 (N_94,In_53,In_30);
and U95 (N_95,In_1265,In_1304);
and U96 (N_96,In_309,In_948);
and U97 (N_97,In_364,In_257);
nand U98 (N_98,In_613,In_1082);
or U99 (N_99,In_650,In_564);
nand U100 (N_100,In_1430,In_874);
and U101 (N_101,In_153,In_732);
or U102 (N_102,In_735,In_1114);
nand U103 (N_103,In_1006,In_1261);
nand U104 (N_104,In_1311,In_324);
nor U105 (N_105,In_1346,In_685);
nand U106 (N_106,In_93,In_987);
nand U107 (N_107,In_283,In_427);
and U108 (N_108,In_204,In_446);
nor U109 (N_109,In_756,In_565);
nor U110 (N_110,In_1113,In_52);
or U111 (N_111,In_498,In_1185);
nand U112 (N_112,In_185,In_541);
or U113 (N_113,In_904,In_718);
and U114 (N_114,In_1215,In_849);
and U115 (N_115,In_118,In_457);
and U116 (N_116,In_773,In_827);
nor U117 (N_117,In_839,In_661);
and U118 (N_118,In_258,In_1295);
nor U119 (N_119,In_840,In_571);
or U120 (N_120,In_266,In_1021);
nand U121 (N_121,In_1310,In_1183);
nor U122 (N_122,In_224,In_38);
and U123 (N_123,In_609,In_537);
or U124 (N_124,In_911,In_937);
nor U125 (N_125,In_432,In_1320);
and U126 (N_126,In_312,In_1314);
or U127 (N_127,In_654,In_1351);
or U128 (N_128,In_454,In_825);
nor U129 (N_129,In_178,In_903);
and U130 (N_130,In_699,In_516);
or U131 (N_131,In_1056,In_293);
or U132 (N_132,In_560,In_69);
nor U133 (N_133,In_1296,In_44);
and U134 (N_134,In_242,In_200);
and U135 (N_135,In_402,In_162);
nand U136 (N_136,In_103,In_1069);
xor U137 (N_137,In_1258,In_383);
and U138 (N_138,In_864,In_317);
and U139 (N_139,In_902,In_483);
nand U140 (N_140,In_1345,In_1300);
nand U141 (N_141,In_1043,In_1111);
nor U142 (N_142,In_447,In_1424);
nand U143 (N_143,In_857,In_462);
or U144 (N_144,In_65,In_16);
nand U145 (N_145,In_1463,In_1283);
nor U146 (N_146,In_529,In_1451);
nor U147 (N_147,In_291,In_763);
nor U148 (N_148,In_628,In_580);
and U149 (N_149,In_376,In_1481);
and U150 (N_150,In_130,In_1243);
xor U151 (N_151,In_1127,In_1278);
nand U152 (N_152,In_1161,In_286);
nand U153 (N_153,In_445,In_112);
and U154 (N_154,In_1004,In_1290);
nand U155 (N_155,In_158,In_269);
nand U156 (N_156,In_538,In_674);
nand U157 (N_157,In_28,In_1318);
nand U158 (N_158,In_202,In_481);
and U159 (N_159,In_368,In_131);
or U160 (N_160,In_1328,In_1368);
nor U161 (N_161,In_241,In_593);
and U162 (N_162,In_579,In_782);
nor U163 (N_163,In_255,In_1007);
nor U164 (N_164,In_1048,In_1405);
nor U165 (N_165,In_87,In_881);
nand U166 (N_166,In_634,In_424);
nand U167 (N_167,In_264,In_666);
nor U168 (N_168,In_789,In_129);
and U169 (N_169,In_1449,In_1096);
nor U170 (N_170,In_998,In_888);
nand U171 (N_171,In_1121,In_754);
nor U172 (N_172,In_616,In_225);
or U173 (N_173,In_254,In_362);
or U174 (N_174,In_943,In_1220);
and U175 (N_175,In_790,In_887);
nand U176 (N_176,In_1498,In_365);
nor U177 (N_177,In_468,In_1381);
and U178 (N_178,In_189,In_544);
nor U179 (N_179,In_1071,In_1459);
and U180 (N_180,In_1209,In_373);
xnor U181 (N_181,In_1471,In_1093);
nand U182 (N_182,In_1026,In_1213);
or U183 (N_183,In_250,In_1194);
nor U184 (N_184,In_1470,In_420);
nand U185 (N_185,In_1267,In_1374);
nand U186 (N_186,In_145,In_1331);
and U187 (N_187,In_81,In_29);
and U188 (N_188,In_1429,In_536);
and U189 (N_189,In_796,In_467);
xor U190 (N_190,In_414,In_619);
nand U191 (N_191,In_152,In_1342);
nor U192 (N_192,In_540,In_633);
nand U193 (N_193,In_426,In_1249);
nor U194 (N_194,In_502,In_1456);
nand U195 (N_195,In_299,In_1067);
and U196 (N_196,In_1058,In_1072);
and U197 (N_197,In_1065,In_1338);
or U198 (N_198,In_523,In_910);
or U199 (N_199,In_1354,In_231);
nand U200 (N_200,In_417,In_1190);
nor U201 (N_201,In_891,In_555);
or U202 (N_202,In_1397,In_181);
nand U203 (N_203,In_1129,In_1418);
or U204 (N_204,In_1337,In_645);
and U205 (N_205,In_1031,In_989);
nand U206 (N_206,In_1159,In_581);
nand U207 (N_207,In_1234,In_73);
nand U208 (N_208,In_505,In_689);
or U209 (N_209,In_1219,In_237);
nor U210 (N_210,In_1028,In_1153);
nor U211 (N_211,In_569,In_392);
and U212 (N_212,In_1324,In_51);
nand U213 (N_213,In_80,In_740);
xnor U214 (N_214,In_1383,In_1068);
and U215 (N_215,In_1488,In_1252);
or U216 (N_216,In_795,In_275);
and U217 (N_217,In_1126,In_378);
nor U218 (N_218,In_1086,In_456);
nand U219 (N_219,In_0,In_905);
or U220 (N_220,In_847,In_549);
or U221 (N_221,In_1232,In_696);
and U222 (N_222,In_658,In_1188);
nor U223 (N_223,In_1353,In_927);
or U224 (N_224,In_956,In_870);
nor U225 (N_225,In_1305,In_528);
or U226 (N_226,In_133,In_669);
or U227 (N_227,In_1390,In_413);
or U228 (N_228,In_853,In_1341);
nor U229 (N_229,In_146,In_461);
nand U230 (N_230,In_1382,In_58);
and U231 (N_231,In_802,In_98);
nor U232 (N_232,In_573,In_48);
nor U233 (N_233,In_422,In_1081);
and U234 (N_234,In_235,In_947);
or U235 (N_235,In_761,In_196);
nor U236 (N_236,In_1075,In_1385);
nor U237 (N_237,In_1484,In_1196);
or U238 (N_238,In_415,In_610);
nor U239 (N_239,In_205,In_558);
and U240 (N_240,In_770,In_1020);
and U241 (N_241,In_199,In_353);
and U242 (N_242,In_366,In_737);
or U243 (N_243,In_1057,In_1443);
and U244 (N_244,In_1109,In_832);
and U245 (N_245,In_75,In_919);
nand U246 (N_246,In_1016,In_1084);
nand U247 (N_247,In_812,In_997);
nor U248 (N_248,In_338,In_501);
and U249 (N_249,In_1034,In_403);
nor U250 (N_250,In_530,In_692);
and U251 (N_251,In_668,In_1203);
nor U252 (N_252,In_34,In_535);
nand U253 (N_253,In_622,In_705);
nor U254 (N_254,In_783,In_217);
nand U255 (N_255,In_466,In_435);
nor U256 (N_256,In_192,In_1330);
and U257 (N_257,In_71,In_688);
nand U258 (N_258,In_958,In_627);
nor U259 (N_259,In_637,In_171);
nand U260 (N_260,In_961,In_36);
or U261 (N_261,In_1132,In_595);
and U262 (N_262,In_1308,In_869);
nand U263 (N_263,In_967,In_909);
and U264 (N_264,In_1402,In_559);
nand U265 (N_265,In_303,In_587);
nor U266 (N_266,In_68,In_355);
and U267 (N_267,In_1134,In_846);
nand U268 (N_268,In_1130,In_140);
nor U269 (N_269,In_751,In_1366);
and U270 (N_270,In_621,In_369);
nor U271 (N_271,In_1259,In_465);
nor U272 (N_272,In_234,In_819);
nand U273 (N_273,In_412,In_632);
or U274 (N_274,In_704,In_391);
nand U275 (N_275,In_942,In_1214);
nor U276 (N_276,In_289,In_682);
nand U277 (N_277,In_1399,In_107);
and U278 (N_278,In_1135,In_298);
nand U279 (N_279,In_267,In_13);
nand U280 (N_280,In_894,In_1005);
xor U281 (N_281,In_354,In_143);
or U282 (N_282,In_1180,In_451);
nor U283 (N_283,In_386,In_404);
and U284 (N_284,In_1317,In_1210);
and U285 (N_285,In_794,In_256);
and U286 (N_286,In_753,In_552);
nor U287 (N_287,In_1033,In_1078);
and U288 (N_288,In_702,In_198);
nor U289 (N_289,In_104,In_1002);
or U290 (N_290,In_175,In_59);
nor U291 (N_291,In_1157,In_617);
and U292 (N_292,In_531,In_228);
and U293 (N_293,In_865,In_42);
nand U294 (N_294,In_390,In_676);
nor U295 (N_295,In_1181,In_798);
and U296 (N_296,In_803,In_216);
and U297 (N_297,In_837,In_1326);
and U298 (N_298,In_917,In_892);
or U299 (N_299,In_429,In_343);
nor U300 (N_300,In_1401,In_742);
or U301 (N_301,In_1292,In_596);
or U302 (N_302,In_1365,In_776);
and U303 (N_303,In_339,In_978);
nor U304 (N_304,In_1066,In_788);
nand U305 (N_305,In_381,In_1460);
nor U306 (N_306,In_900,In_940);
or U307 (N_307,In_409,In_332);
nand U308 (N_308,In_430,In_470);
or U309 (N_309,In_814,In_419);
and U310 (N_310,In_922,In_25);
nor U311 (N_311,In_586,In_842);
and U312 (N_312,In_387,In_698);
nand U313 (N_313,In_188,In_952);
nor U314 (N_314,In_379,In_212);
nand U315 (N_315,In_410,In_1177);
and U316 (N_316,In_810,In_236);
and U317 (N_317,In_1184,In_1313);
nor U318 (N_318,In_981,In_820);
or U319 (N_319,In_485,In_1152);
or U320 (N_320,In_5,In_982);
nand U321 (N_321,In_1204,In_936);
and U322 (N_322,In_1070,In_715);
nor U323 (N_323,In_1207,In_1231);
xnor U324 (N_324,In_635,In_642);
nor U325 (N_325,In_160,In_726);
or U326 (N_326,In_1171,In_335);
nor U327 (N_327,In_868,In_1064);
nor U328 (N_328,In_1417,In_1160);
or U329 (N_329,In_1375,In_1156);
or U330 (N_330,In_582,In_589);
or U331 (N_331,In_752,In_576);
or U332 (N_332,In_1032,In_27);
and U333 (N_333,In_179,In_223);
xnor U334 (N_334,In_652,In_1436);
nor U335 (N_335,In_1307,In_506);
or U336 (N_336,In_921,In_288);
nor U337 (N_337,In_1169,In_1192);
or U338 (N_338,In_363,In_1240);
nand U339 (N_339,In_1468,In_219);
and U340 (N_340,In_1191,In_612);
and U341 (N_341,In_1427,In_482);
and U342 (N_342,In_139,In_463);
nor U343 (N_343,In_1408,In_664);
or U344 (N_344,In_487,In_327);
or U345 (N_345,In_328,In_1361);
nand U346 (N_346,In_290,In_399);
or U347 (N_347,In_17,In_898);
or U348 (N_348,In_1289,In_411);
and U349 (N_349,In_246,In_1019);
or U350 (N_350,In_1286,In_1280);
or U351 (N_351,In_1010,In_1105);
nand U352 (N_352,In_1092,In_1138);
nor U353 (N_353,In_748,In_329);
or U354 (N_354,In_1485,In_813);
or U355 (N_355,In_970,In_1198);
and U356 (N_356,In_739,In_809);
nor U357 (N_357,In_416,In_14);
nor U358 (N_358,In_90,In_88);
and U359 (N_359,In_1097,In_122);
or U360 (N_360,In_954,In_588);
and U361 (N_361,In_170,In_913);
nand U362 (N_362,In_282,In_1143);
nor U363 (N_363,In_33,In_455);
or U364 (N_364,In_137,In_1466);
and U365 (N_365,In_1473,In_1409);
nor U366 (N_366,In_342,In_273);
and U367 (N_367,In_901,In_722);
or U368 (N_368,In_1017,In_657);
nor U369 (N_369,In_106,In_274);
and U370 (N_370,In_834,In_85);
or U371 (N_371,In_268,In_969);
and U372 (N_372,In_1223,In_62);
or U373 (N_373,In_1236,In_1493);
nor U374 (N_374,In_473,In_149);
nand U375 (N_375,In_114,In_144);
nand U376 (N_376,In_1454,In_629);
or U377 (N_377,In_1414,In_360);
or U378 (N_378,In_1085,In_543);
nor U379 (N_379,In_23,In_201);
nor U380 (N_380,In_602,In_1263);
and U381 (N_381,In_1293,In_1490);
and U382 (N_382,In_163,In_21);
and U383 (N_383,In_1323,In_165);
nor U384 (N_384,In_206,In_1012);
nor U385 (N_385,In_1477,In_349);
nand U386 (N_386,In_1435,In_168);
or U387 (N_387,In_777,In_1142);
or U388 (N_388,In_984,In_64);
nor U389 (N_389,In_136,In_1049);
nand U390 (N_390,In_797,In_876);
and U391 (N_391,In_1412,In_497);
and U392 (N_392,In_1095,In_513);
or U393 (N_393,In_811,In_26);
nor U394 (N_394,In_606,In_1410);
nand U395 (N_395,In_1195,In_1238);
or U396 (N_396,In_746,In_60);
and U397 (N_397,In_959,In_843);
or U398 (N_398,In_172,In_1284);
nand U399 (N_399,In_769,In_1139);
and U400 (N_400,In_154,In_1055);
nor U401 (N_401,In_1146,In_1024);
nor U402 (N_402,In_1416,In_1377);
or U403 (N_403,In_515,In_213);
or U404 (N_404,In_1404,In_1358);
nand U405 (N_405,In_1241,In_1106);
nand U406 (N_406,In_1060,In_801);
and U407 (N_407,In_620,In_938);
nand U408 (N_408,In_232,In_532);
nand U409 (N_409,In_96,In_646);
and U410 (N_410,In_845,In_431);
nor U411 (N_411,In_641,In_229);
and U412 (N_412,In_1061,In_251);
and U413 (N_413,In_863,In_831);
nor U414 (N_414,In_486,In_215);
nand U415 (N_415,In_180,In_896);
and U416 (N_416,In_1384,In_1247);
nand U417 (N_417,In_115,In_361);
and U418 (N_418,In_1411,In_882);
nand U419 (N_419,In_1242,In_988);
and U420 (N_420,In_1254,In_563);
and U421 (N_421,In_110,In_1112);
nand U422 (N_422,In_371,In_719);
nor U423 (N_423,In_1110,In_1275);
nand U424 (N_424,In_594,In_675);
or U425 (N_425,In_1144,In_95);
nand U426 (N_426,In_1440,In_655);
nor U427 (N_427,In_1387,In_1379);
and U428 (N_428,In_1122,In_1439);
or U429 (N_429,In_1423,In_974);
nor U430 (N_430,In_434,In_1151);
nor U431 (N_431,In_193,In_1164);
or U432 (N_432,In_962,In_1475);
and U433 (N_433,In_1253,In_1155);
or U434 (N_434,In_1046,In_1117);
or U435 (N_435,In_1483,In_50);
nor U436 (N_436,In_1474,In_1125);
nand U437 (N_437,In_684,In_1348);
nor U438 (N_438,In_713,In_1118);
or U439 (N_439,In_119,In_1150);
nor U440 (N_440,In_855,In_207);
nand U441 (N_441,In_496,In_724);
and U442 (N_442,In_679,In_321);
or U443 (N_443,In_985,In_1287);
and U444 (N_444,In_693,In_452);
or U445 (N_445,In_49,In_105);
nand U446 (N_446,In_1376,In_331);
and U447 (N_447,In_640,In_1051);
and U448 (N_448,In_1217,In_1319);
nor U449 (N_449,In_436,In_310);
and U450 (N_450,In_554,In_1455);
nor U451 (N_451,In_624,In_1009);
and U452 (N_452,In_1137,In_1359);
or U453 (N_453,In_518,In_245);
nor U454 (N_454,In_54,In_1040);
nand U455 (N_455,In_604,In_673);
and U456 (N_456,In_177,In_1325);
nor U457 (N_457,In_1030,In_292);
nor U458 (N_458,In_877,In_1462);
nand U459 (N_459,In_374,In_221);
nor U460 (N_460,In_520,In_836);
nand U461 (N_461,In_1099,In_1035);
or U462 (N_462,In_1492,In_297);
nor U463 (N_463,In_1434,In_1245);
nand U464 (N_464,In_280,In_1264);
nand U465 (N_465,In_1315,In_1274);
nor U466 (N_466,In_829,In_84);
or U467 (N_467,In_598,In_396);
or U468 (N_468,In_592,In_750);
nand U469 (N_469,In_347,In_1212);
or U470 (N_470,In_191,In_663);
and U471 (N_471,In_924,In_623);
nor U472 (N_472,In_1469,In_1187);
nand U473 (N_473,In_156,In_1050);
nor U474 (N_474,In_618,In_714);
or U475 (N_475,In_1486,In_1302);
nor U476 (N_476,In_1497,In_1312);
nor U477 (N_477,In_1420,In_1025);
or U478 (N_478,In_296,In_815);
nor U479 (N_479,In_370,In_511);
nor U480 (N_480,In_1208,In_1332);
nand U481 (N_481,In_499,In_955);
nand U482 (N_482,In_1076,In_1013);
nor U483 (N_483,In_1438,In_475);
nor U484 (N_484,In_2,In_203);
or U485 (N_485,In_1260,In_389);
and U486 (N_486,In_102,In_333);
or U487 (N_487,In_858,In_1128);
nor U488 (N_488,In_340,In_393);
nor U489 (N_489,In_953,In_261);
or U490 (N_490,In_1008,In_944);
nand U491 (N_491,In_807,In_503);
nor U492 (N_492,In_758,In_11);
and U493 (N_493,In_614,In_507);
and U494 (N_494,In_440,In_1205);
or U495 (N_495,In_599,In_771);
nand U496 (N_496,In_680,In_644);
and U497 (N_497,In_733,In_965);
nor U498 (N_498,In_441,In_405);
nand U499 (N_499,In_344,In_238);
and U500 (N_500,In_1200,In_74);
or U501 (N_501,In_182,In_772);
or U502 (N_502,In_398,In_897);
nand U503 (N_503,In_262,In_822);
and U504 (N_504,In_1054,In_643);
nor U505 (N_505,In_99,In_873);
and U506 (N_506,In_861,In_1266);
and U507 (N_507,In_1458,In_871);
and U508 (N_508,In_914,In_590);
nor U509 (N_509,In_488,In_879);
and U510 (N_510,In_960,In_1489);
nand U511 (N_511,In_167,In_294);
nand U512 (N_512,In_999,In_1083);
xor U513 (N_513,In_1446,In_734);
or U514 (N_514,In_1344,In_406);
nand U515 (N_515,In_78,In_157);
and U516 (N_516,In_603,In_315);
nand U517 (N_517,In_1158,In_1445);
and U518 (N_518,In_1228,In_647);
or U519 (N_519,In_667,In_46);
nor U520 (N_520,In_731,In_966);
nand U521 (N_521,In_745,In_1178);
or U522 (N_522,In_841,In_929);
and U523 (N_523,In_526,In_1297);
or U524 (N_524,In_1421,In_709);
and U525 (N_525,In_128,In_991);
and U526 (N_526,In_336,In_1367);
or U527 (N_527,In_1224,In_741);
nand U528 (N_528,In_1380,In_484);
or U529 (N_529,In_7,In_1239);
nor U530 (N_530,In_1133,In_743);
or U531 (N_531,In_826,In_931);
nor U532 (N_532,In_1431,In_678);
or U533 (N_533,In_3,In_690);
and U534 (N_534,In_925,In_109);
nor U535 (N_535,In_649,In_1166);
or U536 (N_536,In_305,In_1179);
nand U537 (N_537,In_1162,In_562);
and U538 (N_538,In_1433,In_67);
nand U539 (N_539,In_1148,In_1059);
nand U540 (N_540,In_1172,In_1472);
and U541 (N_541,In_425,In_823);
and U542 (N_542,In_187,In_1233);
or U543 (N_543,In_983,In_111);
xor U544 (N_544,In_957,In_1413);
nand U545 (N_545,In_749,In_351);
nor U546 (N_546,In_1350,In_183);
or U547 (N_547,In_433,In_895);
nand U548 (N_548,In_885,In_394);
or U549 (N_549,In_493,In_757);
or U550 (N_550,In_77,In_1063);
nor U551 (N_551,In_1167,In_993);
nor U552 (N_552,In_1285,In_1442);
nor U553 (N_553,In_607,In_478);
and U554 (N_554,In_990,In_341);
nor U555 (N_555,In_1173,In_707);
and U556 (N_556,In_142,In_1279);
nor U557 (N_557,In_37,In_575);
and U558 (N_558,In_808,In_1386);
and U559 (N_559,In_975,In_253);
nand U560 (N_560,In_585,In_725);
and U561 (N_561,In_1372,In_730);
or U562 (N_562,In_786,In_1303);
nor U563 (N_563,In_1107,In_1357);
and U564 (N_564,In_1246,In_1182);
nor U565 (N_565,In_557,In_1476);
and U566 (N_566,In_979,In_1335);
nand U567 (N_567,In_444,In_1104);
nor U568 (N_568,In_567,In_279);
and U569 (N_569,In_787,In_367);
nor U570 (N_570,In_630,In_1211);
and U571 (N_571,In_356,In_1045);
nor U572 (N_572,In_1,In_728);
or U573 (N_573,In_884,In_886);
nand U574 (N_574,In_1395,In_1100);
or U575 (N_575,In_438,In_524);
nand U576 (N_576,In_918,In_55);
and U577 (N_577,In_716,In_1189);
nor U578 (N_578,In_584,In_82);
and U579 (N_579,In_1062,In_1452);
nand U580 (N_580,In_866,In_121);
and U581 (N_581,In_45,In_15);
and U582 (N_582,In_683,In_1392);
nand U583 (N_583,In_1322,In_509);
or U584 (N_584,In_437,In_1257);
or U585 (N_585,In_878,In_124);
nor U586 (N_586,In_1001,In_1491);
nand U587 (N_587,In_906,In_322);
and U588 (N_588,In_1176,In_314);
or U589 (N_589,In_108,In_243);
nand U590 (N_590,In_151,In_1227);
and U591 (N_591,In_687,In_583);
nor U592 (N_592,In_916,In_972);
and U593 (N_593,In_835,In_1339);
and U594 (N_594,In_126,In_304);
and U595 (N_595,In_265,In_1398);
nand U596 (N_596,In_1450,In_233);
nor U597 (N_597,In_899,In_1120);
or U598 (N_598,In_1044,In_449);
and U599 (N_599,In_10,In_920);
nor U600 (N_600,In_600,In_926);
nor U601 (N_601,In_908,In_1022);
nor U602 (N_602,In_116,In_56);
and U603 (N_603,In_514,In_1277);
or U604 (N_604,In_66,In_388);
nor U605 (N_605,In_458,In_1170);
nand U606 (N_606,In_1089,In_316);
and U607 (N_607,In_995,In_656);
nand U608 (N_608,In_1403,In_605);
nor U609 (N_609,In_117,In_1141);
or U610 (N_610,In_1147,In_1299);
or U611 (N_611,In_963,In_1422);
or U612 (N_612,In_717,In_941);
and U613 (N_613,In_1131,In_464);
and U614 (N_614,In_729,In_1364);
nand U615 (N_615,In_971,In_285);
nor U616 (N_616,In_764,In_8);
or U617 (N_617,In_1218,In_408);
nor U618 (N_618,In_397,In_850);
and U619 (N_619,In_527,In_1036);
or U620 (N_620,In_334,In_727);
nor U621 (N_621,In_1461,In_566);
or U622 (N_622,In_986,In_127);
or U623 (N_623,In_1087,In_1444);
nor U624 (N_624,In_278,In_767);
nor U625 (N_625,In_542,In_113);
nor U626 (N_626,In_494,In_976);
and U627 (N_627,In_880,In_1406);
nand U628 (N_628,In_720,In_148);
and U629 (N_629,In_281,In_358);
nand U630 (N_630,In_934,In_176);
or U631 (N_631,In_844,In_190);
nor U632 (N_632,In_577,In_1018);
nor U633 (N_633,In_1447,In_591);
nor U634 (N_634,In_311,In_681);
nand U635 (N_635,In_973,In_672);
or U636 (N_636,In_1425,In_1206);
and U637 (N_637,In_1074,In_1123);
nor U638 (N_638,In_1199,In_611);
nor U639 (N_639,In_1400,In_977);
and U640 (N_640,In_448,In_578);
or U641 (N_641,In_407,In_996);
and U642 (N_642,In_816,In_1373);
and U643 (N_643,In_495,In_308);
nor U644 (N_644,In_615,In_608);
nand U645 (N_645,In_61,In_20);
and U646 (N_646,In_276,In_691);
nand U647 (N_647,In_489,In_1480);
and U648 (N_648,In_277,In_775);
nand U649 (N_649,In_76,In_1168);
nor U650 (N_650,In_439,In_1389);
nor U651 (N_651,In_337,In_272);
nand U652 (N_652,In_553,In_135);
or U653 (N_653,In_736,In_1272);
nand U654 (N_654,In_1301,In_1197);
nor U655 (N_655,In_249,In_1495);
and U656 (N_656,In_384,In_774);
nor U657 (N_657,In_1369,In_150);
and U658 (N_658,In_477,In_1276);
xnor U659 (N_659,In_1329,In_533);
nor U660 (N_660,In_818,In_319);
nor U661 (N_661,In_1037,In_671);
and U662 (N_662,In_47,In_1077);
nand U663 (N_663,In_39,In_1428);
or U664 (N_664,In_70,In_766);
and U665 (N_665,In_694,In_459);
and U666 (N_666,In_270,In_1360);
nand U667 (N_667,In_385,In_32);
and U668 (N_668,In_94,In_348);
and U669 (N_669,In_653,In_1482);
nand U670 (N_670,In_1098,In_1140);
and U671 (N_671,In_318,In_320);
nor U672 (N_672,In_1426,In_522);
nand U673 (N_673,In_1419,In_701);
or U674 (N_674,In_780,In_1237);
or U675 (N_675,In_626,In_817);
or U676 (N_676,In_744,In_1256);
nor U677 (N_677,In_1273,In_86);
nand U678 (N_678,In_1437,In_1201);
or U679 (N_679,In_307,In_710);
and U680 (N_680,In_500,In_804);
or U681 (N_681,In_883,In_101);
nand U682 (N_682,In_792,In_352);
nand U683 (N_683,In_1175,In_1407);
nand U684 (N_684,In_800,In_184);
nand U685 (N_685,In_35,In_1306);
nand U686 (N_686,In_252,In_1103);
and U687 (N_687,In_708,In_479);
and U688 (N_688,In_510,In_785);
or U689 (N_689,In_40,In_1288);
or U690 (N_690,In_323,In_372);
and U691 (N_691,In_695,In_1186);
nor U692 (N_692,In_57,In_824);
nand U693 (N_693,In_867,In_147);
nor U694 (N_694,In_89,In_1124);
nor U695 (N_695,In_218,In_244);
and U696 (N_696,In_1221,In_907);
nand U697 (N_697,In_915,In_1041);
nor U698 (N_698,In_791,In_992);
nand U699 (N_699,In_169,In_830);
nand U700 (N_700,In_1108,In_512);
nor U701 (N_701,In_550,In_1388);
and U702 (N_702,In_132,In_525);
nor U703 (N_703,In_856,In_1464);
nand U704 (N_704,In_799,In_935);
nor U705 (N_705,In_1321,In_828);
nand U706 (N_706,In_194,In_1349);
nor U707 (N_707,In_703,In_247);
nor U708 (N_708,In_760,In_1216);
nand U709 (N_709,In_1023,In_197);
xor U710 (N_710,In_1453,In_401);
nand U711 (N_711,In_491,In_821);
nor U712 (N_712,In_357,In_539);
nand U713 (N_713,In_638,In_872);
nand U714 (N_714,In_1465,In_1457);
or U715 (N_715,In_1396,In_239);
nand U716 (N_716,In_784,In_838);
nand U717 (N_717,In_382,In_166);
or U718 (N_718,In_1478,In_134);
nor U719 (N_719,In_778,In_1270);
nor U720 (N_720,In_636,In_24);
and U721 (N_721,In_1000,In_208);
nand U722 (N_722,In_1309,In_545);
and U723 (N_723,In_302,In_173);
nor U724 (N_724,In_226,In_460);
nor U725 (N_725,In_923,In_295);
or U726 (N_726,In_547,In_4);
and U727 (N_727,In_1052,In_706);
or U728 (N_728,In_125,In_1226);
nand U729 (N_729,In_1291,In_601);
nor U730 (N_730,In_1269,In_1101);
and U731 (N_731,In_1038,In_968);
nor U732 (N_732,In_395,In_805);
or U733 (N_733,In_893,In_519);
nand U734 (N_734,In_721,In_712);
xor U735 (N_735,In_1015,In_1268);
nand U736 (N_736,In_1102,In_568);
and U737 (N_737,In_1091,In_930);
and U738 (N_738,In_260,In_1003);
nand U739 (N_739,In_92,In_697);
nand U740 (N_740,In_350,In_561);
nand U741 (N_741,In_859,In_1370);
and U742 (N_742,In_423,In_471);
and U743 (N_743,In_1080,In_651);
or U744 (N_744,In_1394,In_851);
nor U745 (N_745,In_1145,In_227);
and U746 (N_746,In_210,In_1116);
nand U747 (N_747,In_932,In_747);
nand U748 (N_748,In_597,In_442);
or U749 (N_749,In_222,In_951);
nand U750 (N_750,In_963,In_1430);
nand U751 (N_751,In_919,In_545);
nor U752 (N_752,In_1135,In_132);
nor U753 (N_753,In_1097,In_906);
nor U754 (N_754,In_481,In_722);
nand U755 (N_755,In_185,In_707);
nand U756 (N_756,In_794,In_958);
and U757 (N_757,In_837,In_1225);
nor U758 (N_758,In_1236,In_1141);
nand U759 (N_759,In_115,In_1006);
and U760 (N_760,In_263,In_151);
nand U761 (N_761,In_415,In_212);
nor U762 (N_762,In_558,In_1151);
nand U763 (N_763,In_1394,In_310);
or U764 (N_764,In_377,In_929);
nor U765 (N_765,In_440,In_1383);
nor U766 (N_766,In_822,In_85);
or U767 (N_767,In_163,In_724);
nor U768 (N_768,In_646,In_1167);
nor U769 (N_769,In_537,In_364);
nor U770 (N_770,In_1022,In_656);
nand U771 (N_771,In_984,In_1398);
nor U772 (N_772,In_405,In_648);
nor U773 (N_773,In_1016,In_603);
nand U774 (N_774,In_68,In_20);
and U775 (N_775,In_986,In_222);
or U776 (N_776,In_1190,In_231);
and U777 (N_777,In_1225,In_1144);
and U778 (N_778,In_420,In_287);
nor U779 (N_779,In_41,In_1102);
nor U780 (N_780,In_590,In_592);
or U781 (N_781,In_1311,In_1325);
nor U782 (N_782,In_850,In_961);
or U783 (N_783,In_91,In_443);
nand U784 (N_784,In_1151,In_779);
or U785 (N_785,In_1036,In_99);
nor U786 (N_786,In_1133,In_500);
nor U787 (N_787,In_236,In_337);
nor U788 (N_788,In_349,In_1419);
xnor U789 (N_789,In_648,In_1076);
nand U790 (N_790,In_1336,In_359);
nand U791 (N_791,In_486,In_330);
and U792 (N_792,In_588,In_1286);
nand U793 (N_793,In_429,In_837);
xnor U794 (N_794,In_597,In_185);
nor U795 (N_795,In_1417,In_1376);
nand U796 (N_796,In_622,In_734);
nand U797 (N_797,In_808,In_1149);
nand U798 (N_798,In_780,In_771);
nor U799 (N_799,In_1025,In_1417);
nand U800 (N_800,In_1202,In_466);
or U801 (N_801,In_712,In_51);
or U802 (N_802,In_1145,In_956);
nor U803 (N_803,In_1190,In_1096);
nand U804 (N_804,In_618,In_601);
and U805 (N_805,In_1354,In_160);
and U806 (N_806,In_1467,In_974);
nand U807 (N_807,In_83,In_1013);
nor U808 (N_808,In_1141,In_1018);
nor U809 (N_809,In_40,In_1065);
or U810 (N_810,In_896,In_5);
and U811 (N_811,In_182,In_1499);
nor U812 (N_812,In_212,In_1359);
nand U813 (N_813,In_378,In_622);
and U814 (N_814,In_218,In_1333);
nand U815 (N_815,In_910,In_1217);
or U816 (N_816,In_189,In_260);
nor U817 (N_817,In_1059,In_1221);
and U818 (N_818,In_265,In_257);
and U819 (N_819,In_407,In_336);
or U820 (N_820,In_1199,In_699);
and U821 (N_821,In_585,In_302);
nor U822 (N_822,In_1268,In_1146);
nor U823 (N_823,In_1494,In_1363);
nand U824 (N_824,In_320,In_1084);
or U825 (N_825,In_193,In_240);
and U826 (N_826,In_1221,In_1056);
and U827 (N_827,In_405,In_219);
or U828 (N_828,In_1443,In_581);
nand U829 (N_829,In_688,In_652);
and U830 (N_830,In_1345,In_403);
or U831 (N_831,In_47,In_1405);
nand U832 (N_832,In_800,In_700);
nor U833 (N_833,In_699,In_800);
and U834 (N_834,In_501,In_293);
or U835 (N_835,In_1042,In_731);
and U836 (N_836,In_1081,In_431);
and U837 (N_837,In_554,In_575);
nand U838 (N_838,In_590,In_870);
nand U839 (N_839,In_281,In_125);
and U840 (N_840,In_619,In_636);
or U841 (N_841,In_1391,In_1121);
or U842 (N_842,In_1146,In_1417);
nand U843 (N_843,In_1059,In_260);
or U844 (N_844,In_659,In_346);
nand U845 (N_845,In_901,In_91);
nand U846 (N_846,In_1461,In_1015);
or U847 (N_847,In_920,In_817);
and U848 (N_848,In_1125,In_339);
nand U849 (N_849,In_60,In_419);
nand U850 (N_850,In_483,In_316);
or U851 (N_851,In_1366,In_1369);
nand U852 (N_852,In_736,In_477);
or U853 (N_853,In_1476,In_475);
nand U854 (N_854,In_349,In_639);
nor U855 (N_855,In_1295,In_711);
nor U856 (N_856,In_196,In_39);
or U857 (N_857,In_472,In_227);
or U858 (N_858,In_1488,In_525);
and U859 (N_859,In_362,In_622);
nand U860 (N_860,In_111,In_524);
or U861 (N_861,In_317,In_936);
and U862 (N_862,In_1085,In_494);
nand U863 (N_863,In_896,In_739);
nor U864 (N_864,In_227,In_117);
xor U865 (N_865,In_938,In_1167);
nor U866 (N_866,In_273,In_978);
nand U867 (N_867,In_1089,In_355);
and U868 (N_868,In_702,In_1297);
or U869 (N_869,In_705,In_37);
nor U870 (N_870,In_1433,In_469);
and U871 (N_871,In_304,In_1467);
xnor U872 (N_872,In_882,In_1132);
nor U873 (N_873,In_387,In_1235);
and U874 (N_874,In_253,In_1300);
nor U875 (N_875,In_1137,In_175);
and U876 (N_876,In_1494,In_611);
nor U877 (N_877,In_1496,In_671);
or U878 (N_878,In_1003,In_1481);
nand U879 (N_879,In_1178,In_105);
or U880 (N_880,In_1261,In_255);
nand U881 (N_881,In_832,In_549);
or U882 (N_882,In_941,In_1301);
or U883 (N_883,In_973,In_654);
and U884 (N_884,In_639,In_590);
and U885 (N_885,In_1081,In_178);
and U886 (N_886,In_589,In_841);
or U887 (N_887,In_183,In_258);
nand U888 (N_888,In_681,In_1110);
or U889 (N_889,In_1396,In_1268);
nor U890 (N_890,In_803,In_1122);
nor U891 (N_891,In_1380,In_1311);
nor U892 (N_892,In_908,In_1222);
or U893 (N_893,In_1158,In_446);
nand U894 (N_894,In_633,In_459);
nand U895 (N_895,In_796,In_594);
nand U896 (N_896,In_183,In_910);
nand U897 (N_897,In_103,In_350);
nand U898 (N_898,In_1006,In_558);
nand U899 (N_899,In_29,In_707);
nor U900 (N_900,In_803,In_335);
and U901 (N_901,In_394,In_495);
nor U902 (N_902,In_1441,In_1141);
nor U903 (N_903,In_312,In_313);
and U904 (N_904,In_1274,In_1004);
nor U905 (N_905,In_356,In_772);
nand U906 (N_906,In_1074,In_271);
nand U907 (N_907,In_922,In_1367);
nand U908 (N_908,In_1104,In_1188);
nor U909 (N_909,In_1094,In_1397);
and U910 (N_910,In_1116,In_1050);
nor U911 (N_911,In_1000,In_542);
nand U912 (N_912,In_534,In_266);
or U913 (N_913,In_74,In_435);
nand U914 (N_914,In_1112,In_528);
or U915 (N_915,In_2,In_1448);
nand U916 (N_916,In_168,In_826);
or U917 (N_917,In_1430,In_70);
or U918 (N_918,In_647,In_958);
nand U919 (N_919,In_118,In_1471);
and U920 (N_920,In_61,In_695);
nor U921 (N_921,In_1450,In_1092);
or U922 (N_922,In_1400,In_668);
and U923 (N_923,In_1441,In_693);
nor U924 (N_924,In_1049,In_1378);
nand U925 (N_925,In_778,In_1358);
nand U926 (N_926,In_364,In_110);
and U927 (N_927,In_1050,In_597);
nor U928 (N_928,In_619,In_466);
nand U929 (N_929,In_181,In_1262);
or U930 (N_930,In_272,In_973);
or U931 (N_931,In_1333,In_1090);
nand U932 (N_932,In_1239,In_856);
or U933 (N_933,In_918,In_990);
or U934 (N_934,In_1012,In_528);
nand U935 (N_935,In_249,In_362);
and U936 (N_936,In_416,In_520);
nor U937 (N_937,In_546,In_618);
nor U938 (N_938,In_304,In_814);
and U939 (N_939,In_529,In_1146);
or U940 (N_940,In_498,In_1210);
or U941 (N_941,In_1399,In_951);
or U942 (N_942,In_406,In_1247);
nand U943 (N_943,In_977,In_24);
nor U944 (N_944,In_140,In_1074);
or U945 (N_945,In_1452,In_230);
nand U946 (N_946,In_1323,In_1080);
nor U947 (N_947,In_1166,In_627);
nor U948 (N_948,In_1385,In_231);
and U949 (N_949,In_264,In_538);
nand U950 (N_950,In_99,In_105);
nor U951 (N_951,In_1088,In_530);
nand U952 (N_952,In_594,In_329);
nand U953 (N_953,In_173,In_119);
nor U954 (N_954,In_1350,In_1132);
nor U955 (N_955,In_928,In_1309);
or U956 (N_956,In_618,In_1195);
nor U957 (N_957,In_71,In_63);
or U958 (N_958,In_504,In_934);
or U959 (N_959,In_834,In_1160);
or U960 (N_960,In_37,In_789);
nand U961 (N_961,In_456,In_1280);
nand U962 (N_962,In_188,In_822);
nor U963 (N_963,In_1397,In_226);
or U964 (N_964,In_677,In_1248);
or U965 (N_965,In_1422,In_84);
nor U966 (N_966,In_783,In_188);
nand U967 (N_967,In_565,In_237);
nand U968 (N_968,In_179,In_1198);
nor U969 (N_969,In_717,In_1447);
nand U970 (N_970,In_75,In_205);
nor U971 (N_971,In_930,In_1129);
nand U972 (N_972,In_400,In_783);
and U973 (N_973,In_547,In_702);
nor U974 (N_974,In_959,In_943);
nor U975 (N_975,In_372,In_1253);
nor U976 (N_976,In_892,In_1232);
or U977 (N_977,In_526,In_1323);
nand U978 (N_978,In_4,In_567);
and U979 (N_979,In_904,In_954);
or U980 (N_980,In_568,In_320);
nand U981 (N_981,In_83,In_663);
nor U982 (N_982,In_1264,In_80);
and U983 (N_983,In_95,In_1495);
and U984 (N_984,In_575,In_49);
nand U985 (N_985,In_1349,In_71);
nor U986 (N_986,In_1056,In_427);
nor U987 (N_987,In_942,In_446);
or U988 (N_988,In_850,In_990);
or U989 (N_989,In_1103,In_316);
nor U990 (N_990,In_1248,In_459);
nor U991 (N_991,In_641,In_600);
nor U992 (N_992,In_716,In_972);
and U993 (N_993,In_388,In_827);
nand U994 (N_994,In_1205,In_69);
nor U995 (N_995,In_1092,In_475);
or U996 (N_996,In_906,In_498);
nor U997 (N_997,In_397,In_1372);
nand U998 (N_998,In_136,In_111);
or U999 (N_999,In_168,In_1169);
and U1000 (N_1000,In_1047,In_1249);
or U1001 (N_1001,In_908,In_1390);
nand U1002 (N_1002,In_562,In_1342);
nand U1003 (N_1003,In_203,In_184);
or U1004 (N_1004,In_379,In_353);
nand U1005 (N_1005,In_947,In_1081);
and U1006 (N_1006,In_1114,In_980);
and U1007 (N_1007,In_1429,In_995);
nor U1008 (N_1008,In_1019,In_897);
xor U1009 (N_1009,In_938,In_1407);
and U1010 (N_1010,In_591,In_414);
and U1011 (N_1011,In_1265,In_1498);
and U1012 (N_1012,In_1031,In_200);
and U1013 (N_1013,In_984,In_1288);
or U1014 (N_1014,In_1401,In_518);
nand U1015 (N_1015,In_193,In_541);
or U1016 (N_1016,In_1129,In_154);
or U1017 (N_1017,In_1269,In_430);
or U1018 (N_1018,In_301,In_921);
and U1019 (N_1019,In_1229,In_521);
or U1020 (N_1020,In_995,In_650);
and U1021 (N_1021,In_357,In_844);
nand U1022 (N_1022,In_1316,In_990);
or U1023 (N_1023,In_1245,In_912);
nand U1024 (N_1024,In_1031,In_452);
nor U1025 (N_1025,In_423,In_950);
and U1026 (N_1026,In_607,In_637);
nor U1027 (N_1027,In_1399,In_290);
nand U1028 (N_1028,In_339,In_602);
nand U1029 (N_1029,In_888,In_347);
nor U1030 (N_1030,In_327,In_1444);
and U1031 (N_1031,In_381,In_422);
nand U1032 (N_1032,In_1100,In_1421);
nor U1033 (N_1033,In_43,In_225);
nor U1034 (N_1034,In_39,In_1361);
nand U1035 (N_1035,In_1052,In_809);
nand U1036 (N_1036,In_324,In_1059);
and U1037 (N_1037,In_367,In_1002);
and U1038 (N_1038,In_422,In_1089);
nor U1039 (N_1039,In_708,In_221);
or U1040 (N_1040,In_1189,In_1420);
nor U1041 (N_1041,In_1346,In_1459);
and U1042 (N_1042,In_939,In_357);
nand U1043 (N_1043,In_1049,In_1);
or U1044 (N_1044,In_204,In_713);
nand U1045 (N_1045,In_900,In_839);
xor U1046 (N_1046,In_1333,In_175);
and U1047 (N_1047,In_180,In_102);
nor U1048 (N_1048,In_1381,In_616);
and U1049 (N_1049,In_257,In_619);
and U1050 (N_1050,In_742,In_118);
nand U1051 (N_1051,In_1146,In_1411);
nor U1052 (N_1052,In_476,In_651);
nor U1053 (N_1053,In_451,In_203);
and U1054 (N_1054,In_984,In_1472);
or U1055 (N_1055,In_697,In_797);
and U1056 (N_1056,In_167,In_769);
nand U1057 (N_1057,In_978,In_496);
and U1058 (N_1058,In_1249,In_1194);
and U1059 (N_1059,In_1132,In_962);
or U1060 (N_1060,In_1235,In_1221);
and U1061 (N_1061,In_550,In_1148);
nor U1062 (N_1062,In_419,In_630);
and U1063 (N_1063,In_1009,In_4);
nand U1064 (N_1064,In_850,In_1006);
nand U1065 (N_1065,In_201,In_1193);
nand U1066 (N_1066,In_124,In_565);
nor U1067 (N_1067,In_1133,In_272);
and U1068 (N_1068,In_1454,In_1391);
and U1069 (N_1069,In_1295,In_522);
or U1070 (N_1070,In_78,In_573);
and U1071 (N_1071,In_1033,In_516);
nand U1072 (N_1072,In_1321,In_866);
and U1073 (N_1073,In_1158,In_212);
nand U1074 (N_1074,In_263,In_1360);
and U1075 (N_1075,In_1458,In_1379);
and U1076 (N_1076,In_388,In_994);
nor U1077 (N_1077,In_1045,In_467);
nor U1078 (N_1078,In_912,In_1256);
nand U1079 (N_1079,In_415,In_478);
nand U1080 (N_1080,In_728,In_1193);
and U1081 (N_1081,In_1301,In_449);
or U1082 (N_1082,In_144,In_1044);
nor U1083 (N_1083,In_679,In_1336);
nand U1084 (N_1084,In_1483,In_1102);
nor U1085 (N_1085,In_343,In_532);
nor U1086 (N_1086,In_461,In_746);
and U1087 (N_1087,In_1499,In_279);
nand U1088 (N_1088,In_736,In_632);
and U1089 (N_1089,In_251,In_477);
or U1090 (N_1090,In_1185,In_859);
nor U1091 (N_1091,In_706,In_299);
nand U1092 (N_1092,In_1355,In_475);
nor U1093 (N_1093,In_1326,In_461);
nand U1094 (N_1094,In_284,In_1049);
nor U1095 (N_1095,In_619,In_999);
or U1096 (N_1096,In_1041,In_885);
or U1097 (N_1097,In_91,In_1319);
or U1098 (N_1098,In_1449,In_483);
or U1099 (N_1099,In_1235,In_475);
or U1100 (N_1100,In_470,In_912);
or U1101 (N_1101,In_1362,In_1402);
nor U1102 (N_1102,In_1175,In_1238);
and U1103 (N_1103,In_546,In_527);
and U1104 (N_1104,In_261,In_549);
nand U1105 (N_1105,In_644,In_402);
nor U1106 (N_1106,In_1499,In_1496);
nor U1107 (N_1107,In_531,In_656);
and U1108 (N_1108,In_1008,In_1161);
and U1109 (N_1109,In_796,In_862);
nand U1110 (N_1110,In_495,In_959);
nand U1111 (N_1111,In_825,In_504);
nor U1112 (N_1112,In_56,In_836);
and U1113 (N_1113,In_128,In_1276);
nor U1114 (N_1114,In_368,In_1439);
or U1115 (N_1115,In_1402,In_818);
nor U1116 (N_1116,In_1437,In_304);
nor U1117 (N_1117,In_802,In_763);
nand U1118 (N_1118,In_1034,In_833);
nand U1119 (N_1119,In_782,In_882);
and U1120 (N_1120,In_682,In_1288);
nor U1121 (N_1121,In_295,In_735);
and U1122 (N_1122,In_871,In_1354);
nand U1123 (N_1123,In_587,In_771);
and U1124 (N_1124,In_1,In_1353);
and U1125 (N_1125,In_875,In_1113);
nor U1126 (N_1126,In_877,In_66);
nand U1127 (N_1127,In_1133,In_242);
nand U1128 (N_1128,In_1106,In_820);
or U1129 (N_1129,In_1441,In_867);
or U1130 (N_1130,In_1142,In_584);
or U1131 (N_1131,In_937,In_837);
and U1132 (N_1132,In_1036,In_6);
nor U1133 (N_1133,In_20,In_912);
nand U1134 (N_1134,In_940,In_119);
nand U1135 (N_1135,In_225,In_626);
nor U1136 (N_1136,In_246,In_25);
and U1137 (N_1137,In_657,In_301);
nand U1138 (N_1138,In_1186,In_711);
nor U1139 (N_1139,In_1486,In_468);
nand U1140 (N_1140,In_1457,In_1455);
nor U1141 (N_1141,In_1162,In_1124);
nand U1142 (N_1142,In_1289,In_10);
and U1143 (N_1143,In_30,In_1012);
or U1144 (N_1144,In_3,In_787);
nand U1145 (N_1145,In_1008,In_1357);
or U1146 (N_1146,In_852,In_247);
nand U1147 (N_1147,In_1081,In_448);
and U1148 (N_1148,In_1129,In_12);
nand U1149 (N_1149,In_1365,In_622);
or U1150 (N_1150,In_1338,In_1017);
or U1151 (N_1151,In_101,In_975);
and U1152 (N_1152,In_89,In_867);
nor U1153 (N_1153,In_1170,In_380);
nor U1154 (N_1154,In_517,In_761);
nand U1155 (N_1155,In_809,In_1053);
and U1156 (N_1156,In_137,In_166);
nand U1157 (N_1157,In_1408,In_452);
and U1158 (N_1158,In_1015,In_1367);
nor U1159 (N_1159,In_375,In_333);
nor U1160 (N_1160,In_956,In_704);
and U1161 (N_1161,In_818,In_991);
nand U1162 (N_1162,In_1388,In_755);
or U1163 (N_1163,In_254,In_622);
nor U1164 (N_1164,In_1302,In_522);
nor U1165 (N_1165,In_378,In_1011);
and U1166 (N_1166,In_391,In_485);
or U1167 (N_1167,In_1205,In_1250);
nor U1168 (N_1168,In_1230,In_453);
nand U1169 (N_1169,In_1484,In_614);
nor U1170 (N_1170,In_1194,In_560);
nor U1171 (N_1171,In_1074,In_860);
or U1172 (N_1172,In_948,In_291);
nand U1173 (N_1173,In_1441,In_1211);
or U1174 (N_1174,In_524,In_635);
nor U1175 (N_1175,In_403,In_1327);
or U1176 (N_1176,In_1002,In_1093);
xor U1177 (N_1177,In_566,In_667);
and U1178 (N_1178,In_1253,In_905);
or U1179 (N_1179,In_760,In_1333);
or U1180 (N_1180,In_720,In_941);
nor U1181 (N_1181,In_973,In_1087);
nor U1182 (N_1182,In_731,In_904);
nand U1183 (N_1183,In_1360,In_1458);
nor U1184 (N_1184,In_1215,In_1475);
and U1185 (N_1185,In_740,In_467);
nand U1186 (N_1186,In_908,In_923);
and U1187 (N_1187,In_1394,In_1292);
and U1188 (N_1188,In_391,In_1238);
nand U1189 (N_1189,In_1185,In_948);
and U1190 (N_1190,In_224,In_460);
nand U1191 (N_1191,In_132,In_201);
nor U1192 (N_1192,In_785,In_538);
or U1193 (N_1193,In_37,In_1105);
and U1194 (N_1194,In_1167,In_1322);
nand U1195 (N_1195,In_625,In_73);
nor U1196 (N_1196,In_49,In_79);
and U1197 (N_1197,In_154,In_527);
or U1198 (N_1198,In_99,In_841);
or U1199 (N_1199,In_663,In_853);
nand U1200 (N_1200,In_273,In_154);
nand U1201 (N_1201,In_1158,In_1238);
nand U1202 (N_1202,In_637,In_822);
nand U1203 (N_1203,In_1230,In_1358);
nand U1204 (N_1204,In_299,In_102);
nor U1205 (N_1205,In_1469,In_1014);
or U1206 (N_1206,In_1298,In_185);
nand U1207 (N_1207,In_669,In_942);
and U1208 (N_1208,In_647,In_1313);
and U1209 (N_1209,In_1037,In_383);
nand U1210 (N_1210,In_110,In_122);
nor U1211 (N_1211,In_1256,In_1130);
or U1212 (N_1212,In_763,In_390);
and U1213 (N_1213,In_305,In_1104);
or U1214 (N_1214,In_7,In_658);
nor U1215 (N_1215,In_1245,In_1292);
nand U1216 (N_1216,In_638,In_1119);
and U1217 (N_1217,In_235,In_985);
nor U1218 (N_1218,In_98,In_1006);
or U1219 (N_1219,In_614,In_90);
nor U1220 (N_1220,In_51,In_1351);
and U1221 (N_1221,In_30,In_970);
nand U1222 (N_1222,In_1162,In_550);
nor U1223 (N_1223,In_808,In_679);
nand U1224 (N_1224,In_833,In_294);
nor U1225 (N_1225,In_1300,In_918);
nor U1226 (N_1226,In_1000,In_692);
nand U1227 (N_1227,In_790,In_735);
nand U1228 (N_1228,In_1130,In_930);
nand U1229 (N_1229,In_564,In_1335);
nor U1230 (N_1230,In_1265,In_1336);
and U1231 (N_1231,In_1462,In_1452);
or U1232 (N_1232,In_388,In_197);
nor U1233 (N_1233,In_719,In_591);
nand U1234 (N_1234,In_173,In_641);
nor U1235 (N_1235,In_194,In_1306);
or U1236 (N_1236,In_1432,In_401);
and U1237 (N_1237,In_638,In_560);
nand U1238 (N_1238,In_842,In_1486);
nand U1239 (N_1239,In_988,In_1430);
or U1240 (N_1240,In_839,In_116);
nor U1241 (N_1241,In_413,In_93);
nand U1242 (N_1242,In_77,In_952);
and U1243 (N_1243,In_593,In_660);
nand U1244 (N_1244,In_570,In_1128);
nand U1245 (N_1245,In_203,In_983);
nand U1246 (N_1246,In_1003,In_433);
or U1247 (N_1247,In_26,In_629);
nor U1248 (N_1248,In_346,In_1362);
and U1249 (N_1249,In_770,In_1482);
nor U1250 (N_1250,In_1440,In_993);
or U1251 (N_1251,In_413,In_165);
and U1252 (N_1252,In_734,In_403);
nand U1253 (N_1253,In_534,In_787);
or U1254 (N_1254,In_261,In_1333);
or U1255 (N_1255,In_720,In_1080);
xnor U1256 (N_1256,In_226,In_1003);
nor U1257 (N_1257,In_1347,In_111);
and U1258 (N_1258,In_1390,In_423);
nand U1259 (N_1259,In_502,In_807);
nor U1260 (N_1260,In_641,In_1312);
and U1261 (N_1261,In_1010,In_697);
and U1262 (N_1262,In_1475,In_557);
or U1263 (N_1263,In_1481,In_30);
and U1264 (N_1264,In_1460,In_112);
nor U1265 (N_1265,In_783,In_1061);
and U1266 (N_1266,In_627,In_1145);
or U1267 (N_1267,In_682,In_176);
or U1268 (N_1268,In_1020,In_1359);
or U1269 (N_1269,In_1120,In_1198);
or U1270 (N_1270,In_577,In_1115);
and U1271 (N_1271,In_545,In_972);
or U1272 (N_1272,In_754,In_249);
nor U1273 (N_1273,In_333,In_1175);
nand U1274 (N_1274,In_447,In_983);
nand U1275 (N_1275,In_981,In_441);
xor U1276 (N_1276,In_1207,In_5);
or U1277 (N_1277,In_542,In_718);
nor U1278 (N_1278,In_495,In_1042);
or U1279 (N_1279,In_1431,In_751);
and U1280 (N_1280,In_895,In_72);
and U1281 (N_1281,In_557,In_704);
nand U1282 (N_1282,In_37,In_56);
nor U1283 (N_1283,In_30,In_879);
or U1284 (N_1284,In_1347,In_413);
or U1285 (N_1285,In_969,In_222);
nand U1286 (N_1286,In_0,In_994);
nand U1287 (N_1287,In_96,In_1181);
nor U1288 (N_1288,In_963,In_813);
or U1289 (N_1289,In_975,In_37);
or U1290 (N_1290,In_1106,In_1386);
nand U1291 (N_1291,In_1415,In_1295);
or U1292 (N_1292,In_414,In_1339);
nand U1293 (N_1293,In_946,In_288);
and U1294 (N_1294,In_168,In_313);
nand U1295 (N_1295,In_1337,In_578);
nor U1296 (N_1296,In_1375,In_372);
and U1297 (N_1297,In_744,In_832);
or U1298 (N_1298,In_929,In_213);
or U1299 (N_1299,In_515,In_366);
and U1300 (N_1300,In_1283,In_824);
and U1301 (N_1301,In_1012,In_136);
or U1302 (N_1302,In_437,In_766);
nand U1303 (N_1303,In_1156,In_626);
nand U1304 (N_1304,In_1221,In_102);
nor U1305 (N_1305,In_1364,In_987);
or U1306 (N_1306,In_762,In_51);
nand U1307 (N_1307,In_1493,In_431);
or U1308 (N_1308,In_1106,In_262);
and U1309 (N_1309,In_300,In_124);
or U1310 (N_1310,In_1370,In_1454);
and U1311 (N_1311,In_1475,In_605);
and U1312 (N_1312,In_8,In_855);
and U1313 (N_1313,In_1158,In_243);
nor U1314 (N_1314,In_13,In_242);
and U1315 (N_1315,In_921,In_714);
nand U1316 (N_1316,In_1210,In_897);
nor U1317 (N_1317,In_130,In_285);
and U1318 (N_1318,In_856,In_1374);
and U1319 (N_1319,In_450,In_281);
and U1320 (N_1320,In_68,In_932);
and U1321 (N_1321,In_142,In_998);
and U1322 (N_1322,In_144,In_873);
and U1323 (N_1323,In_534,In_1239);
or U1324 (N_1324,In_1341,In_1191);
nand U1325 (N_1325,In_1369,In_1215);
and U1326 (N_1326,In_962,In_556);
nor U1327 (N_1327,In_1229,In_303);
nand U1328 (N_1328,In_1300,In_1394);
nand U1329 (N_1329,In_997,In_1437);
and U1330 (N_1330,In_299,In_60);
or U1331 (N_1331,In_168,In_1010);
or U1332 (N_1332,In_476,In_76);
and U1333 (N_1333,In_1473,In_956);
nand U1334 (N_1334,In_465,In_1165);
or U1335 (N_1335,In_1117,In_182);
or U1336 (N_1336,In_155,In_635);
nor U1337 (N_1337,In_1256,In_635);
nand U1338 (N_1338,In_1205,In_1134);
and U1339 (N_1339,In_604,In_1476);
and U1340 (N_1340,In_840,In_1137);
and U1341 (N_1341,In_1121,In_533);
and U1342 (N_1342,In_239,In_670);
nor U1343 (N_1343,In_741,In_776);
and U1344 (N_1344,In_1272,In_200);
and U1345 (N_1345,In_642,In_672);
and U1346 (N_1346,In_1427,In_664);
or U1347 (N_1347,In_1352,In_381);
xor U1348 (N_1348,In_608,In_780);
nand U1349 (N_1349,In_511,In_689);
nor U1350 (N_1350,In_1450,In_227);
nor U1351 (N_1351,In_342,In_138);
nor U1352 (N_1352,In_184,In_1126);
and U1353 (N_1353,In_1317,In_921);
and U1354 (N_1354,In_1441,In_643);
or U1355 (N_1355,In_1385,In_1088);
or U1356 (N_1356,In_16,In_578);
or U1357 (N_1357,In_669,In_1305);
and U1358 (N_1358,In_573,In_154);
nor U1359 (N_1359,In_634,In_1407);
and U1360 (N_1360,In_131,In_983);
nand U1361 (N_1361,In_388,In_1125);
and U1362 (N_1362,In_1206,In_378);
nor U1363 (N_1363,In_215,In_198);
or U1364 (N_1364,In_1267,In_654);
nand U1365 (N_1365,In_1011,In_691);
and U1366 (N_1366,In_1209,In_968);
and U1367 (N_1367,In_614,In_945);
and U1368 (N_1368,In_944,In_999);
and U1369 (N_1369,In_895,In_31);
and U1370 (N_1370,In_208,In_703);
nor U1371 (N_1371,In_1426,In_886);
or U1372 (N_1372,In_642,In_1476);
and U1373 (N_1373,In_222,In_301);
and U1374 (N_1374,In_725,In_1079);
or U1375 (N_1375,In_1443,In_180);
nor U1376 (N_1376,In_1411,In_1441);
xor U1377 (N_1377,In_367,In_516);
and U1378 (N_1378,In_153,In_977);
or U1379 (N_1379,In_389,In_1166);
nor U1380 (N_1380,In_1178,In_1338);
or U1381 (N_1381,In_1156,In_1444);
and U1382 (N_1382,In_1185,In_262);
and U1383 (N_1383,In_10,In_1068);
nor U1384 (N_1384,In_100,In_398);
nand U1385 (N_1385,In_619,In_776);
nor U1386 (N_1386,In_450,In_25);
nor U1387 (N_1387,In_336,In_49);
nor U1388 (N_1388,In_1308,In_375);
and U1389 (N_1389,In_348,In_69);
and U1390 (N_1390,In_687,In_1249);
nand U1391 (N_1391,In_306,In_1001);
nand U1392 (N_1392,In_688,In_474);
nor U1393 (N_1393,In_201,In_388);
and U1394 (N_1394,In_525,In_689);
nor U1395 (N_1395,In_1049,In_1394);
nand U1396 (N_1396,In_219,In_629);
or U1397 (N_1397,In_1137,In_1418);
or U1398 (N_1398,In_365,In_769);
or U1399 (N_1399,In_508,In_375);
or U1400 (N_1400,In_1228,In_1257);
and U1401 (N_1401,In_1015,In_1428);
and U1402 (N_1402,In_691,In_593);
and U1403 (N_1403,In_459,In_1385);
and U1404 (N_1404,In_576,In_824);
or U1405 (N_1405,In_59,In_460);
and U1406 (N_1406,In_1286,In_463);
and U1407 (N_1407,In_448,In_1269);
and U1408 (N_1408,In_1030,In_114);
or U1409 (N_1409,In_1173,In_56);
nand U1410 (N_1410,In_418,In_38);
nor U1411 (N_1411,In_471,In_732);
nor U1412 (N_1412,In_1243,In_388);
or U1413 (N_1413,In_525,In_1495);
and U1414 (N_1414,In_1111,In_29);
nand U1415 (N_1415,In_599,In_1031);
and U1416 (N_1416,In_276,In_866);
nor U1417 (N_1417,In_468,In_1270);
or U1418 (N_1418,In_1013,In_154);
and U1419 (N_1419,In_921,In_1087);
nor U1420 (N_1420,In_1138,In_1421);
nor U1421 (N_1421,In_485,In_1115);
or U1422 (N_1422,In_643,In_363);
xnor U1423 (N_1423,In_1199,In_1287);
nand U1424 (N_1424,In_241,In_186);
nor U1425 (N_1425,In_656,In_877);
nand U1426 (N_1426,In_213,In_938);
and U1427 (N_1427,In_131,In_1402);
nor U1428 (N_1428,In_1449,In_1433);
and U1429 (N_1429,In_1140,In_1482);
or U1430 (N_1430,In_1198,In_1321);
or U1431 (N_1431,In_110,In_29);
and U1432 (N_1432,In_301,In_1047);
nand U1433 (N_1433,In_809,In_969);
nor U1434 (N_1434,In_905,In_1171);
nand U1435 (N_1435,In_721,In_555);
or U1436 (N_1436,In_1121,In_409);
and U1437 (N_1437,In_888,In_1075);
nand U1438 (N_1438,In_70,In_34);
or U1439 (N_1439,In_262,In_1474);
and U1440 (N_1440,In_147,In_983);
nor U1441 (N_1441,In_1022,In_185);
or U1442 (N_1442,In_609,In_1044);
nand U1443 (N_1443,In_1476,In_1335);
nor U1444 (N_1444,In_1328,In_193);
or U1445 (N_1445,In_711,In_205);
and U1446 (N_1446,In_715,In_81);
or U1447 (N_1447,In_1108,In_1420);
and U1448 (N_1448,In_178,In_1124);
nor U1449 (N_1449,In_906,In_824);
nor U1450 (N_1450,In_511,In_675);
or U1451 (N_1451,In_992,In_537);
and U1452 (N_1452,In_737,In_911);
xor U1453 (N_1453,In_1206,In_1047);
nor U1454 (N_1454,In_318,In_383);
and U1455 (N_1455,In_789,In_567);
and U1456 (N_1456,In_1384,In_815);
xor U1457 (N_1457,In_1338,In_775);
nand U1458 (N_1458,In_668,In_846);
nor U1459 (N_1459,In_878,In_777);
and U1460 (N_1460,In_745,In_1124);
or U1461 (N_1461,In_962,In_365);
or U1462 (N_1462,In_1453,In_411);
nand U1463 (N_1463,In_1494,In_424);
and U1464 (N_1464,In_125,In_1332);
and U1465 (N_1465,In_1284,In_796);
and U1466 (N_1466,In_152,In_508);
nand U1467 (N_1467,In_425,In_282);
nand U1468 (N_1468,In_35,In_400);
nor U1469 (N_1469,In_978,In_702);
or U1470 (N_1470,In_228,In_19);
or U1471 (N_1471,In_279,In_630);
nor U1472 (N_1472,In_326,In_298);
and U1473 (N_1473,In_1171,In_54);
nor U1474 (N_1474,In_1051,In_336);
nand U1475 (N_1475,In_1336,In_1128);
nand U1476 (N_1476,In_169,In_374);
nand U1477 (N_1477,In_1396,In_436);
or U1478 (N_1478,In_95,In_1334);
and U1479 (N_1479,In_1447,In_1034);
nand U1480 (N_1480,In_743,In_1394);
or U1481 (N_1481,In_1480,In_505);
and U1482 (N_1482,In_1370,In_1499);
and U1483 (N_1483,In_817,In_749);
nor U1484 (N_1484,In_20,In_1127);
nor U1485 (N_1485,In_738,In_1221);
and U1486 (N_1486,In_475,In_1039);
or U1487 (N_1487,In_365,In_1442);
and U1488 (N_1488,In_455,In_525);
and U1489 (N_1489,In_717,In_139);
nor U1490 (N_1490,In_1214,In_876);
and U1491 (N_1491,In_391,In_1427);
nand U1492 (N_1492,In_219,In_329);
nor U1493 (N_1493,In_962,In_401);
and U1494 (N_1494,In_445,In_142);
or U1495 (N_1495,In_438,In_103);
or U1496 (N_1496,In_503,In_335);
nor U1497 (N_1497,In_930,In_646);
and U1498 (N_1498,In_85,In_618);
and U1499 (N_1499,In_25,In_524);
or U1500 (N_1500,In_849,In_1068);
nand U1501 (N_1501,In_840,In_924);
and U1502 (N_1502,In_247,In_523);
and U1503 (N_1503,In_1079,In_832);
or U1504 (N_1504,In_1294,In_426);
and U1505 (N_1505,In_56,In_492);
and U1506 (N_1506,In_1476,In_1054);
nand U1507 (N_1507,In_238,In_399);
and U1508 (N_1508,In_1288,In_269);
nand U1509 (N_1509,In_198,In_167);
and U1510 (N_1510,In_987,In_1464);
and U1511 (N_1511,In_1105,In_993);
or U1512 (N_1512,In_207,In_987);
and U1513 (N_1513,In_1223,In_961);
nand U1514 (N_1514,In_1229,In_724);
or U1515 (N_1515,In_410,In_420);
nand U1516 (N_1516,In_1025,In_630);
nor U1517 (N_1517,In_736,In_1204);
or U1518 (N_1518,In_159,In_843);
nor U1519 (N_1519,In_1046,In_1319);
and U1520 (N_1520,In_847,In_790);
and U1521 (N_1521,In_601,In_401);
nand U1522 (N_1522,In_1399,In_1015);
nand U1523 (N_1523,In_752,In_85);
or U1524 (N_1524,In_553,In_1377);
and U1525 (N_1525,In_10,In_1077);
nand U1526 (N_1526,In_999,In_1074);
and U1527 (N_1527,In_1320,In_84);
and U1528 (N_1528,In_405,In_98);
or U1529 (N_1529,In_298,In_900);
nor U1530 (N_1530,In_780,In_571);
or U1531 (N_1531,In_56,In_1381);
or U1532 (N_1532,In_1235,In_964);
or U1533 (N_1533,In_1096,In_1256);
nand U1534 (N_1534,In_828,In_487);
xnor U1535 (N_1535,In_330,In_1325);
or U1536 (N_1536,In_765,In_347);
nand U1537 (N_1537,In_979,In_146);
or U1538 (N_1538,In_447,In_1384);
nand U1539 (N_1539,In_309,In_1356);
or U1540 (N_1540,In_814,In_1189);
nor U1541 (N_1541,In_713,In_1193);
nor U1542 (N_1542,In_833,In_302);
or U1543 (N_1543,In_85,In_592);
nor U1544 (N_1544,In_864,In_170);
or U1545 (N_1545,In_817,In_1109);
or U1546 (N_1546,In_464,In_619);
or U1547 (N_1547,In_573,In_1025);
or U1548 (N_1548,In_31,In_1218);
and U1549 (N_1549,In_468,In_791);
nor U1550 (N_1550,In_239,In_480);
nor U1551 (N_1551,In_1161,In_220);
and U1552 (N_1552,In_540,In_367);
nand U1553 (N_1553,In_1334,In_316);
nor U1554 (N_1554,In_771,In_1358);
and U1555 (N_1555,In_722,In_1391);
and U1556 (N_1556,In_1076,In_1264);
or U1557 (N_1557,In_1091,In_931);
and U1558 (N_1558,In_802,In_1474);
nor U1559 (N_1559,In_524,In_958);
nand U1560 (N_1560,In_673,In_1359);
and U1561 (N_1561,In_1105,In_1021);
nor U1562 (N_1562,In_1122,In_1043);
or U1563 (N_1563,In_635,In_1399);
and U1564 (N_1564,In_77,In_1357);
and U1565 (N_1565,In_1458,In_1464);
nor U1566 (N_1566,In_74,In_952);
and U1567 (N_1567,In_571,In_1028);
nor U1568 (N_1568,In_358,In_377);
and U1569 (N_1569,In_935,In_252);
and U1570 (N_1570,In_303,In_566);
nand U1571 (N_1571,In_506,In_602);
or U1572 (N_1572,In_844,In_1443);
nor U1573 (N_1573,In_22,In_591);
xnor U1574 (N_1574,In_192,In_292);
and U1575 (N_1575,In_1438,In_699);
xnor U1576 (N_1576,In_1035,In_371);
or U1577 (N_1577,In_831,In_761);
and U1578 (N_1578,In_1445,In_1206);
nor U1579 (N_1579,In_145,In_107);
nand U1580 (N_1580,In_1484,In_453);
nor U1581 (N_1581,In_1219,In_268);
and U1582 (N_1582,In_681,In_761);
and U1583 (N_1583,In_145,In_938);
nor U1584 (N_1584,In_537,In_89);
or U1585 (N_1585,In_1138,In_817);
nor U1586 (N_1586,In_859,In_674);
and U1587 (N_1587,In_1392,In_1011);
and U1588 (N_1588,In_515,In_636);
or U1589 (N_1589,In_1259,In_1479);
nand U1590 (N_1590,In_683,In_746);
nor U1591 (N_1591,In_1417,In_384);
or U1592 (N_1592,In_1300,In_469);
or U1593 (N_1593,In_1062,In_836);
or U1594 (N_1594,In_164,In_277);
nor U1595 (N_1595,In_66,In_64);
and U1596 (N_1596,In_1389,In_1171);
nand U1597 (N_1597,In_417,In_1434);
nor U1598 (N_1598,In_854,In_333);
and U1599 (N_1599,In_247,In_1484);
or U1600 (N_1600,In_531,In_8);
or U1601 (N_1601,In_149,In_140);
or U1602 (N_1602,In_805,In_314);
and U1603 (N_1603,In_944,In_1334);
and U1604 (N_1604,In_30,In_1309);
and U1605 (N_1605,In_256,In_248);
nor U1606 (N_1606,In_1051,In_575);
nand U1607 (N_1607,In_733,In_197);
nand U1608 (N_1608,In_249,In_803);
or U1609 (N_1609,In_1499,In_671);
or U1610 (N_1610,In_793,In_822);
and U1611 (N_1611,In_1380,In_771);
nand U1612 (N_1612,In_1496,In_388);
and U1613 (N_1613,In_379,In_1174);
nand U1614 (N_1614,In_734,In_651);
xor U1615 (N_1615,In_373,In_1495);
nor U1616 (N_1616,In_962,In_1226);
and U1617 (N_1617,In_943,In_1335);
and U1618 (N_1618,In_658,In_886);
or U1619 (N_1619,In_557,In_643);
and U1620 (N_1620,In_529,In_905);
nor U1621 (N_1621,In_193,In_664);
and U1622 (N_1622,In_1172,In_91);
or U1623 (N_1623,In_1482,In_1457);
nand U1624 (N_1624,In_1082,In_741);
or U1625 (N_1625,In_800,In_1449);
nand U1626 (N_1626,In_254,In_577);
or U1627 (N_1627,In_834,In_475);
nand U1628 (N_1628,In_877,In_162);
or U1629 (N_1629,In_1290,In_908);
nand U1630 (N_1630,In_638,In_679);
and U1631 (N_1631,In_196,In_1486);
nand U1632 (N_1632,In_190,In_798);
and U1633 (N_1633,In_1154,In_313);
or U1634 (N_1634,In_1304,In_382);
nand U1635 (N_1635,In_1297,In_1036);
and U1636 (N_1636,In_778,In_1413);
or U1637 (N_1637,In_1270,In_1479);
nand U1638 (N_1638,In_1419,In_823);
nor U1639 (N_1639,In_100,In_449);
nor U1640 (N_1640,In_964,In_984);
nor U1641 (N_1641,In_706,In_436);
or U1642 (N_1642,In_1062,In_426);
nor U1643 (N_1643,In_690,In_59);
and U1644 (N_1644,In_162,In_1409);
or U1645 (N_1645,In_1032,In_64);
nand U1646 (N_1646,In_1339,In_1372);
nand U1647 (N_1647,In_90,In_1211);
nand U1648 (N_1648,In_1401,In_185);
or U1649 (N_1649,In_47,In_1368);
and U1650 (N_1650,In_410,In_1174);
nor U1651 (N_1651,In_808,In_1322);
nor U1652 (N_1652,In_556,In_340);
nand U1653 (N_1653,In_1041,In_1128);
nand U1654 (N_1654,In_200,In_1147);
nor U1655 (N_1655,In_342,In_1266);
nand U1656 (N_1656,In_444,In_313);
nor U1657 (N_1657,In_798,In_33);
nor U1658 (N_1658,In_92,In_602);
nand U1659 (N_1659,In_1101,In_970);
nand U1660 (N_1660,In_50,In_657);
or U1661 (N_1661,In_758,In_1285);
or U1662 (N_1662,In_228,In_1035);
and U1663 (N_1663,In_146,In_76);
and U1664 (N_1664,In_247,In_433);
nand U1665 (N_1665,In_1317,In_18);
nand U1666 (N_1666,In_167,In_1401);
nand U1667 (N_1667,In_186,In_844);
and U1668 (N_1668,In_1024,In_1451);
nor U1669 (N_1669,In_672,In_1444);
nand U1670 (N_1670,In_320,In_362);
and U1671 (N_1671,In_401,In_1070);
or U1672 (N_1672,In_1241,In_999);
and U1673 (N_1673,In_155,In_800);
nor U1674 (N_1674,In_578,In_1260);
and U1675 (N_1675,In_587,In_324);
and U1676 (N_1676,In_892,In_496);
nor U1677 (N_1677,In_949,In_51);
nor U1678 (N_1678,In_1361,In_1142);
nor U1679 (N_1679,In_1063,In_215);
or U1680 (N_1680,In_290,In_902);
and U1681 (N_1681,In_441,In_1292);
xnor U1682 (N_1682,In_1174,In_556);
and U1683 (N_1683,In_575,In_1003);
and U1684 (N_1684,In_1024,In_492);
nor U1685 (N_1685,In_1454,In_62);
or U1686 (N_1686,In_332,In_650);
nor U1687 (N_1687,In_126,In_43);
and U1688 (N_1688,In_1086,In_1447);
or U1689 (N_1689,In_408,In_1351);
nand U1690 (N_1690,In_936,In_886);
nor U1691 (N_1691,In_1337,In_1146);
nand U1692 (N_1692,In_10,In_25);
or U1693 (N_1693,In_295,In_1007);
or U1694 (N_1694,In_406,In_407);
nand U1695 (N_1695,In_468,In_672);
nand U1696 (N_1696,In_554,In_1284);
nand U1697 (N_1697,In_1258,In_1088);
and U1698 (N_1698,In_1261,In_552);
nor U1699 (N_1699,In_1181,In_1370);
nand U1700 (N_1700,In_354,In_201);
nor U1701 (N_1701,In_1364,In_868);
nor U1702 (N_1702,In_801,In_654);
or U1703 (N_1703,In_340,In_356);
or U1704 (N_1704,In_17,In_868);
nand U1705 (N_1705,In_1329,In_1167);
nand U1706 (N_1706,In_182,In_655);
nor U1707 (N_1707,In_1459,In_994);
and U1708 (N_1708,In_244,In_192);
and U1709 (N_1709,In_328,In_760);
nand U1710 (N_1710,In_743,In_1291);
nor U1711 (N_1711,In_44,In_1162);
nor U1712 (N_1712,In_260,In_48);
or U1713 (N_1713,In_190,In_244);
or U1714 (N_1714,In_219,In_537);
nand U1715 (N_1715,In_3,In_1363);
or U1716 (N_1716,In_729,In_933);
nor U1717 (N_1717,In_766,In_122);
and U1718 (N_1718,In_932,In_470);
and U1719 (N_1719,In_1360,In_648);
nand U1720 (N_1720,In_645,In_85);
and U1721 (N_1721,In_53,In_106);
nor U1722 (N_1722,In_239,In_396);
nand U1723 (N_1723,In_1378,In_743);
nor U1724 (N_1724,In_1312,In_1095);
nand U1725 (N_1725,In_400,In_747);
nand U1726 (N_1726,In_708,In_505);
nand U1727 (N_1727,In_1360,In_86);
nand U1728 (N_1728,In_66,In_515);
nor U1729 (N_1729,In_1166,In_713);
or U1730 (N_1730,In_1118,In_999);
or U1731 (N_1731,In_692,In_599);
and U1732 (N_1732,In_1422,In_822);
or U1733 (N_1733,In_350,In_365);
and U1734 (N_1734,In_66,In_640);
nor U1735 (N_1735,In_145,In_760);
nand U1736 (N_1736,In_354,In_764);
or U1737 (N_1737,In_1447,In_720);
or U1738 (N_1738,In_511,In_368);
nand U1739 (N_1739,In_1325,In_606);
and U1740 (N_1740,In_1190,In_1360);
and U1741 (N_1741,In_1439,In_242);
and U1742 (N_1742,In_715,In_1246);
and U1743 (N_1743,In_79,In_485);
nor U1744 (N_1744,In_772,In_1476);
nand U1745 (N_1745,In_191,In_953);
nand U1746 (N_1746,In_940,In_276);
nor U1747 (N_1747,In_1387,In_1064);
and U1748 (N_1748,In_721,In_313);
or U1749 (N_1749,In_899,In_373);
or U1750 (N_1750,In_1021,In_1012);
or U1751 (N_1751,In_1010,In_1350);
nand U1752 (N_1752,In_388,In_56);
nand U1753 (N_1753,In_980,In_1202);
nand U1754 (N_1754,In_777,In_268);
or U1755 (N_1755,In_612,In_577);
nand U1756 (N_1756,In_425,In_651);
or U1757 (N_1757,In_1072,In_191);
xor U1758 (N_1758,In_1026,In_542);
nand U1759 (N_1759,In_394,In_332);
or U1760 (N_1760,In_63,In_677);
nor U1761 (N_1761,In_626,In_1331);
nor U1762 (N_1762,In_832,In_1438);
nor U1763 (N_1763,In_1320,In_155);
or U1764 (N_1764,In_1214,In_1095);
nand U1765 (N_1765,In_1176,In_102);
and U1766 (N_1766,In_944,In_273);
or U1767 (N_1767,In_70,In_735);
nor U1768 (N_1768,In_1302,In_747);
and U1769 (N_1769,In_1437,In_671);
or U1770 (N_1770,In_1452,In_18);
or U1771 (N_1771,In_1248,In_1297);
and U1772 (N_1772,In_467,In_391);
and U1773 (N_1773,In_458,In_566);
nor U1774 (N_1774,In_1094,In_1458);
or U1775 (N_1775,In_1383,In_140);
and U1776 (N_1776,In_1230,In_688);
or U1777 (N_1777,In_813,In_831);
nor U1778 (N_1778,In_916,In_49);
nand U1779 (N_1779,In_498,In_464);
and U1780 (N_1780,In_545,In_397);
or U1781 (N_1781,In_459,In_1282);
nor U1782 (N_1782,In_309,In_1378);
nand U1783 (N_1783,In_568,In_806);
or U1784 (N_1784,In_1160,In_804);
or U1785 (N_1785,In_540,In_651);
nor U1786 (N_1786,In_395,In_1488);
nand U1787 (N_1787,In_1146,In_67);
and U1788 (N_1788,In_600,In_924);
nand U1789 (N_1789,In_460,In_260);
or U1790 (N_1790,In_709,In_385);
nor U1791 (N_1791,In_42,In_1467);
nand U1792 (N_1792,In_327,In_1419);
nor U1793 (N_1793,In_1309,In_384);
nor U1794 (N_1794,In_197,In_1383);
nor U1795 (N_1795,In_1327,In_1185);
nor U1796 (N_1796,In_433,In_246);
nor U1797 (N_1797,In_1170,In_1407);
nor U1798 (N_1798,In_635,In_391);
nand U1799 (N_1799,In_336,In_65);
nor U1800 (N_1800,In_594,In_1287);
nor U1801 (N_1801,In_1444,In_153);
nand U1802 (N_1802,In_554,In_309);
nor U1803 (N_1803,In_195,In_654);
or U1804 (N_1804,In_8,In_111);
and U1805 (N_1805,In_780,In_706);
nor U1806 (N_1806,In_674,In_82);
nor U1807 (N_1807,In_287,In_238);
or U1808 (N_1808,In_589,In_1244);
and U1809 (N_1809,In_1214,In_1472);
and U1810 (N_1810,In_470,In_1475);
and U1811 (N_1811,In_27,In_738);
and U1812 (N_1812,In_274,In_828);
nor U1813 (N_1813,In_733,In_639);
nor U1814 (N_1814,In_1186,In_493);
nand U1815 (N_1815,In_652,In_1195);
and U1816 (N_1816,In_124,In_1358);
and U1817 (N_1817,In_1401,In_604);
or U1818 (N_1818,In_120,In_940);
nand U1819 (N_1819,In_1229,In_245);
nand U1820 (N_1820,In_94,In_1298);
and U1821 (N_1821,In_266,In_1010);
nor U1822 (N_1822,In_1306,In_236);
or U1823 (N_1823,In_78,In_286);
or U1824 (N_1824,In_678,In_1035);
nand U1825 (N_1825,In_791,In_443);
and U1826 (N_1826,In_1413,In_861);
nor U1827 (N_1827,In_1311,In_295);
and U1828 (N_1828,In_380,In_758);
nor U1829 (N_1829,In_1418,In_814);
or U1830 (N_1830,In_1481,In_420);
or U1831 (N_1831,In_796,In_1490);
or U1832 (N_1832,In_351,In_1187);
nor U1833 (N_1833,In_388,In_426);
nor U1834 (N_1834,In_598,In_1182);
nand U1835 (N_1835,In_166,In_1169);
nor U1836 (N_1836,In_1380,In_788);
or U1837 (N_1837,In_1301,In_1182);
or U1838 (N_1838,In_421,In_29);
nand U1839 (N_1839,In_121,In_184);
nor U1840 (N_1840,In_193,In_1272);
or U1841 (N_1841,In_396,In_779);
nand U1842 (N_1842,In_1278,In_617);
nor U1843 (N_1843,In_1269,In_1308);
or U1844 (N_1844,In_36,In_773);
nand U1845 (N_1845,In_1302,In_1405);
or U1846 (N_1846,In_1013,In_1356);
nand U1847 (N_1847,In_450,In_309);
nand U1848 (N_1848,In_561,In_1269);
and U1849 (N_1849,In_1030,In_1309);
nor U1850 (N_1850,In_110,In_1327);
and U1851 (N_1851,In_120,In_1030);
nor U1852 (N_1852,In_873,In_1160);
nand U1853 (N_1853,In_693,In_139);
nor U1854 (N_1854,In_243,In_1295);
nand U1855 (N_1855,In_1348,In_186);
nand U1856 (N_1856,In_1043,In_84);
nor U1857 (N_1857,In_1137,In_578);
or U1858 (N_1858,In_6,In_1100);
nand U1859 (N_1859,In_580,In_1182);
or U1860 (N_1860,In_766,In_1102);
and U1861 (N_1861,In_1032,In_241);
or U1862 (N_1862,In_111,In_174);
nand U1863 (N_1863,In_1179,In_78);
or U1864 (N_1864,In_921,In_1268);
or U1865 (N_1865,In_1014,In_835);
nand U1866 (N_1866,In_603,In_1218);
or U1867 (N_1867,In_367,In_224);
nand U1868 (N_1868,In_49,In_1149);
nand U1869 (N_1869,In_241,In_28);
nor U1870 (N_1870,In_1409,In_799);
nor U1871 (N_1871,In_1028,In_449);
nand U1872 (N_1872,In_1038,In_599);
and U1873 (N_1873,In_1083,In_91);
nor U1874 (N_1874,In_1244,In_392);
or U1875 (N_1875,In_117,In_466);
nor U1876 (N_1876,In_504,In_1323);
nand U1877 (N_1877,In_427,In_1296);
nor U1878 (N_1878,In_621,In_1283);
nand U1879 (N_1879,In_851,In_1345);
nor U1880 (N_1880,In_1498,In_495);
nand U1881 (N_1881,In_778,In_576);
or U1882 (N_1882,In_330,In_300);
and U1883 (N_1883,In_582,In_1186);
nand U1884 (N_1884,In_472,In_456);
nand U1885 (N_1885,In_352,In_148);
nand U1886 (N_1886,In_1234,In_586);
nand U1887 (N_1887,In_68,In_258);
nand U1888 (N_1888,In_719,In_40);
or U1889 (N_1889,In_131,In_528);
or U1890 (N_1890,In_1481,In_1387);
and U1891 (N_1891,In_1308,In_171);
or U1892 (N_1892,In_73,In_694);
or U1893 (N_1893,In_1487,In_614);
nor U1894 (N_1894,In_839,In_510);
nor U1895 (N_1895,In_473,In_37);
and U1896 (N_1896,In_1006,In_1227);
nand U1897 (N_1897,In_286,In_900);
or U1898 (N_1898,In_521,In_1137);
nand U1899 (N_1899,In_930,In_457);
nor U1900 (N_1900,In_365,In_1320);
nor U1901 (N_1901,In_1448,In_595);
nand U1902 (N_1902,In_400,In_1235);
nand U1903 (N_1903,In_903,In_96);
nor U1904 (N_1904,In_873,In_1030);
nand U1905 (N_1905,In_607,In_1385);
nor U1906 (N_1906,In_361,In_213);
or U1907 (N_1907,In_1016,In_725);
nand U1908 (N_1908,In_79,In_512);
and U1909 (N_1909,In_372,In_577);
nor U1910 (N_1910,In_451,In_1156);
and U1911 (N_1911,In_480,In_102);
or U1912 (N_1912,In_599,In_780);
nand U1913 (N_1913,In_343,In_846);
nand U1914 (N_1914,In_1094,In_1158);
or U1915 (N_1915,In_28,In_1149);
or U1916 (N_1916,In_836,In_551);
or U1917 (N_1917,In_826,In_1422);
nand U1918 (N_1918,In_1242,In_4);
or U1919 (N_1919,In_1455,In_1306);
and U1920 (N_1920,In_1436,In_458);
nand U1921 (N_1921,In_295,In_493);
nand U1922 (N_1922,In_826,In_331);
nor U1923 (N_1923,In_349,In_1022);
nor U1924 (N_1924,In_751,In_744);
nand U1925 (N_1925,In_334,In_1166);
xor U1926 (N_1926,In_23,In_1273);
nand U1927 (N_1927,In_1245,In_233);
and U1928 (N_1928,In_591,In_1382);
nor U1929 (N_1929,In_1254,In_259);
and U1930 (N_1930,In_221,In_183);
nor U1931 (N_1931,In_156,In_1312);
or U1932 (N_1932,In_198,In_513);
or U1933 (N_1933,In_1469,In_873);
nand U1934 (N_1934,In_855,In_160);
and U1935 (N_1935,In_96,In_822);
and U1936 (N_1936,In_384,In_118);
or U1937 (N_1937,In_663,In_226);
nor U1938 (N_1938,In_21,In_267);
and U1939 (N_1939,In_138,In_274);
or U1940 (N_1940,In_1271,In_155);
and U1941 (N_1941,In_400,In_949);
nand U1942 (N_1942,In_54,In_597);
nand U1943 (N_1943,In_828,In_1122);
or U1944 (N_1944,In_645,In_720);
or U1945 (N_1945,In_730,In_562);
and U1946 (N_1946,In_735,In_1191);
nand U1947 (N_1947,In_1494,In_423);
or U1948 (N_1948,In_101,In_253);
or U1949 (N_1949,In_1148,In_832);
or U1950 (N_1950,In_1330,In_368);
nand U1951 (N_1951,In_1491,In_649);
nor U1952 (N_1952,In_1184,In_81);
or U1953 (N_1953,In_1486,In_438);
nor U1954 (N_1954,In_1317,In_223);
nand U1955 (N_1955,In_766,In_1052);
or U1956 (N_1956,In_1036,In_1064);
xor U1957 (N_1957,In_1343,In_1170);
nor U1958 (N_1958,In_1212,In_487);
xor U1959 (N_1959,In_1381,In_118);
nand U1960 (N_1960,In_1135,In_952);
or U1961 (N_1961,In_1043,In_247);
and U1962 (N_1962,In_1347,In_820);
nand U1963 (N_1963,In_1422,In_169);
and U1964 (N_1964,In_432,In_814);
or U1965 (N_1965,In_608,In_688);
or U1966 (N_1966,In_1197,In_349);
and U1967 (N_1967,In_1101,In_1483);
or U1968 (N_1968,In_795,In_1101);
nor U1969 (N_1969,In_102,In_956);
nor U1970 (N_1970,In_301,In_1265);
nor U1971 (N_1971,In_477,In_227);
or U1972 (N_1972,In_546,In_160);
nor U1973 (N_1973,In_903,In_1196);
nor U1974 (N_1974,In_1408,In_602);
or U1975 (N_1975,In_870,In_439);
or U1976 (N_1976,In_208,In_5);
nand U1977 (N_1977,In_408,In_662);
or U1978 (N_1978,In_1418,In_1128);
or U1979 (N_1979,In_103,In_524);
nand U1980 (N_1980,In_461,In_1233);
nor U1981 (N_1981,In_1007,In_78);
and U1982 (N_1982,In_1173,In_714);
or U1983 (N_1983,In_234,In_239);
xnor U1984 (N_1984,In_206,In_1095);
and U1985 (N_1985,In_310,In_721);
and U1986 (N_1986,In_1379,In_809);
or U1987 (N_1987,In_71,In_257);
nand U1988 (N_1988,In_600,In_801);
nor U1989 (N_1989,In_913,In_16);
nand U1990 (N_1990,In_1321,In_453);
nand U1991 (N_1991,In_604,In_1251);
and U1992 (N_1992,In_817,In_1006);
nor U1993 (N_1993,In_955,In_1203);
nand U1994 (N_1994,In_578,In_745);
nor U1995 (N_1995,In_742,In_33);
or U1996 (N_1996,In_1212,In_552);
and U1997 (N_1997,In_617,In_1047);
and U1998 (N_1998,In_1303,In_1329);
and U1999 (N_1999,In_439,In_741);
nor U2000 (N_2000,In_1246,In_1198);
nor U2001 (N_2001,In_808,In_717);
nor U2002 (N_2002,In_583,In_147);
nand U2003 (N_2003,In_970,In_9);
nor U2004 (N_2004,In_901,In_404);
and U2005 (N_2005,In_986,In_58);
or U2006 (N_2006,In_70,In_520);
or U2007 (N_2007,In_1170,In_706);
nor U2008 (N_2008,In_569,In_747);
nand U2009 (N_2009,In_490,In_1338);
nor U2010 (N_2010,In_266,In_172);
and U2011 (N_2011,In_1027,In_349);
nor U2012 (N_2012,In_1305,In_708);
and U2013 (N_2013,In_440,In_1096);
or U2014 (N_2014,In_625,In_1004);
nand U2015 (N_2015,In_220,In_77);
nand U2016 (N_2016,In_632,In_1271);
and U2017 (N_2017,In_24,In_1223);
nand U2018 (N_2018,In_1277,In_1144);
nand U2019 (N_2019,In_144,In_95);
nor U2020 (N_2020,In_1071,In_187);
and U2021 (N_2021,In_1320,In_654);
or U2022 (N_2022,In_787,In_1139);
nand U2023 (N_2023,In_324,In_319);
nor U2024 (N_2024,In_1481,In_1367);
or U2025 (N_2025,In_96,In_88);
xor U2026 (N_2026,In_1246,In_736);
or U2027 (N_2027,In_1163,In_600);
nor U2028 (N_2028,In_812,In_795);
nand U2029 (N_2029,In_675,In_128);
nor U2030 (N_2030,In_1264,In_508);
nor U2031 (N_2031,In_1073,In_223);
nor U2032 (N_2032,In_220,In_239);
nor U2033 (N_2033,In_1419,In_624);
or U2034 (N_2034,In_145,In_1474);
nor U2035 (N_2035,In_828,In_169);
nor U2036 (N_2036,In_212,In_549);
and U2037 (N_2037,In_1080,In_1116);
or U2038 (N_2038,In_904,In_705);
nor U2039 (N_2039,In_226,In_259);
nand U2040 (N_2040,In_1136,In_461);
or U2041 (N_2041,In_535,In_344);
and U2042 (N_2042,In_173,In_387);
nor U2043 (N_2043,In_403,In_277);
nor U2044 (N_2044,In_1369,In_604);
or U2045 (N_2045,In_1354,In_424);
nand U2046 (N_2046,In_784,In_829);
nor U2047 (N_2047,In_990,In_2);
nand U2048 (N_2048,In_967,In_1138);
or U2049 (N_2049,In_1101,In_971);
xnor U2050 (N_2050,In_874,In_1413);
nand U2051 (N_2051,In_1356,In_18);
and U2052 (N_2052,In_835,In_350);
and U2053 (N_2053,In_634,In_1296);
or U2054 (N_2054,In_1239,In_876);
nand U2055 (N_2055,In_1061,In_767);
nand U2056 (N_2056,In_835,In_607);
or U2057 (N_2057,In_645,In_685);
or U2058 (N_2058,In_342,In_482);
nor U2059 (N_2059,In_165,In_434);
nand U2060 (N_2060,In_1416,In_422);
or U2061 (N_2061,In_821,In_386);
or U2062 (N_2062,In_1230,In_1132);
nand U2063 (N_2063,In_101,In_345);
nor U2064 (N_2064,In_380,In_285);
xnor U2065 (N_2065,In_1108,In_84);
nor U2066 (N_2066,In_367,In_441);
nor U2067 (N_2067,In_1415,In_367);
or U2068 (N_2068,In_965,In_508);
or U2069 (N_2069,In_1431,In_1288);
or U2070 (N_2070,In_1067,In_867);
or U2071 (N_2071,In_266,In_1165);
or U2072 (N_2072,In_499,In_1389);
nor U2073 (N_2073,In_1432,In_210);
or U2074 (N_2074,In_195,In_1126);
nand U2075 (N_2075,In_436,In_79);
and U2076 (N_2076,In_788,In_1265);
and U2077 (N_2077,In_595,In_965);
or U2078 (N_2078,In_1121,In_15);
and U2079 (N_2079,In_908,In_318);
nand U2080 (N_2080,In_1363,In_946);
or U2081 (N_2081,In_55,In_1038);
and U2082 (N_2082,In_480,In_1367);
nand U2083 (N_2083,In_427,In_1208);
or U2084 (N_2084,In_1392,In_1239);
and U2085 (N_2085,In_740,In_1237);
or U2086 (N_2086,In_1364,In_651);
or U2087 (N_2087,In_517,In_2);
nor U2088 (N_2088,In_496,In_1418);
and U2089 (N_2089,In_1119,In_1170);
nor U2090 (N_2090,In_699,In_993);
nor U2091 (N_2091,In_1359,In_233);
nand U2092 (N_2092,In_806,In_823);
or U2093 (N_2093,In_631,In_824);
nand U2094 (N_2094,In_130,In_603);
nand U2095 (N_2095,In_178,In_629);
or U2096 (N_2096,In_52,In_209);
or U2097 (N_2097,In_1074,In_948);
nand U2098 (N_2098,In_292,In_1184);
and U2099 (N_2099,In_849,In_388);
nor U2100 (N_2100,In_1111,In_881);
or U2101 (N_2101,In_118,In_104);
nor U2102 (N_2102,In_648,In_1438);
nor U2103 (N_2103,In_609,In_799);
nand U2104 (N_2104,In_510,In_1384);
nor U2105 (N_2105,In_1145,In_1361);
nand U2106 (N_2106,In_892,In_291);
or U2107 (N_2107,In_390,In_742);
xor U2108 (N_2108,In_714,In_519);
or U2109 (N_2109,In_1409,In_180);
nor U2110 (N_2110,In_1267,In_1104);
or U2111 (N_2111,In_1272,In_854);
xnor U2112 (N_2112,In_3,In_944);
nor U2113 (N_2113,In_192,In_739);
nor U2114 (N_2114,In_74,In_794);
or U2115 (N_2115,In_225,In_1203);
or U2116 (N_2116,In_218,In_840);
nand U2117 (N_2117,In_1278,In_226);
nand U2118 (N_2118,In_336,In_1199);
and U2119 (N_2119,In_1228,In_1396);
nor U2120 (N_2120,In_1397,In_242);
and U2121 (N_2121,In_712,In_898);
nand U2122 (N_2122,In_1066,In_1230);
or U2123 (N_2123,In_602,In_235);
nor U2124 (N_2124,In_953,In_630);
nand U2125 (N_2125,In_1018,In_1121);
xnor U2126 (N_2126,In_531,In_1329);
nand U2127 (N_2127,In_792,In_326);
and U2128 (N_2128,In_670,In_1235);
nand U2129 (N_2129,In_312,In_698);
nor U2130 (N_2130,In_6,In_1077);
nor U2131 (N_2131,In_910,In_265);
nor U2132 (N_2132,In_1499,In_158);
and U2133 (N_2133,In_41,In_1280);
nand U2134 (N_2134,In_387,In_65);
nand U2135 (N_2135,In_628,In_70);
or U2136 (N_2136,In_687,In_215);
nand U2137 (N_2137,In_339,In_521);
and U2138 (N_2138,In_771,In_1166);
and U2139 (N_2139,In_450,In_811);
nand U2140 (N_2140,In_502,In_860);
xor U2141 (N_2141,In_815,In_1231);
and U2142 (N_2142,In_185,In_947);
and U2143 (N_2143,In_1394,In_649);
nor U2144 (N_2144,In_811,In_1098);
nor U2145 (N_2145,In_1121,In_577);
nand U2146 (N_2146,In_1405,In_163);
and U2147 (N_2147,In_589,In_809);
nand U2148 (N_2148,In_391,In_507);
and U2149 (N_2149,In_1271,In_407);
and U2150 (N_2150,In_980,In_57);
and U2151 (N_2151,In_1186,In_1208);
nand U2152 (N_2152,In_202,In_959);
nand U2153 (N_2153,In_561,In_1148);
nor U2154 (N_2154,In_826,In_1266);
nand U2155 (N_2155,In_1479,In_1034);
nand U2156 (N_2156,In_796,In_496);
or U2157 (N_2157,In_463,In_805);
or U2158 (N_2158,In_667,In_330);
or U2159 (N_2159,In_1458,In_1018);
nand U2160 (N_2160,In_1291,In_234);
and U2161 (N_2161,In_946,In_402);
or U2162 (N_2162,In_1352,In_50);
nand U2163 (N_2163,In_1332,In_1156);
nand U2164 (N_2164,In_684,In_1422);
nor U2165 (N_2165,In_562,In_524);
nand U2166 (N_2166,In_1276,In_312);
nor U2167 (N_2167,In_605,In_1061);
nor U2168 (N_2168,In_652,In_1175);
xnor U2169 (N_2169,In_1277,In_43);
nand U2170 (N_2170,In_403,In_731);
or U2171 (N_2171,In_1470,In_1276);
nor U2172 (N_2172,In_127,In_385);
nor U2173 (N_2173,In_1000,In_863);
and U2174 (N_2174,In_393,In_844);
nand U2175 (N_2175,In_1392,In_1286);
nor U2176 (N_2176,In_1369,In_337);
nor U2177 (N_2177,In_1090,In_92);
nand U2178 (N_2178,In_1060,In_416);
nand U2179 (N_2179,In_838,In_519);
and U2180 (N_2180,In_988,In_857);
nand U2181 (N_2181,In_1123,In_850);
nand U2182 (N_2182,In_251,In_861);
nand U2183 (N_2183,In_164,In_8);
or U2184 (N_2184,In_1100,In_313);
nand U2185 (N_2185,In_722,In_924);
nand U2186 (N_2186,In_279,In_931);
nand U2187 (N_2187,In_930,In_171);
and U2188 (N_2188,In_306,In_567);
nor U2189 (N_2189,In_723,In_420);
nand U2190 (N_2190,In_261,In_351);
and U2191 (N_2191,In_198,In_811);
nand U2192 (N_2192,In_620,In_1351);
or U2193 (N_2193,In_1161,In_785);
and U2194 (N_2194,In_862,In_850);
or U2195 (N_2195,In_470,In_1098);
or U2196 (N_2196,In_1289,In_331);
nor U2197 (N_2197,In_988,In_366);
nand U2198 (N_2198,In_944,In_1323);
and U2199 (N_2199,In_1152,In_1258);
and U2200 (N_2200,In_770,In_1056);
and U2201 (N_2201,In_1348,In_841);
nand U2202 (N_2202,In_606,In_33);
nand U2203 (N_2203,In_122,In_866);
or U2204 (N_2204,In_969,In_640);
or U2205 (N_2205,In_1421,In_984);
and U2206 (N_2206,In_1126,In_1023);
nand U2207 (N_2207,In_341,In_613);
or U2208 (N_2208,In_867,In_1478);
nand U2209 (N_2209,In_1319,In_850);
and U2210 (N_2210,In_889,In_363);
and U2211 (N_2211,In_139,In_154);
and U2212 (N_2212,In_970,In_912);
nor U2213 (N_2213,In_1185,In_1139);
nand U2214 (N_2214,In_821,In_1119);
nor U2215 (N_2215,In_473,In_1469);
nand U2216 (N_2216,In_542,In_1060);
or U2217 (N_2217,In_1302,In_386);
and U2218 (N_2218,In_1150,In_1226);
and U2219 (N_2219,In_1084,In_193);
or U2220 (N_2220,In_354,In_989);
nor U2221 (N_2221,In_977,In_245);
and U2222 (N_2222,In_747,In_449);
or U2223 (N_2223,In_538,In_778);
and U2224 (N_2224,In_565,In_1085);
and U2225 (N_2225,In_1350,In_612);
or U2226 (N_2226,In_164,In_909);
or U2227 (N_2227,In_336,In_502);
nand U2228 (N_2228,In_849,In_92);
nor U2229 (N_2229,In_1474,In_679);
or U2230 (N_2230,In_63,In_471);
or U2231 (N_2231,In_698,In_248);
or U2232 (N_2232,In_1342,In_1045);
nand U2233 (N_2233,In_988,In_1375);
or U2234 (N_2234,In_802,In_406);
or U2235 (N_2235,In_1445,In_925);
nand U2236 (N_2236,In_881,In_456);
and U2237 (N_2237,In_640,In_394);
or U2238 (N_2238,In_746,In_1075);
or U2239 (N_2239,In_501,In_162);
nor U2240 (N_2240,In_508,In_669);
nand U2241 (N_2241,In_865,In_971);
or U2242 (N_2242,In_610,In_354);
nor U2243 (N_2243,In_522,In_1058);
and U2244 (N_2244,In_56,In_1024);
nand U2245 (N_2245,In_1130,In_697);
nand U2246 (N_2246,In_1239,In_1300);
or U2247 (N_2247,In_1198,In_394);
nand U2248 (N_2248,In_1220,In_1440);
or U2249 (N_2249,In_683,In_388);
nor U2250 (N_2250,In_1496,In_82);
and U2251 (N_2251,In_1221,In_698);
nand U2252 (N_2252,In_1476,In_1058);
and U2253 (N_2253,In_408,In_633);
or U2254 (N_2254,In_245,In_1217);
nand U2255 (N_2255,In_1075,In_305);
and U2256 (N_2256,In_130,In_1492);
nand U2257 (N_2257,In_528,In_1021);
or U2258 (N_2258,In_316,In_278);
nand U2259 (N_2259,In_1432,In_623);
nand U2260 (N_2260,In_840,In_1299);
and U2261 (N_2261,In_977,In_15);
and U2262 (N_2262,In_324,In_372);
and U2263 (N_2263,In_1119,In_1086);
nor U2264 (N_2264,In_278,In_348);
nand U2265 (N_2265,In_1394,In_370);
or U2266 (N_2266,In_61,In_1365);
nor U2267 (N_2267,In_1164,In_247);
nor U2268 (N_2268,In_596,In_832);
or U2269 (N_2269,In_953,In_1122);
or U2270 (N_2270,In_982,In_501);
and U2271 (N_2271,In_176,In_575);
nor U2272 (N_2272,In_1020,In_79);
xor U2273 (N_2273,In_523,In_1413);
nor U2274 (N_2274,In_983,In_283);
and U2275 (N_2275,In_309,In_726);
nand U2276 (N_2276,In_469,In_1464);
or U2277 (N_2277,In_1057,In_218);
and U2278 (N_2278,In_156,In_346);
and U2279 (N_2279,In_1452,In_145);
and U2280 (N_2280,In_1345,In_446);
or U2281 (N_2281,In_980,In_1047);
or U2282 (N_2282,In_1218,In_910);
or U2283 (N_2283,In_65,In_661);
and U2284 (N_2284,In_985,In_1429);
and U2285 (N_2285,In_292,In_726);
and U2286 (N_2286,In_598,In_443);
nand U2287 (N_2287,In_1313,In_703);
nor U2288 (N_2288,In_186,In_1400);
and U2289 (N_2289,In_668,In_55);
and U2290 (N_2290,In_1075,In_367);
nand U2291 (N_2291,In_883,In_1178);
nor U2292 (N_2292,In_525,In_432);
nand U2293 (N_2293,In_1219,In_809);
or U2294 (N_2294,In_164,In_1324);
or U2295 (N_2295,In_857,In_1366);
nand U2296 (N_2296,In_688,In_1471);
or U2297 (N_2297,In_312,In_1015);
nor U2298 (N_2298,In_1091,In_779);
or U2299 (N_2299,In_592,In_1245);
and U2300 (N_2300,In_858,In_632);
nand U2301 (N_2301,In_232,In_1081);
nor U2302 (N_2302,In_1282,In_607);
nand U2303 (N_2303,In_1166,In_678);
and U2304 (N_2304,In_473,In_1120);
or U2305 (N_2305,In_124,In_454);
nor U2306 (N_2306,In_1237,In_729);
and U2307 (N_2307,In_464,In_1315);
nand U2308 (N_2308,In_197,In_81);
nand U2309 (N_2309,In_184,In_1157);
or U2310 (N_2310,In_563,In_1322);
or U2311 (N_2311,In_1212,In_1358);
or U2312 (N_2312,In_539,In_251);
nand U2313 (N_2313,In_443,In_669);
or U2314 (N_2314,In_1264,In_1294);
nor U2315 (N_2315,In_11,In_1358);
nor U2316 (N_2316,In_1398,In_1152);
nor U2317 (N_2317,In_1329,In_1195);
and U2318 (N_2318,In_1202,In_487);
and U2319 (N_2319,In_50,In_820);
and U2320 (N_2320,In_864,In_550);
and U2321 (N_2321,In_11,In_1110);
and U2322 (N_2322,In_1430,In_494);
nor U2323 (N_2323,In_1174,In_63);
nor U2324 (N_2324,In_1333,In_52);
and U2325 (N_2325,In_836,In_1428);
nand U2326 (N_2326,In_136,In_1175);
and U2327 (N_2327,In_815,In_354);
nand U2328 (N_2328,In_637,In_567);
nor U2329 (N_2329,In_407,In_136);
or U2330 (N_2330,In_227,In_528);
nand U2331 (N_2331,In_1079,In_1468);
and U2332 (N_2332,In_7,In_1158);
or U2333 (N_2333,In_1082,In_1160);
nor U2334 (N_2334,In_632,In_275);
nand U2335 (N_2335,In_1180,In_135);
and U2336 (N_2336,In_1109,In_568);
nor U2337 (N_2337,In_618,In_430);
nand U2338 (N_2338,In_610,In_1083);
nor U2339 (N_2339,In_905,In_1040);
nor U2340 (N_2340,In_1003,In_72);
nand U2341 (N_2341,In_1279,In_1282);
nand U2342 (N_2342,In_1418,In_582);
nor U2343 (N_2343,In_489,In_913);
nand U2344 (N_2344,In_1450,In_1365);
nand U2345 (N_2345,In_647,In_485);
and U2346 (N_2346,In_1371,In_149);
or U2347 (N_2347,In_1117,In_793);
and U2348 (N_2348,In_1244,In_554);
nand U2349 (N_2349,In_2,In_1304);
and U2350 (N_2350,In_1458,In_1025);
or U2351 (N_2351,In_391,In_980);
or U2352 (N_2352,In_224,In_1430);
and U2353 (N_2353,In_1089,In_45);
and U2354 (N_2354,In_1339,In_1483);
nor U2355 (N_2355,In_1123,In_330);
nor U2356 (N_2356,In_298,In_1319);
nand U2357 (N_2357,In_1005,In_480);
and U2358 (N_2358,In_1011,In_522);
nand U2359 (N_2359,In_405,In_896);
and U2360 (N_2360,In_704,In_286);
nor U2361 (N_2361,In_973,In_610);
and U2362 (N_2362,In_1337,In_385);
or U2363 (N_2363,In_1073,In_648);
nand U2364 (N_2364,In_1285,In_200);
nand U2365 (N_2365,In_694,In_331);
xor U2366 (N_2366,In_1150,In_1249);
nor U2367 (N_2367,In_1183,In_298);
and U2368 (N_2368,In_1421,In_631);
nand U2369 (N_2369,In_1138,In_1248);
and U2370 (N_2370,In_792,In_178);
and U2371 (N_2371,In_562,In_544);
nor U2372 (N_2372,In_174,In_1416);
and U2373 (N_2373,In_352,In_614);
nor U2374 (N_2374,In_1004,In_581);
and U2375 (N_2375,In_454,In_1082);
nand U2376 (N_2376,In_357,In_242);
nand U2377 (N_2377,In_1223,In_1183);
nor U2378 (N_2378,In_991,In_420);
nor U2379 (N_2379,In_1384,In_612);
nand U2380 (N_2380,In_8,In_709);
or U2381 (N_2381,In_457,In_569);
or U2382 (N_2382,In_1042,In_1194);
nor U2383 (N_2383,In_754,In_561);
nand U2384 (N_2384,In_1150,In_1074);
nor U2385 (N_2385,In_571,In_97);
or U2386 (N_2386,In_245,In_722);
or U2387 (N_2387,In_1395,In_819);
nor U2388 (N_2388,In_78,In_1103);
or U2389 (N_2389,In_177,In_159);
and U2390 (N_2390,In_667,In_1474);
nor U2391 (N_2391,In_1450,In_979);
nor U2392 (N_2392,In_1220,In_31);
nor U2393 (N_2393,In_1082,In_1011);
nor U2394 (N_2394,In_966,In_1170);
nor U2395 (N_2395,In_114,In_91);
or U2396 (N_2396,In_486,In_1361);
nor U2397 (N_2397,In_1133,In_1404);
nor U2398 (N_2398,In_851,In_475);
nor U2399 (N_2399,In_548,In_329);
and U2400 (N_2400,In_267,In_1166);
nor U2401 (N_2401,In_1144,In_694);
nor U2402 (N_2402,In_900,In_440);
nand U2403 (N_2403,In_1109,In_1496);
and U2404 (N_2404,In_863,In_943);
or U2405 (N_2405,In_1415,In_543);
and U2406 (N_2406,In_1452,In_1370);
nand U2407 (N_2407,In_25,In_377);
or U2408 (N_2408,In_909,In_510);
and U2409 (N_2409,In_782,In_779);
and U2410 (N_2410,In_107,In_987);
or U2411 (N_2411,In_1085,In_117);
and U2412 (N_2412,In_1292,In_1207);
and U2413 (N_2413,In_655,In_745);
and U2414 (N_2414,In_1404,In_267);
nor U2415 (N_2415,In_463,In_1015);
nand U2416 (N_2416,In_264,In_61);
and U2417 (N_2417,In_679,In_627);
nor U2418 (N_2418,In_1173,In_477);
nand U2419 (N_2419,In_232,In_515);
and U2420 (N_2420,In_711,In_337);
or U2421 (N_2421,In_464,In_280);
nand U2422 (N_2422,In_441,In_849);
or U2423 (N_2423,In_522,In_1387);
nand U2424 (N_2424,In_949,In_371);
or U2425 (N_2425,In_1148,In_706);
or U2426 (N_2426,In_796,In_1135);
nand U2427 (N_2427,In_108,In_79);
nand U2428 (N_2428,In_89,In_753);
and U2429 (N_2429,In_492,In_1147);
or U2430 (N_2430,In_1131,In_1277);
nor U2431 (N_2431,In_1269,In_699);
or U2432 (N_2432,In_1416,In_424);
xor U2433 (N_2433,In_1405,In_1279);
or U2434 (N_2434,In_946,In_465);
nor U2435 (N_2435,In_424,In_129);
nor U2436 (N_2436,In_635,In_45);
nand U2437 (N_2437,In_534,In_855);
and U2438 (N_2438,In_20,In_1424);
or U2439 (N_2439,In_895,In_989);
or U2440 (N_2440,In_793,In_62);
and U2441 (N_2441,In_1445,In_315);
and U2442 (N_2442,In_872,In_694);
nand U2443 (N_2443,In_778,In_285);
nor U2444 (N_2444,In_1245,In_1301);
nand U2445 (N_2445,In_620,In_1404);
nor U2446 (N_2446,In_14,In_630);
nor U2447 (N_2447,In_477,In_635);
and U2448 (N_2448,In_119,In_1200);
and U2449 (N_2449,In_237,In_702);
and U2450 (N_2450,In_1392,In_419);
and U2451 (N_2451,In_1292,In_698);
nor U2452 (N_2452,In_818,In_896);
and U2453 (N_2453,In_438,In_1353);
or U2454 (N_2454,In_584,In_504);
nor U2455 (N_2455,In_1470,In_523);
and U2456 (N_2456,In_115,In_299);
nand U2457 (N_2457,In_969,In_1226);
or U2458 (N_2458,In_805,In_217);
nor U2459 (N_2459,In_674,In_49);
or U2460 (N_2460,In_158,In_1141);
nand U2461 (N_2461,In_1044,In_1104);
and U2462 (N_2462,In_62,In_833);
or U2463 (N_2463,In_884,In_1288);
or U2464 (N_2464,In_1371,In_260);
and U2465 (N_2465,In_206,In_633);
nor U2466 (N_2466,In_432,In_827);
nor U2467 (N_2467,In_802,In_1116);
or U2468 (N_2468,In_1112,In_1342);
nand U2469 (N_2469,In_61,In_410);
nor U2470 (N_2470,In_405,In_835);
or U2471 (N_2471,In_1491,In_1370);
nor U2472 (N_2472,In_880,In_386);
and U2473 (N_2473,In_805,In_1306);
or U2474 (N_2474,In_199,In_326);
and U2475 (N_2475,In_1479,In_753);
or U2476 (N_2476,In_1318,In_1175);
nand U2477 (N_2477,In_1000,In_1165);
nand U2478 (N_2478,In_610,In_819);
or U2479 (N_2479,In_298,In_39);
nand U2480 (N_2480,In_0,In_777);
or U2481 (N_2481,In_4,In_1236);
nand U2482 (N_2482,In_892,In_98);
nor U2483 (N_2483,In_1200,In_1413);
nor U2484 (N_2484,In_433,In_798);
and U2485 (N_2485,In_796,In_138);
and U2486 (N_2486,In_1292,In_568);
and U2487 (N_2487,In_1314,In_570);
nor U2488 (N_2488,In_881,In_1032);
nor U2489 (N_2489,In_31,In_332);
or U2490 (N_2490,In_427,In_680);
nand U2491 (N_2491,In_581,In_930);
or U2492 (N_2492,In_328,In_86);
nor U2493 (N_2493,In_437,In_7);
nand U2494 (N_2494,In_910,In_457);
or U2495 (N_2495,In_26,In_470);
nor U2496 (N_2496,In_587,In_95);
or U2497 (N_2497,In_1109,In_272);
nor U2498 (N_2498,In_98,In_1274);
nand U2499 (N_2499,In_447,In_1374);
nand U2500 (N_2500,In_49,In_1044);
or U2501 (N_2501,In_308,In_604);
or U2502 (N_2502,In_1031,In_895);
or U2503 (N_2503,In_473,In_587);
or U2504 (N_2504,In_892,In_20);
or U2505 (N_2505,In_685,In_420);
and U2506 (N_2506,In_178,In_1317);
nor U2507 (N_2507,In_1261,In_1249);
nand U2508 (N_2508,In_359,In_955);
or U2509 (N_2509,In_2,In_1305);
nor U2510 (N_2510,In_563,In_303);
or U2511 (N_2511,In_1112,In_945);
nand U2512 (N_2512,In_147,In_517);
nor U2513 (N_2513,In_806,In_137);
and U2514 (N_2514,In_980,In_1396);
nand U2515 (N_2515,In_235,In_1083);
nand U2516 (N_2516,In_1392,In_159);
nor U2517 (N_2517,In_532,In_337);
or U2518 (N_2518,In_474,In_1281);
nor U2519 (N_2519,In_226,In_787);
and U2520 (N_2520,In_463,In_11);
nor U2521 (N_2521,In_1071,In_547);
or U2522 (N_2522,In_574,In_809);
nor U2523 (N_2523,In_507,In_807);
or U2524 (N_2524,In_1452,In_1412);
and U2525 (N_2525,In_701,In_110);
and U2526 (N_2526,In_315,In_572);
or U2527 (N_2527,In_126,In_118);
or U2528 (N_2528,In_1237,In_1165);
nor U2529 (N_2529,In_952,In_1183);
or U2530 (N_2530,In_1369,In_410);
nor U2531 (N_2531,In_475,In_1157);
or U2532 (N_2532,In_1395,In_854);
and U2533 (N_2533,In_1160,In_1407);
nand U2534 (N_2534,In_457,In_1183);
and U2535 (N_2535,In_1423,In_998);
and U2536 (N_2536,In_65,In_538);
nor U2537 (N_2537,In_730,In_1377);
nor U2538 (N_2538,In_216,In_759);
nand U2539 (N_2539,In_165,In_381);
nor U2540 (N_2540,In_622,In_819);
and U2541 (N_2541,In_174,In_1382);
or U2542 (N_2542,In_576,In_722);
nand U2543 (N_2543,In_523,In_604);
and U2544 (N_2544,In_1057,In_796);
nand U2545 (N_2545,In_533,In_836);
nand U2546 (N_2546,In_1224,In_905);
nor U2547 (N_2547,In_26,In_956);
or U2548 (N_2548,In_647,In_1140);
nand U2549 (N_2549,In_1328,In_966);
and U2550 (N_2550,In_650,In_1019);
and U2551 (N_2551,In_1214,In_754);
nor U2552 (N_2552,In_325,In_703);
nand U2553 (N_2553,In_714,In_44);
nor U2554 (N_2554,In_1137,In_168);
or U2555 (N_2555,In_936,In_1378);
nor U2556 (N_2556,In_991,In_340);
nor U2557 (N_2557,In_664,In_172);
nand U2558 (N_2558,In_1036,In_1113);
nor U2559 (N_2559,In_785,In_1136);
nand U2560 (N_2560,In_660,In_1241);
xnor U2561 (N_2561,In_434,In_215);
nor U2562 (N_2562,In_411,In_1221);
nor U2563 (N_2563,In_166,In_1336);
nor U2564 (N_2564,In_1061,In_914);
and U2565 (N_2565,In_22,In_672);
nand U2566 (N_2566,In_691,In_195);
nand U2567 (N_2567,In_887,In_1301);
and U2568 (N_2568,In_990,In_1001);
nand U2569 (N_2569,In_1445,In_537);
and U2570 (N_2570,In_188,In_1305);
or U2571 (N_2571,In_353,In_671);
and U2572 (N_2572,In_810,In_150);
and U2573 (N_2573,In_386,In_1465);
nor U2574 (N_2574,In_762,In_138);
and U2575 (N_2575,In_1390,In_977);
nor U2576 (N_2576,In_765,In_4);
nor U2577 (N_2577,In_387,In_1265);
or U2578 (N_2578,In_1275,In_248);
nand U2579 (N_2579,In_560,In_504);
nor U2580 (N_2580,In_282,In_841);
nand U2581 (N_2581,In_106,In_475);
or U2582 (N_2582,In_1241,In_1348);
nand U2583 (N_2583,In_975,In_58);
or U2584 (N_2584,In_782,In_714);
nor U2585 (N_2585,In_457,In_485);
and U2586 (N_2586,In_280,In_59);
nor U2587 (N_2587,In_735,In_1108);
nand U2588 (N_2588,In_637,In_825);
nand U2589 (N_2589,In_546,In_488);
nand U2590 (N_2590,In_1286,In_934);
and U2591 (N_2591,In_1225,In_1222);
nor U2592 (N_2592,In_644,In_79);
nand U2593 (N_2593,In_1196,In_1188);
nor U2594 (N_2594,In_498,In_846);
nor U2595 (N_2595,In_1159,In_1339);
or U2596 (N_2596,In_179,In_856);
nand U2597 (N_2597,In_1256,In_590);
nor U2598 (N_2598,In_1443,In_1010);
and U2599 (N_2599,In_1237,In_690);
and U2600 (N_2600,In_1321,In_1415);
and U2601 (N_2601,In_805,In_166);
or U2602 (N_2602,In_1155,In_587);
nor U2603 (N_2603,In_523,In_35);
or U2604 (N_2604,In_857,In_552);
or U2605 (N_2605,In_1067,In_1003);
nand U2606 (N_2606,In_905,In_857);
nor U2607 (N_2607,In_388,In_1459);
and U2608 (N_2608,In_1476,In_1398);
or U2609 (N_2609,In_1290,In_404);
nand U2610 (N_2610,In_729,In_700);
or U2611 (N_2611,In_997,In_1101);
nor U2612 (N_2612,In_245,In_949);
or U2613 (N_2613,In_898,In_766);
nor U2614 (N_2614,In_1233,In_88);
or U2615 (N_2615,In_690,In_757);
nor U2616 (N_2616,In_416,In_1054);
nor U2617 (N_2617,In_1044,In_34);
or U2618 (N_2618,In_514,In_178);
and U2619 (N_2619,In_117,In_549);
or U2620 (N_2620,In_336,In_57);
nor U2621 (N_2621,In_34,In_1020);
and U2622 (N_2622,In_1385,In_575);
nor U2623 (N_2623,In_360,In_90);
nand U2624 (N_2624,In_571,In_839);
nand U2625 (N_2625,In_393,In_420);
or U2626 (N_2626,In_554,In_484);
and U2627 (N_2627,In_1387,In_366);
nand U2628 (N_2628,In_1042,In_354);
and U2629 (N_2629,In_472,In_1313);
nor U2630 (N_2630,In_795,In_1346);
and U2631 (N_2631,In_136,In_441);
nand U2632 (N_2632,In_1131,In_952);
or U2633 (N_2633,In_361,In_206);
and U2634 (N_2634,In_514,In_82);
and U2635 (N_2635,In_1127,In_1468);
nand U2636 (N_2636,In_841,In_378);
or U2637 (N_2637,In_629,In_69);
nor U2638 (N_2638,In_1086,In_260);
or U2639 (N_2639,In_1442,In_272);
nand U2640 (N_2640,In_688,In_1143);
or U2641 (N_2641,In_930,In_745);
nor U2642 (N_2642,In_994,In_160);
or U2643 (N_2643,In_224,In_61);
nor U2644 (N_2644,In_406,In_725);
nor U2645 (N_2645,In_1088,In_522);
xor U2646 (N_2646,In_585,In_1031);
nand U2647 (N_2647,In_101,In_735);
nor U2648 (N_2648,In_431,In_837);
and U2649 (N_2649,In_234,In_157);
xor U2650 (N_2650,In_809,In_1478);
nand U2651 (N_2651,In_519,In_238);
nor U2652 (N_2652,In_877,In_428);
nor U2653 (N_2653,In_793,In_993);
nand U2654 (N_2654,In_418,In_351);
nand U2655 (N_2655,In_193,In_1269);
and U2656 (N_2656,In_1245,In_966);
and U2657 (N_2657,In_61,In_536);
and U2658 (N_2658,In_926,In_1251);
and U2659 (N_2659,In_456,In_164);
nand U2660 (N_2660,In_1395,In_226);
or U2661 (N_2661,In_813,In_507);
or U2662 (N_2662,In_180,In_1074);
or U2663 (N_2663,In_1463,In_441);
and U2664 (N_2664,In_151,In_212);
nand U2665 (N_2665,In_239,In_410);
nand U2666 (N_2666,In_446,In_1458);
nand U2667 (N_2667,In_148,In_1457);
and U2668 (N_2668,In_1375,In_240);
nand U2669 (N_2669,In_1284,In_1267);
and U2670 (N_2670,In_1470,In_512);
nand U2671 (N_2671,In_713,In_944);
nand U2672 (N_2672,In_697,In_1033);
nand U2673 (N_2673,In_920,In_408);
nand U2674 (N_2674,In_736,In_1141);
and U2675 (N_2675,In_1025,In_898);
and U2676 (N_2676,In_1258,In_1256);
nor U2677 (N_2677,In_516,In_1490);
nand U2678 (N_2678,In_1148,In_80);
nor U2679 (N_2679,In_251,In_889);
nor U2680 (N_2680,In_1056,In_1017);
nor U2681 (N_2681,In_467,In_1276);
or U2682 (N_2682,In_1469,In_233);
or U2683 (N_2683,In_1326,In_752);
nor U2684 (N_2684,In_1226,In_1063);
and U2685 (N_2685,In_675,In_196);
nand U2686 (N_2686,In_187,In_549);
nand U2687 (N_2687,In_626,In_1118);
and U2688 (N_2688,In_24,In_466);
or U2689 (N_2689,In_824,In_282);
nor U2690 (N_2690,In_222,In_418);
nand U2691 (N_2691,In_120,In_1307);
and U2692 (N_2692,In_1229,In_1214);
nand U2693 (N_2693,In_470,In_773);
and U2694 (N_2694,In_1290,In_224);
nor U2695 (N_2695,In_1020,In_326);
and U2696 (N_2696,In_384,In_611);
or U2697 (N_2697,In_301,In_1447);
nor U2698 (N_2698,In_742,In_94);
nand U2699 (N_2699,In_690,In_105);
nand U2700 (N_2700,In_1154,In_950);
nor U2701 (N_2701,In_471,In_532);
or U2702 (N_2702,In_940,In_330);
nand U2703 (N_2703,In_1379,In_981);
nand U2704 (N_2704,In_296,In_506);
and U2705 (N_2705,In_504,In_80);
and U2706 (N_2706,In_1188,In_386);
nand U2707 (N_2707,In_941,In_382);
nor U2708 (N_2708,In_715,In_232);
xor U2709 (N_2709,In_1365,In_1269);
or U2710 (N_2710,In_811,In_1291);
and U2711 (N_2711,In_499,In_233);
nor U2712 (N_2712,In_1099,In_284);
or U2713 (N_2713,In_738,In_270);
nor U2714 (N_2714,In_1455,In_334);
xnor U2715 (N_2715,In_557,In_165);
nor U2716 (N_2716,In_1150,In_558);
or U2717 (N_2717,In_410,In_742);
nand U2718 (N_2718,In_472,In_516);
nand U2719 (N_2719,In_997,In_1222);
or U2720 (N_2720,In_377,In_1379);
nand U2721 (N_2721,In_1310,In_935);
nor U2722 (N_2722,In_1389,In_248);
or U2723 (N_2723,In_748,In_824);
nor U2724 (N_2724,In_1239,In_1485);
or U2725 (N_2725,In_741,In_542);
nor U2726 (N_2726,In_832,In_0);
xor U2727 (N_2727,In_1457,In_734);
or U2728 (N_2728,In_452,In_1077);
or U2729 (N_2729,In_1009,In_849);
and U2730 (N_2730,In_591,In_331);
nand U2731 (N_2731,In_895,In_1118);
nor U2732 (N_2732,In_1207,In_925);
and U2733 (N_2733,In_1120,In_1121);
and U2734 (N_2734,In_136,In_686);
or U2735 (N_2735,In_191,In_1067);
nand U2736 (N_2736,In_1485,In_1342);
and U2737 (N_2737,In_907,In_875);
or U2738 (N_2738,In_332,In_509);
nor U2739 (N_2739,In_1402,In_549);
nor U2740 (N_2740,In_237,In_384);
nor U2741 (N_2741,In_448,In_324);
nand U2742 (N_2742,In_787,In_830);
nor U2743 (N_2743,In_201,In_520);
and U2744 (N_2744,In_1224,In_749);
or U2745 (N_2745,In_1411,In_632);
or U2746 (N_2746,In_393,In_313);
and U2747 (N_2747,In_602,In_1485);
nand U2748 (N_2748,In_273,In_1301);
nand U2749 (N_2749,In_412,In_911);
nor U2750 (N_2750,In_978,In_1381);
and U2751 (N_2751,In_1412,In_1390);
and U2752 (N_2752,In_1281,In_1025);
nand U2753 (N_2753,In_62,In_456);
nor U2754 (N_2754,In_1274,In_150);
or U2755 (N_2755,In_751,In_37);
and U2756 (N_2756,In_527,In_818);
nand U2757 (N_2757,In_447,In_153);
nand U2758 (N_2758,In_547,In_43);
nand U2759 (N_2759,In_97,In_1430);
nor U2760 (N_2760,In_917,In_218);
and U2761 (N_2761,In_1304,In_421);
and U2762 (N_2762,In_1261,In_1389);
nor U2763 (N_2763,In_677,In_1311);
nand U2764 (N_2764,In_1030,In_1107);
or U2765 (N_2765,In_1362,In_74);
and U2766 (N_2766,In_1140,In_1265);
nand U2767 (N_2767,In_757,In_336);
nor U2768 (N_2768,In_1081,In_133);
nor U2769 (N_2769,In_529,In_1386);
or U2770 (N_2770,In_690,In_1068);
nor U2771 (N_2771,In_876,In_47);
or U2772 (N_2772,In_669,In_1465);
or U2773 (N_2773,In_309,In_161);
and U2774 (N_2774,In_1211,In_380);
or U2775 (N_2775,In_779,In_1402);
nand U2776 (N_2776,In_117,In_333);
nand U2777 (N_2777,In_427,In_572);
or U2778 (N_2778,In_74,In_390);
nand U2779 (N_2779,In_96,In_545);
or U2780 (N_2780,In_141,In_290);
nor U2781 (N_2781,In_1266,In_61);
and U2782 (N_2782,In_1398,In_1119);
nor U2783 (N_2783,In_546,In_1423);
or U2784 (N_2784,In_1003,In_333);
or U2785 (N_2785,In_136,In_1181);
nand U2786 (N_2786,In_1096,In_632);
nor U2787 (N_2787,In_788,In_1030);
and U2788 (N_2788,In_1147,In_1162);
nor U2789 (N_2789,In_721,In_350);
and U2790 (N_2790,In_680,In_370);
or U2791 (N_2791,In_1397,In_608);
and U2792 (N_2792,In_1249,In_304);
and U2793 (N_2793,In_389,In_1395);
nor U2794 (N_2794,In_826,In_110);
nor U2795 (N_2795,In_1474,In_620);
or U2796 (N_2796,In_1278,In_625);
or U2797 (N_2797,In_312,In_72);
nor U2798 (N_2798,In_1269,In_368);
nand U2799 (N_2799,In_978,In_912);
nand U2800 (N_2800,In_66,In_1017);
nor U2801 (N_2801,In_1496,In_179);
or U2802 (N_2802,In_602,In_596);
nand U2803 (N_2803,In_782,In_1496);
nand U2804 (N_2804,In_699,In_944);
or U2805 (N_2805,In_374,In_1181);
nand U2806 (N_2806,In_838,In_162);
nand U2807 (N_2807,In_272,In_1194);
nor U2808 (N_2808,In_529,In_428);
nor U2809 (N_2809,In_200,In_826);
nor U2810 (N_2810,In_1439,In_483);
nor U2811 (N_2811,In_642,In_479);
nand U2812 (N_2812,In_1272,In_1399);
and U2813 (N_2813,In_910,In_704);
nor U2814 (N_2814,In_852,In_1298);
nor U2815 (N_2815,In_284,In_757);
and U2816 (N_2816,In_12,In_805);
nand U2817 (N_2817,In_272,In_1366);
or U2818 (N_2818,In_1089,In_359);
nand U2819 (N_2819,In_441,In_777);
and U2820 (N_2820,In_972,In_113);
and U2821 (N_2821,In_940,In_458);
or U2822 (N_2822,In_956,In_747);
or U2823 (N_2823,In_604,In_150);
nand U2824 (N_2824,In_1161,In_237);
and U2825 (N_2825,In_1364,In_583);
and U2826 (N_2826,In_516,In_635);
nand U2827 (N_2827,In_489,In_373);
nand U2828 (N_2828,In_311,In_1020);
and U2829 (N_2829,In_632,In_935);
xnor U2830 (N_2830,In_47,In_1144);
nand U2831 (N_2831,In_1365,In_1283);
nor U2832 (N_2832,In_1236,In_358);
nand U2833 (N_2833,In_58,In_1278);
or U2834 (N_2834,In_1405,In_199);
or U2835 (N_2835,In_728,In_1388);
nand U2836 (N_2836,In_1219,In_947);
and U2837 (N_2837,In_1,In_1454);
and U2838 (N_2838,In_397,In_895);
nor U2839 (N_2839,In_90,In_1220);
or U2840 (N_2840,In_220,In_1089);
nor U2841 (N_2841,In_831,In_1279);
or U2842 (N_2842,In_1364,In_354);
nor U2843 (N_2843,In_673,In_804);
or U2844 (N_2844,In_1057,In_1303);
or U2845 (N_2845,In_1486,In_1002);
or U2846 (N_2846,In_202,In_128);
and U2847 (N_2847,In_377,In_1036);
or U2848 (N_2848,In_1489,In_826);
nor U2849 (N_2849,In_1321,In_449);
or U2850 (N_2850,In_802,In_1345);
nor U2851 (N_2851,In_760,In_585);
xor U2852 (N_2852,In_1169,In_1181);
or U2853 (N_2853,In_1450,In_843);
nor U2854 (N_2854,In_610,In_384);
or U2855 (N_2855,In_1475,In_235);
nand U2856 (N_2856,In_527,In_1068);
and U2857 (N_2857,In_1114,In_435);
and U2858 (N_2858,In_178,In_1067);
nand U2859 (N_2859,In_78,In_182);
nor U2860 (N_2860,In_1046,In_1491);
nand U2861 (N_2861,In_31,In_362);
or U2862 (N_2862,In_1022,In_1288);
nand U2863 (N_2863,In_501,In_992);
nor U2864 (N_2864,In_1095,In_725);
and U2865 (N_2865,In_853,In_209);
and U2866 (N_2866,In_776,In_388);
and U2867 (N_2867,In_1209,In_1451);
and U2868 (N_2868,In_1407,In_1422);
nor U2869 (N_2869,In_225,In_1442);
or U2870 (N_2870,In_253,In_988);
or U2871 (N_2871,In_680,In_385);
nand U2872 (N_2872,In_655,In_1205);
and U2873 (N_2873,In_918,In_1375);
and U2874 (N_2874,In_1127,In_678);
and U2875 (N_2875,In_1011,In_477);
and U2876 (N_2876,In_97,In_104);
nor U2877 (N_2877,In_1075,In_1220);
or U2878 (N_2878,In_1060,In_92);
or U2879 (N_2879,In_669,In_1352);
nor U2880 (N_2880,In_1319,In_557);
or U2881 (N_2881,In_9,In_1393);
nand U2882 (N_2882,In_187,In_607);
nand U2883 (N_2883,In_904,In_1337);
nand U2884 (N_2884,In_188,In_1349);
or U2885 (N_2885,In_310,In_58);
and U2886 (N_2886,In_905,In_832);
nand U2887 (N_2887,In_227,In_1258);
or U2888 (N_2888,In_180,In_1145);
nor U2889 (N_2889,In_1350,In_132);
nand U2890 (N_2890,In_265,In_374);
nand U2891 (N_2891,In_1282,In_743);
nand U2892 (N_2892,In_197,In_969);
nor U2893 (N_2893,In_1366,In_227);
nand U2894 (N_2894,In_1463,In_264);
and U2895 (N_2895,In_832,In_1010);
or U2896 (N_2896,In_822,In_534);
or U2897 (N_2897,In_91,In_431);
nand U2898 (N_2898,In_1156,In_1382);
nand U2899 (N_2899,In_926,In_44);
nor U2900 (N_2900,In_302,In_385);
xnor U2901 (N_2901,In_1308,In_356);
nor U2902 (N_2902,In_1175,In_1454);
or U2903 (N_2903,In_593,In_947);
nor U2904 (N_2904,In_588,In_1481);
and U2905 (N_2905,In_135,In_94);
and U2906 (N_2906,In_1457,In_791);
nor U2907 (N_2907,In_999,In_991);
or U2908 (N_2908,In_916,In_504);
and U2909 (N_2909,In_334,In_677);
and U2910 (N_2910,In_484,In_1293);
nor U2911 (N_2911,In_1262,In_1329);
nand U2912 (N_2912,In_659,In_366);
and U2913 (N_2913,In_196,In_759);
nor U2914 (N_2914,In_279,In_781);
nand U2915 (N_2915,In_455,In_90);
nand U2916 (N_2916,In_1319,In_1468);
and U2917 (N_2917,In_477,In_752);
nand U2918 (N_2918,In_1198,In_1367);
nor U2919 (N_2919,In_670,In_483);
nand U2920 (N_2920,In_122,In_155);
nand U2921 (N_2921,In_654,In_522);
nand U2922 (N_2922,In_1187,In_901);
nand U2923 (N_2923,In_860,In_91);
nand U2924 (N_2924,In_330,In_1053);
or U2925 (N_2925,In_551,In_1493);
and U2926 (N_2926,In_136,In_301);
or U2927 (N_2927,In_86,In_1118);
and U2928 (N_2928,In_1112,In_503);
nor U2929 (N_2929,In_444,In_749);
nor U2930 (N_2930,In_1372,In_1471);
nor U2931 (N_2931,In_1150,In_1266);
or U2932 (N_2932,In_413,In_476);
nor U2933 (N_2933,In_1054,In_706);
or U2934 (N_2934,In_1091,In_881);
and U2935 (N_2935,In_606,In_672);
and U2936 (N_2936,In_148,In_1286);
nor U2937 (N_2937,In_744,In_224);
and U2938 (N_2938,In_319,In_381);
or U2939 (N_2939,In_573,In_9);
nor U2940 (N_2940,In_380,In_71);
and U2941 (N_2941,In_1059,In_830);
nor U2942 (N_2942,In_120,In_1161);
or U2943 (N_2943,In_354,In_1339);
or U2944 (N_2944,In_49,In_1233);
or U2945 (N_2945,In_476,In_210);
nor U2946 (N_2946,In_293,In_820);
nand U2947 (N_2947,In_1381,In_973);
or U2948 (N_2948,In_1252,In_466);
or U2949 (N_2949,In_278,In_476);
nor U2950 (N_2950,In_96,In_1130);
nor U2951 (N_2951,In_264,In_369);
and U2952 (N_2952,In_852,In_96);
or U2953 (N_2953,In_795,In_1076);
and U2954 (N_2954,In_120,In_1434);
and U2955 (N_2955,In_432,In_1223);
and U2956 (N_2956,In_29,In_90);
and U2957 (N_2957,In_959,In_1271);
nor U2958 (N_2958,In_1457,In_192);
and U2959 (N_2959,In_845,In_149);
or U2960 (N_2960,In_16,In_682);
nor U2961 (N_2961,In_921,In_806);
and U2962 (N_2962,In_1279,In_408);
or U2963 (N_2963,In_917,In_1011);
and U2964 (N_2964,In_1077,In_1240);
nor U2965 (N_2965,In_306,In_1164);
nand U2966 (N_2966,In_607,In_1401);
or U2967 (N_2967,In_1417,In_391);
nand U2968 (N_2968,In_410,In_338);
or U2969 (N_2969,In_258,In_1004);
nand U2970 (N_2970,In_216,In_20);
or U2971 (N_2971,In_674,In_634);
and U2972 (N_2972,In_471,In_272);
and U2973 (N_2973,In_997,In_386);
or U2974 (N_2974,In_768,In_1199);
nand U2975 (N_2975,In_411,In_525);
nor U2976 (N_2976,In_30,In_606);
nand U2977 (N_2977,In_809,In_306);
nor U2978 (N_2978,In_273,In_1042);
or U2979 (N_2979,In_327,In_1492);
or U2980 (N_2980,In_1100,In_1136);
and U2981 (N_2981,In_57,In_32);
and U2982 (N_2982,In_457,In_819);
nor U2983 (N_2983,In_925,In_1429);
nor U2984 (N_2984,In_306,In_1240);
or U2985 (N_2985,In_866,In_1352);
and U2986 (N_2986,In_809,In_41);
xnor U2987 (N_2987,In_165,In_409);
nand U2988 (N_2988,In_87,In_48);
and U2989 (N_2989,In_369,In_1104);
nor U2990 (N_2990,In_1428,In_1300);
and U2991 (N_2991,In_713,In_276);
nand U2992 (N_2992,In_541,In_845);
or U2993 (N_2993,In_1429,In_798);
or U2994 (N_2994,In_308,In_696);
nor U2995 (N_2995,In_615,In_442);
xnor U2996 (N_2996,In_957,In_369);
and U2997 (N_2997,In_52,In_459);
nor U2998 (N_2998,In_168,In_1484);
or U2999 (N_2999,In_856,In_102);
nand U3000 (N_3000,N_1889,N_2353);
nor U3001 (N_3001,N_1974,N_2879);
nand U3002 (N_3002,N_2478,N_522);
nand U3003 (N_3003,N_858,N_2578);
nand U3004 (N_3004,N_870,N_785);
or U3005 (N_3005,N_87,N_1755);
and U3006 (N_3006,N_2800,N_1830);
nor U3007 (N_3007,N_1058,N_2477);
nand U3008 (N_3008,N_1206,N_2395);
nand U3009 (N_3009,N_1170,N_2877);
nor U3010 (N_3010,N_2699,N_66);
and U3011 (N_3011,N_67,N_1727);
or U3012 (N_3012,N_49,N_400);
and U3013 (N_3013,N_2845,N_2666);
or U3014 (N_3014,N_1386,N_2871);
or U3015 (N_3015,N_1975,N_947);
nand U3016 (N_3016,N_2865,N_2282);
nand U3017 (N_3017,N_1185,N_1722);
and U3018 (N_3018,N_1420,N_2721);
and U3019 (N_3019,N_876,N_1355);
nor U3020 (N_3020,N_1071,N_1231);
and U3021 (N_3021,N_651,N_948);
nand U3022 (N_3022,N_1546,N_2708);
nor U3023 (N_3023,N_2911,N_2499);
or U3024 (N_3024,N_1258,N_1073);
and U3025 (N_3025,N_2894,N_2370);
nand U3026 (N_3026,N_2133,N_2029);
or U3027 (N_3027,N_1048,N_145);
nand U3028 (N_3028,N_728,N_850);
or U3029 (N_3029,N_1262,N_1280);
and U3030 (N_3030,N_1610,N_226);
or U3031 (N_3031,N_1516,N_1772);
nand U3032 (N_3032,N_410,N_559);
nor U3033 (N_3033,N_177,N_2585);
nand U3034 (N_3034,N_2461,N_2050);
or U3035 (N_3035,N_1271,N_756);
and U3036 (N_3036,N_2648,N_926);
and U3037 (N_3037,N_196,N_761);
nand U3038 (N_3038,N_332,N_2143);
nand U3039 (N_3039,N_1899,N_442);
and U3040 (N_3040,N_1393,N_1898);
nor U3041 (N_3041,N_1362,N_1462);
or U3042 (N_3042,N_2259,N_1587);
or U3043 (N_3043,N_1200,N_1857);
nand U3044 (N_3044,N_816,N_1361);
nand U3045 (N_3045,N_1490,N_626);
nand U3046 (N_3046,N_1669,N_313);
nand U3047 (N_3047,N_152,N_2434);
nand U3048 (N_3048,N_1695,N_1913);
and U3049 (N_3049,N_1756,N_1227);
nor U3050 (N_3050,N_1652,N_999);
and U3051 (N_3051,N_781,N_2175);
or U3052 (N_3052,N_923,N_264);
or U3053 (N_3053,N_2298,N_757);
nor U3054 (N_3054,N_1173,N_2681);
xor U3055 (N_3055,N_2830,N_810);
or U3056 (N_3056,N_1298,N_2092);
or U3057 (N_3057,N_1762,N_1665);
nor U3058 (N_3058,N_1860,N_978);
nand U3059 (N_3059,N_298,N_979);
or U3060 (N_3060,N_1731,N_981);
and U3061 (N_3061,N_603,N_358);
nand U3062 (N_3062,N_1395,N_1670);
nor U3063 (N_3063,N_1633,N_2854);
and U3064 (N_3064,N_2178,N_1525);
and U3065 (N_3065,N_2159,N_1673);
nand U3066 (N_3066,N_1667,N_2073);
nand U3067 (N_3067,N_1703,N_581);
or U3068 (N_3068,N_1776,N_753);
or U3069 (N_3069,N_153,N_782);
nand U3070 (N_3070,N_17,N_2437);
nor U3071 (N_3071,N_2527,N_1149);
nand U3072 (N_3072,N_2546,N_1216);
and U3073 (N_3073,N_1916,N_2669);
or U3074 (N_3074,N_470,N_63);
nand U3075 (N_3075,N_1981,N_1246);
nand U3076 (N_3076,N_1556,N_2943);
or U3077 (N_3077,N_2561,N_1907);
and U3078 (N_3078,N_174,N_2025);
nor U3079 (N_3079,N_1557,N_2064);
nor U3080 (N_3080,N_92,N_157);
and U3081 (N_3081,N_2179,N_959);
nand U3082 (N_3082,N_2704,N_563);
and U3083 (N_3083,N_2797,N_2947);
nand U3084 (N_3084,N_1661,N_2929);
nand U3085 (N_3085,N_2422,N_1145);
or U3086 (N_3086,N_1708,N_2433);
and U3087 (N_3087,N_593,N_1492);
and U3088 (N_3088,N_1630,N_2827);
nor U3089 (N_3089,N_875,N_2731);
or U3090 (N_3090,N_1010,N_57);
nor U3091 (N_3091,N_510,N_1896);
nor U3092 (N_3092,N_2058,N_2835);
and U3093 (N_3093,N_282,N_1915);
and U3094 (N_3094,N_2631,N_2195);
and U3095 (N_3095,N_2791,N_2022);
nand U3096 (N_3096,N_1653,N_1162);
nand U3097 (N_3097,N_2444,N_2331);
nand U3098 (N_3098,N_369,N_2120);
nor U3099 (N_3099,N_1549,N_241);
or U3100 (N_3100,N_121,N_1107);
nand U3101 (N_3101,N_5,N_2200);
nor U3102 (N_3102,N_2584,N_279);
and U3103 (N_3103,N_1257,N_300);
and U3104 (N_3104,N_2861,N_740);
nor U3105 (N_3105,N_1991,N_2095);
or U3106 (N_3106,N_420,N_597);
or U3107 (N_3107,N_1187,N_840);
or U3108 (N_3108,N_129,N_1690);
nor U3109 (N_3109,N_1779,N_2644);
and U3110 (N_3110,N_1958,N_1956);
nand U3111 (N_3111,N_221,N_1158);
nor U3112 (N_3112,N_819,N_1802);
nand U3113 (N_3113,N_2608,N_443);
nor U3114 (N_3114,N_1485,N_1237);
or U3115 (N_3115,N_2933,N_1963);
and U3116 (N_3116,N_1303,N_336);
nand U3117 (N_3117,N_1848,N_835);
or U3118 (N_3118,N_2295,N_565);
nand U3119 (N_3119,N_2512,N_1521);
and U3120 (N_3120,N_582,N_2198);
or U3121 (N_3121,N_1182,N_454);
nor U3122 (N_3122,N_1012,N_898);
or U3123 (N_3123,N_992,N_1276);
or U3124 (N_3124,N_382,N_1259);
nand U3125 (N_3125,N_1918,N_186);
nand U3126 (N_3126,N_552,N_708);
nand U3127 (N_3127,N_1183,N_2606);
or U3128 (N_3128,N_2937,N_1838);
nand U3129 (N_3129,N_921,N_1438);
nor U3130 (N_3130,N_2513,N_2408);
nand U3131 (N_3131,N_1191,N_2051);
and U3132 (N_3132,N_1030,N_2128);
and U3133 (N_3133,N_422,N_2919);
nor U3134 (N_3134,N_644,N_861);
nand U3135 (N_3135,N_2878,N_2390);
or U3136 (N_3136,N_2418,N_222);
and U3137 (N_3137,N_1637,N_2296);
and U3138 (N_3138,N_633,N_2468);
nand U3139 (N_3139,N_14,N_1548);
nor U3140 (N_3140,N_2132,N_2172);
and U3141 (N_3141,N_623,N_2785);
nor U3142 (N_3142,N_2983,N_2490);
and U3143 (N_3143,N_2221,N_368);
or U3144 (N_3144,N_913,N_668);
nor U3145 (N_3145,N_2743,N_546);
or U3146 (N_3146,N_2326,N_2484);
and U3147 (N_3147,N_1657,N_2890);
and U3148 (N_3148,N_1108,N_1202);
nor U3149 (N_3149,N_726,N_2735);
nand U3150 (N_3150,N_1207,N_705);
and U3151 (N_3151,N_138,N_931);
or U3152 (N_3152,N_415,N_886);
nor U3153 (N_3153,N_1424,N_354);
or U3154 (N_3154,N_229,N_2057);
nand U3155 (N_3155,N_692,N_1301);
or U3156 (N_3156,N_1687,N_2416);
or U3157 (N_3157,N_2424,N_2385);
and U3158 (N_3158,N_1363,N_1510);
or U3159 (N_3159,N_2403,N_1810);
or U3160 (N_3160,N_2944,N_1478);
nand U3161 (N_3161,N_1486,N_1384);
nor U3162 (N_3162,N_440,N_2473);
and U3163 (N_3163,N_1847,N_2246);
nand U3164 (N_3164,N_1558,N_945);
nand U3165 (N_3165,N_854,N_2149);
and U3166 (N_3166,N_1319,N_1423);
nor U3167 (N_3167,N_398,N_2375);
nand U3168 (N_3168,N_2528,N_102);
nor U3169 (N_3169,N_2469,N_2517);
and U3170 (N_3170,N_1564,N_845);
nor U3171 (N_3171,N_918,N_862);
nor U3172 (N_3172,N_2253,N_1960);
nand U3173 (N_3173,N_2849,N_419);
nor U3174 (N_3174,N_1534,N_637);
and U3175 (N_3175,N_2828,N_492);
nor U3176 (N_3176,N_1150,N_1225);
nand U3177 (N_3177,N_1938,N_169);
and U3178 (N_3178,N_215,N_2237);
nor U3179 (N_3179,N_339,N_2448);
and U3180 (N_3180,N_796,N_1201);
nor U3181 (N_3181,N_54,N_2601);
nor U3182 (N_3182,N_1452,N_2746);
nand U3183 (N_3183,N_2376,N_2244);
nand U3184 (N_3184,N_2492,N_1003);
or U3185 (N_3185,N_2641,N_1948);
or U3186 (N_3186,N_455,N_0);
and U3187 (N_3187,N_2667,N_908);
nor U3188 (N_3188,N_2479,N_1013);
nand U3189 (N_3189,N_749,N_334);
and U3190 (N_3190,N_1748,N_1935);
nor U3191 (N_3191,N_2323,N_2303);
and U3192 (N_3192,N_162,N_1563);
or U3193 (N_3193,N_1582,N_1055);
nand U3194 (N_3194,N_89,N_2124);
or U3195 (N_3195,N_137,N_930);
nor U3196 (N_3196,N_2851,N_1575);
nor U3197 (N_3197,N_1087,N_319);
nand U3198 (N_3198,N_2536,N_2062);
and U3199 (N_3199,N_317,N_2779);
and U3200 (N_3200,N_2278,N_2084);
or U3201 (N_3201,N_2700,N_905);
or U3202 (N_3202,N_1160,N_122);
nor U3203 (N_3203,N_1815,N_78);
nor U3204 (N_3204,N_2491,N_1577);
nor U3205 (N_3205,N_2355,N_1743);
nor U3206 (N_3206,N_1904,N_402);
or U3207 (N_3207,N_2640,N_2060);
nand U3208 (N_3208,N_1944,N_1518);
or U3209 (N_3209,N_343,N_961);
or U3210 (N_3210,N_1936,N_950);
or U3211 (N_3211,N_1451,N_537);
nand U3212 (N_3212,N_2948,N_2297);
and U3213 (N_3213,N_715,N_1103);
and U3214 (N_3214,N_34,N_2284);
and U3215 (N_3215,N_276,N_1953);
and U3216 (N_3216,N_718,N_1950);
and U3217 (N_3217,N_1494,N_1052);
and U3218 (N_3218,N_1072,N_399);
or U3219 (N_3219,N_2466,N_101);
nor U3220 (N_3220,N_268,N_2405);
nand U3221 (N_3221,N_2428,N_526);
nand U3222 (N_3222,N_1428,N_1900);
nand U3223 (N_3223,N_2262,N_1647);
nand U3224 (N_3224,N_1537,N_736);
or U3225 (N_3225,N_2472,N_2519);
and U3226 (N_3226,N_887,N_325);
and U3227 (N_3227,N_1120,N_1374);
and U3228 (N_3228,N_2410,N_2141);
and U3229 (N_3229,N_1749,N_2985);
or U3230 (N_3230,N_2264,N_2888);
or U3231 (N_3231,N_2191,N_1672);
or U3232 (N_3232,N_1870,N_1837);
nand U3233 (N_3233,N_2327,N_857);
nor U3234 (N_3234,N_249,N_1268);
nand U3235 (N_3235,N_2104,N_1193);
nor U3236 (N_3236,N_1260,N_344);
nand U3237 (N_3237,N_2006,N_780);
nand U3238 (N_3238,N_2995,N_1952);
and U3239 (N_3239,N_949,N_2151);
nand U3240 (N_3240,N_1400,N_2949);
nand U3241 (N_3241,N_386,N_706);
nor U3242 (N_3242,N_1750,N_2197);
nand U3243 (N_3243,N_2841,N_1228);
and U3244 (N_3244,N_1240,N_449);
and U3245 (N_3245,N_613,N_1562);
and U3246 (N_3246,N_306,N_2567);
nand U3247 (N_3247,N_2824,N_484);
and U3248 (N_3248,N_451,N_1514);
or U3249 (N_3249,N_2885,N_1371);
nor U3250 (N_3250,N_864,N_2599);
and U3251 (N_3251,N_2440,N_573);
or U3252 (N_3252,N_1224,N_2308);
and U3253 (N_3253,N_1942,N_1538);
or U3254 (N_3254,N_1157,N_2842);
nand U3255 (N_3255,N_2127,N_444);
nor U3256 (N_3256,N_1382,N_2624);
or U3257 (N_3257,N_481,N_1972);
and U3258 (N_3258,N_1794,N_2533);
nor U3259 (N_3259,N_1329,N_2286);
nor U3260 (N_3260,N_280,N_647);
and U3261 (N_3261,N_700,N_1891);
or U3262 (N_3262,N_2635,N_837);
nor U3263 (N_3263,N_2347,N_250);
or U3264 (N_3264,N_2103,N_2320);
nand U3265 (N_3265,N_2153,N_189);
xnor U3266 (N_3266,N_1014,N_2125);
nand U3267 (N_3267,N_760,N_2531);
nor U3268 (N_3268,N_889,N_1528);
nand U3269 (N_3269,N_534,N_826);
and U3270 (N_3270,N_2928,N_2381);
nor U3271 (N_3271,N_1926,N_1914);
nand U3272 (N_3272,N_2116,N_2652);
or U3273 (N_3273,N_355,N_1310);
nand U3274 (N_3274,N_925,N_480);
nand U3275 (N_3275,N_1666,N_624);
nor U3276 (N_3276,N_823,N_1807);
nor U3277 (N_3277,N_2031,N_2692);
and U3278 (N_3278,N_2660,N_1739);
nor U3279 (N_3279,N_192,N_535);
nand U3280 (N_3280,N_664,N_496);
and U3281 (N_3281,N_1504,N_427);
or U3282 (N_3282,N_920,N_397);
nand U3283 (N_3283,N_1990,N_2001);
nand U3284 (N_3284,N_1385,N_2958);
or U3285 (N_3285,N_97,N_424);
and U3286 (N_3286,N_487,N_634);
and U3287 (N_3287,N_2535,N_1892);
nor U3288 (N_3288,N_2532,N_1047);
nor U3289 (N_3289,N_435,N_1317);
or U3290 (N_3290,N_2754,N_1982);
nand U3291 (N_3291,N_2497,N_1497);
nand U3292 (N_3292,N_119,N_2275);
nor U3293 (N_3293,N_2110,N_1316);
and U3294 (N_3294,N_1442,N_232);
nor U3295 (N_3295,N_1897,N_2974);
and U3296 (N_3296,N_2065,N_2993);
nor U3297 (N_3297,N_163,N_860);
or U3298 (N_3298,N_1941,N_769);
or U3299 (N_3299,N_236,N_969);
and U3300 (N_3300,N_612,N_1281);
and U3301 (N_3301,N_1234,N_778);
nand U3302 (N_3302,N_1080,N_1894);
or U3303 (N_3303,N_1997,N_271);
or U3304 (N_3304,N_562,N_1861);
or U3305 (N_3305,N_1311,N_1463);
and U3306 (N_3306,N_1920,N_323);
nor U3307 (N_3307,N_606,N_1226);
or U3308 (N_3308,N_373,N_523);
nand U3309 (N_3309,N_2138,N_18);
nand U3310 (N_3310,N_2054,N_880);
nor U3311 (N_3311,N_1621,N_1416);
or U3312 (N_3312,N_902,N_2024);
or U3313 (N_3313,N_1279,N_431);
nand U3314 (N_3314,N_40,N_1684);
or U3315 (N_3315,N_1314,N_1369);
and U3316 (N_3316,N_2679,N_204);
and U3317 (N_3317,N_791,N_2514);
or U3318 (N_3318,N_1426,N_2579);
or U3319 (N_3319,N_2285,N_10);
or U3320 (N_3320,N_2097,N_305);
or U3321 (N_3321,N_1778,N_790);
and U3322 (N_3322,N_594,N_2653);
or U3323 (N_3323,N_1152,N_2088);
or U3324 (N_3324,N_1979,N_730);
or U3325 (N_3325,N_1509,N_517);
and U3326 (N_3326,N_1906,N_91);
and U3327 (N_3327,N_805,N_2122);
nor U3328 (N_3328,N_2494,N_2654);
or U3329 (N_3329,N_2174,N_1741);
nand U3330 (N_3330,N_1836,N_659);
nor U3331 (N_3331,N_2926,N_1996);
and U3332 (N_3332,N_1334,N_1378);
nor U3333 (N_3333,N_2611,N_1984);
and U3334 (N_3334,N_2615,N_2118);
nor U3335 (N_3335,N_787,N_1931);
nor U3336 (N_3336,N_472,N_2836);
or U3337 (N_3337,N_2475,N_1269);
nand U3338 (N_3338,N_2977,N_916);
nor U3339 (N_3339,N_1589,N_2881);
nor U3340 (N_3340,N_425,N_1024);
nor U3341 (N_3341,N_1088,N_669);
nand U3342 (N_3342,N_1406,N_1542);
or U3343 (N_3343,N_1817,N_672);
nand U3344 (N_3344,N_1590,N_2619);
or U3345 (N_3345,N_493,N_1023);
and U3346 (N_3346,N_338,N_2866);
nand U3347 (N_3347,N_1214,N_1685);
and U3348 (N_3348,N_1598,N_783);
nand U3349 (N_3349,N_1039,N_2657);
nor U3350 (N_3350,N_863,N_2167);
and U3351 (N_3351,N_883,N_2239);
nor U3352 (N_3352,N_108,N_2821);
nand U3353 (N_3353,N_1218,N_795);
and U3354 (N_3354,N_1694,N_2598);
nor U3355 (N_3355,N_497,N_1128);
xnor U3356 (N_3356,N_2157,N_463);
nand U3357 (N_3357,N_909,N_2566);
nor U3358 (N_3358,N_698,N_2117);
nor U3359 (N_3359,N_1089,N_642);
nand U3360 (N_3360,N_1714,N_1874);
nand U3361 (N_3361,N_2554,N_235);
nor U3362 (N_3362,N_1219,N_2685);
or U3363 (N_3363,N_246,N_2794);
nor U3364 (N_3364,N_2719,N_2511);
nor U3365 (N_3365,N_15,N_2233);
nand U3366 (N_3366,N_2155,N_245);
or U3367 (N_3367,N_1713,N_2720);
nor U3368 (N_3368,N_813,N_1266);
nand U3369 (N_3369,N_846,N_971);
nand U3370 (N_3370,N_311,N_190);
nand U3371 (N_3371,N_1069,N_2306);
or U3372 (N_3372,N_670,N_2753);
nand U3373 (N_3373,N_1844,N_1354);
or U3374 (N_3374,N_2504,N_2569);
xnor U3375 (N_3375,N_1761,N_1964);
and U3376 (N_3376,N_1866,N_123);
nor U3377 (N_3377,N_1040,N_2377);
or U3378 (N_3378,N_1640,N_2850);
or U3379 (N_3379,N_1342,N_2789);
nor U3380 (N_3380,N_2238,N_1278);
nand U3381 (N_3381,N_1284,N_1196);
nor U3382 (N_3382,N_1181,N_1768);
and U3383 (N_3383,N_662,N_699);
nand U3384 (N_3384,N_966,N_627);
xor U3385 (N_3385,N_2603,N_746);
and U3386 (N_3386,N_1238,N_1360);
or U3387 (N_3387,N_1554,N_2371);
nand U3388 (N_3388,N_1131,N_935);
nand U3389 (N_3389,N_2391,N_1007);
or U3390 (N_3390,N_166,N_2177);
or U3391 (N_3391,N_2651,N_2819);
and U3392 (N_3392,N_2560,N_2939);
nor U3393 (N_3393,N_2904,N_893);
or U3394 (N_3394,N_86,N_1033);
nor U3395 (N_3395,N_2814,N_2623);
nor U3396 (N_3396,N_2730,N_2212);
and U3397 (N_3397,N_515,N_1458);
and U3398 (N_3398,N_641,N_2452);
nand U3399 (N_3399,N_2781,N_2425);
and U3400 (N_3400,N_1068,N_963);
nor U3401 (N_3401,N_2963,N_366);
nand U3402 (N_3402,N_1507,N_75);
xor U3403 (N_3403,N_2843,N_172);
nor U3404 (N_3404,N_441,N_1300);
nand U3405 (N_3405,N_1883,N_297);
nor U3406 (N_3406,N_944,N_1992);
or U3407 (N_3407,N_460,N_2067);
nor U3408 (N_3408,N_1567,N_1327);
nand U3409 (N_3409,N_2261,N_116);
nand U3410 (N_3410,N_1511,N_1951);
or U3411 (N_3411,N_2301,N_148);
and U3412 (N_3412,N_259,N_2277);
and U3413 (N_3413,N_495,N_1512);
nor U3414 (N_3414,N_1774,N_2208);
and U3415 (N_3415,N_622,N_1878);
or U3416 (N_3416,N_743,N_302);
or U3417 (N_3417,N_1432,N_1985);
or U3418 (N_3418,N_2248,N_1176);
nor U3419 (N_3419,N_147,N_1011);
nor U3420 (N_3420,N_434,N_2417);
nor U3421 (N_3421,N_1102,N_389);
nor U3422 (N_3422,N_173,N_486);
and U3423 (N_3423,N_1292,N_541);
and U3424 (N_3424,N_1862,N_2094);
nor U3425 (N_3425,N_2279,N_2485);
nor U3426 (N_3426,N_2017,N_1308);
and U3427 (N_3427,N_680,N_1345);
and U3428 (N_3428,N_792,N_134);
and U3429 (N_3429,N_1184,N_2898);
and U3430 (N_3430,N_1328,N_2137);
nand U3431 (N_3431,N_910,N_1403);
or U3432 (N_3432,N_1675,N_2364);
nand U3433 (N_3433,N_2729,N_195);
nor U3434 (N_3434,N_2336,N_136);
nor U3435 (N_3435,N_1453,N_2252);
nor U3436 (N_3436,N_114,N_661);
or U3437 (N_3437,N_2576,N_2581);
nand U3438 (N_3438,N_2972,N_1759);
or U3439 (N_3439,N_1352,N_2852);
nor U3440 (N_3440,N_50,N_142);
nor U3441 (N_3441,N_2673,N_2604);
and U3442 (N_3442,N_2696,N_1045);
nand U3443 (N_3443,N_2691,N_2450);
xor U3444 (N_3444,N_834,N_2883);
nand U3445 (N_3445,N_1457,N_508);
nand U3446 (N_3446,N_2190,N_1656);
nor U3447 (N_3447,N_2243,N_821);
nand U3448 (N_3448,N_1489,N_798);
nor U3449 (N_3449,N_19,N_2792);
nand U3450 (N_3450,N_2610,N_105);
nor U3451 (N_3451,N_2906,N_557);
or U3452 (N_3452,N_2047,N_2021);
nand U3453 (N_3453,N_2161,N_640);
and U3454 (N_3454,N_786,N_1050);
and U3455 (N_3455,N_2053,N_1884);
or U3456 (N_3456,N_1121,N_2069);
and U3457 (N_3457,N_299,N_1454);
and U3458 (N_3458,N_665,N_1295);
or U3459 (N_3459,N_1732,N_1387);
or U3460 (N_3460,N_1042,N_309);
nand U3461 (N_3461,N_2056,N_1429);
and U3462 (N_3462,N_2136,N_2123);
and U3463 (N_3463,N_1026,N_1947);
nand U3464 (N_3464,N_1127,N_877);
nand U3465 (N_3465,N_1074,N_2938);
nor U3466 (N_3466,N_2369,N_1882);
or U3467 (N_3467,N_1811,N_2413);
nor U3468 (N_3468,N_2987,N_2530);
and U3469 (N_3469,N_2107,N_709);
and U3470 (N_3470,N_206,N_135);
or U3471 (N_3471,N_2351,N_303);
or U3472 (N_3472,N_1816,N_1709);
or U3473 (N_3473,N_2209,N_2036);
nor U3474 (N_3474,N_1496,N_1165);
nor U3475 (N_3475,N_912,N_491);
nand U3476 (N_3476,N_1912,N_2981);
or U3477 (N_3477,N_381,N_2358);
and U3478 (N_3478,N_658,N_892);
nor U3479 (N_3479,N_251,N_1283);
nand U3480 (N_3480,N_1998,N_418);
or U3481 (N_3481,N_2488,N_1767);
nor U3482 (N_3482,N_839,N_2634);
or U3483 (N_3483,N_747,N_1287);
nand U3484 (N_3484,N_155,N_531);
nor U3485 (N_3485,N_1044,N_1570);
and U3486 (N_3486,N_2384,N_1795);
nor U3487 (N_3487,N_41,N_1491);
or U3488 (N_3488,N_2379,N_1095);
or U3489 (N_3489,N_2333,N_2897);
or U3490 (N_3490,N_1609,N_1254);
or U3491 (N_3491,N_2962,N_1523);
and U3492 (N_3492,N_2266,N_1006);
nand U3493 (N_3493,N_1500,N_1414);
nor U3494 (N_3494,N_1626,N_1336);
and U3495 (N_3495,N_103,N_1605);
or U3496 (N_3496,N_1976,N_1728);
and U3497 (N_3497,N_2609,N_762);
and U3498 (N_3498,N_836,N_878);
or U3499 (N_3499,N_149,N_733);
and U3500 (N_3500,N_2858,N_1468);
and U3501 (N_3501,N_243,N_1204);
or U3502 (N_3502,N_2749,N_304);
and U3503 (N_3503,N_2171,N_1066);
and U3504 (N_3504,N_1053,N_779);
nand U3505 (N_3505,N_112,N_727);
nand U3506 (N_3506,N_2196,N_2020);
nand U3507 (N_3507,N_1651,N_869);
and U3508 (N_3508,N_227,N_2950);
and U3509 (N_3509,N_802,N_2927);
or U3510 (N_3510,N_988,N_2368);
nand U3511 (N_3511,N_1879,N_296);
nand U3512 (N_3512,N_2147,N_77);
and U3513 (N_3513,N_652,N_673);
or U3514 (N_3514,N_1455,N_2189);
nor U3515 (N_3515,N_2105,N_689);
and U3516 (N_3516,N_1801,N_2955);
and U3517 (N_3517,N_617,N_2205);
and U3518 (N_3518,N_678,N_253);
nand U3519 (N_3519,N_266,N_503);
nor U3520 (N_3520,N_1547,N_1602);
nor U3521 (N_3521,N_527,N_2510);
or U3522 (N_3522,N_281,N_1890);
or U3523 (N_3523,N_2637,N_2052);
nand U3524 (N_3524,N_48,N_750);
or U3525 (N_3525,N_248,N_1330);
nand U3526 (N_3526,N_2755,N_2803);
nor U3527 (N_3527,N_1380,N_540);
and U3528 (N_3528,N_4,N_2255);
or U3529 (N_3529,N_1814,N_499);
nand U3530 (N_3530,N_1388,N_2414);
or U3531 (N_3531,N_1119,N_742);
and U3532 (N_3532,N_1771,N_974);
nand U3533 (N_3533,N_2365,N_2689);
and U3534 (N_3534,N_378,N_532);
nor U3535 (N_3535,N_1773,N_1404);
or U3536 (N_3536,N_2242,N_2495);
or U3537 (N_3537,N_1106,N_2734);
nor U3538 (N_3538,N_842,N_632);
and U3539 (N_3539,N_23,N_2573);
nor U3540 (N_3540,N_71,N_2042);
nand U3541 (N_3541,N_1639,N_2388);
nor U3542 (N_3542,N_506,N_1339);
and U3543 (N_3543,N_198,N_2033);
nand U3544 (N_3544,N_1391,N_409);
nor U3545 (N_3545,N_2675,N_2967);
or U3546 (N_3546,N_514,N_543);
nor U3547 (N_3547,N_849,N_1338);
nor U3548 (N_3548,N_1658,N_85);
nand U3549 (N_3549,N_2760,N_2718);
or U3550 (N_3550,N_489,N_1051);
nor U3551 (N_3551,N_1718,N_1849);
or U3552 (N_3552,N_2330,N_8);
and U3553 (N_3553,N_1909,N_124);
or U3554 (N_3554,N_896,N_2726);
nand U3555 (N_3555,N_1249,N_2961);
or U3556 (N_3556,N_2763,N_2762);
nand U3557 (N_3557,N_1954,N_216);
or U3558 (N_3558,N_2441,N_561);
and U3559 (N_3559,N_2895,N_567);
nand U3560 (N_3560,N_2192,N_474);
nor U3561 (N_3561,N_1169,N_252);
and U3562 (N_3562,N_1635,N_2522);
nand U3563 (N_3563,N_772,N_1480);
nor U3564 (N_3564,N_2896,N_90);
nor U3565 (N_3565,N_1410,N_504);
nor U3566 (N_3566,N_748,N_426);
nor U3567 (N_3567,N_1966,N_1502);
nand U3568 (N_3568,N_345,N_2091);
nand U3569 (N_3569,N_1796,N_2357);
nor U3570 (N_3570,N_738,N_853);
and U3571 (N_3571,N_1584,N_2294);
or U3572 (N_3572,N_1326,N_1190);
nand U3573 (N_3573,N_775,N_994);
nand U3574 (N_3574,N_500,N_566);
and U3575 (N_3575,N_2682,N_392);
or U3576 (N_3576,N_2728,N_1843);
or U3577 (N_3577,N_873,N_2304);
or U3578 (N_3578,N_2975,N_1057);
nand U3579 (N_3579,N_2039,N_2250);
nand U3580 (N_3580,N_2217,N_285);
nand U3581 (N_3581,N_205,N_11);
nand U3582 (N_3582,N_256,N_2582);
nor U3583 (N_3583,N_1986,N_167);
or U3584 (N_3584,N_881,N_1);
nor U3585 (N_3585,N_2335,N_2934);
or U3586 (N_3586,N_2831,N_1545);
nor U3587 (N_3587,N_723,N_62);
or U3588 (N_3588,N_2010,N_1751);
nand U3589 (N_3589,N_571,N_704);
nor U3590 (N_3590,N_833,N_1929);
nor U3591 (N_3591,N_621,N_1501);
or U3592 (N_3592,N_871,N_851);
and U3593 (N_3593,N_653,N_2270);
nand U3594 (N_3594,N_675,N_1725);
nand U3595 (N_3595,N_2586,N_2345);
nor U3596 (N_3596,N_494,N_636);
nor U3597 (N_3597,N_1402,N_2725);
and U3598 (N_3598,N_1681,N_478);
and U3599 (N_3599,N_1090,N_2423);
or U3600 (N_3600,N_1812,N_2483);
nor U3601 (N_3601,N_1934,N_1138);
and U3602 (N_3602,N_2942,N_1729);
or U3603 (N_3603,N_639,N_2957);
and U3604 (N_3604,N_1075,N_716);
nand U3605 (N_3605,N_1076,N_284);
and U3606 (N_3606,N_1302,N_2925);
nor U3607 (N_3607,N_231,N_1965);
nand U3608 (N_3608,N_44,N_1002);
and U3609 (N_3609,N_586,N_1142);
nor U3610 (N_3610,N_884,N_35);
and U3611 (N_3611,N_2748,N_2622);
nand U3612 (N_3612,N_269,N_1677);
nor U3613 (N_3613,N_973,N_2783);
or U3614 (N_3614,N_872,N_1835);
and U3615 (N_3615,N_2770,N_316);
or U3616 (N_3616,N_179,N_1994);
nor U3617 (N_3617,N_754,N_2741);
nor U3618 (N_3618,N_2616,N_1118);
nor U3619 (N_3619,N_1620,N_2230);
nor U3620 (N_3620,N_720,N_2638);
or U3621 (N_3621,N_1818,N_1307);
nor U3622 (N_3622,N_1376,N_1433);
and U3623 (N_3623,N_1484,N_927);
and U3624 (N_3624,N_2283,N_1565);
and U3625 (N_3625,N_310,N_2078);
nand U3626 (N_3626,N_1648,N_712);
nor U3627 (N_3627,N_2193,N_2360);
or U3628 (N_3628,N_53,N_1845);
nor U3629 (N_3629,N_687,N_997);
nor U3630 (N_3630,N_1519,N_784);
or U3631 (N_3631,N_501,N_1146);
nor U3632 (N_3632,N_585,N_879);
nand U3633 (N_3633,N_598,N_224);
nor U3634 (N_3634,N_2325,N_1591);
and U3635 (N_3635,N_1720,N_2886);
nand U3636 (N_3636,N_2817,N_2629);
or U3637 (N_3637,N_550,N_1726);
or U3638 (N_3638,N_1659,N_1241);
and U3639 (N_3639,N_768,N_657);
and U3640 (N_3640,N_2184,N_1806);
nand U3641 (N_3641,N_645,N_439);
and U3642 (N_3642,N_751,N_9);
nor U3643 (N_3643,N_469,N_357);
or U3644 (N_3644,N_1636,N_1389);
nand U3645 (N_3645,N_2612,N_2923);
nor U3646 (N_3646,N_1770,N_2354);
and U3647 (N_3647,N_807,N_43);
nor U3648 (N_3648,N_2361,N_258);
or U3649 (N_3649,N_2130,N_2639);
and U3650 (N_3650,N_1601,N_1353);
nor U3651 (N_3651,N_212,N_1217);
or U3652 (N_3652,N_2562,N_611);
nand U3653 (N_3653,N_26,N_1524);
nor U3654 (N_3654,N_437,N_674);
or U3655 (N_3655,N_2589,N_131);
xnor U3656 (N_3656,N_777,N_2633);
nor U3657 (N_3657,N_314,N_1742);
and U3658 (N_3658,N_407,N_695);
or U3659 (N_3659,N_2313,N_1349);
nand U3660 (N_3660,N_2953,N_1340);
nor U3661 (N_3661,N_1366,N_1790);
nor U3662 (N_3662,N_957,N_2663);
and U3663 (N_3663,N_2035,N_164);
nor U3664 (N_3664,N_2240,N_1717);
or U3665 (N_3665,N_793,N_1025);
or U3666 (N_3666,N_1662,N_1032);
nor U3667 (N_3667,N_383,N_2705);
or U3668 (N_3668,N_380,N_2458);
nand U3669 (N_3669,N_2541,N_2917);
nand U3670 (N_3670,N_2665,N_1561);
or U3671 (N_3671,N_2338,N_2907);
nand U3672 (N_3672,N_2342,N_618);
nor U3673 (N_3673,N_1569,N_578);
and U3674 (N_3674,N_1247,N_2015);
nand U3675 (N_3675,N_838,N_2548);
and U3676 (N_3676,N_548,N_1737);
nand U3677 (N_3677,N_1377,N_1208);
or U3678 (N_3678,N_160,N_2856);
and U3679 (N_3679,N_2899,N_1437);
and U3680 (N_3680,N_1820,N_391);
and U3681 (N_3681,N_2112,N_2818);
or U3682 (N_3682,N_2148,N_2337);
nand U3683 (N_3683,N_2799,N_2218);
xor U3684 (N_3684,N_724,N_208);
or U3685 (N_3685,N_2658,N_2520);
and U3686 (N_3686,N_263,N_2108);
or U3687 (N_3687,N_1466,N_1905);
nand U3688 (N_3688,N_2101,N_722);
and U3689 (N_3689,N_2628,N_2185);
nand U3690 (N_3690,N_2378,N_575);
nand U3691 (N_3691,N_2834,N_2709);
and U3692 (N_3692,N_1198,N_1881);
nor U3693 (N_3693,N_815,N_2100);
and U3694 (N_3694,N_2254,N_2563);
and U3695 (N_3695,N_2971,N_1244);
or U3696 (N_3696,N_2767,N_891);
and U3697 (N_3697,N_326,N_599);
or U3698 (N_3698,N_2509,N_1797);
nor U3699 (N_3699,N_2839,N_371);
or U3700 (N_3700,N_2213,N_2588);
or U3701 (N_3701,N_2046,N_165);
nor U3702 (N_3702,N_2595,N_1733);
nor U3703 (N_3703,N_2014,N_2960);
or U3704 (N_3704,N_800,N_516);
nor U3705 (N_3705,N_2543,N_2324);
and U3706 (N_3706,N_907,N_2627);
nor U3707 (N_3707,N_619,N_1412);
and U3708 (N_3708,N_865,N_2921);
nor U3709 (N_3709,N_1611,N_242);
nor U3710 (N_3710,N_1256,N_2876);
and U3711 (N_3711,N_1230,N_530);
and U3712 (N_3712,N_450,N_1171);
or U3713 (N_3713,N_2702,N_744);
nand U3714 (N_3714,N_1540,N_1296);
or U3715 (N_3715,N_2087,N_2419);
and U3716 (N_3716,N_2901,N_2727);
or U3717 (N_3717,N_178,N_1099);
or U3718 (N_3718,N_2041,N_2471);
nor U3719 (N_3719,N_2593,N_2202);
and U3720 (N_3720,N_1373,N_666);
nor U3721 (N_3721,N_1472,N_1716);
nor U3722 (N_3722,N_2332,N_2026);
nor U3723 (N_3723,N_2570,N_2965);
nor U3724 (N_3724,N_2862,N_1864);
or U3725 (N_3725,N_2397,N_2973);
nor U3726 (N_3726,N_1248,N_1627);
or U3727 (N_3727,N_1046,N_353);
xnor U3728 (N_3728,N_1137,N_2694);
and U3729 (N_3729,N_106,N_2089);
and U3730 (N_3730,N_333,N_2063);
nand U3731 (N_3731,N_1350,N_694);
and U3732 (N_3732,N_1105,N_1348);
nor U3733 (N_3733,N_2346,N_656);
xnor U3734 (N_3734,N_812,N_1643);
nand U3735 (N_3735,N_1399,N_2258);
xnor U3736 (N_3736,N_1775,N_521);
or U3737 (N_3737,N_2150,N_1983);
nand U3738 (N_3738,N_1553,N_2864);
and U3739 (N_3739,N_1117,N_140);
nand U3740 (N_3740,N_1592,N_1959);
nor U3741 (N_3741,N_1337,N_714);
nor U3742 (N_3742,N_1593,N_962);
nor U3743 (N_3743,N_203,N_615);
nand U3744 (N_3744,N_2559,N_2825);
or U3745 (N_3745,N_2085,N_2070);
nor U3746 (N_3746,N_2111,N_73);
or U3747 (N_3747,N_2493,N_2547);
nor U3748 (N_3748,N_968,N_322);
nand U3749 (N_3749,N_2625,N_518);
and U3750 (N_3750,N_1222,N_1143);
or U3751 (N_3751,N_938,N_987);
nor U3752 (N_3752,N_1305,N_1608);
or U3753 (N_3753,N_677,N_2432);
nand U3754 (N_3754,N_1957,N_1766);
and U3755 (N_3755,N_590,N_650);
and U3756 (N_3756,N_1034,N_404);
nor U3757 (N_3757,N_2146,N_2312);
nor U3758 (N_3758,N_555,N_2011);
and U3759 (N_3759,N_824,N_2788);
nor U3760 (N_3760,N_1448,N_341);
and U3761 (N_3761,N_2525,N_2758);
and U3762 (N_3762,N_2545,N_2572);
and U3763 (N_3763,N_2180,N_2232);
or U3764 (N_3764,N_1671,N_447);
and U3765 (N_3765,N_2671,N_1679);
nand U3766 (N_3766,N_1628,N_2404);
nand U3767 (N_3767,N_150,N_1868);
nand U3768 (N_3768,N_697,N_2287);
nand U3769 (N_3769,N_12,N_1147);
or U3770 (N_3770,N_1513,N_868);
nand U3771 (N_3771,N_614,N_752);
or U3772 (N_3772,N_1674,N_377);
nor U3773 (N_3773,N_2018,N_602);
and U3774 (N_3774,N_2659,N_2918);
nand U3775 (N_3775,N_1129,N_1522);
or U3776 (N_3776,N_2080,N_3);
nor U3777 (N_3777,N_2181,N_2446);
nor U3778 (N_3778,N_476,N_1482);
nor U3779 (N_3779,N_79,N_1808);
nand U3780 (N_3780,N_1022,N_265);
nor U3781 (N_3781,N_1791,N_2427);
nand U3782 (N_3782,N_257,N_1474);
nor U3783 (N_3783,N_1922,N_654);
and U3784 (N_3784,N_181,N_2832);
nand U3785 (N_3785,N_1660,N_1852);
nand U3786 (N_3786,N_107,N_1008);
nand U3787 (N_3787,N_976,N_2500);
or U3788 (N_3788,N_801,N_1498);
or U3789 (N_3789,N_2214,N_88);
nor U3790 (N_3790,N_423,N_2840);
nor U3791 (N_3791,N_1370,N_579);
and U3792 (N_3792,N_2645,N_2291);
and U3793 (N_3793,N_2526,N_773);
nor U3794 (N_3794,N_1746,N_975);
or U3795 (N_3795,N_2131,N_1928);
or U3796 (N_3796,N_301,N_385);
or U3797 (N_3797,N_2034,N_663);
and U3798 (N_3798,N_2807,N_2004);
and U3799 (N_3799,N_2859,N_82);
or U3800 (N_3800,N_1664,N_576);
nor U3801 (N_3801,N_1083,N_200);
or U3802 (N_3802,N_1764,N_2736);
nand U3803 (N_3803,N_2464,N_556);
nor U3804 (N_3804,N_1347,N_2847);
or U3805 (N_3805,N_2406,N_2096);
and U3806 (N_3806,N_2231,N_843);
and U3807 (N_3807,N_512,N_703);
and U3808 (N_3808,N_324,N_98);
nor U3809 (N_3809,N_2442,N_2837);
nand U3810 (N_3810,N_655,N_685);
nand U3811 (N_3811,N_1745,N_1282);
or U3812 (N_3812,N_2863,N_848);
xnor U3813 (N_3813,N_1821,N_1615);
or U3814 (N_3814,N_468,N_1809);
or U3815 (N_3815,N_1578,N_1368);
or U3816 (N_3816,N_2396,N_342);
or U3817 (N_3817,N_376,N_1065);
nand U3818 (N_3818,N_289,N_1955);
nand U3819 (N_3819,N_856,N_2083);
or U3820 (N_3820,N_1415,N_225);
or U3821 (N_3821,N_2650,N_1505);
or U3822 (N_3822,N_2954,N_1093);
or U3823 (N_3823,N_1939,N_274);
or U3824 (N_3824,N_2235,N_1159);
nand U3825 (N_3825,N_1744,N_133);
or U3826 (N_3826,N_367,N_1290);
and U3827 (N_3827,N_2564,N_348);
nand U3828 (N_3828,N_2032,N_725);
and U3829 (N_3829,N_1595,N_194);
nand U3830 (N_3830,N_2027,N_1822);
nor U3831 (N_3831,N_132,N_1568);
and U3832 (N_3832,N_1527,N_788);
and U3833 (N_3833,N_917,N_977);
or U3834 (N_3834,N_688,N_1471);
nor U3835 (N_3835,N_2257,N_185);
nand U3836 (N_3836,N_2348,N_2793);
or U3837 (N_3837,N_2970,N_2990);
nand U3838 (N_3838,N_1195,N_2747);
nand U3839 (N_3839,N_118,N_2114);
nor U3840 (N_3840,N_589,N_1440);
and U3841 (N_3841,N_1421,N_2521);
nor U3842 (N_3842,N_1277,N_2445);
xnor U3843 (N_3843,N_2274,N_1753);
xnor U3844 (N_3844,N_331,N_1824);
or U3845 (N_3845,N_2941,N_941);
xor U3846 (N_3846,N_1449,N_1740);
and U3847 (N_3847,N_1213,N_2765);
and U3848 (N_3848,N_551,N_2998);
nor U3849 (N_3849,N_2529,N_681);
nand U3850 (N_3850,N_855,N_1826);
or U3851 (N_3851,N_1780,N_117);
nand U3852 (N_3852,N_421,N_1109);
nand U3853 (N_3853,N_485,N_1961);
nand U3854 (N_3854,N_741,N_1734);
or U3855 (N_3855,N_1243,N_36);
or U3856 (N_3856,N_1115,N_629);
nand U3857 (N_3857,N_1623,N_388);
nor U3858 (N_3858,N_558,N_2798);
nor U3859 (N_3859,N_465,N_61);
nor U3860 (N_3860,N_1819,N_1445);
nor U3861 (N_3861,N_1566,N_1082);
or U3862 (N_3862,N_1341,N_1144);
or U3863 (N_3863,N_2162,N_2946);
nand U3864 (N_3864,N_2932,N_2268);
and U3865 (N_3865,N_1700,N_2909);
or U3866 (N_3866,N_2764,N_2999);
or U3867 (N_3867,N_2516,N_408);
nor U3868 (N_3868,N_2976,N_1154);
and U3869 (N_3869,N_825,N_1641);
or U3870 (N_3870,N_2701,N_453);
nand U3871 (N_3871,N_584,N_417);
and U3872 (N_3872,N_1614,N_1654);
or U3873 (N_3873,N_1417,N_2402);
nor U3874 (N_3874,N_1418,N_1698);
or U3875 (N_3875,N_1969,N_187);
nor U3876 (N_3876,N_852,N_2199);
or U3877 (N_3877,N_2276,N_1872);
and U3878 (N_3878,N_30,N_1803);
nor U3879 (N_3879,N_2055,N_482);
or U3880 (N_3880,N_2695,N_2684);
or U3881 (N_3881,N_1865,N_649);
or U3882 (N_3882,N_1495,N_1763);
and U3883 (N_3883,N_182,N_693);
nand U3884 (N_3884,N_1029,N_1946);
nand U3885 (N_3885,N_2773,N_625);
nand U3886 (N_3886,N_520,N_1588);
nor U3887 (N_3887,N_2407,N_2838);
nor U3888 (N_3888,N_330,N_2805);
or U3889 (N_3889,N_2882,N_524);
nor U3890 (N_3890,N_1600,N_2207);
and U3891 (N_3891,N_22,N_956);
nor U3892 (N_3892,N_1834,N_953);
and U3893 (N_3893,N_509,N_1422);
nor U3894 (N_3894,N_1447,N_1136);
nor U3895 (N_3895,N_2210,N_2613);
or U3896 (N_3896,N_288,N_660);
and U3897 (N_3897,N_2870,N_1153);
nor U3898 (N_3898,N_943,N_2183);
and U3899 (N_3899,N_2672,N_1923);
nor U3900 (N_3900,N_570,N_457);
nor U3901 (N_3901,N_832,N_2398);
nand U3902 (N_3902,N_2867,N_2206);
or U3903 (N_3903,N_2226,N_428);
nor U3904 (N_3904,N_2980,N_1242);
or U3905 (N_3905,N_1427,N_1949);
nand U3906 (N_3906,N_1503,N_2373);
nand U3907 (N_3907,N_2077,N_2194);
and U3908 (N_3908,N_154,N_1333);
and U3909 (N_3909,N_2016,N_818);
nand U3910 (N_3910,N_789,N_829);
nor U3911 (N_3911,N_83,N_2480);
or U3912 (N_3912,N_1921,N_1459);
or U3913 (N_3913,N_811,N_100);
nand U3914 (N_3914,N_1696,N_1711);
or U3915 (N_3915,N_1539,N_1604);
and U3916 (N_3916,N_2607,N_2649);
nor U3917 (N_3917,N_2643,N_940);
or U3918 (N_3918,N_2030,N_1441);
nand U3919 (N_3919,N_290,N_601);
nor U3920 (N_3920,N_1164,N_1536);
and U3921 (N_3921,N_1968,N_1715);
and U3922 (N_3922,N_980,N_2594);
nor U3923 (N_3923,N_1617,N_1552);
nor U3924 (N_3924,N_1712,N_1625);
or U3925 (N_3925,N_361,N_2994);
nor U3926 (N_3926,N_998,N_2714);
or U3927 (N_3927,N_1062,N_2872);
nor U3928 (N_3928,N_2142,N_564);
and U3929 (N_3929,N_2912,N_2227);
or U3930 (N_3930,N_2455,N_2537);
and U3931 (N_3931,N_2188,N_844);
and U3932 (N_3932,N_2487,N_2317);
and U3933 (N_3933,N_1846,N_808);
and U3934 (N_3934,N_1461,N_2086);
and U3935 (N_3935,N_93,N_2372);
and U3936 (N_3936,N_1618,N_1686);
or U3937 (N_3937,N_1833,N_1324);
nand U3938 (N_3938,N_519,N_2597);
nand U3939 (N_3939,N_1829,N_59);
nor U3940 (N_3940,N_1397,N_1887);
nand U3941 (N_3941,N_218,N_2356);
or U3942 (N_3942,N_2908,N_170);
and U3943 (N_3943,N_1793,N_770);
nor U3944 (N_3944,N_1911,N_900);
and U3945 (N_3945,N_739,N_2722);
nor U3946 (N_3946,N_180,N_104);
nand U3947 (N_3947,N_1250,N_464);
and U3948 (N_3948,N_2778,N_2802);
or U3949 (N_3949,N_372,N_151);
or U3950 (N_3950,N_1346,N_1430);
and U3951 (N_3951,N_2984,N_247);
and U3952 (N_3952,N_1576,N_2752);
nor U3953 (N_3953,N_1799,N_2224);
or U3954 (N_3954,N_1372,N_65);
nor U3955 (N_3955,N_2712,N_2642);
and U3956 (N_3956,N_906,N_538);
or U3957 (N_3957,N_1443,N_2884);
nor U3958 (N_3958,N_2986,N_2887);
nand U3959 (N_3959,N_507,N_2676);
nor U3960 (N_3960,N_1264,N_1855);
or U3961 (N_3961,N_1331,N_2848);
and U3962 (N_3962,N_448,N_1475);
and U3963 (N_3963,N_2272,N_2430);
and U3964 (N_3964,N_2916,N_2647);
or U3965 (N_3965,N_1239,N_2457);
or U3966 (N_3966,N_94,N_885);
nand U3967 (N_3967,N_2061,N_21);
or U3968 (N_3968,N_2399,N_1094);
and U3969 (N_3969,N_1483,N_1529);
and U3970 (N_3970,N_2382,N_2833);
nor U3971 (N_3971,N_2914,N_2081);
and U3972 (N_3972,N_113,N_1413);
and U3973 (N_3973,N_2315,N_2544);
nor U3974 (N_3974,N_513,N_951);
nor U3975 (N_3975,N_350,N_797);
nand U3976 (N_3976,N_436,N_996);
nor U3977 (N_3977,N_1436,N_610);
and U3978 (N_3978,N_1987,N_233);
nand U3979 (N_3979,N_2902,N_2808);
nand U3980 (N_3980,N_533,N_2964);
nand U3981 (N_3981,N_2186,N_96);
and U3982 (N_3982,N_1086,N_1096);
nand U3983 (N_3983,N_2677,N_220);
or U3984 (N_3984,N_1877,N_2037);
nand U3985 (N_3985,N_365,N_1460);
and U3986 (N_3986,N_2201,N_701);
or U3987 (N_3987,N_1581,N_1365);
xnor U3988 (N_3988,N_964,N_321);
nor U3989 (N_3989,N_2687,N_2245);
nand U3990 (N_3990,N_628,N_1585);
nor U3991 (N_3991,N_707,N_934);
nor U3992 (N_3992,N_2454,N_1594);
and U3993 (N_3993,N_2889,N_1782);
nor U3994 (N_3994,N_2288,N_729);
nand U3995 (N_3995,N_2234,N_1730);
nor U3996 (N_3996,N_737,N_1038);
nor U3997 (N_3997,N_1125,N_1707);
nand U3998 (N_3998,N_2732,N_458);
nand U3999 (N_3999,N_2777,N_1383);
or U4000 (N_4000,N_1786,N_671);
nor U4001 (N_4001,N_2810,N_308);
nand U4002 (N_4002,N_989,N_2160);
or U4003 (N_4003,N_1995,N_175);
or U4004 (N_4004,N_2307,N_2524);
or U4005 (N_4005,N_207,N_2182);
nor U4006 (N_4006,N_1757,N_488);
and U4007 (N_4007,N_1873,N_1506);
and U4008 (N_4008,N_240,N_2144);
xnor U4009 (N_4009,N_32,N_620);
nand U4010 (N_4010,N_2707,N_2812);
nand U4011 (N_4011,N_2134,N_1335);
or U4012 (N_4012,N_1683,N_547);
nor U4013 (N_4013,N_471,N_2716);
or U4014 (N_4014,N_1028,N_2680);
and U4015 (N_4015,N_2269,N_60);
or U4016 (N_4016,N_1613,N_25);
or U4017 (N_4017,N_2044,N_1840);
or U4018 (N_4018,N_1060,N_2222);
nand U4019 (N_4019,N_2557,N_2966);
nor U4020 (N_4020,N_209,N_2674);
and U4021 (N_4021,N_1970,N_115);
and U4022 (N_4022,N_2900,N_2826);
or U4023 (N_4023,N_2706,N_2568);
nor U4024 (N_4024,N_2829,N_1680);
nor U4025 (N_4025,N_2415,N_2565);
nor U4026 (N_4026,N_1473,N_630);
nor U4027 (N_4027,N_2621,N_2439);
nor U4028 (N_4028,N_2341,N_2256);
or U4029 (N_4029,N_2670,N_277);
and U4030 (N_4030,N_1312,N_2605);
or U4031 (N_4031,N_1344,N_1978);
or U4032 (N_4032,N_2903,N_2119);
nand U4033 (N_4033,N_2583,N_1785);
nor U4034 (N_4034,N_1091,N_2459);
or U4035 (N_4035,N_109,N_806);
and U4036 (N_4036,N_1988,N_648);
or U4037 (N_4037,N_1017,N_384);
nand U4038 (N_4038,N_2539,N_2710);
nor U4039 (N_4039,N_1783,N_239);
nand U4040 (N_4040,N_1446,N_1064);
or U4041 (N_4041,N_1270,N_2309);
or U4042 (N_4042,N_1738,N_1526);
nor U4043 (N_4043,N_631,N_2059);
nor U4044 (N_4044,N_1551,N_1535);
nand U4045 (N_4045,N_197,N_2211);
nand U4046 (N_4046,N_1236,N_2711);
nor U4047 (N_4047,N_2498,N_2474);
nor U4048 (N_4048,N_2165,N_2698);
or U4049 (N_4049,N_2813,N_2968);
and U4050 (N_4050,N_2715,N_1550);
xnor U4051 (N_4051,N_2319,N_2152);
and U4052 (N_4052,N_1079,N_1828);
and U4053 (N_4053,N_2005,N_735);
or U4054 (N_4054,N_193,N_1304);
nand U4055 (N_4055,N_438,N_1356);
and U4056 (N_4056,N_2553,N_2737);
and U4057 (N_4057,N_346,N_830);
and U4058 (N_4058,N_1409,N_2811);
nand U4059 (N_4059,N_456,N_364);
and U4060 (N_4060,N_2173,N_2614);
nand U4061 (N_4061,N_1320,N_937);
and U4062 (N_4062,N_475,N_188);
nand U4063 (N_4063,N_1135,N_2790);
nor U4064 (N_4064,N_970,N_1603);
or U4065 (N_4065,N_1488,N_1210);
or U4066 (N_4066,N_1179,N_1054);
nor U4067 (N_4067,N_1245,N_1009);
and U4068 (N_4068,N_2806,N_1701);
and U4069 (N_4069,N_110,N_2299);
nand U4070 (N_4070,N_2776,N_2109);
and U4071 (N_4071,N_2043,N_1932);
nand U4072 (N_4072,N_1560,N_587);
or U4073 (N_4073,N_1945,N_2421);
and U4074 (N_4074,N_1036,N_933);
nor U4075 (N_4075,N_2740,N_1856);
and U4076 (N_4076,N_2575,N_2009);
or U4077 (N_4077,N_1682,N_1599);
and U4078 (N_4078,N_1188,N_2745);
or U4079 (N_4079,N_2447,N_1114);
nor U4080 (N_4080,N_238,N_1943);
nand U4081 (N_4081,N_2956,N_1020);
nand U4082 (N_4082,N_2074,N_1294);
nand U4083 (N_4083,N_405,N_2225);
or U4084 (N_4084,N_74,N_2636);
and U4085 (N_4085,N_2846,N_1933);
and U4086 (N_4086,N_2686,N_529);
or U4087 (N_4087,N_2426,N_318);
or U4088 (N_4088,N_2873,N_2759);
and U4089 (N_4089,N_511,N_2305);
or U4090 (N_4090,N_1924,N_2989);
and U4091 (N_4091,N_1233,N_2467);
and U4092 (N_4092,N_2322,N_349);
nand U4093 (N_4093,N_2090,N_2380);
and U4094 (N_4094,N_2796,N_1155);
and U4095 (N_4095,N_1359,N_2724);
and U4096 (N_4096,N_1607,N_2552);
or U4097 (N_4097,N_932,N_745);
nand U4098 (N_4098,N_2540,N_2482);
nand U4099 (N_4099,N_28,N_2988);
nor U4100 (N_4100,N_774,N_1398);
and U4101 (N_4101,N_2362,N_2470);
nand U4102 (N_4102,N_2757,N_1110);
nand U4103 (N_4103,N_1263,N_605);
nand U4104 (N_4104,N_291,N_1586);
nand U4105 (N_4105,N_2394,N_1005);
and U4106 (N_4106,N_1869,N_1758);
nor U4107 (N_4107,N_983,N_416);
and U4108 (N_4108,N_68,N_396);
and U4109 (N_4109,N_406,N_2804);
nand U4110 (N_4110,N_1597,N_275);
and U4111 (N_4111,N_2113,N_936);
and U4112 (N_4112,N_1697,N_1063);
nor U4113 (N_4113,N_1893,N_696);
nor U4114 (N_4114,N_80,N_2066);
nor U4115 (N_4115,N_1309,N_1596);
and U4116 (N_4116,N_76,N_1544);
nand U4117 (N_4117,N_1583,N_2756);
and U4118 (N_4118,N_542,N_1161);
and U4119 (N_4119,N_2697,N_952);
or U4120 (N_4120,N_841,N_1832);
or U4121 (N_4121,N_2506,N_2518);
and U4122 (N_4122,N_2555,N_2121);
or U4123 (N_4123,N_2668,N_717);
nand U4124 (N_4124,N_211,N_2271);
or U4125 (N_4125,N_569,N_2656);
nor U4126 (N_4126,N_1177,N_1823);
or U4127 (N_4127,N_2508,N_2343);
or U4128 (N_4128,N_954,N_882);
nand U4129 (N_4129,N_1396,N_817);
nor U4130 (N_4130,N_922,N_2098);
or U4131 (N_4131,N_2166,N_847);
nand U4132 (N_4132,N_1067,N_1937);
nor U4133 (N_4133,N_403,N_2922);
nor U4134 (N_4134,N_2875,N_184);
and U4135 (N_4135,N_1364,N_2996);
nand U4136 (N_4136,N_820,N_1917);
or U4137 (N_4137,N_1487,N_609);
and U4138 (N_4138,N_1172,N_2997);
or U4139 (N_4139,N_2982,N_411);
and U4140 (N_4140,N_1325,N_2389);
nand U4141 (N_4141,N_2072,N_1888);
nand U4142 (N_4142,N_684,N_2507);
nor U4143 (N_4143,N_1101,N_2930);
nor U4144 (N_4144,N_1760,N_2969);
or U4145 (N_4145,N_1655,N_2486);
nor U4146 (N_4146,N_928,N_171);
or U4147 (N_4147,N_1286,N_1493);
and U4148 (N_4148,N_1723,N_1902);
nor U4149 (N_4149,N_972,N_2263);
or U4150 (N_4150,N_1973,N_1139);
xor U4151 (N_4151,N_158,N_2815);
nor U4152 (N_4152,N_2273,N_2400);
or U4153 (N_4153,N_64,N_1543);
nor U4154 (N_4154,N_1439,N_2156);
or U4155 (N_4155,N_2892,N_340);
or U4156 (N_4156,N_2596,N_2340);
nor U4157 (N_4157,N_1719,N_1358);
nor U4158 (N_4158,N_2387,N_2135);
nand U4159 (N_4159,N_990,N_2880);
nor U4160 (N_4160,N_2920,N_721);
or U4161 (N_4161,N_924,N_202);
or U4162 (N_4162,N_794,N_2768);
and U4163 (N_4163,N_2534,N_1141);
nor U4164 (N_4164,N_539,N_1706);
and U4165 (N_4165,N_370,N_84);
or U4166 (N_4166,N_1842,N_1019);
and U4167 (N_4167,N_1077,N_1962);
and U4168 (N_4168,N_595,N_2311);
nand U4169 (N_4169,N_2438,N_1116);
xnor U4170 (N_4170,N_1788,N_183);
nor U4171 (N_4171,N_394,N_2766);
and U4172 (N_4172,N_545,N_2693);
nand U4173 (N_4173,N_2187,N_1419);
or U4174 (N_4174,N_7,N_544);
and U4175 (N_4175,N_1464,N_2316);
nand U4176 (N_4176,N_2267,N_690);
or U4177 (N_4177,N_2328,N_1343);
nand U4178 (N_4178,N_1148,N_2751);
and U4179 (N_4179,N_2761,N_1407);
nand U4180 (N_4180,N_191,N_1133);
and U4181 (N_4181,N_1215,N_1642);
or U4182 (N_4182,N_1124,N_1515);
nand U4183 (N_4183,N_2496,N_2228);
nor U4184 (N_4184,N_315,N_286);
nand U4185 (N_4185,N_352,N_2463);
nor U4186 (N_4186,N_2008,N_414);
or U4187 (N_4187,N_360,N_502);
nand U4188 (N_4188,N_2503,N_2129);
nand U4189 (N_4189,N_223,N_2204);
or U4190 (N_4190,N_2158,N_362);
nand U4191 (N_4191,N_588,N_2991);
nand U4192 (N_4192,N_1678,N_2265);
nor U4193 (N_4193,N_1481,N_911);
and U4194 (N_4194,N_1859,N_176);
or U4195 (N_4195,N_2145,N_1619);
nand U4196 (N_4196,N_1035,N_2139);
or U4197 (N_4197,N_2048,N_356);
or U4198 (N_4198,N_919,N_1854);
and U4199 (N_4199,N_866,N_2590);
or U4200 (N_4200,N_312,N_42);
nor U4201 (N_4201,N_2844,N_646);
or U4202 (N_4202,N_432,N_894);
or U4203 (N_4203,N_553,N_141);
and U4204 (N_4204,N_70,N_1175);
nor U4205 (N_4205,N_1435,N_1411);
and U4206 (N_4206,N_2646,N_1151);
or U4207 (N_4207,N_2321,N_2401);
or U4208 (N_4208,N_1477,N_2003);
nor U4209 (N_4209,N_1132,N_126);
xor U4210 (N_4210,N_1880,N_1126);
nor U4211 (N_4211,N_429,N_1927);
or U4212 (N_4212,N_267,N_1841);
nand U4213 (N_4213,N_2769,N_37);
nor U4214 (N_4214,N_809,N_711);
nand U4215 (N_4215,N_1375,N_1140);
or U4216 (N_4216,N_607,N_2979);
nor U4217 (N_4217,N_667,N_2289);
or U4218 (N_4218,N_1688,N_554);
or U4219 (N_4219,N_2703,N_2772);
nor U4220 (N_4220,N_2170,N_1178);
nand U4221 (N_4221,N_260,N_1691);
or U4222 (N_4222,N_764,N_254);
or U4223 (N_4223,N_1265,N_536);
and U4224 (N_4224,N_955,N_446);
or U4225 (N_4225,N_676,N_1321);
and U4226 (N_4226,N_2664,N_2106);
or U4227 (N_4227,N_1111,N_2489);
nor U4228 (N_4228,N_2855,N_1194);
or U4229 (N_4229,N_1122,N_2251);
and U4230 (N_4230,N_1624,N_144);
nand U4231 (N_4231,N_2002,N_2374);
and U4232 (N_4232,N_2869,N_1573);
or U4233 (N_4233,N_1967,N_1097);
or U4234 (N_4234,N_283,N_413);
or U4235 (N_4235,N_337,N_2868);
nand U4236 (N_4236,N_1993,N_111);
nor U4237 (N_4237,N_2823,N_2549);
nor U4238 (N_4238,N_467,N_1113);
or U4239 (N_4239,N_549,N_2951);
nor U4240 (N_4240,N_461,N_1467);
or U4241 (N_4241,N_2292,N_1223);
or U4242 (N_4242,N_1689,N_525);
nor U4243 (N_4243,N_1858,N_1533);
and U4244 (N_4244,N_1789,N_1805);
or U4245 (N_4245,N_638,N_591);
xor U4246 (N_4246,N_2891,N_1018);
or U4247 (N_4247,N_2786,N_393);
or U4248 (N_4248,N_1919,N_2352);
and U4249 (N_4249,N_2076,N_2386);
and U4250 (N_4250,N_498,N_2771);
and U4251 (N_4251,N_1357,N_759);
nand U4252 (N_4252,N_1104,N_33);
and U4253 (N_4253,N_1800,N_1444);
nor U4254 (N_4254,N_2678,N_1704);
and U4255 (N_4255,N_505,N_1408);
or U4256 (N_4256,N_1541,N_143);
or U4257 (N_4257,N_2068,N_95);
or U4258 (N_4258,N_2481,N_2574);
nand U4259 (N_4259,N_2007,N_1332);
nor U4260 (N_4260,N_2558,N_2591);
and U4261 (N_4261,N_1632,N_2140);
or U4262 (N_4262,N_1616,N_213);
and U4263 (N_4263,N_1016,N_244);
nand U4264 (N_4264,N_58,N_2550);
nor U4265 (N_4265,N_2661,N_1134);
or U4266 (N_4266,N_1999,N_2443);
nand U4267 (N_4267,N_1702,N_958);
nand U4268 (N_4268,N_1571,N_1721);
nor U4269 (N_4269,N_2945,N_2075);
nand U4270 (N_4270,N_895,N_29);
or U4271 (N_4271,N_156,N_2924);
or U4272 (N_4272,N_2462,N_1886);
nand U4273 (N_4273,N_2505,N_1792);
nand U4274 (N_4274,N_1693,N_2857);
nor U4275 (N_4275,N_1520,N_1297);
nand U4276 (N_4276,N_804,N_490);
and U4277 (N_4277,N_234,N_2476);
nand U4278 (N_4278,N_1517,N_2913);
and U4279 (N_4279,N_1163,N_327);
and U4280 (N_4280,N_395,N_293);
nand U4281 (N_4281,N_2318,N_2931);
or U4282 (N_4282,N_379,N_2082);
nand U4283 (N_4283,N_2738,N_2893);
and U4284 (N_4284,N_2013,N_452);
or U4285 (N_4285,N_2816,N_1253);
and U4286 (N_4286,N_462,N_125);
nor U4287 (N_4287,N_1532,N_1168);
nand U4288 (N_4288,N_1000,N_1041);
nand U4289 (N_4289,N_2236,N_2329);
and U4290 (N_4290,N_1925,N_47);
nand U4291 (N_4291,N_1197,N_2630);
and U4292 (N_4292,N_2750,N_1291);
or U4293 (N_4293,N_2784,N_608);
xnor U4294 (N_4294,N_568,N_2571);
or U4295 (N_4295,N_1205,N_2451);
and U4296 (N_4296,N_1092,N_1787);
nand U4297 (N_4297,N_604,N_2683);
nor U4298 (N_4298,N_2115,N_99);
nand U4299 (N_4299,N_2632,N_2538);
or U4300 (N_4300,N_583,N_2154);
nor U4301 (N_4301,N_2429,N_2860);
nand U4302 (N_4302,N_643,N_2);
or U4303 (N_4303,N_874,N_985);
and U4304 (N_4304,N_771,N_1211);
or U4305 (N_4305,N_2431,N_2618);
or U4306 (N_4306,N_1299,N_1798);
nor U4307 (N_4307,N_2293,N_986);
nor U4308 (N_4308,N_2409,N_1804);
nor U4309 (N_4309,N_261,N_2344);
and U4310 (N_4310,N_2587,N_1229);
or U4311 (N_4311,N_2952,N_828);
nor U4312 (N_4312,N_466,N_1980);
and U4313 (N_4313,N_2688,N_1289);
nand U4314 (N_4314,N_1056,N_2164);
nand U4315 (N_4315,N_56,N_295);
nor U4316 (N_4316,N_1251,N_710);
nor U4317 (N_4317,N_2216,N_1903);
nand U4318 (N_4318,N_1499,N_2620);
and U4319 (N_4319,N_81,N_2795);
and U4320 (N_4320,N_1130,N_1777);
nand U4321 (N_4321,N_1001,N_347);
and U4322 (N_4322,N_351,N_38);
nand U4323 (N_4323,N_329,N_702);
and U4324 (N_4324,N_1405,N_430);
or U4325 (N_4325,N_814,N_2079);
nor U4326 (N_4326,N_1971,N_776);
and U4327 (N_4327,N_2281,N_1650);
nand U4328 (N_4328,N_2820,N_2822);
and U4329 (N_4329,N_1885,N_635);
or U4330 (N_4330,N_2910,N_1275);
or U4331 (N_4331,N_1724,N_1199);
and U4332 (N_4332,N_1061,N_965);
nor U4333 (N_4333,N_1940,N_1180);
nand U4334 (N_4334,N_1572,N_1867);
or U4335 (N_4335,N_1752,N_45);
nand U4336 (N_4336,N_1313,N_2655);
and U4337 (N_4337,N_2038,N_2717);
nor U4338 (N_4338,N_1910,N_292);
and U4339 (N_4339,N_2334,N_1876);
nand U4340 (N_4340,N_1450,N_2383);
or U4341 (N_4341,N_1070,N_960);
or U4342 (N_4342,N_2302,N_2915);
and U4343 (N_4343,N_2099,N_1174);
and U4344 (N_4344,N_1084,N_387);
or U4345 (N_4345,N_1579,N_686);
nor U4346 (N_4346,N_217,N_2241);
nand U4347 (N_4347,N_2617,N_929);
or U4348 (N_4348,N_2436,N_401);
nand U4349 (N_4349,N_890,N_2662);
nand U4350 (N_4350,N_799,N_1559);
and U4351 (N_4351,N_1367,N_2713);
or U4352 (N_4352,N_2435,N_219);
nand U4353 (N_4353,N_2723,N_1784);
nor U4354 (N_4354,N_230,N_592);
nor U4355 (N_4355,N_2465,N_580);
and U4356 (N_4356,N_831,N_596);
nor U4357 (N_4357,N_127,N_270);
or U4358 (N_4358,N_2515,N_31);
nor U4359 (N_4359,N_731,N_228);
nor U4360 (N_4360,N_1825,N_1895);
and U4361 (N_4361,N_2290,N_1508);
nand U4362 (N_4362,N_2542,N_2905);
and U4363 (N_4363,N_2367,N_2163);
nand U4364 (N_4364,N_967,N_237);
or U4365 (N_4365,N_1765,N_577);
nor U4366 (N_4366,N_1850,N_262);
nor U4367 (N_4367,N_867,N_1930);
nand U4368 (N_4368,N_1901,N_2775);
nand U4369 (N_4369,N_1530,N_1431);
nand U4370 (N_4370,N_1646,N_2093);
and U4371 (N_4371,N_1098,N_1434);
and U4372 (N_4372,N_2577,N_2260);
nand U4373 (N_4373,N_1479,N_2809);
nand U4374 (N_4374,N_1649,N_2392);
or U4375 (N_4375,N_1612,N_161);
and U4376 (N_4376,N_1232,N_2782);
or U4377 (N_4377,N_168,N_2959);
or U4378 (N_4378,N_1470,N_477);
nand U4379 (N_4379,N_294,N_903);
or U4380 (N_4380,N_1220,N_822);
and U4381 (N_4381,N_1323,N_897);
and U4382 (N_4382,N_1476,N_993);
or U4383 (N_4383,N_946,N_2940);
and U4384 (N_4384,N_1390,N_1634);
or U4385 (N_4385,N_2359,N_374);
and U4386 (N_4386,N_363,N_433);
or U4387 (N_4387,N_1221,N_1851);
and U4388 (N_4388,N_683,N_2310);
or U4389 (N_4389,N_1908,N_2411);
or U4390 (N_4390,N_1606,N_1379);
nor U4391 (N_4391,N_199,N_1123);
or U4392 (N_4392,N_307,N_2935);
nand U4393 (N_4393,N_1555,N_1112);
or U4394 (N_4394,N_901,N_767);
nor U4395 (N_4395,N_2801,N_763);
or U4396 (N_4396,N_1629,N_2203);
nor U4397 (N_4397,N_255,N_2602);
nor U4398 (N_4398,N_1827,N_69);
nand U4399 (N_4399,N_146,N_1381);
or U4400 (N_4400,N_55,N_1004);
nand U4401 (N_4401,N_2412,N_1186);
nor U4402 (N_4402,N_328,N_1735);
nor U4403 (N_4403,N_1644,N_128);
nor U4404 (N_4404,N_904,N_201);
or U4405 (N_4405,N_755,N_2742);
or U4406 (N_4406,N_375,N_287);
nor U4407 (N_4407,N_1059,N_1710);
nor U4408 (N_4408,N_899,N_1037);
nand U4409 (N_4409,N_214,N_39);
or U4410 (N_4410,N_2936,N_888);
nand U4411 (N_4411,N_2229,N_1699);
nand U4412 (N_4412,N_1465,N_758);
nor U4413 (N_4413,N_2028,N_2219);
nor U4414 (N_4414,N_859,N_1813);
nand U4415 (N_4415,N_359,N_2215);
nand U4416 (N_4416,N_2874,N_16);
or U4417 (N_4417,N_600,N_335);
nor U4418 (N_4418,N_1043,N_1638);
nor U4419 (N_4419,N_2023,N_1235);
and U4420 (N_4420,N_1267,N_995);
and U4421 (N_4421,N_984,N_2300);
xnor U4422 (N_4422,N_139,N_1645);
and U4423 (N_4423,N_2600,N_2739);
nor U4424 (N_4424,N_765,N_572);
nor U4425 (N_4425,N_1580,N_1831);
xnor U4426 (N_4426,N_1027,N_2393);
nand U4427 (N_4427,N_272,N_479);
and U4428 (N_4428,N_1285,N_2314);
nor U4429 (N_4429,N_1081,N_991);
and U4430 (N_4430,N_159,N_2000);
or U4431 (N_4431,N_1631,N_2176);
and U4432 (N_4432,N_1469,N_1212);
nor U4433 (N_4433,N_1322,N_2523);
or U4434 (N_4434,N_2349,N_827);
and U4435 (N_4435,N_682,N_2449);
or U4436 (N_4436,N_1705,N_2502);
and U4437 (N_4437,N_1166,N_2992);
nor U4438 (N_4438,N_2551,N_2040);
and U4439 (N_4439,N_1977,N_27);
nor U4440 (N_4440,N_2169,N_2102);
nor U4441 (N_4441,N_20,N_1293);
or U4442 (N_4442,N_2733,N_210);
nor U4443 (N_4443,N_2220,N_120);
nor U4444 (N_4444,N_6,N_2501);
nand U4445 (N_4445,N_1203,N_1261);
nand U4446 (N_4446,N_2045,N_1736);
or U4447 (N_4447,N_1871,N_1863);
nand U4448 (N_4448,N_2626,N_2690);
nand U4449 (N_4449,N_732,N_1209);
nand U4450 (N_4450,N_2453,N_2019);
or U4451 (N_4451,N_1747,N_1769);
or U4452 (N_4452,N_2420,N_1078);
and U4453 (N_4453,N_1781,N_1853);
and U4454 (N_4454,N_1189,N_2853);
and U4455 (N_4455,N_528,N_713);
and U4456 (N_4456,N_914,N_1456);
and U4457 (N_4457,N_2350,N_2012);
nor U4458 (N_4458,N_412,N_46);
nor U4459 (N_4459,N_1252,N_52);
or U4460 (N_4460,N_2366,N_1875);
nand U4461 (N_4461,N_691,N_560);
nor U4462 (N_4462,N_1156,N_1288);
or U4463 (N_4463,N_2592,N_278);
and U4464 (N_4464,N_273,N_1192);
or U4465 (N_4465,N_1255,N_320);
or U4466 (N_4466,N_574,N_1754);
nor U4467 (N_4467,N_1015,N_2456);
nor U4468 (N_4468,N_1085,N_390);
and U4469 (N_4469,N_2787,N_1574);
nor U4470 (N_4470,N_719,N_459);
and U4471 (N_4471,N_473,N_2363);
nor U4472 (N_4472,N_2223,N_1031);
nor U4473 (N_4473,N_1692,N_1663);
nor U4474 (N_4474,N_2774,N_1315);
or U4475 (N_4475,N_483,N_1622);
nand U4476 (N_4476,N_1394,N_2168);
xnor U4477 (N_4477,N_1351,N_2126);
and U4478 (N_4478,N_1668,N_24);
and U4479 (N_4479,N_1274,N_982);
or U4480 (N_4480,N_1392,N_2249);
nor U4481 (N_4481,N_1272,N_2978);
nor U4482 (N_4482,N_803,N_679);
nor U4483 (N_4483,N_1401,N_2556);
nand U4484 (N_4484,N_130,N_2744);
and U4485 (N_4485,N_2780,N_2071);
and U4486 (N_4486,N_2460,N_51);
xnor U4487 (N_4487,N_2580,N_2049);
or U4488 (N_4488,N_1318,N_445);
nand U4489 (N_4489,N_1306,N_915);
nor U4490 (N_4490,N_766,N_1989);
nand U4491 (N_4491,N_939,N_1049);
nand U4492 (N_4492,N_1021,N_2339);
nor U4493 (N_4493,N_1100,N_2280);
or U4494 (N_4494,N_734,N_1676);
and U4495 (N_4495,N_72,N_1839);
or U4496 (N_4496,N_616,N_942);
or U4497 (N_4497,N_1167,N_13);
nand U4498 (N_4498,N_1425,N_1531);
or U4499 (N_4499,N_2247,N_1273);
and U4500 (N_4500,N_959,N_1092);
nand U4501 (N_4501,N_993,N_311);
nand U4502 (N_4502,N_1166,N_2754);
nor U4503 (N_4503,N_1202,N_119);
nand U4504 (N_4504,N_2106,N_406);
nor U4505 (N_4505,N_71,N_1572);
or U4506 (N_4506,N_390,N_1827);
and U4507 (N_4507,N_1221,N_2415);
nand U4508 (N_4508,N_421,N_1031);
or U4509 (N_4509,N_2469,N_971);
nand U4510 (N_4510,N_1295,N_987);
or U4511 (N_4511,N_35,N_1994);
or U4512 (N_4512,N_1766,N_1158);
nand U4513 (N_4513,N_2899,N_1522);
or U4514 (N_4514,N_2638,N_1718);
nand U4515 (N_4515,N_2351,N_353);
or U4516 (N_4516,N_1751,N_451);
or U4517 (N_4517,N_1865,N_1529);
nand U4518 (N_4518,N_2254,N_46);
nor U4519 (N_4519,N_2746,N_1606);
and U4520 (N_4520,N_2157,N_2952);
nand U4521 (N_4521,N_2758,N_2947);
nor U4522 (N_4522,N_1367,N_2589);
and U4523 (N_4523,N_2015,N_2239);
and U4524 (N_4524,N_31,N_923);
nor U4525 (N_4525,N_1407,N_142);
or U4526 (N_4526,N_1143,N_1444);
and U4527 (N_4527,N_2316,N_1521);
nor U4528 (N_4528,N_1098,N_747);
nand U4529 (N_4529,N_2270,N_2149);
xor U4530 (N_4530,N_944,N_1460);
nand U4531 (N_4531,N_2059,N_1559);
or U4532 (N_4532,N_2205,N_2611);
and U4533 (N_4533,N_990,N_1902);
xnor U4534 (N_4534,N_1287,N_2023);
nor U4535 (N_4535,N_266,N_759);
and U4536 (N_4536,N_1497,N_2636);
nand U4537 (N_4537,N_1569,N_2272);
and U4538 (N_4538,N_2514,N_1498);
or U4539 (N_4539,N_2025,N_1988);
and U4540 (N_4540,N_1491,N_2543);
nand U4541 (N_4541,N_2396,N_2882);
nor U4542 (N_4542,N_1873,N_1716);
nand U4543 (N_4543,N_78,N_1578);
and U4544 (N_4544,N_2580,N_2066);
and U4545 (N_4545,N_1005,N_2705);
and U4546 (N_4546,N_701,N_2625);
and U4547 (N_4547,N_2729,N_1750);
or U4548 (N_4548,N_1259,N_1816);
or U4549 (N_4549,N_239,N_1447);
and U4550 (N_4550,N_2653,N_1341);
and U4551 (N_4551,N_355,N_824);
or U4552 (N_4552,N_2047,N_1282);
nor U4553 (N_4553,N_1482,N_2431);
or U4554 (N_4554,N_2141,N_450);
nand U4555 (N_4555,N_1378,N_849);
nand U4556 (N_4556,N_2477,N_639);
or U4557 (N_4557,N_259,N_2735);
and U4558 (N_4558,N_753,N_647);
nor U4559 (N_4559,N_1654,N_295);
nor U4560 (N_4560,N_1379,N_1483);
nor U4561 (N_4561,N_2150,N_796);
or U4562 (N_4562,N_236,N_1936);
or U4563 (N_4563,N_2136,N_436);
nand U4564 (N_4564,N_1569,N_1990);
nand U4565 (N_4565,N_2862,N_436);
and U4566 (N_4566,N_2411,N_2356);
nor U4567 (N_4567,N_2511,N_379);
nor U4568 (N_4568,N_2081,N_167);
xor U4569 (N_4569,N_2903,N_1055);
nand U4570 (N_4570,N_462,N_1449);
or U4571 (N_4571,N_119,N_358);
and U4572 (N_4572,N_1638,N_1961);
nand U4573 (N_4573,N_776,N_704);
and U4574 (N_4574,N_211,N_2525);
and U4575 (N_4575,N_1841,N_482);
nand U4576 (N_4576,N_65,N_1945);
and U4577 (N_4577,N_349,N_579);
and U4578 (N_4578,N_31,N_1770);
and U4579 (N_4579,N_1510,N_2132);
and U4580 (N_4580,N_2285,N_839);
nor U4581 (N_4581,N_1145,N_641);
and U4582 (N_4582,N_2518,N_2453);
nor U4583 (N_4583,N_2778,N_1898);
nor U4584 (N_4584,N_2866,N_1127);
nor U4585 (N_4585,N_462,N_209);
or U4586 (N_4586,N_2298,N_282);
nand U4587 (N_4587,N_1156,N_65);
or U4588 (N_4588,N_1831,N_2007);
and U4589 (N_4589,N_2473,N_2859);
or U4590 (N_4590,N_586,N_696);
nor U4591 (N_4591,N_1340,N_917);
nor U4592 (N_4592,N_2361,N_2567);
and U4593 (N_4593,N_121,N_77);
or U4594 (N_4594,N_2926,N_1413);
or U4595 (N_4595,N_1150,N_838);
or U4596 (N_4596,N_1180,N_538);
nand U4597 (N_4597,N_2021,N_942);
nand U4598 (N_4598,N_1644,N_998);
and U4599 (N_4599,N_1696,N_681);
or U4600 (N_4600,N_1798,N_27);
nand U4601 (N_4601,N_173,N_122);
nor U4602 (N_4602,N_80,N_455);
nand U4603 (N_4603,N_279,N_2149);
nand U4604 (N_4604,N_2960,N_1387);
nor U4605 (N_4605,N_2348,N_206);
nor U4606 (N_4606,N_1202,N_2070);
and U4607 (N_4607,N_2324,N_1739);
nor U4608 (N_4608,N_1007,N_175);
nand U4609 (N_4609,N_911,N_2361);
or U4610 (N_4610,N_763,N_2907);
nor U4611 (N_4611,N_2407,N_1318);
and U4612 (N_4612,N_2036,N_1406);
and U4613 (N_4613,N_2609,N_1586);
nand U4614 (N_4614,N_2964,N_252);
nor U4615 (N_4615,N_1840,N_749);
and U4616 (N_4616,N_1591,N_1566);
and U4617 (N_4617,N_2634,N_1178);
and U4618 (N_4618,N_2874,N_1512);
nor U4619 (N_4619,N_2530,N_1582);
or U4620 (N_4620,N_2064,N_655);
and U4621 (N_4621,N_2903,N_552);
nand U4622 (N_4622,N_2346,N_246);
and U4623 (N_4623,N_356,N_2862);
nand U4624 (N_4624,N_535,N_558);
or U4625 (N_4625,N_42,N_750);
or U4626 (N_4626,N_2838,N_338);
nor U4627 (N_4627,N_2373,N_1052);
or U4628 (N_4628,N_2921,N_1062);
nor U4629 (N_4629,N_903,N_881);
nor U4630 (N_4630,N_771,N_2181);
nand U4631 (N_4631,N_497,N_2420);
nor U4632 (N_4632,N_156,N_55);
or U4633 (N_4633,N_1396,N_1400);
and U4634 (N_4634,N_1250,N_2051);
or U4635 (N_4635,N_2859,N_1157);
or U4636 (N_4636,N_2025,N_870);
nor U4637 (N_4637,N_2849,N_1492);
or U4638 (N_4638,N_2022,N_2292);
nor U4639 (N_4639,N_2597,N_984);
nor U4640 (N_4640,N_1212,N_1889);
or U4641 (N_4641,N_2197,N_2022);
and U4642 (N_4642,N_535,N_256);
nand U4643 (N_4643,N_1580,N_1686);
nand U4644 (N_4644,N_1727,N_619);
nand U4645 (N_4645,N_1457,N_2855);
nor U4646 (N_4646,N_393,N_220);
nand U4647 (N_4647,N_1921,N_238);
or U4648 (N_4648,N_1549,N_2507);
nor U4649 (N_4649,N_1074,N_267);
nand U4650 (N_4650,N_2452,N_1937);
nand U4651 (N_4651,N_1816,N_2908);
or U4652 (N_4652,N_2686,N_1834);
or U4653 (N_4653,N_1915,N_1005);
nand U4654 (N_4654,N_1073,N_2862);
nand U4655 (N_4655,N_2051,N_856);
nand U4656 (N_4656,N_2240,N_1850);
or U4657 (N_4657,N_1003,N_1612);
or U4658 (N_4658,N_797,N_1764);
nand U4659 (N_4659,N_2154,N_722);
nand U4660 (N_4660,N_2957,N_20);
nor U4661 (N_4661,N_774,N_2194);
nor U4662 (N_4662,N_1580,N_2466);
nor U4663 (N_4663,N_434,N_1870);
or U4664 (N_4664,N_432,N_1649);
xor U4665 (N_4665,N_1625,N_579);
and U4666 (N_4666,N_1908,N_1791);
nand U4667 (N_4667,N_317,N_2561);
and U4668 (N_4668,N_505,N_2790);
nand U4669 (N_4669,N_2041,N_47);
and U4670 (N_4670,N_35,N_1699);
xnor U4671 (N_4671,N_2697,N_172);
nor U4672 (N_4672,N_2465,N_1499);
and U4673 (N_4673,N_1840,N_2160);
nand U4674 (N_4674,N_2856,N_326);
nor U4675 (N_4675,N_1587,N_120);
nor U4676 (N_4676,N_2999,N_2052);
xnor U4677 (N_4677,N_220,N_965);
and U4678 (N_4678,N_2707,N_287);
or U4679 (N_4679,N_1579,N_2298);
and U4680 (N_4680,N_2693,N_1502);
nand U4681 (N_4681,N_683,N_1031);
or U4682 (N_4682,N_1370,N_1976);
and U4683 (N_4683,N_269,N_2041);
and U4684 (N_4684,N_2098,N_825);
and U4685 (N_4685,N_1129,N_2453);
nand U4686 (N_4686,N_1846,N_406);
nand U4687 (N_4687,N_1199,N_2992);
nor U4688 (N_4688,N_13,N_2169);
and U4689 (N_4689,N_1891,N_738);
and U4690 (N_4690,N_1279,N_2983);
and U4691 (N_4691,N_2536,N_600);
or U4692 (N_4692,N_251,N_1968);
and U4693 (N_4693,N_1354,N_2919);
or U4694 (N_4694,N_1999,N_1738);
nand U4695 (N_4695,N_1772,N_145);
nand U4696 (N_4696,N_2787,N_307);
nand U4697 (N_4697,N_1740,N_607);
and U4698 (N_4698,N_910,N_2593);
nor U4699 (N_4699,N_557,N_1776);
nand U4700 (N_4700,N_2900,N_2093);
or U4701 (N_4701,N_2056,N_1390);
nand U4702 (N_4702,N_2926,N_21);
or U4703 (N_4703,N_1705,N_365);
or U4704 (N_4704,N_2566,N_1825);
nand U4705 (N_4705,N_2210,N_617);
xnor U4706 (N_4706,N_1572,N_1456);
nor U4707 (N_4707,N_1890,N_1281);
nor U4708 (N_4708,N_10,N_1999);
and U4709 (N_4709,N_2338,N_1924);
nand U4710 (N_4710,N_1679,N_1359);
and U4711 (N_4711,N_1869,N_398);
and U4712 (N_4712,N_1938,N_2105);
nor U4713 (N_4713,N_2014,N_1992);
xor U4714 (N_4714,N_731,N_1631);
nand U4715 (N_4715,N_1125,N_83);
nand U4716 (N_4716,N_2572,N_1906);
nor U4717 (N_4717,N_54,N_2459);
nand U4718 (N_4718,N_614,N_527);
nor U4719 (N_4719,N_710,N_2785);
and U4720 (N_4720,N_1509,N_395);
nand U4721 (N_4721,N_2217,N_2902);
nor U4722 (N_4722,N_2393,N_1490);
nand U4723 (N_4723,N_744,N_285);
nor U4724 (N_4724,N_975,N_1347);
nand U4725 (N_4725,N_2886,N_714);
nor U4726 (N_4726,N_192,N_1191);
and U4727 (N_4727,N_1047,N_2388);
and U4728 (N_4728,N_484,N_280);
and U4729 (N_4729,N_229,N_1792);
or U4730 (N_4730,N_746,N_772);
nand U4731 (N_4731,N_591,N_1254);
or U4732 (N_4732,N_1727,N_2646);
nor U4733 (N_4733,N_1098,N_1555);
and U4734 (N_4734,N_2551,N_2363);
nand U4735 (N_4735,N_2661,N_2404);
nand U4736 (N_4736,N_2043,N_835);
nand U4737 (N_4737,N_452,N_1951);
nand U4738 (N_4738,N_2444,N_2243);
nand U4739 (N_4739,N_1001,N_1091);
nor U4740 (N_4740,N_2358,N_2487);
nor U4741 (N_4741,N_1058,N_2647);
nand U4742 (N_4742,N_2993,N_1078);
or U4743 (N_4743,N_1229,N_690);
nand U4744 (N_4744,N_1607,N_194);
nand U4745 (N_4745,N_2239,N_2061);
or U4746 (N_4746,N_2098,N_2534);
and U4747 (N_4747,N_1813,N_25);
or U4748 (N_4748,N_1535,N_2246);
nand U4749 (N_4749,N_2391,N_179);
and U4750 (N_4750,N_1144,N_2775);
or U4751 (N_4751,N_887,N_2944);
and U4752 (N_4752,N_33,N_1668);
nand U4753 (N_4753,N_606,N_2975);
nand U4754 (N_4754,N_2947,N_189);
and U4755 (N_4755,N_1664,N_2902);
nor U4756 (N_4756,N_330,N_688);
or U4757 (N_4757,N_560,N_1080);
nor U4758 (N_4758,N_1209,N_1700);
and U4759 (N_4759,N_380,N_762);
or U4760 (N_4760,N_629,N_1090);
nand U4761 (N_4761,N_1276,N_972);
nor U4762 (N_4762,N_2688,N_2948);
and U4763 (N_4763,N_2952,N_916);
nor U4764 (N_4764,N_266,N_588);
and U4765 (N_4765,N_677,N_2223);
nor U4766 (N_4766,N_192,N_2179);
nor U4767 (N_4767,N_718,N_2676);
nand U4768 (N_4768,N_125,N_1710);
and U4769 (N_4769,N_1104,N_2972);
and U4770 (N_4770,N_782,N_1889);
nor U4771 (N_4771,N_737,N_417);
nor U4772 (N_4772,N_1077,N_685);
nand U4773 (N_4773,N_2445,N_2060);
and U4774 (N_4774,N_2161,N_1322);
nand U4775 (N_4775,N_2576,N_1815);
xor U4776 (N_4776,N_2865,N_1543);
and U4777 (N_4777,N_2019,N_975);
and U4778 (N_4778,N_2283,N_1032);
and U4779 (N_4779,N_2461,N_850);
and U4780 (N_4780,N_1729,N_2855);
nor U4781 (N_4781,N_1451,N_1984);
and U4782 (N_4782,N_2502,N_333);
and U4783 (N_4783,N_2329,N_2915);
nor U4784 (N_4784,N_543,N_2012);
or U4785 (N_4785,N_2971,N_1941);
or U4786 (N_4786,N_874,N_66);
nor U4787 (N_4787,N_1271,N_1562);
nor U4788 (N_4788,N_2777,N_944);
nor U4789 (N_4789,N_1321,N_1941);
nand U4790 (N_4790,N_1027,N_77);
nor U4791 (N_4791,N_2308,N_1253);
nor U4792 (N_4792,N_2367,N_1076);
nand U4793 (N_4793,N_2583,N_1751);
nand U4794 (N_4794,N_2211,N_2025);
and U4795 (N_4795,N_2756,N_608);
nor U4796 (N_4796,N_2477,N_1132);
nand U4797 (N_4797,N_1780,N_1490);
and U4798 (N_4798,N_2672,N_2944);
and U4799 (N_4799,N_1194,N_1930);
and U4800 (N_4800,N_2868,N_675);
or U4801 (N_4801,N_133,N_2438);
or U4802 (N_4802,N_2038,N_2680);
and U4803 (N_4803,N_2049,N_1701);
xnor U4804 (N_4804,N_2939,N_1544);
nand U4805 (N_4805,N_441,N_2649);
nand U4806 (N_4806,N_2095,N_1884);
and U4807 (N_4807,N_1163,N_1677);
nor U4808 (N_4808,N_1968,N_1872);
or U4809 (N_4809,N_2442,N_2127);
and U4810 (N_4810,N_2289,N_1068);
nand U4811 (N_4811,N_1965,N_2113);
nand U4812 (N_4812,N_1016,N_408);
nand U4813 (N_4813,N_124,N_747);
or U4814 (N_4814,N_143,N_1548);
or U4815 (N_4815,N_1566,N_414);
and U4816 (N_4816,N_495,N_2542);
and U4817 (N_4817,N_1089,N_2475);
and U4818 (N_4818,N_2173,N_971);
nand U4819 (N_4819,N_2026,N_2633);
nor U4820 (N_4820,N_730,N_1174);
and U4821 (N_4821,N_646,N_1931);
and U4822 (N_4822,N_1529,N_1537);
or U4823 (N_4823,N_1915,N_96);
or U4824 (N_4824,N_281,N_2815);
and U4825 (N_4825,N_171,N_2577);
nand U4826 (N_4826,N_1127,N_2863);
nand U4827 (N_4827,N_1699,N_1618);
and U4828 (N_4828,N_1610,N_2112);
nand U4829 (N_4829,N_272,N_1527);
and U4830 (N_4830,N_914,N_186);
and U4831 (N_4831,N_935,N_409);
nor U4832 (N_4832,N_217,N_2650);
nand U4833 (N_4833,N_1211,N_1640);
xnor U4834 (N_4834,N_1130,N_2104);
nand U4835 (N_4835,N_118,N_1978);
or U4836 (N_4836,N_2343,N_945);
nand U4837 (N_4837,N_164,N_2703);
and U4838 (N_4838,N_1355,N_1168);
and U4839 (N_4839,N_484,N_1327);
and U4840 (N_4840,N_1351,N_2125);
or U4841 (N_4841,N_1486,N_508);
nor U4842 (N_4842,N_2615,N_1910);
or U4843 (N_4843,N_1320,N_790);
nand U4844 (N_4844,N_261,N_62);
or U4845 (N_4845,N_788,N_845);
nand U4846 (N_4846,N_1131,N_1332);
nand U4847 (N_4847,N_1051,N_1454);
nor U4848 (N_4848,N_2513,N_1883);
and U4849 (N_4849,N_2986,N_2204);
or U4850 (N_4850,N_1488,N_490);
and U4851 (N_4851,N_573,N_1157);
xor U4852 (N_4852,N_1963,N_1398);
nor U4853 (N_4853,N_844,N_1699);
and U4854 (N_4854,N_1327,N_2773);
nand U4855 (N_4855,N_1928,N_2557);
xnor U4856 (N_4856,N_2755,N_977);
nand U4857 (N_4857,N_924,N_2874);
and U4858 (N_4858,N_1057,N_376);
or U4859 (N_4859,N_300,N_401);
and U4860 (N_4860,N_2862,N_692);
nand U4861 (N_4861,N_2652,N_899);
nor U4862 (N_4862,N_1198,N_1640);
or U4863 (N_4863,N_1580,N_768);
nand U4864 (N_4864,N_2583,N_708);
and U4865 (N_4865,N_752,N_1930);
nand U4866 (N_4866,N_1847,N_2784);
nand U4867 (N_4867,N_1435,N_2696);
nand U4868 (N_4868,N_2759,N_273);
and U4869 (N_4869,N_2962,N_37);
and U4870 (N_4870,N_2260,N_1169);
nor U4871 (N_4871,N_1919,N_445);
or U4872 (N_4872,N_2264,N_227);
and U4873 (N_4873,N_211,N_138);
nor U4874 (N_4874,N_2272,N_2818);
and U4875 (N_4875,N_2065,N_1432);
nand U4876 (N_4876,N_2902,N_1133);
and U4877 (N_4877,N_2606,N_1170);
nand U4878 (N_4878,N_2687,N_1522);
or U4879 (N_4879,N_64,N_1499);
nor U4880 (N_4880,N_1660,N_2497);
or U4881 (N_4881,N_372,N_1118);
and U4882 (N_4882,N_2515,N_2336);
nand U4883 (N_4883,N_2169,N_1156);
and U4884 (N_4884,N_2654,N_1368);
and U4885 (N_4885,N_1702,N_2700);
nor U4886 (N_4886,N_996,N_1060);
or U4887 (N_4887,N_589,N_2553);
and U4888 (N_4888,N_1465,N_1002);
nor U4889 (N_4889,N_946,N_1868);
and U4890 (N_4890,N_676,N_1249);
nor U4891 (N_4891,N_676,N_1664);
nor U4892 (N_4892,N_2303,N_1508);
nand U4893 (N_4893,N_1899,N_2986);
nor U4894 (N_4894,N_1205,N_2511);
nand U4895 (N_4895,N_120,N_996);
or U4896 (N_4896,N_231,N_703);
xor U4897 (N_4897,N_2557,N_881);
nor U4898 (N_4898,N_696,N_2574);
nand U4899 (N_4899,N_227,N_2806);
nor U4900 (N_4900,N_1303,N_1213);
nor U4901 (N_4901,N_66,N_1150);
or U4902 (N_4902,N_753,N_1356);
nand U4903 (N_4903,N_2076,N_2083);
or U4904 (N_4904,N_2494,N_762);
or U4905 (N_4905,N_380,N_1516);
nand U4906 (N_4906,N_1828,N_2428);
and U4907 (N_4907,N_1124,N_1833);
nor U4908 (N_4908,N_84,N_361);
or U4909 (N_4909,N_2524,N_2246);
and U4910 (N_4910,N_2261,N_2066);
xnor U4911 (N_4911,N_435,N_2547);
and U4912 (N_4912,N_2644,N_1427);
nand U4913 (N_4913,N_2135,N_2416);
nand U4914 (N_4914,N_167,N_1298);
nor U4915 (N_4915,N_1612,N_1122);
and U4916 (N_4916,N_145,N_241);
and U4917 (N_4917,N_656,N_691);
or U4918 (N_4918,N_600,N_1800);
nor U4919 (N_4919,N_1998,N_1316);
and U4920 (N_4920,N_1635,N_211);
nand U4921 (N_4921,N_337,N_537);
and U4922 (N_4922,N_342,N_356);
and U4923 (N_4923,N_2264,N_1129);
nor U4924 (N_4924,N_623,N_2469);
and U4925 (N_4925,N_1023,N_1844);
nor U4926 (N_4926,N_1844,N_1119);
nor U4927 (N_4927,N_407,N_1438);
nor U4928 (N_4928,N_1393,N_2833);
nand U4929 (N_4929,N_1362,N_1662);
nor U4930 (N_4930,N_2410,N_1328);
nor U4931 (N_4931,N_1244,N_421);
and U4932 (N_4932,N_2182,N_2063);
or U4933 (N_4933,N_693,N_870);
nor U4934 (N_4934,N_1232,N_2191);
nor U4935 (N_4935,N_1558,N_399);
or U4936 (N_4936,N_1989,N_427);
nand U4937 (N_4937,N_2397,N_259);
nand U4938 (N_4938,N_1008,N_2276);
and U4939 (N_4939,N_683,N_2014);
or U4940 (N_4940,N_1129,N_479);
and U4941 (N_4941,N_31,N_1447);
nand U4942 (N_4942,N_2206,N_1859);
or U4943 (N_4943,N_2742,N_2971);
nor U4944 (N_4944,N_117,N_152);
and U4945 (N_4945,N_758,N_121);
nor U4946 (N_4946,N_97,N_2931);
or U4947 (N_4947,N_1419,N_946);
and U4948 (N_4948,N_808,N_425);
or U4949 (N_4949,N_2465,N_528);
nor U4950 (N_4950,N_2355,N_1189);
nor U4951 (N_4951,N_216,N_2575);
nand U4952 (N_4952,N_2186,N_2720);
or U4953 (N_4953,N_361,N_553);
nor U4954 (N_4954,N_1299,N_641);
and U4955 (N_4955,N_2176,N_2537);
nor U4956 (N_4956,N_921,N_2423);
nand U4957 (N_4957,N_375,N_396);
nor U4958 (N_4958,N_1531,N_2941);
nand U4959 (N_4959,N_1925,N_1177);
nor U4960 (N_4960,N_1204,N_1829);
nor U4961 (N_4961,N_808,N_446);
or U4962 (N_4962,N_1073,N_852);
nor U4963 (N_4963,N_1382,N_2906);
and U4964 (N_4964,N_112,N_1080);
nor U4965 (N_4965,N_2410,N_2744);
nand U4966 (N_4966,N_2255,N_2424);
and U4967 (N_4967,N_1862,N_2647);
and U4968 (N_4968,N_2583,N_2745);
or U4969 (N_4969,N_923,N_2561);
and U4970 (N_4970,N_1066,N_151);
or U4971 (N_4971,N_424,N_1241);
nor U4972 (N_4972,N_2529,N_1243);
nand U4973 (N_4973,N_2028,N_2316);
nand U4974 (N_4974,N_1726,N_1971);
or U4975 (N_4975,N_1268,N_370);
and U4976 (N_4976,N_253,N_2481);
and U4977 (N_4977,N_2471,N_1778);
nor U4978 (N_4978,N_1225,N_1040);
nand U4979 (N_4979,N_514,N_1579);
or U4980 (N_4980,N_2944,N_1387);
nand U4981 (N_4981,N_39,N_2927);
nor U4982 (N_4982,N_1364,N_100);
nand U4983 (N_4983,N_2831,N_493);
or U4984 (N_4984,N_413,N_2728);
or U4985 (N_4985,N_1658,N_449);
nor U4986 (N_4986,N_1542,N_2836);
and U4987 (N_4987,N_2646,N_585);
nand U4988 (N_4988,N_67,N_1232);
nand U4989 (N_4989,N_1503,N_2490);
nand U4990 (N_4990,N_2970,N_1107);
nor U4991 (N_4991,N_2398,N_1066);
nand U4992 (N_4992,N_2801,N_2970);
and U4993 (N_4993,N_2200,N_1263);
nand U4994 (N_4994,N_2909,N_902);
or U4995 (N_4995,N_1908,N_1474);
or U4996 (N_4996,N_2580,N_1674);
nor U4997 (N_4997,N_1370,N_454);
nand U4998 (N_4998,N_986,N_357);
nor U4999 (N_4999,N_426,N_355);
nand U5000 (N_5000,N_2457,N_2592);
nor U5001 (N_5001,N_735,N_647);
and U5002 (N_5002,N_38,N_828);
and U5003 (N_5003,N_2198,N_2429);
nor U5004 (N_5004,N_1233,N_1637);
or U5005 (N_5005,N_331,N_1676);
nand U5006 (N_5006,N_1822,N_707);
nor U5007 (N_5007,N_1687,N_757);
nand U5008 (N_5008,N_2720,N_2058);
and U5009 (N_5009,N_2123,N_2809);
nor U5010 (N_5010,N_1951,N_2396);
or U5011 (N_5011,N_204,N_897);
or U5012 (N_5012,N_1927,N_2293);
or U5013 (N_5013,N_122,N_2918);
nor U5014 (N_5014,N_1013,N_2901);
nand U5015 (N_5015,N_861,N_765);
xnor U5016 (N_5016,N_272,N_849);
and U5017 (N_5017,N_1648,N_1310);
nand U5018 (N_5018,N_2459,N_1275);
nand U5019 (N_5019,N_2302,N_1747);
and U5020 (N_5020,N_1504,N_1260);
or U5021 (N_5021,N_2007,N_158);
nand U5022 (N_5022,N_2182,N_1626);
or U5023 (N_5023,N_1274,N_219);
or U5024 (N_5024,N_2818,N_2957);
nor U5025 (N_5025,N_531,N_2390);
and U5026 (N_5026,N_1509,N_1672);
or U5027 (N_5027,N_2110,N_2134);
nor U5028 (N_5028,N_764,N_2307);
nand U5029 (N_5029,N_711,N_2482);
nand U5030 (N_5030,N_57,N_1950);
nand U5031 (N_5031,N_1790,N_2955);
or U5032 (N_5032,N_1724,N_2179);
and U5033 (N_5033,N_2586,N_2106);
and U5034 (N_5034,N_2891,N_1576);
or U5035 (N_5035,N_2934,N_522);
nand U5036 (N_5036,N_774,N_1347);
nand U5037 (N_5037,N_2130,N_1010);
or U5038 (N_5038,N_2352,N_2715);
or U5039 (N_5039,N_876,N_2047);
and U5040 (N_5040,N_2014,N_2936);
or U5041 (N_5041,N_722,N_1986);
nor U5042 (N_5042,N_2636,N_2352);
nand U5043 (N_5043,N_1012,N_2472);
and U5044 (N_5044,N_2201,N_2574);
or U5045 (N_5045,N_774,N_2707);
nand U5046 (N_5046,N_892,N_2270);
nor U5047 (N_5047,N_1353,N_1713);
and U5048 (N_5048,N_2067,N_2884);
xor U5049 (N_5049,N_2098,N_787);
and U5050 (N_5050,N_1962,N_327);
and U5051 (N_5051,N_1306,N_1353);
and U5052 (N_5052,N_1505,N_1513);
and U5053 (N_5053,N_409,N_1696);
and U5054 (N_5054,N_2701,N_1969);
nand U5055 (N_5055,N_2160,N_750);
nor U5056 (N_5056,N_537,N_1932);
or U5057 (N_5057,N_2743,N_348);
and U5058 (N_5058,N_2573,N_376);
or U5059 (N_5059,N_2303,N_2666);
nand U5060 (N_5060,N_1197,N_2301);
nand U5061 (N_5061,N_2756,N_2016);
nor U5062 (N_5062,N_974,N_419);
nand U5063 (N_5063,N_1146,N_2641);
nand U5064 (N_5064,N_2666,N_2375);
nor U5065 (N_5065,N_2170,N_1216);
nor U5066 (N_5066,N_287,N_2493);
or U5067 (N_5067,N_2504,N_1447);
nand U5068 (N_5068,N_1456,N_1083);
xnor U5069 (N_5069,N_1608,N_554);
or U5070 (N_5070,N_355,N_1377);
nor U5071 (N_5071,N_2016,N_1801);
and U5072 (N_5072,N_1829,N_914);
nand U5073 (N_5073,N_1301,N_1298);
and U5074 (N_5074,N_960,N_2521);
or U5075 (N_5075,N_2731,N_618);
nand U5076 (N_5076,N_2331,N_2993);
nand U5077 (N_5077,N_1748,N_2833);
nor U5078 (N_5078,N_657,N_1819);
nand U5079 (N_5079,N_910,N_1847);
nand U5080 (N_5080,N_859,N_544);
nand U5081 (N_5081,N_19,N_2548);
nor U5082 (N_5082,N_2155,N_2030);
nor U5083 (N_5083,N_1362,N_631);
and U5084 (N_5084,N_312,N_728);
and U5085 (N_5085,N_1359,N_722);
or U5086 (N_5086,N_1284,N_1263);
nand U5087 (N_5087,N_1735,N_2637);
nor U5088 (N_5088,N_2667,N_919);
and U5089 (N_5089,N_2681,N_1998);
and U5090 (N_5090,N_2930,N_2726);
and U5091 (N_5091,N_113,N_2767);
nand U5092 (N_5092,N_531,N_936);
nand U5093 (N_5093,N_2092,N_1428);
or U5094 (N_5094,N_192,N_510);
nor U5095 (N_5095,N_2794,N_2103);
nor U5096 (N_5096,N_865,N_398);
or U5097 (N_5097,N_1893,N_1831);
and U5098 (N_5098,N_477,N_2745);
nor U5099 (N_5099,N_1411,N_2302);
nand U5100 (N_5100,N_1857,N_2521);
nand U5101 (N_5101,N_1248,N_2564);
or U5102 (N_5102,N_2204,N_637);
nor U5103 (N_5103,N_1854,N_2472);
nor U5104 (N_5104,N_1523,N_153);
or U5105 (N_5105,N_2875,N_1143);
or U5106 (N_5106,N_980,N_2723);
nand U5107 (N_5107,N_1401,N_2422);
nand U5108 (N_5108,N_394,N_734);
nand U5109 (N_5109,N_2846,N_2594);
nor U5110 (N_5110,N_2431,N_1809);
nand U5111 (N_5111,N_2508,N_954);
nor U5112 (N_5112,N_628,N_885);
or U5113 (N_5113,N_2753,N_2414);
and U5114 (N_5114,N_1555,N_787);
nand U5115 (N_5115,N_2498,N_721);
nor U5116 (N_5116,N_426,N_2916);
nand U5117 (N_5117,N_2810,N_2812);
or U5118 (N_5118,N_2099,N_1215);
and U5119 (N_5119,N_1027,N_7);
and U5120 (N_5120,N_1567,N_1848);
nor U5121 (N_5121,N_713,N_1127);
and U5122 (N_5122,N_2124,N_189);
nor U5123 (N_5123,N_598,N_2770);
nand U5124 (N_5124,N_687,N_1886);
and U5125 (N_5125,N_204,N_2896);
or U5126 (N_5126,N_2628,N_909);
or U5127 (N_5127,N_2100,N_507);
nand U5128 (N_5128,N_627,N_2484);
and U5129 (N_5129,N_2361,N_1741);
or U5130 (N_5130,N_468,N_2999);
or U5131 (N_5131,N_2459,N_2552);
nand U5132 (N_5132,N_1486,N_1019);
nand U5133 (N_5133,N_241,N_1414);
nor U5134 (N_5134,N_1707,N_2421);
and U5135 (N_5135,N_484,N_2375);
nor U5136 (N_5136,N_2094,N_1781);
nor U5137 (N_5137,N_174,N_1487);
nor U5138 (N_5138,N_1406,N_785);
or U5139 (N_5139,N_2717,N_577);
or U5140 (N_5140,N_1258,N_2585);
nor U5141 (N_5141,N_1127,N_2293);
nor U5142 (N_5142,N_2765,N_1335);
or U5143 (N_5143,N_1044,N_1845);
nand U5144 (N_5144,N_2196,N_1691);
nor U5145 (N_5145,N_323,N_2353);
and U5146 (N_5146,N_1614,N_2269);
nor U5147 (N_5147,N_60,N_587);
nand U5148 (N_5148,N_464,N_1701);
or U5149 (N_5149,N_1640,N_1681);
or U5150 (N_5150,N_1011,N_2726);
nor U5151 (N_5151,N_1786,N_334);
and U5152 (N_5152,N_2180,N_977);
and U5153 (N_5153,N_1065,N_409);
nand U5154 (N_5154,N_465,N_1328);
and U5155 (N_5155,N_1522,N_2440);
and U5156 (N_5156,N_1591,N_133);
or U5157 (N_5157,N_2097,N_2069);
nand U5158 (N_5158,N_1107,N_2999);
or U5159 (N_5159,N_2340,N_542);
and U5160 (N_5160,N_2390,N_410);
nor U5161 (N_5161,N_2944,N_718);
or U5162 (N_5162,N_1981,N_591);
nand U5163 (N_5163,N_2384,N_1707);
nand U5164 (N_5164,N_2685,N_1088);
nor U5165 (N_5165,N_126,N_2255);
nor U5166 (N_5166,N_703,N_1795);
nand U5167 (N_5167,N_1766,N_2191);
or U5168 (N_5168,N_1249,N_929);
nand U5169 (N_5169,N_2801,N_71);
or U5170 (N_5170,N_2206,N_101);
nand U5171 (N_5171,N_651,N_2911);
and U5172 (N_5172,N_547,N_261);
and U5173 (N_5173,N_2592,N_1630);
or U5174 (N_5174,N_1184,N_1737);
nor U5175 (N_5175,N_735,N_857);
nand U5176 (N_5176,N_2435,N_1893);
nand U5177 (N_5177,N_1007,N_1365);
and U5178 (N_5178,N_892,N_459);
or U5179 (N_5179,N_596,N_674);
or U5180 (N_5180,N_5,N_1136);
or U5181 (N_5181,N_210,N_1363);
or U5182 (N_5182,N_2819,N_659);
and U5183 (N_5183,N_2248,N_1047);
and U5184 (N_5184,N_1479,N_224);
and U5185 (N_5185,N_17,N_1440);
and U5186 (N_5186,N_2682,N_218);
or U5187 (N_5187,N_2890,N_846);
nand U5188 (N_5188,N_2280,N_878);
nor U5189 (N_5189,N_615,N_1737);
nor U5190 (N_5190,N_1217,N_2540);
nand U5191 (N_5191,N_563,N_920);
nor U5192 (N_5192,N_1562,N_2874);
nand U5193 (N_5193,N_70,N_280);
nor U5194 (N_5194,N_1792,N_689);
nand U5195 (N_5195,N_1726,N_1999);
and U5196 (N_5196,N_1161,N_2990);
or U5197 (N_5197,N_1149,N_2540);
nor U5198 (N_5198,N_2584,N_964);
nor U5199 (N_5199,N_1207,N_2308);
nand U5200 (N_5200,N_797,N_46);
and U5201 (N_5201,N_1422,N_2523);
or U5202 (N_5202,N_1201,N_1609);
and U5203 (N_5203,N_2774,N_828);
and U5204 (N_5204,N_2409,N_579);
and U5205 (N_5205,N_1098,N_920);
nand U5206 (N_5206,N_849,N_1377);
nor U5207 (N_5207,N_1437,N_2081);
or U5208 (N_5208,N_1208,N_848);
and U5209 (N_5209,N_754,N_1981);
and U5210 (N_5210,N_1848,N_2975);
and U5211 (N_5211,N_588,N_2095);
nand U5212 (N_5212,N_2083,N_1715);
or U5213 (N_5213,N_2760,N_2352);
xnor U5214 (N_5214,N_134,N_198);
nor U5215 (N_5215,N_1816,N_2541);
or U5216 (N_5216,N_234,N_876);
or U5217 (N_5217,N_657,N_1377);
or U5218 (N_5218,N_266,N_1432);
or U5219 (N_5219,N_2419,N_1973);
or U5220 (N_5220,N_2399,N_2262);
nand U5221 (N_5221,N_1915,N_1894);
and U5222 (N_5222,N_2015,N_2732);
and U5223 (N_5223,N_1625,N_1737);
or U5224 (N_5224,N_1988,N_1133);
and U5225 (N_5225,N_1881,N_519);
nand U5226 (N_5226,N_2477,N_1714);
nor U5227 (N_5227,N_1018,N_1802);
or U5228 (N_5228,N_2156,N_2164);
nand U5229 (N_5229,N_2442,N_2358);
nor U5230 (N_5230,N_419,N_1099);
nor U5231 (N_5231,N_2248,N_1402);
and U5232 (N_5232,N_2457,N_1874);
nand U5233 (N_5233,N_19,N_2159);
and U5234 (N_5234,N_86,N_1998);
nor U5235 (N_5235,N_1988,N_2012);
nor U5236 (N_5236,N_2505,N_2146);
or U5237 (N_5237,N_2592,N_1793);
nand U5238 (N_5238,N_115,N_2003);
and U5239 (N_5239,N_1983,N_814);
or U5240 (N_5240,N_2810,N_2526);
nand U5241 (N_5241,N_2130,N_745);
and U5242 (N_5242,N_389,N_810);
nand U5243 (N_5243,N_809,N_2386);
and U5244 (N_5244,N_236,N_765);
or U5245 (N_5245,N_1043,N_1655);
or U5246 (N_5246,N_2501,N_2211);
nand U5247 (N_5247,N_2915,N_1194);
nor U5248 (N_5248,N_1653,N_1710);
nand U5249 (N_5249,N_1672,N_2511);
nor U5250 (N_5250,N_2140,N_2978);
and U5251 (N_5251,N_342,N_2651);
and U5252 (N_5252,N_1674,N_984);
nor U5253 (N_5253,N_1331,N_451);
or U5254 (N_5254,N_1918,N_1941);
nand U5255 (N_5255,N_161,N_124);
or U5256 (N_5256,N_1983,N_1202);
or U5257 (N_5257,N_1274,N_1397);
or U5258 (N_5258,N_1383,N_1113);
and U5259 (N_5259,N_970,N_272);
nor U5260 (N_5260,N_2273,N_2037);
nor U5261 (N_5261,N_1207,N_1913);
and U5262 (N_5262,N_371,N_1116);
nand U5263 (N_5263,N_2878,N_1994);
nand U5264 (N_5264,N_2759,N_2589);
nand U5265 (N_5265,N_2511,N_1591);
nand U5266 (N_5266,N_1903,N_2874);
xnor U5267 (N_5267,N_1486,N_2212);
or U5268 (N_5268,N_1049,N_1217);
nor U5269 (N_5269,N_1783,N_523);
and U5270 (N_5270,N_1014,N_1738);
and U5271 (N_5271,N_1329,N_2439);
and U5272 (N_5272,N_1010,N_1332);
nand U5273 (N_5273,N_2573,N_1459);
or U5274 (N_5274,N_2555,N_1076);
or U5275 (N_5275,N_1159,N_2795);
nor U5276 (N_5276,N_711,N_274);
nand U5277 (N_5277,N_1181,N_977);
and U5278 (N_5278,N_1032,N_2383);
or U5279 (N_5279,N_2965,N_484);
or U5280 (N_5280,N_2877,N_2499);
or U5281 (N_5281,N_2048,N_2170);
and U5282 (N_5282,N_1014,N_1453);
or U5283 (N_5283,N_1150,N_2094);
nand U5284 (N_5284,N_1886,N_205);
nor U5285 (N_5285,N_346,N_1514);
and U5286 (N_5286,N_2450,N_256);
nand U5287 (N_5287,N_923,N_627);
nand U5288 (N_5288,N_1730,N_798);
nor U5289 (N_5289,N_881,N_1013);
nand U5290 (N_5290,N_1552,N_4);
nor U5291 (N_5291,N_1902,N_215);
and U5292 (N_5292,N_275,N_2738);
nor U5293 (N_5293,N_2588,N_1480);
nor U5294 (N_5294,N_943,N_2375);
nand U5295 (N_5295,N_457,N_1930);
or U5296 (N_5296,N_1145,N_500);
nor U5297 (N_5297,N_2781,N_487);
nor U5298 (N_5298,N_1504,N_1212);
nand U5299 (N_5299,N_2378,N_1200);
or U5300 (N_5300,N_737,N_700);
or U5301 (N_5301,N_910,N_1858);
nor U5302 (N_5302,N_583,N_2280);
nand U5303 (N_5303,N_2891,N_1763);
and U5304 (N_5304,N_2229,N_1202);
nor U5305 (N_5305,N_1524,N_157);
or U5306 (N_5306,N_2389,N_316);
or U5307 (N_5307,N_2241,N_2467);
nand U5308 (N_5308,N_1644,N_2615);
and U5309 (N_5309,N_2798,N_986);
and U5310 (N_5310,N_2024,N_2905);
and U5311 (N_5311,N_1201,N_317);
nand U5312 (N_5312,N_2088,N_1975);
nand U5313 (N_5313,N_438,N_1575);
or U5314 (N_5314,N_2886,N_1009);
or U5315 (N_5315,N_2254,N_494);
nand U5316 (N_5316,N_105,N_939);
or U5317 (N_5317,N_1976,N_888);
nand U5318 (N_5318,N_1033,N_2590);
or U5319 (N_5319,N_2357,N_2902);
and U5320 (N_5320,N_2395,N_1285);
nand U5321 (N_5321,N_1546,N_2688);
nor U5322 (N_5322,N_229,N_570);
nor U5323 (N_5323,N_416,N_1040);
and U5324 (N_5324,N_2983,N_2401);
nor U5325 (N_5325,N_1949,N_1377);
nand U5326 (N_5326,N_1165,N_1978);
and U5327 (N_5327,N_2980,N_17);
nor U5328 (N_5328,N_2112,N_774);
nor U5329 (N_5329,N_1044,N_90);
and U5330 (N_5330,N_2262,N_690);
nor U5331 (N_5331,N_654,N_2634);
and U5332 (N_5332,N_2709,N_1526);
nor U5333 (N_5333,N_1,N_1089);
nor U5334 (N_5334,N_1940,N_1176);
nand U5335 (N_5335,N_1961,N_2681);
nor U5336 (N_5336,N_257,N_915);
nand U5337 (N_5337,N_2749,N_1051);
nand U5338 (N_5338,N_2567,N_1033);
or U5339 (N_5339,N_2501,N_1597);
and U5340 (N_5340,N_1775,N_1719);
nor U5341 (N_5341,N_2011,N_2782);
and U5342 (N_5342,N_2998,N_979);
and U5343 (N_5343,N_2641,N_847);
nor U5344 (N_5344,N_2019,N_505);
and U5345 (N_5345,N_1856,N_5);
nor U5346 (N_5346,N_141,N_1244);
nor U5347 (N_5347,N_157,N_1330);
and U5348 (N_5348,N_1325,N_1145);
and U5349 (N_5349,N_714,N_975);
nor U5350 (N_5350,N_111,N_462);
and U5351 (N_5351,N_1151,N_1871);
or U5352 (N_5352,N_977,N_2514);
or U5353 (N_5353,N_2029,N_2858);
nand U5354 (N_5354,N_2024,N_1286);
or U5355 (N_5355,N_1117,N_731);
and U5356 (N_5356,N_358,N_120);
and U5357 (N_5357,N_1294,N_1336);
and U5358 (N_5358,N_726,N_981);
nand U5359 (N_5359,N_1020,N_2516);
nor U5360 (N_5360,N_1450,N_1036);
and U5361 (N_5361,N_2086,N_431);
nand U5362 (N_5362,N_2488,N_1731);
and U5363 (N_5363,N_2592,N_1037);
nor U5364 (N_5364,N_1401,N_1627);
nor U5365 (N_5365,N_1296,N_1854);
or U5366 (N_5366,N_604,N_526);
nand U5367 (N_5367,N_574,N_1182);
or U5368 (N_5368,N_881,N_2212);
nand U5369 (N_5369,N_2428,N_2829);
nor U5370 (N_5370,N_1864,N_504);
and U5371 (N_5371,N_2284,N_1955);
nand U5372 (N_5372,N_2695,N_2847);
or U5373 (N_5373,N_2531,N_2148);
or U5374 (N_5374,N_1401,N_1102);
or U5375 (N_5375,N_576,N_2819);
and U5376 (N_5376,N_382,N_2703);
or U5377 (N_5377,N_298,N_2893);
or U5378 (N_5378,N_1124,N_404);
and U5379 (N_5379,N_1321,N_47);
nand U5380 (N_5380,N_1821,N_1628);
or U5381 (N_5381,N_1022,N_1086);
nor U5382 (N_5382,N_698,N_2422);
nor U5383 (N_5383,N_491,N_2271);
or U5384 (N_5384,N_608,N_1688);
and U5385 (N_5385,N_1720,N_2280);
and U5386 (N_5386,N_858,N_1830);
nand U5387 (N_5387,N_2962,N_2812);
and U5388 (N_5388,N_2147,N_1571);
or U5389 (N_5389,N_78,N_2477);
nor U5390 (N_5390,N_169,N_240);
nor U5391 (N_5391,N_982,N_1686);
and U5392 (N_5392,N_202,N_2382);
nor U5393 (N_5393,N_2253,N_1197);
nor U5394 (N_5394,N_1934,N_262);
nor U5395 (N_5395,N_17,N_788);
or U5396 (N_5396,N_2466,N_1599);
and U5397 (N_5397,N_138,N_2997);
nand U5398 (N_5398,N_2048,N_1296);
and U5399 (N_5399,N_1301,N_1497);
nor U5400 (N_5400,N_2213,N_2016);
nor U5401 (N_5401,N_449,N_2305);
nand U5402 (N_5402,N_1081,N_227);
and U5403 (N_5403,N_1312,N_2861);
nor U5404 (N_5404,N_1045,N_1041);
xnor U5405 (N_5405,N_369,N_2722);
nand U5406 (N_5406,N_88,N_280);
nor U5407 (N_5407,N_155,N_1161);
nand U5408 (N_5408,N_2020,N_2478);
nor U5409 (N_5409,N_280,N_1886);
nor U5410 (N_5410,N_684,N_1236);
or U5411 (N_5411,N_284,N_2500);
or U5412 (N_5412,N_426,N_2975);
and U5413 (N_5413,N_1386,N_1409);
and U5414 (N_5414,N_1397,N_1486);
and U5415 (N_5415,N_594,N_162);
or U5416 (N_5416,N_1533,N_2027);
or U5417 (N_5417,N_447,N_1);
or U5418 (N_5418,N_290,N_2237);
or U5419 (N_5419,N_33,N_264);
nand U5420 (N_5420,N_98,N_534);
and U5421 (N_5421,N_1167,N_248);
nor U5422 (N_5422,N_1492,N_2294);
or U5423 (N_5423,N_2753,N_1522);
or U5424 (N_5424,N_882,N_2793);
or U5425 (N_5425,N_297,N_1895);
nand U5426 (N_5426,N_2423,N_2067);
and U5427 (N_5427,N_927,N_1604);
nand U5428 (N_5428,N_2826,N_970);
and U5429 (N_5429,N_356,N_1267);
and U5430 (N_5430,N_1833,N_575);
nand U5431 (N_5431,N_2403,N_2973);
or U5432 (N_5432,N_2204,N_1538);
nand U5433 (N_5433,N_384,N_1231);
nor U5434 (N_5434,N_2796,N_1744);
and U5435 (N_5435,N_802,N_1510);
and U5436 (N_5436,N_2307,N_1064);
and U5437 (N_5437,N_297,N_47);
or U5438 (N_5438,N_2467,N_1283);
or U5439 (N_5439,N_1429,N_1463);
nor U5440 (N_5440,N_2686,N_2655);
or U5441 (N_5441,N_2777,N_424);
nand U5442 (N_5442,N_1440,N_1346);
and U5443 (N_5443,N_2542,N_1567);
or U5444 (N_5444,N_547,N_2227);
nand U5445 (N_5445,N_2832,N_1666);
nand U5446 (N_5446,N_1550,N_974);
and U5447 (N_5447,N_1788,N_1644);
or U5448 (N_5448,N_2141,N_80);
and U5449 (N_5449,N_2011,N_740);
and U5450 (N_5450,N_1134,N_2218);
nand U5451 (N_5451,N_2760,N_736);
and U5452 (N_5452,N_275,N_1101);
nor U5453 (N_5453,N_1690,N_1944);
and U5454 (N_5454,N_686,N_616);
nor U5455 (N_5455,N_1958,N_408);
or U5456 (N_5456,N_744,N_2890);
and U5457 (N_5457,N_2859,N_2401);
nand U5458 (N_5458,N_2151,N_2570);
xor U5459 (N_5459,N_2193,N_2354);
or U5460 (N_5460,N_1148,N_264);
and U5461 (N_5461,N_2565,N_2928);
and U5462 (N_5462,N_851,N_92);
and U5463 (N_5463,N_1200,N_1296);
nor U5464 (N_5464,N_2485,N_469);
or U5465 (N_5465,N_310,N_818);
nand U5466 (N_5466,N_588,N_1466);
or U5467 (N_5467,N_936,N_1197);
or U5468 (N_5468,N_410,N_2922);
or U5469 (N_5469,N_2303,N_1144);
and U5470 (N_5470,N_1276,N_1375);
and U5471 (N_5471,N_2779,N_2494);
nor U5472 (N_5472,N_125,N_1275);
or U5473 (N_5473,N_601,N_2145);
nand U5474 (N_5474,N_2325,N_2426);
or U5475 (N_5475,N_648,N_2592);
nor U5476 (N_5476,N_474,N_1585);
or U5477 (N_5477,N_504,N_223);
nor U5478 (N_5478,N_2093,N_611);
nor U5479 (N_5479,N_1433,N_1182);
or U5480 (N_5480,N_2683,N_1046);
and U5481 (N_5481,N_1889,N_1640);
nor U5482 (N_5482,N_2896,N_2240);
nand U5483 (N_5483,N_2666,N_1306);
nor U5484 (N_5484,N_1169,N_2911);
or U5485 (N_5485,N_1770,N_724);
nand U5486 (N_5486,N_2683,N_2614);
or U5487 (N_5487,N_2159,N_515);
nor U5488 (N_5488,N_2095,N_93);
nand U5489 (N_5489,N_1673,N_2856);
nor U5490 (N_5490,N_1391,N_1976);
nand U5491 (N_5491,N_1218,N_509);
nand U5492 (N_5492,N_430,N_792);
or U5493 (N_5493,N_2070,N_653);
and U5494 (N_5494,N_2962,N_2168);
nand U5495 (N_5495,N_2410,N_2698);
nand U5496 (N_5496,N_206,N_2494);
nor U5497 (N_5497,N_1874,N_2062);
nor U5498 (N_5498,N_2598,N_2293);
or U5499 (N_5499,N_1408,N_1518);
and U5500 (N_5500,N_2675,N_2927);
nand U5501 (N_5501,N_267,N_2295);
nor U5502 (N_5502,N_2199,N_2282);
or U5503 (N_5503,N_1070,N_2378);
nand U5504 (N_5504,N_373,N_1967);
and U5505 (N_5505,N_2524,N_1552);
and U5506 (N_5506,N_853,N_496);
or U5507 (N_5507,N_2035,N_2092);
nor U5508 (N_5508,N_1425,N_2147);
nand U5509 (N_5509,N_150,N_330);
or U5510 (N_5510,N_835,N_96);
nand U5511 (N_5511,N_1362,N_2364);
and U5512 (N_5512,N_2832,N_2494);
and U5513 (N_5513,N_32,N_875);
and U5514 (N_5514,N_2226,N_2886);
nand U5515 (N_5515,N_2476,N_1823);
or U5516 (N_5516,N_551,N_2398);
nor U5517 (N_5517,N_1138,N_1850);
and U5518 (N_5518,N_1136,N_1284);
nand U5519 (N_5519,N_1209,N_88);
or U5520 (N_5520,N_577,N_1280);
nor U5521 (N_5521,N_2261,N_1074);
and U5522 (N_5522,N_1536,N_2464);
or U5523 (N_5523,N_180,N_2601);
and U5524 (N_5524,N_1927,N_754);
nand U5525 (N_5525,N_2113,N_2544);
or U5526 (N_5526,N_2681,N_1464);
or U5527 (N_5527,N_1347,N_2951);
and U5528 (N_5528,N_2269,N_2380);
nand U5529 (N_5529,N_152,N_1447);
and U5530 (N_5530,N_736,N_1320);
or U5531 (N_5531,N_1978,N_508);
nand U5532 (N_5532,N_2064,N_2964);
or U5533 (N_5533,N_2896,N_209);
or U5534 (N_5534,N_1794,N_1699);
or U5535 (N_5535,N_494,N_1425);
nor U5536 (N_5536,N_1161,N_2216);
or U5537 (N_5537,N_1747,N_594);
nand U5538 (N_5538,N_1643,N_2953);
or U5539 (N_5539,N_1976,N_1472);
nor U5540 (N_5540,N_815,N_130);
or U5541 (N_5541,N_89,N_298);
nor U5542 (N_5542,N_1435,N_2107);
or U5543 (N_5543,N_2788,N_1943);
nand U5544 (N_5544,N_2578,N_1346);
or U5545 (N_5545,N_1702,N_937);
nor U5546 (N_5546,N_2297,N_2399);
nand U5547 (N_5547,N_260,N_487);
nor U5548 (N_5548,N_2966,N_551);
and U5549 (N_5549,N_137,N_2592);
nor U5550 (N_5550,N_220,N_2355);
or U5551 (N_5551,N_385,N_2559);
nand U5552 (N_5552,N_1361,N_1844);
nand U5553 (N_5553,N_1458,N_2211);
nor U5554 (N_5554,N_561,N_1182);
xor U5555 (N_5555,N_877,N_491);
nand U5556 (N_5556,N_1153,N_2413);
and U5557 (N_5557,N_2878,N_1470);
nor U5558 (N_5558,N_2275,N_1403);
nor U5559 (N_5559,N_2173,N_2446);
or U5560 (N_5560,N_545,N_1808);
nor U5561 (N_5561,N_2042,N_731);
or U5562 (N_5562,N_533,N_382);
or U5563 (N_5563,N_2505,N_454);
or U5564 (N_5564,N_1249,N_2620);
and U5565 (N_5565,N_265,N_605);
nand U5566 (N_5566,N_1511,N_2935);
xnor U5567 (N_5567,N_1531,N_2343);
and U5568 (N_5568,N_2436,N_1475);
nand U5569 (N_5569,N_1947,N_490);
nand U5570 (N_5570,N_1817,N_1980);
and U5571 (N_5571,N_1600,N_2100);
nand U5572 (N_5572,N_602,N_2722);
and U5573 (N_5573,N_2476,N_909);
and U5574 (N_5574,N_2494,N_951);
nor U5575 (N_5575,N_1749,N_965);
or U5576 (N_5576,N_370,N_1046);
or U5577 (N_5577,N_530,N_2320);
or U5578 (N_5578,N_2459,N_2833);
nand U5579 (N_5579,N_2301,N_2760);
nand U5580 (N_5580,N_451,N_2391);
nor U5581 (N_5581,N_906,N_1035);
nor U5582 (N_5582,N_143,N_1979);
and U5583 (N_5583,N_1990,N_1298);
nand U5584 (N_5584,N_2769,N_289);
nor U5585 (N_5585,N_1256,N_1950);
and U5586 (N_5586,N_2875,N_1911);
and U5587 (N_5587,N_2663,N_137);
and U5588 (N_5588,N_2872,N_2519);
or U5589 (N_5589,N_2950,N_2927);
nand U5590 (N_5590,N_2631,N_2913);
or U5591 (N_5591,N_40,N_2589);
or U5592 (N_5592,N_137,N_1823);
or U5593 (N_5593,N_1329,N_1170);
and U5594 (N_5594,N_1854,N_2531);
nor U5595 (N_5595,N_771,N_231);
nor U5596 (N_5596,N_1505,N_958);
nor U5597 (N_5597,N_409,N_975);
nand U5598 (N_5598,N_2880,N_511);
and U5599 (N_5599,N_1996,N_2674);
nand U5600 (N_5600,N_2205,N_2207);
or U5601 (N_5601,N_1211,N_1573);
and U5602 (N_5602,N_872,N_1309);
xnor U5603 (N_5603,N_780,N_2275);
and U5604 (N_5604,N_720,N_1020);
and U5605 (N_5605,N_1386,N_1987);
or U5606 (N_5606,N_2149,N_2958);
nand U5607 (N_5607,N_1196,N_2964);
or U5608 (N_5608,N_2753,N_1610);
nand U5609 (N_5609,N_759,N_716);
and U5610 (N_5610,N_1327,N_1428);
or U5611 (N_5611,N_867,N_2447);
nor U5612 (N_5612,N_2917,N_2378);
nand U5613 (N_5613,N_1883,N_2516);
or U5614 (N_5614,N_1,N_1190);
nand U5615 (N_5615,N_387,N_366);
and U5616 (N_5616,N_1087,N_942);
or U5617 (N_5617,N_2236,N_1056);
and U5618 (N_5618,N_1778,N_734);
nor U5619 (N_5619,N_25,N_1620);
or U5620 (N_5620,N_2539,N_2561);
nand U5621 (N_5621,N_1298,N_2008);
or U5622 (N_5622,N_2723,N_448);
nor U5623 (N_5623,N_812,N_1345);
and U5624 (N_5624,N_249,N_1438);
nor U5625 (N_5625,N_1587,N_1645);
nand U5626 (N_5626,N_2117,N_2423);
or U5627 (N_5627,N_1950,N_2802);
nor U5628 (N_5628,N_2968,N_1442);
and U5629 (N_5629,N_1689,N_819);
or U5630 (N_5630,N_562,N_1025);
nand U5631 (N_5631,N_1809,N_1138);
and U5632 (N_5632,N_306,N_954);
nand U5633 (N_5633,N_2079,N_2573);
nor U5634 (N_5634,N_462,N_1878);
nor U5635 (N_5635,N_729,N_2317);
and U5636 (N_5636,N_897,N_116);
or U5637 (N_5637,N_844,N_796);
and U5638 (N_5638,N_1236,N_1071);
or U5639 (N_5639,N_78,N_908);
or U5640 (N_5640,N_2202,N_923);
nand U5641 (N_5641,N_100,N_94);
and U5642 (N_5642,N_1534,N_1606);
and U5643 (N_5643,N_1758,N_647);
nand U5644 (N_5644,N_1828,N_22);
nand U5645 (N_5645,N_736,N_1900);
nor U5646 (N_5646,N_1127,N_1752);
nor U5647 (N_5647,N_2191,N_1062);
or U5648 (N_5648,N_1931,N_981);
and U5649 (N_5649,N_2872,N_202);
nand U5650 (N_5650,N_2611,N_291);
nor U5651 (N_5651,N_2661,N_840);
and U5652 (N_5652,N_181,N_937);
nand U5653 (N_5653,N_1377,N_2775);
or U5654 (N_5654,N_2620,N_2718);
nor U5655 (N_5655,N_2226,N_2076);
xor U5656 (N_5656,N_207,N_1274);
nand U5657 (N_5657,N_2477,N_1739);
nor U5658 (N_5658,N_648,N_1661);
and U5659 (N_5659,N_2766,N_240);
nor U5660 (N_5660,N_1553,N_1674);
or U5661 (N_5661,N_2071,N_1068);
or U5662 (N_5662,N_578,N_746);
nand U5663 (N_5663,N_1276,N_2740);
or U5664 (N_5664,N_1553,N_1943);
or U5665 (N_5665,N_2429,N_1210);
nand U5666 (N_5666,N_2462,N_980);
and U5667 (N_5667,N_1272,N_2902);
or U5668 (N_5668,N_625,N_1012);
or U5669 (N_5669,N_2631,N_577);
or U5670 (N_5670,N_1656,N_1588);
or U5671 (N_5671,N_1665,N_2288);
or U5672 (N_5672,N_823,N_2995);
and U5673 (N_5673,N_2097,N_2956);
nand U5674 (N_5674,N_1944,N_1322);
and U5675 (N_5675,N_344,N_2661);
nor U5676 (N_5676,N_2706,N_2156);
nor U5677 (N_5677,N_389,N_1906);
and U5678 (N_5678,N_2438,N_2824);
and U5679 (N_5679,N_2469,N_2866);
or U5680 (N_5680,N_1398,N_277);
or U5681 (N_5681,N_162,N_274);
or U5682 (N_5682,N_2950,N_998);
or U5683 (N_5683,N_942,N_2534);
or U5684 (N_5684,N_2551,N_433);
nand U5685 (N_5685,N_1573,N_264);
and U5686 (N_5686,N_1386,N_1568);
or U5687 (N_5687,N_459,N_1183);
or U5688 (N_5688,N_1407,N_2878);
or U5689 (N_5689,N_1008,N_2771);
or U5690 (N_5690,N_2953,N_2445);
or U5691 (N_5691,N_500,N_2936);
or U5692 (N_5692,N_2023,N_1476);
or U5693 (N_5693,N_1601,N_1028);
nor U5694 (N_5694,N_851,N_1690);
nand U5695 (N_5695,N_2532,N_413);
or U5696 (N_5696,N_1561,N_1382);
or U5697 (N_5697,N_1969,N_858);
nor U5698 (N_5698,N_2748,N_2078);
or U5699 (N_5699,N_2364,N_179);
and U5700 (N_5700,N_2642,N_2556);
nor U5701 (N_5701,N_1814,N_1329);
and U5702 (N_5702,N_769,N_453);
and U5703 (N_5703,N_2280,N_1634);
nor U5704 (N_5704,N_685,N_2609);
nor U5705 (N_5705,N_2685,N_1357);
nand U5706 (N_5706,N_1923,N_1595);
or U5707 (N_5707,N_564,N_2542);
nand U5708 (N_5708,N_1344,N_1393);
nor U5709 (N_5709,N_2961,N_2286);
or U5710 (N_5710,N_981,N_689);
nor U5711 (N_5711,N_1862,N_528);
and U5712 (N_5712,N_1824,N_1152);
and U5713 (N_5713,N_1589,N_1618);
nand U5714 (N_5714,N_1810,N_1699);
or U5715 (N_5715,N_2833,N_751);
or U5716 (N_5716,N_1651,N_2650);
nand U5717 (N_5717,N_1347,N_1737);
nand U5718 (N_5718,N_251,N_2380);
or U5719 (N_5719,N_1191,N_901);
nand U5720 (N_5720,N_2500,N_2111);
nand U5721 (N_5721,N_2578,N_1825);
nor U5722 (N_5722,N_1690,N_203);
or U5723 (N_5723,N_790,N_1525);
nand U5724 (N_5724,N_1047,N_1558);
nor U5725 (N_5725,N_1223,N_2110);
xnor U5726 (N_5726,N_1529,N_2548);
and U5727 (N_5727,N_219,N_2199);
or U5728 (N_5728,N_1110,N_1692);
nand U5729 (N_5729,N_2100,N_948);
or U5730 (N_5730,N_2128,N_528);
nor U5731 (N_5731,N_2071,N_1928);
nor U5732 (N_5732,N_1181,N_504);
or U5733 (N_5733,N_711,N_687);
or U5734 (N_5734,N_1803,N_2456);
nor U5735 (N_5735,N_1310,N_747);
and U5736 (N_5736,N_1666,N_598);
nand U5737 (N_5737,N_1941,N_2238);
or U5738 (N_5738,N_274,N_1078);
and U5739 (N_5739,N_153,N_793);
nor U5740 (N_5740,N_893,N_2779);
or U5741 (N_5741,N_2444,N_1461);
or U5742 (N_5742,N_1803,N_1900);
nand U5743 (N_5743,N_2502,N_2433);
nand U5744 (N_5744,N_2854,N_2937);
nor U5745 (N_5745,N_640,N_2542);
nand U5746 (N_5746,N_2892,N_2156);
nor U5747 (N_5747,N_2202,N_412);
or U5748 (N_5748,N_2362,N_1539);
nor U5749 (N_5749,N_658,N_1684);
or U5750 (N_5750,N_2384,N_496);
and U5751 (N_5751,N_1459,N_2890);
nor U5752 (N_5752,N_1968,N_629);
and U5753 (N_5753,N_2095,N_1994);
nand U5754 (N_5754,N_2921,N_663);
nand U5755 (N_5755,N_2101,N_1809);
nand U5756 (N_5756,N_581,N_235);
or U5757 (N_5757,N_459,N_2164);
and U5758 (N_5758,N_2692,N_1754);
or U5759 (N_5759,N_1928,N_18);
nor U5760 (N_5760,N_4,N_708);
nor U5761 (N_5761,N_1181,N_1171);
nor U5762 (N_5762,N_404,N_2105);
nand U5763 (N_5763,N_2772,N_870);
or U5764 (N_5764,N_1851,N_1643);
nor U5765 (N_5765,N_311,N_2608);
nand U5766 (N_5766,N_1109,N_1778);
nor U5767 (N_5767,N_1178,N_467);
nor U5768 (N_5768,N_208,N_2696);
or U5769 (N_5769,N_1890,N_1342);
nand U5770 (N_5770,N_2781,N_854);
or U5771 (N_5771,N_2260,N_1477);
and U5772 (N_5772,N_585,N_2552);
nand U5773 (N_5773,N_2225,N_2082);
xnor U5774 (N_5774,N_2150,N_1633);
xor U5775 (N_5775,N_660,N_1779);
nor U5776 (N_5776,N_1780,N_1065);
or U5777 (N_5777,N_1841,N_1646);
nand U5778 (N_5778,N_2206,N_758);
nor U5779 (N_5779,N_1595,N_2073);
and U5780 (N_5780,N_1863,N_302);
nor U5781 (N_5781,N_1967,N_456);
nand U5782 (N_5782,N_668,N_2526);
or U5783 (N_5783,N_2,N_603);
or U5784 (N_5784,N_2052,N_1598);
nand U5785 (N_5785,N_116,N_1692);
and U5786 (N_5786,N_2661,N_763);
and U5787 (N_5787,N_892,N_999);
nor U5788 (N_5788,N_703,N_212);
nor U5789 (N_5789,N_1160,N_2438);
nor U5790 (N_5790,N_1975,N_930);
nor U5791 (N_5791,N_618,N_75);
nand U5792 (N_5792,N_572,N_1702);
nand U5793 (N_5793,N_839,N_2653);
nor U5794 (N_5794,N_1678,N_2785);
and U5795 (N_5795,N_2424,N_230);
nand U5796 (N_5796,N_650,N_1133);
and U5797 (N_5797,N_365,N_957);
and U5798 (N_5798,N_1095,N_2695);
and U5799 (N_5799,N_1830,N_1205);
nand U5800 (N_5800,N_690,N_2495);
nand U5801 (N_5801,N_2926,N_651);
or U5802 (N_5802,N_86,N_1508);
nand U5803 (N_5803,N_2324,N_792);
nand U5804 (N_5804,N_1119,N_2239);
nor U5805 (N_5805,N_534,N_807);
and U5806 (N_5806,N_1456,N_2614);
nand U5807 (N_5807,N_2625,N_1825);
nand U5808 (N_5808,N_1203,N_2910);
and U5809 (N_5809,N_656,N_686);
nand U5810 (N_5810,N_955,N_2692);
or U5811 (N_5811,N_1761,N_455);
or U5812 (N_5812,N_1166,N_1937);
or U5813 (N_5813,N_1264,N_1418);
and U5814 (N_5814,N_1497,N_2687);
and U5815 (N_5815,N_1456,N_1644);
nand U5816 (N_5816,N_703,N_40);
and U5817 (N_5817,N_1622,N_572);
nand U5818 (N_5818,N_1792,N_503);
nand U5819 (N_5819,N_1035,N_2543);
or U5820 (N_5820,N_409,N_2338);
nor U5821 (N_5821,N_68,N_175);
nand U5822 (N_5822,N_1440,N_1936);
nand U5823 (N_5823,N_2617,N_782);
and U5824 (N_5824,N_2136,N_895);
nor U5825 (N_5825,N_1800,N_1136);
nor U5826 (N_5826,N_271,N_1356);
and U5827 (N_5827,N_131,N_2096);
nor U5828 (N_5828,N_223,N_1944);
nand U5829 (N_5829,N_1858,N_2538);
nand U5830 (N_5830,N_2896,N_2671);
nand U5831 (N_5831,N_2843,N_2042);
and U5832 (N_5832,N_2862,N_2035);
or U5833 (N_5833,N_2649,N_1967);
nor U5834 (N_5834,N_2499,N_2570);
or U5835 (N_5835,N_2904,N_946);
nor U5836 (N_5836,N_1852,N_214);
and U5837 (N_5837,N_2139,N_1236);
nor U5838 (N_5838,N_1748,N_1699);
nor U5839 (N_5839,N_1433,N_2796);
or U5840 (N_5840,N_306,N_2272);
or U5841 (N_5841,N_765,N_416);
or U5842 (N_5842,N_61,N_2931);
nand U5843 (N_5843,N_1644,N_144);
nand U5844 (N_5844,N_1818,N_1408);
nand U5845 (N_5845,N_1162,N_1721);
nor U5846 (N_5846,N_1437,N_633);
and U5847 (N_5847,N_557,N_318);
or U5848 (N_5848,N_457,N_535);
nor U5849 (N_5849,N_551,N_1697);
and U5850 (N_5850,N_1918,N_1317);
xnor U5851 (N_5851,N_2456,N_1938);
nor U5852 (N_5852,N_674,N_333);
or U5853 (N_5853,N_2026,N_206);
and U5854 (N_5854,N_256,N_197);
xor U5855 (N_5855,N_2687,N_1299);
or U5856 (N_5856,N_1339,N_1928);
and U5857 (N_5857,N_2639,N_1340);
nand U5858 (N_5858,N_2040,N_987);
nor U5859 (N_5859,N_1264,N_1762);
or U5860 (N_5860,N_2198,N_1118);
nand U5861 (N_5861,N_657,N_1734);
nand U5862 (N_5862,N_1963,N_295);
nand U5863 (N_5863,N_2266,N_175);
nor U5864 (N_5864,N_1848,N_2288);
xnor U5865 (N_5865,N_2011,N_2638);
nor U5866 (N_5866,N_1686,N_440);
and U5867 (N_5867,N_1064,N_2177);
nand U5868 (N_5868,N_1573,N_943);
and U5869 (N_5869,N_1361,N_2149);
or U5870 (N_5870,N_1759,N_1541);
nand U5871 (N_5871,N_126,N_28);
and U5872 (N_5872,N_1273,N_2736);
and U5873 (N_5873,N_1845,N_998);
nor U5874 (N_5874,N_1885,N_1063);
nand U5875 (N_5875,N_2948,N_2347);
nand U5876 (N_5876,N_450,N_329);
and U5877 (N_5877,N_903,N_1180);
nand U5878 (N_5878,N_2649,N_2635);
nand U5879 (N_5879,N_1840,N_513);
or U5880 (N_5880,N_2768,N_2884);
or U5881 (N_5881,N_876,N_1483);
and U5882 (N_5882,N_1757,N_2144);
nand U5883 (N_5883,N_108,N_1904);
xnor U5884 (N_5884,N_745,N_1742);
nand U5885 (N_5885,N_926,N_251);
or U5886 (N_5886,N_1672,N_2486);
and U5887 (N_5887,N_1056,N_1308);
nor U5888 (N_5888,N_2345,N_2764);
and U5889 (N_5889,N_516,N_683);
nand U5890 (N_5890,N_212,N_291);
nand U5891 (N_5891,N_1130,N_2203);
and U5892 (N_5892,N_345,N_1001);
nor U5893 (N_5893,N_197,N_296);
nor U5894 (N_5894,N_2053,N_806);
nand U5895 (N_5895,N_911,N_1149);
nor U5896 (N_5896,N_2880,N_1483);
or U5897 (N_5897,N_2262,N_2362);
nor U5898 (N_5898,N_2506,N_2905);
and U5899 (N_5899,N_945,N_2584);
and U5900 (N_5900,N_408,N_675);
nand U5901 (N_5901,N_159,N_773);
nand U5902 (N_5902,N_2514,N_978);
and U5903 (N_5903,N_1266,N_3);
and U5904 (N_5904,N_377,N_438);
nor U5905 (N_5905,N_691,N_924);
or U5906 (N_5906,N_39,N_239);
nand U5907 (N_5907,N_323,N_1659);
nor U5908 (N_5908,N_342,N_1990);
nand U5909 (N_5909,N_2894,N_2032);
nand U5910 (N_5910,N_425,N_2128);
nor U5911 (N_5911,N_84,N_2957);
or U5912 (N_5912,N_262,N_2417);
nor U5913 (N_5913,N_2898,N_975);
or U5914 (N_5914,N_1724,N_2755);
nor U5915 (N_5915,N_716,N_1112);
nand U5916 (N_5916,N_2141,N_1579);
and U5917 (N_5917,N_1484,N_2675);
and U5918 (N_5918,N_2315,N_1113);
or U5919 (N_5919,N_1621,N_2625);
and U5920 (N_5920,N_2415,N_1074);
nand U5921 (N_5921,N_2880,N_789);
nand U5922 (N_5922,N_158,N_1529);
and U5923 (N_5923,N_2509,N_209);
nor U5924 (N_5924,N_425,N_1373);
nand U5925 (N_5925,N_222,N_959);
and U5926 (N_5926,N_1229,N_827);
nor U5927 (N_5927,N_735,N_486);
or U5928 (N_5928,N_370,N_2388);
or U5929 (N_5929,N_2082,N_1336);
and U5930 (N_5930,N_2871,N_2106);
and U5931 (N_5931,N_2259,N_193);
nor U5932 (N_5932,N_1948,N_634);
nor U5933 (N_5933,N_2088,N_2496);
or U5934 (N_5934,N_2493,N_1689);
nor U5935 (N_5935,N_1268,N_1691);
and U5936 (N_5936,N_1644,N_1936);
nor U5937 (N_5937,N_2875,N_1538);
nor U5938 (N_5938,N_783,N_2621);
or U5939 (N_5939,N_292,N_2799);
or U5940 (N_5940,N_2695,N_1587);
or U5941 (N_5941,N_280,N_1843);
and U5942 (N_5942,N_160,N_613);
nand U5943 (N_5943,N_574,N_1893);
nand U5944 (N_5944,N_1374,N_831);
and U5945 (N_5945,N_1323,N_468);
nor U5946 (N_5946,N_2886,N_1724);
nand U5947 (N_5947,N_627,N_892);
and U5948 (N_5948,N_2236,N_1698);
xnor U5949 (N_5949,N_2851,N_1902);
or U5950 (N_5950,N_1006,N_306);
and U5951 (N_5951,N_1865,N_807);
xnor U5952 (N_5952,N_2458,N_2889);
nor U5953 (N_5953,N_61,N_1556);
nand U5954 (N_5954,N_2265,N_1235);
nand U5955 (N_5955,N_2245,N_314);
or U5956 (N_5956,N_233,N_1708);
or U5957 (N_5957,N_1109,N_666);
and U5958 (N_5958,N_59,N_323);
nand U5959 (N_5959,N_2399,N_1495);
nand U5960 (N_5960,N_2944,N_393);
or U5961 (N_5961,N_211,N_1182);
and U5962 (N_5962,N_975,N_1985);
and U5963 (N_5963,N_1753,N_1593);
nor U5964 (N_5964,N_2457,N_2174);
nand U5965 (N_5965,N_2962,N_2815);
or U5966 (N_5966,N_2063,N_515);
or U5967 (N_5967,N_1578,N_965);
nor U5968 (N_5968,N_2431,N_1624);
and U5969 (N_5969,N_2136,N_2210);
and U5970 (N_5970,N_496,N_1148);
and U5971 (N_5971,N_2733,N_2392);
or U5972 (N_5972,N_1277,N_2789);
nand U5973 (N_5973,N_2263,N_2335);
and U5974 (N_5974,N_434,N_2860);
nand U5975 (N_5975,N_2550,N_1606);
and U5976 (N_5976,N_2045,N_144);
nand U5977 (N_5977,N_2813,N_925);
nor U5978 (N_5978,N_258,N_1842);
nand U5979 (N_5979,N_2910,N_2009);
nor U5980 (N_5980,N_1383,N_2150);
nand U5981 (N_5981,N_1309,N_2048);
nor U5982 (N_5982,N_763,N_1566);
or U5983 (N_5983,N_772,N_1427);
and U5984 (N_5984,N_2834,N_265);
and U5985 (N_5985,N_2756,N_332);
nor U5986 (N_5986,N_1263,N_49);
and U5987 (N_5987,N_2150,N_1019);
nor U5988 (N_5988,N_561,N_2286);
nand U5989 (N_5989,N_1737,N_588);
or U5990 (N_5990,N_2911,N_271);
or U5991 (N_5991,N_2615,N_499);
nand U5992 (N_5992,N_262,N_257);
and U5993 (N_5993,N_954,N_1700);
nand U5994 (N_5994,N_1306,N_470);
and U5995 (N_5995,N_153,N_2044);
or U5996 (N_5996,N_2752,N_2977);
or U5997 (N_5997,N_1826,N_268);
nor U5998 (N_5998,N_886,N_817);
nand U5999 (N_5999,N_461,N_1953);
or U6000 (N_6000,N_4023,N_4487);
or U6001 (N_6001,N_3772,N_4674);
nand U6002 (N_6002,N_4097,N_4806);
nor U6003 (N_6003,N_5984,N_5830);
or U6004 (N_6004,N_5923,N_5922);
or U6005 (N_6005,N_5309,N_5260);
and U6006 (N_6006,N_5913,N_5064);
nand U6007 (N_6007,N_4496,N_5137);
or U6008 (N_6008,N_3502,N_4515);
nor U6009 (N_6009,N_4316,N_5340);
nand U6010 (N_6010,N_4732,N_4885);
and U6011 (N_6011,N_3987,N_5669);
nand U6012 (N_6012,N_3775,N_3033);
and U6013 (N_6013,N_3169,N_3481);
or U6014 (N_6014,N_5865,N_4767);
and U6015 (N_6015,N_5039,N_4943);
and U6016 (N_6016,N_3439,N_5912);
nor U6017 (N_6017,N_5595,N_4893);
nor U6018 (N_6018,N_3803,N_5970);
or U6019 (N_6019,N_5818,N_5573);
and U6020 (N_6020,N_4070,N_3098);
nand U6021 (N_6021,N_3851,N_3570);
and U6022 (N_6022,N_4296,N_4998);
nand U6023 (N_6023,N_4176,N_3349);
and U6024 (N_6024,N_5797,N_3245);
or U6025 (N_6025,N_3348,N_5578);
and U6026 (N_6026,N_4925,N_4388);
or U6027 (N_6027,N_3027,N_5894);
nand U6028 (N_6028,N_3638,N_5386);
or U6029 (N_6029,N_4059,N_5085);
or U6030 (N_6030,N_5046,N_4094);
nand U6031 (N_6031,N_5798,N_5537);
nor U6032 (N_6032,N_5028,N_3694);
or U6033 (N_6033,N_3103,N_3361);
nor U6034 (N_6034,N_4877,N_5475);
and U6035 (N_6035,N_5559,N_3531);
or U6036 (N_6036,N_3629,N_4864);
and U6037 (N_6037,N_4154,N_3170);
and U6038 (N_6038,N_5479,N_5054);
nand U6039 (N_6039,N_4556,N_4549);
and U6040 (N_6040,N_5090,N_5400);
and U6041 (N_6041,N_5388,N_5393);
or U6042 (N_6042,N_5843,N_5379);
nand U6043 (N_6043,N_4051,N_4466);
and U6044 (N_6044,N_3087,N_4685);
xnor U6045 (N_6045,N_3028,N_5483);
and U6046 (N_6046,N_4262,N_5633);
nand U6047 (N_6047,N_4448,N_3300);
nand U6048 (N_6048,N_4841,N_5859);
nand U6049 (N_6049,N_3492,N_4259);
nand U6050 (N_6050,N_3143,N_3672);
nor U6051 (N_6051,N_3509,N_5642);
nor U6052 (N_6052,N_4571,N_5273);
or U6053 (N_6053,N_5957,N_5193);
and U6054 (N_6054,N_4505,N_3689);
nand U6055 (N_6055,N_4566,N_3206);
nor U6056 (N_6056,N_4681,N_3845);
nor U6057 (N_6057,N_4174,N_3462);
nand U6058 (N_6058,N_3903,N_4078);
or U6059 (N_6059,N_3266,N_4425);
nand U6060 (N_6060,N_3681,N_3271);
or U6061 (N_6061,N_3709,N_3830);
and U6062 (N_6062,N_4553,N_5574);
or U6063 (N_6063,N_5891,N_5766);
nand U6064 (N_6064,N_5493,N_3227);
xnor U6065 (N_6065,N_5083,N_3196);
nand U6066 (N_6066,N_3594,N_4802);
nand U6067 (N_6067,N_4382,N_4532);
nand U6068 (N_6068,N_5436,N_5285);
nor U6069 (N_6069,N_3399,N_4874);
nor U6070 (N_6070,N_3628,N_3096);
and U6071 (N_6071,N_5697,N_3343);
nand U6072 (N_6072,N_5211,N_3603);
or U6073 (N_6073,N_5422,N_4853);
nor U6074 (N_6074,N_4611,N_5986);
or U6075 (N_6075,N_4481,N_4246);
nand U6076 (N_6076,N_4062,N_3797);
nand U6077 (N_6077,N_5666,N_3102);
and U6078 (N_6078,N_4828,N_5074);
or U6079 (N_6079,N_3994,N_5895);
nor U6080 (N_6080,N_5394,N_5514);
nand U6081 (N_6081,N_3060,N_3303);
nand U6082 (N_6082,N_5786,N_4748);
and U6083 (N_6083,N_4695,N_3374);
and U6084 (N_6084,N_3036,N_5034);
nor U6085 (N_6085,N_5002,N_5238);
nand U6086 (N_6086,N_5860,N_5881);
nand U6087 (N_6087,N_4507,N_5529);
nor U6088 (N_6088,N_3981,N_5163);
nor U6089 (N_6089,N_5598,N_3781);
nor U6090 (N_6090,N_5761,N_5696);
nor U6091 (N_6091,N_3950,N_4536);
nor U6092 (N_6092,N_3722,N_5960);
nor U6093 (N_6093,N_4033,N_3770);
or U6094 (N_6094,N_5096,N_4380);
nor U6095 (N_6095,N_4441,N_4552);
and U6096 (N_6096,N_4095,N_3866);
nor U6097 (N_6097,N_3649,N_3560);
nand U6098 (N_6098,N_4029,N_3476);
or U6099 (N_6099,N_3010,N_5954);
and U6100 (N_6100,N_4191,N_5440);
and U6101 (N_6101,N_4288,N_5835);
nor U6102 (N_6102,N_3933,N_4941);
and U6103 (N_6103,N_5066,N_3634);
and U6104 (N_6104,N_4541,N_3274);
or U6105 (N_6105,N_5252,N_5177);
or U6106 (N_6106,N_3217,N_3575);
nand U6107 (N_6107,N_4865,N_5173);
nor U6108 (N_6108,N_5175,N_4689);
and U6109 (N_6109,N_5065,N_3627);
and U6110 (N_6110,N_5426,N_5180);
nor U6111 (N_6111,N_5992,N_4283);
nand U6112 (N_6112,N_4131,N_3872);
and U6113 (N_6113,N_4546,N_4432);
and U6114 (N_6114,N_5668,N_4445);
and U6115 (N_6115,N_3524,N_3061);
nor U6116 (N_6116,N_5239,N_3004);
or U6117 (N_6117,N_4821,N_3517);
or U6118 (N_6118,N_5369,N_5908);
nor U6119 (N_6119,N_4431,N_4374);
and U6120 (N_6120,N_3069,N_4212);
or U6121 (N_6121,N_5858,N_4135);
nand U6122 (N_6122,N_5953,N_4794);
and U6123 (N_6123,N_3841,N_4535);
nor U6124 (N_6124,N_3580,N_4780);
nand U6125 (N_6125,N_4114,N_4774);
nor U6126 (N_6126,N_4126,N_4121);
nor U6127 (N_6127,N_5518,N_5225);
and U6128 (N_6128,N_3717,N_4658);
nand U6129 (N_6129,N_4929,N_5741);
nor U6130 (N_6130,N_3136,N_3510);
or U6131 (N_6131,N_5032,N_3716);
and U6132 (N_6132,N_3958,N_5276);
nor U6133 (N_6133,N_5888,N_3112);
nor U6134 (N_6134,N_3937,N_3491);
and U6135 (N_6135,N_3949,N_3537);
and U6136 (N_6136,N_5156,N_5263);
and U6137 (N_6137,N_4547,N_3090);
and U6138 (N_6138,N_5435,N_4488);
nor U6139 (N_6139,N_4714,N_4285);
and U6140 (N_6140,N_3766,N_3968);
nand U6141 (N_6141,N_4851,N_5326);
nor U6142 (N_6142,N_5490,N_4087);
and U6143 (N_6143,N_4111,N_4236);
nand U6144 (N_6144,N_3359,N_3955);
and U6145 (N_6145,N_5725,N_5325);
nand U6146 (N_6146,N_3287,N_3768);
nor U6147 (N_6147,N_3737,N_4887);
nand U6148 (N_6148,N_4548,N_3615);
and U6149 (N_6149,N_4447,N_4254);
nand U6150 (N_6150,N_5628,N_3832);
nand U6151 (N_6151,N_4580,N_4719);
and U6152 (N_6152,N_3423,N_4103);
or U6153 (N_6153,N_4314,N_3870);
or U6154 (N_6154,N_4698,N_4178);
and U6155 (N_6155,N_3183,N_4971);
and U6156 (N_6156,N_5374,N_5773);
nor U6157 (N_6157,N_4902,N_5084);
and U6158 (N_6158,N_5370,N_4871);
nand U6159 (N_6159,N_3367,N_5680);
nor U6160 (N_6160,N_3003,N_4184);
or U6161 (N_6161,N_3424,N_3201);
nand U6162 (N_6162,N_3425,N_5763);
nor U6163 (N_6163,N_3504,N_4061);
nor U6164 (N_6164,N_3104,N_5407);
or U6165 (N_6165,N_5507,N_4733);
nand U6166 (N_6166,N_4644,N_3974);
or U6167 (N_6167,N_5201,N_5372);
and U6168 (N_6168,N_4579,N_5815);
and U6169 (N_6169,N_5900,N_3881);
nand U6170 (N_6170,N_5817,N_4375);
or U6171 (N_6171,N_5380,N_4915);
nand U6172 (N_6172,N_5148,N_5503);
or U6173 (N_6173,N_5232,N_3728);
or U6174 (N_6174,N_5994,N_5358);
or U6175 (N_6175,N_3602,N_4506);
and U6176 (N_6176,N_3733,N_5128);
or U6177 (N_6177,N_4589,N_3489);
or U6178 (N_6178,N_5088,N_3199);
and U6179 (N_6179,N_4758,N_4833);
nand U6180 (N_6180,N_5571,N_3801);
or U6181 (N_6181,N_3650,N_3444);
nand U6182 (N_6182,N_3308,N_4817);
or U6183 (N_6183,N_4083,N_4778);
xnor U6184 (N_6184,N_4226,N_3187);
and U6185 (N_6185,N_5760,N_4753);
nor U6186 (N_6186,N_5321,N_3880);
nand U6187 (N_6187,N_5251,N_4967);
and U6188 (N_6188,N_3472,N_5471);
nand U6189 (N_6189,N_3135,N_3166);
nand U6190 (N_6190,N_4798,N_5893);
nor U6191 (N_6191,N_4878,N_3970);
nor U6192 (N_6192,N_5233,N_3350);
nand U6193 (N_6193,N_5550,N_4002);
or U6194 (N_6194,N_5771,N_5496);
and U6195 (N_6195,N_3320,N_5676);
nor U6196 (N_6196,N_3018,N_3192);
nand U6197 (N_6197,N_3831,N_4215);
nor U6198 (N_6198,N_4010,N_4730);
nor U6199 (N_6199,N_3511,N_5863);
nand U6200 (N_6200,N_3918,N_5594);
nor U6201 (N_6201,N_4561,N_5318);
nor U6202 (N_6202,N_5467,N_3920);
and U6203 (N_6203,N_3683,N_3662);
or U6204 (N_6204,N_3236,N_3704);
or U6205 (N_6205,N_4771,N_3212);
or U6206 (N_6206,N_3333,N_5873);
nor U6207 (N_6207,N_5896,N_4735);
or U6208 (N_6208,N_3579,N_3820);
nor U6209 (N_6209,N_3805,N_3647);
nand U6210 (N_6210,N_3777,N_3487);
or U6211 (N_6211,N_5719,N_3268);
nor U6212 (N_6212,N_3860,N_5820);
and U6213 (N_6213,N_3473,N_4026);
nor U6214 (N_6214,N_3583,N_5008);
and U6215 (N_6215,N_4334,N_5995);
nor U6216 (N_6216,N_4075,N_4707);
nor U6217 (N_6217,N_3807,N_4227);
nand U6218 (N_6218,N_3743,N_3262);
and U6219 (N_6219,N_4142,N_4079);
nand U6220 (N_6220,N_3893,N_3241);
or U6221 (N_6221,N_4493,N_4870);
and U6222 (N_6222,N_4290,N_3248);
and U6223 (N_6223,N_3392,N_3942);
nor U6224 (N_6224,N_5807,N_5317);
or U6225 (N_6225,N_3284,N_4993);
nand U6226 (N_6226,N_3835,N_5538);
nand U6227 (N_6227,N_4233,N_5844);
xnor U6228 (N_6228,N_4945,N_3859);
or U6229 (N_6229,N_5651,N_4660);
nor U6230 (N_6230,N_4291,N_3152);
or U6231 (N_6231,N_4350,N_5653);
or U6232 (N_6232,N_4757,N_5051);
and U6233 (N_6233,N_4444,N_4298);
nor U6234 (N_6234,N_5183,N_5621);
nand U6235 (N_6235,N_4203,N_3815);
nor U6236 (N_6236,N_5919,N_4930);
nor U6237 (N_6237,N_5015,N_3309);
nor U6238 (N_6238,N_5799,N_3754);
nand U6239 (N_6239,N_5782,N_5434);
nand U6240 (N_6240,N_3984,N_3892);
or U6241 (N_6241,N_5904,N_5425);
nor U6242 (N_6242,N_3454,N_4610);
and U6243 (N_6243,N_5124,N_5781);
and U6244 (N_6244,N_3611,N_4472);
or U6245 (N_6245,N_3025,N_5087);
nor U6246 (N_6246,N_4020,N_4179);
and U6247 (N_6247,N_3895,N_5591);
nor U6248 (N_6248,N_5024,N_3837);
nor U6249 (N_6249,N_3175,N_5758);
nor U6250 (N_6250,N_3631,N_5498);
and U6251 (N_6251,N_4210,N_4725);
nor U6252 (N_6252,N_4844,N_4838);
nand U6253 (N_6253,N_5929,N_5775);
nor U6254 (N_6254,N_3637,N_3286);
nand U6255 (N_6255,N_3635,N_5772);
and U6256 (N_6256,N_3259,N_3936);
or U6257 (N_6257,N_4381,N_3393);
nand U6258 (N_6258,N_4934,N_4146);
or U6259 (N_6259,N_5816,N_5733);
nor U6260 (N_6260,N_5728,N_3547);
nor U6261 (N_6261,N_3549,N_4022);
or U6262 (N_6262,N_5041,N_3072);
nor U6263 (N_6263,N_5437,N_5332);
or U6264 (N_6264,N_3419,N_3500);
and U6265 (N_6265,N_5588,N_5787);
or U6266 (N_6266,N_5948,N_5966);
or U6267 (N_6267,N_5169,N_4379);
nand U6268 (N_6268,N_3989,N_3455);
nand U6269 (N_6269,N_3701,N_3324);
nor U6270 (N_6270,N_4608,N_4045);
nand U6271 (N_6271,N_4130,N_3769);
and U6272 (N_6272,N_3985,N_5940);
nor U6273 (N_6273,N_5840,N_5584);
and U6274 (N_6274,N_3301,N_5135);
nor U6275 (N_6275,N_3257,N_5445);
or U6276 (N_6276,N_5103,N_3493);
nor U6277 (N_6277,N_3605,N_5376);
or U6278 (N_6278,N_3999,N_3732);
or U6279 (N_6279,N_3179,N_3237);
and U6280 (N_6280,N_3412,N_5720);
and U6281 (N_6281,N_5679,N_4682);
nor U6282 (N_6282,N_5997,N_5266);
nand U6283 (N_6283,N_5981,N_3078);
and U6284 (N_6284,N_5967,N_4096);
or U6285 (N_6285,N_5812,N_4756);
nand U6286 (N_6286,N_5109,N_5810);
nor U6287 (N_6287,N_4152,N_4407);
and U6288 (N_6288,N_5298,N_3404);
nor U6289 (N_6289,N_5293,N_5911);
or U6290 (N_6290,N_4752,N_5539);
or U6291 (N_6291,N_3375,N_4139);
nor U6292 (N_6292,N_5833,N_4568);
nor U6293 (N_6293,N_4138,N_4718);
and U6294 (N_6294,N_3092,N_4416);
nand U6295 (N_6295,N_4105,N_5656);
or U6296 (N_6296,N_4906,N_5469);
nor U6297 (N_6297,N_5756,N_5557);
and U6298 (N_6298,N_5409,N_5737);
nor U6299 (N_6299,N_4463,N_4376);
or U6300 (N_6300,N_4462,N_3752);
and U6301 (N_6301,N_4976,N_5631);
nand U6302 (N_6302,N_4855,N_3868);
nand U6303 (N_6303,N_4265,N_5987);
nor U6304 (N_6304,N_4351,N_4005);
nand U6305 (N_6305,N_4827,N_5592);
and U6306 (N_6306,N_3558,N_5466);
nor U6307 (N_6307,N_5999,N_3120);
and U6308 (N_6308,N_4238,N_3244);
nor U6309 (N_6309,N_3313,N_4764);
nor U6310 (N_6310,N_3220,N_4413);
or U6311 (N_6311,N_4245,N_3535);
or U6312 (N_6312,N_4882,N_5307);
nand U6313 (N_6313,N_5226,N_5885);
nor U6314 (N_6314,N_4636,N_4517);
nand U6315 (N_6315,N_4908,N_4897);
and U6316 (N_6316,N_5164,N_3063);
and U6317 (N_6317,N_3787,N_5053);
nor U6318 (N_6318,N_3630,N_3038);
and U6319 (N_6319,N_4905,N_5221);
or U6320 (N_6320,N_4199,N_4795);
nand U6321 (N_6321,N_3661,N_5357);
nor U6322 (N_6322,N_4697,N_3840);
or U6323 (N_6323,N_3724,N_5520);
and U6324 (N_6324,N_5007,N_3198);
or U6325 (N_6325,N_4183,N_4938);
and U6326 (N_6326,N_5917,N_3031);
xor U6327 (N_6327,N_4072,N_5314);
and U6328 (N_6328,N_4560,N_4500);
nor U6329 (N_6329,N_4297,N_4286);
and U6330 (N_6330,N_4770,N_5724);
nand U6331 (N_6331,N_4522,N_4872);
and U6332 (N_6332,N_4955,N_3954);
nor U6333 (N_6333,N_5254,N_4278);
and U6334 (N_6334,N_4165,N_5459);
and U6335 (N_6335,N_3878,N_5921);
nand U6336 (N_6336,N_4516,N_4613);
nand U6337 (N_6337,N_3734,N_4836);
and U6338 (N_6338,N_4229,N_3572);
nor U6339 (N_6339,N_3026,N_5576);
or U6340 (N_6340,N_4692,N_4326);
nand U6341 (N_6341,N_5715,N_5387);
and U6342 (N_6342,N_5336,N_4504);
nor U6343 (N_6343,N_3358,N_4281);
nor U6344 (N_6344,N_5067,N_5670);
nand U6345 (N_6345,N_3645,N_3589);
nand U6346 (N_6346,N_3742,N_5202);
nor U6347 (N_6347,N_3821,N_5022);
xnor U6348 (N_6348,N_5077,N_3930);
nand U6349 (N_6349,N_4195,N_3048);
and U6350 (N_6350,N_5611,N_5218);
nor U6351 (N_6351,N_5274,N_3819);
or U6352 (N_6352,N_4663,N_5528);
and U6353 (N_6353,N_5246,N_4459);
or U6354 (N_6354,N_4875,N_5880);
and U6355 (N_6355,N_4973,N_4329);
and U6356 (N_6356,N_3883,N_5058);
or U6357 (N_6357,N_5916,N_3865);
nand U6358 (N_6358,N_4391,N_5602);
or U6359 (N_6359,N_5553,N_4703);
or U6360 (N_6360,N_3882,N_4578);
or U6361 (N_6361,N_3601,N_5448);
nor U6362 (N_6362,N_4442,N_3290);
nor U6363 (N_6363,N_3788,N_3746);
nor U6364 (N_6364,N_5214,N_5335);
nor U6365 (N_6365,N_3447,N_3402);
nor U6366 (N_6366,N_5794,N_4761);
nor U6367 (N_6367,N_4056,N_3624);
nor U6368 (N_6368,N_3600,N_5629);
nor U6369 (N_6369,N_4373,N_3996);
or U6370 (N_6370,N_3396,N_4551);
nor U6371 (N_6371,N_3824,N_3216);
or U6372 (N_6372,N_4662,N_5284);
or U6373 (N_6373,N_3543,N_4559);
nor U6374 (N_6374,N_3486,N_3713);
and U6375 (N_6375,N_5389,N_5215);
nor U6376 (N_6376,N_5489,N_4651);
and U6377 (N_6377,N_3498,N_5976);
nand U6378 (N_6378,N_5220,N_5521);
or U6379 (N_6379,N_5950,N_4918);
and U6380 (N_6380,N_3691,N_3180);
and U6381 (N_6381,N_5879,N_3867);
and U6382 (N_6382,N_3091,N_5207);
and U6383 (N_6383,N_4569,N_3520);
or U6384 (N_6384,N_4762,N_4818);
nor U6385 (N_6385,N_5410,N_4804);
nand U6386 (N_6386,N_3029,N_4016);
and U6387 (N_6387,N_4324,N_5412);
nor U6388 (N_6388,N_4687,N_3673);
or U6389 (N_6389,N_5461,N_3280);
nand U6390 (N_6390,N_5964,N_4922);
and U6391 (N_6391,N_4469,N_5726);
nand U6392 (N_6392,N_5150,N_4558);
or U6393 (N_6393,N_5308,N_3464);
and U6394 (N_6394,N_4498,N_5151);
and U6395 (N_6395,N_3696,N_3202);
nand U6396 (N_6396,N_5014,N_5470);
nor U6397 (N_6397,N_4367,N_4711);
or U6398 (N_6398,N_5925,N_4585);
nand U6399 (N_6399,N_3416,N_4881);
or U6400 (N_6400,N_5959,N_3363);
or U6401 (N_6401,N_5542,N_3850);
or U6402 (N_6402,N_4287,N_4228);
or U6403 (N_6403,N_3998,N_5327);
and U6404 (N_6404,N_3334,N_3298);
nand U6405 (N_6405,N_3101,N_4098);
nand U6406 (N_6406,N_5829,N_3478);
nand U6407 (N_6407,N_4230,N_4117);
and U6408 (N_6408,N_5564,N_4282);
and U6409 (N_6409,N_4502,N_5262);
nand U6410 (N_6410,N_4321,N_5158);
nor U6411 (N_6411,N_5581,N_4204);
nand U6412 (N_6412,N_3552,N_4599);
nand U6413 (N_6413,N_5117,N_4348);
and U6414 (N_6414,N_5431,N_4232);
nor U6415 (N_6415,N_3456,N_3430);
nand U6416 (N_6416,N_5005,N_4859);
or U6417 (N_6417,N_4653,N_3813);
and U6418 (N_6418,N_5482,N_5745);
or U6419 (N_6419,N_5453,N_4514);
or U6420 (N_6420,N_5295,N_3484);
and U6421 (N_6421,N_3762,N_4355);
or U6422 (N_6422,N_4039,N_5236);
and U6423 (N_6423,N_3686,N_3929);
or U6424 (N_6424,N_5013,N_5244);
nand U6425 (N_6425,N_5397,N_5938);
nand U6426 (N_6426,N_5228,N_5230);
nor U6427 (N_6427,N_3338,N_4073);
or U6428 (N_6428,N_5543,N_4899);
and U6429 (N_6429,N_5590,N_3723);
or U6430 (N_6430,N_5190,N_5035);
and U6431 (N_6431,N_3071,N_4418);
or U6432 (N_6432,N_3745,N_4605);
nor U6433 (N_6433,N_4144,N_5095);
nor U6434 (N_6434,N_4345,N_3826);
and U6435 (N_6435,N_5990,N_3928);
or U6436 (N_6436,N_4007,N_4995);
nand U6437 (N_6437,N_5749,N_5778);
nor U6438 (N_6438,N_5635,N_4429);
nand U6439 (N_6439,N_3014,N_5094);
nor U6440 (N_6440,N_3587,N_3213);
or U6441 (N_6441,N_5572,N_4276);
or U6442 (N_6442,N_4526,N_4582);
or U6443 (N_6443,N_4041,N_3794);
or U6444 (N_6444,N_5566,N_5416);
and U6445 (N_6445,N_3007,N_4940);
nor U6446 (N_6446,N_5497,N_3142);
nand U6447 (N_6447,N_4107,N_5905);
nor U6448 (N_6448,N_4977,N_5191);
xnor U6449 (N_6449,N_5777,N_4954);
or U6450 (N_6450,N_5918,N_4729);
and U6451 (N_6451,N_3253,N_3483);
nand U6452 (N_6452,N_4331,N_5439);
and U6453 (N_6453,N_4784,N_4615);
nand U6454 (N_6454,N_3879,N_5577);
or U6455 (N_6455,N_5910,N_3431);
nand U6456 (N_6456,N_3906,N_4596);
nand U6457 (N_6457,N_5750,N_4801);
or U6458 (N_6458,N_4337,N_4119);
and U6459 (N_6459,N_5256,N_5132);
nor U6460 (N_6460,N_4294,N_3032);
or U6461 (N_6461,N_4829,N_5890);
and U6462 (N_6462,N_5206,N_3506);
nor U6463 (N_6463,N_5296,N_3751);
or U6464 (N_6464,N_5324,N_4318);
nor U6465 (N_6465,N_4508,N_5247);
xnor U6466 (N_6466,N_3005,N_4034);
nand U6467 (N_6467,N_3076,N_5746);
nor U6468 (N_6468,N_3855,N_3049);
nor U6469 (N_6469,N_3773,N_4581);
nor U6470 (N_6470,N_4963,N_3222);
and U6471 (N_6471,N_5508,N_4303);
nand U6472 (N_6472,N_5029,N_3283);
nand U6473 (N_6473,N_4120,N_3362);
nor U6474 (N_6474,N_5160,N_5121);
nor U6475 (N_6475,N_4673,N_5650);
or U6476 (N_6476,N_3951,N_3780);
and U6477 (N_6477,N_3783,N_5418);
xnor U6478 (N_6478,N_4312,N_3158);
nor U6479 (N_6479,N_4437,N_4645);
and U6480 (N_6480,N_5433,N_4225);
or U6481 (N_6481,N_4339,N_4132);
nor U6482 (N_6482,N_3978,N_3767);
nor U6483 (N_6483,N_5362,N_5764);
or U6484 (N_6484,N_4724,N_3512);
nor U6485 (N_6485,N_5850,N_4340);
and U6486 (N_6486,N_5678,N_5849);
and U6487 (N_6487,N_5072,N_3708);
or U6488 (N_6488,N_3791,N_4793);
nand U6489 (N_6489,N_4216,N_3626);
nand U6490 (N_6490,N_3680,N_4598);
nand U6491 (N_6491,N_3771,N_3622);
and U6492 (N_6492,N_3731,N_3086);
and U6493 (N_6493,N_5612,N_4370);
and U6494 (N_6494,N_4792,N_4066);
nand U6495 (N_6495,N_3155,N_4606);
nand U6496 (N_6496,N_5037,N_3263);
nor U6497 (N_6497,N_4632,N_4365);
nand U6498 (N_6498,N_5610,N_4521);
or U6499 (N_6499,N_4177,N_5316);
or U6500 (N_6500,N_4538,N_5811);
nand U6501 (N_6501,N_5139,N_5546);
nand U6502 (N_6502,N_3051,N_5313);
nand U6503 (N_6503,N_4511,N_4457);
or U6504 (N_6504,N_5826,N_4788);
and U6505 (N_6505,N_3132,N_3501);
and U6506 (N_6506,N_3532,N_4361);
nor U6507 (N_6507,N_5854,N_4819);
and U6508 (N_6508,N_3138,N_4573);
or U6509 (N_6509,N_5579,N_3411);
and U6510 (N_6510,N_4439,N_3039);
xnor U6511 (N_6511,N_4832,N_4202);
or U6512 (N_6512,N_4394,N_5530);
or U6513 (N_6513,N_4654,N_4161);
nand U6514 (N_6514,N_5115,N_5257);
and U6515 (N_6515,N_5038,N_5375);
nand U6516 (N_6516,N_5455,N_3172);
nand U6517 (N_6517,N_3100,N_5017);
or U6518 (N_6518,N_3058,N_4395);
nor U6519 (N_6519,N_4019,N_4341);
nand U6520 (N_6520,N_4555,N_4058);
nand U6521 (N_6521,N_5060,N_4626);
and U6522 (N_6522,N_5189,N_3563);
and U6523 (N_6523,N_3931,N_3677);
nor U6524 (N_6524,N_3559,N_4475);
or U6525 (N_6525,N_3130,N_4602);
nand U6526 (N_6526,N_4933,N_4453);
and U6527 (N_6527,N_5457,N_3496);
nand U6528 (N_6528,N_4856,N_5305);
nor U6529 (N_6529,N_4055,N_3546);
nor U6530 (N_6530,N_5198,N_3385);
and U6531 (N_6531,N_3479,N_3068);
and U6532 (N_6532,N_3319,N_4134);
nor U6533 (N_6533,N_3093,N_5632);
nor U6534 (N_6534,N_5098,N_3621);
nor U6535 (N_6535,N_3946,N_4200);
nand U6536 (N_6536,N_5930,N_5162);
nand U6537 (N_6537,N_5702,N_5869);
nand U6538 (N_6538,N_3561,N_5998);
or U6539 (N_6539,N_3064,N_5499);
nor U6540 (N_6540,N_5451,N_5743);
or U6541 (N_6541,N_4972,N_4222);
and U6542 (N_6542,N_5971,N_4150);
and U6543 (N_6543,N_3381,N_4401);
or U6544 (N_6544,N_3000,N_3967);
and U6545 (N_6545,N_4251,N_5874);
and U6546 (N_6546,N_4627,N_4704);
and U6547 (N_6547,N_5876,N_3808);
nor U6548 (N_6548,N_3802,N_3551);
or U6549 (N_6549,N_3008,N_4525);
nand U6550 (N_6550,N_4570,N_5985);
or U6551 (N_6551,N_5286,N_4686);
nand U6552 (N_6552,N_3162,N_4797);
or U6553 (N_6553,N_3513,N_3668);
and U6554 (N_6554,N_3122,N_5946);
or U6555 (N_6555,N_4984,N_4846);
nor U6556 (N_6556,N_4402,N_3438);
or U6557 (N_6557,N_5078,N_4417);
nand U6558 (N_6558,N_5462,N_5277);
or U6559 (N_6559,N_3997,N_4478);
or U6560 (N_6560,N_3869,N_3642);
and U6561 (N_6561,N_5803,N_4389);
or U6562 (N_6562,N_4825,N_3299);
nand U6563 (N_6563,N_3659,N_4068);
nand U6564 (N_6564,N_3578,N_4313);
xnor U6565 (N_6565,N_5449,N_4182);
nand U6566 (N_6566,N_3796,N_5302);
nand U6567 (N_6567,N_3604,N_4562);
nor U6568 (N_6568,N_3962,N_5989);
and U6569 (N_6569,N_5655,N_4791);
nor U6570 (N_6570,N_5928,N_3089);
and U6571 (N_6571,N_5785,N_5235);
or U6572 (N_6572,N_4679,N_3593);
nand U6573 (N_6573,N_4641,N_4776);
nor U6574 (N_6574,N_4156,N_4700);
nand U6575 (N_6575,N_4968,N_5082);
nor U6576 (N_6576,N_3584,N_3530);
or U6577 (N_6577,N_3186,N_5603);
nand U6578 (N_6578,N_3368,N_5654);
nor U6579 (N_6579,N_5505,N_3034);
nor U6580 (N_6580,N_3469,N_4273);
or U6581 (N_6581,N_3674,N_5323);
nand U6582 (N_6582,N_4065,N_5188);
or U6583 (N_6583,N_4054,N_3853);
nand U6584 (N_6584,N_3226,N_3782);
nand U6585 (N_6585,N_3441,N_4385);
and U6586 (N_6586,N_5770,N_3526);
or U6587 (N_6587,N_4620,N_3065);
nand U6588 (N_6588,N_5730,N_4149);
nor U6589 (N_6589,N_4928,N_4163);
nor U6590 (N_6590,N_3934,N_5626);
or U6591 (N_6591,N_5933,N_5119);
nor U6592 (N_6592,N_4731,N_3176);
nor U6593 (N_6593,N_4647,N_3814);
nor U6594 (N_6594,N_4779,N_5381);
or U6595 (N_6595,N_4424,N_5345);
and U6596 (N_6596,N_4006,N_3988);
nand U6597 (N_6597,N_3239,N_3285);
nand U6598 (N_6598,N_4008,N_4952);
or U6599 (N_6599,N_3296,N_4812);
nor U6600 (N_6600,N_4001,N_3159);
or U6601 (N_6601,N_5937,N_4706);
or U6602 (N_6602,N_5243,N_4155);
and U6603 (N_6603,N_5662,N_5073);
nand U6604 (N_6604,N_5861,N_3718);
nor U6605 (N_6605,N_5774,N_3806);
and U6606 (N_6606,N_3311,N_5857);
or U6607 (N_6607,N_5338,N_4991);
or U6608 (N_6608,N_4497,N_3816);
nand U6609 (N_6609,N_4741,N_4076);
nand U6610 (N_6610,N_3596,N_4944);
nand U6611 (N_6611,N_5837,N_3682);
nand U6612 (N_6612,N_5329,N_5685);
or U6613 (N_6613,N_4648,N_3606);
and U6614 (N_6614,N_5601,N_5561);
nand U6615 (N_6615,N_5605,N_5665);
or U6616 (N_6616,N_3864,N_4064);
nand U6617 (N_6617,N_5753,N_4092);
nand U6618 (N_6618,N_3917,N_5924);
and U6619 (N_6619,N_4414,N_5597);
and U6620 (N_6620,N_3927,N_5776);
and U6621 (N_6621,N_4890,N_5171);
nor U6622 (N_6622,N_5645,N_3332);
nand U6623 (N_6623,N_4715,N_3926);
nand U6624 (N_6624,N_5502,N_4037);
nand U6625 (N_6625,N_5568,N_5618);
nor U6626 (N_6626,N_3157,N_3856);
and U6627 (N_6627,N_5884,N_3466);
nand U6628 (N_6628,N_4272,N_5047);
nand U6629 (N_6629,N_3658,N_4322);
nand U6630 (N_6630,N_4004,N_5902);
nand U6631 (N_6631,N_3203,N_3846);
and U6632 (N_6632,N_5149,N_5118);
nand U6633 (N_6633,N_3417,N_5209);
and U6634 (N_6634,N_3519,N_5570);
nand U6635 (N_6635,N_4950,N_4106);
nand U6636 (N_6636,N_3586,N_3884);
nor U6637 (N_6637,N_4520,N_5993);
and U6638 (N_6638,N_4289,N_3294);
nor U6639 (N_6639,N_5159,N_5973);
nor U6640 (N_6640,N_5889,N_5691);
and U6641 (N_6641,N_5961,N_4513);
or U6642 (N_6642,N_4306,N_3249);
nand U6643 (N_6643,N_5185,N_5903);
nor U6644 (N_6644,N_4428,N_5747);
and U6645 (N_6645,N_4249,N_4912);
nand U6646 (N_6646,N_3410,N_4518);
and U6647 (N_6647,N_3041,N_3514);
nand U6648 (N_6648,N_3002,N_3119);
or U6649 (N_6649,N_5800,N_5155);
or U6650 (N_6650,N_3118,N_4482);
and U6651 (N_6651,N_4965,N_4100);
nor U6652 (N_6652,N_3490,N_4122);
nor U6653 (N_6653,N_4990,N_5341);
or U6654 (N_6654,N_4649,N_5056);
nand U6655 (N_6655,N_5333,N_3074);
nand U6656 (N_6656,N_3957,N_4777);
and U6657 (N_6657,N_3125,N_5551);
nand U6658 (N_6658,N_3127,N_5727);
or U6659 (N_6659,N_5701,N_5447);
xor U6660 (N_6660,N_4713,N_4612);
nand U6661 (N_6661,N_3177,N_3685);
nor U6662 (N_6662,N_3907,N_5033);
nor U6663 (N_6663,N_3654,N_4529);
or U6664 (N_6664,N_4358,N_3790);
or U6665 (N_6665,N_3115,N_5147);
or U6666 (N_6666,N_4837,N_5130);
nand U6667 (N_6667,N_3304,N_4970);
and U6668 (N_6668,N_5134,N_3429);
or U6669 (N_6669,N_3288,N_4261);
and U6670 (N_6670,N_3597,N_3541);
nor U6671 (N_6671,N_3800,N_3983);
or U6672 (N_6672,N_3160,N_5839);
or U6673 (N_6673,N_4604,N_5009);
or U6674 (N_6674,N_3421,N_5825);
nand U6675 (N_6675,N_5703,N_3700);
nor U6676 (N_6676,N_4145,N_4720);
nor U6677 (N_6677,N_5101,N_3852);
and U6678 (N_6678,N_5853,N_3407);
or U6679 (N_6679,N_3042,N_4594);
xor U6680 (N_6680,N_5391,N_3670);
or U6681 (N_6681,N_3693,N_5176);
or U6682 (N_6682,N_4721,N_3269);
and U6683 (N_6683,N_5949,N_4390);
nand U6684 (N_6684,N_5951,N_4208);
nor U6685 (N_6685,N_3240,N_3529);
nand U6686 (N_6686,N_5759,N_3095);
nand U6687 (N_6687,N_3282,N_3938);
and U6688 (N_6688,N_3017,N_3264);
nand U6689 (N_6689,N_4167,N_3953);
nand U6690 (N_6690,N_3566,N_3088);
nand U6691 (N_6691,N_4888,N_5062);
nor U6692 (N_6692,N_3291,N_3747);
and U6693 (N_6693,N_5330,N_4173);
and U6694 (N_6694,N_3250,N_3252);
nor U6695 (N_6695,N_3312,N_5531);
and U6696 (N_6696,N_3795,N_4260);
and U6697 (N_6697,N_4637,N_5474);
and U6698 (N_6698,N_4979,N_5767);
nand U6699 (N_6699,N_4694,N_4465);
nand U6700 (N_6700,N_4067,N_5477);
or U6701 (N_6701,N_3167,N_5823);
or U6702 (N_6702,N_5501,N_3947);
and U6703 (N_6703,N_3990,N_5634);
or U6704 (N_6704,N_3533,N_3434);
nor U6705 (N_6705,N_5123,N_5718);
or U6706 (N_6706,N_4642,N_4275);
nor U6707 (N_6707,N_5677,N_3620);
or U6708 (N_6708,N_4850,N_5395);
or U6709 (N_6709,N_4292,N_5205);
or U6710 (N_6710,N_3215,N_4883);
and U6711 (N_6711,N_5516,N_4398);
or U6712 (N_6712,N_4869,N_4557);
nor U6713 (N_6713,N_3161,N_5417);
and U6714 (N_6714,N_4857,N_4985);
or U6715 (N_6715,N_3377,N_4916);
and U6716 (N_6716,N_4542,N_5871);
nand U6717 (N_6717,N_4790,N_3640);
and U6718 (N_6718,N_3448,N_3753);
or U6719 (N_6719,N_5805,N_4621);
nand U6720 (N_6720,N_3505,N_3341);
and U6721 (N_6721,N_3973,N_3016);
nor U6722 (N_6722,N_5347,N_5383);
nand U6723 (N_6723,N_3494,N_3825);
nor U6724 (N_6724,N_5614,N_5264);
or U6725 (N_6725,N_5714,N_4601);
nand U6726 (N_6726,N_5901,N_4307);
or U6727 (N_6727,N_4031,N_5567);
and U6728 (N_6728,N_5143,N_5301);
nor U6729 (N_6729,N_4247,N_5100);
or U6730 (N_6730,N_5882,N_5947);
xor U6731 (N_6731,N_4823,N_3225);
and U6732 (N_6732,N_5780,N_5907);
or U6733 (N_6733,N_5649,N_5287);
or U6734 (N_6734,N_5695,N_4343);
nand U6735 (N_6735,N_5692,N_5140);
and U6736 (N_6736,N_4239,N_5086);
nor U6737 (N_6737,N_5988,N_4223);
xor U6738 (N_6738,N_4523,N_4533);
nand U6739 (N_6739,N_3281,N_4267);
nand U6740 (N_6740,N_4409,N_5616);
nand U6741 (N_6741,N_4659,N_3608);
or U6742 (N_6742,N_3475,N_4592);
or U6743 (N_6743,N_4108,N_4939);
nand U6744 (N_6744,N_5554,N_5290);
nor U6745 (N_6745,N_5562,N_5018);
or U6746 (N_6746,N_3571,N_3314);
and U6747 (N_6747,N_3067,N_5112);
and U6748 (N_6748,N_5122,N_4907);
or U6749 (N_6749,N_3141,N_5010);
nor U6750 (N_6750,N_4088,N_5864);
or U6751 (N_6751,N_3963,N_3193);
or U6752 (N_6752,N_4931,N_3139);
nor U6753 (N_6753,N_4545,N_3123);
or U6754 (N_6754,N_5956,N_4102);
nor U6755 (N_6755,N_5059,N_5027);
or U6756 (N_6756,N_4860,N_4896);
nand U6757 (N_6757,N_3912,N_5965);
nand U6758 (N_6758,N_5227,N_5509);
or U6759 (N_6759,N_4270,N_5089);
or U6760 (N_6760,N_3279,N_3085);
nor U6761 (N_6761,N_5575,N_5279);
or U6762 (N_6762,N_5334,N_5755);
and U6763 (N_6763,N_3449,N_3910);
or U6764 (N_6764,N_3372,N_4125);
nand U6765 (N_6765,N_3099,N_4047);
or U6766 (N_6766,N_3465,N_5789);
or U6767 (N_6767,N_5558,N_4652);
and U6768 (N_6768,N_4765,N_4109);
nor U6769 (N_6769,N_3557,N_3113);
nor U6770 (N_6770,N_5569,N_3420);
or U6771 (N_6771,N_4858,N_5672);
nand U6772 (N_6772,N_4914,N_3258);
nor U6773 (N_6773,N_3474,N_4271);
or U6774 (N_6774,N_3941,N_3550);
nand U6775 (N_6775,N_5941,N_4450);
or U6776 (N_6776,N_3789,N_3675);
or U6777 (N_6777,N_3305,N_3565);
nor U6778 (N_6778,N_5687,N_3246);
nor U6779 (N_6779,N_4951,N_5361);
nand U6780 (N_6780,N_4243,N_3902);
and U6781 (N_6781,N_4629,N_4994);
nor U6782 (N_6782,N_4737,N_4000);
and U6783 (N_6783,N_4277,N_3522);
nor U6784 (N_6784,N_4492,N_3242);
or U6785 (N_6785,N_4323,N_5738);
nor U6786 (N_6786,N_4728,N_3664);
nor U6787 (N_6787,N_3261,N_3406);
and U6788 (N_6788,N_3891,N_3786);
nor U6789 (N_6789,N_5184,N_4490);
nor U6790 (N_6790,N_4396,N_5748);
and U6791 (N_6791,N_3657,N_4253);
nand U6792 (N_6792,N_3922,N_3585);
xnor U6793 (N_6793,N_4044,N_4595);
nor U6794 (N_6794,N_4953,N_3323);
or U6795 (N_6795,N_5092,N_5620);
nor U6796 (N_6796,N_3914,N_4090);
nand U6797 (N_6797,N_5404,N_3890);
and U6798 (N_6798,N_5791,N_5977);
and U6799 (N_6799,N_5282,N_5261);
and U6800 (N_6800,N_4057,N_4781);
nand U6801 (N_6801,N_4766,N_5872);
nor U6802 (N_6802,N_5411,N_4258);
and U6803 (N_6803,N_3727,N_5399);
or U6804 (N_6804,N_4664,N_3255);
nor U6805 (N_6805,N_3898,N_4327);
or U6806 (N_6806,N_5472,N_3340);
and U6807 (N_6807,N_3371,N_3435);
and U6808 (N_6808,N_3075,N_4477);
nand U6809 (N_6809,N_4722,N_5630);
nand U6810 (N_6810,N_4479,N_3386);
nor U6811 (N_6811,N_4330,N_4196);
and U6812 (N_6812,N_5845,N_3229);
and U6813 (N_6813,N_5657,N_5061);
or U6814 (N_6814,N_3969,N_3184);
nor U6815 (N_6815,N_3389,N_3418);
or U6816 (N_6816,N_4369,N_5127);
and U6817 (N_6817,N_5710,N_3741);
and U6818 (N_6818,N_4880,N_5717);
or U6819 (N_6819,N_5711,N_3687);
or U6820 (N_6820,N_4190,N_4911);
nor U6821 (N_6821,N_4809,N_4597);
or U6822 (N_6822,N_4891,N_5485);
nor U6823 (N_6823,N_4900,N_3916);
or U6824 (N_6824,N_4333,N_4876);
and U6825 (N_6825,N_5356,N_4153);
or U6826 (N_6826,N_5486,N_5915);
nand U6827 (N_6827,N_4796,N_3944);
or U6828 (N_6828,N_4727,N_5197);
nand U6829 (N_6829,N_5867,N_5025);
or U6830 (N_6830,N_4691,N_5420);
nor U6831 (N_6831,N_5432,N_4510);
xor U6832 (N_6832,N_5000,N_5129);
or U6833 (N_6833,N_4667,N_4027);
or U6834 (N_6834,N_4255,N_5875);
nand U6835 (N_6835,N_3760,N_5487);
or U6836 (N_6836,N_3121,N_5796);
nand U6837 (N_6837,N_3702,N_5105);
or U6838 (N_6838,N_5515,N_3564);
or U6839 (N_6839,N_4974,N_5693);
nand U6840 (N_6840,N_3209,N_4509);
and U6841 (N_6841,N_4577,N_3415);
nand U6842 (N_6842,N_4734,N_5042);
nor U6843 (N_6843,N_3289,N_4964);
nand U6844 (N_6844,N_4252,N_3995);
or U6845 (N_6845,N_3982,N_5351);
and U6846 (N_6846,N_3452,N_4360);
nor U6847 (N_6847,N_4661,N_5713);
nor U6848 (N_6848,N_5637,N_3024);
or U6849 (N_6849,N_5690,N_5212);
nand U6850 (N_6850,N_5204,N_5136);
nor U6851 (N_6851,N_4785,N_3886);
nor U6852 (N_6852,N_5640,N_5108);
or U6853 (N_6853,N_3582,N_4861);
or U6854 (N_6854,N_5802,N_3485);
nand U6855 (N_6855,N_4738,N_5643);
nor U6856 (N_6856,N_3171,N_4158);
nor U6857 (N_6857,N_4936,N_3663);
nor U6858 (N_6858,N_4603,N_5878);
and U6859 (N_6859,N_3919,N_5586);
or U6860 (N_6860,N_5080,N_4194);
and U6861 (N_6861,N_3738,N_3182);
nand U6862 (N_6862,N_5732,N_3804);
or U6863 (N_6863,N_3200,N_4839);
nand U6864 (N_6864,N_5684,N_4403);
nand U6865 (N_6865,N_3208,N_4115);
and U6866 (N_6866,N_4143,N_4787);
nor U6867 (N_6867,N_3843,N_3292);
nor U6868 (N_6868,N_5208,N_3276);
nand U6869 (N_6869,N_5834,N_5161);
and U6870 (N_6870,N_5887,N_5707);
nor U6871 (N_6871,N_3178,N_5958);
or U6872 (N_6872,N_5070,N_4530);
or U6873 (N_6873,N_4268,N_3915);
or U6874 (N_6874,N_4235,N_3965);
nand U6875 (N_6875,N_4123,N_4300);
and U6876 (N_6876,N_4822,N_4617);
or U6877 (N_6877,N_3345,N_4430);
nor U6878 (N_6878,N_5352,N_4166);
and U6879 (N_6879,N_4198,N_4726);
nor U6880 (N_6880,N_3909,N_3619);
nor U6881 (N_6881,N_3470,N_3899);
or U6882 (N_6882,N_4845,N_5740);
and U6883 (N_6883,N_5138,N_4609);
and U6884 (N_6884,N_5667,N_5076);
nor U6885 (N_6885,N_5481,N_4805);
nor U6886 (N_6886,N_4133,N_5996);
nor U6887 (N_6887,N_5392,N_5049);
or U6888 (N_6888,N_5698,N_5639);
or U6889 (N_6889,N_5480,N_5031);
nand U6890 (N_6890,N_4811,N_3714);
and U6891 (N_6891,N_4989,N_5442);
nand U6892 (N_6892,N_3019,N_3316);
nand U6893 (N_6893,N_5428,N_3451);
nand U6894 (N_6894,N_3330,N_4074);
and U6895 (N_6895,N_4634,N_3799);
nand U6896 (N_6896,N_3336,N_5600);
or U6897 (N_6897,N_5320,N_4759);
or U6898 (N_6898,N_3690,N_3730);
and U6899 (N_6899,N_3706,N_3669);
nand U6900 (N_6900,N_4946,N_4028);
nand U6901 (N_6901,N_4338,N_3105);
nor U6902 (N_6902,N_4426,N_4224);
or U6903 (N_6903,N_3528,N_4093);
nor U6904 (N_6904,N_3144,N_5920);
nor U6905 (N_6905,N_3581,N_4042);
nor U6906 (N_6906,N_3648,N_4018);
nor U6907 (N_6907,N_4847,N_3836);
or U6908 (N_6908,N_3440,N_3956);
and U6909 (N_6909,N_5441,N_4269);
nand U6910 (N_6910,N_4567,N_3633);
and U6911 (N_6911,N_4392,N_3084);
nor U6912 (N_6912,N_3194,N_3721);
and U6913 (N_6913,N_3616,N_3467);
nor U6914 (N_6914,N_3387,N_4843);
nor U6915 (N_6915,N_5438,N_3618);
nor U6916 (N_6916,N_5504,N_4474);
xnor U6917 (N_6917,N_3327,N_4256);
or U6918 (N_6918,N_3887,N_3574);
or U6919 (N_6919,N_5708,N_3347);
nor U6920 (N_6920,N_4910,N_4274);
nand U6921 (N_6921,N_3015,N_3562);
and U6922 (N_6922,N_3390,N_5343);
or U6923 (N_6923,N_5991,N_4186);
or U6924 (N_6924,N_5331,N_3329);
or U6925 (N_6925,N_5731,N_5196);
or U6926 (N_6926,N_3652,N_5291);
nand U6927 (N_6927,N_4942,N_5589);
nor U6928 (N_6928,N_3971,N_3360);
or U6929 (N_6929,N_4960,N_5978);
and U6930 (N_6930,N_5862,N_3376);
nor U6931 (N_6931,N_3020,N_5460);
and U6932 (N_6932,N_5217,N_4359);
or U6933 (N_6933,N_5267,N_4151);
nor U6934 (N_6934,N_5240,N_3726);
nand U6935 (N_6935,N_5886,N_3939);
nor U6936 (N_6936,N_3450,N_4786);
or U6937 (N_6937,N_3223,N_4813);
and U6938 (N_6938,N_4308,N_4310);
nand U6939 (N_6939,N_4588,N_4404);
or U6940 (N_6940,N_4600,N_5237);
nand U6941 (N_6941,N_5739,N_5673);
and U6942 (N_6942,N_5248,N_4614);
or U6943 (N_6943,N_5165,N_4863);
and U6944 (N_6944,N_3885,N_3538);
or U6945 (N_6945,N_5522,N_5914);
and U6946 (N_6946,N_4923,N_3595);
nor U6947 (N_6947,N_3081,N_3863);
nor U6948 (N_6948,N_5752,N_4052);
or U6949 (N_6949,N_4032,N_3607);
and U6950 (N_6950,N_4455,N_4206);
and U6951 (N_6951,N_3426,N_5319);
and U6952 (N_6952,N_4769,N_3293);
and U6953 (N_6953,N_4242,N_3943);
nor U6954 (N_6954,N_5762,N_4304);
and U6955 (N_6955,N_3163,N_3838);
nor U6956 (N_6956,N_3335,N_5294);
nor U6957 (N_6957,N_5982,N_4655);
nand U6958 (N_6958,N_3617,N_3297);
nand U6959 (N_6959,N_5415,N_3632);
and U6960 (N_6960,N_5478,N_4221);
nor U6961 (N_6961,N_4816,N_3066);
nand U6962 (N_6962,N_5346,N_4315);
or U6963 (N_6963,N_4584,N_5199);
or U6964 (N_6964,N_5792,N_5344);
xor U6965 (N_6965,N_5868,N_4554);
and U6966 (N_6966,N_5942,N_5401);
nor U6967 (N_6967,N_4384,N_5048);
or U6968 (N_6968,N_4624,N_4140);
nor U6969 (N_6969,N_3749,N_4820);
or U6970 (N_6970,N_5856,N_4201);
and U6971 (N_6971,N_5660,N_5952);
and U6972 (N_6972,N_5040,N_4118);
nor U6973 (N_6973,N_3542,N_3134);
or U6974 (N_6974,N_4397,N_4091);
nand U6975 (N_6975,N_5979,N_3011);
and U6976 (N_6976,N_3671,N_4467);
nand U6977 (N_6977,N_3353,N_3515);
and U6978 (N_6978,N_5234,N_4772);
nand U6979 (N_6979,N_3056,N_4709);
and U6980 (N_6980,N_4618,N_5450);
or U6981 (N_6981,N_5897,N_3030);
and U6982 (N_6982,N_5757,N_3488);
nand U6983 (N_6983,N_4319,N_5795);
or U6984 (N_6984,N_5446,N_3521);
and U6985 (N_6985,N_4116,N_3331);
nor U6986 (N_6986,N_4248,N_5339);
or U6987 (N_6987,N_4366,N_5744);
and U6988 (N_6988,N_5126,N_3712);
nor U6989 (N_6989,N_5271,N_5377);
nor U6990 (N_6990,N_4978,N_3720);
or U6991 (N_6991,N_3567,N_3109);
or U6992 (N_6992,N_4716,N_3445);
and U6993 (N_6993,N_5300,N_3477);
or U6994 (N_6994,N_3979,N_5001);
or U6995 (N_6995,N_3818,N_4625);
or U6996 (N_6996,N_5378,N_5663);
and U6997 (N_6997,N_5468,N_3554);
nand U6998 (N_6998,N_5519,N_4543);
nand U6999 (N_6999,N_5722,N_4024);
nor U7000 (N_7000,N_4480,N_4354);
or U7001 (N_7001,N_3822,N_5809);
and U7002 (N_7002,N_5484,N_5500);
nor U7003 (N_7003,N_3149,N_3428);
or U7004 (N_7004,N_5582,N_3021);
and U7005 (N_7005,N_3900,N_4279);
and U7006 (N_7006,N_5398,N_3839);
and U7007 (N_7007,N_3116,N_5712);
nand U7008 (N_7008,N_5683,N_4213);
nor U7009 (N_7009,N_3351,N_5641);
or U7010 (N_7010,N_4996,N_4852);
nand U7011 (N_7011,N_3352,N_4932);
nand U7012 (N_7012,N_3073,N_4356);
and U7013 (N_7013,N_4017,N_3785);
or U7014 (N_7014,N_3405,N_5544);
nor U7015 (N_7015,N_4676,N_3678);
or U7016 (N_7016,N_5021,N_4240);
nor U7017 (N_7017,N_4808,N_3471);
nor U7018 (N_7018,N_4148,N_3765);
nand U7019 (N_7019,N_3960,N_3639);
or U7020 (N_7020,N_5454,N_4113);
or U7021 (N_7021,N_4408,N_5625);
and U7022 (N_7022,N_5648,N_3925);
or U7023 (N_7023,N_5222,N_5104);
nor U7024 (N_7024,N_5142,N_3740);
nor U7025 (N_7025,N_3043,N_3729);
nand U7026 (N_7026,N_3395,N_4280);
nand U7027 (N_7027,N_4293,N_4393);
nor U7028 (N_7028,N_3364,N_4884);
nand U7029 (N_7029,N_4081,N_5646);
and U7030 (N_7030,N_3463,N_3453);
nand U7031 (N_7031,N_3556,N_5583);
and U7032 (N_7032,N_4747,N_5364);
or U7033 (N_7033,N_3888,N_3408);
nand U7034 (N_7034,N_5079,N_5229);
or U7035 (N_7035,N_4739,N_5716);
or U7036 (N_7036,N_5855,N_5131);
nand U7037 (N_7037,N_3896,N_5604);
nand U7038 (N_7038,N_4745,N_3339);
nand U7039 (N_7039,N_5661,N_5609);
nor U7040 (N_7040,N_3151,N_3211);
or U7041 (N_7041,N_3413,N_3400);
or U7042 (N_7042,N_3715,N_4666);
nand U7043 (N_7043,N_3964,N_3854);
and U7044 (N_7044,N_5192,N_3373);
and U7045 (N_7045,N_5194,N_5819);
nor U7046 (N_7046,N_4362,N_3219);
nor U7047 (N_7047,N_3037,N_4491);
or U7048 (N_7048,N_4080,N_4344);
nand U7049 (N_7049,N_3401,N_5488);
and U7050 (N_7050,N_4962,N_4531);
and U7051 (N_7051,N_4129,N_5847);
nor U7052 (N_7052,N_3461,N_4440);
or U7053 (N_7053,N_5342,N_5203);
nand U7054 (N_7054,N_4063,N_4583);
or U7055 (N_7055,N_4175,N_3842);
nor U7056 (N_7056,N_4053,N_4710);
nor U7057 (N_7057,N_4638,N_3154);
nor U7058 (N_7058,N_4656,N_5458);
nor U7059 (N_7059,N_3643,N_5524);
or U7060 (N_7060,N_5371,N_5644);
nor U7061 (N_7061,N_5627,N_3383);
nand U7062 (N_7062,N_5742,N_4436);
nand U7063 (N_7063,N_4622,N_3711);
and U7064 (N_7064,N_3908,N_3409);
and U7065 (N_7065,N_5962,N_3610);
or U7066 (N_7066,N_5963,N_4128);
and U7067 (N_7067,N_5617,N_3082);
and U7068 (N_7068,N_5560,N_5268);
and U7069 (N_7069,N_3235,N_3862);
nand U7070 (N_7070,N_4141,N_3858);
or U7071 (N_7071,N_3321,N_3948);
and U7072 (N_7072,N_4420,N_4011);
or U7073 (N_7073,N_5694,N_3905);
nor U7074 (N_7074,N_3646,N_3079);
and U7075 (N_7075,N_5241,N_3499);
and U7076 (N_7076,N_3188,N_4009);
and U7077 (N_7077,N_3233,N_5382);
and U7078 (N_7078,N_5729,N_3623);
nand U7079 (N_7079,N_5306,N_4494);
nor U7080 (N_7080,N_3544,N_3277);
nor U7081 (N_7081,N_3055,N_5157);
and U7082 (N_7082,N_5186,N_3054);
nand U7083 (N_7083,N_4476,N_5983);
or U7084 (N_7084,N_4800,N_3503);
nor U7085 (N_7085,N_3828,N_3273);
or U7086 (N_7086,N_3388,N_3097);
nor U7087 (N_7087,N_4783,N_5270);
nand U7088 (N_7088,N_3224,N_5216);
nand U7089 (N_7089,N_3398,N_4961);
or U7090 (N_7090,N_4591,N_3536);
nor U7091 (N_7091,N_5167,N_5456);
nand U7092 (N_7092,N_3555,N_3342);
nor U7093 (N_7093,N_5784,N_5975);
nand U7094 (N_7094,N_3736,N_4705);
nor U7095 (N_7095,N_4982,N_4927);
or U7096 (N_7096,N_3495,N_4332);
nand U7097 (N_7097,N_3776,N_5366);
and U7098 (N_7098,N_4631,N_5182);
nor U7099 (N_7099,N_4537,N_4746);
and U7100 (N_7100,N_4030,N_3710);
xor U7101 (N_7101,N_3165,N_5540);
or U7102 (N_7102,N_4755,N_3961);
nand U7103 (N_7103,N_3045,N_5224);
and U7104 (N_7104,N_5619,N_3397);
and U7105 (N_7105,N_4688,N_4736);
nand U7106 (N_7106,N_5272,N_3614);
or U7107 (N_7107,N_5328,N_5898);
or U7108 (N_7108,N_5075,N_5510);
xnor U7109 (N_7109,N_5355,N_4458);
and U7110 (N_7110,N_3976,N_5367);
nor U7111 (N_7111,N_3114,N_3370);
nor U7112 (N_7112,N_3365,N_4640);
or U7113 (N_7113,N_5052,N_5599);
or U7114 (N_7114,N_4371,N_4668);
or U7115 (N_7115,N_4773,N_3810);
nand U7116 (N_7116,N_3059,N_5723);
nand U7117 (N_7117,N_4421,N_4842);
and U7118 (N_7118,N_4237,N_5421);
or U7119 (N_7119,N_3346,N_5927);
and U7120 (N_7120,N_5304,N_4680);
or U7121 (N_7121,N_5071,N_5245);
nor U7122 (N_7122,N_5408,N_4412);
or U7123 (N_7123,N_4244,N_5682);
nand U7124 (N_7124,N_4471,N_3636);
or U7125 (N_7125,N_4220,N_3146);
or U7126 (N_7126,N_4464,N_4003);
nor U7127 (N_7127,N_5133,N_4895);
and U7128 (N_7128,N_3553,N_5624);
and U7129 (N_7129,N_4563,N_4590);
or U7130 (N_7130,N_4815,N_5664);
or U7131 (N_7131,N_3873,N_3315);
or U7132 (N_7132,N_3798,N_5322);
or U7133 (N_7133,N_4035,N_4460);
or U7134 (N_7134,N_5297,N_3480);
nand U7135 (N_7135,N_3817,N_4539);
nand U7136 (N_7136,N_5045,N_5935);
nor U7137 (N_7137,N_4473,N_4049);
nor U7138 (N_7138,N_3205,N_3695);
or U7139 (N_7139,N_4751,N_3260);
or U7140 (N_7140,N_3414,N_3057);
and U7141 (N_7141,N_5443,N_3750);
or U7142 (N_7142,N_4241,N_4483);
or U7143 (N_7143,N_5671,N_3231);
nor U7144 (N_7144,N_3904,N_4082);
nand U7145 (N_7145,N_4712,N_5709);
and U7146 (N_7146,N_5020,N_3379);
and U7147 (N_7147,N_4947,N_4683);
and U7148 (N_7148,N_3975,N_3525);
nor U7149 (N_7149,N_5870,N_3197);
nor U7150 (N_7150,N_4342,N_5303);
or U7151 (N_7151,N_5545,N_5906);
and U7152 (N_7152,N_5636,N_4435);
and U7153 (N_7153,N_4986,N_4633);
and U7154 (N_7154,N_5292,N_5231);
or U7155 (N_7155,N_3759,N_4486);
nand U7156 (N_7156,N_4349,N_4699);
and U7157 (N_7157,N_4449,N_3083);
nand U7158 (N_7158,N_4760,N_3875);
nor U7159 (N_7159,N_4188,N_5174);
nand U7160 (N_7160,N_5464,N_5473);
and U7161 (N_7161,N_5511,N_3189);
nor U7162 (N_7162,N_5223,N_4670);
nor U7163 (N_7163,N_3009,N_4835);
nor U7164 (N_7164,N_5934,N_5099);
nand U7165 (N_7165,N_5832,N_5373);
nand U7166 (N_7166,N_5429,N_4616);
nand U7167 (N_7167,N_3871,N_4101);
nor U7168 (N_7168,N_5170,N_3436);
and U7169 (N_7169,N_5836,N_5402);
nand U7170 (N_7170,N_3940,N_3307);
nand U7171 (N_7171,N_5525,N_5106);
or U7172 (N_7172,N_3569,N_4071);
or U7173 (N_7173,N_3861,N_3676);
xnor U7174 (N_7174,N_3913,N_3748);
or U7175 (N_7175,N_5793,N_3204);
nand U7176 (N_7176,N_4920,N_5463);
or U7177 (N_7177,N_5116,N_4048);
and U7178 (N_7178,N_5735,N_3369);
or U7179 (N_7179,N_4399,N_5006);
and U7180 (N_7180,N_4935,N_4519);
or U7181 (N_7181,N_4377,N_4892);
nand U7182 (N_7182,N_3725,N_3318);
and U7183 (N_7183,N_4422,N_4160);
and U7184 (N_7184,N_5699,N_3124);
or U7185 (N_7185,N_4489,N_4452);
or U7186 (N_7186,N_5824,N_5427);
or U7187 (N_7187,N_3518,N_3432);
nor U7188 (N_7188,N_3267,N_5178);
nand U7189 (N_7189,N_5283,N_4415);
and U7190 (N_7190,N_4368,N_4485);
or U7191 (N_7191,N_3901,N_3592);
nor U7192 (N_7192,N_4320,N_3666);
or U7193 (N_7193,N_3705,N_4112);
nand U7194 (N_7194,N_5146,N_3959);
or U7195 (N_7195,N_3757,N_4992);
and U7196 (N_7196,N_4099,N_5955);
or U7197 (N_7197,N_3609,N_3847);
and U7198 (N_7198,N_5003,N_5419);
nand U7199 (N_7199,N_3110,N_5705);
or U7200 (N_7200,N_5721,N_4038);
nand U7201 (N_7201,N_3923,N_3935);
nor U7202 (N_7202,N_4854,N_4084);
or U7203 (N_7203,N_5019,N_5390);
xnor U7204 (N_7204,N_5806,N_4219);
or U7205 (N_7205,N_5838,N_5932);
nand U7206 (N_7206,N_5494,N_3023);
nand U7207 (N_7207,N_4077,N_5275);
and U7208 (N_7208,N_4069,N_5153);
nand U7209 (N_7209,N_4386,N_3779);
and U7210 (N_7210,N_3001,N_5036);
nand U7211 (N_7211,N_5312,N_5265);
and U7212 (N_7212,N_3446,N_4575);
and U7213 (N_7213,N_4461,N_5848);
nand U7214 (N_7214,N_4501,N_5563);
nor U7215 (N_7215,N_3644,N_5596);
or U7216 (N_7216,N_5608,N_3106);
or U7217 (N_7217,N_3844,N_5754);
and U7218 (N_7218,N_3133,N_5533);
and U7219 (N_7219,N_4364,N_4060);
nand U7220 (N_7220,N_3874,N_3591);
and U7221 (N_7221,N_5091,N_5405);
and U7222 (N_7222,N_3823,N_5548);
nand U7223 (N_7223,N_4309,N_3459);
or U7224 (N_7224,N_4147,N_5250);
nor U7225 (N_7225,N_3534,N_3612);
and U7226 (N_7226,N_3442,N_3827);
nor U7227 (N_7227,N_4137,N_5788);
nor U7228 (N_7228,N_4124,N_3889);
nand U7229 (N_7229,N_3458,N_5972);
or U7230 (N_7230,N_3214,N_3047);
nand U7231 (N_7231,N_4919,N_5011);
and U7232 (N_7232,N_4646,N_4171);
nand U7233 (N_7233,N_3684,N_3107);
nor U7234 (N_7234,N_4214,N_4999);
nor U7235 (N_7235,N_3326,N_4948);
nand U7236 (N_7236,N_4997,N_4587);
nor U7237 (N_7237,N_5187,N_3337);
nand U7238 (N_7238,N_5790,N_4427);
nor U7239 (N_7239,N_3756,N_3357);
or U7240 (N_7240,N_4607,N_4372);
or U7241 (N_7241,N_4043,N_5686);
or U7242 (N_7242,N_3656,N_4406);
nand U7243 (N_7243,N_4528,N_3022);
and U7244 (N_7244,N_3433,N_4572);
or U7245 (N_7245,N_5842,N_4301);
or U7246 (N_7246,N_3295,N_5288);
nand U7247 (N_7247,N_5168,N_3210);
and U7248 (N_7248,N_3207,N_5883);
nand U7249 (N_7249,N_3040,N_5931);
and U7250 (N_7250,N_5659,N_5219);
or U7251 (N_7251,N_3897,N_5044);
nor U7252 (N_7252,N_4503,N_4744);
xor U7253 (N_7253,N_5213,N_4635);
or U7254 (N_7254,N_5779,N_5523);
or U7255 (N_7255,N_5120,N_5110);
nand U7256 (N_7256,N_4917,N_4207);
and U7257 (N_7257,N_5822,N_3764);
nor U7258 (N_7258,N_5414,N_4684);
nand U7259 (N_7259,N_5255,N_5831);
nor U7260 (N_7260,N_3548,N_3857);
nor U7261 (N_7261,N_5936,N_5093);
nand U7262 (N_7262,N_3653,N_4586);
nand U7263 (N_7263,N_5613,N_4352);
and U7264 (N_7264,N_3128,N_5506);
nor U7265 (N_7265,N_4454,N_4593);
nand U7266 (N_7266,N_4189,N_5030);
and U7267 (N_7267,N_4894,N_4383);
or U7268 (N_7268,N_4924,N_4346);
nand U7269 (N_7269,N_5359,N_5113);
and U7270 (N_7270,N_5622,N_5851);
or U7271 (N_7271,N_3077,N_4740);
nand U7272 (N_7272,N_5166,N_5926);
nor U7273 (N_7273,N_3655,N_3238);
nand U7274 (N_7274,N_3568,N_5349);
and U7275 (N_7275,N_5704,N_4419);
nand U7276 (N_7276,N_3508,N_5615);
or U7277 (N_7277,N_3809,N_5315);
nor U7278 (N_7278,N_5424,N_4904);
nand U7279 (N_7279,N_3540,N_4898);
and U7280 (N_7280,N_4702,N_4499);
nor U7281 (N_7281,N_4040,N_3168);
or U7282 (N_7282,N_4387,N_3641);
nand U7283 (N_7283,N_4180,N_4086);
nand U7284 (N_7284,N_3829,N_5536);
nand U7285 (N_7285,N_5866,N_5026);
nor U7286 (N_7286,N_5638,N_5969);
or U7287 (N_7287,N_5403,N_5179);
nor U7288 (N_7288,N_3173,N_5348);
nand U7289 (N_7289,N_4782,N_5154);
or U7290 (N_7290,N_3894,N_4335);
nand U7291 (N_7291,N_3306,N_3046);
or U7292 (N_7292,N_5877,N_4628);
nand U7293 (N_7293,N_3932,N_3758);
or U7294 (N_7294,N_5353,N_3117);
and U7295 (N_7295,N_5688,N_5384);
nor U7296 (N_7296,N_5549,N_5430);
or U7297 (N_7297,N_5783,N_4266);
nor U7298 (N_7298,N_5337,N_5258);
nor U7299 (N_7299,N_4185,N_4886);
nand U7300 (N_7300,N_3784,N_3848);
nand U7301 (N_7301,N_3577,N_3126);
xnor U7302 (N_7302,N_3539,N_4834);
nor U7303 (N_7303,N_4311,N_4675);
nand U7304 (N_7304,N_4127,N_5269);
nor U7305 (N_7305,N_3164,N_3972);
and U7306 (N_7306,N_3230,N_3625);
nor U7307 (N_7307,N_5674,N_3774);
nand U7308 (N_7308,N_5310,N_5114);
or U7309 (N_7309,N_3437,N_4231);
nor U7310 (N_7310,N_4540,N_4534);
and U7311 (N_7311,N_3849,N_3482);
and U7312 (N_7312,N_4958,N_5801);
nand U7313 (N_7313,N_4423,N_3497);
nand U7314 (N_7314,N_4840,N_3545);
nor U7315 (N_7315,N_3150,N_5768);
nand U7316 (N_7316,N_4981,N_5368);
nor U7317 (N_7317,N_3744,N_3131);
or U7318 (N_7318,N_5658,N_3945);
or U7319 (N_7319,N_5808,N_5681);
or U7320 (N_7320,N_3977,N_4468);
or U7321 (N_7321,N_4438,N_5909);
and U7322 (N_7322,N_5587,N_3328);
or U7323 (N_7323,N_5452,N_5465);
nand U7324 (N_7324,N_4754,N_4456);
or U7325 (N_7325,N_3050,N_5892);
nand U7326 (N_7326,N_4623,N_5513);
and U7327 (N_7327,N_4763,N_5814);
and U7328 (N_7328,N_4110,N_5552);
and U7329 (N_7329,N_4325,N_5259);
nand U7330 (N_7330,N_3992,N_4302);
and U7331 (N_7331,N_5172,N_3427);
nand U7332 (N_7332,N_4742,N_3966);
or U7333 (N_7333,N_4937,N_4305);
and U7334 (N_7334,N_4901,N_4169);
and U7335 (N_7335,N_4550,N_3812);
nand U7336 (N_7336,N_3153,N_5736);
nand U7337 (N_7337,N_4446,N_3006);
nand U7338 (N_7338,N_3660,N_5200);
nand U7339 (N_7339,N_3613,N_5413);
nand U7340 (N_7340,N_4197,N_3527);
or U7341 (N_7341,N_3254,N_5004);
and U7342 (N_7342,N_4677,N_4181);
nand U7343 (N_7343,N_5607,N_5125);
nor U7344 (N_7344,N_4527,N_5012);
nand U7345 (N_7345,N_4903,N_4495);
nor U7346 (N_7346,N_3980,N_4696);
and U7347 (N_7347,N_4678,N_4749);
xnor U7348 (N_7348,N_5491,N_4576);
and U7349 (N_7349,N_4701,N_4085);
xnor U7350 (N_7350,N_5102,N_3012);
nand U7351 (N_7351,N_4162,N_3588);
nand U7352 (N_7352,N_4926,N_4263);
and U7353 (N_7353,N_5107,N_4831);
nand U7354 (N_7354,N_5069,N_3013);
and U7355 (N_7355,N_5406,N_5363);
nand U7356 (N_7356,N_4157,N_4889);
nand U7357 (N_7357,N_4810,N_3354);
nor U7358 (N_7358,N_4959,N_4564);
and U7359 (N_7359,N_5097,N_4743);
or U7360 (N_7360,N_5751,N_4879);
and U7361 (N_7361,N_4250,N_5535);
and U7362 (N_7362,N_4807,N_3181);
nand U7363 (N_7363,N_3094,N_4723);
nor U7364 (N_7364,N_5623,N_4021);
or U7365 (N_7365,N_5593,N_3380);
and U7366 (N_7366,N_3507,N_5023);
and U7367 (N_7367,N_5354,N_5057);
nor U7368 (N_7368,N_5396,N_5980);
nor U7369 (N_7369,N_3062,N_4665);
and U7370 (N_7370,N_4172,N_4013);
or U7371 (N_7371,N_4672,N_4357);
or U7372 (N_7372,N_3698,N_3108);
or U7373 (N_7373,N_4347,N_5517);
nor U7374 (N_7374,N_4512,N_3719);
nand U7375 (N_7375,N_3044,N_4980);
nand U7376 (N_7376,N_4630,N_3317);
nand U7377 (N_7377,N_4159,N_5769);
or U7378 (N_7378,N_3679,N_3811);
nand U7379 (N_7379,N_4650,N_4192);
nor U7380 (N_7380,N_4400,N_3344);
nor U7381 (N_7381,N_3599,N_3129);
nor U7382 (N_7382,N_3707,N_4036);
and U7383 (N_7383,N_4750,N_4913);
or U7384 (N_7384,N_5526,N_5055);
or U7385 (N_7385,N_4956,N_3140);
nand U7386 (N_7386,N_5016,N_3792);
nand U7387 (N_7387,N_3573,N_4803);
or U7388 (N_7388,N_5111,N_4690);
nand U7389 (N_7389,N_3302,N_5281);
and U7390 (N_7390,N_3921,N_3325);
nand U7391 (N_7391,N_4966,N_5652);
nand U7392 (N_7392,N_3174,N_4657);
nand U7393 (N_7393,N_4484,N_3218);
and U7394 (N_7394,N_3366,N_5280);
nor U7395 (N_7395,N_5804,N_3247);
or U7396 (N_7396,N_3755,N_3195);
nor U7397 (N_7397,N_4168,N_3145);
and U7398 (N_7398,N_5945,N_3598);
nor U7399 (N_7399,N_3763,N_4975);
and U7400 (N_7400,N_4257,N_4211);
or U7401 (N_7401,N_5852,N_5841);
or U7402 (N_7402,N_4987,N_4295);
nor U7403 (N_7403,N_5476,N_5541);
or U7404 (N_7404,N_4988,N_5242);
and U7405 (N_7405,N_3378,N_5495);
or U7406 (N_7406,N_4693,N_3651);
nand U7407 (N_7407,N_3877,N_3665);
or U7408 (N_7408,N_3156,N_5385);
nand U7409 (N_7409,N_5253,N_5813);
nand U7410 (N_7410,N_5944,N_4363);
nand U7411 (N_7411,N_4524,N_5152);
or U7412 (N_7412,N_5299,N_5943);
and U7413 (N_7413,N_5210,N_4218);
or U7414 (N_7414,N_4234,N_3275);
or U7415 (N_7415,N_3793,N_5565);
nand U7416 (N_7416,N_5556,N_3137);
or U7417 (N_7417,N_4264,N_5512);
and U7418 (N_7418,N_4909,N_3191);
or U7419 (N_7419,N_4799,N_3703);
nand U7420 (N_7420,N_3356,N_4284);
or U7421 (N_7421,N_5765,N_4574);
nor U7422 (N_7422,N_3185,N_4433);
and U7423 (N_7423,N_4868,N_4104);
nor U7424 (N_7424,N_5043,N_4170);
nor U7425 (N_7425,N_5647,N_4873);
or U7426 (N_7426,N_5585,N_4671);
nand U7427 (N_7427,N_5555,N_4708);
xnor U7428 (N_7428,N_3080,N_4849);
nor U7429 (N_7429,N_4378,N_5675);
or U7430 (N_7430,N_3035,N_4983);
or U7431 (N_7431,N_3924,N_5700);
nand U7432 (N_7432,N_5181,N_5580);
or U7433 (N_7433,N_4217,N_4949);
or U7434 (N_7434,N_4410,N_4015);
and U7435 (N_7435,N_3739,N_4789);
and U7436 (N_7436,N_5734,N_4405);
or U7437 (N_7437,N_5939,N_3221);
and U7438 (N_7438,N_3699,N_4544);
or U7439 (N_7439,N_3251,N_3692);
nor U7440 (N_7440,N_3355,N_3278);
and U7441 (N_7441,N_4826,N_5050);
nand U7442 (N_7442,N_5706,N_3148);
and U7443 (N_7443,N_5828,N_3688);
nor U7444 (N_7444,N_3391,N_5689);
and U7445 (N_7445,N_3778,N_4012);
nand U7446 (N_7446,N_3310,N_5144);
nor U7447 (N_7447,N_4643,N_4824);
nand U7448 (N_7448,N_3590,N_4619);
and U7449 (N_7449,N_4336,N_3147);
and U7450 (N_7450,N_4434,N_5068);
xor U7451 (N_7451,N_5423,N_3516);
or U7452 (N_7452,N_3232,N_5063);
nor U7453 (N_7453,N_4443,N_5311);
and U7454 (N_7454,N_4969,N_3228);
nor U7455 (N_7455,N_4848,N_3243);
nand U7456 (N_7456,N_4866,N_4299);
or U7457 (N_7457,N_5195,N_3322);
and U7458 (N_7458,N_4451,N_3697);
or U7459 (N_7459,N_5278,N_5532);
nor U7460 (N_7460,N_4669,N_4187);
or U7461 (N_7461,N_3834,N_4089);
or U7462 (N_7462,N_4565,N_3468);
nand U7463 (N_7463,N_5365,N_3272);
nand U7464 (N_7464,N_3993,N_4411);
or U7465 (N_7465,N_5289,N_4209);
or U7466 (N_7466,N_5606,N_5547);
nor U7467 (N_7467,N_5974,N_4717);
and U7468 (N_7468,N_5141,N_4136);
nand U7469 (N_7469,N_3460,N_3190);
nand U7470 (N_7470,N_5350,N_4193);
or U7471 (N_7471,N_3384,N_3876);
nor U7472 (N_7472,N_5145,N_3052);
nand U7473 (N_7473,N_3911,N_3761);
nand U7474 (N_7474,N_4046,N_3833);
or U7475 (N_7475,N_3403,N_5444);
nand U7476 (N_7476,N_4639,N_3234);
nand U7477 (N_7477,N_5821,N_4014);
and U7478 (N_7478,N_3523,N_4317);
and U7479 (N_7479,N_4775,N_4025);
xnor U7480 (N_7480,N_3443,N_3576);
or U7481 (N_7481,N_3735,N_3111);
or U7482 (N_7482,N_4328,N_3952);
nor U7483 (N_7483,N_5846,N_3991);
and U7484 (N_7484,N_5534,N_3422);
or U7485 (N_7485,N_5527,N_5492);
and U7486 (N_7486,N_4814,N_5081);
and U7487 (N_7487,N_3667,N_5249);
or U7488 (N_7488,N_4862,N_4470);
nor U7489 (N_7489,N_3265,N_5968);
nor U7490 (N_7490,N_4164,N_3270);
nor U7491 (N_7491,N_4205,N_4830);
nor U7492 (N_7492,N_3053,N_5360);
nand U7493 (N_7493,N_4768,N_3457);
or U7494 (N_7494,N_3394,N_4353);
nor U7495 (N_7495,N_4921,N_4867);
and U7496 (N_7496,N_4050,N_3382);
nand U7497 (N_7497,N_3070,N_3256);
nand U7498 (N_7498,N_5899,N_5827);
nand U7499 (N_7499,N_3986,N_4957);
nand U7500 (N_7500,N_5856,N_4450);
nor U7501 (N_7501,N_5468,N_3565);
nor U7502 (N_7502,N_5633,N_5005);
and U7503 (N_7503,N_3958,N_5351);
or U7504 (N_7504,N_5757,N_4126);
nor U7505 (N_7505,N_4983,N_4763);
and U7506 (N_7506,N_5790,N_5242);
nand U7507 (N_7507,N_5955,N_3072);
or U7508 (N_7508,N_5168,N_4947);
nand U7509 (N_7509,N_4108,N_5189);
nand U7510 (N_7510,N_5323,N_4532);
nand U7511 (N_7511,N_5592,N_3333);
or U7512 (N_7512,N_4455,N_4648);
or U7513 (N_7513,N_3278,N_5807);
and U7514 (N_7514,N_5838,N_5449);
and U7515 (N_7515,N_5026,N_5024);
or U7516 (N_7516,N_5417,N_3792);
and U7517 (N_7517,N_3515,N_5585);
or U7518 (N_7518,N_4554,N_4238);
or U7519 (N_7519,N_5738,N_5743);
or U7520 (N_7520,N_3054,N_4228);
nand U7521 (N_7521,N_5835,N_5789);
nor U7522 (N_7522,N_3256,N_5309);
nor U7523 (N_7523,N_4845,N_4811);
and U7524 (N_7524,N_5756,N_4239);
and U7525 (N_7525,N_3203,N_5215);
nor U7526 (N_7526,N_3347,N_3683);
or U7527 (N_7527,N_4253,N_4980);
and U7528 (N_7528,N_5975,N_5643);
nor U7529 (N_7529,N_4612,N_5589);
nor U7530 (N_7530,N_3562,N_5446);
nor U7531 (N_7531,N_5173,N_5805);
and U7532 (N_7532,N_5247,N_3723);
nand U7533 (N_7533,N_3808,N_4257);
nand U7534 (N_7534,N_3812,N_5828);
nor U7535 (N_7535,N_3391,N_4443);
and U7536 (N_7536,N_5322,N_4484);
nand U7537 (N_7537,N_5862,N_4935);
nor U7538 (N_7538,N_4828,N_4491);
and U7539 (N_7539,N_3294,N_5179);
and U7540 (N_7540,N_3259,N_5561);
nor U7541 (N_7541,N_3097,N_4971);
or U7542 (N_7542,N_4680,N_4530);
or U7543 (N_7543,N_5635,N_3116);
and U7544 (N_7544,N_5671,N_3204);
nand U7545 (N_7545,N_4874,N_5383);
or U7546 (N_7546,N_4934,N_5866);
or U7547 (N_7547,N_3020,N_3805);
and U7548 (N_7548,N_3280,N_5018);
nor U7549 (N_7549,N_3237,N_3431);
and U7550 (N_7550,N_3109,N_4495);
xnor U7551 (N_7551,N_3441,N_5580);
nor U7552 (N_7552,N_5192,N_3857);
or U7553 (N_7553,N_3094,N_3764);
and U7554 (N_7554,N_3081,N_3524);
and U7555 (N_7555,N_5739,N_4160);
nand U7556 (N_7556,N_5099,N_3126);
nor U7557 (N_7557,N_3660,N_5683);
nand U7558 (N_7558,N_5066,N_3947);
or U7559 (N_7559,N_3843,N_4389);
and U7560 (N_7560,N_3851,N_4482);
nand U7561 (N_7561,N_5468,N_4492);
nand U7562 (N_7562,N_5725,N_4577);
nand U7563 (N_7563,N_4174,N_5855);
or U7564 (N_7564,N_5687,N_3974);
nand U7565 (N_7565,N_4364,N_5891);
or U7566 (N_7566,N_4456,N_3689);
and U7567 (N_7567,N_5764,N_3533);
nand U7568 (N_7568,N_5685,N_3044);
nor U7569 (N_7569,N_5801,N_5298);
and U7570 (N_7570,N_5844,N_4989);
or U7571 (N_7571,N_5660,N_3847);
and U7572 (N_7572,N_5220,N_4343);
or U7573 (N_7573,N_5480,N_4589);
and U7574 (N_7574,N_4125,N_4131);
nand U7575 (N_7575,N_3991,N_4640);
and U7576 (N_7576,N_5612,N_4593);
or U7577 (N_7577,N_5449,N_4343);
or U7578 (N_7578,N_5371,N_4718);
nor U7579 (N_7579,N_4776,N_4700);
nor U7580 (N_7580,N_3461,N_3559);
and U7581 (N_7581,N_5528,N_3743);
or U7582 (N_7582,N_4362,N_5439);
nor U7583 (N_7583,N_4320,N_5196);
nor U7584 (N_7584,N_4354,N_4837);
nand U7585 (N_7585,N_3626,N_4510);
nand U7586 (N_7586,N_5492,N_4805);
nand U7587 (N_7587,N_3540,N_5445);
and U7588 (N_7588,N_5518,N_5958);
nor U7589 (N_7589,N_4848,N_5531);
nor U7590 (N_7590,N_4275,N_4188);
nand U7591 (N_7591,N_3854,N_5702);
nor U7592 (N_7592,N_3867,N_4464);
nor U7593 (N_7593,N_3331,N_4598);
nand U7594 (N_7594,N_3917,N_5187);
nand U7595 (N_7595,N_4236,N_3314);
nor U7596 (N_7596,N_5217,N_3756);
nand U7597 (N_7597,N_5596,N_5857);
or U7598 (N_7598,N_3876,N_4801);
nand U7599 (N_7599,N_4080,N_3212);
nor U7600 (N_7600,N_5778,N_3836);
and U7601 (N_7601,N_3300,N_5496);
nor U7602 (N_7602,N_4250,N_4127);
and U7603 (N_7603,N_4855,N_5974);
nand U7604 (N_7604,N_4852,N_4058);
and U7605 (N_7605,N_4701,N_3602);
nor U7606 (N_7606,N_5206,N_4750);
nand U7607 (N_7607,N_4678,N_3499);
and U7608 (N_7608,N_5611,N_4660);
or U7609 (N_7609,N_4116,N_4529);
nor U7610 (N_7610,N_3721,N_3521);
and U7611 (N_7611,N_3815,N_5508);
nor U7612 (N_7612,N_4868,N_4600);
and U7613 (N_7613,N_5803,N_5438);
or U7614 (N_7614,N_4781,N_3426);
nand U7615 (N_7615,N_3285,N_5395);
and U7616 (N_7616,N_5330,N_3166);
or U7617 (N_7617,N_5541,N_4797);
nand U7618 (N_7618,N_3959,N_4755);
nand U7619 (N_7619,N_5934,N_3313);
xor U7620 (N_7620,N_4534,N_5344);
or U7621 (N_7621,N_4987,N_3408);
nor U7622 (N_7622,N_5156,N_5675);
xor U7623 (N_7623,N_4825,N_3408);
nor U7624 (N_7624,N_3853,N_4116);
nor U7625 (N_7625,N_5674,N_3739);
and U7626 (N_7626,N_5208,N_5323);
and U7627 (N_7627,N_4587,N_4435);
and U7628 (N_7628,N_3769,N_3586);
nand U7629 (N_7629,N_4557,N_4636);
nand U7630 (N_7630,N_5924,N_5619);
or U7631 (N_7631,N_5825,N_5536);
nor U7632 (N_7632,N_3132,N_5104);
nand U7633 (N_7633,N_5441,N_4752);
or U7634 (N_7634,N_3391,N_5642);
or U7635 (N_7635,N_3311,N_5764);
nand U7636 (N_7636,N_4768,N_4790);
and U7637 (N_7637,N_4443,N_5551);
and U7638 (N_7638,N_4770,N_3482);
nand U7639 (N_7639,N_3648,N_4057);
nand U7640 (N_7640,N_5770,N_3824);
nor U7641 (N_7641,N_4043,N_4523);
or U7642 (N_7642,N_5079,N_5408);
and U7643 (N_7643,N_3830,N_4091);
nor U7644 (N_7644,N_5349,N_5259);
nor U7645 (N_7645,N_5046,N_4460);
and U7646 (N_7646,N_3262,N_3038);
and U7647 (N_7647,N_3596,N_4076);
and U7648 (N_7648,N_4774,N_3369);
nor U7649 (N_7649,N_4407,N_5043);
and U7650 (N_7650,N_4646,N_4308);
nand U7651 (N_7651,N_3024,N_3631);
and U7652 (N_7652,N_5253,N_5031);
nand U7653 (N_7653,N_4430,N_3997);
nand U7654 (N_7654,N_3324,N_5919);
and U7655 (N_7655,N_5082,N_3827);
or U7656 (N_7656,N_3391,N_3492);
or U7657 (N_7657,N_4660,N_4027);
nor U7658 (N_7658,N_5851,N_4942);
nand U7659 (N_7659,N_5083,N_5369);
nand U7660 (N_7660,N_4522,N_3842);
nand U7661 (N_7661,N_3816,N_5740);
nand U7662 (N_7662,N_3651,N_4951);
xnor U7663 (N_7663,N_5598,N_4208);
nor U7664 (N_7664,N_4285,N_3074);
or U7665 (N_7665,N_3359,N_5615);
and U7666 (N_7666,N_3953,N_4648);
and U7667 (N_7667,N_4965,N_4015);
or U7668 (N_7668,N_4083,N_5527);
nor U7669 (N_7669,N_5840,N_5081);
or U7670 (N_7670,N_3475,N_5647);
or U7671 (N_7671,N_5721,N_4864);
and U7672 (N_7672,N_5234,N_5031);
and U7673 (N_7673,N_4807,N_5149);
nand U7674 (N_7674,N_5965,N_4201);
nor U7675 (N_7675,N_4014,N_4575);
and U7676 (N_7676,N_3111,N_4983);
xnor U7677 (N_7677,N_5318,N_4793);
and U7678 (N_7678,N_5532,N_4590);
nand U7679 (N_7679,N_3928,N_5921);
nor U7680 (N_7680,N_3219,N_4081);
nand U7681 (N_7681,N_5688,N_4747);
nand U7682 (N_7682,N_5643,N_3305);
nand U7683 (N_7683,N_3309,N_3454);
or U7684 (N_7684,N_4076,N_4520);
or U7685 (N_7685,N_5923,N_3766);
or U7686 (N_7686,N_4717,N_3187);
nor U7687 (N_7687,N_3033,N_5893);
and U7688 (N_7688,N_4392,N_5698);
or U7689 (N_7689,N_3103,N_5499);
or U7690 (N_7690,N_4984,N_5324);
and U7691 (N_7691,N_5359,N_4489);
nand U7692 (N_7692,N_5024,N_4181);
or U7693 (N_7693,N_5310,N_5925);
nor U7694 (N_7694,N_4790,N_3885);
nor U7695 (N_7695,N_3730,N_4735);
or U7696 (N_7696,N_5687,N_3608);
and U7697 (N_7697,N_4170,N_4650);
nand U7698 (N_7698,N_5968,N_3458);
nor U7699 (N_7699,N_3113,N_4470);
nand U7700 (N_7700,N_4712,N_4891);
nand U7701 (N_7701,N_4260,N_5091);
or U7702 (N_7702,N_3261,N_4415);
nand U7703 (N_7703,N_3334,N_3350);
nand U7704 (N_7704,N_4420,N_4631);
nand U7705 (N_7705,N_3866,N_3066);
nand U7706 (N_7706,N_4552,N_4963);
nand U7707 (N_7707,N_3967,N_3175);
or U7708 (N_7708,N_5774,N_3528);
nand U7709 (N_7709,N_3171,N_5662);
nor U7710 (N_7710,N_5220,N_4492);
nor U7711 (N_7711,N_4989,N_4777);
nand U7712 (N_7712,N_3680,N_3085);
and U7713 (N_7713,N_3598,N_3346);
and U7714 (N_7714,N_3158,N_3052);
nor U7715 (N_7715,N_4784,N_5731);
and U7716 (N_7716,N_4519,N_3451);
or U7717 (N_7717,N_3217,N_4601);
and U7718 (N_7718,N_3819,N_3967);
or U7719 (N_7719,N_5287,N_5405);
nand U7720 (N_7720,N_4083,N_4435);
and U7721 (N_7721,N_5796,N_3085);
nor U7722 (N_7722,N_3750,N_3063);
and U7723 (N_7723,N_5505,N_3132);
nor U7724 (N_7724,N_4124,N_5577);
or U7725 (N_7725,N_5195,N_3985);
or U7726 (N_7726,N_4588,N_4538);
or U7727 (N_7727,N_3199,N_5880);
and U7728 (N_7728,N_4507,N_5270);
nor U7729 (N_7729,N_4029,N_5581);
and U7730 (N_7730,N_4059,N_4485);
or U7731 (N_7731,N_5739,N_4761);
or U7732 (N_7732,N_3970,N_5291);
or U7733 (N_7733,N_5810,N_4356);
nand U7734 (N_7734,N_4730,N_5582);
nand U7735 (N_7735,N_5056,N_4713);
and U7736 (N_7736,N_4890,N_3237);
nand U7737 (N_7737,N_3248,N_5701);
nand U7738 (N_7738,N_5107,N_4489);
nor U7739 (N_7739,N_5496,N_4793);
or U7740 (N_7740,N_3844,N_3200);
or U7741 (N_7741,N_3988,N_5602);
nand U7742 (N_7742,N_4828,N_5730);
nor U7743 (N_7743,N_3538,N_4936);
nand U7744 (N_7744,N_4301,N_5099);
and U7745 (N_7745,N_4486,N_4540);
nor U7746 (N_7746,N_5912,N_3728);
nor U7747 (N_7747,N_5350,N_4417);
and U7748 (N_7748,N_5814,N_5064);
nand U7749 (N_7749,N_4743,N_4255);
nand U7750 (N_7750,N_4339,N_5506);
nor U7751 (N_7751,N_3841,N_4334);
and U7752 (N_7752,N_5085,N_4727);
nor U7753 (N_7753,N_3589,N_5061);
nor U7754 (N_7754,N_4485,N_3623);
or U7755 (N_7755,N_5225,N_5320);
nand U7756 (N_7756,N_4437,N_4348);
nor U7757 (N_7757,N_4318,N_5449);
nor U7758 (N_7758,N_3794,N_3862);
nand U7759 (N_7759,N_5632,N_5195);
or U7760 (N_7760,N_4241,N_5186);
nor U7761 (N_7761,N_4642,N_3372);
nand U7762 (N_7762,N_5277,N_3360);
or U7763 (N_7763,N_3881,N_3120);
nand U7764 (N_7764,N_5702,N_4988);
xor U7765 (N_7765,N_4414,N_5051);
or U7766 (N_7766,N_5340,N_4061);
or U7767 (N_7767,N_4465,N_3403);
and U7768 (N_7768,N_4547,N_4627);
nand U7769 (N_7769,N_4656,N_3432);
nor U7770 (N_7770,N_3359,N_5873);
nor U7771 (N_7771,N_3605,N_3363);
nor U7772 (N_7772,N_4176,N_5585);
xor U7773 (N_7773,N_3487,N_5355);
and U7774 (N_7774,N_3069,N_4485);
nor U7775 (N_7775,N_5365,N_3019);
nor U7776 (N_7776,N_5828,N_5415);
or U7777 (N_7777,N_4736,N_5026);
or U7778 (N_7778,N_5386,N_5883);
nand U7779 (N_7779,N_3645,N_5023);
or U7780 (N_7780,N_5869,N_3922);
and U7781 (N_7781,N_5360,N_3758);
nand U7782 (N_7782,N_5615,N_3491);
or U7783 (N_7783,N_5288,N_3469);
nor U7784 (N_7784,N_4604,N_4750);
or U7785 (N_7785,N_4210,N_3863);
nor U7786 (N_7786,N_5391,N_5050);
nor U7787 (N_7787,N_4592,N_4729);
and U7788 (N_7788,N_3438,N_4221);
nor U7789 (N_7789,N_3750,N_5857);
nand U7790 (N_7790,N_4778,N_5252);
or U7791 (N_7791,N_5835,N_3147);
or U7792 (N_7792,N_4065,N_5380);
and U7793 (N_7793,N_4261,N_4400);
nand U7794 (N_7794,N_5745,N_4793);
nand U7795 (N_7795,N_3005,N_5615);
or U7796 (N_7796,N_3753,N_3714);
nor U7797 (N_7797,N_3722,N_4865);
or U7798 (N_7798,N_3692,N_5470);
and U7799 (N_7799,N_5242,N_4479);
nand U7800 (N_7800,N_3658,N_3621);
nor U7801 (N_7801,N_4947,N_3933);
nand U7802 (N_7802,N_5986,N_5843);
nor U7803 (N_7803,N_5757,N_4025);
or U7804 (N_7804,N_3956,N_3066);
and U7805 (N_7805,N_5532,N_3378);
xnor U7806 (N_7806,N_5785,N_4864);
nor U7807 (N_7807,N_3030,N_4250);
or U7808 (N_7808,N_5842,N_3170);
nor U7809 (N_7809,N_5409,N_3377);
nor U7810 (N_7810,N_5369,N_4192);
and U7811 (N_7811,N_3653,N_3442);
and U7812 (N_7812,N_3368,N_4619);
or U7813 (N_7813,N_3410,N_3095);
nand U7814 (N_7814,N_3665,N_3486);
nor U7815 (N_7815,N_5997,N_5370);
or U7816 (N_7816,N_5409,N_3083);
nand U7817 (N_7817,N_4226,N_5449);
or U7818 (N_7818,N_4840,N_5067);
nor U7819 (N_7819,N_3881,N_5950);
and U7820 (N_7820,N_3907,N_3011);
nand U7821 (N_7821,N_3512,N_3092);
nor U7822 (N_7822,N_4455,N_5833);
nor U7823 (N_7823,N_4012,N_4543);
nor U7824 (N_7824,N_4662,N_5706);
nand U7825 (N_7825,N_3028,N_5039);
nor U7826 (N_7826,N_3008,N_5237);
nand U7827 (N_7827,N_4287,N_5733);
and U7828 (N_7828,N_5457,N_5949);
nor U7829 (N_7829,N_3654,N_5071);
and U7830 (N_7830,N_5822,N_4289);
nor U7831 (N_7831,N_5491,N_5051);
nand U7832 (N_7832,N_5819,N_4330);
nand U7833 (N_7833,N_5684,N_3235);
nand U7834 (N_7834,N_4727,N_4947);
nand U7835 (N_7835,N_3500,N_5623);
and U7836 (N_7836,N_4671,N_4003);
nand U7837 (N_7837,N_4762,N_3884);
nor U7838 (N_7838,N_5835,N_5729);
and U7839 (N_7839,N_4627,N_5159);
nand U7840 (N_7840,N_5502,N_5777);
nand U7841 (N_7841,N_5908,N_5738);
nor U7842 (N_7842,N_5184,N_4250);
nor U7843 (N_7843,N_4495,N_4107);
and U7844 (N_7844,N_4410,N_4541);
nor U7845 (N_7845,N_5139,N_3842);
nor U7846 (N_7846,N_3347,N_4508);
and U7847 (N_7847,N_4620,N_4178);
nand U7848 (N_7848,N_5340,N_5831);
nand U7849 (N_7849,N_3018,N_3290);
nor U7850 (N_7850,N_5394,N_5408);
xnor U7851 (N_7851,N_4016,N_4526);
nor U7852 (N_7852,N_3667,N_3145);
nand U7853 (N_7853,N_5703,N_5603);
nor U7854 (N_7854,N_4354,N_3673);
or U7855 (N_7855,N_4470,N_3943);
and U7856 (N_7856,N_5955,N_4688);
and U7857 (N_7857,N_5591,N_3925);
and U7858 (N_7858,N_4710,N_5578);
nand U7859 (N_7859,N_3182,N_3258);
or U7860 (N_7860,N_5452,N_3702);
nor U7861 (N_7861,N_3590,N_4369);
or U7862 (N_7862,N_5368,N_4180);
and U7863 (N_7863,N_5348,N_4878);
or U7864 (N_7864,N_4261,N_5339);
or U7865 (N_7865,N_4500,N_4355);
or U7866 (N_7866,N_4483,N_4377);
and U7867 (N_7867,N_3203,N_4245);
nor U7868 (N_7868,N_5103,N_3817);
nor U7869 (N_7869,N_5014,N_4570);
nor U7870 (N_7870,N_4117,N_4916);
or U7871 (N_7871,N_3773,N_3896);
or U7872 (N_7872,N_5777,N_3958);
or U7873 (N_7873,N_5056,N_3584);
or U7874 (N_7874,N_5533,N_3213);
or U7875 (N_7875,N_3977,N_5411);
nor U7876 (N_7876,N_5901,N_3604);
nand U7877 (N_7877,N_3285,N_4060);
nor U7878 (N_7878,N_4321,N_4934);
or U7879 (N_7879,N_5459,N_5250);
or U7880 (N_7880,N_3965,N_3326);
nor U7881 (N_7881,N_4025,N_4741);
or U7882 (N_7882,N_4650,N_4437);
and U7883 (N_7883,N_4189,N_5676);
or U7884 (N_7884,N_4120,N_5917);
and U7885 (N_7885,N_4577,N_3969);
nand U7886 (N_7886,N_5313,N_5121);
nor U7887 (N_7887,N_5671,N_3308);
nand U7888 (N_7888,N_3462,N_5438);
or U7889 (N_7889,N_5476,N_4866);
and U7890 (N_7890,N_5010,N_4155);
and U7891 (N_7891,N_3405,N_5421);
nor U7892 (N_7892,N_4559,N_4062);
or U7893 (N_7893,N_4672,N_3149);
or U7894 (N_7894,N_5132,N_4156);
xnor U7895 (N_7895,N_5520,N_3959);
nand U7896 (N_7896,N_4962,N_3998);
and U7897 (N_7897,N_4186,N_5277);
nand U7898 (N_7898,N_5487,N_4949);
and U7899 (N_7899,N_4447,N_5769);
nor U7900 (N_7900,N_3948,N_3345);
or U7901 (N_7901,N_5636,N_4139);
nor U7902 (N_7902,N_3802,N_5359);
or U7903 (N_7903,N_4714,N_4938);
nor U7904 (N_7904,N_3446,N_5972);
or U7905 (N_7905,N_3346,N_4679);
nand U7906 (N_7906,N_4328,N_3638);
or U7907 (N_7907,N_5265,N_5486);
or U7908 (N_7908,N_4465,N_3825);
and U7909 (N_7909,N_5026,N_5042);
or U7910 (N_7910,N_5734,N_4901);
nand U7911 (N_7911,N_3938,N_5761);
or U7912 (N_7912,N_3644,N_4965);
and U7913 (N_7913,N_5898,N_5382);
nand U7914 (N_7914,N_3416,N_4915);
and U7915 (N_7915,N_4880,N_3067);
nor U7916 (N_7916,N_3357,N_4596);
and U7917 (N_7917,N_4479,N_5885);
and U7918 (N_7918,N_5551,N_4125);
nand U7919 (N_7919,N_3741,N_3048);
nor U7920 (N_7920,N_4865,N_5469);
or U7921 (N_7921,N_5947,N_3396);
xor U7922 (N_7922,N_3773,N_4980);
and U7923 (N_7923,N_3790,N_3073);
xnor U7924 (N_7924,N_5176,N_5733);
or U7925 (N_7925,N_4231,N_5200);
or U7926 (N_7926,N_5985,N_4266);
or U7927 (N_7927,N_5076,N_4436);
or U7928 (N_7928,N_4140,N_4778);
nand U7929 (N_7929,N_3259,N_5574);
or U7930 (N_7930,N_5466,N_4546);
nand U7931 (N_7931,N_4857,N_3967);
or U7932 (N_7932,N_4014,N_4294);
or U7933 (N_7933,N_3967,N_4965);
nand U7934 (N_7934,N_3172,N_5038);
nand U7935 (N_7935,N_3001,N_3372);
and U7936 (N_7936,N_3546,N_5487);
and U7937 (N_7937,N_4237,N_4937);
or U7938 (N_7938,N_3161,N_4117);
and U7939 (N_7939,N_4712,N_3481);
and U7940 (N_7940,N_4118,N_3673);
or U7941 (N_7941,N_3459,N_3243);
and U7942 (N_7942,N_4534,N_4343);
or U7943 (N_7943,N_3634,N_5168);
nor U7944 (N_7944,N_3833,N_4711);
and U7945 (N_7945,N_4110,N_4127);
nor U7946 (N_7946,N_4864,N_3128);
and U7947 (N_7947,N_5710,N_5939);
nand U7948 (N_7948,N_4981,N_5674);
nand U7949 (N_7949,N_3281,N_5882);
nand U7950 (N_7950,N_3631,N_3904);
nor U7951 (N_7951,N_5682,N_5890);
nor U7952 (N_7952,N_3848,N_3891);
and U7953 (N_7953,N_4537,N_5040);
and U7954 (N_7954,N_3403,N_5439);
nor U7955 (N_7955,N_5751,N_5430);
or U7956 (N_7956,N_4282,N_4377);
and U7957 (N_7957,N_5228,N_3408);
or U7958 (N_7958,N_3508,N_4046);
nand U7959 (N_7959,N_4622,N_5045);
nor U7960 (N_7960,N_5453,N_4076);
or U7961 (N_7961,N_5918,N_4832);
and U7962 (N_7962,N_3081,N_4857);
and U7963 (N_7963,N_3050,N_5235);
or U7964 (N_7964,N_5038,N_3619);
nand U7965 (N_7965,N_3954,N_4976);
or U7966 (N_7966,N_3672,N_4658);
nand U7967 (N_7967,N_4238,N_3882);
and U7968 (N_7968,N_5411,N_3998);
or U7969 (N_7969,N_4297,N_3113);
and U7970 (N_7970,N_5850,N_3825);
nor U7971 (N_7971,N_4659,N_5745);
nor U7972 (N_7972,N_5532,N_3028);
nand U7973 (N_7973,N_4053,N_3321);
or U7974 (N_7974,N_4673,N_5277);
nand U7975 (N_7975,N_4590,N_4520);
or U7976 (N_7976,N_3294,N_5379);
and U7977 (N_7977,N_3512,N_5571);
nor U7978 (N_7978,N_5674,N_3081);
and U7979 (N_7979,N_3221,N_5993);
nor U7980 (N_7980,N_3614,N_5829);
nor U7981 (N_7981,N_4320,N_5545);
or U7982 (N_7982,N_3561,N_4957);
or U7983 (N_7983,N_5749,N_4367);
nor U7984 (N_7984,N_4496,N_3837);
nand U7985 (N_7985,N_5167,N_4523);
nor U7986 (N_7986,N_5937,N_4156);
and U7987 (N_7987,N_3503,N_3043);
nor U7988 (N_7988,N_5264,N_4157);
nand U7989 (N_7989,N_5177,N_3364);
nand U7990 (N_7990,N_4200,N_5981);
or U7991 (N_7991,N_3723,N_5347);
and U7992 (N_7992,N_4465,N_5041);
or U7993 (N_7993,N_3324,N_3040);
nor U7994 (N_7994,N_5357,N_5980);
nor U7995 (N_7995,N_3072,N_3169);
nor U7996 (N_7996,N_3995,N_3957);
nor U7997 (N_7997,N_3876,N_4600);
nor U7998 (N_7998,N_5383,N_3721);
nand U7999 (N_7999,N_5319,N_3582);
or U8000 (N_8000,N_5918,N_4090);
nor U8001 (N_8001,N_3275,N_4262);
or U8002 (N_8002,N_4245,N_3387);
and U8003 (N_8003,N_3435,N_4357);
nor U8004 (N_8004,N_3962,N_3992);
or U8005 (N_8005,N_3193,N_5807);
or U8006 (N_8006,N_5823,N_3852);
and U8007 (N_8007,N_3771,N_4576);
or U8008 (N_8008,N_3172,N_3296);
and U8009 (N_8009,N_5428,N_3629);
and U8010 (N_8010,N_4051,N_4279);
and U8011 (N_8011,N_5212,N_4763);
nand U8012 (N_8012,N_3106,N_4953);
or U8013 (N_8013,N_5438,N_5406);
nor U8014 (N_8014,N_3191,N_5082);
nand U8015 (N_8015,N_5100,N_4139);
and U8016 (N_8016,N_3807,N_3938);
nor U8017 (N_8017,N_3831,N_3983);
and U8018 (N_8018,N_4801,N_3904);
nor U8019 (N_8019,N_3763,N_3448);
nor U8020 (N_8020,N_4451,N_3043);
nor U8021 (N_8021,N_4824,N_5199);
nor U8022 (N_8022,N_5833,N_5737);
and U8023 (N_8023,N_5723,N_4222);
nand U8024 (N_8024,N_5200,N_5531);
and U8025 (N_8025,N_4111,N_5190);
nor U8026 (N_8026,N_3611,N_3673);
or U8027 (N_8027,N_4272,N_4368);
and U8028 (N_8028,N_4384,N_5314);
nor U8029 (N_8029,N_5509,N_5146);
and U8030 (N_8030,N_5488,N_5933);
nor U8031 (N_8031,N_5327,N_5618);
and U8032 (N_8032,N_3671,N_5443);
nor U8033 (N_8033,N_5803,N_4478);
and U8034 (N_8034,N_5607,N_5286);
and U8035 (N_8035,N_5674,N_5531);
or U8036 (N_8036,N_4364,N_5967);
nand U8037 (N_8037,N_3364,N_3320);
and U8038 (N_8038,N_5838,N_3027);
nand U8039 (N_8039,N_3627,N_3201);
nor U8040 (N_8040,N_4233,N_4511);
and U8041 (N_8041,N_5074,N_4597);
nor U8042 (N_8042,N_3833,N_3270);
nor U8043 (N_8043,N_5756,N_3601);
and U8044 (N_8044,N_5192,N_3593);
nand U8045 (N_8045,N_3302,N_5845);
nor U8046 (N_8046,N_4477,N_3963);
and U8047 (N_8047,N_3714,N_3694);
or U8048 (N_8048,N_5373,N_4896);
or U8049 (N_8049,N_3939,N_5315);
nor U8050 (N_8050,N_5606,N_5347);
nor U8051 (N_8051,N_3591,N_3333);
or U8052 (N_8052,N_4298,N_4280);
nand U8053 (N_8053,N_5137,N_5085);
nor U8054 (N_8054,N_4379,N_5023);
nand U8055 (N_8055,N_5979,N_4185);
nor U8056 (N_8056,N_4969,N_3945);
or U8057 (N_8057,N_5210,N_3836);
nand U8058 (N_8058,N_3263,N_4367);
and U8059 (N_8059,N_4452,N_3801);
and U8060 (N_8060,N_3825,N_5223);
or U8061 (N_8061,N_5895,N_3282);
or U8062 (N_8062,N_3340,N_3136);
nand U8063 (N_8063,N_5539,N_4057);
nor U8064 (N_8064,N_3062,N_4399);
and U8065 (N_8065,N_3908,N_3345);
or U8066 (N_8066,N_3973,N_5276);
nor U8067 (N_8067,N_3579,N_5371);
nand U8068 (N_8068,N_4691,N_3247);
nor U8069 (N_8069,N_5862,N_4151);
nor U8070 (N_8070,N_3028,N_5569);
nor U8071 (N_8071,N_3223,N_3908);
and U8072 (N_8072,N_4988,N_5079);
nand U8073 (N_8073,N_4682,N_3663);
nor U8074 (N_8074,N_3448,N_4247);
or U8075 (N_8075,N_5343,N_4838);
and U8076 (N_8076,N_4182,N_4704);
and U8077 (N_8077,N_5787,N_3429);
nand U8078 (N_8078,N_3526,N_5546);
nand U8079 (N_8079,N_3130,N_4493);
or U8080 (N_8080,N_5757,N_3283);
or U8081 (N_8081,N_3097,N_3347);
nand U8082 (N_8082,N_5841,N_3818);
and U8083 (N_8083,N_5972,N_4296);
nor U8084 (N_8084,N_5327,N_4078);
and U8085 (N_8085,N_3458,N_5320);
or U8086 (N_8086,N_5631,N_5326);
nor U8087 (N_8087,N_3553,N_4287);
and U8088 (N_8088,N_5231,N_4250);
and U8089 (N_8089,N_5679,N_3079);
nand U8090 (N_8090,N_4109,N_3114);
and U8091 (N_8091,N_5366,N_5597);
nor U8092 (N_8092,N_3043,N_3733);
nand U8093 (N_8093,N_4785,N_3597);
and U8094 (N_8094,N_5643,N_3267);
and U8095 (N_8095,N_4514,N_3763);
nand U8096 (N_8096,N_4246,N_5662);
nor U8097 (N_8097,N_3967,N_4945);
and U8098 (N_8098,N_3460,N_3669);
or U8099 (N_8099,N_3547,N_3606);
nand U8100 (N_8100,N_4374,N_4504);
nor U8101 (N_8101,N_5475,N_5036);
nor U8102 (N_8102,N_4950,N_3868);
nor U8103 (N_8103,N_5497,N_3093);
nor U8104 (N_8104,N_5465,N_5558);
nor U8105 (N_8105,N_3771,N_4186);
nand U8106 (N_8106,N_3506,N_4744);
nor U8107 (N_8107,N_3170,N_4613);
nor U8108 (N_8108,N_3428,N_5341);
nand U8109 (N_8109,N_5381,N_5105);
and U8110 (N_8110,N_5186,N_4890);
or U8111 (N_8111,N_4232,N_5962);
and U8112 (N_8112,N_4486,N_3319);
or U8113 (N_8113,N_4113,N_3811);
nand U8114 (N_8114,N_3521,N_3709);
nor U8115 (N_8115,N_3252,N_5131);
nand U8116 (N_8116,N_4906,N_3430);
and U8117 (N_8117,N_4120,N_4567);
or U8118 (N_8118,N_3857,N_3250);
nand U8119 (N_8119,N_3227,N_3496);
or U8120 (N_8120,N_3580,N_3017);
and U8121 (N_8121,N_4426,N_4612);
or U8122 (N_8122,N_4693,N_4664);
and U8123 (N_8123,N_4752,N_5693);
nand U8124 (N_8124,N_5540,N_5110);
nand U8125 (N_8125,N_4659,N_4074);
nor U8126 (N_8126,N_4112,N_5256);
or U8127 (N_8127,N_5498,N_3931);
nand U8128 (N_8128,N_5267,N_4617);
or U8129 (N_8129,N_5821,N_4931);
or U8130 (N_8130,N_3890,N_5624);
nand U8131 (N_8131,N_4942,N_3452);
or U8132 (N_8132,N_4747,N_4254);
or U8133 (N_8133,N_4334,N_3183);
and U8134 (N_8134,N_3072,N_3069);
and U8135 (N_8135,N_5338,N_3779);
nor U8136 (N_8136,N_4742,N_5702);
xnor U8137 (N_8137,N_3289,N_3059);
nor U8138 (N_8138,N_4602,N_3685);
or U8139 (N_8139,N_3606,N_4946);
or U8140 (N_8140,N_5756,N_3611);
nor U8141 (N_8141,N_4913,N_5856);
nand U8142 (N_8142,N_5006,N_3042);
nor U8143 (N_8143,N_5491,N_3957);
xor U8144 (N_8144,N_5327,N_5573);
nor U8145 (N_8145,N_4296,N_5046);
nor U8146 (N_8146,N_3290,N_3780);
or U8147 (N_8147,N_5598,N_4835);
or U8148 (N_8148,N_5779,N_3675);
and U8149 (N_8149,N_5673,N_3596);
xnor U8150 (N_8150,N_5463,N_5125);
or U8151 (N_8151,N_3077,N_3217);
nor U8152 (N_8152,N_5527,N_5309);
nor U8153 (N_8153,N_3544,N_3171);
nand U8154 (N_8154,N_3829,N_3700);
or U8155 (N_8155,N_3674,N_4453);
nand U8156 (N_8156,N_4673,N_3922);
nand U8157 (N_8157,N_4982,N_3749);
nor U8158 (N_8158,N_3859,N_4557);
nand U8159 (N_8159,N_3028,N_5111);
and U8160 (N_8160,N_3748,N_5418);
nand U8161 (N_8161,N_5340,N_5287);
or U8162 (N_8162,N_4633,N_4125);
nor U8163 (N_8163,N_3263,N_3602);
nor U8164 (N_8164,N_4683,N_3051);
and U8165 (N_8165,N_4466,N_3018);
and U8166 (N_8166,N_3647,N_3343);
nand U8167 (N_8167,N_5751,N_4015);
or U8168 (N_8168,N_5551,N_3870);
or U8169 (N_8169,N_3292,N_3888);
or U8170 (N_8170,N_4082,N_3712);
nor U8171 (N_8171,N_3696,N_4385);
and U8172 (N_8172,N_4461,N_5999);
and U8173 (N_8173,N_4251,N_3395);
or U8174 (N_8174,N_4025,N_5457);
nand U8175 (N_8175,N_3517,N_3745);
or U8176 (N_8176,N_5742,N_5087);
or U8177 (N_8177,N_4344,N_4826);
or U8178 (N_8178,N_3384,N_3365);
or U8179 (N_8179,N_5972,N_3653);
nor U8180 (N_8180,N_3360,N_3656);
nor U8181 (N_8181,N_4391,N_3433);
nor U8182 (N_8182,N_3421,N_5637);
and U8183 (N_8183,N_4689,N_4351);
nor U8184 (N_8184,N_4709,N_5236);
or U8185 (N_8185,N_5017,N_4386);
nor U8186 (N_8186,N_3923,N_4549);
nand U8187 (N_8187,N_3025,N_5705);
nor U8188 (N_8188,N_4198,N_3068);
nand U8189 (N_8189,N_4152,N_4272);
or U8190 (N_8190,N_3439,N_5239);
nor U8191 (N_8191,N_5800,N_5215);
or U8192 (N_8192,N_3955,N_4062);
or U8193 (N_8193,N_3848,N_4828);
or U8194 (N_8194,N_5769,N_5267);
nand U8195 (N_8195,N_3631,N_5904);
nand U8196 (N_8196,N_4853,N_3459);
and U8197 (N_8197,N_4629,N_4957);
and U8198 (N_8198,N_5929,N_4189);
nand U8199 (N_8199,N_3413,N_3010);
nand U8200 (N_8200,N_4225,N_3478);
or U8201 (N_8201,N_3203,N_5753);
and U8202 (N_8202,N_3623,N_5353);
nor U8203 (N_8203,N_4552,N_3547);
and U8204 (N_8204,N_5616,N_3919);
or U8205 (N_8205,N_5423,N_4161);
or U8206 (N_8206,N_5633,N_5537);
nor U8207 (N_8207,N_4236,N_5495);
nand U8208 (N_8208,N_4521,N_3053);
nand U8209 (N_8209,N_3685,N_5625);
or U8210 (N_8210,N_3568,N_5674);
or U8211 (N_8211,N_4875,N_4445);
nand U8212 (N_8212,N_5234,N_5005);
or U8213 (N_8213,N_4260,N_3143);
nor U8214 (N_8214,N_4287,N_3576);
and U8215 (N_8215,N_5761,N_3657);
and U8216 (N_8216,N_4232,N_5927);
or U8217 (N_8217,N_3405,N_3214);
and U8218 (N_8218,N_5058,N_4947);
nand U8219 (N_8219,N_4483,N_5688);
nor U8220 (N_8220,N_3638,N_3326);
nand U8221 (N_8221,N_4081,N_3968);
nor U8222 (N_8222,N_4120,N_4384);
nor U8223 (N_8223,N_3538,N_4269);
or U8224 (N_8224,N_4677,N_4147);
nand U8225 (N_8225,N_5159,N_4633);
nor U8226 (N_8226,N_3436,N_5188);
and U8227 (N_8227,N_5689,N_4757);
and U8228 (N_8228,N_4159,N_3337);
or U8229 (N_8229,N_4892,N_5136);
or U8230 (N_8230,N_5394,N_4308);
and U8231 (N_8231,N_4847,N_4631);
and U8232 (N_8232,N_3913,N_4377);
nand U8233 (N_8233,N_5241,N_4190);
and U8234 (N_8234,N_3906,N_3352);
nor U8235 (N_8235,N_3840,N_5004);
and U8236 (N_8236,N_5757,N_5911);
nand U8237 (N_8237,N_4481,N_5141);
nand U8238 (N_8238,N_4306,N_4090);
nand U8239 (N_8239,N_5347,N_5279);
nand U8240 (N_8240,N_3498,N_4190);
and U8241 (N_8241,N_5348,N_5155);
and U8242 (N_8242,N_5140,N_5725);
nor U8243 (N_8243,N_4460,N_5585);
or U8244 (N_8244,N_3146,N_5488);
nand U8245 (N_8245,N_5503,N_5228);
nand U8246 (N_8246,N_4900,N_5446);
and U8247 (N_8247,N_3273,N_3972);
nor U8248 (N_8248,N_4224,N_4210);
or U8249 (N_8249,N_5912,N_3838);
nor U8250 (N_8250,N_3287,N_4211);
and U8251 (N_8251,N_4486,N_3420);
nand U8252 (N_8252,N_5244,N_5030);
nor U8253 (N_8253,N_5272,N_5220);
nand U8254 (N_8254,N_4162,N_4887);
and U8255 (N_8255,N_4445,N_4117);
or U8256 (N_8256,N_5146,N_3656);
and U8257 (N_8257,N_4187,N_5997);
nand U8258 (N_8258,N_5394,N_4241);
and U8259 (N_8259,N_3463,N_5192);
nor U8260 (N_8260,N_5404,N_5884);
nor U8261 (N_8261,N_3117,N_5674);
and U8262 (N_8262,N_5540,N_5957);
nor U8263 (N_8263,N_5522,N_4174);
and U8264 (N_8264,N_5128,N_4343);
nand U8265 (N_8265,N_3387,N_4354);
or U8266 (N_8266,N_4006,N_3609);
nand U8267 (N_8267,N_4511,N_4236);
and U8268 (N_8268,N_5227,N_4430);
and U8269 (N_8269,N_5429,N_4393);
nor U8270 (N_8270,N_5239,N_5943);
and U8271 (N_8271,N_3068,N_4716);
nor U8272 (N_8272,N_4318,N_5762);
nor U8273 (N_8273,N_5989,N_5067);
and U8274 (N_8274,N_3854,N_4667);
and U8275 (N_8275,N_4452,N_5689);
or U8276 (N_8276,N_4488,N_5075);
nor U8277 (N_8277,N_4331,N_4908);
nand U8278 (N_8278,N_5974,N_5423);
nand U8279 (N_8279,N_3710,N_3584);
or U8280 (N_8280,N_5680,N_4211);
and U8281 (N_8281,N_4058,N_3961);
and U8282 (N_8282,N_3706,N_4662);
nor U8283 (N_8283,N_3157,N_5760);
nor U8284 (N_8284,N_5680,N_3331);
or U8285 (N_8285,N_4583,N_5841);
nand U8286 (N_8286,N_5631,N_4866);
xor U8287 (N_8287,N_3550,N_4708);
or U8288 (N_8288,N_3396,N_3786);
or U8289 (N_8289,N_4302,N_3295);
and U8290 (N_8290,N_4656,N_4529);
or U8291 (N_8291,N_4925,N_3820);
nor U8292 (N_8292,N_5636,N_3704);
nor U8293 (N_8293,N_3212,N_5750);
nor U8294 (N_8294,N_4293,N_5283);
or U8295 (N_8295,N_5048,N_4137);
or U8296 (N_8296,N_3417,N_3339);
nor U8297 (N_8297,N_5440,N_3209);
nor U8298 (N_8298,N_4662,N_5772);
nand U8299 (N_8299,N_5938,N_5331);
and U8300 (N_8300,N_4526,N_3387);
or U8301 (N_8301,N_4994,N_3561);
or U8302 (N_8302,N_5247,N_3775);
nor U8303 (N_8303,N_5139,N_3314);
nor U8304 (N_8304,N_4313,N_5068);
or U8305 (N_8305,N_4375,N_5675);
or U8306 (N_8306,N_4684,N_3236);
nor U8307 (N_8307,N_4277,N_5794);
and U8308 (N_8308,N_4427,N_5038);
or U8309 (N_8309,N_5255,N_3223);
and U8310 (N_8310,N_4666,N_5395);
or U8311 (N_8311,N_4102,N_3874);
nor U8312 (N_8312,N_3615,N_3426);
and U8313 (N_8313,N_4280,N_4336);
or U8314 (N_8314,N_3255,N_5969);
and U8315 (N_8315,N_5825,N_3409);
and U8316 (N_8316,N_3686,N_4931);
nor U8317 (N_8317,N_5274,N_4343);
nand U8318 (N_8318,N_4387,N_3409);
or U8319 (N_8319,N_4434,N_4512);
nand U8320 (N_8320,N_4997,N_3750);
or U8321 (N_8321,N_4839,N_4389);
and U8322 (N_8322,N_3597,N_4546);
and U8323 (N_8323,N_5088,N_5058);
or U8324 (N_8324,N_3519,N_3593);
nand U8325 (N_8325,N_4597,N_5974);
or U8326 (N_8326,N_5108,N_3497);
nand U8327 (N_8327,N_3706,N_3985);
or U8328 (N_8328,N_5032,N_5789);
or U8329 (N_8329,N_3216,N_4518);
nand U8330 (N_8330,N_3385,N_3134);
and U8331 (N_8331,N_5167,N_3832);
or U8332 (N_8332,N_5181,N_4351);
or U8333 (N_8333,N_3173,N_5888);
and U8334 (N_8334,N_3087,N_3699);
nand U8335 (N_8335,N_4861,N_5343);
or U8336 (N_8336,N_5303,N_5035);
xor U8337 (N_8337,N_5095,N_3737);
and U8338 (N_8338,N_3320,N_3434);
and U8339 (N_8339,N_5461,N_5593);
and U8340 (N_8340,N_4913,N_3915);
or U8341 (N_8341,N_4128,N_3311);
nor U8342 (N_8342,N_4913,N_4338);
nor U8343 (N_8343,N_3540,N_4288);
and U8344 (N_8344,N_4111,N_5666);
and U8345 (N_8345,N_5408,N_4533);
xnor U8346 (N_8346,N_4897,N_5104);
or U8347 (N_8347,N_4983,N_3950);
and U8348 (N_8348,N_4532,N_4048);
and U8349 (N_8349,N_5379,N_3356);
nor U8350 (N_8350,N_3648,N_4519);
nand U8351 (N_8351,N_3782,N_3988);
nand U8352 (N_8352,N_3541,N_4397);
nor U8353 (N_8353,N_5334,N_5395);
nand U8354 (N_8354,N_4222,N_3923);
nor U8355 (N_8355,N_3439,N_4344);
nand U8356 (N_8356,N_5197,N_4303);
or U8357 (N_8357,N_4183,N_5590);
or U8358 (N_8358,N_4151,N_4098);
nor U8359 (N_8359,N_5897,N_3373);
or U8360 (N_8360,N_4525,N_5708);
and U8361 (N_8361,N_4601,N_3767);
nor U8362 (N_8362,N_5808,N_3110);
and U8363 (N_8363,N_3696,N_3109);
and U8364 (N_8364,N_3735,N_4065);
and U8365 (N_8365,N_3818,N_3364);
or U8366 (N_8366,N_4033,N_4219);
nand U8367 (N_8367,N_4245,N_4278);
and U8368 (N_8368,N_5059,N_5523);
nor U8369 (N_8369,N_5708,N_3861);
nand U8370 (N_8370,N_3808,N_3780);
nor U8371 (N_8371,N_4017,N_4385);
nand U8372 (N_8372,N_5734,N_3424);
nor U8373 (N_8373,N_3771,N_3578);
or U8374 (N_8374,N_5992,N_3575);
nor U8375 (N_8375,N_5155,N_5046);
nor U8376 (N_8376,N_4604,N_4315);
and U8377 (N_8377,N_4806,N_4942);
nand U8378 (N_8378,N_3539,N_4088);
nand U8379 (N_8379,N_4834,N_3393);
or U8380 (N_8380,N_4614,N_3545);
nor U8381 (N_8381,N_3506,N_3554);
xor U8382 (N_8382,N_3963,N_3124);
nand U8383 (N_8383,N_5354,N_5887);
or U8384 (N_8384,N_4926,N_3741);
nor U8385 (N_8385,N_4823,N_4431);
nor U8386 (N_8386,N_4099,N_5168);
nor U8387 (N_8387,N_5054,N_3403);
nor U8388 (N_8388,N_3473,N_3280);
nor U8389 (N_8389,N_3630,N_3858);
and U8390 (N_8390,N_3772,N_5713);
or U8391 (N_8391,N_5802,N_5969);
or U8392 (N_8392,N_4124,N_5931);
nand U8393 (N_8393,N_5886,N_5656);
nor U8394 (N_8394,N_4701,N_4452);
and U8395 (N_8395,N_5591,N_5652);
or U8396 (N_8396,N_5987,N_3696);
nand U8397 (N_8397,N_5029,N_5229);
nand U8398 (N_8398,N_3191,N_4435);
and U8399 (N_8399,N_4286,N_4917);
and U8400 (N_8400,N_3146,N_4382);
nand U8401 (N_8401,N_5762,N_3589);
and U8402 (N_8402,N_5787,N_4855);
and U8403 (N_8403,N_3029,N_3650);
nand U8404 (N_8404,N_5615,N_3626);
nand U8405 (N_8405,N_5686,N_3714);
and U8406 (N_8406,N_4074,N_4261);
nand U8407 (N_8407,N_3062,N_5543);
nor U8408 (N_8408,N_4168,N_5346);
or U8409 (N_8409,N_5434,N_3324);
nand U8410 (N_8410,N_5474,N_5042);
nor U8411 (N_8411,N_5210,N_4678);
nand U8412 (N_8412,N_5576,N_3674);
nor U8413 (N_8413,N_3751,N_3463);
or U8414 (N_8414,N_3784,N_5357);
nand U8415 (N_8415,N_5593,N_4991);
nor U8416 (N_8416,N_3108,N_3564);
or U8417 (N_8417,N_4068,N_3776);
nand U8418 (N_8418,N_5530,N_5119);
and U8419 (N_8419,N_5365,N_5514);
or U8420 (N_8420,N_5454,N_5891);
or U8421 (N_8421,N_4198,N_3957);
nor U8422 (N_8422,N_4209,N_3432);
and U8423 (N_8423,N_3581,N_5517);
or U8424 (N_8424,N_3620,N_4447);
nor U8425 (N_8425,N_3290,N_4568);
nor U8426 (N_8426,N_4218,N_4431);
nand U8427 (N_8427,N_4778,N_5623);
and U8428 (N_8428,N_3771,N_5999);
and U8429 (N_8429,N_3236,N_5786);
and U8430 (N_8430,N_4654,N_4506);
or U8431 (N_8431,N_5574,N_4270);
or U8432 (N_8432,N_5958,N_4743);
nor U8433 (N_8433,N_4746,N_5149);
and U8434 (N_8434,N_3190,N_3710);
or U8435 (N_8435,N_4395,N_3608);
nand U8436 (N_8436,N_3983,N_5202);
or U8437 (N_8437,N_5963,N_4712);
and U8438 (N_8438,N_4466,N_4284);
nand U8439 (N_8439,N_3060,N_5250);
and U8440 (N_8440,N_3023,N_4741);
and U8441 (N_8441,N_5169,N_5298);
and U8442 (N_8442,N_3269,N_5269);
nor U8443 (N_8443,N_3410,N_5890);
or U8444 (N_8444,N_4256,N_4664);
and U8445 (N_8445,N_4888,N_4781);
nand U8446 (N_8446,N_5181,N_3303);
nand U8447 (N_8447,N_3846,N_4088);
and U8448 (N_8448,N_5678,N_4638);
and U8449 (N_8449,N_4191,N_5134);
and U8450 (N_8450,N_4136,N_3400);
and U8451 (N_8451,N_3739,N_4756);
nand U8452 (N_8452,N_5820,N_3713);
and U8453 (N_8453,N_4821,N_5974);
and U8454 (N_8454,N_4223,N_4530);
nor U8455 (N_8455,N_3497,N_5477);
nor U8456 (N_8456,N_4427,N_3123);
nand U8457 (N_8457,N_4348,N_3946);
nor U8458 (N_8458,N_3219,N_5483);
nor U8459 (N_8459,N_5561,N_5797);
nand U8460 (N_8460,N_5883,N_5572);
or U8461 (N_8461,N_3617,N_3915);
nand U8462 (N_8462,N_4223,N_4332);
and U8463 (N_8463,N_5580,N_3924);
nor U8464 (N_8464,N_5147,N_3995);
or U8465 (N_8465,N_5476,N_5220);
nor U8466 (N_8466,N_5856,N_3827);
and U8467 (N_8467,N_5896,N_5704);
and U8468 (N_8468,N_5096,N_3517);
nand U8469 (N_8469,N_5887,N_3968);
or U8470 (N_8470,N_4476,N_5862);
nor U8471 (N_8471,N_5182,N_4486);
nor U8472 (N_8472,N_3551,N_5941);
or U8473 (N_8473,N_5616,N_4008);
xor U8474 (N_8474,N_3890,N_5991);
nor U8475 (N_8475,N_5131,N_3776);
and U8476 (N_8476,N_5602,N_5858);
nor U8477 (N_8477,N_3579,N_3295);
nor U8478 (N_8478,N_5544,N_5525);
nor U8479 (N_8479,N_4364,N_3490);
nand U8480 (N_8480,N_3242,N_5849);
nand U8481 (N_8481,N_4780,N_4726);
and U8482 (N_8482,N_3437,N_5131);
and U8483 (N_8483,N_5781,N_4799);
nand U8484 (N_8484,N_3861,N_3771);
nand U8485 (N_8485,N_5527,N_3808);
and U8486 (N_8486,N_5657,N_5731);
or U8487 (N_8487,N_5360,N_3543);
and U8488 (N_8488,N_3791,N_3108);
nor U8489 (N_8489,N_5802,N_5929);
nor U8490 (N_8490,N_4521,N_3885);
nand U8491 (N_8491,N_4689,N_4814);
or U8492 (N_8492,N_4363,N_5698);
and U8493 (N_8493,N_3406,N_4296);
and U8494 (N_8494,N_5619,N_5208);
and U8495 (N_8495,N_3819,N_3502);
or U8496 (N_8496,N_3038,N_3257);
or U8497 (N_8497,N_5487,N_4801);
xor U8498 (N_8498,N_5226,N_3893);
and U8499 (N_8499,N_5624,N_3978);
nor U8500 (N_8500,N_5879,N_3996);
nor U8501 (N_8501,N_3203,N_5784);
nand U8502 (N_8502,N_4511,N_3257);
and U8503 (N_8503,N_4704,N_4484);
and U8504 (N_8504,N_3439,N_5169);
and U8505 (N_8505,N_3161,N_4805);
nor U8506 (N_8506,N_3646,N_4481);
or U8507 (N_8507,N_4302,N_5934);
xor U8508 (N_8508,N_5839,N_4257);
or U8509 (N_8509,N_5179,N_3866);
nor U8510 (N_8510,N_5895,N_4222);
nor U8511 (N_8511,N_4974,N_4635);
nand U8512 (N_8512,N_4280,N_4224);
or U8513 (N_8513,N_5817,N_5737);
nand U8514 (N_8514,N_5794,N_5511);
and U8515 (N_8515,N_4575,N_3655);
nand U8516 (N_8516,N_3962,N_5580);
nand U8517 (N_8517,N_3334,N_5254);
nor U8518 (N_8518,N_5396,N_4799);
nand U8519 (N_8519,N_4987,N_3785);
nor U8520 (N_8520,N_5785,N_5689);
nand U8521 (N_8521,N_4588,N_3254);
and U8522 (N_8522,N_3221,N_5244);
nor U8523 (N_8523,N_3086,N_4219);
nor U8524 (N_8524,N_4603,N_3209);
and U8525 (N_8525,N_5699,N_4946);
or U8526 (N_8526,N_3348,N_4951);
nand U8527 (N_8527,N_3905,N_4689);
and U8528 (N_8528,N_4302,N_4956);
and U8529 (N_8529,N_3805,N_4065);
and U8530 (N_8530,N_4540,N_5272);
nand U8531 (N_8531,N_3757,N_4190);
nand U8532 (N_8532,N_4080,N_4045);
and U8533 (N_8533,N_4329,N_3716);
or U8534 (N_8534,N_3927,N_3221);
nor U8535 (N_8535,N_5571,N_5916);
and U8536 (N_8536,N_5170,N_3089);
and U8537 (N_8537,N_5395,N_4538);
and U8538 (N_8538,N_3841,N_5122);
xor U8539 (N_8539,N_4181,N_5025);
nor U8540 (N_8540,N_3241,N_3911);
and U8541 (N_8541,N_4589,N_4251);
and U8542 (N_8542,N_4096,N_4033);
nand U8543 (N_8543,N_5867,N_3771);
nor U8544 (N_8544,N_3982,N_4475);
nor U8545 (N_8545,N_5318,N_4316);
or U8546 (N_8546,N_5981,N_4676);
nand U8547 (N_8547,N_5069,N_4384);
or U8548 (N_8548,N_5090,N_4693);
nor U8549 (N_8549,N_5374,N_4037);
nand U8550 (N_8550,N_4891,N_4890);
and U8551 (N_8551,N_5896,N_4195);
nand U8552 (N_8552,N_5658,N_3841);
nor U8553 (N_8553,N_4658,N_3382);
and U8554 (N_8554,N_5152,N_4928);
nand U8555 (N_8555,N_5234,N_4913);
or U8556 (N_8556,N_3036,N_5538);
or U8557 (N_8557,N_4302,N_4384);
or U8558 (N_8558,N_3019,N_5750);
and U8559 (N_8559,N_3824,N_5700);
nand U8560 (N_8560,N_5769,N_3959);
and U8561 (N_8561,N_4530,N_5965);
nor U8562 (N_8562,N_4181,N_3696);
xor U8563 (N_8563,N_4866,N_5732);
nor U8564 (N_8564,N_5862,N_5031);
and U8565 (N_8565,N_4575,N_4247);
xor U8566 (N_8566,N_5101,N_5812);
and U8567 (N_8567,N_3479,N_3326);
nor U8568 (N_8568,N_3196,N_4880);
nand U8569 (N_8569,N_3530,N_3676);
xor U8570 (N_8570,N_4898,N_5467);
nor U8571 (N_8571,N_5602,N_5259);
nand U8572 (N_8572,N_4543,N_5122);
or U8573 (N_8573,N_4539,N_4176);
nor U8574 (N_8574,N_3820,N_3595);
and U8575 (N_8575,N_4396,N_4135);
nor U8576 (N_8576,N_5486,N_3690);
or U8577 (N_8577,N_4117,N_4391);
nand U8578 (N_8578,N_5882,N_4078);
nor U8579 (N_8579,N_5800,N_5092);
or U8580 (N_8580,N_3540,N_4904);
or U8581 (N_8581,N_3666,N_3095);
nand U8582 (N_8582,N_4768,N_4576);
or U8583 (N_8583,N_4268,N_5915);
and U8584 (N_8584,N_3448,N_3244);
nor U8585 (N_8585,N_4144,N_4158);
or U8586 (N_8586,N_5217,N_5000);
and U8587 (N_8587,N_3307,N_4600);
and U8588 (N_8588,N_4712,N_3713);
and U8589 (N_8589,N_3458,N_3487);
nor U8590 (N_8590,N_4688,N_5050);
or U8591 (N_8591,N_3015,N_5770);
xor U8592 (N_8592,N_5497,N_4581);
nor U8593 (N_8593,N_4255,N_5912);
nor U8594 (N_8594,N_4930,N_3743);
or U8595 (N_8595,N_3626,N_3177);
nor U8596 (N_8596,N_3391,N_3121);
and U8597 (N_8597,N_3645,N_3385);
nand U8598 (N_8598,N_4466,N_5538);
nor U8599 (N_8599,N_5299,N_5392);
and U8600 (N_8600,N_4679,N_4616);
nand U8601 (N_8601,N_3003,N_3427);
nor U8602 (N_8602,N_3792,N_3693);
nand U8603 (N_8603,N_3842,N_3901);
and U8604 (N_8604,N_3239,N_3746);
and U8605 (N_8605,N_4353,N_5496);
or U8606 (N_8606,N_4366,N_3793);
nor U8607 (N_8607,N_4831,N_3831);
nor U8608 (N_8608,N_4044,N_4601);
nand U8609 (N_8609,N_5365,N_5063);
or U8610 (N_8610,N_4628,N_3236);
and U8611 (N_8611,N_5546,N_4921);
nor U8612 (N_8612,N_3270,N_3668);
nor U8613 (N_8613,N_3175,N_5302);
nor U8614 (N_8614,N_4881,N_4728);
and U8615 (N_8615,N_4670,N_3800);
or U8616 (N_8616,N_5497,N_4044);
and U8617 (N_8617,N_4556,N_3874);
and U8618 (N_8618,N_5245,N_5270);
or U8619 (N_8619,N_3914,N_5800);
nor U8620 (N_8620,N_3563,N_4482);
and U8621 (N_8621,N_5689,N_3899);
nand U8622 (N_8622,N_3684,N_3335);
and U8623 (N_8623,N_4708,N_4568);
nor U8624 (N_8624,N_4145,N_4070);
nor U8625 (N_8625,N_4714,N_5193);
nor U8626 (N_8626,N_5354,N_4665);
nor U8627 (N_8627,N_3887,N_3174);
nor U8628 (N_8628,N_4472,N_4892);
nand U8629 (N_8629,N_5860,N_3351);
nor U8630 (N_8630,N_4192,N_5941);
nand U8631 (N_8631,N_5616,N_4557);
nor U8632 (N_8632,N_5164,N_4904);
nand U8633 (N_8633,N_5235,N_4092);
or U8634 (N_8634,N_3322,N_5926);
or U8635 (N_8635,N_4018,N_3198);
or U8636 (N_8636,N_3934,N_5334);
nor U8637 (N_8637,N_3641,N_3091);
nand U8638 (N_8638,N_5898,N_5908);
or U8639 (N_8639,N_3144,N_3825);
nand U8640 (N_8640,N_5518,N_3400);
nor U8641 (N_8641,N_4614,N_3727);
and U8642 (N_8642,N_3091,N_3953);
nand U8643 (N_8643,N_5089,N_5327);
nor U8644 (N_8644,N_4319,N_4012);
xnor U8645 (N_8645,N_5405,N_3165);
nor U8646 (N_8646,N_4711,N_4340);
or U8647 (N_8647,N_4365,N_3727);
or U8648 (N_8648,N_5228,N_4104);
nand U8649 (N_8649,N_5026,N_4711);
nand U8650 (N_8650,N_4816,N_4331);
and U8651 (N_8651,N_3004,N_4153);
and U8652 (N_8652,N_4408,N_4728);
and U8653 (N_8653,N_5973,N_3054);
nand U8654 (N_8654,N_3424,N_5303);
and U8655 (N_8655,N_4080,N_5597);
and U8656 (N_8656,N_3783,N_4215);
nand U8657 (N_8657,N_4831,N_5953);
nand U8658 (N_8658,N_3549,N_4356);
or U8659 (N_8659,N_3207,N_3564);
nor U8660 (N_8660,N_5424,N_5084);
and U8661 (N_8661,N_3950,N_3834);
nor U8662 (N_8662,N_4017,N_5197);
or U8663 (N_8663,N_4677,N_5983);
nand U8664 (N_8664,N_4965,N_3537);
and U8665 (N_8665,N_3950,N_4594);
or U8666 (N_8666,N_3662,N_4820);
nor U8667 (N_8667,N_4193,N_4415);
and U8668 (N_8668,N_5576,N_3097);
nand U8669 (N_8669,N_5179,N_3753);
nand U8670 (N_8670,N_5045,N_4998);
or U8671 (N_8671,N_4644,N_3008);
nand U8672 (N_8672,N_3699,N_3580);
nand U8673 (N_8673,N_5522,N_5448);
or U8674 (N_8674,N_3149,N_3548);
or U8675 (N_8675,N_5422,N_4342);
or U8676 (N_8676,N_5527,N_5509);
nand U8677 (N_8677,N_5882,N_3913);
and U8678 (N_8678,N_3531,N_5925);
xnor U8679 (N_8679,N_5363,N_4788);
or U8680 (N_8680,N_3422,N_3796);
or U8681 (N_8681,N_3178,N_3983);
or U8682 (N_8682,N_4506,N_5869);
or U8683 (N_8683,N_4439,N_4645);
nor U8684 (N_8684,N_4578,N_3272);
or U8685 (N_8685,N_4359,N_5538);
nand U8686 (N_8686,N_5129,N_4554);
nor U8687 (N_8687,N_4537,N_5679);
and U8688 (N_8688,N_5626,N_4544);
or U8689 (N_8689,N_5906,N_3288);
nand U8690 (N_8690,N_4295,N_5869);
or U8691 (N_8691,N_3323,N_3091);
nand U8692 (N_8692,N_4892,N_4722);
nand U8693 (N_8693,N_5040,N_3307);
and U8694 (N_8694,N_5696,N_5578);
nand U8695 (N_8695,N_3331,N_3582);
nor U8696 (N_8696,N_4713,N_4029);
nand U8697 (N_8697,N_4997,N_3414);
or U8698 (N_8698,N_3596,N_4956);
and U8699 (N_8699,N_4443,N_3902);
nand U8700 (N_8700,N_3359,N_5381);
nand U8701 (N_8701,N_5409,N_4730);
nor U8702 (N_8702,N_4027,N_3082);
and U8703 (N_8703,N_3077,N_3581);
or U8704 (N_8704,N_3634,N_5614);
and U8705 (N_8705,N_5203,N_4712);
or U8706 (N_8706,N_3524,N_4040);
nor U8707 (N_8707,N_4937,N_3208);
and U8708 (N_8708,N_5173,N_3322);
nand U8709 (N_8709,N_4665,N_3267);
nor U8710 (N_8710,N_4043,N_4818);
and U8711 (N_8711,N_5918,N_5077);
nand U8712 (N_8712,N_5654,N_3584);
nor U8713 (N_8713,N_3608,N_3498);
nor U8714 (N_8714,N_4291,N_4007);
and U8715 (N_8715,N_4067,N_5459);
nand U8716 (N_8716,N_4718,N_4284);
nor U8717 (N_8717,N_4127,N_3234);
or U8718 (N_8718,N_3745,N_3133);
nor U8719 (N_8719,N_5625,N_3693);
and U8720 (N_8720,N_3361,N_4253);
nand U8721 (N_8721,N_4503,N_5408);
nand U8722 (N_8722,N_5770,N_3245);
nand U8723 (N_8723,N_3825,N_4001);
and U8724 (N_8724,N_3488,N_5924);
or U8725 (N_8725,N_4098,N_3969);
nor U8726 (N_8726,N_5226,N_4383);
nor U8727 (N_8727,N_3690,N_5677);
or U8728 (N_8728,N_5335,N_3120);
nand U8729 (N_8729,N_3840,N_5371);
nand U8730 (N_8730,N_4914,N_4045);
nand U8731 (N_8731,N_4860,N_3966);
nand U8732 (N_8732,N_5090,N_4190);
nand U8733 (N_8733,N_3151,N_5077);
nand U8734 (N_8734,N_3231,N_3671);
and U8735 (N_8735,N_5584,N_4582);
nor U8736 (N_8736,N_3451,N_3154);
or U8737 (N_8737,N_5657,N_5459);
nor U8738 (N_8738,N_4331,N_4722);
or U8739 (N_8739,N_3567,N_5623);
nor U8740 (N_8740,N_5301,N_3692);
nand U8741 (N_8741,N_5713,N_4163);
nand U8742 (N_8742,N_5931,N_4428);
or U8743 (N_8743,N_3779,N_5832);
nor U8744 (N_8744,N_4302,N_5152);
or U8745 (N_8745,N_5507,N_4030);
nor U8746 (N_8746,N_4749,N_3914);
nor U8747 (N_8747,N_4116,N_3448);
nand U8748 (N_8748,N_3982,N_4484);
nor U8749 (N_8749,N_4772,N_4785);
nor U8750 (N_8750,N_4526,N_3493);
nand U8751 (N_8751,N_4706,N_4723);
or U8752 (N_8752,N_4827,N_5996);
or U8753 (N_8753,N_3700,N_5610);
and U8754 (N_8754,N_4714,N_5698);
or U8755 (N_8755,N_3377,N_4590);
and U8756 (N_8756,N_5188,N_5501);
or U8757 (N_8757,N_5653,N_5835);
nand U8758 (N_8758,N_5965,N_5344);
nor U8759 (N_8759,N_5516,N_5278);
or U8760 (N_8760,N_3710,N_5017);
xor U8761 (N_8761,N_3545,N_4000);
or U8762 (N_8762,N_3119,N_3309);
or U8763 (N_8763,N_4794,N_3079);
and U8764 (N_8764,N_4348,N_5558);
or U8765 (N_8765,N_3108,N_4767);
or U8766 (N_8766,N_5516,N_4278);
or U8767 (N_8767,N_4687,N_5430);
nor U8768 (N_8768,N_5595,N_4474);
or U8769 (N_8769,N_3098,N_4183);
nand U8770 (N_8770,N_4169,N_5304);
nand U8771 (N_8771,N_5553,N_5898);
or U8772 (N_8772,N_3490,N_3273);
and U8773 (N_8773,N_4050,N_5594);
and U8774 (N_8774,N_4997,N_3250);
and U8775 (N_8775,N_4171,N_5723);
nor U8776 (N_8776,N_3809,N_4183);
or U8777 (N_8777,N_5843,N_5815);
and U8778 (N_8778,N_5965,N_3848);
nor U8779 (N_8779,N_5840,N_3140);
and U8780 (N_8780,N_5369,N_4221);
or U8781 (N_8781,N_3069,N_4452);
or U8782 (N_8782,N_5895,N_3247);
and U8783 (N_8783,N_3992,N_4485);
or U8784 (N_8784,N_4695,N_4428);
and U8785 (N_8785,N_5748,N_4474);
and U8786 (N_8786,N_3751,N_4211);
nor U8787 (N_8787,N_3918,N_3129);
or U8788 (N_8788,N_5240,N_3267);
and U8789 (N_8789,N_5354,N_4833);
nand U8790 (N_8790,N_4509,N_5806);
nand U8791 (N_8791,N_5356,N_5842);
nand U8792 (N_8792,N_4564,N_5867);
and U8793 (N_8793,N_5270,N_5769);
nand U8794 (N_8794,N_5115,N_5186);
or U8795 (N_8795,N_4107,N_4843);
or U8796 (N_8796,N_5342,N_3791);
nand U8797 (N_8797,N_4331,N_5234);
nor U8798 (N_8798,N_5843,N_4782);
nor U8799 (N_8799,N_5803,N_5683);
and U8800 (N_8800,N_4890,N_4486);
nand U8801 (N_8801,N_5304,N_3957);
or U8802 (N_8802,N_4729,N_5197);
nand U8803 (N_8803,N_3869,N_4248);
and U8804 (N_8804,N_4275,N_4244);
and U8805 (N_8805,N_5223,N_5174);
or U8806 (N_8806,N_4879,N_3362);
nand U8807 (N_8807,N_5197,N_5268);
or U8808 (N_8808,N_5951,N_3718);
nand U8809 (N_8809,N_4611,N_5542);
and U8810 (N_8810,N_3963,N_4267);
or U8811 (N_8811,N_3282,N_3801);
and U8812 (N_8812,N_5440,N_4360);
or U8813 (N_8813,N_3114,N_3395);
and U8814 (N_8814,N_4163,N_4151);
or U8815 (N_8815,N_5469,N_5179);
or U8816 (N_8816,N_3375,N_4951);
nand U8817 (N_8817,N_4389,N_4055);
or U8818 (N_8818,N_3645,N_3206);
and U8819 (N_8819,N_3115,N_4590);
nand U8820 (N_8820,N_5265,N_5688);
nand U8821 (N_8821,N_3874,N_4487);
and U8822 (N_8822,N_4435,N_3968);
nand U8823 (N_8823,N_4423,N_3703);
nor U8824 (N_8824,N_3330,N_3725);
and U8825 (N_8825,N_3440,N_4077);
nor U8826 (N_8826,N_3043,N_5171);
nor U8827 (N_8827,N_3901,N_3474);
or U8828 (N_8828,N_4467,N_3612);
and U8829 (N_8829,N_3176,N_5721);
or U8830 (N_8830,N_5871,N_4251);
and U8831 (N_8831,N_4616,N_3583);
and U8832 (N_8832,N_5746,N_3509);
nor U8833 (N_8833,N_5925,N_4631);
and U8834 (N_8834,N_3146,N_3618);
nor U8835 (N_8835,N_3618,N_3042);
and U8836 (N_8836,N_5327,N_3598);
nand U8837 (N_8837,N_5243,N_4983);
nand U8838 (N_8838,N_4699,N_3724);
and U8839 (N_8839,N_3151,N_5852);
nor U8840 (N_8840,N_4747,N_4908);
nor U8841 (N_8841,N_4285,N_5787);
and U8842 (N_8842,N_5986,N_4845);
and U8843 (N_8843,N_4248,N_3424);
and U8844 (N_8844,N_4625,N_4735);
and U8845 (N_8845,N_4014,N_4327);
nand U8846 (N_8846,N_5622,N_3021);
nor U8847 (N_8847,N_5746,N_4093);
and U8848 (N_8848,N_3876,N_3744);
or U8849 (N_8849,N_4837,N_4307);
nand U8850 (N_8850,N_4639,N_4635);
and U8851 (N_8851,N_4793,N_3686);
or U8852 (N_8852,N_5640,N_3185);
nor U8853 (N_8853,N_3381,N_3426);
nor U8854 (N_8854,N_4469,N_4765);
nand U8855 (N_8855,N_5911,N_4094);
and U8856 (N_8856,N_5002,N_5046);
nor U8857 (N_8857,N_4089,N_5381);
nand U8858 (N_8858,N_4957,N_4984);
and U8859 (N_8859,N_5958,N_3440);
or U8860 (N_8860,N_3705,N_5476);
and U8861 (N_8861,N_3403,N_3524);
nand U8862 (N_8862,N_3908,N_3319);
nand U8863 (N_8863,N_4536,N_5282);
nor U8864 (N_8864,N_4893,N_5008);
or U8865 (N_8865,N_4153,N_4459);
and U8866 (N_8866,N_4005,N_4765);
nand U8867 (N_8867,N_3503,N_3289);
nand U8868 (N_8868,N_4393,N_5138);
or U8869 (N_8869,N_4747,N_5392);
or U8870 (N_8870,N_5883,N_3276);
nand U8871 (N_8871,N_5111,N_4808);
and U8872 (N_8872,N_3500,N_4153);
and U8873 (N_8873,N_5259,N_4035);
nor U8874 (N_8874,N_3198,N_3963);
nor U8875 (N_8875,N_4586,N_4914);
and U8876 (N_8876,N_5843,N_4083);
and U8877 (N_8877,N_4152,N_4351);
or U8878 (N_8878,N_3293,N_3928);
and U8879 (N_8879,N_5892,N_3266);
nand U8880 (N_8880,N_3439,N_5340);
and U8881 (N_8881,N_5307,N_3675);
or U8882 (N_8882,N_3484,N_3443);
nand U8883 (N_8883,N_4106,N_5079);
or U8884 (N_8884,N_4980,N_3127);
and U8885 (N_8885,N_4301,N_4095);
nand U8886 (N_8886,N_4315,N_3770);
and U8887 (N_8887,N_5880,N_3325);
nor U8888 (N_8888,N_5899,N_5433);
and U8889 (N_8889,N_4732,N_3757);
nand U8890 (N_8890,N_4214,N_3588);
nor U8891 (N_8891,N_5736,N_3164);
or U8892 (N_8892,N_3547,N_3056);
and U8893 (N_8893,N_5024,N_4819);
nor U8894 (N_8894,N_5062,N_5619);
and U8895 (N_8895,N_5457,N_4389);
nand U8896 (N_8896,N_5874,N_5104);
or U8897 (N_8897,N_4618,N_5722);
nand U8898 (N_8898,N_3340,N_4097);
nor U8899 (N_8899,N_3232,N_4369);
and U8900 (N_8900,N_5532,N_4136);
nand U8901 (N_8901,N_4355,N_3703);
and U8902 (N_8902,N_3157,N_5223);
or U8903 (N_8903,N_3915,N_4379);
and U8904 (N_8904,N_5935,N_4435);
nand U8905 (N_8905,N_3063,N_4178);
xnor U8906 (N_8906,N_3981,N_4305);
nand U8907 (N_8907,N_3039,N_3116);
and U8908 (N_8908,N_5347,N_5754);
and U8909 (N_8909,N_5737,N_5327);
and U8910 (N_8910,N_3360,N_5567);
xnor U8911 (N_8911,N_3699,N_5990);
nor U8912 (N_8912,N_4331,N_5980);
or U8913 (N_8913,N_3498,N_5672);
and U8914 (N_8914,N_3632,N_5362);
nor U8915 (N_8915,N_5849,N_5554);
nor U8916 (N_8916,N_5307,N_5104);
and U8917 (N_8917,N_4571,N_5205);
nand U8918 (N_8918,N_4428,N_3615);
or U8919 (N_8919,N_5465,N_4171);
nor U8920 (N_8920,N_4704,N_5445);
nand U8921 (N_8921,N_5490,N_4751);
nand U8922 (N_8922,N_5560,N_3477);
xnor U8923 (N_8923,N_3463,N_4365);
or U8924 (N_8924,N_5928,N_5542);
or U8925 (N_8925,N_4529,N_5324);
nor U8926 (N_8926,N_5159,N_4494);
or U8927 (N_8927,N_5082,N_5191);
nor U8928 (N_8928,N_4173,N_3578);
and U8929 (N_8929,N_4279,N_3543);
nand U8930 (N_8930,N_4498,N_5999);
nand U8931 (N_8931,N_4558,N_5432);
or U8932 (N_8932,N_3629,N_4231);
or U8933 (N_8933,N_5719,N_4489);
and U8934 (N_8934,N_3145,N_5829);
nor U8935 (N_8935,N_5520,N_3363);
and U8936 (N_8936,N_3932,N_4780);
or U8937 (N_8937,N_4555,N_5648);
nand U8938 (N_8938,N_5534,N_3548);
or U8939 (N_8939,N_4440,N_5903);
and U8940 (N_8940,N_5363,N_3075);
nor U8941 (N_8941,N_4187,N_4330);
nor U8942 (N_8942,N_4365,N_5188);
nor U8943 (N_8943,N_5062,N_4636);
nand U8944 (N_8944,N_4376,N_4818);
nor U8945 (N_8945,N_4639,N_4281);
or U8946 (N_8946,N_5736,N_5920);
or U8947 (N_8947,N_4592,N_5721);
nor U8948 (N_8948,N_4706,N_4869);
nor U8949 (N_8949,N_4206,N_5857);
nor U8950 (N_8950,N_5505,N_3022);
nor U8951 (N_8951,N_3242,N_3559);
and U8952 (N_8952,N_3962,N_5594);
and U8953 (N_8953,N_3574,N_5547);
or U8954 (N_8954,N_3550,N_3006);
or U8955 (N_8955,N_4630,N_5723);
and U8956 (N_8956,N_4316,N_5386);
and U8957 (N_8957,N_4133,N_3905);
nor U8958 (N_8958,N_4989,N_4324);
nor U8959 (N_8959,N_4411,N_3328);
nor U8960 (N_8960,N_3397,N_5315);
nand U8961 (N_8961,N_4575,N_3481);
and U8962 (N_8962,N_4445,N_3912);
and U8963 (N_8963,N_4611,N_4037);
or U8964 (N_8964,N_3106,N_3802);
nor U8965 (N_8965,N_4631,N_5143);
and U8966 (N_8966,N_5114,N_5716);
nand U8967 (N_8967,N_3920,N_3941);
nor U8968 (N_8968,N_5460,N_4101);
nor U8969 (N_8969,N_5259,N_5546);
nor U8970 (N_8970,N_3796,N_3040);
and U8971 (N_8971,N_4802,N_3192);
nor U8972 (N_8972,N_3540,N_5577);
nand U8973 (N_8973,N_4936,N_5925);
or U8974 (N_8974,N_5483,N_4574);
nor U8975 (N_8975,N_4990,N_3263);
and U8976 (N_8976,N_5855,N_5587);
nor U8977 (N_8977,N_4147,N_5053);
nand U8978 (N_8978,N_4844,N_5352);
nor U8979 (N_8979,N_5582,N_4821);
and U8980 (N_8980,N_3190,N_5586);
or U8981 (N_8981,N_3632,N_3700);
nand U8982 (N_8982,N_5340,N_3279);
and U8983 (N_8983,N_3443,N_3004);
and U8984 (N_8984,N_4231,N_5710);
and U8985 (N_8985,N_3117,N_3959);
nand U8986 (N_8986,N_3730,N_3027);
nor U8987 (N_8987,N_5336,N_3056);
or U8988 (N_8988,N_3561,N_5579);
nor U8989 (N_8989,N_3659,N_4928);
or U8990 (N_8990,N_5626,N_3501);
or U8991 (N_8991,N_5135,N_4045);
nand U8992 (N_8992,N_3189,N_3802);
nor U8993 (N_8993,N_4562,N_3069);
nand U8994 (N_8994,N_5264,N_5484);
or U8995 (N_8995,N_3758,N_4601);
and U8996 (N_8996,N_4655,N_3730);
and U8997 (N_8997,N_3804,N_4435);
and U8998 (N_8998,N_5744,N_5606);
or U8999 (N_8999,N_5741,N_4457);
nor U9000 (N_9000,N_8893,N_7710);
or U9001 (N_9001,N_8385,N_6901);
nor U9002 (N_9002,N_8989,N_7147);
and U9003 (N_9003,N_6375,N_8520);
or U9004 (N_9004,N_7155,N_7808);
and U9005 (N_9005,N_6224,N_7583);
nand U9006 (N_9006,N_6282,N_8930);
nand U9007 (N_9007,N_6364,N_8505);
nor U9008 (N_9008,N_7036,N_6144);
nor U9009 (N_9009,N_8288,N_7639);
and U9010 (N_9010,N_8066,N_7796);
nand U9011 (N_9011,N_8920,N_8702);
nor U9012 (N_9012,N_6138,N_7196);
and U9013 (N_9013,N_7383,N_8118);
or U9014 (N_9014,N_8231,N_7663);
and U9015 (N_9015,N_6530,N_6640);
nand U9016 (N_9016,N_6365,N_7990);
nand U9017 (N_9017,N_7223,N_7231);
nand U9018 (N_9018,N_8701,N_8349);
or U9019 (N_9019,N_6992,N_8194);
or U9020 (N_9020,N_7309,N_8939);
or U9021 (N_9021,N_8403,N_7982);
nor U9022 (N_9022,N_8183,N_6795);
or U9023 (N_9023,N_7989,N_8020);
and U9024 (N_9024,N_8190,N_8793);
or U9025 (N_9025,N_8658,N_8299);
nor U9026 (N_9026,N_8218,N_7740);
nor U9027 (N_9027,N_7855,N_6082);
nand U9028 (N_9028,N_6918,N_8142);
nor U9029 (N_9029,N_8398,N_6195);
nand U9030 (N_9030,N_6738,N_7974);
nor U9031 (N_9031,N_7074,N_8728);
nor U9032 (N_9032,N_7322,N_6917);
nand U9033 (N_9033,N_8377,N_6476);
or U9034 (N_9034,N_6499,N_7872);
or U9035 (N_9035,N_8139,N_7542);
or U9036 (N_9036,N_6656,N_8626);
nand U9037 (N_9037,N_8119,N_6950);
nor U9038 (N_9038,N_8980,N_8443);
nand U9039 (N_9039,N_6725,N_7133);
or U9040 (N_9040,N_8446,N_8228);
and U9041 (N_9041,N_8102,N_7550);
and U9042 (N_9042,N_6077,N_7308);
or U9043 (N_9043,N_8061,N_8570);
and U9044 (N_9044,N_6426,N_6264);
nor U9045 (N_9045,N_6785,N_8192);
or U9046 (N_9046,N_8226,N_6033);
and U9047 (N_9047,N_8411,N_6178);
nand U9048 (N_9048,N_6019,N_6047);
nor U9049 (N_9049,N_8749,N_7441);
or U9050 (N_9050,N_8967,N_8327);
nor U9051 (N_9051,N_7830,N_8365);
or U9052 (N_9052,N_6261,N_7859);
or U9053 (N_9053,N_8912,N_8915);
or U9054 (N_9054,N_7464,N_7827);
nor U9055 (N_9055,N_6602,N_8393);
and U9056 (N_9056,N_7081,N_6312);
or U9057 (N_9057,N_8290,N_8618);
nor U9058 (N_9058,N_6865,N_7554);
and U9059 (N_9059,N_6230,N_8986);
xor U9060 (N_9060,N_6971,N_7440);
or U9061 (N_9061,N_6354,N_8925);
or U9062 (N_9062,N_8379,N_8448);
nor U9063 (N_9063,N_6863,N_6319);
or U9064 (N_9064,N_6960,N_7613);
or U9065 (N_9065,N_8207,N_7871);
or U9066 (N_9066,N_7140,N_8597);
nand U9067 (N_9067,N_6808,N_8491);
and U9068 (N_9068,N_6652,N_8851);
nand U9069 (N_9069,N_7296,N_8787);
nor U9070 (N_9070,N_8017,N_6616);
nand U9071 (N_9071,N_8865,N_8117);
or U9072 (N_9072,N_8179,N_7574);
nand U9073 (N_9073,N_8496,N_6356);
nor U9074 (N_9074,N_7173,N_7065);
or U9075 (N_9075,N_6945,N_8014);
and U9076 (N_9076,N_6828,N_6151);
or U9077 (N_9077,N_6043,N_7466);
nand U9078 (N_9078,N_7046,N_7992);
nand U9079 (N_9079,N_6956,N_6205);
and U9080 (N_9080,N_7237,N_6843);
nand U9081 (N_9081,N_7163,N_8441);
and U9082 (N_9082,N_8069,N_6078);
xor U9083 (N_9083,N_8503,N_8331);
or U9084 (N_9084,N_8741,N_6771);
nor U9085 (N_9085,N_8959,N_6131);
and U9086 (N_9086,N_7080,N_6957);
nor U9087 (N_9087,N_6542,N_6632);
nand U9088 (N_9088,N_6050,N_6774);
xor U9089 (N_9089,N_8303,N_6366);
nor U9090 (N_9090,N_8631,N_8193);
nor U9091 (N_9091,N_6804,N_6601);
nor U9092 (N_9092,N_6471,N_8455);
and U9093 (N_9093,N_7653,N_8896);
nor U9094 (N_9094,N_7731,N_8601);
and U9095 (N_9095,N_8333,N_6904);
nand U9096 (N_9096,N_6288,N_8780);
and U9097 (N_9097,N_8151,N_8525);
nand U9098 (N_9098,N_7443,N_8990);
xor U9099 (N_9099,N_6496,N_8350);
or U9100 (N_9100,N_7953,N_7528);
and U9101 (N_9101,N_6767,N_7183);
xor U9102 (N_9102,N_6299,N_7136);
and U9103 (N_9103,N_8033,N_8425);
nand U9104 (N_9104,N_7555,N_6036);
nor U9105 (N_9105,N_6812,N_8090);
and U9106 (N_9106,N_6528,N_8673);
nand U9107 (N_9107,N_7540,N_8273);
nor U9108 (N_9108,N_8308,N_8733);
nor U9109 (N_9109,N_8594,N_6381);
and U9110 (N_9110,N_7134,N_8846);
or U9111 (N_9111,N_8616,N_7750);
nand U9112 (N_9112,N_6141,N_7465);
nand U9113 (N_9113,N_7190,N_7626);
nand U9114 (N_9114,N_6126,N_7253);
nor U9115 (N_9115,N_7338,N_6711);
nand U9116 (N_9116,N_6715,N_6815);
or U9117 (N_9117,N_8278,N_7592);
or U9118 (N_9118,N_8711,N_7543);
and U9119 (N_9119,N_7432,N_8531);
nor U9120 (N_9120,N_6959,N_6636);
or U9121 (N_9121,N_7130,N_8312);
or U9122 (N_9122,N_8497,N_6493);
or U9123 (N_9123,N_8382,N_6085);
or U9124 (N_9124,N_8633,N_7558);
and U9125 (N_9125,N_6521,N_6799);
and U9126 (N_9126,N_6820,N_6106);
nand U9127 (N_9127,N_8129,N_7460);
nand U9128 (N_9128,N_7960,N_7525);
nor U9129 (N_9129,N_6645,N_8574);
and U9130 (N_9130,N_8575,N_8074);
or U9131 (N_9131,N_8970,N_7354);
nor U9132 (N_9132,N_7670,N_8929);
nor U9133 (N_9133,N_8806,N_6534);
nand U9134 (N_9134,N_6630,N_8763);
or U9135 (N_9135,N_7621,N_6765);
and U9136 (N_9136,N_6303,N_8748);
or U9137 (N_9137,N_8271,N_6497);
nor U9138 (N_9138,N_7851,N_8470);
nor U9139 (N_9139,N_6407,N_6213);
or U9140 (N_9140,N_7415,N_7283);
and U9141 (N_9141,N_7531,N_7204);
nor U9142 (N_9142,N_6218,N_8072);
and U9143 (N_9143,N_7921,N_6900);
nor U9144 (N_9144,N_8814,N_6679);
nand U9145 (N_9145,N_6995,N_7243);
nor U9146 (N_9146,N_8461,N_6391);
or U9147 (N_9147,N_8241,N_7222);
nand U9148 (N_9148,N_6245,N_6096);
nand U9149 (N_9149,N_8250,N_6981);
or U9150 (N_9150,N_7366,N_7300);
nand U9151 (N_9151,N_7552,N_7735);
nand U9152 (N_9152,N_8945,N_7025);
and U9153 (N_9153,N_6897,N_8751);
nor U9154 (N_9154,N_6739,N_7180);
and U9155 (N_9155,N_6545,N_8084);
or U9156 (N_9156,N_8623,N_7291);
nand U9157 (N_9157,N_8657,N_6993);
nand U9158 (N_9158,N_7629,N_6017);
nor U9159 (N_9159,N_8589,N_6349);
nand U9160 (N_9160,N_7676,N_7571);
or U9161 (N_9161,N_6851,N_8395);
nand U9162 (N_9162,N_8434,N_6063);
nor U9163 (N_9163,N_7593,N_8476);
or U9164 (N_9164,N_7251,N_6609);
or U9165 (N_9165,N_8164,N_6886);
and U9166 (N_9166,N_7514,N_6726);
nor U9167 (N_9167,N_8484,N_8988);
or U9168 (N_9168,N_8720,N_7430);
nor U9169 (N_9169,N_7813,N_7567);
or U9170 (N_9170,N_6729,N_6223);
nand U9171 (N_9171,N_8849,N_7882);
nor U9172 (N_9172,N_7809,N_7482);
nor U9173 (N_9173,N_6667,N_7433);
nor U9174 (N_9174,N_8962,N_6604);
and U9175 (N_9175,N_6395,N_8855);
or U9176 (N_9176,N_7556,N_7193);
nand U9177 (N_9177,N_8059,N_7880);
nand U9178 (N_9178,N_7890,N_8977);
or U9179 (N_9179,N_6403,N_8955);
or U9180 (N_9180,N_7759,N_8895);
nor U9181 (N_9181,N_7245,N_6177);
or U9182 (N_9182,N_7779,N_6776);
or U9183 (N_9183,N_7927,N_7491);
nand U9184 (N_9184,N_6332,N_7776);
or U9185 (N_9185,N_8794,N_8115);
nor U9186 (N_9186,N_7801,N_7067);
nor U9187 (N_9187,N_6583,N_7449);
nor U9188 (N_9188,N_6919,N_6143);
nor U9189 (N_9189,N_8902,N_6589);
xor U9190 (N_9190,N_7211,N_8202);
nand U9191 (N_9191,N_8901,N_8587);
and U9192 (N_9192,N_7764,N_8219);
nand U9193 (N_9193,N_8807,N_7458);
or U9194 (N_9194,N_7631,N_7993);
or U9195 (N_9195,N_8454,N_6859);
and U9196 (N_9196,N_8847,N_6340);
nor U9197 (N_9197,N_8857,N_8176);
nor U9198 (N_9198,N_8705,N_7568);
or U9199 (N_9199,N_7429,N_6631);
or U9200 (N_9200,N_8622,N_8289);
nand U9201 (N_9201,N_6121,N_8602);
nand U9202 (N_9202,N_8905,N_7703);
or U9203 (N_9203,N_7050,N_6116);
and U9204 (N_9204,N_7368,N_8047);
or U9205 (N_9205,N_7785,N_7185);
and U9206 (N_9206,N_6049,N_8285);
and U9207 (N_9207,N_7461,N_7697);
nand U9208 (N_9208,N_7869,N_7124);
or U9209 (N_9209,N_8573,N_7701);
nand U9210 (N_9210,N_8511,N_8991);
or U9211 (N_9211,N_8146,N_8405);
nor U9212 (N_9212,N_7945,N_7055);
nand U9213 (N_9213,N_8076,N_8783);
nor U9214 (N_9214,N_6228,N_7382);
or U9215 (N_9215,N_8615,N_7267);
nand U9216 (N_9216,N_6461,N_8105);
nand U9217 (N_9217,N_8255,N_7570);
or U9218 (N_9218,N_8931,N_7339);
and U9219 (N_9219,N_8042,N_7478);
xnor U9220 (N_9220,N_8707,N_7395);
nor U9221 (N_9221,N_8655,N_7535);
nand U9222 (N_9222,N_6650,N_6281);
or U9223 (N_9223,N_8824,N_7580);
or U9224 (N_9224,N_6582,N_6701);
nor U9225 (N_9225,N_7889,N_6302);
or U9226 (N_9226,N_7634,N_7043);
and U9227 (N_9227,N_8532,N_7011);
nor U9228 (N_9228,N_8956,N_8029);
and U9229 (N_9229,N_7792,N_8843);
nor U9230 (N_9230,N_6953,N_8314);
or U9231 (N_9231,N_8325,N_8736);
and U9232 (N_9232,N_7874,N_7757);
or U9233 (N_9233,N_6973,N_6201);
nand U9234 (N_9234,N_8709,N_7506);
or U9235 (N_9235,N_8232,N_6994);
nor U9236 (N_9236,N_8892,N_6814);
nor U9237 (N_9237,N_7729,N_6980);
nand U9238 (N_9238,N_6662,N_8798);
nor U9239 (N_9239,N_6501,N_6301);
nor U9240 (N_9240,N_7840,N_8433);
or U9241 (N_9241,N_6028,N_7484);
nand U9242 (N_9242,N_7344,N_6753);
and U9243 (N_9243,N_8872,N_6044);
and U9244 (N_9244,N_6067,N_6089);
nor U9245 (N_9245,N_6690,N_7157);
and U9246 (N_9246,N_6517,N_8914);
or U9247 (N_9247,N_7746,N_7797);
nand U9248 (N_9248,N_8717,N_6452);
or U9249 (N_9249,N_8442,N_7380);
and U9250 (N_9250,N_6551,N_6833);
nand U9251 (N_9251,N_6238,N_7501);
and U9252 (N_9252,N_7643,N_6877);
nor U9253 (N_9253,N_7557,N_6405);
or U9254 (N_9254,N_6194,N_7700);
nand U9255 (N_9255,N_6084,N_6259);
nor U9256 (N_9256,N_8121,N_6117);
and U9257 (N_9257,N_6304,N_7452);
nor U9258 (N_9258,N_8721,N_6346);
or U9259 (N_9259,N_7837,N_6253);
and U9260 (N_9260,N_6578,N_8187);
or U9261 (N_9261,N_8800,N_7958);
or U9262 (N_9262,N_6884,N_8863);
nor U9263 (N_9263,N_7563,N_7044);
nand U9264 (N_9264,N_8553,N_7728);
and U9265 (N_9265,N_8269,N_6844);
and U9266 (N_9266,N_6665,N_7161);
nand U9267 (N_9267,N_6511,N_7708);
and U9268 (N_9268,N_7475,N_8435);
or U9269 (N_9269,N_8521,N_7814);
nor U9270 (N_9270,N_6781,N_7790);
nor U9271 (N_9271,N_6835,N_7118);
nor U9272 (N_9272,N_8781,N_6465);
or U9273 (N_9273,N_6010,N_8514);
or U9274 (N_9274,N_7864,N_7146);
nor U9275 (N_9275,N_6286,N_6698);
and U9276 (N_9276,N_7793,N_7726);
nand U9277 (N_9277,N_7347,N_8910);
nor U9278 (N_9278,N_8404,N_6355);
nor U9279 (N_9279,N_6484,N_6289);
or U9280 (N_9280,N_8884,N_6896);
xnor U9281 (N_9281,N_8300,N_7538);
and U9282 (N_9282,N_7226,N_8362);
nor U9283 (N_9283,N_6780,N_7633);
and U9284 (N_9284,N_6587,N_7206);
nor U9285 (N_9285,N_8704,N_7416);
nor U9286 (N_9286,N_6892,N_7879);
nand U9287 (N_9287,N_8171,N_6983);
nand U9288 (N_9288,N_6758,N_8624);
nand U9289 (N_9289,N_6794,N_7600);
and U9290 (N_9290,N_6415,N_6977);
and U9291 (N_9291,N_8465,N_6459);
nand U9292 (N_9292,N_8025,N_6412);
or U9293 (N_9293,N_6934,N_7182);
and U9294 (N_9294,N_8887,N_8257);
nand U9295 (N_9295,N_8013,N_8997);
or U9296 (N_9296,N_7317,N_6635);
or U9297 (N_9297,N_8170,N_6825);
and U9298 (N_9298,N_6233,N_7214);
nor U9299 (N_9299,N_8094,N_7422);
and U9300 (N_9300,N_7208,N_7867);
nand U9301 (N_9301,N_8621,N_8100);
or U9302 (N_9302,N_8667,N_6716);
nor U9303 (N_9303,N_7692,N_7737);
or U9304 (N_9304,N_6849,N_8674);
and U9305 (N_9305,N_6720,N_6054);
and U9306 (N_9306,N_8666,N_8483);
nor U9307 (N_9307,N_6941,N_7363);
nor U9308 (N_9308,N_8739,N_7032);
or U9309 (N_9309,N_6670,N_7337);
nor U9310 (N_9310,N_7678,N_7014);
or U9311 (N_9311,N_8188,N_6704);
and U9312 (N_9312,N_6246,N_7356);
nand U9313 (N_9313,N_8254,N_6987);
nor U9314 (N_9314,N_8610,N_8453);
and U9315 (N_9315,N_8055,N_7730);
or U9316 (N_9316,N_6928,N_8880);
nand U9317 (N_9317,N_7381,N_8046);
and U9318 (N_9318,N_8552,N_8782);
and U9319 (N_9319,N_8963,N_8488);
nand U9320 (N_9320,N_8378,N_6595);
or U9321 (N_9321,N_7329,N_7821);
nand U9322 (N_9322,N_7604,N_6095);
nand U9323 (N_9323,N_8840,N_8252);
nor U9324 (N_9324,N_6477,N_7786);
or U9325 (N_9325,N_6359,N_7372);
or U9326 (N_9326,N_8466,N_8545);
xnor U9327 (N_9327,N_7899,N_6805);
or U9328 (N_9328,N_8002,N_6699);
or U9329 (N_9329,N_7051,N_8856);
nand U9330 (N_9330,N_7419,N_6997);
and U9331 (N_9331,N_8675,N_6134);
nor U9332 (N_9332,N_7174,N_8942);
nor U9333 (N_9333,N_7693,N_7655);
or U9334 (N_9334,N_6165,N_8946);
nand U9335 (N_9335,N_6572,N_6864);
nand U9336 (N_9336,N_7277,N_7352);
nor U9337 (N_9337,N_6350,N_7152);
nand U9338 (N_9338,N_7495,N_8714);
nand U9339 (N_9339,N_6514,N_8791);
and U9340 (N_9340,N_8035,N_7642);
nor U9341 (N_9341,N_6167,N_6661);
xor U9342 (N_9342,N_8813,N_8003);
and U9343 (N_9343,N_7490,N_7195);
nand U9344 (N_9344,N_7929,N_7765);
nand U9345 (N_9345,N_8515,N_8315);
nor U9346 (N_9346,N_8523,N_6681);
nor U9347 (N_9347,N_8472,N_6086);
nand U9348 (N_9348,N_7636,N_8339);
nor U9349 (N_9349,N_8746,N_6345);
and U9350 (N_9350,N_6293,N_8152);
nand U9351 (N_9351,N_7333,N_8016);
and U9352 (N_9352,N_6806,N_8049);
and U9353 (N_9353,N_8900,N_6554);
and U9354 (N_9354,N_7153,N_8544);
nor U9355 (N_9355,N_8063,N_8352);
nand U9356 (N_9356,N_7532,N_7127);
nand U9357 (N_9357,N_6087,N_8644);
nor U9358 (N_9358,N_7075,N_7559);
and U9359 (N_9359,N_6796,N_6417);
and U9360 (N_9360,N_6750,N_7751);
and U9361 (N_9361,N_8295,N_7885);
nand U9362 (N_9362,N_7915,N_8668);
nand U9363 (N_9363,N_6473,N_7273);
and U9364 (N_9364,N_6685,N_7199);
and U9365 (N_9365,N_7940,N_6873);
nor U9366 (N_9366,N_7254,N_6013);
nor U9367 (N_9367,N_7717,N_8630);
or U9368 (N_9368,N_7048,N_6597);
nor U9369 (N_9369,N_7160,N_8274);
and U9370 (N_9370,N_7284,N_6564);
or U9371 (N_9371,N_8985,N_7541);
nor U9372 (N_9372,N_6102,N_7828);
and U9373 (N_9373,N_8661,N_8862);
nor U9374 (N_9374,N_8951,N_6408);
or U9375 (N_9375,N_6618,N_7129);
or U9376 (N_9376,N_6791,N_8175);
nand U9377 (N_9377,N_7811,N_7454);
nor U9378 (N_9378,N_7881,N_7686);
nand U9379 (N_9379,N_6533,N_7520);
and U9380 (N_9380,N_8400,N_7261);
or U9381 (N_9381,N_8085,N_6414);
xnor U9382 (N_9382,N_8012,N_6672);
and U9383 (N_9383,N_8297,N_6413);
nor U9384 (N_9384,N_8397,N_8369);
and U9385 (N_9385,N_7572,N_6940);
nand U9386 (N_9386,N_8984,N_8820);
or U9387 (N_9387,N_8771,N_8124);
nor U9388 (N_9388,N_6483,N_6136);
or U9389 (N_9389,N_8270,N_8860);
nor U9390 (N_9390,N_8147,N_7720);
or U9391 (N_9391,N_8752,N_8802);
or U9392 (N_9392,N_8916,N_7695);
nand U9393 (N_9393,N_8430,N_7219);
or U9394 (N_9394,N_7954,N_8145);
or U9395 (N_9395,N_6673,N_7280);
nor U9396 (N_9396,N_7232,N_6211);
and U9397 (N_9397,N_8394,N_8492);
nand U9398 (N_9398,N_7355,N_7950);
xor U9399 (N_9399,N_7427,N_8127);
nand U9400 (N_9400,N_6600,N_7121);
and U9401 (N_9401,N_7376,N_7016);
nor U9402 (N_9402,N_7090,N_6324);
or U9403 (N_9403,N_6031,N_6926);
or U9404 (N_9404,N_6999,N_8409);
and U9405 (N_9405,N_7902,N_6000);
and U9406 (N_9406,N_8535,N_8261);
nand U9407 (N_9407,N_7229,N_7898);
nand U9408 (N_9408,N_8144,N_7524);
or U9409 (N_9409,N_8660,N_7264);
and U9410 (N_9410,N_6649,N_8537);
nand U9411 (N_9411,N_8789,N_6881);
nor U9412 (N_9412,N_8564,N_8027);
nor U9413 (N_9413,N_6042,N_7783);
nor U9414 (N_9414,N_8897,N_6721);
nand U9415 (N_9415,N_6916,N_8160);
or U9416 (N_9416,N_8508,N_6216);
or U9417 (N_9417,N_6674,N_6985);
and U9418 (N_9418,N_7224,N_7933);
nor U9419 (N_9419,N_6494,N_8801);
and U9420 (N_9420,N_8209,N_7961);
nor U9421 (N_9421,N_6816,N_8375);
nand U9422 (N_9422,N_6932,N_7396);
nand U9423 (N_9423,N_8678,N_8592);
nand U9424 (N_9424,N_8550,N_6016);
nand U9425 (N_9425,N_7113,N_6219);
nand U9426 (N_9426,N_6651,N_8494);
nand U9427 (N_9427,N_6768,N_7038);
nor U9428 (N_9428,N_6298,N_8185);
nor U9429 (N_9429,N_8994,N_7723);
nor U9430 (N_9430,N_8993,N_6586);
and U9431 (N_9431,N_8506,N_6512);
or U9432 (N_9432,N_6443,N_8507);
or U9433 (N_9433,N_6374,N_7893);
xnor U9434 (N_9434,N_8236,N_6939);
nand U9435 (N_9435,N_8670,N_8417);
nor U9436 (N_9436,N_7216,N_8215);
nor U9437 (N_9437,N_6500,N_8286);
nand U9438 (N_9438,N_6428,N_8992);
nor U9439 (N_9439,N_8210,N_8342);
and U9440 (N_9440,N_7578,N_8543);
or U9441 (N_9441,N_8960,N_8475);
nor U9442 (N_9442,N_6387,N_6308);
and U9443 (N_9443,N_6377,N_8716);
nor U9444 (N_9444,N_6955,N_6666);
nor U9445 (N_9445,N_7418,N_7034);
nor U9446 (N_9446,N_7705,N_6541);
nand U9447 (N_9447,N_8845,N_8264);
nand U9448 (N_9448,N_6710,N_7564);
nor U9449 (N_9449,N_7012,N_6241);
or U9450 (N_9450,N_8165,N_7934);
nand U9451 (N_9451,N_7551,N_7834);
or U9452 (N_9452,N_6606,N_7228);
and U9453 (N_9453,N_8619,N_6482);
nor U9454 (N_9454,N_6552,N_8444);
nand U9455 (N_9455,N_7470,N_7637);
and U9456 (N_9456,N_8357,N_8449);
nor U9457 (N_9457,N_7769,N_8635);
and U9458 (N_9458,N_8891,N_7230);
nor U9459 (N_9459,N_8811,N_7288);
or U9460 (N_9460,N_8099,N_6487);
or U9461 (N_9461,N_7184,N_7627);
or U9462 (N_9462,N_6066,N_8605);
or U9463 (N_9463,N_8275,N_7863);
nor U9464 (N_9464,N_6826,N_6237);
nand U9465 (N_9465,N_8866,N_8534);
and U9466 (N_9466,N_7838,N_7165);
or U9467 (N_9467,N_7622,N_6127);
nor U9468 (N_9468,N_6015,N_8211);
or U9469 (N_9469,N_6588,N_8030);
nor U9470 (N_9470,N_7620,N_6603);
nand U9471 (N_9471,N_7447,N_8087);
nand U9472 (N_9472,N_8664,N_8593);
nand U9473 (N_9473,N_8899,N_6027);
nand U9474 (N_9474,N_6495,N_7675);
or U9475 (N_9475,N_6613,N_6208);
nand U9476 (N_9476,N_7200,N_7379);
or U9477 (N_9477,N_7238,N_6757);
and U9478 (N_9478,N_7428,N_8918);
or U9479 (N_9479,N_6179,N_7758);
and U9480 (N_9480,N_7772,N_8563);
nor U9481 (N_9481,N_7159,N_6173);
nand U9482 (N_9482,N_7164,N_7682);
nor U9483 (N_9483,N_6852,N_6614);
or U9484 (N_9484,N_6416,N_6936);
nor U9485 (N_9485,N_6906,N_6437);
and U9486 (N_9486,N_7649,N_6637);
nor U9487 (N_9487,N_7132,N_8198);
and U9488 (N_9488,N_8387,N_7054);
nand U9489 (N_9489,N_8979,N_6492);
nor U9490 (N_9490,N_6480,N_8518);
nand U9491 (N_9491,N_8388,N_6829);
or U9492 (N_9492,N_7605,N_6214);
nand U9493 (N_9493,N_6561,N_6607);
nand U9494 (N_9494,N_6441,N_6344);
nor U9495 (N_9495,N_7819,N_6745);
and U9496 (N_9496,N_6633,N_6429);
nor U9497 (N_9497,N_6438,N_6074);
or U9498 (N_9498,N_8428,N_7210);
nand U9499 (N_9499,N_6161,N_6591);
nand U9500 (N_9500,N_8478,N_6700);
or U9501 (N_9501,N_7852,N_7925);
nor U9502 (N_9502,N_6148,N_6341);
nor U9503 (N_9503,N_7117,N_6529);
and U9504 (N_9504,N_8859,N_8065);
nand U9505 (N_9505,N_6307,N_7496);
and U9506 (N_9506,N_8745,N_7062);
nand U9507 (N_9507,N_6435,N_6693);
xnor U9508 (N_9508,N_6809,N_7894);
and U9509 (N_9509,N_6824,N_8214);
and U9510 (N_9510,N_6204,N_6579);
nor U9511 (N_9511,N_8873,N_8473);
and U9512 (N_9512,N_6122,N_6760);
nand U9513 (N_9513,N_7217,N_8712);
nand U9514 (N_9514,N_8927,N_7691);
nand U9515 (N_9515,N_8096,N_6737);
nand U9516 (N_9516,N_8513,N_6654);
and U9517 (N_9517,N_8343,N_6566);
and U9518 (N_9518,N_8561,N_8961);
nand U9519 (N_9519,N_7289,N_8560);
nor U9520 (N_9520,N_6543,N_7348);
nand U9521 (N_9521,N_6118,N_6068);
or U9522 (N_9522,N_7619,N_7088);
nor U9523 (N_9523,N_8045,N_7569);
or U9524 (N_9524,N_8885,N_8415);
nand U9525 (N_9525,N_6778,N_7526);
and U9526 (N_9526,N_7752,N_7533);
nor U9527 (N_9527,N_7143,N_6052);
nor U9528 (N_9528,N_8406,N_6990);
or U9529 (N_9529,N_6425,N_6813);
nor U9530 (N_9530,N_6269,N_7544);
or U9531 (N_9531,N_7369,N_6059);
or U9532 (N_9532,N_6498,N_6185);
or U9533 (N_9533,N_7548,N_8420);
nor U9534 (N_9534,N_7853,N_7517);
nor U9535 (N_9535,N_8652,N_7711);
nor U9536 (N_9536,N_6988,N_6872);
nand U9537 (N_9537,N_7188,N_8848);
nand U9538 (N_9538,N_7718,N_8489);
and U9539 (N_9539,N_7017,N_7385);
and U9540 (N_9540,N_8784,N_6647);
and U9541 (N_9541,N_6880,N_7714);
nor U9542 (N_9542,N_8640,N_7698);
nor U9543 (N_9543,N_8161,N_8468);
nor U9544 (N_9544,N_6199,N_7500);
or U9545 (N_9545,N_7137,N_6516);
nand U9546 (N_9546,N_7917,N_6335);
or U9547 (N_9547,N_6076,N_6021);
or U9548 (N_9548,N_6200,N_7023);
nand U9549 (N_9549,N_6444,N_8501);
and U9550 (N_9550,N_8011,N_7259);
or U9551 (N_9551,N_7877,N_7983);
nor U9552 (N_9552,N_8834,N_7312);
and U9553 (N_9553,N_7768,N_7802);
nand U9554 (N_9554,N_8287,N_6921);
and U9555 (N_9555,N_8718,N_8422);
nand U9556 (N_9556,N_7292,N_8493);
and U9557 (N_9557,N_8177,N_6090);
and U9558 (N_9558,N_8071,N_6316);
nor U9559 (N_9559,N_6128,N_6845);
nor U9560 (N_9560,N_8355,N_7343);
nand U9561 (N_9561,N_7389,N_6446);
nand U9562 (N_9562,N_8562,N_7350);
or U9563 (N_9563,N_8740,N_8335);
nor U9564 (N_9564,N_8839,N_8340);
nand U9565 (N_9565,N_6902,N_6206);
nor U9566 (N_9566,N_6318,N_7450);
nor U9567 (N_9567,N_8722,N_8367);
nor U9568 (N_9568,N_6914,N_8869);
nand U9569 (N_9569,N_6235,N_8677);
nand U9570 (N_9570,N_8982,N_8547);
nor U9571 (N_9571,N_7364,N_8909);
nor U9572 (N_9572,N_7212,N_7144);
and U9573 (N_9573,N_7257,N_7736);
nor U9574 (N_9574,N_7402,N_8058);
nor U9575 (N_9575,N_6466,N_8148);
nand U9576 (N_9576,N_6574,N_7995);
nor U9577 (N_9577,N_6527,N_8296);
or U9578 (N_9578,N_7358,N_6295);
and U9579 (N_9579,N_6832,N_8212);
or U9580 (N_9580,N_8345,N_8135);
nor U9581 (N_9581,N_7721,N_7805);
nand U9582 (N_9582,N_8251,N_6142);
or U9583 (N_9583,N_8853,N_6638);
nor U9584 (N_9584,N_7064,N_8246);
nor U9585 (N_9585,N_7362,N_6149);
and U9586 (N_9586,N_7901,N_6460);
or U9587 (N_9587,N_6276,N_7448);
or U9588 (N_9588,N_7781,N_6634);
xnor U9589 (N_9589,N_7241,N_7777);
nand U9590 (N_9590,N_7299,N_8996);
nor U9591 (N_9591,N_8978,N_7606);
or U9592 (N_9592,N_6718,N_8376);
nand U9593 (N_9593,N_6759,N_7497);
nor U9594 (N_9594,N_8447,N_8366);
and U9595 (N_9595,N_7468,N_6585);
or U9596 (N_9596,N_8078,N_8186);
and U9597 (N_9597,N_6676,N_8169);
or U9598 (N_9598,N_7628,N_8328);
or U9599 (N_9599,N_7712,N_8804);
and U9600 (N_9600,N_6402,N_8645);
nor U9601 (N_9601,N_7788,N_6020);
or U9602 (N_9602,N_6798,N_7984);
and U9603 (N_9603,N_7795,N_7357);
and U9604 (N_9604,N_7086,N_7022);
or U9605 (N_9605,N_6584,N_6272);
or U9606 (N_9606,N_7209,N_6507);
and U9607 (N_9607,N_8973,N_7865);
nand U9608 (N_9608,N_6968,N_7082);
or U9609 (N_9609,N_8944,N_6119);
or U9610 (N_9610,N_7573,N_8026);
nor U9611 (N_9611,N_7666,N_7749);
or U9612 (N_9612,N_7680,N_7952);
nor U9613 (N_9613,N_7015,N_6751);
or U9614 (N_9614,N_6065,N_6255);
and U9615 (N_9615,N_7305,N_7002);
xor U9616 (N_9616,N_8571,N_8617);
or U9617 (N_9617,N_8917,N_7803);
or U9618 (N_9618,N_7778,N_7141);
and U9619 (N_9619,N_6310,N_8075);
nor U9620 (N_9620,N_8391,N_6559);
or U9621 (N_9621,N_7316,N_7800);
or U9622 (N_9622,N_7755,N_7888);
or U9623 (N_9623,N_6445,N_6688);
xnor U9624 (N_9624,N_7401,N_6653);
and U9625 (N_9625,N_8625,N_7150);
nor U9626 (N_9626,N_6989,N_6581);
nand U9627 (N_9627,N_7262,N_8037);
nand U9628 (N_9628,N_7459,N_7530);
nor U9629 (N_9629,N_6014,N_7325);
nor U9630 (N_9630,N_6510,N_6278);
nor U9631 (N_9631,N_8904,N_7194);
and U9632 (N_9632,N_6256,N_8603);
nand U9633 (N_9633,N_6440,N_8048);
or U9634 (N_9634,N_6436,N_7773);
nand U9635 (N_9635,N_7504,N_8669);
nor U9636 (N_9636,N_8208,N_8309);
and U9637 (N_9637,N_6722,N_7026);
nor U9638 (N_9638,N_7084,N_6008);
nand U9639 (N_9639,N_6184,N_6882);
or U9640 (N_9640,N_7546,N_6629);
nand U9641 (N_9641,N_6088,N_8233);
and U9642 (N_9642,N_6125,N_7999);
nand U9643 (N_9643,N_6624,N_6292);
nor U9644 (N_9644,N_7240,N_8197);
or U9645 (N_9645,N_6120,N_7058);
and U9646 (N_9646,N_7172,N_8240);
nand U9647 (N_9647,N_8754,N_6041);
and U9648 (N_9648,N_8381,N_7351);
or U9649 (N_9649,N_6369,N_8599);
or U9650 (N_9650,N_6546,N_8647);
or U9651 (N_9651,N_8158,N_8110);
or U9652 (N_9652,N_7932,N_7908);
nand U9653 (N_9653,N_6080,N_8818);
or U9654 (N_9654,N_7473,N_6942);
or U9655 (N_9655,N_6296,N_6970);
or U9656 (N_9656,N_8768,N_8450);
and U9657 (N_9657,N_6056,N_8600);
nand U9658 (N_9658,N_8089,N_7331);
or U9659 (N_9659,N_8195,N_8596);
and U9660 (N_9660,N_6196,N_8427);
or U9661 (N_9661,N_6124,N_6129);
nand U9662 (N_9662,N_8258,N_6888);
nor U9663 (N_9663,N_7906,N_7285);
and U9664 (N_9664,N_8143,N_7651);
or U9665 (N_9665,N_6221,N_8685);
nand U9666 (N_9666,N_6713,N_6363);
and U9667 (N_9667,N_7027,N_6002);
and U9668 (N_9668,N_8765,N_6001);
nand U9669 (N_9669,N_8082,N_6147);
nor U9670 (N_9670,N_7110,N_8412);
or U9671 (N_9671,N_6283,N_6594);
or U9672 (N_9672,N_7035,N_6617);
nand U9673 (N_9673,N_6717,N_6389);
nand U9674 (N_9674,N_6046,N_6180);
or U9675 (N_9675,N_6508,N_7644);
or U9676 (N_9676,N_7635,N_6409);
and U9677 (N_9677,N_6394,N_7895);
or U9678 (N_9678,N_7179,N_6708);
or U9679 (N_9679,N_7816,N_7033);
or U9680 (N_9680,N_7077,N_7561);
and U9681 (N_9681,N_7919,N_8044);
nand U9682 (N_9682,N_6485,N_7846);
nor U9683 (N_9683,N_7839,N_7242);
nand U9684 (N_9684,N_6150,N_7089);
nor U9685 (N_9685,N_7298,N_8206);
nor U9686 (N_9686,N_6730,N_7761);
and U9687 (N_9687,N_7976,N_8363);
nor U9688 (N_9688,N_8792,N_7310);
and U9689 (N_9689,N_7480,N_8064);
and U9690 (N_9690,N_6958,N_7641);
and U9691 (N_9691,N_7093,N_8199);
and U9692 (N_9692,N_7097,N_6763);
or U9693 (N_9693,N_7166,N_7847);
or U9694 (N_9694,N_7125,N_7102);
nand U9695 (N_9695,N_6406,N_6348);
or U9696 (N_9696,N_7103,N_7303);
and U9697 (N_9697,N_8460,N_6777);
or U9698 (N_9698,N_7630,N_8348);
or U9699 (N_9699,N_8731,N_6135);
or U9700 (N_9700,N_7937,N_6290);
and U9701 (N_9701,N_6857,N_6232);
nor U9702 (N_9702,N_6462,N_7104);
nor U9703 (N_9703,N_7122,N_8154);
and U9704 (N_9704,N_8586,N_7685);
nor U9705 (N_9705,N_8542,N_7716);
nor U9706 (N_9706,N_6447,N_6924);
nor U9707 (N_9707,N_6434,N_6334);
and U9708 (N_9708,N_7313,N_8032);
nor U9709 (N_9709,N_6615,N_8744);
nand U9710 (N_9710,N_8911,N_8687);
and U9711 (N_9711,N_7263,N_8414);
nand U9712 (N_9712,N_7412,N_8696);
and U9713 (N_9713,N_8580,N_8182);
nand U9714 (N_9714,N_8665,N_8324);
or U9715 (N_9715,N_7031,N_8426);
or U9716 (N_9716,N_6168,N_8954);
nor U9717 (N_9717,N_7658,N_7085);
nor U9718 (N_9718,N_6937,N_8043);
nand U9719 (N_9719,N_8548,N_8380);
nand U9720 (N_9720,N_7905,N_7713);
nor U9721 (N_9721,N_7939,N_6250);
or U9722 (N_9722,N_8576,N_7671);
nand U9723 (N_9723,N_7754,N_7311);
and U9724 (N_9724,N_7876,N_8053);
or U9725 (N_9725,N_8924,N_6724);
nor U9726 (N_9726,N_6427,N_7892);
nor U9727 (N_9727,N_7664,N_8298);
nor U9728 (N_9728,N_6682,N_7341);
xnor U9729 (N_9729,N_7063,N_8577);
nand U9730 (N_9730,N_7522,N_8060);
nand U9731 (N_9731,N_6899,N_8868);
nor U9732 (N_9732,N_7903,N_7281);
and U9733 (N_9733,N_6668,N_7502);
nor U9734 (N_9734,N_6911,N_7866);
or U9735 (N_9735,N_6371,N_7602);
nand U9736 (N_9736,N_7771,N_6764);
or U9737 (N_9737,N_6105,N_6625);
nand U9738 (N_9738,N_8762,N_7610);
nand U9739 (N_9739,N_8173,N_6163);
and U9740 (N_9740,N_8495,N_6039);
and U9741 (N_9741,N_8023,N_6866);
nand U9742 (N_9742,N_6097,N_8608);
nor U9743 (N_9743,N_7467,N_8120);
nand U9744 (N_9744,N_8057,N_6626);
nor U9745 (N_9745,N_6222,N_8557);
or U9746 (N_9746,N_6174,N_7962);
or U9747 (N_9747,N_7804,N_7001);
and U9748 (N_9748,N_6252,N_6696);
and U9749 (N_9749,N_7171,N_6030);
nor U9750 (N_9750,N_8823,N_8360);
nand U9751 (N_9751,N_7061,N_8612);
nand U9752 (N_9752,N_8456,N_8772);
nand U9753 (N_9753,N_7799,N_7202);
or U9754 (N_9754,N_7393,N_7207);
and U9755 (N_9755,N_8737,N_7910);
nor U9756 (N_9756,N_7030,N_6420);
nor U9757 (N_9757,N_6562,N_6938);
or U9758 (N_9758,N_7941,N_7463);
and U9759 (N_9759,N_8953,N_7167);
nand U9760 (N_9760,N_8788,N_7767);
or U9761 (N_9761,N_8019,N_8549);
nor U9762 (N_9762,N_7825,N_6130);
nor U9763 (N_9763,N_7435,N_8952);
nand U9764 (N_9764,N_7965,N_6839);
or U9765 (N_9765,N_7590,N_8256);
nand U9766 (N_9766,N_7233,N_6576);
nand U9767 (N_9767,N_7101,N_8267);
nand U9768 (N_9768,N_6962,N_8079);
nand U9769 (N_9769,N_6657,N_8747);
and U9770 (N_9770,N_8968,N_7286);
nor U9771 (N_9771,N_7886,N_8227);
and U9772 (N_9772,N_6110,N_8611);
nor U9773 (N_9773,N_7744,N_8326);
or U9774 (N_9774,N_6433,N_6522);
nor U9775 (N_9775,N_8588,N_6193);
nor U9776 (N_9776,N_6592,N_7072);
nor U9777 (N_9777,N_8572,N_6840);
or U9778 (N_9778,N_8077,N_6948);
nor U9779 (N_9779,N_7963,N_6506);
nand U9780 (N_9780,N_6537,N_7078);
nand U9781 (N_9781,N_7996,N_6164);
or U9782 (N_9782,N_8581,N_7986);
and U9783 (N_9783,N_7335,N_6159);
nand U9784 (N_9784,N_8928,N_6905);
nor U9785 (N_9785,N_6943,N_6741);
or U9786 (N_9786,N_8948,N_6166);
and U9787 (N_9787,N_6104,N_8833);
and U9788 (N_9788,N_6890,N_8972);
and U9789 (N_9789,N_8168,N_7487);
and U9790 (N_9790,N_8156,N_8390);
nand U9791 (N_9791,N_8132,N_8009);
or U9792 (N_9792,N_8584,N_6876);
and U9793 (N_9793,N_7431,N_8894);
or U9794 (N_9794,N_7437,N_6524);
or U9795 (N_9795,N_7815,N_6802);
or U9796 (N_9796,N_6797,N_8282);
nand U9797 (N_9797,N_6599,N_7654);
or U9798 (N_9798,N_8330,N_7092);
nor U9799 (N_9799,N_6867,N_7922);
nor U9800 (N_9800,N_8850,N_7715);
or U9801 (N_9801,N_7486,N_8107);
nor U9802 (N_9802,N_8263,N_6927);
or U9803 (N_9803,N_8238,N_6284);
nand U9804 (N_9804,N_6842,N_7266);
nor U9805 (N_9805,N_8086,N_6337);
nor U9806 (N_9806,N_8816,N_7539);
and U9807 (N_9807,N_8440,N_6605);
or U9808 (N_9808,N_7774,N_7883);
nor U9809 (N_9809,N_7321,N_8590);
and U9810 (N_9810,N_6338,N_8680);
nor U9811 (N_9811,N_7920,N_7469);
nor U9812 (N_9812,N_8730,N_7914);
nand U9813 (N_9813,N_7734,N_8715);
and U9814 (N_9814,N_7762,N_8101);
or U9815 (N_9815,N_6114,N_8812);
nor U9816 (N_9816,N_8583,N_6432);
or U9817 (N_9817,N_6736,N_6113);
nor U9818 (N_9818,N_6553,N_8957);
or U9819 (N_9819,N_6556,N_7971);
nand U9820 (N_9820,N_6982,N_6053);
nor U9821 (N_9821,N_8436,N_7301);
nand U9822 (N_9822,N_7873,N_8569);
or U9823 (N_9823,N_7706,N_8926);
nand U9824 (N_9824,N_8729,N_8216);
and U9825 (N_9825,N_7112,N_6254);
xor U9826 (N_9826,N_7747,N_7008);
and U9827 (N_9827,N_8401,N_6470);
and U9828 (N_9828,N_6285,N_6258);
nand U9829 (N_9829,N_6858,N_6789);
or U9830 (N_9830,N_6038,N_6570);
or U9831 (N_9831,N_7249,N_6979);
nor U9832 (N_9832,N_8874,N_8764);
nand U9833 (N_9833,N_7683,N_6464);
nand U9834 (N_9834,N_8266,N_7585);
nand U9835 (N_9835,N_8949,N_7413);
or U9836 (N_9836,N_6399,N_8329);
or U9837 (N_9837,N_7408,N_7045);
or U9838 (N_9838,N_6558,N_7410);
xor U9839 (N_9839,N_7624,N_6287);
and U9840 (N_9840,N_6836,N_8201);
nor U9841 (N_9841,N_8181,N_8725);
or U9842 (N_9842,N_7087,N_7826);
nor U9843 (N_9843,N_6675,N_8606);
nand U9844 (N_9844,N_6215,N_7052);
nand U9845 (N_9845,N_8527,N_8852);
or U9846 (N_9846,N_7056,N_6766);
nor U9847 (N_9847,N_8389,N_7123);
and U9848 (N_9848,N_7823,N_6819);
or U9849 (N_9849,N_6454,N_8975);
nor U9850 (N_9850,N_8217,N_7968);
nand U9851 (N_9851,N_8826,N_8424);
nor U9852 (N_9852,N_6111,N_7294);
and U9853 (N_9853,N_7878,N_7861);
and U9854 (N_9854,N_8068,N_7411);
nor U9855 (N_9855,N_7979,N_8429);
nand U9856 (N_9856,N_8062,N_6642);
and U9857 (N_9857,N_8533,N_6358);
nand U9858 (N_9858,N_7057,N_7519);
nand U9859 (N_9859,N_8903,N_6868);
nor U9860 (N_9860,N_6612,N_7386);
nor U9861 (N_9861,N_6565,N_8125);
nor U9862 (N_9862,N_7601,N_7227);
nand U9863 (N_9863,N_7483,N_7926);
nor U9864 (N_9864,N_7456,N_8706);
nand U9865 (N_9865,N_6862,N_7936);
or U9866 (N_9866,N_6683,N_8502);
nor U9867 (N_9867,N_7668,N_8108);
and U9868 (N_9868,N_6856,N_7059);
or U9869 (N_9869,N_7924,N_6188);
nor U9870 (N_9870,N_8073,N_8196);
and U9871 (N_9871,N_8106,N_7269);
nand U9872 (N_9872,N_8734,N_7964);
nand U9873 (N_9873,N_6035,N_7608);
or U9874 (N_9874,N_6518,N_8123);
nand U9875 (N_9875,N_6055,N_7494);
nand U9876 (N_9876,N_8480,N_6160);
or U9877 (N_9877,N_8056,N_8753);
nand U9878 (N_9878,N_7003,N_7887);
or U9879 (N_9879,N_7201,N_6782);
nor U9880 (N_9880,N_7791,N_7451);
or U9881 (N_9881,N_6644,N_7536);
or U9882 (N_9882,N_6123,N_6153);
nor U9883 (N_9883,N_6242,N_8316);
nand U9884 (N_9884,N_7732,N_7942);
or U9885 (N_9885,N_7115,N_8280);
or U9886 (N_9886,N_8116,N_6079);
nand U9887 (N_9887,N_7987,N_6458);
or U9888 (N_9888,N_6012,N_6315);
and U9889 (N_9889,N_6677,N_6678);
nand U9890 (N_9890,N_8464,N_7997);
nand U9891 (N_9891,N_8469,N_7189);
or U9892 (N_9892,N_7139,N_6263);
nand U9893 (N_9893,N_7420,N_6850);
nor U9894 (N_9894,N_6397,N_8416);
or U9895 (N_9895,N_7445,N_7935);
or U9896 (N_9896,N_7256,N_6396);
nand U9897 (N_9897,N_7975,N_8244);
and U9898 (N_9898,N_6202,N_8613);
or U9899 (N_9899,N_6593,N_7236);
nand U9900 (N_9900,N_7947,N_8248);
nand U9901 (N_9901,N_8679,N_7302);
nand U9902 (N_9902,N_6893,N_6680);
nand U9903 (N_9903,N_8878,N_6061);
or U9904 (N_9904,N_7255,N_8092);
nand U9905 (N_9905,N_6870,N_6140);
nor U9906 (N_9906,N_6267,N_7810);
or U9907 (N_9907,N_8691,N_7969);
and U9908 (N_9908,N_6538,N_6930);
nor U9909 (N_9909,N_8499,N_7168);
nand U9910 (N_9910,N_7073,N_8795);
nand U9911 (N_9911,N_6367,N_6769);
or U9912 (N_9912,N_7275,N_8692);
nand U9913 (N_9913,N_8827,N_8934);
or U9914 (N_9914,N_7534,N_6329);
nor U9915 (N_9915,N_8467,N_7258);
nor U9916 (N_9916,N_8755,N_8083);
nor U9917 (N_9917,N_8831,N_7900);
nand U9918 (N_9918,N_8935,N_7854);
nor U9919 (N_9919,N_8607,N_6733);
or U9920 (N_9920,N_8481,N_6234);
nand U9921 (N_9921,N_6608,N_8922);
and U9922 (N_9922,N_7687,N_7120);
or U9923 (N_9923,N_6577,N_8098);
nor U9924 (N_9924,N_7323,N_8008);
or U9925 (N_9925,N_7004,N_6325);
or U9926 (N_9926,N_6342,N_6251);
nand U9927 (N_9927,N_6071,N_7576);
or U9928 (N_9928,N_7623,N_6029);
nor U9929 (N_9929,N_8604,N_8541);
nor U9930 (N_9930,N_8653,N_7060);
nand U9931 (N_9931,N_7946,N_6646);
nand U9932 (N_9932,N_8969,N_8301);
or U9933 (N_9933,N_6658,N_7897);
nand U9934 (N_9934,N_6182,N_6784);
and U9935 (N_9935,N_7272,N_7414);
nand U9936 (N_9936,N_8137,N_7221);
or U9937 (N_9937,N_7234,N_6203);
nand U9938 (N_9938,N_7007,N_8490);
xor U9939 (N_9939,N_6489,N_8374);
nor U9940 (N_9940,N_6419,N_8383);
nor U9941 (N_9941,N_7049,N_8150);
nand U9942 (N_9942,N_8637,N_7738);
nor U9943 (N_9943,N_7000,N_8038);
or U9944 (N_9944,N_6742,N_7278);
or U9945 (N_9945,N_6382,N_7079);
and U9946 (N_9946,N_6373,N_8530);
nor U9947 (N_9947,N_6525,N_7471);
or U9948 (N_9948,N_8881,N_7529);
or U9949 (N_9949,N_6848,N_6175);
nand U9950 (N_9950,N_8402,N_7457);
nand U9951 (N_9951,N_8786,N_8200);
and U9952 (N_9952,N_7099,N_7156);
or U9953 (N_9953,N_8344,N_7560);
or U9954 (N_9954,N_7297,N_6689);
nand U9955 (N_9955,N_7400,N_7138);
or U9956 (N_9956,N_8114,N_6540);
nor U9957 (N_9957,N_8439,N_8836);
or U9958 (N_9958,N_8015,N_8656);
or U9959 (N_9959,N_8293,N_8940);
nor U9960 (N_9960,N_7306,N_8695);
and U9961 (N_9961,N_7586,N_8882);
or U9962 (N_9962,N_7991,N_7114);
nand U9963 (N_9963,N_8767,N_6695);
nor U9964 (N_9964,N_8779,N_6491);
nor U9965 (N_9965,N_6978,N_7868);
nor U9966 (N_9966,N_6410,N_8235);
and U9967 (N_9967,N_8259,N_6311);
nand U9968 (N_9968,N_6567,N_7377);
nand U9969 (N_9969,N_7743,N_6555);
nor U9970 (N_9970,N_8636,N_6513);
or U9971 (N_9971,N_8642,N_6669);
or U9972 (N_9972,N_8410,N_8620);
nor U9973 (N_9973,N_6170,N_8437);
nor U9974 (N_9974,N_7699,N_7594);
nor U9975 (N_9975,N_8566,N_7612);
or U9976 (N_9976,N_8776,N_6996);
nand U9977 (N_9977,N_6472,N_6947);
nand U9978 (N_9978,N_6557,N_7438);
or U9979 (N_9979,N_6229,N_7488);
and U9980 (N_9980,N_6309,N_8136);
or U9981 (N_9981,N_6424,N_7404);
or U9982 (N_9982,N_6515,N_7858);
and U9983 (N_9983,N_8277,N_7545);
and U9984 (N_9984,N_6051,N_8890);
nand U9985 (N_9985,N_7453,N_8841);
nand U9986 (N_9986,N_6209,N_8260);
nand U9987 (N_9987,N_7426,N_8815);
nor U9988 (N_9988,N_6503,N_8654);
and U9989 (N_9989,N_8766,N_7009);
nor U9990 (N_9990,N_8719,N_8006);
nand U9991 (N_9991,N_7896,N_6262);
nor U9992 (N_9992,N_6155,N_8112);
or U9993 (N_9993,N_8021,N_8932);
nor U9994 (N_9994,N_6991,N_7394);
nor U9995 (N_9995,N_6083,N_6563);
or U9996 (N_9996,N_6831,N_6746);
or U9997 (N_9997,N_8486,N_7587);
nor U9998 (N_9998,N_6322,N_6974);
nand U9999 (N_9999,N_8054,N_8938);
nor U10000 (N_10000,N_8338,N_6456);
nor U10001 (N_10001,N_7010,N_8104);
and U10002 (N_10002,N_7798,N_6171);
nand U10003 (N_10003,N_6081,N_8671);
and U10004 (N_10004,N_8423,N_7918);
nand U10005 (N_10005,N_8756,N_6773);
and U10006 (N_10006,N_6064,N_8694);
and U10007 (N_10007,N_8742,N_7069);
and U10008 (N_10008,N_6749,N_6475);
nand U10009 (N_10009,N_6004,N_6788);
nor U10010 (N_10010,N_7831,N_7290);
or U10011 (N_10011,N_6317,N_8822);
and U10012 (N_10012,N_7472,N_7346);
or U10013 (N_10013,N_8861,N_8031);
and U10014 (N_10014,N_6388,N_8837);
nand U10015 (N_10015,N_8307,N_6838);
and U10016 (N_10016,N_8162,N_7549);
and U10017 (N_10017,N_8284,N_6735);
and U10018 (N_10018,N_7913,N_8743);
or U10019 (N_10019,N_6535,N_7515);
or U10020 (N_10020,N_7595,N_6627);
nor U10021 (N_10021,N_8512,N_7591);
or U10022 (N_10022,N_7998,N_8322);
xnor U10023 (N_10023,N_8180,N_7353);
nand U10024 (N_10024,N_6172,N_8921);
and U10025 (N_10025,N_7907,N_6421);
and U10026 (N_10026,N_7944,N_6811);
xor U10027 (N_10027,N_7444,N_6620);
and U10028 (N_10028,N_7244,N_8317);
nor U10029 (N_10029,N_7181,N_8790);
nand U10030 (N_10030,N_8018,N_8875);
or U10031 (N_10031,N_6305,N_7053);
nand U10032 (N_10032,N_8672,N_6401);
or U10033 (N_10033,N_7724,N_8262);
and U10034 (N_10034,N_8690,N_6040);
and U10035 (N_10035,N_7722,N_8585);
nor U10036 (N_10036,N_7835,N_6351);
nand U10037 (N_10037,N_7066,N_6550);
or U10038 (N_10038,N_6257,N_8159);
and U10039 (N_10039,N_6547,N_8445);
nor U10040 (N_10040,N_6092,N_8998);
and U10041 (N_10041,N_7994,N_7041);
and U10042 (N_10042,N_8272,N_7856);
and U10043 (N_10043,N_8516,N_6018);
and U10044 (N_10044,N_7978,N_7753);
nand U10045 (N_10045,N_8760,N_6754);
or U10046 (N_10046,N_6622,N_7417);
nand U10047 (N_10047,N_8713,N_7916);
nand U10048 (N_10048,N_8770,N_8471);
or U10049 (N_10049,N_7304,N_7360);
or U10050 (N_10050,N_7439,N_6225);
nand U10051 (N_10051,N_8796,N_8222);
nor U10052 (N_10052,N_8245,N_7688);
or U10053 (N_10053,N_6861,N_6869);
or U10054 (N_10054,N_7523,N_7246);
or U10055 (N_10055,N_7748,N_8109);
and U10056 (N_10056,N_7672,N_6009);
or U10057 (N_10057,N_6821,N_8097);
and U10058 (N_10058,N_7833,N_7739);
nor U10059 (N_10059,N_6326,N_6240);
nand U10060 (N_10060,N_7039,N_8682);
or U10061 (N_10061,N_7047,N_6946);
nand U10062 (N_10062,N_7287,N_6384);
nor U10063 (N_10063,N_6479,N_6623);
nor U10064 (N_10064,N_8735,N_7931);
or U10065 (N_10065,N_6659,N_6400);
and U10066 (N_10066,N_6660,N_6108);
or U10067 (N_10067,N_8524,N_8650);
nand U10068 (N_10068,N_6692,N_7625);
nor U10069 (N_10069,N_6596,N_6772);
or U10070 (N_10070,N_8224,N_8128);
nor U10071 (N_10071,N_8399,N_8225);
nand U10072 (N_10072,N_8923,N_7516);
nor U10073 (N_10073,N_8649,N_7492);
and U10074 (N_10074,N_7220,N_8080);
nor U10075 (N_10075,N_8871,N_6431);
nor U10076 (N_10076,N_7733,N_6779);
or U10077 (N_10077,N_6321,N_6469);
or U10078 (N_10078,N_6404,N_8028);
or U10079 (N_10079,N_8396,N_7553);
and U10080 (N_10080,N_6523,N_7326);
nor U10081 (N_10081,N_8372,N_7318);
nand U10082 (N_10082,N_8091,N_7912);
and U10083 (N_10083,N_7293,N_6519);
and U10084 (N_10084,N_6509,N_8292);
nor U10085 (N_10085,N_8663,N_7977);
and U10086 (N_10086,N_6368,N_6874);
nand U10087 (N_10087,N_8040,N_8639);
nor U10088 (N_10088,N_6115,N_8203);
nand U10089 (N_10089,N_6705,N_6664);
nor U10090 (N_10090,N_8482,N_6210);
nand U10091 (N_10091,N_8321,N_6093);
or U10092 (N_10092,N_7959,N_6422);
nor U10093 (N_10093,N_6488,N_8785);
nand U10094 (N_10094,N_8609,N_7985);
nand U10095 (N_10095,N_7037,N_8888);
nor U10096 (N_10096,N_6744,N_7527);
and U10097 (N_10097,N_7499,N_7374);
nor U10098 (N_10098,N_8697,N_8628);
nand U10099 (N_10099,N_8559,N_8001);
nor U10100 (N_10100,N_8551,N_7684);
nor U10101 (N_10101,N_6922,N_8689);
and U10102 (N_10102,N_7235,N_8646);
nand U10103 (N_10103,N_7745,N_7191);
nor U10104 (N_10104,N_8627,N_7175);
nor U10105 (N_10105,N_8229,N_8913);
and U10106 (N_10106,N_8155,N_6352);
and U10107 (N_10107,N_7481,N_8022);
and U10108 (N_10108,N_6265,N_8708);
and U10109 (N_10109,N_7149,N_8937);
nor U10110 (N_10110,N_7848,N_7349);
nor U10111 (N_10111,N_6935,N_7328);
nor U10112 (N_10112,N_6006,N_7829);
or U10113 (N_10113,N_8458,N_6270);
or U10114 (N_10114,N_8452,N_8000);
or U10115 (N_10115,N_8965,N_6834);
or U10116 (N_10116,N_6965,N_7681);
nand U10117 (N_10117,N_7197,N_7845);
nand U10118 (N_10118,N_8565,N_7507);
and U10119 (N_10119,N_8867,N_6022);
nand U10120 (N_10120,N_6145,N_8632);
nor U10121 (N_10121,N_8291,N_8877);
or U10122 (N_10122,N_8582,N_8337);
and U10123 (N_10123,N_7268,N_6714);
or U10124 (N_10124,N_7131,N_7949);
or U10125 (N_10125,N_8829,N_7332);
nand U10126 (N_10126,N_8828,N_6756);
and U10127 (N_10127,N_6931,N_8769);
and U10128 (N_10128,N_6898,N_8294);
or U10129 (N_10129,N_7760,N_8648);
nor U10130 (N_10130,N_7021,N_6297);
and U10131 (N_10131,N_7518,N_6827);
and U10132 (N_10132,N_8341,N_8346);
and U10133 (N_10133,N_8526,N_7820);
nand U10134 (N_10134,N_7782,N_6158);
and U10135 (N_10135,N_6639,N_8976);
or U10136 (N_10136,N_7462,N_8149);
nor U10137 (N_10137,N_6702,N_8803);
nand U10138 (N_10138,N_6455,N_6841);
nor U10139 (N_10139,N_6243,N_8036);
nand U10140 (N_10140,N_7162,N_8024);
or U10141 (N_10141,N_8249,N_8041);
nor U10142 (N_10142,N_6383,N_8050);
nor U10143 (N_10143,N_7108,N_6837);
nor U10144 (N_10144,N_6007,N_6327);
xor U10145 (N_10145,N_6107,N_6091);
nand U10146 (N_10146,N_8141,N_8974);
and U10147 (N_10147,N_7029,N_7646);
and U10148 (N_10148,N_8408,N_8359);
or U10149 (N_10149,N_8641,N_7390);
nor U10150 (N_10150,N_7904,N_8778);
or U10151 (N_10151,N_7070,N_7119);
nand U10152 (N_10152,N_6045,N_7973);
or U10153 (N_10153,N_7169,N_6526);
or U10154 (N_10154,N_8336,N_6457);
nand U10155 (N_10155,N_6986,N_8898);
nand U10156 (N_10156,N_6691,N_6026);
nand U10157 (N_10157,N_7135,N_8651);
and U10158 (N_10158,N_7505,N_6357);
nor U10159 (N_10159,N_7128,N_8681);
nand U10160 (N_10160,N_7474,N_8629);
nor U10161 (N_10161,N_7616,N_7656);
or U10162 (N_10162,N_6294,N_8958);
nand U10163 (N_10163,N_8384,N_7260);
nor U10164 (N_10164,N_6801,N_8243);
or U10165 (N_10165,N_8479,N_8451);
nand U10166 (N_10166,N_7270,N_6187);
or U10167 (N_10167,N_7239,N_7596);
nor U10168 (N_10168,N_6706,N_6719);
nand U10169 (N_10169,N_7388,N_6360);
or U10170 (N_10170,N_6732,N_6099);
nor U10171 (N_10171,N_6966,N_7763);
nand U10172 (N_10172,N_7403,N_6648);
and U10173 (N_10173,N_7340,N_7096);
nand U10174 (N_10174,N_6169,N_7770);
nor U10175 (N_10175,N_8184,N_8178);
or U10176 (N_10176,N_7493,N_7607);
and U10177 (N_10177,N_8568,N_6571);
or U10178 (N_10178,N_6853,N_7923);
or U10179 (N_10179,N_6818,N_7434);
and U10180 (N_10180,N_7577,N_6005);
nand U10181 (N_10181,N_6112,N_8432);
and U10182 (N_10182,N_6450,N_8983);
and U10183 (N_10183,N_8509,N_7367);
and U10184 (N_10184,N_7794,N_6154);
and U10185 (N_10185,N_6011,N_6504);
nand U10186 (N_10186,N_7615,N_8908);
and U10187 (N_10187,N_7406,N_8361);
or U10188 (N_10188,N_6239,N_8323);
or U10189 (N_10189,N_7673,N_6569);
nor U10190 (N_10190,N_6353,N_8242);
nand U10191 (N_10191,N_7784,N_7780);
or U10192 (N_10192,N_6687,N_8643);
and U10193 (N_10193,N_7841,N_7213);
and U10194 (N_10194,N_7018,N_8253);
nor U10195 (N_10195,N_8500,N_6137);
and U10196 (N_10196,N_8809,N_8131);
xnor U10197 (N_10197,N_6972,N_8364);
and U10198 (N_10198,N_6490,N_7365);
nor U10199 (N_10199,N_8230,N_6048);
nand U10200 (N_10200,N_7106,N_8684);
nor U10201 (N_10201,N_6775,N_8556);
nor U10202 (N_10202,N_6034,N_6998);
nor U10203 (N_10203,N_7509,N_7373);
and U10204 (N_10204,N_6423,N_6328);
nand U10205 (N_10205,N_6075,N_6728);
and U10206 (N_10206,N_6975,N_7198);
or U10207 (N_10207,N_7565,N_6520);
nand U10208 (N_10208,N_7250,N_7928);
or U10209 (N_10209,N_6070,N_8842);
nor U10210 (N_10210,N_6984,N_6963);
nor U10211 (N_10211,N_8950,N_8838);
nand U10212 (N_10212,N_7789,N_7661);
nand U10213 (N_10213,N_7407,N_6684);
and U10214 (N_10214,N_8305,N_8320);
and U10215 (N_10215,N_7988,N_6448);
and U10216 (N_10216,N_7005,N_8700);
nor U10217 (N_10217,N_8373,N_6385);
and U10218 (N_10218,N_6770,N_7909);
or U10219 (N_10219,N_6920,N_7276);
and U10220 (N_10220,N_6610,N_6313);
and U10221 (N_10221,N_7660,N_7315);
nand U10222 (N_10222,N_8174,N_8941);
nor U10223 (N_10223,N_8204,N_6362);
and U10224 (N_10224,N_6058,N_7640);
nor U10225 (N_10225,N_6376,N_7704);
or U10226 (N_10226,N_8347,N_6393);
nor U10227 (N_10227,N_6740,N_6247);
or U10228 (N_10228,N_8907,N_6390);
nand U10229 (N_10229,N_6548,N_6463);
and U10230 (N_10230,N_6933,N_6854);
and U10231 (N_10231,N_8810,N_8510);
nor U10232 (N_10232,N_8797,N_7972);
or U10233 (N_10233,N_7151,N_6560);
or U10234 (N_10234,N_8889,N_6398);
nor U10235 (N_10235,N_7455,N_8971);
and U10236 (N_10236,N_6062,N_7446);
and U10237 (N_10237,N_6846,N_6101);
nor U10238 (N_10238,N_6291,N_8005);
and U10239 (N_10239,N_6847,N_7512);
or U10240 (N_10240,N_7579,N_8738);
nand U10241 (N_10241,N_7955,N_6671);
xnor U10242 (N_10242,N_8163,N_8368);
or U10243 (N_10243,N_8870,N_7371);
and U10244 (N_10244,N_6621,N_7702);
nand U10245 (N_10245,N_7489,N_7307);
or U10246 (N_10246,N_7943,N_6146);
nand U10247 (N_10247,N_8306,N_7824);
xor U10248 (N_10248,N_6889,N_6903);
nor U10249 (N_10249,N_6192,N_6248);
or U10250 (N_10250,N_7588,N_6976);
and U10251 (N_10251,N_7582,N_8213);
nor U10252 (N_10252,N_7320,N_6951);
nor U10253 (N_10253,N_7657,N_8281);
nand U10254 (N_10254,N_6830,N_6807);
nor U10255 (N_10255,N_8138,N_6109);
nand U10256 (N_10256,N_7870,N_6025);
nand U10257 (N_10257,N_7019,N_6003);
nand U10258 (N_10258,N_6910,N_7694);
or U10259 (N_10259,N_6069,N_8688);
nor U10260 (N_10260,N_7707,N_6969);
nand U10261 (N_10261,N_7279,N_6925);
and U10262 (N_10262,N_6217,N_8356);
nand U10263 (N_10263,N_6590,N_8724);
and U10264 (N_10264,N_8332,N_6954);
nand U10265 (N_10265,N_6207,N_6544);
nand U10266 (N_10266,N_7562,N_8419);
and U10267 (N_10267,N_7648,N_7756);
and U10268 (N_10268,N_6418,N_7424);
and U10269 (N_10269,N_8567,N_7513);
nand U10270 (N_10270,N_7911,N_7178);
or U10271 (N_10271,N_8750,N_6073);
or U10272 (N_10272,N_7832,N_8854);
or U10273 (N_10273,N_7677,N_6411);
and U10274 (N_10274,N_6032,N_7980);
nand U10275 (N_10275,N_7806,N_6372);
or U10276 (N_10276,N_6786,N_6152);
or U10277 (N_10277,N_8283,N_8358);
nor U10278 (N_10278,N_8936,N_6370);
and U10279 (N_10279,N_7225,N_6944);
nand U10280 (N_10280,N_7378,N_6189);
or U10281 (N_10281,N_7215,N_6879);
or U10282 (N_10282,N_6619,N_7966);
nor U10283 (N_10283,N_7617,N_8528);
nor U10284 (N_10284,N_8614,N_8392);
or U10285 (N_10285,N_7862,N_8223);
nor U10286 (N_10286,N_8485,N_6712);
or U10287 (N_10287,N_7485,N_6502);
nand U10288 (N_10288,N_7028,N_8595);
or U10289 (N_10289,N_6783,N_7566);
nor U10290 (N_10290,N_8463,N_8538);
and U10291 (N_10291,N_6481,N_8591);
and U10292 (N_10292,N_8808,N_7956);
nor U10293 (N_10293,N_7891,N_7334);
or U10294 (N_10294,N_8504,N_8153);
nand U10295 (N_10295,N_7154,N_8351);
and U10296 (N_10296,N_6273,N_8313);
or U10297 (N_10297,N_7599,N_6575);
and U10298 (N_10298,N_6568,N_6198);
nand U10299 (N_10299,N_7192,N_8999);
and U10300 (N_10300,N_8134,N_6822);
nor U10301 (N_10301,N_7652,N_6887);
or U10302 (N_10302,N_8234,N_8727);
nand U10303 (N_10303,N_7142,N_7109);
and U10304 (N_10304,N_6380,N_8418);
or U10305 (N_10305,N_7632,N_8052);
and U10306 (N_10306,N_8699,N_6952);
or U10307 (N_10307,N_7696,N_7040);
nand U10308 (N_10308,N_6176,N_6755);
nor U10309 (N_10309,N_7766,N_7071);
or U10310 (N_10310,N_8805,N_8703);
nor U10311 (N_10311,N_7421,N_7930);
and U10312 (N_10312,N_6611,N_6894);
nor U10313 (N_10313,N_8817,N_6734);
nand U10314 (N_10314,N_8133,N_6339);
nor U10315 (N_10315,N_6330,N_6686);
nor U10316 (N_10316,N_6279,N_7013);
nor U10317 (N_10317,N_8757,N_6156);
and U10318 (N_10318,N_8353,N_8775);
xnor U10319 (N_10319,N_7100,N_8906);
and U10320 (N_10320,N_7091,N_6183);
or U10321 (N_10321,N_6793,N_7547);
or U10322 (N_10322,N_8334,N_8067);
or U10323 (N_10323,N_6531,N_8830);
nand U10324 (N_10324,N_7614,N_8438);
or U10325 (N_10325,N_6505,N_6803);
nand U10326 (N_10326,N_8034,N_6787);
and U10327 (N_10327,N_7330,N_6961);
nor U10328 (N_10328,N_7158,N_7618);
nor U10329 (N_10329,N_8088,N_6817);
and U10330 (N_10330,N_6762,N_7042);
nor U10331 (N_10331,N_8172,N_7967);
nand U10332 (N_10332,N_7884,N_7405);
and U10333 (N_10333,N_7094,N_6855);
nand U10334 (N_10334,N_7176,N_8370);
xnor U10335 (N_10335,N_7442,N_7817);
and U10336 (N_10336,N_8858,N_8407);
or U10337 (N_10337,N_6643,N_7725);
or U10338 (N_10338,N_8598,N_7265);
nand U10339 (N_10339,N_7589,N_7342);
nor U10340 (N_10340,N_8758,N_8237);
nor U10341 (N_10341,N_8883,N_7024);
or U10342 (N_10342,N_6628,N_6883);
or U10343 (N_10343,N_8265,N_6580);
nand U10344 (N_10344,N_6468,N_7970);
and U10345 (N_10345,N_7295,N_7282);
or U10346 (N_10346,N_6539,N_6249);
xnor U10347 (N_10347,N_8093,N_6072);
nand U10348 (N_10348,N_8268,N_8683);
or U10349 (N_10349,N_7510,N_8710);
nand U10350 (N_10350,N_7314,N_8638);
nor U10351 (N_10351,N_8191,N_6915);
and U10352 (N_10352,N_6790,N_8311);
or U10353 (N_10353,N_6236,N_7359);
or U10354 (N_10354,N_7849,N_7020);
nor U10355 (N_10355,N_8774,N_7836);
and U10356 (N_10356,N_7006,N_6186);
nor U10357 (N_10357,N_8522,N_7248);
nand U10358 (N_10358,N_7787,N_7951);
nand U10359 (N_10359,N_6132,N_7436);
and U10360 (N_10360,N_7274,N_7938);
and U10361 (N_10361,N_7148,N_8844);
nand U10362 (N_10362,N_7203,N_8723);
nor U10363 (N_10363,N_8221,N_7098);
nand U10364 (N_10364,N_6244,N_8431);
nor U10365 (N_10365,N_8835,N_8879);
or U10366 (N_10366,N_6094,N_8004);
or U10367 (N_10367,N_7107,N_6871);
nand U10368 (N_10368,N_7598,N_7397);
nor U10369 (N_10369,N_7679,N_7498);
nand U10370 (N_10370,N_7638,N_7719);
nand U10371 (N_10371,N_8981,N_8821);
nor U10372 (N_10372,N_6098,N_6923);
nand U10373 (N_10373,N_6895,N_8205);
nand U10374 (N_10374,N_6709,N_7818);
and U10375 (N_10375,N_6743,N_7187);
and U10376 (N_10376,N_6949,N_8081);
and U10377 (N_10377,N_6878,N_8517);
nor U10378 (N_10378,N_7669,N_7603);
nand U10379 (N_10379,N_6197,N_6275);
or U10380 (N_10380,N_6761,N_6453);
and U10381 (N_10381,N_8761,N_8662);
nand U10382 (N_10382,N_7105,N_7647);
nor U10383 (N_10383,N_6810,N_8578);
or U10384 (N_10384,N_7503,N_7177);
nor U10385 (N_10385,N_6133,N_8421);
and U10386 (N_10386,N_7095,N_6190);
or U10387 (N_10387,N_7575,N_8319);
or U10388 (N_10388,N_7398,N_8477);
nor U10389 (N_10389,N_7186,N_7650);
nand U10390 (N_10390,N_7076,N_7511);
and U10391 (N_10391,N_8558,N_6474);
nor U10392 (N_10392,N_8536,N_7170);
or U10393 (N_10393,N_8189,N_7425);
nor U10394 (N_10394,N_7370,N_6268);
or U10395 (N_10395,N_6220,N_6274);
nand U10396 (N_10396,N_8457,N_7387);
nor U10397 (N_10397,N_7391,N_8634);
nor U10398 (N_10398,N_8498,N_8995);
or U10399 (N_10399,N_6280,N_8876);
nand U10400 (N_10400,N_7477,N_7145);
or U10401 (N_10401,N_8413,N_6598);
nor U10402 (N_10402,N_6907,N_8546);
or U10403 (N_10403,N_6913,N_6641);
and U10404 (N_10404,N_6723,N_8276);
nand U10405 (N_10405,N_8759,N_8095);
nand U10406 (N_10406,N_6277,N_6057);
nor U10407 (N_10407,N_7126,N_6266);
nand U10408 (N_10408,N_8676,N_6439);
or U10409 (N_10409,N_7345,N_7384);
nand U10410 (N_10410,N_8166,N_6912);
nand U10411 (N_10411,N_7741,N_7252);
nand U10412 (N_10412,N_8773,N_6697);
or U10413 (N_10413,N_8371,N_6747);
nor U10414 (N_10414,N_7205,N_6891);
nand U10415 (N_10415,N_6023,N_6486);
nor U10416 (N_10416,N_7844,N_7609);
nand U10417 (N_10417,N_8777,N_8474);
nor U10418 (N_10418,N_8947,N_6231);
nand U10419 (N_10419,N_7597,N_8726);
or U10420 (N_10420,N_7674,N_6386);
nand U10421 (N_10421,N_6103,N_6227);
nand U10422 (N_10422,N_8579,N_8487);
or U10423 (N_10423,N_8825,N_8279);
nor U10424 (N_10424,N_8554,N_8659);
and U10425 (N_10425,N_7116,N_6752);
and U10426 (N_10426,N_8130,N_6478);
nand U10427 (N_10427,N_8966,N_8964);
and U10428 (N_10428,N_8310,N_8157);
nor U10429 (N_10429,N_7822,N_6306);
or U10430 (N_10430,N_7319,N_7812);
nand U10431 (N_10431,N_8111,N_6655);
and U10432 (N_10432,N_8919,N_7665);
and U10433 (N_10433,N_6536,N_6323);
or U10434 (N_10434,N_6727,N_7479);
or U10435 (N_10435,N_6430,N_6157);
nand U10436 (N_10436,N_6823,N_7581);
nand U10437 (N_10437,N_6037,N_8122);
and U10438 (N_10438,N_8167,N_8051);
nand U10439 (N_10439,N_8140,N_7327);
and U10440 (N_10440,N_7508,N_7842);
nor U10441 (N_10441,N_7423,N_7247);
nand U10442 (N_10442,N_8126,N_7690);
nand U10443 (N_10443,N_7476,N_8220);
nand U10444 (N_10444,N_6162,N_8819);
nand U10445 (N_10445,N_8886,N_7857);
nand U10446 (N_10446,N_7611,N_7218);
nor U10447 (N_10447,N_8354,N_8864);
nand U10448 (N_10448,N_7742,N_8686);
and U10449 (N_10449,N_8943,N_7336);
and U10450 (N_10450,N_6800,N_6885);
and U10451 (N_10451,N_6467,N_6549);
and U10452 (N_10452,N_7537,N_7361);
nand U10453 (N_10453,N_6314,N_6212);
nand U10454 (N_10454,N_7709,N_7399);
nor U10455 (N_10455,N_8555,N_6663);
nor U10456 (N_10456,N_8987,N_8103);
or U10457 (N_10457,N_8459,N_7875);
nand U10458 (N_10458,N_6703,N_6964);
nor U10459 (N_10459,N_7667,N_6449);
nand U10460 (N_10460,N_6860,N_7409);
and U10461 (N_10461,N_6929,N_8239);
or U10462 (N_10462,N_6707,N_8540);
and U10463 (N_10463,N_7324,N_7645);
or U10464 (N_10464,N_8070,N_8462);
nor U10465 (N_10465,N_6875,N_7689);
nand U10466 (N_10466,N_6181,N_6967);
or U10467 (N_10467,N_8113,N_7392);
and U10468 (N_10468,N_6300,N_6379);
and U10469 (N_10469,N_8304,N_8732);
or U10470 (N_10470,N_7775,N_8832);
or U10471 (N_10471,N_6060,N_8529);
and U10472 (N_10472,N_6392,N_6333);
nand U10473 (N_10473,N_6908,N_8698);
nand U10474 (N_10474,N_7860,N_8519);
and U10475 (N_10475,N_7068,N_6361);
nor U10476 (N_10476,N_7083,N_6731);
nor U10477 (N_10477,N_8693,N_6343);
and U10478 (N_10478,N_7375,N_8539);
or U10479 (N_10479,N_8010,N_7271);
and U10480 (N_10480,N_7850,N_7727);
nand U10481 (N_10481,N_6271,N_7981);
nor U10482 (N_10482,N_7521,N_7662);
and U10483 (N_10483,N_8302,N_6226);
and U10484 (N_10484,N_6748,N_7111);
and U10485 (N_10485,N_6100,N_6024);
nor U10486 (N_10486,N_6909,N_6347);
or U10487 (N_10487,N_6331,N_6573);
and U10488 (N_10488,N_8386,N_6139);
nor U10489 (N_10489,N_7659,N_6191);
nor U10490 (N_10490,N_6378,N_8039);
nor U10491 (N_10491,N_7948,N_7584);
nor U10492 (N_10492,N_6260,N_8933);
nor U10493 (N_10493,N_6532,N_6694);
nand U10494 (N_10494,N_6442,N_8247);
nand U10495 (N_10495,N_7957,N_6451);
or U10496 (N_10496,N_8007,N_7843);
or U10497 (N_10497,N_6792,N_6336);
or U10498 (N_10498,N_8799,N_6320);
nand U10499 (N_10499,N_8318,N_7807);
and U10500 (N_10500,N_7008,N_6912);
nand U10501 (N_10501,N_6896,N_7808);
and U10502 (N_10502,N_8887,N_7302);
or U10503 (N_10503,N_6551,N_6287);
or U10504 (N_10504,N_8574,N_7572);
or U10505 (N_10505,N_8219,N_8720);
nor U10506 (N_10506,N_6821,N_6817);
or U10507 (N_10507,N_7949,N_6474);
and U10508 (N_10508,N_6559,N_8893);
or U10509 (N_10509,N_7477,N_7623);
nor U10510 (N_10510,N_8897,N_8737);
nor U10511 (N_10511,N_8862,N_8131);
or U10512 (N_10512,N_6941,N_7205);
nor U10513 (N_10513,N_8025,N_6269);
and U10514 (N_10514,N_6417,N_8340);
nand U10515 (N_10515,N_6936,N_7120);
and U10516 (N_10516,N_6191,N_6545);
nand U10517 (N_10517,N_8550,N_6138);
or U10518 (N_10518,N_8930,N_6590);
or U10519 (N_10519,N_7416,N_8236);
and U10520 (N_10520,N_7379,N_8761);
nor U10521 (N_10521,N_8258,N_8262);
and U10522 (N_10522,N_7944,N_8312);
nand U10523 (N_10523,N_8121,N_7706);
nand U10524 (N_10524,N_8709,N_8529);
or U10525 (N_10525,N_7147,N_8695);
or U10526 (N_10526,N_8658,N_7559);
nor U10527 (N_10527,N_6689,N_8560);
and U10528 (N_10528,N_6710,N_8298);
nand U10529 (N_10529,N_6244,N_7898);
nor U10530 (N_10530,N_6646,N_8255);
and U10531 (N_10531,N_8289,N_6593);
nand U10532 (N_10532,N_6331,N_7245);
or U10533 (N_10533,N_6578,N_8972);
or U10534 (N_10534,N_8576,N_7551);
and U10535 (N_10535,N_7209,N_8161);
nor U10536 (N_10536,N_6644,N_7100);
or U10537 (N_10537,N_6309,N_7813);
and U10538 (N_10538,N_6876,N_8208);
nand U10539 (N_10539,N_6458,N_6950);
or U10540 (N_10540,N_7651,N_8347);
and U10541 (N_10541,N_7832,N_6502);
nor U10542 (N_10542,N_6298,N_6951);
nor U10543 (N_10543,N_8755,N_8664);
nand U10544 (N_10544,N_8199,N_8555);
nor U10545 (N_10545,N_8333,N_8778);
and U10546 (N_10546,N_7257,N_7462);
nand U10547 (N_10547,N_8189,N_6575);
nand U10548 (N_10548,N_6205,N_6459);
nand U10549 (N_10549,N_7567,N_7575);
and U10550 (N_10550,N_8129,N_8866);
or U10551 (N_10551,N_7844,N_6382);
nand U10552 (N_10552,N_8273,N_6591);
or U10553 (N_10553,N_6947,N_7664);
nand U10554 (N_10554,N_8565,N_7874);
or U10555 (N_10555,N_6441,N_6790);
nand U10556 (N_10556,N_6626,N_7380);
nor U10557 (N_10557,N_6096,N_7242);
nor U10558 (N_10558,N_6659,N_6785);
nand U10559 (N_10559,N_6507,N_6734);
or U10560 (N_10560,N_6160,N_8720);
or U10561 (N_10561,N_8672,N_8311);
or U10562 (N_10562,N_6685,N_6059);
and U10563 (N_10563,N_8096,N_6948);
or U10564 (N_10564,N_6865,N_7261);
nor U10565 (N_10565,N_8200,N_6995);
nor U10566 (N_10566,N_7430,N_7583);
and U10567 (N_10567,N_6758,N_8097);
and U10568 (N_10568,N_6624,N_7584);
nand U10569 (N_10569,N_6909,N_6373);
and U10570 (N_10570,N_8865,N_8125);
and U10571 (N_10571,N_8713,N_7760);
nor U10572 (N_10572,N_6120,N_8524);
nand U10573 (N_10573,N_7975,N_7181);
nand U10574 (N_10574,N_7969,N_6872);
or U10575 (N_10575,N_8477,N_8267);
nor U10576 (N_10576,N_7228,N_6207);
or U10577 (N_10577,N_7973,N_8946);
nand U10578 (N_10578,N_6725,N_8970);
nand U10579 (N_10579,N_7347,N_7290);
nand U10580 (N_10580,N_7587,N_7103);
and U10581 (N_10581,N_7131,N_6412);
nand U10582 (N_10582,N_7051,N_7897);
or U10583 (N_10583,N_6866,N_8135);
or U10584 (N_10584,N_7515,N_6800);
nor U10585 (N_10585,N_8252,N_7384);
nor U10586 (N_10586,N_6647,N_7722);
or U10587 (N_10587,N_6833,N_8354);
and U10588 (N_10588,N_6220,N_6195);
nor U10589 (N_10589,N_8197,N_7556);
or U10590 (N_10590,N_8054,N_7727);
and U10591 (N_10591,N_6950,N_8312);
nand U10592 (N_10592,N_7711,N_7440);
xor U10593 (N_10593,N_6041,N_8131);
nand U10594 (N_10594,N_7183,N_8692);
and U10595 (N_10595,N_7321,N_8299);
nor U10596 (N_10596,N_8058,N_6550);
and U10597 (N_10597,N_6722,N_6300);
nand U10598 (N_10598,N_7058,N_7794);
and U10599 (N_10599,N_7271,N_8301);
nand U10600 (N_10600,N_8047,N_7808);
nand U10601 (N_10601,N_7409,N_6943);
or U10602 (N_10602,N_8336,N_8164);
and U10603 (N_10603,N_8893,N_6606);
nand U10604 (N_10604,N_7149,N_8696);
or U10605 (N_10605,N_7764,N_6301);
nand U10606 (N_10606,N_8206,N_6164);
nor U10607 (N_10607,N_6746,N_7400);
and U10608 (N_10608,N_6816,N_7389);
nor U10609 (N_10609,N_6266,N_6051);
nand U10610 (N_10610,N_8592,N_8663);
and U10611 (N_10611,N_6807,N_6327);
nand U10612 (N_10612,N_8672,N_6187);
or U10613 (N_10613,N_7661,N_8102);
or U10614 (N_10614,N_6612,N_8463);
nand U10615 (N_10615,N_7982,N_7670);
and U10616 (N_10616,N_6551,N_8149);
and U10617 (N_10617,N_6154,N_6226);
nor U10618 (N_10618,N_8916,N_6697);
or U10619 (N_10619,N_7471,N_7766);
nand U10620 (N_10620,N_8966,N_8561);
nor U10621 (N_10621,N_6868,N_7245);
nor U10622 (N_10622,N_7533,N_8540);
and U10623 (N_10623,N_8558,N_7311);
nor U10624 (N_10624,N_7294,N_6680);
or U10625 (N_10625,N_6438,N_7050);
and U10626 (N_10626,N_8095,N_6442);
nand U10627 (N_10627,N_7607,N_7946);
or U10628 (N_10628,N_8101,N_8814);
nand U10629 (N_10629,N_8647,N_6112);
and U10630 (N_10630,N_6778,N_6617);
nand U10631 (N_10631,N_6808,N_7142);
and U10632 (N_10632,N_6930,N_6957);
or U10633 (N_10633,N_7778,N_8592);
and U10634 (N_10634,N_7757,N_6657);
or U10635 (N_10635,N_7869,N_7353);
nand U10636 (N_10636,N_6355,N_6559);
nor U10637 (N_10637,N_6466,N_7276);
or U10638 (N_10638,N_7082,N_6166);
and U10639 (N_10639,N_8676,N_8938);
nand U10640 (N_10640,N_7363,N_7036);
nand U10641 (N_10641,N_6538,N_8596);
or U10642 (N_10642,N_8346,N_7413);
nand U10643 (N_10643,N_8414,N_7424);
and U10644 (N_10644,N_7867,N_8064);
nand U10645 (N_10645,N_7019,N_7835);
nor U10646 (N_10646,N_8110,N_6845);
and U10647 (N_10647,N_6337,N_7664);
and U10648 (N_10648,N_7590,N_6472);
or U10649 (N_10649,N_8875,N_6805);
nor U10650 (N_10650,N_6486,N_6348);
and U10651 (N_10651,N_6865,N_6562);
xor U10652 (N_10652,N_8053,N_7514);
nor U10653 (N_10653,N_8894,N_7339);
and U10654 (N_10654,N_8944,N_8976);
nor U10655 (N_10655,N_8689,N_7877);
nand U10656 (N_10656,N_8760,N_7862);
or U10657 (N_10657,N_7366,N_8668);
nor U10658 (N_10658,N_6126,N_6554);
nand U10659 (N_10659,N_7731,N_6353);
or U10660 (N_10660,N_8059,N_6330);
nand U10661 (N_10661,N_6525,N_8913);
nand U10662 (N_10662,N_6885,N_7549);
nand U10663 (N_10663,N_6258,N_7473);
and U10664 (N_10664,N_6166,N_6064);
and U10665 (N_10665,N_7261,N_8091);
or U10666 (N_10666,N_8654,N_8411);
or U10667 (N_10667,N_8708,N_6643);
and U10668 (N_10668,N_6400,N_8501);
and U10669 (N_10669,N_7718,N_6975);
and U10670 (N_10670,N_8158,N_7659);
nor U10671 (N_10671,N_8543,N_7140);
nand U10672 (N_10672,N_8249,N_7905);
nor U10673 (N_10673,N_7963,N_8978);
nor U10674 (N_10674,N_6246,N_8223);
or U10675 (N_10675,N_7067,N_7380);
or U10676 (N_10676,N_6422,N_6132);
and U10677 (N_10677,N_7872,N_6781);
and U10678 (N_10678,N_6077,N_8727);
or U10679 (N_10679,N_7852,N_8335);
and U10680 (N_10680,N_7788,N_8620);
nand U10681 (N_10681,N_7900,N_7046);
nand U10682 (N_10682,N_8535,N_7679);
nand U10683 (N_10683,N_8817,N_7638);
or U10684 (N_10684,N_8599,N_8374);
or U10685 (N_10685,N_8535,N_6777);
or U10686 (N_10686,N_6752,N_8165);
nand U10687 (N_10687,N_8549,N_7211);
nand U10688 (N_10688,N_8019,N_6511);
xnor U10689 (N_10689,N_8575,N_7400);
nor U10690 (N_10690,N_6311,N_6544);
nand U10691 (N_10691,N_7245,N_7857);
nor U10692 (N_10692,N_6765,N_7653);
nor U10693 (N_10693,N_7087,N_7138);
nand U10694 (N_10694,N_8672,N_7199);
nand U10695 (N_10695,N_8007,N_8235);
nand U10696 (N_10696,N_6677,N_7424);
nor U10697 (N_10697,N_6715,N_7800);
and U10698 (N_10698,N_6517,N_8574);
and U10699 (N_10699,N_7410,N_6398);
xnor U10700 (N_10700,N_6453,N_6465);
xnor U10701 (N_10701,N_8089,N_8290);
or U10702 (N_10702,N_8936,N_8698);
and U10703 (N_10703,N_7943,N_8080);
nand U10704 (N_10704,N_6883,N_8050);
nand U10705 (N_10705,N_7624,N_6764);
or U10706 (N_10706,N_8423,N_6836);
nand U10707 (N_10707,N_8488,N_6926);
nor U10708 (N_10708,N_7673,N_6640);
nand U10709 (N_10709,N_8224,N_7343);
and U10710 (N_10710,N_7824,N_8704);
nor U10711 (N_10711,N_7637,N_8118);
nand U10712 (N_10712,N_8236,N_8312);
nand U10713 (N_10713,N_7605,N_8116);
or U10714 (N_10714,N_6216,N_7126);
nand U10715 (N_10715,N_8200,N_6844);
nand U10716 (N_10716,N_7964,N_6591);
nand U10717 (N_10717,N_6258,N_6987);
nor U10718 (N_10718,N_8732,N_6814);
or U10719 (N_10719,N_7773,N_7219);
nand U10720 (N_10720,N_6505,N_6687);
or U10721 (N_10721,N_8380,N_8694);
nor U10722 (N_10722,N_8149,N_8583);
and U10723 (N_10723,N_7664,N_6810);
and U10724 (N_10724,N_6370,N_6057);
nand U10725 (N_10725,N_7901,N_6916);
nor U10726 (N_10726,N_7008,N_6303);
nand U10727 (N_10727,N_8323,N_8536);
xor U10728 (N_10728,N_7409,N_8815);
and U10729 (N_10729,N_8216,N_7358);
nor U10730 (N_10730,N_8241,N_8326);
nand U10731 (N_10731,N_8386,N_7445);
nor U10732 (N_10732,N_6087,N_8625);
nor U10733 (N_10733,N_6150,N_8142);
or U10734 (N_10734,N_7257,N_7074);
or U10735 (N_10735,N_7054,N_8485);
or U10736 (N_10736,N_8854,N_7726);
and U10737 (N_10737,N_6398,N_8618);
or U10738 (N_10738,N_8321,N_7692);
and U10739 (N_10739,N_7871,N_7851);
or U10740 (N_10740,N_7221,N_8466);
and U10741 (N_10741,N_7212,N_8005);
or U10742 (N_10742,N_7153,N_8021);
and U10743 (N_10743,N_7925,N_7828);
nand U10744 (N_10744,N_6153,N_7961);
and U10745 (N_10745,N_7671,N_6198);
and U10746 (N_10746,N_7663,N_8603);
or U10747 (N_10747,N_7286,N_8038);
xor U10748 (N_10748,N_8551,N_7618);
and U10749 (N_10749,N_6120,N_8357);
or U10750 (N_10750,N_7796,N_8114);
nor U10751 (N_10751,N_7222,N_7711);
nor U10752 (N_10752,N_6423,N_6794);
or U10753 (N_10753,N_8979,N_8100);
nor U10754 (N_10754,N_8869,N_8633);
nand U10755 (N_10755,N_7737,N_8469);
nand U10756 (N_10756,N_7751,N_8747);
and U10757 (N_10757,N_6956,N_7218);
nand U10758 (N_10758,N_8288,N_6259);
nand U10759 (N_10759,N_8629,N_7451);
or U10760 (N_10760,N_6028,N_8891);
nor U10761 (N_10761,N_8448,N_6899);
nor U10762 (N_10762,N_7833,N_8748);
nand U10763 (N_10763,N_6508,N_7601);
or U10764 (N_10764,N_8591,N_7028);
and U10765 (N_10765,N_6057,N_6010);
and U10766 (N_10766,N_6868,N_8922);
nor U10767 (N_10767,N_6717,N_7773);
and U10768 (N_10768,N_8343,N_7509);
or U10769 (N_10769,N_6059,N_8572);
nor U10770 (N_10770,N_8867,N_8459);
nor U10771 (N_10771,N_8213,N_8532);
and U10772 (N_10772,N_7262,N_8776);
nand U10773 (N_10773,N_6857,N_7440);
or U10774 (N_10774,N_8555,N_6973);
nand U10775 (N_10775,N_8946,N_7494);
nor U10776 (N_10776,N_7215,N_8457);
nand U10777 (N_10777,N_6904,N_8462);
nand U10778 (N_10778,N_8241,N_6683);
or U10779 (N_10779,N_8673,N_8785);
nand U10780 (N_10780,N_7528,N_6372);
and U10781 (N_10781,N_8313,N_6709);
and U10782 (N_10782,N_6978,N_6499);
or U10783 (N_10783,N_6708,N_8518);
nor U10784 (N_10784,N_7865,N_7450);
nor U10785 (N_10785,N_6636,N_8006);
and U10786 (N_10786,N_7104,N_7198);
nor U10787 (N_10787,N_7015,N_6150);
nand U10788 (N_10788,N_6791,N_7564);
nor U10789 (N_10789,N_6410,N_6683);
nand U10790 (N_10790,N_6700,N_7794);
nor U10791 (N_10791,N_6062,N_7620);
or U10792 (N_10792,N_7746,N_7221);
nand U10793 (N_10793,N_8905,N_8565);
nand U10794 (N_10794,N_7208,N_8572);
or U10795 (N_10795,N_8167,N_6107);
nor U10796 (N_10796,N_6794,N_8964);
nor U10797 (N_10797,N_6940,N_7575);
nand U10798 (N_10798,N_6288,N_6981);
nor U10799 (N_10799,N_8295,N_8140);
or U10800 (N_10800,N_6748,N_8038);
nor U10801 (N_10801,N_6882,N_7406);
nand U10802 (N_10802,N_8648,N_7610);
and U10803 (N_10803,N_6507,N_7297);
or U10804 (N_10804,N_6986,N_8607);
nand U10805 (N_10805,N_7007,N_8384);
or U10806 (N_10806,N_8344,N_7645);
nand U10807 (N_10807,N_6304,N_6458);
and U10808 (N_10808,N_6835,N_7126);
and U10809 (N_10809,N_8845,N_8459);
or U10810 (N_10810,N_7412,N_8242);
nand U10811 (N_10811,N_8813,N_7009);
and U10812 (N_10812,N_6847,N_7747);
or U10813 (N_10813,N_7403,N_6380);
nor U10814 (N_10814,N_8570,N_7397);
and U10815 (N_10815,N_7093,N_6040);
nand U10816 (N_10816,N_8095,N_8486);
nand U10817 (N_10817,N_7120,N_8158);
or U10818 (N_10818,N_8082,N_8292);
nand U10819 (N_10819,N_8385,N_8008);
and U10820 (N_10820,N_7228,N_6932);
nand U10821 (N_10821,N_7837,N_8499);
or U10822 (N_10822,N_8042,N_6749);
nor U10823 (N_10823,N_8667,N_6893);
nand U10824 (N_10824,N_6648,N_6424);
or U10825 (N_10825,N_6286,N_8313);
nor U10826 (N_10826,N_6220,N_7690);
nor U10827 (N_10827,N_6123,N_8357);
or U10828 (N_10828,N_7530,N_7444);
and U10829 (N_10829,N_6480,N_7861);
nand U10830 (N_10830,N_6763,N_6022);
nor U10831 (N_10831,N_6656,N_8866);
nand U10832 (N_10832,N_7668,N_6600);
nor U10833 (N_10833,N_8734,N_7411);
xor U10834 (N_10834,N_6024,N_8298);
nor U10835 (N_10835,N_6305,N_8386);
or U10836 (N_10836,N_7653,N_6539);
or U10837 (N_10837,N_6356,N_6011);
or U10838 (N_10838,N_8492,N_8140);
or U10839 (N_10839,N_7893,N_8315);
nand U10840 (N_10840,N_6197,N_7536);
nand U10841 (N_10841,N_6414,N_8644);
xnor U10842 (N_10842,N_6527,N_7872);
nand U10843 (N_10843,N_7940,N_7794);
or U10844 (N_10844,N_6134,N_6903);
or U10845 (N_10845,N_6959,N_8007);
or U10846 (N_10846,N_7334,N_6021);
nor U10847 (N_10847,N_8911,N_7353);
and U10848 (N_10848,N_6465,N_8373);
nor U10849 (N_10849,N_8116,N_6472);
nand U10850 (N_10850,N_7592,N_8507);
nand U10851 (N_10851,N_8750,N_6768);
nand U10852 (N_10852,N_7801,N_7811);
or U10853 (N_10853,N_7567,N_6513);
or U10854 (N_10854,N_6862,N_8392);
nand U10855 (N_10855,N_8834,N_8360);
or U10856 (N_10856,N_6526,N_8648);
or U10857 (N_10857,N_8283,N_7553);
nor U10858 (N_10858,N_8139,N_7282);
nor U10859 (N_10859,N_7683,N_8605);
nand U10860 (N_10860,N_7303,N_8616);
nand U10861 (N_10861,N_7244,N_7752);
nor U10862 (N_10862,N_7377,N_7818);
nand U10863 (N_10863,N_8426,N_6759);
and U10864 (N_10864,N_8179,N_6599);
or U10865 (N_10865,N_8874,N_6748);
and U10866 (N_10866,N_7210,N_7924);
nor U10867 (N_10867,N_7721,N_7727);
nor U10868 (N_10868,N_8490,N_8508);
nor U10869 (N_10869,N_8705,N_6851);
nand U10870 (N_10870,N_6496,N_8382);
and U10871 (N_10871,N_8940,N_7515);
or U10872 (N_10872,N_8428,N_6491);
nand U10873 (N_10873,N_8780,N_7243);
or U10874 (N_10874,N_6744,N_6372);
and U10875 (N_10875,N_8882,N_7217);
or U10876 (N_10876,N_7350,N_7049);
nand U10877 (N_10877,N_7782,N_7961);
and U10878 (N_10878,N_7975,N_8047);
or U10879 (N_10879,N_8194,N_8037);
or U10880 (N_10880,N_7433,N_7149);
and U10881 (N_10881,N_7618,N_6269);
nand U10882 (N_10882,N_8047,N_7537);
or U10883 (N_10883,N_8400,N_6230);
nand U10884 (N_10884,N_6257,N_7300);
nand U10885 (N_10885,N_6601,N_7245);
nand U10886 (N_10886,N_6456,N_6701);
and U10887 (N_10887,N_7658,N_7653);
and U10888 (N_10888,N_7955,N_7709);
nor U10889 (N_10889,N_6559,N_7029);
nand U10890 (N_10890,N_8350,N_7945);
or U10891 (N_10891,N_7614,N_6456);
or U10892 (N_10892,N_6514,N_6921);
nand U10893 (N_10893,N_8505,N_6982);
nand U10894 (N_10894,N_6036,N_6797);
nand U10895 (N_10895,N_7647,N_8832);
or U10896 (N_10896,N_7689,N_7524);
nor U10897 (N_10897,N_8442,N_7536);
nand U10898 (N_10898,N_8209,N_7532);
or U10899 (N_10899,N_8490,N_7669);
and U10900 (N_10900,N_7290,N_6656);
nand U10901 (N_10901,N_7949,N_7920);
or U10902 (N_10902,N_7723,N_6285);
or U10903 (N_10903,N_6845,N_8613);
nor U10904 (N_10904,N_6277,N_7441);
and U10905 (N_10905,N_6173,N_7240);
or U10906 (N_10906,N_6557,N_8420);
nor U10907 (N_10907,N_8962,N_8940);
and U10908 (N_10908,N_6886,N_7683);
nor U10909 (N_10909,N_6176,N_6275);
or U10910 (N_10910,N_7379,N_8158);
nand U10911 (N_10911,N_6914,N_6040);
and U10912 (N_10912,N_7552,N_6443);
and U10913 (N_10913,N_7012,N_6861);
nor U10914 (N_10914,N_7640,N_6409);
or U10915 (N_10915,N_7782,N_6391);
nand U10916 (N_10916,N_6777,N_8420);
and U10917 (N_10917,N_7705,N_7638);
nand U10918 (N_10918,N_7054,N_8656);
nor U10919 (N_10919,N_8332,N_7717);
or U10920 (N_10920,N_8294,N_7572);
nor U10921 (N_10921,N_6484,N_8935);
and U10922 (N_10922,N_8458,N_6890);
and U10923 (N_10923,N_7492,N_8450);
nand U10924 (N_10924,N_7960,N_8061);
and U10925 (N_10925,N_6329,N_8779);
nand U10926 (N_10926,N_6666,N_7528);
or U10927 (N_10927,N_8886,N_7780);
or U10928 (N_10928,N_6604,N_6581);
and U10929 (N_10929,N_8953,N_8006);
nor U10930 (N_10930,N_7191,N_7874);
or U10931 (N_10931,N_8516,N_6880);
and U10932 (N_10932,N_7619,N_6293);
or U10933 (N_10933,N_8133,N_6746);
nor U10934 (N_10934,N_8502,N_6116);
nor U10935 (N_10935,N_8090,N_6218);
nor U10936 (N_10936,N_7851,N_7795);
or U10937 (N_10937,N_6445,N_7567);
nand U10938 (N_10938,N_8469,N_7926);
or U10939 (N_10939,N_8792,N_8712);
nor U10940 (N_10940,N_8892,N_7468);
and U10941 (N_10941,N_8203,N_8034);
nor U10942 (N_10942,N_7666,N_7176);
nor U10943 (N_10943,N_6639,N_8588);
nand U10944 (N_10944,N_6114,N_7350);
or U10945 (N_10945,N_8034,N_8771);
and U10946 (N_10946,N_8277,N_6839);
and U10947 (N_10947,N_8464,N_8253);
nor U10948 (N_10948,N_8079,N_8403);
and U10949 (N_10949,N_7427,N_8326);
and U10950 (N_10950,N_8037,N_6879);
or U10951 (N_10951,N_6207,N_8809);
and U10952 (N_10952,N_6770,N_6415);
nor U10953 (N_10953,N_8472,N_7280);
or U10954 (N_10954,N_7338,N_7096);
nand U10955 (N_10955,N_6768,N_6183);
and U10956 (N_10956,N_6433,N_8872);
nor U10957 (N_10957,N_6016,N_8185);
nor U10958 (N_10958,N_7643,N_7389);
nor U10959 (N_10959,N_8084,N_6991);
and U10960 (N_10960,N_8297,N_7115);
and U10961 (N_10961,N_8980,N_7804);
nand U10962 (N_10962,N_6705,N_7755);
and U10963 (N_10963,N_6428,N_8392);
and U10964 (N_10964,N_8353,N_6565);
nand U10965 (N_10965,N_7093,N_7946);
or U10966 (N_10966,N_8081,N_8723);
nor U10967 (N_10967,N_7825,N_7744);
and U10968 (N_10968,N_7715,N_8841);
nor U10969 (N_10969,N_7444,N_6635);
or U10970 (N_10970,N_8576,N_6798);
and U10971 (N_10971,N_8569,N_8170);
and U10972 (N_10972,N_7084,N_8532);
nor U10973 (N_10973,N_6281,N_7058);
and U10974 (N_10974,N_7870,N_6011);
or U10975 (N_10975,N_8101,N_8971);
nor U10976 (N_10976,N_7533,N_7332);
nand U10977 (N_10977,N_7226,N_6096);
nor U10978 (N_10978,N_7639,N_8806);
or U10979 (N_10979,N_7288,N_6064);
and U10980 (N_10980,N_8983,N_8932);
nand U10981 (N_10981,N_6868,N_7271);
and U10982 (N_10982,N_6315,N_8915);
and U10983 (N_10983,N_7018,N_6224);
nor U10984 (N_10984,N_8376,N_8869);
and U10985 (N_10985,N_8196,N_7016);
or U10986 (N_10986,N_7033,N_6163);
or U10987 (N_10987,N_7481,N_6029);
and U10988 (N_10988,N_6669,N_6405);
nor U10989 (N_10989,N_8884,N_7400);
nand U10990 (N_10990,N_7205,N_7948);
or U10991 (N_10991,N_7859,N_6632);
nor U10992 (N_10992,N_8751,N_6184);
nor U10993 (N_10993,N_7260,N_8648);
or U10994 (N_10994,N_6839,N_7367);
nor U10995 (N_10995,N_7704,N_7515);
nor U10996 (N_10996,N_7060,N_8558);
and U10997 (N_10997,N_6703,N_8652);
and U10998 (N_10998,N_6751,N_7368);
or U10999 (N_10999,N_6753,N_7930);
and U11000 (N_11000,N_8269,N_8485);
xnor U11001 (N_11001,N_6717,N_7345);
nor U11002 (N_11002,N_8481,N_6337);
nor U11003 (N_11003,N_8764,N_8590);
nor U11004 (N_11004,N_7989,N_7947);
nand U11005 (N_11005,N_8223,N_8978);
nand U11006 (N_11006,N_7635,N_8578);
nand U11007 (N_11007,N_7836,N_7218);
nor U11008 (N_11008,N_8481,N_8785);
nor U11009 (N_11009,N_8432,N_6545);
and U11010 (N_11010,N_7093,N_7173);
nand U11011 (N_11011,N_6413,N_6808);
xnor U11012 (N_11012,N_6679,N_8465);
nor U11013 (N_11013,N_6654,N_8982);
and U11014 (N_11014,N_8446,N_6365);
or U11015 (N_11015,N_7657,N_8460);
or U11016 (N_11016,N_7446,N_6660);
and U11017 (N_11017,N_7024,N_7787);
and U11018 (N_11018,N_7704,N_8329);
and U11019 (N_11019,N_8679,N_7046);
or U11020 (N_11020,N_7281,N_6794);
nand U11021 (N_11021,N_8205,N_8273);
and U11022 (N_11022,N_7549,N_8956);
and U11023 (N_11023,N_6430,N_7303);
or U11024 (N_11024,N_8138,N_7837);
or U11025 (N_11025,N_7071,N_6861);
nor U11026 (N_11026,N_6111,N_8619);
nor U11027 (N_11027,N_6461,N_7460);
nand U11028 (N_11028,N_8707,N_7119);
and U11029 (N_11029,N_7946,N_6278);
or U11030 (N_11030,N_6637,N_8800);
or U11031 (N_11031,N_6303,N_7443);
nor U11032 (N_11032,N_7477,N_8971);
and U11033 (N_11033,N_8097,N_6514);
or U11034 (N_11034,N_6219,N_8928);
and U11035 (N_11035,N_8287,N_6825);
nand U11036 (N_11036,N_8487,N_7147);
nor U11037 (N_11037,N_6118,N_6278);
and U11038 (N_11038,N_8767,N_8619);
nor U11039 (N_11039,N_7023,N_7650);
nand U11040 (N_11040,N_7053,N_8020);
or U11041 (N_11041,N_7134,N_8414);
nor U11042 (N_11042,N_6978,N_7050);
nor U11043 (N_11043,N_6939,N_7933);
nand U11044 (N_11044,N_6704,N_7740);
or U11045 (N_11045,N_6818,N_7102);
nand U11046 (N_11046,N_6051,N_6668);
and U11047 (N_11047,N_6736,N_7435);
nor U11048 (N_11048,N_7996,N_8669);
and U11049 (N_11049,N_6343,N_7772);
and U11050 (N_11050,N_7859,N_8736);
nand U11051 (N_11051,N_7246,N_8010);
nand U11052 (N_11052,N_7189,N_7684);
nor U11053 (N_11053,N_7427,N_8000);
or U11054 (N_11054,N_6336,N_7175);
or U11055 (N_11055,N_6331,N_6426);
nand U11056 (N_11056,N_6277,N_8407);
nor U11057 (N_11057,N_8045,N_6130);
and U11058 (N_11058,N_7240,N_8109);
nor U11059 (N_11059,N_8980,N_8507);
nand U11060 (N_11060,N_7375,N_6900);
nand U11061 (N_11061,N_8575,N_6713);
nand U11062 (N_11062,N_6457,N_7604);
and U11063 (N_11063,N_7283,N_6494);
and U11064 (N_11064,N_7675,N_6553);
nand U11065 (N_11065,N_6685,N_7979);
nor U11066 (N_11066,N_8379,N_7658);
and U11067 (N_11067,N_8625,N_6189);
nand U11068 (N_11068,N_8956,N_8487);
nor U11069 (N_11069,N_6818,N_8978);
nor U11070 (N_11070,N_6904,N_7283);
nor U11071 (N_11071,N_6328,N_7369);
or U11072 (N_11072,N_7665,N_8008);
nor U11073 (N_11073,N_7484,N_7315);
nor U11074 (N_11074,N_6058,N_8803);
or U11075 (N_11075,N_6965,N_7041);
or U11076 (N_11076,N_7039,N_7714);
and U11077 (N_11077,N_8377,N_6858);
nand U11078 (N_11078,N_8583,N_7513);
and U11079 (N_11079,N_7668,N_7979);
and U11080 (N_11080,N_6099,N_6246);
nand U11081 (N_11081,N_6951,N_8712);
or U11082 (N_11082,N_6792,N_7335);
and U11083 (N_11083,N_8087,N_8628);
nand U11084 (N_11084,N_6970,N_8248);
nor U11085 (N_11085,N_6741,N_6558);
nor U11086 (N_11086,N_6111,N_8270);
and U11087 (N_11087,N_7486,N_8163);
nor U11088 (N_11088,N_8730,N_8554);
nor U11089 (N_11089,N_8373,N_7335);
nor U11090 (N_11090,N_8323,N_8851);
xor U11091 (N_11091,N_7865,N_6530);
or U11092 (N_11092,N_7784,N_6254);
nand U11093 (N_11093,N_6789,N_7923);
and U11094 (N_11094,N_7402,N_7387);
nand U11095 (N_11095,N_6968,N_7194);
or U11096 (N_11096,N_7708,N_7464);
or U11097 (N_11097,N_7402,N_8162);
nor U11098 (N_11098,N_6310,N_6841);
nor U11099 (N_11099,N_8757,N_8595);
or U11100 (N_11100,N_7333,N_7579);
or U11101 (N_11101,N_8867,N_7801);
or U11102 (N_11102,N_8270,N_7146);
nand U11103 (N_11103,N_8427,N_7846);
nor U11104 (N_11104,N_7503,N_7642);
and U11105 (N_11105,N_7349,N_7203);
and U11106 (N_11106,N_7248,N_7360);
nand U11107 (N_11107,N_6570,N_7652);
or U11108 (N_11108,N_6250,N_6882);
nor U11109 (N_11109,N_8824,N_7687);
or U11110 (N_11110,N_8785,N_7685);
and U11111 (N_11111,N_8181,N_7368);
and U11112 (N_11112,N_7623,N_8629);
or U11113 (N_11113,N_8462,N_7389);
nor U11114 (N_11114,N_7510,N_8592);
or U11115 (N_11115,N_6087,N_7800);
nor U11116 (N_11116,N_6045,N_7389);
and U11117 (N_11117,N_7871,N_7615);
nor U11118 (N_11118,N_7308,N_7724);
and U11119 (N_11119,N_8846,N_8882);
and U11120 (N_11120,N_7363,N_7489);
and U11121 (N_11121,N_6144,N_8871);
and U11122 (N_11122,N_7888,N_8133);
and U11123 (N_11123,N_7687,N_8347);
and U11124 (N_11124,N_6641,N_7760);
nor U11125 (N_11125,N_7224,N_6685);
nor U11126 (N_11126,N_8634,N_8685);
and U11127 (N_11127,N_6291,N_7722);
or U11128 (N_11128,N_8027,N_6531);
nor U11129 (N_11129,N_6631,N_6767);
nor U11130 (N_11130,N_8154,N_8012);
and U11131 (N_11131,N_6997,N_8869);
or U11132 (N_11132,N_6583,N_8321);
nor U11133 (N_11133,N_8086,N_8577);
nor U11134 (N_11134,N_8257,N_8706);
nor U11135 (N_11135,N_8867,N_6626);
and U11136 (N_11136,N_7345,N_7511);
nand U11137 (N_11137,N_7325,N_7334);
or U11138 (N_11138,N_8206,N_7646);
or U11139 (N_11139,N_7869,N_8848);
nor U11140 (N_11140,N_6486,N_7911);
or U11141 (N_11141,N_7811,N_6393);
and U11142 (N_11142,N_8332,N_8480);
nor U11143 (N_11143,N_7632,N_7983);
or U11144 (N_11144,N_8368,N_7130);
nor U11145 (N_11145,N_8893,N_8212);
and U11146 (N_11146,N_8072,N_6537);
or U11147 (N_11147,N_8047,N_8104);
nand U11148 (N_11148,N_7059,N_8954);
and U11149 (N_11149,N_6896,N_8720);
or U11150 (N_11150,N_8834,N_6770);
and U11151 (N_11151,N_7426,N_7189);
and U11152 (N_11152,N_8698,N_6590);
and U11153 (N_11153,N_8243,N_8404);
and U11154 (N_11154,N_8904,N_8779);
nor U11155 (N_11155,N_7440,N_7500);
and U11156 (N_11156,N_7928,N_7518);
or U11157 (N_11157,N_8669,N_8509);
nor U11158 (N_11158,N_6204,N_8029);
nand U11159 (N_11159,N_8273,N_8069);
and U11160 (N_11160,N_8754,N_7581);
and U11161 (N_11161,N_6847,N_7090);
nor U11162 (N_11162,N_7172,N_6597);
nand U11163 (N_11163,N_7247,N_8700);
and U11164 (N_11164,N_8955,N_8117);
nor U11165 (N_11165,N_8913,N_6240);
and U11166 (N_11166,N_7607,N_7057);
nand U11167 (N_11167,N_8028,N_6651);
or U11168 (N_11168,N_7931,N_6762);
nand U11169 (N_11169,N_7275,N_8759);
nand U11170 (N_11170,N_7385,N_6268);
or U11171 (N_11171,N_7979,N_6139);
and U11172 (N_11172,N_6715,N_6917);
nand U11173 (N_11173,N_7285,N_8630);
or U11174 (N_11174,N_6184,N_7065);
and U11175 (N_11175,N_6230,N_6922);
and U11176 (N_11176,N_7420,N_6597);
and U11177 (N_11177,N_8275,N_7211);
xor U11178 (N_11178,N_7911,N_7069);
or U11179 (N_11179,N_7217,N_8907);
nand U11180 (N_11180,N_6020,N_6510);
or U11181 (N_11181,N_8132,N_7338);
and U11182 (N_11182,N_7953,N_8954);
and U11183 (N_11183,N_8312,N_8963);
or U11184 (N_11184,N_6002,N_7267);
nand U11185 (N_11185,N_6144,N_7165);
nand U11186 (N_11186,N_6490,N_6588);
or U11187 (N_11187,N_8729,N_6863);
and U11188 (N_11188,N_7696,N_8246);
nand U11189 (N_11189,N_6587,N_7647);
or U11190 (N_11190,N_8995,N_7602);
nand U11191 (N_11191,N_8726,N_6257);
nor U11192 (N_11192,N_7635,N_8704);
and U11193 (N_11193,N_7534,N_7980);
nand U11194 (N_11194,N_6064,N_6982);
nor U11195 (N_11195,N_6740,N_8138);
nor U11196 (N_11196,N_7938,N_6366);
and U11197 (N_11197,N_6017,N_7648);
and U11198 (N_11198,N_6403,N_6767);
nand U11199 (N_11199,N_8175,N_8021);
nand U11200 (N_11200,N_8304,N_6792);
nand U11201 (N_11201,N_8909,N_7863);
or U11202 (N_11202,N_8005,N_7492);
nand U11203 (N_11203,N_7769,N_7207);
and U11204 (N_11204,N_7233,N_8774);
nor U11205 (N_11205,N_7462,N_7195);
and U11206 (N_11206,N_7251,N_7857);
or U11207 (N_11207,N_8220,N_6718);
nor U11208 (N_11208,N_6140,N_8542);
nor U11209 (N_11209,N_7994,N_8099);
nand U11210 (N_11210,N_6224,N_7816);
nand U11211 (N_11211,N_8289,N_6782);
nor U11212 (N_11212,N_8434,N_8664);
and U11213 (N_11213,N_6121,N_8768);
nor U11214 (N_11214,N_8875,N_6645);
nor U11215 (N_11215,N_7565,N_8700);
and U11216 (N_11216,N_8246,N_6090);
and U11217 (N_11217,N_7738,N_8591);
and U11218 (N_11218,N_8449,N_6448);
nor U11219 (N_11219,N_8259,N_8382);
or U11220 (N_11220,N_8800,N_7057);
or U11221 (N_11221,N_8839,N_8812);
or U11222 (N_11222,N_7592,N_7202);
nand U11223 (N_11223,N_8524,N_6440);
and U11224 (N_11224,N_8815,N_7811);
nor U11225 (N_11225,N_6439,N_7912);
nand U11226 (N_11226,N_8167,N_6361);
and U11227 (N_11227,N_7282,N_8995);
nand U11228 (N_11228,N_8327,N_8265);
nand U11229 (N_11229,N_7165,N_7049);
and U11230 (N_11230,N_6995,N_6709);
or U11231 (N_11231,N_6536,N_8524);
and U11232 (N_11232,N_8536,N_7041);
nor U11233 (N_11233,N_8478,N_6526);
xnor U11234 (N_11234,N_7098,N_6409);
nor U11235 (N_11235,N_8053,N_6218);
nor U11236 (N_11236,N_8315,N_7418);
nand U11237 (N_11237,N_8531,N_6878);
nor U11238 (N_11238,N_6521,N_6085);
nor U11239 (N_11239,N_8117,N_7958);
or U11240 (N_11240,N_6064,N_8746);
or U11241 (N_11241,N_7146,N_8017);
or U11242 (N_11242,N_7311,N_7332);
or U11243 (N_11243,N_7767,N_8308);
and U11244 (N_11244,N_8294,N_6516);
nand U11245 (N_11245,N_6326,N_8181);
nor U11246 (N_11246,N_6308,N_6913);
and U11247 (N_11247,N_8895,N_8795);
nor U11248 (N_11248,N_8042,N_7872);
or U11249 (N_11249,N_7064,N_8335);
nor U11250 (N_11250,N_7770,N_8324);
nor U11251 (N_11251,N_7945,N_8540);
and U11252 (N_11252,N_8318,N_7583);
or U11253 (N_11253,N_7597,N_7206);
or U11254 (N_11254,N_8953,N_6377);
or U11255 (N_11255,N_6484,N_8400);
and U11256 (N_11256,N_8721,N_8496);
and U11257 (N_11257,N_7675,N_6722);
nor U11258 (N_11258,N_7566,N_7576);
or U11259 (N_11259,N_7547,N_7431);
nor U11260 (N_11260,N_8244,N_6681);
and U11261 (N_11261,N_8031,N_6695);
nor U11262 (N_11262,N_6435,N_7592);
or U11263 (N_11263,N_7389,N_8214);
and U11264 (N_11264,N_7088,N_8733);
nor U11265 (N_11265,N_7478,N_6585);
nand U11266 (N_11266,N_6142,N_7633);
nor U11267 (N_11267,N_8284,N_7651);
and U11268 (N_11268,N_7080,N_6870);
nor U11269 (N_11269,N_6773,N_7092);
and U11270 (N_11270,N_8103,N_7951);
nand U11271 (N_11271,N_8626,N_6895);
and U11272 (N_11272,N_7746,N_7025);
or U11273 (N_11273,N_8007,N_7908);
nor U11274 (N_11274,N_7294,N_7072);
nor U11275 (N_11275,N_8023,N_6354);
and U11276 (N_11276,N_7111,N_6485);
or U11277 (N_11277,N_8963,N_7943);
nor U11278 (N_11278,N_6447,N_7813);
nand U11279 (N_11279,N_6297,N_6038);
nor U11280 (N_11280,N_6138,N_7321);
or U11281 (N_11281,N_6833,N_6658);
nor U11282 (N_11282,N_7478,N_7437);
or U11283 (N_11283,N_6128,N_7214);
or U11284 (N_11284,N_6765,N_6663);
nor U11285 (N_11285,N_6053,N_8424);
nor U11286 (N_11286,N_8158,N_7702);
or U11287 (N_11287,N_7219,N_6741);
and U11288 (N_11288,N_8151,N_7148);
xnor U11289 (N_11289,N_8677,N_8699);
and U11290 (N_11290,N_6914,N_7509);
nand U11291 (N_11291,N_7957,N_8962);
or U11292 (N_11292,N_8902,N_6976);
nand U11293 (N_11293,N_6014,N_8379);
nand U11294 (N_11294,N_6497,N_7749);
or U11295 (N_11295,N_7568,N_7438);
or U11296 (N_11296,N_6344,N_6131);
nand U11297 (N_11297,N_7130,N_6845);
nand U11298 (N_11298,N_7595,N_7937);
or U11299 (N_11299,N_8975,N_7866);
nand U11300 (N_11300,N_7935,N_6711);
nor U11301 (N_11301,N_7859,N_8025);
and U11302 (N_11302,N_7378,N_8850);
nor U11303 (N_11303,N_8121,N_6994);
nor U11304 (N_11304,N_7098,N_6195);
and U11305 (N_11305,N_8146,N_6571);
or U11306 (N_11306,N_7133,N_8368);
nand U11307 (N_11307,N_8017,N_8301);
nand U11308 (N_11308,N_8065,N_7850);
nand U11309 (N_11309,N_8600,N_8705);
nor U11310 (N_11310,N_6990,N_6939);
nand U11311 (N_11311,N_7386,N_6432);
and U11312 (N_11312,N_7581,N_6451);
nand U11313 (N_11313,N_7531,N_8608);
nor U11314 (N_11314,N_7211,N_8390);
nor U11315 (N_11315,N_6974,N_8480);
and U11316 (N_11316,N_7205,N_7876);
nand U11317 (N_11317,N_8958,N_7905);
nand U11318 (N_11318,N_8484,N_6461);
nor U11319 (N_11319,N_7668,N_8881);
nor U11320 (N_11320,N_6546,N_8126);
nor U11321 (N_11321,N_7260,N_7348);
and U11322 (N_11322,N_7474,N_6627);
nor U11323 (N_11323,N_8872,N_6068);
nor U11324 (N_11324,N_7000,N_7956);
nor U11325 (N_11325,N_6982,N_8771);
nand U11326 (N_11326,N_7475,N_6924);
nand U11327 (N_11327,N_6429,N_8891);
nand U11328 (N_11328,N_8846,N_8445);
or U11329 (N_11329,N_8027,N_8247);
nor U11330 (N_11330,N_8484,N_6792);
and U11331 (N_11331,N_6693,N_7066);
xor U11332 (N_11332,N_7536,N_8804);
or U11333 (N_11333,N_7885,N_8859);
or U11334 (N_11334,N_6058,N_6268);
or U11335 (N_11335,N_6313,N_8013);
and U11336 (N_11336,N_8351,N_7513);
nand U11337 (N_11337,N_8294,N_6272);
nor U11338 (N_11338,N_6839,N_7167);
or U11339 (N_11339,N_8617,N_8722);
nor U11340 (N_11340,N_8627,N_8538);
and U11341 (N_11341,N_8033,N_6180);
nor U11342 (N_11342,N_6683,N_7649);
or U11343 (N_11343,N_6805,N_7727);
nand U11344 (N_11344,N_6660,N_7453);
nor U11345 (N_11345,N_6731,N_8727);
or U11346 (N_11346,N_6347,N_6435);
nand U11347 (N_11347,N_8110,N_7325);
nor U11348 (N_11348,N_8089,N_7868);
nor U11349 (N_11349,N_7263,N_8643);
or U11350 (N_11350,N_7987,N_6927);
nor U11351 (N_11351,N_6628,N_7274);
and U11352 (N_11352,N_8050,N_8786);
or U11353 (N_11353,N_7110,N_7225);
or U11354 (N_11354,N_7126,N_6114);
nand U11355 (N_11355,N_7426,N_8591);
or U11356 (N_11356,N_6042,N_6655);
and U11357 (N_11357,N_8549,N_7707);
nand U11358 (N_11358,N_8061,N_7667);
nor U11359 (N_11359,N_7045,N_8765);
or U11360 (N_11360,N_8623,N_7701);
nor U11361 (N_11361,N_7217,N_7255);
nand U11362 (N_11362,N_8810,N_8303);
and U11363 (N_11363,N_8419,N_7689);
or U11364 (N_11364,N_7627,N_7947);
or U11365 (N_11365,N_7422,N_7630);
or U11366 (N_11366,N_6640,N_8312);
nor U11367 (N_11367,N_6198,N_8633);
or U11368 (N_11368,N_6264,N_7607);
or U11369 (N_11369,N_7621,N_7528);
nand U11370 (N_11370,N_7475,N_7220);
and U11371 (N_11371,N_7594,N_8172);
nor U11372 (N_11372,N_7140,N_8514);
xnor U11373 (N_11373,N_8085,N_8225);
and U11374 (N_11374,N_7017,N_6006);
and U11375 (N_11375,N_6521,N_8605);
or U11376 (N_11376,N_6256,N_7227);
and U11377 (N_11377,N_7632,N_8773);
and U11378 (N_11378,N_8520,N_6448);
nor U11379 (N_11379,N_7142,N_7837);
or U11380 (N_11380,N_8227,N_6837);
and U11381 (N_11381,N_7306,N_8381);
nand U11382 (N_11382,N_8425,N_7840);
nor U11383 (N_11383,N_7620,N_8266);
nor U11384 (N_11384,N_6543,N_8420);
nand U11385 (N_11385,N_7763,N_7487);
and U11386 (N_11386,N_8285,N_7047);
nor U11387 (N_11387,N_8245,N_7625);
nand U11388 (N_11388,N_6139,N_8606);
and U11389 (N_11389,N_8637,N_8488);
nor U11390 (N_11390,N_6782,N_7191);
and U11391 (N_11391,N_8018,N_6045);
or U11392 (N_11392,N_8417,N_7913);
or U11393 (N_11393,N_8551,N_7556);
or U11394 (N_11394,N_7847,N_6876);
or U11395 (N_11395,N_7097,N_7358);
nor U11396 (N_11396,N_7159,N_8376);
and U11397 (N_11397,N_7964,N_8009);
nor U11398 (N_11398,N_6003,N_8750);
nand U11399 (N_11399,N_6136,N_7503);
nand U11400 (N_11400,N_6925,N_6693);
nand U11401 (N_11401,N_7052,N_7033);
and U11402 (N_11402,N_8347,N_8399);
or U11403 (N_11403,N_6275,N_7459);
nor U11404 (N_11404,N_6942,N_7499);
nor U11405 (N_11405,N_6192,N_7810);
and U11406 (N_11406,N_8467,N_7359);
nor U11407 (N_11407,N_6466,N_6826);
nor U11408 (N_11408,N_7312,N_7659);
and U11409 (N_11409,N_7327,N_8980);
nand U11410 (N_11410,N_6288,N_8212);
nand U11411 (N_11411,N_7827,N_6219);
nand U11412 (N_11412,N_8863,N_7595);
nor U11413 (N_11413,N_8696,N_7570);
nor U11414 (N_11414,N_7747,N_8793);
nor U11415 (N_11415,N_7948,N_7215);
and U11416 (N_11416,N_6062,N_8096);
nor U11417 (N_11417,N_7072,N_8660);
or U11418 (N_11418,N_7427,N_6739);
nand U11419 (N_11419,N_8582,N_7643);
and U11420 (N_11420,N_8361,N_6225);
and U11421 (N_11421,N_6063,N_8401);
and U11422 (N_11422,N_8318,N_8122);
nand U11423 (N_11423,N_6264,N_6297);
or U11424 (N_11424,N_6321,N_7077);
nor U11425 (N_11425,N_7920,N_6043);
nand U11426 (N_11426,N_6040,N_8126);
and U11427 (N_11427,N_6968,N_8102);
or U11428 (N_11428,N_6244,N_6521);
or U11429 (N_11429,N_8457,N_8481);
nor U11430 (N_11430,N_8248,N_8027);
nor U11431 (N_11431,N_6822,N_6867);
and U11432 (N_11432,N_7468,N_6731);
nor U11433 (N_11433,N_6332,N_7369);
and U11434 (N_11434,N_6337,N_6401);
and U11435 (N_11435,N_8304,N_7390);
or U11436 (N_11436,N_7298,N_6985);
and U11437 (N_11437,N_7086,N_7640);
or U11438 (N_11438,N_6074,N_6143);
nand U11439 (N_11439,N_8864,N_7066);
or U11440 (N_11440,N_8110,N_6861);
or U11441 (N_11441,N_7880,N_7636);
and U11442 (N_11442,N_8162,N_8386);
nand U11443 (N_11443,N_8902,N_6042);
nor U11444 (N_11444,N_6282,N_7707);
and U11445 (N_11445,N_6829,N_6537);
or U11446 (N_11446,N_7355,N_6836);
and U11447 (N_11447,N_7901,N_7470);
nand U11448 (N_11448,N_6935,N_7065);
or U11449 (N_11449,N_8882,N_7694);
or U11450 (N_11450,N_7411,N_7511);
nand U11451 (N_11451,N_7682,N_7961);
nor U11452 (N_11452,N_8449,N_8990);
and U11453 (N_11453,N_8173,N_8566);
xor U11454 (N_11454,N_6222,N_6461);
and U11455 (N_11455,N_6023,N_7118);
nand U11456 (N_11456,N_7907,N_6401);
xor U11457 (N_11457,N_8232,N_6719);
nand U11458 (N_11458,N_6480,N_6285);
nand U11459 (N_11459,N_6164,N_7451);
nand U11460 (N_11460,N_7406,N_8262);
nand U11461 (N_11461,N_6028,N_7020);
nor U11462 (N_11462,N_7722,N_8971);
or U11463 (N_11463,N_6917,N_7103);
nand U11464 (N_11464,N_6187,N_7949);
or U11465 (N_11465,N_7504,N_7633);
and U11466 (N_11466,N_6835,N_8158);
nand U11467 (N_11467,N_8493,N_6929);
nor U11468 (N_11468,N_8272,N_6976);
nand U11469 (N_11469,N_8998,N_8570);
or U11470 (N_11470,N_8440,N_8301);
or U11471 (N_11471,N_6046,N_6771);
and U11472 (N_11472,N_7595,N_8154);
and U11473 (N_11473,N_7395,N_6317);
or U11474 (N_11474,N_8417,N_8155);
nand U11475 (N_11475,N_7516,N_8485);
or U11476 (N_11476,N_6466,N_6908);
and U11477 (N_11477,N_7012,N_8921);
xnor U11478 (N_11478,N_8641,N_7865);
nand U11479 (N_11479,N_8147,N_7210);
or U11480 (N_11480,N_7515,N_7723);
or U11481 (N_11481,N_7516,N_8868);
nor U11482 (N_11482,N_6203,N_6610);
nand U11483 (N_11483,N_7692,N_7630);
nand U11484 (N_11484,N_8471,N_6213);
nand U11485 (N_11485,N_7180,N_7904);
or U11486 (N_11486,N_7504,N_6992);
nand U11487 (N_11487,N_8144,N_8297);
nand U11488 (N_11488,N_6479,N_8972);
or U11489 (N_11489,N_7755,N_6535);
and U11490 (N_11490,N_8598,N_7538);
and U11491 (N_11491,N_6229,N_6536);
nor U11492 (N_11492,N_8028,N_8772);
nand U11493 (N_11493,N_8277,N_7220);
nor U11494 (N_11494,N_8821,N_7056);
nand U11495 (N_11495,N_8436,N_8257);
or U11496 (N_11496,N_7197,N_7309);
or U11497 (N_11497,N_7474,N_8009);
nor U11498 (N_11498,N_7219,N_7488);
nand U11499 (N_11499,N_6003,N_8955);
nor U11500 (N_11500,N_7861,N_7656);
nor U11501 (N_11501,N_6590,N_8589);
nand U11502 (N_11502,N_7425,N_8784);
nand U11503 (N_11503,N_6998,N_7379);
and U11504 (N_11504,N_7124,N_6049);
or U11505 (N_11505,N_8602,N_8925);
nand U11506 (N_11506,N_7003,N_7363);
xnor U11507 (N_11507,N_8976,N_6779);
nand U11508 (N_11508,N_7222,N_7293);
nor U11509 (N_11509,N_8480,N_6039);
nor U11510 (N_11510,N_6258,N_7950);
or U11511 (N_11511,N_8729,N_6300);
and U11512 (N_11512,N_8618,N_8184);
and U11513 (N_11513,N_7429,N_8439);
nor U11514 (N_11514,N_7280,N_6340);
nor U11515 (N_11515,N_6426,N_8884);
nand U11516 (N_11516,N_6006,N_7729);
or U11517 (N_11517,N_7220,N_8854);
and U11518 (N_11518,N_7782,N_6838);
nand U11519 (N_11519,N_6537,N_7752);
or U11520 (N_11520,N_6234,N_8115);
and U11521 (N_11521,N_7835,N_7605);
nand U11522 (N_11522,N_8681,N_8255);
and U11523 (N_11523,N_8184,N_8013);
and U11524 (N_11524,N_8945,N_7899);
or U11525 (N_11525,N_7549,N_7599);
or U11526 (N_11526,N_6703,N_6239);
nor U11527 (N_11527,N_8427,N_7991);
nor U11528 (N_11528,N_7243,N_7858);
nand U11529 (N_11529,N_7596,N_8650);
and U11530 (N_11530,N_7919,N_6491);
and U11531 (N_11531,N_6759,N_6658);
or U11532 (N_11532,N_6621,N_7668);
nand U11533 (N_11533,N_8588,N_7402);
and U11534 (N_11534,N_7667,N_8212);
or U11535 (N_11535,N_6842,N_6544);
nor U11536 (N_11536,N_7788,N_8834);
nand U11537 (N_11537,N_8657,N_6336);
or U11538 (N_11538,N_7481,N_6916);
nand U11539 (N_11539,N_6339,N_8700);
nand U11540 (N_11540,N_8519,N_6181);
or U11541 (N_11541,N_7012,N_8386);
nand U11542 (N_11542,N_7616,N_8324);
nand U11543 (N_11543,N_7985,N_8837);
or U11544 (N_11544,N_8028,N_7198);
nand U11545 (N_11545,N_8342,N_8204);
and U11546 (N_11546,N_8833,N_8985);
and U11547 (N_11547,N_6529,N_6187);
nand U11548 (N_11548,N_6536,N_7682);
nand U11549 (N_11549,N_8650,N_6044);
nand U11550 (N_11550,N_6021,N_7403);
nand U11551 (N_11551,N_6578,N_7987);
and U11552 (N_11552,N_6637,N_6414);
or U11553 (N_11553,N_7787,N_6059);
nor U11554 (N_11554,N_6216,N_6783);
nand U11555 (N_11555,N_7623,N_7843);
or U11556 (N_11556,N_6875,N_8386);
and U11557 (N_11557,N_8457,N_8625);
or U11558 (N_11558,N_8715,N_7873);
or U11559 (N_11559,N_8815,N_7761);
or U11560 (N_11560,N_7414,N_8497);
nand U11561 (N_11561,N_8661,N_6527);
nor U11562 (N_11562,N_6388,N_8896);
or U11563 (N_11563,N_7535,N_6253);
and U11564 (N_11564,N_6745,N_6268);
and U11565 (N_11565,N_6302,N_7516);
nand U11566 (N_11566,N_6231,N_8129);
and U11567 (N_11567,N_7647,N_6019);
and U11568 (N_11568,N_8686,N_7239);
nor U11569 (N_11569,N_7126,N_6568);
or U11570 (N_11570,N_7436,N_6924);
nor U11571 (N_11571,N_7025,N_6231);
nand U11572 (N_11572,N_6362,N_7125);
or U11573 (N_11573,N_8234,N_8500);
and U11574 (N_11574,N_6978,N_8472);
nand U11575 (N_11575,N_7734,N_8039);
and U11576 (N_11576,N_7074,N_7674);
or U11577 (N_11577,N_8455,N_7007);
nand U11578 (N_11578,N_6738,N_7871);
or U11579 (N_11579,N_7068,N_8718);
and U11580 (N_11580,N_7998,N_8353);
nand U11581 (N_11581,N_6523,N_7739);
and U11582 (N_11582,N_8675,N_8891);
and U11583 (N_11583,N_8793,N_8439);
or U11584 (N_11584,N_7149,N_8034);
nor U11585 (N_11585,N_8132,N_7070);
or U11586 (N_11586,N_8026,N_6988);
and U11587 (N_11587,N_6546,N_6248);
and U11588 (N_11588,N_7776,N_8594);
and U11589 (N_11589,N_7053,N_6195);
and U11590 (N_11590,N_6236,N_7324);
or U11591 (N_11591,N_7159,N_8452);
and U11592 (N_11592,N_8460,N_6697);
nor U11593 (N_11593,N_8313,N_7610);
nor U11594 (N_11594,N_8431,N_6864);
or U11595 (N_11595,N_8621,N_7577);
nor U11596 (N_11596,N_6706,N_7808);
nand U11597 (N_11597,N_7886,N_8702);
nor U11598 (N_11598,N_7013,N_6196);
nor U11599 (N_11599,N_8941,N_8969);
or U11600 (N_11600,N_6579,N_8698);
nand U11601 (N_11601,N_6397,N_8925);
or U11602 (N_11602,N_6557,N_8858);
or U11603 (N_11603,N_6364,N_7024);
or U11604 (N_11604,N_8518,N_6358);
or U11605 (N_11605,N_7897,N_6485);
nand U11606 (N_11606,N_6132,N_8758);
nand U11607 (N_11607,N_7464,N_7532);
nand U11608 (N_11608,N_7215,N_8383);
nand U11609 (N_11609,N_7827,N_6822);
nor U11610 (N_11610,N_6161,N_6183);
nor U11611 (N_11611,N_8714,N_6281);
nand U11612 (N_11612,N_6038,N_7661);
and U11613 (N_11613,N_8048,N_8802);
and U11614 (N_11614,N_8148,N_7618);
and U11615 (N_11615,N_7699,N_7199);
nand U11616 (N_11616,N_6258,N_7325);
nor U11617 (N_11617,N_6899,N_7341);
and U11618 (N_11618,N_7934,N_7396);
and U11619 (N_11619,N_8026,N_6818);
or U11620 (N_11620,N_7778,N_7280);
and U11621 (N_11621,N_7723,N_8703);
and U11622 (N_11622,N_8793,N_7946);
nand U11623 (N_11623,N_7506,N_8430);
nor U11624 (N_11624,N_8804,N_7812);
and U11625 (N_11625,N_7611,N_6143);
or U11626 (N_11626,N_6949,N_8903);
nand U11627 (N_11627,N_8483,N_8041);
nor U11628 (N_11628,N_7708,N_6047);
or U11629 (N_11629,N_6568,N_7244);
nor U11630 (N_11630,N_7706,N_8165);
or U11631 (N_11631,N_8899,N_8813);
or U11632 (N_11632,N_6701,N_7876);
nor U11633 (N_11633,N_6329,N_6833);
and U11634 (N_11634,N_8311,N_8769);
nand U11635 (N_11635,N_6326,N_8953);
nand U11636 (N_11636,N_7457,N_8679);
nand U11637 (N_11637,N_7927,N_8993);
nor U11638 (N_11638,N_8482,N_8046);
or U11639 (N_11639,N_6164,N_7876);
and U11640 (N_11640,N_7149,N_7342);
or U11641 (N_11641,N_7915,N_7080);
or U11642 (N_11642,N_6420,N_7743);
nand U11643 (N_11643,N_8228,N_8002);
nor U11644 (N_11644,N_8781,N_7181);
or U11645 (N_11645,N_7464,N_6291);
nor U11646 (N_11646,N_7997,N_8430);
and U11647 (N_11647,N_6861,N_6380);
nor U11648 (N_11648,N_7412,N_7353);
nor U11649 (N_11649,N_6559,N_6431);
nand U11650 (N_11650,N_7247,N_7075);
nor U11651 (N_11651,N_6405,N_8713);
and U11652 (N_11652,N_8260,N_8257);
and U11653 (N_11653,N_6618,N_8896);
nor U11654 (N_11654,N_6032,N_8304);
nand U11655 (N_11655,N_8740,N_7295);
nor U11656 (N_11656,N_8093,N_6063);
nand U11657 (N_11657,N_8938,N_7913);
or U11658 (N_11658,N_7914,N_8511);
or U11659 (N_11659,N_8336,N_6157);
and U11660 (N_11660,N_7563,N_6934);
nor U11661 (N_11661,N_8482,N_7687);
nor U11662 (N_11662,N_6365,N_7039);
or U11663 (N_11663,N_8309,N_7252);
and U11664 (N_11664,N_7774,N_7988);
and U11665 (N_11665,N_8912,N_7052);
or U11666 (N_11666,N_8902,N_8581);
and U11667 (N_11667,N_7488,N_8926);
or U11668 (N_11668,N_8319,N_7350);
nand U11669 (N_11669,N_8230,N_6198);
nor U11670 (N_11670,N_8217,N_6347);
nand U11671 (N_11671,N_7670,N_7355);
nor U11672 (N_11672,N_6679,N_6041);
nand U11673 (N_11673,N_8533,N_6948);
nor U11674 (N_11674,N_7588,N_7085);
nor U11675 (N_11675,N_6503,N_7435);
or U11676 (N_11676,N_8762,N_7005);
or U11677 (N_11677,N_7999,N_7438);
nand U11678 (N_11678,N_6392,N_8708);
nand U11679 (N_11679,N_8575,N_8150);
nand U11680 (N_11680,N_6589,N_6252);
nor U11681 (N_11681,N_8599,N_7792);
or U11682 (N_11682,N_7181,N_8754);
xnor U11683 (N_11683,N_7101,N_6517);
or U11684 (N_11684,N_7498,N_6660);
nor U11685 (N_11685,N_8359,N_8773);
nor U11686 (N_11686,N_8140,N_6931);
nor U11687 (N_11687,N_7336,N_6131);
nand U11688 (N_11688,N_8380,N_7021);
and U11689 (N_11689,N_6168,N_7188);
nor U11690 (N_11690,N_7562,N_6626);
or U11691 (N_11691,N_7544,N_6284);
and U11692 (N_11692,N_6158,N_8516);
and U11693 (N_11693,N_7381,N_6931);
nand U11694 (N_11694,N_8070,N_8038);
nand U11695 (N_11695,N_6278,N_7810);
or U11696 (N_11696,N_6680,N_8661);
or U11697 (N_11697,N_8358,N_7765);
nand U11698 (N_11698,N_6474,N_6499);
or U11699 (N_11699,N_6962,N_6833);
nor U11700 (N_11700,N_8120,N_8932);
and U11701 (N_11701,N_7951,N_6060);
nor U11702 (N_11702,N_6903,N_8817);
and U11703 (N_11703,N_6081,N_6529);
and U11704 (N_11704,N_6582,N_8101);
or U11705 (N_11705,N_8229,N_7962);
nor U11706 (N_11706,N_7059,N_7856);
nand U11707 (N_11707,N_7582,N_7354);
nand U11708 (N_11708,N_6905,N_8751);
nand U11709 (N_11709,N_7910,N_6871);
and U11710 (N_11710,N_6532,N_7923);
nor U11711 (N_11711,N_6635,N_7527);
and U11712 (N_11712,N_7112,N_7491);
nor U11713 (N_11713,N_8218,N_7852);
or U11714 (N_11714,N_8988,N_7504);
and U11715 (N_11715,N_8678,N_6217);
and U11716 (N_11716,N_6081,N_8997);
and U11717 (N_11717,N_7926,N_6339);
and U11718 (N_11718,N_7273,N_7659);
or U11719 (N_11719,N_8645,N_7237);
nor U11720 (N_11720,N_6396,N_8912);
and U11721 (N_11721,N_6443,N_6834);
or U11722 (N_11722,N_8523,N_6242);
nor U11723 (N_11723,N_7785,N_8355);
or U11724 (N_11724,N_8695,N_6542);
and U11725 (N_11725,N_6139,N_7233);
and U11726 (N_11726,N_7777,N_8325);
xor U11727 (N_11727,N_8346,N_7909);
nor U11728 (N_11728,N_7447,N_8648);
nor U11729 (N_11729,N_8144,N_6994);
or U11730 (N_11730,N_8901,N_6935);
nand U11731 (N_11731,N_7096,N_6353);
nand U11732 (N_11732,N_7770,N_6643);
nor U11733 (N_11733,N_7218,N_7869);
nor U11734 (N_11734,N_6694,N_7827);
nor U11735 (N_11735,N_8906,N_8039);
and U11736 (N_11736,N_6901,N_7357);
nand U11737 (N_11737,N_7480,N_8096);
and U11738 (N_11738,N_7271,N_8513);
and U11739 (N_11739,N_7026,N_8316);
or U11740 (N_11740,N_6681,N_6082);
and U11741 (N_11741,N_6041,N_8253);
or U11742 (N_11742,N_7466,N_7848);
or U11743 (N_11743,N_6023,N_7273);
and U11744 (N_11744,N_7199,N_7634);
nor U11745 (N_11745,N_8483,N_7684);
nand U11746 (N_11746,N_8342,N_6929);
nor U11747 (N_11747,N_8182,N_8092);
and U11748 (N_11748,N_6439,N_8810);
nand U11749 (N_11749,N_7164,N_6671);
nand U11750 (N_11750,N_8214,N_6862);
nand U11751 (N_11751,N_6405,N_6782);
or U11752 (N_11752,N_8735,N_6958);
nand U11753 (N_11753,N_8144,N_7452);
or U11754 (N_11754,N_7729,N_8987);
and U11755 (N_11755,N_7054,N_8253);
nand U11756 (N_11756,N_8532,N_6359);
or U11757 (N_11757,N_7592,N_8856);
and U11758 (N_11758,N_7574,N_7956);
nor U11759 (N_11759,N_8885,N_8206);
nand U11760 (N_11760,N_8083,N_7127);
nor U11761 (N_11761,N_7641,N_7008);
nand U11762 (N_11762,N_6065,N_8122);
or U11763 (N_11763,N_8627,N_8734);
and U11764 (N_11764,N_8032,N_7842);
nand U11765 (N_11765,N_6827,N_7146);
and U11766 (N_11766,N_6720,N_8807);
and U11767 (N_11767,N_6736,N_6888);
and U11768 (N_11768,N_7344,N_7998);
nor U11769 (N_11769,N_7993,N_8507);
and U11770 (N_11770,N_7026,N_8178);
and U11771 (N_11771,N_8324,N_8268);
or U11772 (N_11772,N_6943,N_7670);
or U11773 (N_11773,N_7950,N_6864);
and U11774 (N_11774,N_6213,N_6968);
or U11775 (N_11775,N_8917,N_6125);
or U11776 (N_11776,N_6032,N_6325);
and U11777 (N_11777,N_8580,N_7483);
nor U11778 (N_11778,N_7613,N_7432);
and U11779 (N_11779,N_8503,N_8312);
nor U11780 (N_11780,N_7671,N_6715);
or U11781 (N_11781,N_8687,N_7563);
or U11782 (N_11782,N_8668,N_6694);
and U11783 (N_11783,N_6832,N_6219);
nand U11784 (N_11784,N_7102,N_7939);
or U11785 (N_11785,N_6320,N_8303);
xnor U11786 (N_11786,N_8898,N_8581);
and U11787 (N_11787,N_6094,N_8481);
nand U11788 (N_11788,N_6538,N_6579);
nand U11789 (N_11789,N_6844,N_6318);
or U11790 (N_11790,N_6633,N_6794);
nor U11791 (N_11791,N_7593,N_7791);
nand U11792 (N_11792,N_8338,N_6106);
nand U11793 (N_11793,N_7353,N_7690);
nor U11794 (N_11794,N_7575,N_7441);
xnor U11795 (N_11795,N_6696,N_8633);
or U11796 (N_11796,N_7392,N_7519);
nor U11797 (N_11797,N_7777,N_7290);
nor U11798 (N_11798,N_6981,N_7081);
or U11799 (N_11799,N_7213,N_8606);
and U11800 (N_11800,N_7770,N_6794);
or U11801 (N_11801,N_7253,N_8304);
nand U11802 (N_11802,N_7932,N_8172);
nor U11803 (N_11803,N_8352,N_8935);
nor U11804 (N_11804,N_8917,N_7274);
nand U11805 (N_11805,N_8522,N_6570);
or U11806 (N_11806,N_7930,N_7619);
and U11807 (N_11807,N_7716,N_7951);
nor U11808 (N_11808,N_8472,N_6930);
or U11809 (N_11809,N_6274,N_7396);
nand U11810 (N_11810,N_8034,N_7746);
nor U11811 (N_11811,N_8060,N_8019);
and U11812 (N_11812,N_7901,N_6797);
nor U11813 (N_11813,N_8178,N_8710);
nand U11814 (N_11814,N_8297,N_8749);
nand U11815 (N_11815,N_7840,N_8018);
or U11816 (N_11816,N_6145,N_8963);
or U11817 (N_11817,N_6218,N_8564);
and U11818 (N_11818,N_6548,N_8454);
nand U11819 (N_11819,N_6084,N_8973);
and U11820 (N_11820,N_6933,N_8055);
nor U11821 (N_11821,N_7773,N_6058);
and U11822 (N_11822,N_7309,N_6806);
or U11823 (N_11823,N_8430,N_6661);
or U11824 (N_11824,N_7754,N_6149);
xor U11825 (N_11825,N_8279,N_7198);
nor U11826 (N_11826,N_8132,N_8565);
and U11827 (N_11827,N_7670,N_8216);
nor U11828 (N_11828,N_7087,N_7292);
nand U11829 (N_11829,N_6547,N_8418);
or U11830 (N_11830,N_6023,N_6571);
nand U11831 (N_11831,N_7081,N_6987);
or U11832 (N_11832,N_8513,N_6689);
nor U11833 (N_11833,N_8229,N_8211);
or U11834 (N_11834,N_7092,N_8245);
nand U11835 (N_11835,N_6457,N_7242);
nand U11836 (N_11836,N_6167,N_6991);
or U11837 (N_11837,N_6536,N_6467);
nand U11838 (N_11838,N_8483,N_6589);
or U11839 (N_11839,N_6927,N_6977);
nor U11840 (N_11840,N_6168,N_6516);
or U11841 (N_11841,N_6798,N_6634);
nor U11842 (N_11842,N_6337,N_8807);
or U11843 (N_11843,N_8747,N_7709);
and U11844 (N_11844,N_8919,N_8507);
or U11845 (N_11845,N_6166,N_7189);
and U11846 (N_11846,N_6431,N_6843);
and U11847 (N_11847,N_8826,N_8937);
and U11848 (N_11848,N_6971,N_6626);
and U11849 (N_11849,N_6085,N_7875);
and U11850 (N_11850,N_7059,N_8347);
or U11851 (N_11851,N_8174,N_7350);
nor U11852 (N_11852,N_6350,N_8428);
nor U11853 (N_11853,N_7575,N_6561);
or U11854 (N_11854,N_8707,N_6356);
xor U11855 (N_11855,N_8546,N_6179);
nand U11856 (N_11856,N_6363,N_7127);
or U11857 (N_11857,N_6441,N_8457);
and U11858 (N_11858,N_8078,N_7200);
nand U11859 (N_11859,N_7839,N_8545);
and U11860 (N_11860,N_8417,N_7003);
or U11861 (N_11861,N_8978,N_7957);
nor U11862 (N_11862,N_6030,N_6397);
and U11863 (N_11863,N_6728,N_8596);
nor U11864 (N_11864,N_7142,N_6622);
nor U11865 (N_11865,N_7859,N_8172);
nand U11866 (N_11866,N_8961,N_6349);
or U11867 (N_11867,N_8845,N_8272);
nor U11868 (N_11868,N_8432,N_8109);
and U11869 (N_11869,N_6523,N_6818);
or U11870 (N_11870,N_6978,N_6577);
or U11871 (N_11871,N_7905,N_8890);
or U11872 (N_11872,N_7043,N_7825);
nand U11873 (N_11873,N_6837,N_6887);
nor U11874 (N_11874,N_7269,N_7744);
and U11875 (N_11875,N_8448,N_8285);
nor U11876 (N_11876,N_7502,N_7674);
or U11877 (N_11877,N_8204,N_7974);
nor U11878 (N_11878,N_7751,N_8012);
nor U11879 (N_11879,N_7932,N_7158);
or U11880 (N_11880,N_6550,N_6068);
and U11881 (N_11881,N_7865,N_8134);
or U11882 (N_11882,N_8208,N_6464);
nand U11883 (N_11883,N_7215,N_7187);
nand U11884 (N_11884,N_6965,N_6754);
nand U11885 (N_11885,N_6313,N_8520);
nand U11886 (N_11886,N_7204,N_7537);
and U11887 (N_11887,N_8777,N_7790);
nor U11888 (N_11888,N_7669,N_8557);
nand U11889 (N_11889,N_7845,N_8824);
nor U11890 (N_11890,N_7470,N_6571);
nand U11891 (N_11891,N_6638,N_7224);
or U11892 (N_11892,N_7081,N_8735);
or U11893 (N_11893,N_7453,N_8057);
or U11894 (N_11894,N_6205,N_7217);
nand U11895 (N_11895,N_8608,N_8241);
or U11896 (N_11896,N_6821,N_7279);
nand U11897 (N_11897,N_8250,N_7446);
and U11898 (N_11898,N_8672,N_8613);
nor U11899 (N_11899,N_6626,N_6654);
nor U11900 (N_11900,N_6780,N_8905);
nor U11901 (N_11901,N_7625,N_7330);
and U11902 (N_11902,N_8159,N_7239);
or U11903 (N_11903,N_6643,N_6566);
or U11904 (N_11904,N_6445,N_8716);
and U11905 (N_11905,N_6785,N_7967);
nor U11906 (N_11906,N_6003,N_8262);
and U11907 (N_11907,N_6269,N_7515);
nor U11908 (N_11908,N_8939,N_8593);
or U11909 (N_11909,N_6510,N_8089);
nand U11910 (N_11910,N_6209,N_7860);
nor U11911 (N_11911,N_6720,N_6472);
and U11912 (N_11912,N_6536,N_6928);
or U11913 (N_11913,N_6698,N_8248);
or U11914 (N_11914,N_7670,N_7557);
nor U11915 (N_11915,N_7580,N_7420);
or U11916 (N_11916,N_8067,N_7676);
or U11917 (N_11917,N_7131,N_8160);
nand U11918 (N_11918,N_6281,N_8394);
and U11919 (N_11919,N_8497,N_6291);
nand U11920 (N_11920,N_8617,N_6317);
or U11921 (N_11921,N_8900,N_8859);
and U11922 (N_11922,N_7260,N_8904);
and U11923 (N_11923,N_8324,N_8290);
nor U11924 (N_11924,N_7286,N_8106);
or U11925 (N_11925,N_7213,N_8633);
nor U11926 (N_11926,N_8674,N_8801);
or U11927 (N_11927,N_6583,N_7356);
nor U11928 (N_11928,N_7113,N_8882);
and U11929 (N_11929,N_8609,N_7484);
nor U11930 (N_11930,N_8293,N_7232);
nor U11931 (N_11931,N_7528,N_7196);
or U11932 (N_11932,N_8352,N_6437);
nor U11933 (N_11933,N_8138,N_8413);
xnor U11934 (N_11934,N_8626,N_7015);
or U11935 (N_11935,N_6982,N_7867);
or U11936 (N_11936,N_6004,N_7304);
or U11937 (N_11937,N_8856,N_6659);
nor U11938 (N_11938,N_8554,N_8532);
xor U11939 (N_11939,N_6382,N_6781);
and U11940 (N_11940,N_6190,N_6214);
nand U11941 (N_11941,N_7120,N_7623);
and U11942 (N_11942,N_7014,N_7121);
and U11943 (N_11943,N_7177,N_8491);
nor U11944 (N_11944,N_7361,N_6385);
or U11945 (N_11945,N_8533,N_6277);
nand U11946 (N_11946,N_7945,N_8509);
nand U11947 (N_11947,N_7020,N_6779);
nor U11948 (N_11948,N_8267,N_8254);
nand U11949 (N_11949,N_8562,N_8982);
or U11950 (N_11950,N_6659,N_8299);
nand U11951 (N_11951,N_7615,N_8883);
or U11952 (N_11952,N_8237,N_7669);
nand U11953 (N_11953,N_8793,N_8163);
or U11954 (N_11954,N_7535,N_8349);
or U11955 (N_11955,N_7888,N_8066);
nor U11956 (N_11956,N_6395,N_6049);
and U11957 (N_11957,N_8946,N_8377);
and U11958 (N_11958,N_8501,N_6028);
nor U11959 (N_11959,N_6367,N_7466);
nand U11960 (N_11960,N_7882,N_7612);
and U11961 (N_11961,N_8260,N_8825);
nor U11962 (N_11962,N_6490,N_8186);
nand U11963 (N_11963,N_6919,N_7787);
nand U11964 (N_11964,N_6012,N_7825);
and U11965 (N_11965,N_6416,N_6616);
xnor U11966 (N_11966,N_6717,N_8005);
nand U11967 (N_11967,N_8355,N_8412);
nand U11968 (N_11968,N_8640,N_8321);
or U11969 (N_11969,N_7464,N_8831);
nor U11970 (N_11970,N_6992,N_6014);
and U11971 (N_11971,N_8376,N_8637);
nor U11972 (N_11972,N_7276,N_8428);
or U11973 (N_11973,N_8438,N_7087);
or U11974 (N_11974,N_8022,N_6245);
and U11975 (N_11975,N_7647,N_8228);
or U11976 (N_11976,N_6296,N_6407);
or U11977 (N_11977,N_6632,N_8804);
nor U11978 (N_11978,N_6595,N_6828);
and U11979 (N_11979,N_7452,N_6574);
nand U11980 (N_11980,N_7481,N_8555);
nand U11981 (N_11981,N_7503,N_8154);
and U11982 (N_11982,N_7779,N_6961);
and U11983 (N_11983,N_8859,N_8366);
or U11984 (N_11984,N_8545,N_6717);
or U11985 (N_11985,N_8108,N_7167);
and U11986 (N_11986,N_6862,N_7606);
or U11987 (N_11987,N_7282,N_8012);
and U11988 (N_11988,N_6226,N_7157);
nor U11989 (N_11989,N_8319,N_7892);
nand U11990 (N_11990,N_8989,N_6275);
nor U11991 (N_11991,N_6373,N_6218);
or U11992 (N_11992,N_7582,N_7682);
or U11993 (N_11993,N_8809,N_6064);
and U11994 (N_11994,N_8567,N_8593);
nand U11995 (N_11995,N_7492,N_6753);
or U11996 (N_11996,N_6049,N_6452);
nand U11997 (N_11997,N_7841,N_6624);
and U11998 (N_11998,N_6786,N_7521);
nand U11999 (N_11999,N_8700,N_6095);
nand U12000 (N_12000,N_9910,N_11996);
nor U12001 (N_12001,N_9971,N_10147);
nor U12002 (N_12002,N_11323,N_10717);
nor U12003 (N_12003,N_10188,N_10863);
nor U12004 (N_12004,N_10042,N_11967);
or U12005 (N_12005,N_11050,N_9493);
and U12006 (N_12006,N_10230,N_9585);
nand U12007 (N_12007,N_10872,N_11742);
nor U12008 (N_12008,N_11704,N_11374);
and U12009 (N_12009,N_11043,N_11919);
and U12010 (N_12010,N_11526,N_11238);
nand U12011 (N_12011,N_11133,N_11095);
or U12012 (N_12012,N_11462,N_11661);
nand U12013 (N_12013,N_11191,N_11453);
nor U12014 (N_12014,N_10319,N_11950);
nand U12015 (N_12015,N_9334,N_9641);
and U12016 (N_12016,N_9582,N_11606);
and U12017 (N_12017,N_11454,N_10472);
and U12018 (N_12018,N_10272,N_11074);
nor U12019 (N_12019,N_10043,N_9777);
nand U12020 (N_12020,N_9982,N_10412);
nor U12021 (N_12021,N_10489,N_10049);
nor U12022 (N_12022,N_11787,N_9681);
nand U12023 (N_12023,N_10249,N_11507);
nand U12024 (N_12024,N_10628,N_10607);
nor U12025 (N_12025,N_9770,N_9924);
and U12026 (N_12026,N_11944,N_10587);
or U12027 (N_12027,N_9616,N_10906);
nand U12028 (N_12028,N_10307,N_11219);
nand U12029 (N_12029,N_9675,N_11156);
and U12030 (N_12030,N_10434,N_11502);
and U12031 (N_12031,N_9541,N_9726);
or U12032 (N_12032,N_9066,N_11817);
and U12033 (N_12033,N_9399,N_10217);
nor U12034 (N_12034,N_9504,N_9759);
or U12035 (N_12035,N_9513,N_11332);
nand U12036 (N_12036,N_10975,N_11296);
nor U12037 (N_12037,N_11913,N_10842);
nor U12038 (N_12038,N_11062,N_10321);
or U12039 (N_12039,N_9783,N_10942);
nor U12040 (N_12040,N_11932,N_11153);
and U12041 (N_12041,N_11623,N_10559);
and U12042 (N_12042,N_10294,N_11487);
and U12043 (N_12043,N_9596,N_10564);
nor U12044 (N_12044,N_10347,N_9124);
and U12045 (N_12045,N_9395,N_9037);
and U12046 (N_12046,N_10600,N_10422);
nand U12047 (N_12047,N_9220,N_10457);
nor U12048 (N_12048,N_10391,N_10828);
and U12049 (N_12049,N_11549,N_10405);
nand U12050 (N_12050,N_9986,N_9444);
or U12051 (N_12051,N_9791,N_10380);
nand U12052 (N_12052,N_9741,N_10162);
or U12053 (N_12053,N_11670,N_10428);
and U12054 (N_12054,N_10464,N_9572);
and U12055 (N_12055,N_9191,N_9902);
nand U12056 (N_12056,N_9202,N_9677);
and U12057 (N_12057,N_10550,N_9417);
and U12058 (N_12058,N_11885,N_10511);
and U12059 (N_12059,N_10327,N_10661);
nor U12060 (N_12060,N_9315,N_10030);
nand U12061 (N_12061,N_11873,N_9861);
or U12062 (N_12062,N_10664,N_11566);
and U12063 (N_12063,N_10078,N_9915);
and U12064 (N_12064,N_10096,N_10088);
nand U12065 (N_12065,N_9438,N_10917);
nor U12066 (N_12066,N_10022,N_11647);
nand U12067 (N_12067,N_11884,N_9656);
nor U12068 (N_12068,N_9031,N_11038);
nand U12069 (N_12069,N_11975,N_9969);
nor U12070 (N_12070,N_10337,N_9146);
or U12071 (N_12071,N_11535,N_11791);
or U12072 (N_12072,N_10393,N_11151);
nand U12073 (N_12073,N_11018,N_11053);
and U12074 (N_12074,N_11115,N_11337);
and U12075 (N_12075,N_10077,N_10884);
nor U12076 (N_12076,N_10366,N_9743);
and U12077 (N_12077,N_9440,N_9758);
nor U12078 (N_12078,N_10614,N_10224);
nor U12079 (N_12079,N_11049,N_9344);
or U12080 (N_12080,N_9203,N_11278);
and U12081 (N_12081,N_10996,N_9631);
and U12082 (N_12082,N_10617,N_10362);
nor U12083 (N_12083,N_9524,N_10844);
nor U12084 (N_12084,N_10971,N_11784);
and U12085 (N_12085,N_9486,N_10107);
or U12086 (N_12086,N_10885,N_10952);
or U12087 (N_12087,N_9548,N_11363);
or U12088 (N_12088,N_9101,N_11294);
nand U12089 (N_12089,N_11421,N_9721);
nor U12090 (N_12090,N_10868,N_11710);
nor U12091 (N_12091,N_11551,N_10845);
nand U12092 (N_12092,N_10447,N_11200);
nand U12093 (N_12093,N_11856,N_11665);
nor U12094 (N_12094,N_11673,N_11061);
nor U12095 (N_12095,N_11226,N_10915);
and U12096 (N_12096,N_10331,N_9539);
and U12097 (N_12097,N_9680,N_9970);
or U12098 (N_12098,N_10252,N_9615);
or U12099 (N_12099,N_11359,N_10704);
or U12100 (N_12100,N_9566,N_10069);
nand U12101 (N_12101,N_10601,N_11953);
and U12102 (N_12102,N_10718,N_11654);
nand U12103 (N_12103,N_11700,N_10445);
or U12104 (N_12104,N_9893,N_9457);
or U12105 (N_12105,N_9560,N_9150);
nand U12106 (N_12106,N_9697,N_9727);
or U12107 (N_12107,N_11940,N_9254);
or U12108 (N_12108,N_9612,N_10357);
nor U12109 (N_12109,N_11703,N_9333);
and U12110 (N_12110,N_9209,N_9782);
and U12111 (N_12111,N_11290,N_9657);
nand U12112 (N_12112,N_10411,N_10988);
or U12113 (N_12113,N_11045,N_10560);
nand U12114 (N_12114,N_11047,N_10072);
and U12115 (N_12115,N_10935,N_9421);
nand U12116 (N_12116,N_10314,N_9495);
nor U12117 (N_12117,N_10303,N_11065);
or U12118 (N_12118,N_11772,N_11746);
nand U12119 (N_12119,N_10288,N_9478);
and U12120 (N_12120,N_9581,N_11974);
and U12121 (N_12121,N_11773,N_9323);
or U12122 (N_12122,N_9480,N_11761);
or U12123 (N_12123,N_9933,N_10467);
nand U12124 (N_12124,N_10295,N_10378);
or U12125 (N_12125,N_10806,N_11271);
nor U12126 (N_12126,N_9255,N_11792);
or U12127 (N_12127,N_9637,N_11508);
nand U12128 (N_12128,N_11128,N_9604);
or U12129 (N_12129,N_10974,N_11447);
nor U12130 (N_12130,N_9038,N_11331);
nand U12131 (N_12131,N_10106,N_11517);
and U12132 (N_12132,N_9174,N_10274);
and U12133 (N_12133,N_9055,N_10115);
and U12134 (N_12134,N_11215,N_11938);
or U12135 (N_12135,N_11531,N_11829);
nor U12136 (N_12136,N_9165,N_11064);
nand U12137 (N_12137,N_11099,N_9356);
nor U12138 (N_12138,N_9898,N_9733);
and U12139 (N_12139,N_10883,N_9739);
or U12140 (N_12140,N_9089,N_11450);
or U12141 (N_12141,N_10984,N_11329);
nor U12142 (N_12142,N_9502,N_11336);
nand U12143 (N_12143,N_10210,N_11106);
or U12144 (N_12144,N_10625,N_9114);
nor U12145 (N_12145,N_11528,N_10758);
nand U12146 (N_12146,N_9967,N_9947);
or U12147 (N_12147,N_11154,N_11883);
nand U12148 (N_12148,N_11930,N_10655);
and U12149 (N_12149,N_9723,N_9303);
and U12150 (N_12150,N_11912,N_9455);
or U12151 (N_12151,N_10871,N_11165);
nor U12152 (N_12152,N_9251,N_9109);
or U12153 (N_12153,N_9278,N_9400);
and U12154 (N_12154,N_10719,N_11457);
or U12155 (N_12155,N_11619,N_9128);
and U12156 (N_12156,N_10207,N_9229);
nand U12157 (N_12157,N_9588,N_11512);
and U12158 (N_12158,N_9434,N_9242);
nor U12159 (N_12159,N_10399,N_9980);
nand U12160 (N_12160,N_10205,N_10978);
and U12161 (N_12161,N_10619,N_9270);
nand U12162 (N_12162,N_9266,N_9143);
nor U12163 (N_12163,N_11832,N_10199);
or U12164 (N_12164,N_11183,N_9184);
or U12165 (N_12165,N_11922,N_11197);
nor U12166 (N_12166,N_11845,N_10375);
or U12167 (N_12167,N_9005,N_10181);
and U12168 (N_12168,N_11306,N_10371);
nand U12169 (N_12169,N_11970,N_11721);
or U12170 (N_12170,N_9979,N_11889);
nor U12171 (N_12171,N_10090,N_9145);
and U12172 (N_12172,N_11185,N_10134);
nand U12173 (N_12173,N_10169,N_9082);
or U12174 (N_12174,N_10540,N_10258);
nor U12175 (N_12175,N_9877,N_9887);
nor U12176 (N_12176,N_11625,N_10418);
nand U12177 (N_12177,N_10754,N_9019);
or U12178 (N_12178,N_11287,N_9832);
or U12179 (N_12179,N_11840,N_11574);
nand U12180 (N_12180,N_9685,N_10116);
nor U12181 (N_12181,N_10015,N_11385);
nor U12182 (N_12182,N_11167,N_11173);
nand U12183 (N_12183,N_11389,N_11699);
and U12184 (N_12184,N_9911,N_11486);
nor U12185 (N_12185,N_11663,N_11866);
nand U12186 (N_12186,N_10150,N_9067);
and U12187 (N_12187,N_9827,N_10306);
and U12188 (N_12188,N_11893,N_11790);
nor U12189 (N_12189,N_10913,N_9406);
or U12190 (N_12190,N_11190,N_10908);
nand U12191 (N_12191,N_11342,N_11155);
nand U12192 (N_12192,N_9773,N_11322);
or U12193 (N_12193,N_9611,N_11078);
and U12194 (N_12194,N_10992,N_11992);
nor U12195 (N_12195,N_10712,N_11776);
nand U12196 (N_12196,N_10632,N_11240);
nor U12197 (N_12197,N_10603,N_11069);
and U12198 (N_12198,N_10241,N_11552);
nand U12199 (N_12199,N_9941,N_11785);
nor U12200 (N_12200,N_10735,N_9992);
nor U12201 (N_12201,N_10960,N_10963);
nand U12202 (N_12202,N_9000,N_10002);
nand U12203 (N_12203,N_11004,N_11333);
nor U12204 (N_12204,N_11616,N_9245);
and U12205 (N_12205,N_10178,N_11231);
and U12206 (N_12206,N_11463,N_9022);
nand U12207 (N_12207,N_9413,N_11474);
nor U12208 (N_12208,N_9643,N_11230);
and U12209 (N_12209,N_9899,N_10175);
or U12210 (N_12210,N_10056,N_11514);
or U12211 (N_12211,N_11591,N_9466);
and U12212 (N_12212,N_10648,N_9219);
nor U12213 (N_12213,N_10736,N_9144);
and U12214 (N_12214,N_9593,N_10584);
nand U12215 (N_12215,N_11113,N_10263);
nor U12216 (N_12216,N_11779,N_11426);
nor U12217 (N_12217,N_11117,N_10204);
nor U12218 (N_12218,N_9852,N_9071);
nor U12219 (N_12219,N_9286,N_9594);
nand U12220 (N_12220,N_11534,N_9807);
nor U12221 (N_12221,N_9408,N_11533);
or U12222 (N_12222,N_9218,N_10865);
xor U12223 (N_12223,N_10866,N_10710);
or U12224 (N_12224,N_9802,N_9574);
and U12225 (N_12225,N_10360,N_11142);
and U12226 (N_12226,N_9891,N_9573);
nor U12227 (N_12227,N_11926,N_11221);
nor U12228 (N_12228,N_10186,N_10976);
and U12229 (N_12229,N_10983,N_11989);
nand U12230 (N_12230,N_9989,N_11725);
and U12231 (N_12231,N_9954,N_10171);
nand U12232 (N_12232,N_11478,N_10642);
or U12233 (N_12233,N_9557,N_9017);
nand U12234 (N_12234,N_11499,N_11291);
nor U12235 (N_12235,N_11554,N_11434);
nand U12236 (N_12236,N_11163,N_11650);
nand U12237 (N_12237,N_9694,N_10521);
or U12238 (N_12238,N_10462,N_11695);
nor U12239 (N_12239,N_11983,N_11403);
and U12240 (N_12240,N_11448,N_10959);
and U12241 (N_12241,N_10951,N_9234);
or U12242 (N_12242,N_9569,N_11316);
and U12243 (N_12243,N_11545,N_9401);
nand U12244 (N_12244,N_11923,N_10697);
and U12245 (N_12245,N_10262,N_9301);
nor U12246 (N_12246,N_11058,N_10849);
or U12247 (N_12247,N_11079,N_9647);
nand U12248 (N_12248,N_11734,N_10568);
and U12249 (N_12249,N_10683,N_11916);
and U12250 (N_12250,N_11402,N_9096);
nor U12251 (N_12251,N_9650,N_10752);
or U12252 (N_12252,N_11862,N_9760);
or U12253 (N_12253,N_10195,N_11419);
nand U12254 (N_12254,N_10456,N_10739);
nor U12255 (N_12255,N_9993,N_9195);
nand U12256 (N_12256,N_9385,N_11380);
or U12257 (N_12257,N_9994,N_9884);
and U12258 (N_12258,N_11174,N_9774);
nand U12259 (N_12259,N_9142,N_11556);
and U12260 (N_12260,N_9917,N_10962);
and U12261 (N_12261,N_9431,N_11601);
and U12262 (N_12262,N_10918,N_11494);
nor U12263 (N_12263,N_11266,N_11994);
and U12264 (N_12264,N_10370,N_9630);
nand U12265 (N_12265,N_9320,N_9181);
nand U12266 (N_12266,N_11460,N_9439);
and U12267 (N_12267,N_10082,N_9757);
nand U12268 (N_12268,N_9873,N_10479);
nand U12269 (N_12269,N_9169,N_9649);
or U12270 (N_12270,N_11971,N_9415);
nand U12271 (N_12271,N_11990,N_10046);
or U12272 (N_12272,N_9208,N_10440);
and U12273 (N_12273,N_11760,N_11091);
nor U12274 (N_12274,N_11080,N_9805);
or U12275 (N_12275,N_9343,N_11366);
nor U12276 (N_12276,N_11475,N_9359);
or U12277 (N_12277,N_10458,N_9667);
nor U12278 (N_12278,N_9492,N_11059);
or U12279 (N_12279,N_11878,N_9968);
and U12280 (N_12280,N_10157,N_9349);
and U12281 (N_12281,N_9603,N_11850);
nand U12282 (N_12282,N_11222,N_11087);
nand U12283 (N_12283,N_10964,N_11060);
and U12284 (N_12284,N_10334,N_11777);
or U12285 (N_12285,N_9227,N_9821);
nand U12286 (N_12286,N_11339,N_11918);
nor U12287 (N_12287,N_9118,N_9583);
nand U12288 (N_12288,N_9332,N_9942);
and U12289 (N_12289,N_9407,N_9776);
or U12290 (N_12290,N_11892,N_10510);
nand U12291 (N_12291,N_11657,N_9151);
nand U12292 (N_12292,N_11749,N_11073);
and U12293 (N_12293,N_9272,N_10981);
and U12294 (N_12294,N_9370,N_10410);
nor U12295 (N_12295,N_11481,N_9238);
nor U12296 (N_12296,N_9053,N_10494);
or U12297 (N_12297,N_10499,N_9060);
or U12298 (N_12298,N_9830,N_11655);
nand U12299 (N_12299,N_11881,N_10894);
nand U12300 (N_12300,N_11691,N_10417);
nor U12301 (N_12301,N_9163,N_9012);
nor U12302 (N_12302,N_10796,N_9461);
and U12303 (N_12303,N_9295,N_11801);
or U12304 (N_12304,N_9479,N_11604);
nor U12305 (N_12305,N_11543,N_11648);
and U12306 (N_12306,N_11598,N_9023);
nand U12307 (N_12307,N_9606,N_11867);
nor U12308 (N_12308,N_9404,N_9375);
and U12309 (N_12309,N_10566,N_11658);
and U12310 (N_12310,N_11755,N_9010);
and U12311 (N_12311,N_10497,N_9059);
nor U12312 (N_12312,N_10737,N_11660);
nor U12313 (N_12313,N_9462,N_9753);
nor U12314 (N_12314,N_10825,N_10565);
nand U12315 (N_12315,N_10563,N_11954);
nor U12316 (N_12316,N_11175,N_11455);
nor U12317 (N_12317,N_10359,N_11269);
nand U12318 (N_12318,N_10986,N_9808);
or U12319 (N_12319,N_9500,N_9056);
or U12320 (N_12320,N_11887,N_11805);
xnor U12321 (N_12321,N_11644,N_9983);
or U12322 (N_12322,N_10649,N_10136);
or U12323 (N_12323,N_10747,N_11877);
or U12324 (N_12324,N_9691,N_11548);
nor U12325 (N_12325,N_9900,N_9475);
or U12326 (N_12326,N_11247,N_10933);
and U12327 (N_12327,N_9926,N_11067);
nand U12328 (N_12328,N_10676,N_10782);
or U12329 (N_12329,N_11224,N_10197);
or U12330 (N_12330,N_9886,N_9883);
and U12331 (N_12331,N_11284,N_10376);
and U12332 (N_12332,N_10524,N_9182);
nor U12333 (N_12333,N_9347,N_10439);
or U12334 (N_12334,N_9903,N_9083);
or U12335 (N_12335,N_9390,N_10823);
nand U12336 (N_12336,N_11754,N_10356);
nand U12337 (N_12337,N_11645,N_11869);
and U12338 (N_12338,N_11007,N_11468);
or U12339 (N_12339,N_9014,N_9798);
nor U12340 (N_12340,N_10048,N_9384);
nor U12341 (N_12341,N_9291,N_9073);
or U12342 (N_12342,N_9951,N_11304);
nand U12343 (N_12343,N_10878,N_10010);
nor U12344 (N_12344,N_10170,N_11594);
and U12345 (N_12345,N_11443,N_9609);
nor U12346 (N_12346,N_9396,N_9939);
nor U12347 (N_12347,N_9171,N_9365);
and U12348 (N_12348,N_11125,N_11308);
nor U12349 (N_12349,N_9925,N_11281);
and U12350 (N_12350,N_10490,N_11236);
and U12351 (N_12351,N_10816,N_10164);
nand U12352 (N_12352,N_9977,N_9510);
nand U12353 (N_12353,N_10688,N_9722);
and U12354 (N_12354,N_11620,N_9695);
nor U12355 (N_12355,N_10117,N_11608);
nor U12356 (N_12356,N_9020,N_9080);
and U12357 (N_12357,N_9872,N_10932);
or U12358 (N_12358,N_10220,N_10998);
nor U12359 (N_12359,N_9578,N_9806);
nand U12360 (N_12360,N_11192,N_9125);
or U12361 (N_12361,N_9004,N_10335);
nand U12362 (N_12362,N_9355,N_9904);
and U12363 (N_12363,N_9689,N_10629);
nor U12364 (N_12364,N_10593,N_10223);
and U12365 (N_12365,N_10153,N_9134);
nor U12366 (N_12366,N_9389,N_10338);
nor U12367 (N_12367,N_10189,N_10451);
nor U12368 (N_12368,N_10012,N_10093);
nand U12369 (N_12369,N_9644,N_10592);
nand U12370 (N_12370,N_9546,N_9654);
nor U12371 (N_12371,N_11157,N_10322);
nor U12372 (N_12372,N_10921,N_9374);
xnor U12373 (N_12373,N_10315,N_11243);
nand U12374 (N_12374,N_9187,N_11521);
or U12375 (N_12375,N_10547,N_10343);
and U12376 (N_12376,N_10260,N_10937);
or U12377 (N_12377,N_11086,N_10953);
and U12378 (N_12378,N_9833,N_9442);
nand U12379 (N_12379,N_9011,N_10123);
or U12380 (N_12380,N_11748,N_11998);
nand U12381 (N_12381,N_10855,N_9686);
nand U12382 (N_12382,N_11980,N_10973);
and U12383 (N_12383,N_11076,N_9354);
xor U12384 (N_12384,N_9232,N_9558);
or U12385 (N_12385,N_9523,N_9257);
nor U12386 (N_12386,N_10000,N_11147);
and U12387 (N_12387,N_10398,N_9090);
nand U12388 (N_12388,N_11097,N_9838);
nand U12389 (N_12389,N_9794,N_10749);
nor U12390 (N_12390,N_9450,N_11234);
and U12391 (N_12391,N_10192,N_9411);
or U12392 (N_12392,N_10812,N_9831);
nor U12393 (N_12393,N_11977,N_9561);
and U12394 (N_12394,N_11516,N_10846);
nand U12395 (N_12395,N_10856,N_9820);
nor U12396 (N_12396,N_11570,N_9953);
nor U12397 (N_12397,N_9050,N_11627);
nor U12398 (N_12398,N_9247,N_9263);
or U12399 (N_12399,N_11622,N_9788);
and U12400 (N_12400,N_10530,N_10858);
nand U12401 (N_12401,N_11618,N_9525);
nand U12402 (N_12402,N_11041,N_11706);
nor U12403 (N_12403,N_11571,N_9908);
nor U12404 (N_12404,N_11202,N_10805);
nor U12405 (N_12405,N_11522,N_9966);
and U12406 (N_12406,N_10250,N_11781);
and U12407 (N_12407,N_10874,N_9714);
xor U12408 (N_12408,N_10837,N_10145);
xnor U12409 (N_12409,N_11327,N_9366);
or U12410 (N_12410,N_10527,N_9129);
and U12411 (N_12411,N_10124,N_10811);
and U12412 (N_12412,N_9912,N_10453);
nor U12413 (N_12413,N_10892,N_9030);
nor U12414 (N_12414,N_11498,N_10528);
nor U12415 (N_12415,N_11206,N_11044);
or U12416 (N_12416,N_11144,N_11324);
nor U12417 (N_12417,N_9405,N_10695);
and U12418 (N_12418,N_11567,N_11633);
nor U12419 (N_12419,N_9664,N_11250);
nand U12420 (N_12420,N_9472,N_11199);
nand U12421 (N_12421,N_10897,N_10087);
and U12422 (N_12422,N_10243,N_10038);
nand U12423 (N_12423,N_9666,N_11635);
and U12424 (N_12424,N_10196,N_11229);
or U12425 (N_12425,N_10656,N_9081);
nor U12426 (N_12426,N_11799,N_11634);
and U12427 (N_12427,N_10626,N_11435);
or U12428 (N_12428,N_10122,N_9063);
or U12429 (N_12429,N_10214,N_9288);
or U12430 (N_12430,N_9447,N_9771);
nor U12431 (N_12431,N_11529,N_11480);
nand U12432 (N_12432,N_9568,N_11582);
nor U12433 (N_12433,N_11607,N_9882);
nor U12434 (N_12434,N_11260,N_11015);
nand U12435 (N_12435,N_9709,N_9509);
nand U12436 (N_12436,N_10966,N_10045);
and U12437 (N_12437,N_11251,N_10995);
nand U12438 (N_12438,N_9981,N_10008);
nand U12439 (N_12439,N_9522,N_11943);
and U12440 (N_12440,N_9460,N_11798);
nand U12441 (N_12441,N_10353,N_9635);
nand U12442 (N_12442,N_9551,N_10029);
and U12443 (N_12443,N_9819,N_11212);
or U12444 (N_12444,N_9314,N_9331);
or U12445 (N_12445,N_10910,N_10280);
and U12446 (N_12446,N_10218,N_9372);
nand U12447 (N_12447,N_11265,N_9671);
and U12448 (N_12448,N_9698,N_10242);
nand U12449 (N_12449,N_10244,N_9533);
and U12450 (N_12450,N_9829,N_10947);
and U12451 (N_12451,N_11979,N_10616);
and U12452 (N_12452,N_10923,N_9784);
or U12453 (N_12453,N_10179,N_9536);
nor U12454 (N_12454,N_9264,N_9136);
nor U12455 (N_12455,N_9088,N_9490);
or U12456 (N_12456,N_10316,N_10832);
or U12457 (N_12457,N_10860,N_10427);
nand U12458 (N_12458,N_11613,N_11629);
and U12459 (N_12459,N_10114,N_10604);
or U12460 (N_12460,N_9324,N_10429);
nor U12461 (N_12461,N_11292,N_9707);
or U12462 (N_12462,N_9274,N_9589);
nand U12463 (N_12463,N_10687,N_11149);
or U12464 (N_12464,N_11587,N_10830);
nor U12465 (N_12465,N_10501,N_10231);
or U12466 (N_12466,N_9617,N_9237);
nor U12467 (N_12467,N_9342,N_9985);
nand U12468 (N_12468,N_10443,N_10141);
nor U12469 (N_12469,N_9197,N_11684);
nand U12470 (N_12470,N_11577,N_11417);
nand U12471 (N_12471,N_10623,N_10113);
and U12472 (N_12472,N_10425,N_10054);
nand U12473 (N_12473,N_10095,N_10351);
nor U12474 (N_12474,N_11640,N_10597);
nand U12475 (N_12475,N_10377,N_10586);
or U12476 (N_12476,N_9840,N_10914);
nor U12477 (N_12477,N_11656,N_9132);
and U12478 (N_12478,N_9795,N_10817);
nand U12479 (N_12479,N_11299,N_10075);
or U12480 (N_12480,N_9640,N_9294);
and U12481 (N_12481,N_9549,N_11028);
nor U12482 (N_12482,N_10624,N_11112);
or U12483 (N_12483,N_10146,N_11579);
nor U12484 (N_12484,N_9244,N_9960);
and U12485 (N_12485,N_10140,N_10571);
nor U12486 (N_12486,N_11035,N_9043);
nor U12487 (N_12487,N_9039,N_9418);
and U12488 (N_12488,N_9319,N_9468);
or U12489 (N_12489,N_11709,N_11063);
and U12490 (N_12490,N_9634,N_10081);
nand U12491 (N_12491,N_11909,N_10588);
and U12492 (N_12492,N_11711,N_9717);
or U12493 (N_12493,N_11836,N_10763);
or U12494 (N_12494,N_11248,N_11961);
or U12495 (N_12495,N_11575,N_9179);
or U12496 (N_12496,N_10156,N_10738);
or U12497 (N_12497,N_11318,N_11871);
nor U12498 (N_12498,N_11811,N_11201);
nand U12499 (N_12499,N_9972,N_9668);
nor U12500 (N_12500,N_10302,N_9537);
and U12501 (N_12501,N_9962,N_11542);
or U12502 (N_12502,N_9608,N_9765);
and U12503 (N_12503,N_10459,N_11172);
nor U12504 (N_12504,N_9087,N_10714);
and U12505 (N_12505,N_9684,N_11581);
nor U12506 (N_12506,N_10163,N_10483);
or U12507 (N_12507,N_9859,N_11904);
nor U12508 (N_12508,N_9046,N_11213);
nor U12509 (N_12509,N_10066,N_10006);
nor U12510 (N_12510,N_10235,N_10415);
nand U12511 (N_12511,N_9141,N_10783);
or U12512 (N_12512,N_9007,N_11437);
or U12513 (N_12513,N_9521,N_11241);
nor U12514 (N_12514,N_10076,N_11991);
nor U12515 (N_12515,N_9044,N_9422);
nand U12516 (N_12516,N_9896,N_10167);
or U12517 (N_12517,N_10047,N_11268);
nor U12518 (N_12518,N_9489,N_11841);
and U12519 (N_12519,N_11712,N_11479);
nor U12520 (N_12520,N_9213,N_9944);
and U12521 (N_12521,N_11894,N_10397);
or U12522 (N_12522,N_10441,N_10151);
nor U12523 (N_12523,N_11143,N_9281);
and U12524 (N_12524,N_9946,N_11838);
and U12525 (N_12525,N_9275,N_10080);
and U12526 (N_12526,N_11789,N_11048);
nand U12527 (N_12527,N_9397,N_9731);
and U12528 (N_12528,N_9474,N_9736);
and U12529 (N_12529,N_9430,N_9297);
or U12530 (N_12530,N_10034,N_9813);
and U12531 (N_12531,N_9720,N_10662);
or U12532 (N_12532,N_11539,N_9346);
nor U12533 (N_12533,N_9547,N_10663);
and U12534 (N_12534,N_9761,N_9380);
or U12535 (N_12535,N_9287,N_10916);
and U12536 (N_12536,N_10793,N_11678);
and U12537 (N_12537,N_11679,N_10305);
nand U12538 (N_12538,N_11524,N_10552);
nor U12539 (N_12539,N_11546,N_10298);
nand U12540 (N_12540,N_10641,N_10254);
nor U12541 (N_12541,N_10814,N_11993);
and U12542 (N_12542,N_9398,N_10730);
nand U12543 (N_12543,N_11906,N_10009);
or U12544 (N_12544,N_9619,N_11947);
nand U12545 (N_12545,N_9351,N_10361);
and U12546 (N_12546,N_10620,N_10948);
nor U12547 (N_12547,N_9373,N_9869);
nor U12548 (N_12548,N_9498,N_9660);
and U12549 (N_12549,N_10092,N_11626);
or U12550 (N_12550,N_10039,N_10446);
and U12551 (N_12551,N_9337,N_9094);
and U12552 (N_12552,N_9168,N_11510);
or U12553 (N_12553,N_11134,N_11057);
nor U12554 (N_12554,N_10901,N_10198);
or U12555 (N_12555,N_11227,N_10621);
nand U12556 (N_12556,N_11104,N_10373);
or U12557 (N_12557,N_11936,N_10779);
nor U12558 (N_12558,N_11491,N_10007);
and U12559 (N_12559,N_11010,N_9527);
nand U12560 (N_12560,N_11261,N_10344);
nor U12561 (N_12561,N_11075,N_9290);
nand U12562 (N_12562,N_9133,N_9867);
or U12563 (N_12563,N_9716,N_10919);
nor U12564 (N_12564,N_9035,N_10653);
and U12565 (N_12565,N_9496,N_11753);
nor U12566 (N_12566,N_10561,N_11505);
nor U12567 (N_12567,N_10651,N_10631);
nor U12568 (N_12568,N_10310,N_11423);
or U12569 (N_12569,N_11714,N_10019);
or U12570 (N_12570,N_10493,N_10339);
nor U12571 (N_12571,N_10455,N_11483);
nand U12572 (N_12572,N_11664,N_9228);
or U12573 (N_12573,N_11051,N_9543);
or U12574 (N_12574,N_11334,N_9692);
or U12575 (N_12575,N_9190,N_10707);
nor U12576 (N_12576,N_11189,N_11459);
and U12577 (N_12577,N_10486,N_9535);
nor U12578 (N_12578,N_10471,N_9825);
and U12579 (N_12579,N_9064,N_11020);
and U12580 (N_12580,N_11765,N_9880);
nand U12581 (N_12581,N_11055,N_9298);
and U12582 (N_12582,N_11325,N_10221);
nand U12583 (N_12583,N_10102,N_9780);
or U12584 (N_12584,N_9293,N_9084);
nand U12585 (N_12585,N_9026,N_11696);
or U12586 (N_12586,N_10606,N_9183);
and U12587 (N_12587,N_11289,N_9214);
and U12588 (N_12588,N_10599,N_10554);
nand U12589 (N_12589,N_9249,N_10386);
and U12590 (N_12590,N_11252,N_9383);
nor U12591 (N_12591,N_11795,N_9212);
and U12592 (N_12592,N_11409,N_11758);
nand U12593 (N_12593,N_10051,N_10291);
and U12594 (N_12594,N_10927,N_10079);
and U12595 (N_12595,N_11599,N_11258);
nand U12596 (N_12596,N_10672,N_10127);
or U12597 (N_12597,N_10317,N_11818);
and U12598 (N_12598,N_10535,N_11823);
nor U12599 (N_12599,N_11972,N_11180);
and U12600 (N_12600,N_10813,N_10744);
and U12601 (N_12601,N_9273,N_11612);
and U12602 (N_12602,N_11365,N_9850);
nand U12603 (N_12603,N_9764,N_11341);
xor U12604 (N_12604,N_11563,N_11273);
or U12605 (N_12605,N_10278,N_10911);
or U12606 (N_12606,N_9598,N_10345);
nand U12607 (N_12607,N_11039,N_10276);
nand U12608 (N_12608,N_10934,N_10589);
and U12609 (N_12609,N_10505,N_11303);
nand U12610 (N_12610,N_11724,N_9853);
or U12611 (N_12611,N_10067,N_10109);
nand U12612 (N_12612,N_11123,N_9126);
nor U12613 (N_12613,N_10696,N_9008);
and U12614 (N_12614,N_10001,N_9048);
or U12615 (N_12615,N_10728,N_11186);
nand U12616 (N_12616,N_10063,N_10551);
and U12617 (N_12617,N_9162,N_9897);
nand U12618 (N_12618,N_9211,N_10861);
nand U12619 (N_12619,N_11693,N_10745);
nor U12620 (N_12620,N_10301,N_9700);
and U12621 (N_12621,N_11270,N_11911);
and U12622 (N_12622,N_9874,N_9565);
xnor U12623 (N_12623,N_11733,N_10734);
nand U12624 (N_12624,N_10228,N_9927);
nand U12625 (N_12625,N_11782,N_11870);
nand U12626 (N_12626,N_9070,N_11405);
nand U12627 (N_12627,N_10772,N_10602);
and U12628 (N_12628,N_10746,N_9613);
and U12629 (N_12629,N_10675,N_11121);
nor U12630 (N_12630,N_11259,N_10982);
or U12631 (N_12631,N_11401,N_9577);
nand U12632 (N_12632,N_11178,N_10792);
and U12633 (N_12633,N_11429,N_9016);
nand U12634 (N_12634,N_11023,N_11586);
or U12635 (N_12635,N_11858,N_9655);
or U12636 (N_12636,N_10575,N_9458);
and U12637 (N_12637,N_9531,N_9379);
nand U12638 (N_12638,N_9651,N_9312);
and U12639 (N_12639,N_11560,N_9708);
and U12640 (N_12640,N_10529,N_11794);
or U12641 (N_12641,N_9940,N_11518);
nand U12642 (N_12642,N_11921,N_9076);
nor U12643 (N_12643,N_11864,N_11244);
or U12644 (N_12644,N_11756,N_11962);
or U12645 (N_12645,N_9984,N_11707);
nand U12646 (N_12646,N_11948,N_9027);
and U12647 (N_12647,N_10516,N_9514);
nand U12648 (N_12648,N_10898,N_11008);
or U12649 (N_12649,N_10541,N_11573);
nand U12650 (N_12650,N_11723,N_11344);
or U12651 (N_12651,N_9216,N_10994);
nand U12652 (N_12652,N_10383,N_11934);
and U12653 (N_12653,N_11132,N_10658);
and U12654 (N_12654,N_10308,N_10534);
nand U12655 (N_12655,N_11353,N_11077);
nor U12656 (N_12656,N_11564,N_10126);
nand U12657 (N_12657,N_11515,N_11682);
or U12658 (N_12658,N_9482,N_10702);
and U12659 (N_12659,N_9534,N_10591);
and U12660 (N_12660,N_10670,N_9262);
nand U12661 (N_12661,N_9160,N_11690);
and U12662 (N_12662,N_10333,N_11343);
or U12663 (N_12663,N_11731,N_9368);
and U12664 (N_12664,N_9545,N_11362);
or U12665 (N_12665,N_10634,N_10610);
or U12666 (N_12666,N_10074,N_10105);
nand U12667 (N_12667,N_11931,N_9402);
nor U12668 (N_12668,N_11228,N_10950);
nand U12669 (N_12669,N_11430,N_11771);
and U12670 (N_12670,N_10595,N_9045);
and U12671 (N_12671,N_11210,N_10881);
and U12672 (N_12672,N_11066,N_10903);
and U12673 (N_12673,N_11609,N_11367);
nor U12674 (N_12674,N_11915,N_9464);
and U12675 (N_12675,N_11330,N_9079);
xnor U12676 (N_12676,N_11743,N_9069);
nand U12677 (N_12677,N_10064,N_10485);
nor U12678 (N_12678,N_9112,N_11003);
nand U12679 (N_12679,N_11744,N_11527);
and U12680 (N_12680,N_9282,N_10299);
nand U12681 (N_12681,N_11615,N_10484);
xnor U12682 (N_12682,N_9499,N_10287);
nand U12683 (N_12683,N_10543,N_11624);
nor U12684 (N_12684,N_10036,N_10944);
nand U12685 (N_12685,N_11506,N_11399);
nor U12686 (N_12686,N_11966,N_11029);
xnor U12687 (N_12687,N_11017,N_9878);
or U12688 (N_12688,N_9308,N_11686);
nor U12689 (N_12689,N_9104,N_10831);
and U12690 (N_12690,N_11346,N_11032);
and U12691 (N_12691,N_10533,N_9719);
or U12692 (N_12692,N_9528,N_9834);
nor U12693 (N_12693,N_11879,N_11637);
or U12694 (N_12694,N_9948,N_10701);
nand U12695 (N_12695,N_10778,N_9352);
and U12696 (N_12696,N_11503,N_11488);
nand U12697 (N_12697,N_10166,N_9567);
nor U12698 (N_12698,N_10537,N_10677);
and U12699 (N_12699,N_9215,N_10759);
nand U12700 (N_12700,N_10275,N_11398);
xor U12701 (N_12701,N_9147,N_10808);
and U12702 (N_12702,N_9906,N_9796);
and U12703 (N_12703,N_10686,N_11131);
or U12704 (N_12704,N_9817,N_10068);
and U12705 (N_12705,N_9391,N_11891);
or U12706 (N_12706,N_9003,N_10519);
nor U12707 (N_12707,N_10437,N_10419);
nand U12708 (N_12708,N_10850,N_9988);
nand U12709 (N_12709,N_11846,N_11778);
or U12710 (N_12710,N_10909,N_10864);
nand U12711 (N_12711,N_11585,N_10503);
or U12712 (N_12712,N_10765,N_11413);
nor U12713 (N_12713,N_11649,N_11169);
and U12714 (N_12714,N_11471,N_10251);
nand U12715 (N_12715,N_11070,N_11796);
or U12716 (N_12716,N_10945,N_9909);
or U12717 (N_12717,N_9285,N_9628);
nor U12718 (N_12718,N_10358,N_11747);
or U12719 (N_12719,N_11999,N_11844);
nand U12720 (N_12720,N_10890,N_9724);
nor U12721 (N_12721,N_9837,N_11988);
and U12722 (N_12722,N_11082,N_11621);
nand U12723 (N_12723,N_9120,N_9116);
nand U12724 (N_12724,N_10857,N_10682);
nand U12725 (N_12725,N_11317,N_11927);
or U12726 (N_12726,N_11302,N_10605);
nand U12727 (N_12727,N_9358,N_11298);
nand U12728 (N_12728,N_9934,N_11732);
nor U12729 (N_12729,N_9866,N_10413);
or U12730 (N_12730,N_11902,N_9786);
nand U12731 (N_12731,N_10286,N_11824);
or U12732 (N_12732,N_11369,N_10757);
nor U12733 (N_12733,N_9338,N_10323);
or U12734 (N_12734,N_10583,N_10416);
nor U12735 (N_12735,N_11933,N_10526);
nor U12736 (N_12736,N_9284,N_9949);
or U12737 (N_12737,N_9075,N_11083);
or U12738 (N_12738,N_9943,N_11600);
and U12739 (N_12739,N_9276,N_11875);
nor U12740 (N_12740,N_11305,N_11851);
nand U12741 (N_12741,N_10423,N_10144);
nand U12742 (N_12742,N_9463,N_11000);
and U12743 (N_12743,N_9481,N_10509);
or U12744 (N_12744,N_11012,N_10128);
or U12745 (N_12745,N_11458,N_9327);
and U12746 (N_12746,N_11752,N_9092);
xor U12747 (N_12747,N_9835,N_10237);
or U12748 (N_12748,N_10790,N_10647);
or U12749 (N_12749,N_11072,N_9627);
nor U12750 (N_12750,N_11692,N_9772);
nand U12751 (N_12751,N_10466,N_9130);
or U12752 (N_12752,N_11854,N_10432);
nand U12753 (N_12753,N_11489,N_10660);
and U12754 (N_12754,N_10929,N_10748);
or U12755 (N_12755,N_11681,N_10852);
nand U12756 (N_12756,N_10740,N_11839);
nand U12757 (N_12757,N_9730,N_9477);
or U12758 (N_12758,N_11319,N_9746);
nor U12759 (N_12759,N_9205,N_9888);
nand U12760 (N_12760,N_9576,N_11808);
nand U12761 (N_12761,N_11081,N_10525);
and U12762 (N_12762,N_10936,N_11935);
or U12763 (N_12763,N_9822,N_10495);
nand U12764 (N_12764,N_11328,N_11924);
or U12765 (N_12765,N_9470,N_9336);
nor U12766 (N_12766,N_10121,N_9041);
or U12767 (N_12767,N_11701,N_9363);
and U12768 (N_12768,N_10346,N_11676);
and U12769 (N_12769,N_9653,N_11451);
and U12770 (N_12770,N_9618,N_11804);
and U12771 (N_12771,N_11646,N_10498);
or U12772 (N_12772,N_10956,N_11769);
or U12773 (N_12773,N_11449,N_10158);
and U12774 (N_12774,N_11098,N_10245);
and U12775 (N_12775,N_11279,N_11162);
or U12776 (N_12776,N_9221,N_9231);
and U12777 (N_12777,N_11662,N_10222);
nor U12778 (N_12778,N_9241,N_9111);
nand U12779 (N_12779,N_10340,N_10819);
and U12780 (N_12780,N_10637,N_10028);
and U12781 (N_12781,N_11951,N_11738);
and U12782 (N_12782,N_9538,N_10523);
or U12783 (N_12783,N_11272,N_11987);
nand U12784 (N_12784,N_10281,N_11559);
nand U12785 (N_12785,N_11698,N_11208);
or U12786 (N_12786,N_9013,N_10836);
nand U12787 (N_12787,N_9683,N_10133);
or U12788 (N_12788,N_11013,N_11550);
or U12789 (N_12789,N_10421,N_11726);
or U12790 (N_12790,N_9740,N_9905);
nor U12791 (N_12791,N_9879,N_9542);
and U12792 (N_12792,N_10352,N_10118);
and U12793 (N_12793,N_9170,N_9674);
or U12794 (N_12794,N_9443,N_9503);
nand U12795 (N_12795,N_9473,N_11641);
and U12796 (N_12796,N_11540,N_10993);
nor U12797 (N_12797,N_11720,N_10021);
and U12798 (N_12798,N_11446,N_9789);
and U12799 (N_12799,N_10762,N_10086);
or U12800 (N_12800,N_10426,N_11349);
and U12801 (N_12801,N_9353,N_10609);
and U12802 (N_12802,N_9963,N_9448);
nor U12803 (N_12803,N_10853,N_11350);
nor U12804 (N_12804,N_11910,N_9662);
nand U12805 (N_12805,N_11610,N_11719);
nand U12806 (N_12806,N_10794,N_10448);
nand U12807 (N_12807,N_11848,N_9367);
or U12808 (N_12808,N_10055,N_10155);
or U12809 (N_12809,N_11031,N_9224);
nand U12810 (N_12810,N_10408,N_10279);
nor U12811 (N_12811,N_10889,N_10802);
nor U12812 (N_12812,N_11187,N_9658);
and U12813 (N_12813,N_11960,N_9790);
or U12814 (N_12814,N_10854,N_10309);
nor U12815 (N_12815,N_10733,N_11170);
or U12816 (N_12816,N_9313,N_11002);
nand U12817 (N_12817,N_9987,N_11863);
nand U12818 (N_12818,N_9002,N_11351);
or U12819 (N_12819,N_9678,N_9998);
or U12820 (N_12820,N_11828,N_11204);
nand U12821 (N_12821,N_10154,N_10643);
nor U12822 (N_12822,N_11372,N_11118);
nand U12823 (N_12823,N_10402,N_11907);
nor U12824 (N_12824,N_10104,N_9225);
nor U12825 (N_12825,N_11116,N_10137);
or U12826 (N_12826,N_11360,N_9688);
or U12827 (N_12827,N_10476,N_11166);
nand U12828 (N_12828,N_9929,N_9895);
or U12829 (N_12829,N_10753,N_9516);
nor U12830 (N_12830,N_9454,N_9703);
and U12831 (N_12831,N_9836,N_9155);
and U12832 (N_12832,N_10848,N_10253);
nand U12833 (N_12833,N_9178,N_10392);
nand U12834 (N_12834,N_11718,N_11880);
nand U12835 (N_12835,N_11590,N_11022);
or U12836 (N_12836,N_10681,N_11842);
nor U12837 (N_12837,N_10257,N_11815);
and U12838 (N_12838,N_11384,N_11275);
xor U12839 (N_12839,N_10465,N_10775);
and U12840 (N_12840,N_11963,N_11643);
or U12841 (N_12841,N_10539,N_9393);
nand U12842 (N_12842,N_10703,N_11418);
nor U12843 (N_12843,N_9103,N_9310);
or U12844 (N_12844,N_9100,N_9029);
nand U12845 (N_12845,N_10692,N_9369);
and U12846 (N_12846,N_11865,N_10184);
and U12847 (N_12847,N_11256,N_11900);
and U12848 (N_12848,N_9269,N_10991);
nor U12849 (N_12849,N_10555,N_11253);
or U12850 (N_12850,N_11688,N_10292);
and U12851 (N_12851,N_9226,N_10264);
nor U12852 (N_12852,N_10827,N_11397);
nor U12853 (N_12853,N_9892,N_9930);
and U12854 (N_12854,N_10247,N_10435);
nor U12855 (N_12855,N_10277,N_11544);
nand U12856 (N_12856,N_9175,N_9077);
nor U12857 (N_12857,N_11146,N_10480);
or U12858 (N_12858,N_10355,N_11672);
nand U12859 (N_12859,N_11037,N_10463);
or U12860 (N_12860,N_10018,N_9483);
and U12861 (N_12861,N_9289,N_11847);
and U12862 (N_12862,N_10073,N_11557);
and U12863 (N_12863,N_10354,N_9452);
nor U12864 (N_12864,N_9259,N_11352);
or U12865 (N_12865,N_9515,N_9106);
and U12866 (N_12866,N_11232,N_9704);
and U12867 (N_12867,N_11182,N_10538);
or U12868 (N_12868,N_10125,N_10052);
nor U12869 (N_12869,N_9855,N_11391);
xor U12870 (N_12870,N_9429,N_11014);
nor U12871 (N_12871,N_10268,N_9518);
nand U12872 (N_12872,N_11807,N_9846);
xnor U12873 (N_12873,N_9901,N_11312);
or U12874 (N_12874,N_11759,N_10176);
nand U12875 (N_12875,N_9036,N_11831);
or U12876 (N_12876,N_11825,N_10450);
or U12877 (N_12877,N_9809,N_11427);
or U12878 (N_12878,N_9420,N_11908);
nor U12879 (N_12879,N_10005,N_11216);
nor U12880 (N_12880,N_11898,N_10905);
and U12881 (N_12881,N_9881,N_11465);
or U12882 (N_12882,N_11952,N_9328);
or U12883 (N_12883,N_10972,N_11786);
and U12884 (N_12884,N_9392,N_10460);
and U12885 (N_12885,N_9506,N_10161);
nor U12886 (N_12886,N_10870,N_11809);
and U12887 (N_12887,N_11826,N_11768);
or U12888 (N_12888,N_10569,N_9467);
or U12889 (N_12889,N_10152,N_11713);
nand U12890 (N_12890,N_11442,N_9449);
nand U12891 (N_12891,N_10820,N_9702);
or U12892 (N_12892,N_11301,N_10904);
nand U12893 (N_12893,N_10259,N_10481);
nor U12894 (N_12894,N_11997,N_9403);
and U12895 (N_12895,N_10369,N_9824);
or U12896 (N_12896,N_10668,N_9436);
nor U12897 (N_12897,N_11141,N_9376);
nor U12898 (N_12898,N_11377,N_11148);
nand U12899 (N_12899,N_11394,N_9696);
nand U12900 (N_12900,N_9261,N_11751);
or U12901 (N_12901,N_10667,N_11861);
or U12902 (N_12902,N_11177,N_11669);
nand U12903 (N_12903,N_11589,N_10261);
and U12904 (N_12904,N_11424,N_10654);
and U12905 (N_12905,N_9919,N_11986);
nand U12906 (N_12906,N_9735,N_10094);
and U12907 (N_12907,N_11356,N_10804);
nand U12908 (N_12908,N_10193,N_10027);
nor U12909 (N_12909,N_9279,N_9157);
nor U12910 (N_12910,N_9061,N_11456);
nand U12911 (N_12911,N_10729,N_11274);
nand U12912 (N_12912,N_10579,N_9517);
and U12913 (N_12913,N_9778,N_10896);
nor U12914 (N_12914,N_9918,N_9729);
nor U12915 (N_12915,N_9024,N_11019);
nand U12916 (N_12916,N_11764,N_11555);
and U12917 (N_12917,N_10388,N_11628);
or U12918 (N_12918,N_10342,N_9149);
nor U12919 (N_12919,N_10822,N_9217);
nor U12920 (N_12920,N_9137,N_9277);
and U12921 (N_12921,N_10912,N_9745);
and U12922 (N_12922,N_11636,N_11130);
and U12923 (N_12923,N_11145,N_10800);
nor U12924 (N_12924,N_9095,N_10517);
nand U12925 (N_12925,N_9093,N_11476);
xor U12926 (N_12926,N_9629,N_10798);
nand U12927 (N_12927,N_11774,N_9159);
nor U12928 (N_12928,N_9799,N_9033);
nor U12929 (N_12929,N_9938,N_10961);
and U12930 (N_12930,N_11981,N_11114);
and U12931 (N_12931,N_11027,N_11472);
and U12932 (N_12932,N_11257,N_11415);
or U12933 (N_12933,N_10999,N_10016);
and U12934 (N_12934,N_9127,N_11242);
or U12935 (N_12935,N_10741,N_10233);
or U12936 (N_12936,N_10880,N_10496);
or U12937 (N_12937,N_9316,N_10549);
and U12938 (N_12938,N_10283,N_9435);
nor U12939 (N_12939,N_10888,N_11428);
and U12940 (N_12940,N_11857,N_11547);
and U12941 (N_12941,N_11473,N_9913);
nand U12942 (N_12942,N_9253,N_10679);
nor U12943 (N_12943,N_11209,N_9768);
or U12944 (N_12944,N_10615,N_9526);
nand U12945 (N_12945,N_11603,N_9839);
and U12946 (N_12946,N_9646,N_9554);
nand U12947 (N_12947,N_9762,N_10711);
or U12948 (N_12948,N_9311,N_9364);
or U12949 (N_12949,N_9280,N_10454);
nor U12950 (N_12950,N_11054,N_11803);
nor U12951 (N_12951,N_11957,N_11393);
and U12952 (N_12952,N_10239,N_9570);
nand U12953 (N_12953,N_9590,N_11520);
or U12954 (N_12954,N_10070,N_11181);
or U12955 (N_12955,N_11968,N_10020);
nand U12956 (N_12956,N_11511,N_9858);
or U12957 (N_12957,N_11245,N_10190);
nand U12958 (N_12958,N_10473,N_9296);
or U12959 (N_12959,N_9599,N_9520);
or U12960 (N_12960,N_9115,N_9158);
nand U12961 (N_12961,N_9592,N_10520);
and U12962 (N_12962,N_11404,N_10875);
nor U12963 (N_12963,N_11583,N_9755);
nor U12964 (N_12964,N_10390,N_9738);
nand U12965 (N_12965,N_11300,N_11235);
nand U12966 (N_12966,N_9164,N_10887);
and U12967 (N_12967,N_10341,N_11493);
nor U12968 (N_12968,N_9935,N_9200);
or U12969 (N_12969,N_11011,N_11820);
nand U12970 (N_12970,N_9818,N_11929);
nor U12971 (N_12971,N_11697,N_10033);
nand U12972 (N_12972,N_11396,N_10895);
nand U12973 (N_12973,N_11874,N_9326);
nand U12974 (N_12974,N_11770,N_11920);
and U12975 (N_12975,N_10590,N_11985);
nand U12976 (N_12976,N_9787,N_9386);
and U12977 (N_12977,N_10722,N_10720);
nand U12978 (N_12978,N_11320,N_11914);
nor U12979 (N_12979,N_10225,N_11370);
and U12980 (N_12980,N_11249,N_9152);
nor U12981 (N_12981,N_11347,N_10099);
nor U12982 (N_12982,N_10149,N_11100);
or U12983 (N_12983,N_11876,N_9459);
nor U12984 (N_12984,N_10771,N_9562);
and U12985 (N_12985,N_11762,N_10727);
nand U12986 (N_12986,N_10234,N_11532);
and U12987 (N_12987,N_11750,N_11164);
or U12988 (N_12988,N_9811,N_11107);
or U12989 (N_12989,N_9591,N_11406);
or U12990 (N_12990,N_9922,N_11376);
and U12991 (N_12991,N_9889,N_9571);
and U12992 (N_12992,N_9995,N_9107);
and U12993 (N_12993,N_10367,N_11523);
or U12994 (N_12994,N_10269,N_9682);
or U12995 (N_12995,N_9999,N_10949);
nand U12996 (N_12996,N_10639,N_10726);
or U12997 (N_12997,N_10562,N_10928);
and U12998 (N_12998,N_10142,N_11945);
nand U12999 (N_12999,N_10925,N_9042);
nand U13000 (N_13000,N_11685,N_11509);
and U13001 (N_13001,N_11939,N_11689);
and U13002 (N_13002,N_11040,N_11482);
xnor U13003 (N_13003,N_11492,N_10678);
nor U13004 (N_13004,N_10789,N_11614);
and U13005 (N_13005,N_10312,N_10512);
nand U13006 (N_13006,N_9744,N_10403);
nand U13007 (N_13007,N_10131,N_10120);
nor U13008 (N_13008,N_9065,N_10689);
nand U13009 (N_13009,N_9113,N_10795);
nor U13010 (N_13010,N_11102,N_11959);
nor U13011 (N_13011,N_9345,N_10930);
and U13012 (N_13012,N_11411,N_10977);
and U13013 (N_13013,N_9625,N_9189);
or U13014 (N_13014,N_11562,N_10743);
or U13015 (N_13015,N_9339,N_11903);
nand U13016 (N_13016,N_10172,N_9699);
and U13017 (N_13017,N_10799,N_11297);
nor U13018 (N_13018,N_9633,N_10955);
or U13019 (N_13019,N_9097,N_10477);
nand U13020 (N_13020,N_9427,N_9652);
nor U13021 (N_13021,N_11680,N_10851);
nand U13022 (N_13022,N_9062,N_11357);
nand U13023 (N_13023,N_10011,N_9710);
nor U13024 (N_13024,N_10183,N_9663);
nand U13025 (N_13025,N_11135,N_9258);
nand U13026 (N_13026,N_9488,N_9961);
and U13027 (N_13027,N_11088,N_10461);
and U13028 (N_13028,N_10847,N_10026);
nand U13029 (N_13029,N_11119,N_11757);
or U13030 (N_13030,N_10414,N_11530);
nor U13031 (N_13031,N_11833,N_11288);
nand U13032 (N_13032,N_11469,N_9485);
nor U13033 (N_13033,N_9122,N_9958);
or U13034 (N_13034,N_10185,N_9348);
nor U13035 (N_13035,N_9419,N_11408);
and U13036 (N_13036,N_9519,N_11917);
nor U13037 (N_13037,N_11225,N_9602);
or U13038 (N_13038,N_11034,N_10508);
and U13039 (N_13039,N_9550,N_9679);
or U13040 (N_13040,N_9330,N_9997);
nor U13041 (N_13041,N_10400,N_11595);
or U13042 (N_13042,N_11395,N_9718);
nor U13043 (N_13043,N_11504,N_9377);
and U13044 (N_13044,N_10267,N_9335);
and U13045 (N_13045,N_10594,N_9600);
and U13046 (N_13046,N_11179,N_11129);
and U13047 (N_13047,N_9177,N_9793);
or U13048 (N_13048,N_9185,N_11371);
nand U13049 (N_13049,N_11716,N_10203);
and U13050 (N_13050,N_10089,N_10041);
nand U13051 (N_13051,N_11675,N_9052);
nor U13052 (N_13052,N_10103,N_10100);
or U13053 (N_13053,N_10129,N_9001);
nor U13054 (N_13054,N_11666,N_11025);
and U13055 (N_13055,N_10438,N_10194);
and U13056 (N_13056,N_9956,N_10329);
or U13057 (N_13057,N_10470,N_9243);
and U13058 (N_13058,N_9645,N_9445);
or U13059 (N_13059,N_9412,N_9705);
nor U13060 (N_13060,N_9844,N_10580);
nand U13061 (N_13061,N_9497,N_10328);
or U13062 (N_13062,N_9865,N_10401);
and U13063 (N_13063,N_9605,N_9845);
and U13064 (N_13064,N_10770,N_9747);
nor U13065 (N_13065,N_9341,N_10468);
nor U13066 (N_13066,N_11321,N_11651);
nand U13067 (N_13067,N_10177,N_11834);
and U13068 (N_13068,N_11381,N_11176);
or U13069 (N_13069,N_10553,N_10025);
and U13070 (N_13070,N_11246,N_10542);
or U13071 (N_13071,N_10969,N_11467);
nor U13072 (N_13072,N_9135,N_10965);
and U13073 (N_13073,N_9950,N_10760);
nor U13074 (N_13074,N_10926,N_10289);
and U13075 (N_13075,N_11422,N_10014);
and U13076 (N_13076,N_10801,N_9317);
or U13077 (N_13077,N_10130,N_10050);
nor U13078 (N_13078,N_9098,N_10311);
and U13079 (N_13079,N_11263,N_9749);
nand U13080 (N_13080,N_10174,N_11722);
nor U13081 (N_13081,N_9797,N_9860);
nand U13082 (N_13082,N_10053,N_10546);
or U13083 (N_13083,N_10502,N_9529);
or U13084 (N_13084,N_11466,N_10173);
or U13085 (N_13085,N_9661,N_11578);
nor U13086 (N_13086,N_9268,N_9505);
and U13087 (N_13087,N_10997,N_11715);
nand U13088 (N_13088,N_11736,N_9728);
and U13089 (N_13089,N_11956,N_9622);
or U13090 (N_13090,N_11264,N_9530);
or U13091 (N_13091,N_11111,N_11314);
nand U13092 (N_13092,N_11580,N_9446);
nand U13093 (N_13093,N_10168,N_9283);
or U13094 (N_13094,N_10112,N_11565);
nand U13095 (N_13095,N_11414,N_11195);
and U13096 (N_13096,N_10040,N_10954);
nor U13097 (N_13097,N_9321,N_11484);
nand U13098 (N_13098,N_9309,N_9842);
or U13099 (N_13099,N_10803,N_10879);
and U13100 (N_13100,N_9201,N_10787);
nand U13101 (N_13101,N_10444,N_10475);
nand U13102 (N_13102,N_11497,N_10023);
and U13103 (N_13103,N_11085,N_11837);
nor U13104 (N_13104,N_9465,N_11611);
nor U13105 (N_13105,N_10148,N_9507);
nor U13106 (N_13106,N_11124,N_11068);
nand U13107 (N_13107,N_9816,N_9032);
nor U13108 (N_13108,N_10867,N_10807);
and U13109 (N_13109,N_9597,N_9823);
and U13110 (N_13110,N_10716,N_11500);
or U13111 (N_13111,N_10980,N_9800);
nand U13112 (N_13112,N_10091,N_11593);
nand U13113 (N_13113,N_10098,N_11819);
nand U13114 (N_13114,N_10940,N_9196);
nor U13115 (N_13115,N_10684,N_9172);
and U13116 (N_13116,N_10059,N_10843);
nor U13117 (N_13117,N_10769,N_9199);
nor U13118 (N_13118,N_11090,N_9756);
and U13119 (N_13119,N_11872,N_9511);
nor U13120 (N_13120,N_10060,N_10970);
and U13121 (N_13121,N_10436,N_10514);
and U13122 (N_13122,N_11597,N_9804);
nand U13123 (N_13123,N_11501,N_9815);
nand U13124 (N_13124,N_10420,N_10841);
and U13125 (N_13125,N_9712,N_11958);
nand U13126 (N_13126,N_9428,N_9552);
or U13127 (N_13127,N_9959,N_10382);
nand U13128 (N_13128,N_10797,N_11513);
or U13129 (N_13129,N_10491,N_10941);
nor U13130 (N_13130,N_9371,N_9973);
nor U13131 (N_13131,N_11445,N_9154);
and U13132 (N_13132,N_11596,N_10394);
and U13133 (N_13133,N_11345,N_10732);
or U13134 (N_13134,N_9223,N_10349);
nor U13135 (N_13135,N_9848,N_9193);
and U13136 (N_13136,N_11536,N_10320);
nand U13137 (N_13137,N_9156,N_10492);
nand U13138 (N_13138,N_10622,N_10379);
nor U13139 (N_13139,N_10213,N_9173);
and U13140 (N_13140,N_9072,N_10724);
nor U13141 (N_13141,N_10680,N_11378);
or U13142 (N_13142,N_10821,N_10285);
and U13143 (N_13143,N_10004,N_11410);
nand U13144 (N_13144,N_11285,N_9706);
nor U13145 (N_13145,N_11775,N_9676);
nor U13146 (N_13146,N_10449,N_9639);
and U13147 (N_13147,N_9167,N_10433);
or U13148 (N_13148,N_10557,N_10300);
nand U13149 (N_13149,N_9140,N_10618);
nand U13150 (N_13150,N_9975,N_10581);
and U13151 (N_13151,N_10318,N_11730);
xor U13152 (N_13152,N_10931,N_9579);
and U13153 (N_13153,N_9501,N_9964);
and U13154 (N_13154,N_11237,N_11338);
nor U13155 (N_13155,N_10644,N_10598);
nand U13156 (N_13156,N_11431,N_11152);
and U13157 (N_13157,N_9307,N_9207);
nand U13158 (N_13158,N_11159,N_11767);
or U13159 (N_13159,N_11464,N_9826);
nor U13160 (N_13160,N_10044,N_10699);
nand U13161 (N_13161,N_9086,N_11745);
xnor U13162 (N_13162,N_10781,N_10673);
or U13163 (N_13163,N_10985,N_11160);
xor U13164 (N_13164,N_11400,N_9945);
nor U13165 (N_13165,N_10119,N_11901);
and U13166 (N_13166,N_11361,N_9928);
nor U13167 (N_13167,N_9166,N_9559);
nand U13168 (N_13168,N_11425,N_9085);
or U13169 (N_13169,N_9715,N_11605);
nor U13170 (N_13170,N_11843,N_11207);
or U13171 (N_13171,N_11158,N_10024);
and U13172 (N_13172,N_10665,N_9907);
and U13173 (N_13173,N_10296,N_9734);
or U13174 (N_13174,N_11026,N_9624);
nor U13175 (N_13175,N_9117,N_11139);
nand U13176 (N_13176,N_10374,N_9409);
nor U13177 (N_13177,N_11905,N_11254);
and U13178 (N_13178,N_11094,N_11277);
nor U13179 (N_13179,N_11969,N_10669);
nand U13180 (N_13180,N_9123,N_11105);
and U13181 (N_13181,N_10815,N_10326);
nor U13182 (N_13182,N_9732,N_10271);
nand U13183 (N_13183,N_11101,N_9176);
and U13184 (N_13184,N_11218,N_10824);
nand U13185 (N_13185,N_11766,N_10899);
and U13186 (N_13186,N_10325,N_10290);
nand U13187 (N_13187,N_9057,N_11282);
and U13188 (N_13188,N_9388,N_9870);
nor U13189 (N_13189,N_9876,N_11436);
nand U13190 (N_13190,N_10700,N_10774);
and U13191 (N_13191,N_9921,N_9299);
nor U13192 (N_13192,N_11852,N_10385);
and U13193 (N_13193,N_10132,N_9854);
or U13194 (N_13194,N_11822,N_11313);
nor U13195 (N_13195,N_11255,N_11708);
nand U13196 (N_13196,N_10313,N_9843);
nor U13197 (N_13197,N_11071,N_11433);
or U13198 (N_13198,N_10545,N_11233);
nor U13199 (N_13199,N_9690,N_11978);
and U13200 (N_13200,N_9847,N_11668);
nand U13201 (N_13201,N_10958,N_10835);
nor U13202 (N_13202,N_11976,N_11223);
and U13203 (N_13203,N_11203,N_9378);
or U13204 (N_13204,N_9916,N_11899);
nand U13205 (N_13205,N_10372,N_9769);
nand U13206 (N_13206,N_9575,N_10829);
nor U13207 (N_13207,N_9974,N_9381);
or U13208 (N_13208,N_9091,N_9713);
nor U13209 (N_13209,N_9785,N_9532);
nand U13210 (N_13210,N_9669,N_9632);
nor U13211 (N_13211,N_9491,N_11485);
nand U13212 (N_13212,N_10265,N_11444);
or U13213 (N_13213,N_11196,N_9192);
and U13214 (N_13214,N_10182,N_9198);
or U13215 (N_13215,N_11364,N_11702);
or U13216 (N_13216,N_10482,N_11853);
or U13217 (N_13217,N_9306,N_10635);
nand U13218 (N_13218,N_9849,N_10531);
nand U13219 (N_13219,N_10788,N_9957);
and U13220 (N_13220,N_10330,N_10363);
nor U13221 (N_13221,N_11311,N_9626);
nand U13222 (N_13222,N_9387,N_10165);
and U13223 (N_13223,N_9416,N_9426);
nand U13224 (N_13224,N_9180,N_10409);
nor U13225 (N_13225,N_11639,N_9188);
and U13226 (N_13226,N_11588,N_10756);
or U13227 (N_13227,N_11326,N_9701);
or U13228 (N_13228,N_10705,N_10574);
and U13229 (N_13229,N_10786,N_10572);
nand U13230 (N_13230,N_10135,N_9058);
or U13231 (N_13231,N_10900,N_11729);
or U13232 (N_13232,N_10893,N_9673);
nor U13233 (N_13233,N_9139,N_10003);
nor U13234 (N_13234,N_11420,N_10645);
nand U13235 (N_13235,N_9766,N_11335);
nor U13236 (N_13236,N_9737,N_10206);
and U13237 (N_13237,N_10187,N_10532);
or U13238 (N_13238,N_10938,N_11973);
nor U13239 (N_13239,N_9955,N_9803);
nand U13240 (N_13240,N_10652,N_11056);
nor U13241 (N_13241,N_10061,N_11188);
nand U13242 (N_13242,N_10638,N_11315);
nand U13243 (N_13243,N_10826,N_9236);
nor U13244 (N_13244,N_10685,N_10979);
nor U13245 (N_13245,N_11295,N_11220);
or U13246 (N_13246,N_11802,N_11630);
or U13247 (N_13247,N_11687,N_10659);
or U13248 (N_13248,N_11631,N_10085);
nor U13249 (N_13249,N_9006,N_9410);
nand U13250 (N_13250,N_9636,N_10548);
nor U13251 (N_13251,N_9614,N_9148);
or U13252 (N_13252,N_9814,N_11382);
and U13253 (N_13253,N_9487,N_10873);
nand U13254 (N_13254,N_10200,N_11016);
nor U13255 (N_13255,N_11558,N_11440);
and U13256 (N_13256,N_9875,N_11214);
or U13257 (N_13257,N_11659,N_11089);
nor U13258 (N_13258,N_10240,N_11995);
nor U13259 (N_13259,N_9862,N_10227);
nand U13260 (N_13260,N_10902,N_11136);
and U13261 (N_13261,N_11184,N_9754);
or U13262 (N_13262,N_10336,N_9108);
or U13263 (N_13263,N_11568,N_10839);
and U13264 (N_13264,N_11830,N_9752);
nand U13265 (N_13265,N_9894,N_9350);
and U13266 (N_13266,N_10518,N_10723);
nand U13267 (N_13267,N_11941,N_11375);
nor U13268 (N_13268,N_10139,N_10957);
and U13269 (N_13269,N_11093,N_9563);
nor U13270 (N_13270,N_10159,N_11009);
or U13271 (N_13271,N_10761,N_11109);
nor U13272 (N_13272,N_11694,N_10404);
and U13273 (N_13273,N_11211,N_9868);
and U13274 (N_13274,N_9260,N_10246);
or U13275 (N_13275,N_9292,N_11592);
nand U13276 (N_13276,N_10407,N_11021);
nor U13277 (N_13277,N_11392,N_11496);
and U13278 (N_13278,N_9642,N_9074);
or U13279 (N_13279,N_11276,N_9587);
nand U13280 (N_13280,N_11470,N_11632);
nand U13281 (N_13281,N_9936,N_9931);
nand U13282 (N_13282,N_9239,N_10430);
or U13283 (N_13283,N_9665,N_11982);
nor U13284 (N_13284,N_11783,N_10585);
or U13285 (N_13285,N_11541,N_10671);
and U13286 (N_13286,N_10693,N_10611);
nand U13287 (N_13287,N_10396,N_10990);
nand U13288 (N_13288,N_11895,N_11886);
nor U13289 (N_13289,N_10488,N_11103);
or U13290 (N_13290,N_9648,N_10058);
and U13291 (N_13291,N_9508,N_10513);
nand U13292 (N_13292,N_10776,N_10365);
nand U13293 (N_13293,N_11984,N_9256);
or U13294 (N_13294,N_9233,N_10946);
nand U13295 (N_13295,N_11096,N_11717);
nand U13296 (N_13296,N_11683,N_11737);
nor U13297 (N_13297,N_10709,N_10777);
and U13298 (N_13298,N_10731,N_11108);
and U13299 (N_13299,N_11441,N_10708);
nand U13300 (N_13300,N_10751,N_11001);
and U13301 (N_13301,N_9110,N_10256);
nor U13302 (N_13302,N_9810,N_9476);
nand U13303 (N_13303,N_10627,N_10515);
and U13304 (N_13304,N_9693,N_9978);
nor U13305 (N_13305,N_11267,N_10987);
or U13306 (N_13306,N_11495,N_9453);
and U13307 (N_13307,N_10886,N_9801);
nor U13308 (N_13308,N_11788,N_9885);
nand U13309 (N_13309,N_10536,N_11110);
or U13310 (N_13310,N_11052,N_11810);
nand U13311 (N_13311,N_9432,N_9318);
nand U13312 (N_13312,N_9018,N_11860);
nand U13313 (N_13313,N_11388,N_9711);
and U13314 (N_13314,N_10478,N_10111);
xnor U13315 (N_13315,N_9841,N_10698);
nor U13316 (N_13316,N_9054,N_9687);
nor U13317 (N_13317,N_9751,N_10834);
and U13318 (N_13318,N_9471,N_10577);
and U13319 (N_13319,N_10368,N_9494);
nand U13320 (N_13320,N_10143,N_9564);
or U13321 (N_13321,N_9991,N_11092);
nand U13322 (N_13322,N_11490,N_10646);
or U13323 (N_13323,N_9920,N_11653);
nand U13324 (N_13324,N_11354,N_9610);
nor U13325 (N_13325,N_9812,N_11280);
or U13326 (N_13326,N_9556,N_11741);
nand U13327 (N_13327,N_11890,N_11538);
and U13328 (N_13328,N_11283,N_9424);
and U13329 (N_13329,N_11827,N_10666);
and U13330 (N_13330,N_9914,N_9267);
nand U13331 (N_13331,N_10876,N_11193);
nand U13332 (N_13332,N_9265,N_11006);
nor U13333 (N_13333,N_9051,N_10582);
and U13334 (N_13334,N_9302,N_9329);
nand U13335 (N_13335,N_10924,N_11036);
nor U13336 (N_13336,N_9138,N_11735);
nand U13337 (N_13337,N_9828,N_9555);
nand U13338 (N_13338,N_9414,N_11358);
nor U13339 (N_13339,N_11965,N_11194);
nand U13340 (N_13340,N_10212,N_10764);
nand U13341 (N_13341,N_10229,N_11638);
nand U13342 (N_13342,N_10474,N_10922);
nand U13343 (N_13343,N_10273,N_10596);
nor U13344 (N_13344,N_11407,N_10395);
or U13345 (N_13345,N_9028,N_9034);
or U13346 (N_13346,N_10469,N_11859);
or U13347 (N_13347,N_9601,N_9340);
nor U13348 (N_13348,N_9025,N_9357);
or U13349 (N_13349,N_10180,N_10304);
and U13350 (N_13350,N_11763,N_10013);
nand U13351 (N_13351,N_11030,N_10766);
or U13352 (N_13352,N_9638,N_9742);
nand U13353 (N_13353,N_10110,N_9670);
and U13354 (N_13354,N_10691,N_11739);
and U13355 (N_13355,N_9851,N_11793);
or U13356 (N_13356,N_10083,N_11868);
and U13357 (N_13357,N_11140,N_9204);
nand U13358 (N_13358,N_10452,N_9194);
nand U13359 (N_13359,N_11432,N_9361);
and U13360 (N_13360,N_10160,N_10266);
or U13361 (N_13361,N_11412,N_9584);
or U13362 (N_13362,N_9792,N_10578);
nor U13363 (N_13363,N_10209,N_9102);
xor U13364 (N_13364,N_10943,N_11150);
nor U13365 (N_13365,N_10809,N_10694);
nor U13366 (N_13366,N_11477,N_10017);
and U13367 (N_13367,N_11383,N_9623);
xor U13368 (N_13368,N_10608,N_10062);
or U13369 (N_13369,N_9009,N_10713);
or U13370 (N_13370,N_10442,N_11368);
nor U13371 (N_13371,N_10202,N_10862);
or U13372 (N_13372,N_9763,N_11942);
and U13373 (N_13373,N_9222,N_9047);
nand U13374 (N_13374,N_10891,N_10657);
nand U13375 (N_13375,N_9394,N_11198);
or U13376 (N_13376,N_9305,N_11033);
and U13377 (N_13377,N_10348,N_10138);
nor U13378 (N_13378,N_10101,N_11576);
and U13379 (N_13379,N_10640,N_11642);
and U13380 (N_13380,N_10387,N_10297);
nor U13381 (N_13381,N_11888,N_10389);
or U13382 (N_13382,N_10191,N_9621);
nand U13383 (N_13383,N_10108,N_9252);
or U13384 (N_13384,N_9210,N_9382);
or U13385 (N_13385,N_9952,N_11005);
xor U13386 (N_13386,N_11849,N_9750);
or U13387 (N_13387,N_10869,N_9451);
and U13388 (N_13388,N_10785,N_9863);
and U13389 (N_13389,N_10558,N_10613);
nand U13390 (N_13390,N_9425,N_10630);
nor U13391 (N_13391,N_10636,N_9206);
or U13392 (N_13392,N_9781,N_10544);
nand U13393 (N_13393,N_11835,N_11727);
nand U13394 (N_13394,N_11667,N_11671);
and U13395 (N_13395,N_11127,N_9153);
nor U13396 (N_13396,N_10706,N_11309);
nand U13397 (N_13397,N_10833,N_9923);
and U13398 (N_13398,N_9540,N_11355);
nand U13399 (N_13399,N_9235,N_11584);
or U13400 (N_13400,N_10248,N_10939);
nor U13401 (N_13401,N_10506,N_10725);
nor U13402 (N_13402,N_9996,N_10032);
and U13403 (N_13403,N_11882,N_9105);
or U13404 (N_13404,N_10721,N_10037);
nor U13405 (N_13405,N_11572,N_10576);
nor U13406 (N_13406,N_10507,N_9068);
nor U13407 (N_13407,N_11024,N_11925);
nor U13408 (N_13408,N_11379,N_11937);
nor U13409 (N_13409,N_11239,N_10406);
nor U13410 (N_13410,N_9240,N_10570);
and U13411 (N_13411,N_9322,N_10270);
nand U13412 (N_13412,N_10226,N_11348);
or U13413 (N_13413,N_10364,N_10742);
nor U13414 (N_13414,N_10612,N_11677);
or U13415 (N_13415,N_10791,N_11084);
nand U13416 (N_13416,N_9300,N_10211);
nand U13417 (N_13417,N_9078,N_11205);
and U13418 (N_13418,N_11812,N_11386);
nand U13419 (N_13419,N_9161,N_10818);
or U13420 (N_13420,N_9544,N_9748);
nand U13421 (N_13421,N_9937,N_9362);
nor U13422 (N_13422,N_11897,N_11217);
nor U13423 (N_13423,N_11705,N_9976);
nor U13424 (N_13424,N_9725,N_9856);
or U13425 (N_13425,N_11780,N_11120);
nor U13426 (N_13426,N_10773,N_9775);
nor U13427 (N_13427,N_10920,N_10232);
nor U13428 (N_13428,N_9553,N_9512);
and U13429 (N_13429,N_11813,N_9932);
xor U13430 (N_13430,N_9456,N_11946);
and U13431 (N_13431,N_10556,N_10838);
nor U13432 (N_13432,N_10384,N_10057);
and U13433 (N_13433,N_11452,N_11171);
nor U13434 (N_13434,N_11569,N_10768);
or U13435 (N_13435,N_10284,N_10208);
and U13436 (N_13436,N_11955,N_9767);
or U13437 (N_13437,N_10840,N_9131);
nand U13438 (N_13438,N_10431,N_10968);
nor U13439 (N_13439,N_11797,N_9437);
nor U13440 (N_13440,N_9119,N_10324);
nand U13441 (N_13441,N_11525,N_9250);
nand U13442 (N_13442,N_11964,N_10035);
and U13443 (N_13443,N_11561,N_11439);
or U13444 (N_13444,N_9586,N_11553);
nand U13445 (N_13445,N_9423,N_9659);
or U13446 (N_13446,N_9890,N_11949);
nor U13447 (N_13447,N_10065,N_11387);
or U13448 (N_13448,N_11928,N_10201);
or U13449 (N_13449,N_10350,N_11617);
and U13450 (N_13450,N_9021,N_10784);
and U13451 (N_13451,N_10750,N_10293);
or U13452 (N_13452,N_10071,N_9620);
nor U13453 (N_13453,N_11390,N_11674);
and U13454 (N_13454,N_10097,N_11168);
nor U13455 (N_13455,N_11537,N_11438);
nor U13456 (N_13456,N_11816,N_10859);
and U13457 (N_13457,N_11461,N_11602);
nor U13458 (N_13458,N_9325,N_9015);
or U13459 (N_13459,N_11310,N_9304);
nor U13460 (N_13460,N_9672,N_10767);
nor U13461 (N_13461,N_11126,N_10882);
nor U13462 (N_13462,N_10031,N_10967);
or U13463 (N_13463,N_10215,N_9484);
or U13464 (N_13464,N_9441,N_9607);
and U13465 (N_13465,N_11800,N_11122);
or U13466 (N_13466,N_11728,N_11855);
nor U13467 (N_13467,N_9469,N_11307);
nand U13468 (N_13468,N_10567,N_10084);
and U13469 (N_13469,N_10715,N_10522);
or U13470 (N_13470,N_10282,N_11896);
nand U13471 (N_13471,N_10674,N_11161);
or U13472 (N_13472,N_9246,N_9360);
and U13473 (N_13473,N_10780,N_11137);
nor U13474 (N_13474,N_10500,N_10332);
and U13475 (N_13475,N_10877,N_11262);
nand U13476 (N_13476,N_9595,N_11814);
nor U13477 (N_13477,N_11286,N_9990);
and U13478 (N_13478,N_9230,N_9121);
or U13479 (N_13479,N_11740,N_9857);
or U13480 (N_13480,N_10650,N_11821);
or U13481 (N_13481,N_10381,N_10236);
nand U13482 (N_13482,N_10504,N_10487);
nand U13483 (N_13483,N_9779,N_11652);
nor U13484 (N_13484,N_10755,N_9049);
and U13485 (N_13485,N_9433,N_10907);
nor U13486 (N_13486,N_9186,N_9965);
nand U13487 (N_13487,N_10219,N_10690);
or U13488 (N_13488,N_11519,N_9248);
and U13489 (N_13489,N_10633,N_10238);
and U13490 (N_13490,N_11138,N_9271);
or U13491 (N_13491,N_10989,N_9864);
nand U13492 (N_13492,N_9099,N_11806);
or U13493 (N_13493,N_11416,N_11293);
and U13494 (N_13494,N_11340,N_9040);
or U13495 (N_13495,N_10573,N_10810);
nand U13496 (N_13496,N_11373,N_11046);
nand U13497 (N_13497,N_10255,N_11042);
or U13498 (N_13498,N_9580,N_9871);
nor U13499 (N_13499,N_10216,N_10424);
nor U13500 (N_13500,N_10457,N_9830);
nand U13501 (N_13501,N_11502,N_10085);
and U13502 (N_13502,N_11452,N_11985);
nand U13503 (N_13503,N_11961,N_11216);
or U13504 (N_13504,N_9950,N_11182);
nand U13505 (N_13505,N_11466,N_11968);
nand U13506 (N_13506,N_11725,N_11332);
nor U13507 (N_13507,N_11500,N_10230);
nand U13508 (N_13508,N_11780,N_11128);
nor U13509 (N_13509,N_9348,N_10482);
and U13510 (N_13510,N_10598,N_11354);
nand U13511 (N_13511,N_9116,N_9064);
nor U13512 (N_13512,N_11910,N_10904);
or U13513 (N_13513,N_11151,N_9703);
and U13514 (N_13514,N_11271,N_11346);
nand U13515 (N_13515,N_9496,N_11318);
nor U13516 (N_13516,N_9987,N_9276);
or U13517 (N_13517,N_11297,N_10270);
nor U13518 (N_13518,N_11864,N_11053);
or U13519 (N_13519,N_10462,N_9165);
and U13520 (N_13520,N_9179,N_10818);
nand U13521 (N_13521,N_11293,N_9061);
nor U13522 (N_13522,N_11145,N_9627);
nand U13523 (N_13523,N_10711,N_10614);
and U13524 (N_13524,N_9905,N_9223);
nor U13525 (N_13525,N_11752,N_11960);
nor U13526 (N_13526,N_9995,N_9499);
nor U13527 (N_13527,N_9496,N_9042);
nor U13528 (N_13528,N_10326,N_10281);
xnor U13529 (N_13529,N_10485,N_9413);
and U13530 (N_13530,N_9445,N_9967);
or U13531 (N_13531,N_9743,N_9476);
or U13532 (N_13532,N_9813,N_11643);
and U13533 (N_13533,N_9745,N_9183);
or U13534 (N_13534,N_10512,N_11870);
or U13535 (N_13535,N_11817,N_10012);
nor U13536 (N_13536,N_10536,N_10785);
and U13537 (N_13537,N_10305,N_10322);
nand U13538 (N_13538,N_11703,N_10395);
nand U13539 (N_13539,N_11584,N_9420);
nor U13540 (N_13540,N_9717,N_11954);
nand U13541 (N_13541,N_11738,N_10863);
and U13542 (N_13542,N_10177,N_10530);
and U13543 (N_13543,N_9693,N_9851);
nor U13544 (N_13544,N_10007,N_9239);
and U13545 (N_13545,N_10038,N_9123);
nand U13546 (N_13546,N_9867,N_10890);
nor U13547 (N_13547,N_11405,N_9334);
nor U13548 (N_13548,N_9383,N_9406);
nand U13549 (N_13549,N_9577,N_9075);
or U13550 (N_13550,N_10329,N_10961);
or U13551 (N_13551,N_11209,N_11034);
and U13552 (N_13552,N_11995,N_11615);
or U13553 (N_13553,N_11320,N_11801);
nand U13554 (N_13554,N_11444,N_10284);
nor U13555 (N_13555,N_9256,N_9904);
nand U13556 (N_13556,N_9509,N_11435);
nand U13557 (N_13557,N_11083,N_10196);
nand U13558 (N_13558,N_11708,N_9983);
nand U13559 (N_13559,N_9802,N_11128);
nand U13560 (N_13560,N_9414,N_10429);
nor U13561 (N_13561,N_10041,N_9314);
and U13562 (N_13562,N_11174,N_11286);
or U13563 (N_13563,N_10382,N_10503);
nor U13564 (N_13564,N_11710,N_10537);
and U13565 (N_13565,N_10922,N_10544);
and U13566 (N_13566,N_11605,N_10454);
and U13567 (N_13567,N_9278,N_10084);
and U13568 (N_13568,N_10098,N_11871);
nor U13569 (N_13569,N_10855,N_10740);
and U13570 (N_13570,N_11591,N_11982);
or U13571 (N_13571,N_10521,N_11081);
or U13572 (N_13572,N_10604,N_9947);
or U13573 (N_13573,N_9434,N_10019);
nor U13574 (N_13574,N_11520,N_10475);
and U13575 (N_13575,N_11760,N_11429);
and U13576 (N_13576,N_9706,N_11876);
nand U13577 (N_13577,N_11236,N_10104);
and U13578 (N_13578,N_9197,N_10561);
nor U13579 (N_13579,N_10682,N_10077);
or U13580 (N_13580,N_11247,N_11311);
and U13581 (N_13581,N_10748,N_11256);
nand U13582 (N_13582,N_9262,N_11689);
nor U13583 (N_13583,N_11769,N_9199);
nand U13584 (N_13584,N_9003,N_10886);
or U13585 (N_13585,N_10365,N_9146);
nand U13586 (N_13586,N_10213,N_11920);
nor U13587 (N_13587,N_9281,N_11855);
or U13588 (N_13588,N_9707,N_10170);
xor U13589 (N_13589,N_10605,N_9430);
or U13590 (N_13590,N_9301,N_10995);
nor U13591 (N_13591,N_9255,N_9809);
nor U13592 (N_13592,N_10127,N_11395);
nand U13593 (N_13593,N_10129,N_9403);
nor U13594 (N_13594,N_11886,N_11632);
nand U13595 (N_13595,N_11173,N_11663);
nor U13596 (N_13596,N_11412,N_9909);
or U13597 (N_13597,N_11084,N_10502);
or U13598 (N_13598,N_10587,N_10330);
and U13599 (N_13599,N_10157,N_9050);
and U13600 (N_13600,N_10127,N_9577);
and U13601 (N_13601,N_11413,N_11631);
and U13602 (N_13602,N_9196,N_10581);
xnor U13603 (N_13603,N_11707,N_9410);
nor U13604 (N_13604,N_11676,N_9216);
and U13605 (N_13605,N_9921,N_9941);
and U13606 (N_13606,N_10098,N_10341);
nand U13607 (N_13607,N_9700,N_9847);
and U13608 (N_13608,N_11927,N_11163);
and U13609 (N_13609,N_9302,N_9480);
and U13610 (N_13610,N_9540,N_11840);
or U13611 (N_13611,N_10377,N_10802);
and U13612 (N_13612,N_11428,N_9528);
nor U13613 (N_13613,N_10764,N_9863);
and U13614 (N_13614,N_11759,N_9131);
or U13615 (N_13615,N_9580,N_9596);
nor U13616 (N_13616,N_11641,N_9060);
or U13617 (N_13617,N_10621,N_9417);
and U13618 (N_13618,N_10292,N_11826);
nor U13619 (N_13619,N_9847,N_9879);
nand U13620 (N_13620,N_9278,N_9200);
or U13621 (N_13621,N_10346,N_10200);
nand U13622 (N_13622,N_11226,N_9525);
and U13623 (N_13623,N_9303,N_9688);
and U13624 (N_13624,N_9534,N_11573);
nand U13625 (N_13625,N_11684,N_11237);
and U13626 (N_13626,N_10663,N_11617);
nor U13627 (N_13627,N_9665,N_11428);
or U13628 (N_13628,N_9178,N_9013);
nor U13629 (N_13629,N_9088,N_11053);
or U13630 (N_13630,N_11197,N_11218);
nor U13631 (N_13631,N_11266,N_10512);
or U13632 (N_13632,N_10697,N_9816);
nor U13633 (N_13633,N_9662,N_10731);
nand U13634 (N_13634,N_10525,N_9135);
nand U13635 (N_13635,N_11804,N_9484);
nand U13636 (N_13636,N_9953,N_11667);
nand U13637 (N_13637,N_9397,N_9076);
and U13638 (N_13638,N_10698,N_11038);
or U13639 (N_13639,N_11170,N_10443);
or U13640 (N_13640,N_10294,N_10939);
or U13641 (N_13641,N_11490,N_11984);
nand U13642 (N_13642,N_10366,N_9280);
or U13643 (N_13643,N_9827,N_9521);
or U13644 (N_13644,N_11364,N_9771);
nand U13645 (N_13645,N_10510,N_10937);
or U13646 (N_13646,N_9120,N_9417);
nor U13647 (N_13647,N_11949,N_11381);
nor U13648 (N_13648,N_9853,N_11997);
and U13649 (N_13649,N_9555,N_11821);
and U13650 (N_13650,N_10648,N_10056);
nand U13651 (N_13651,N_11364,N_11016);
nand U13652 (N_13652,N_11361,N_9464);
nor U13653 (N_13653,N_11511,N_9123);
nand U13654 (N_13654,N_9981,N_11317);
or U13655 (N_13655,N_11790,N_9186);
or U13656 (N_13656,N_10800,N_11531);
nor U13657 (N_13657,N_9619,N_11436);
nor U13658 (N_13658,N_11617,N_9409);
or U13659 (N_13659,N_9006,N_9610);
and U13660 (N_13660,N_10823,N_10133);
or U13661 (N_13661,N_9056,N_10417);
nand U13662 (N_13662,N_9013,N_10607);
and U13663 (N_13663,N_11547,N_9339);
or U13664 (N_13664,N_11664,N_11901);
nor U13665 (N_13665,N_9395,N_11887);
or U13666 (N_13666,N_10841,N_10131);
nand U13667 (N_13667,N_9420,N_10296);
nor U13668 (N_13668,N_11508,N_10348);
or U13669 (N_13669,N_11922,N_11577);
nand U13670 (N_13670,N_10377,N_9606);
nand U13671 (N_13671,N_10298,N_9369);
and U13672 (N_13672,N_11221,N_10876);
nor U13673 (N_13673,N_11192,N_9792);
or U13674 (N_13674,N_10246,N_11997);
or U13675 (N_13675,N_9914,N_10203);
or U13676 (N_13676,N_9053,N_11280);
nor U13677 (N_13677,N_9260,N_9293);
nor U13678 (N_13678,N_10855,N_11443);
nand U13679 (N_13679,N_11231,N_10353);
nand U13680 (N_13680,N_9217,N_11164);
nor U13681 (N_13681,N_10494,N_10896);
nor U13682 (N_13682,N_10502,N_9341);
or U13683 (N_13683,N_9559,N_9164);
nand U13684 (N_13684,N_10057,N_11465);
and U13685 (N_13685,N_11575,N_10917);
and U13686 (N_13686,N_11561,N_11903);
or U13687 (N_13687,N_9712,N_9355);
or U13688 (N_13688,N_11053,N_9704);
nor U13689 (N_13689,N_11379,N_9573);
nor U13690 (N_13690,N_9257,N_10634);
and U13691 (N_13691,N_10406,N_11128);
nand U13692 (N_13692,N_10812,N_11237);
nor U13693 (N_13693,N_11777,N_9246);
nand U13694 (N_13694,N_11129,N_10897);
nand U13695 (N_13695,N_9802,N_10249);
or U13696 (N_13696,N_11312,N_11560);
or U13697 (N_13697,N_9287,N_10136);
xnor U13698 (N_13698,N_11245,N_11037);
nand U13699 (N_13699,N_11869,N_10219);
nand U13700 (N_13700,N_10610,N_11718);
nand U13701 (N_13701,N_9710,N_9329);
or U13702 (N_13702,N_11905,N_11145);
nand U13703 (N_13703,N_9642,N_11100);
nor U13704 (N_13704,N_11224,N_11789);
and U13705 (N_13705,N_9182,N_10681);
nor U13706 (N_13706,N_9982,N_9478);
and U13707 (N_13707,N_11308,N_9540);
and U13708 (N_13708,N_9192,N_10808);
nand U13709 (N_13709,N_9158,N_11873);
and U13710 (N_13710,N_9451,N_11822);
and U13711 (N_13711,N_10365,N_11764);
nand U13712 (N_13712,N_10183,N_9299);
or U13713 (N_13713,N_10164,N_9420);
nor U13714 (N_13714,N_9266,N_10230);
nand U13715 (N_13715,N_9639,N_11078);
nor U13716 (N_13716,N_9301,N_11009);
nor U13717 (N_13717,N_9676,N_10926);
or U13718 (N_13718,N_11668,N_11893);
nor U13719 (N_13719,N_11299,N_11729);
nand U13720 (N_13720,N_10159,N_9397);
nand U13721 (N_13721,N_10454,N_11526);
nand U13722 (N_13722,N_9218,N_10830);
nor U13723 (N_13723,N_11536,N_9339);
nor U13724 (N_13724,N_11125,N_9050);
and U13725 (N_13725,N_9923,N_11616);
or U13726 (N_13726,N_9931,N_10255);
and U13727 (N_13727,N_10554,N_11578);
or U13728 (N_13728,N_10928,N_10888);
nor U13729 (N_13729,N_9851,N_9514);
nor U13730 (N_13730,N_10261,N_10380);
or U13731 (N_13731,N_10076,N_11246);
nand U13732 (N_13732,N_10929,N_9112);
or U13733 (N_13733,N_11421,N_10577);
or U13734 (N_13734,N_10656,N_11099);
xor U13735 (N_13735,N_10526,N_11592);
nor U13736 (N_13736,N_10368,N_10707);
and U13737 (N_13737,N_10870,N_10461);
nor U13738 (N_13738,N_11047,N_11763);
or U13739 (N_13739,N_9073,N_10185);
or U13740 (N_13740,N_10257,N_11272);
nor U13741 (N_13741,N_10859,N_10698);
and U13742 (N_13742,N_10128,N_11359);
and U13743 (N_13743,N_10317,N_11273);
nand U13744 (N_13744,N_10739,N_10845);
or U13745 (N_13745,N_10327,N_11232);
nand U13746 (N_13746,N_10138,N_9667);
or U13747 (N_13747,N_11986,N_10659);
and U13748 (N_13748,N_9239,N_9535);
nor U13749 (N_13749,N_10833,N_11581);
and U13750 (N_13750,N_11811,N_11818);
or U13751 (N_13751,N_9493,N_10041);
nor U13752 (N_13752,N_9046,N_10770);
nor U13753 (N_13753,N_9528,N_11206);
nand U13754 (N_13754,N_10148,N_10508);
and U13755 (N_13755,N_9037,N_9848);
or U13756 (N_13756,N_9995,N_11414);
xnor U13757 (N_13757,N_10494,N_11259);
xor U13758 (N_13758,N_9878,N_10103);
nand U13759 (N_13759,N_10548,N_9486);
and U13760 (N_13760,N_11399,N_10579);
or U13761 (N_13761,N_11495,N_11205);
or U13762 (N_13762,N_11774,N_11596);
or U13763 (N_13763,N_10166,N_10953);
or U13764 (N_13764,N_9322,N_11576);
nand U13765 (N_13765,N_10364,N_9465);
and U13766 (N_13766,N_10411,N_10919);
or U13767 (N_13767,N_9016,N_10680);
nor U13768 (N_13768,N_11484,N_10222);
or U13769 (N_13769,N_11628,N_11926);
nand U13770 (N_13770,N_10068,N_11759);
nand U13771 (N_13771,N_9990,N_9241);
or U13772 (N_13772,N_11417,N_9483);
or U13773 (N_13773,N_9093,N_10597);
nand U13774 (N_13774,N_10682,N_10705);
or U13775 (N_13775,N_9487,N_9587);
nor U13776 (N_13776,N_10611,N_9481);
and U13777 (N_13777,N_9217,N_9440);
nand U13778 (N_13778,N_10433,N_11886);
nor U13779 (N_13779,N_11349,N_9687);
or U13780 (N_13780,N_9741,N_11981);
and U13781 (N_13781,N_11801,N_10581);
and U13782 (N_13782,N_11856,N_9563);
nand U13783 (N_13783,N_9274,N_11522);
and U13784 (N_13784,N_10979,N_10015);
and U13785 (N_13785,N_11289,N_10714);
and U13786 (N_13786,N_10189,N_10588);
nor U13787 (N_13787,N_11072,N_11411);
and U13788 (N_13788,N_9753,N_9301);
or U13789 (N_13789,N_11014,N_9116);
nor U13790 (N_13790,N_10801,N_10147);
or U13791 (N_13791,N_10389,N_11939);
or U13792 (N_13792,N_10753,N_10500);
nor U13793 (N_13793,N_9260,N_11948);
and U13794 (N_13794,N_10402,N_9013);
nand U13795 (N_13795,N_10965,N_9235);
nand U13796 (N_13796,N_10172,N_9726);
nand U13797 (N_13797,N_10820,N_10779);
and U13798 (N_13798,N_10338,N_10722);
or U13799 (N_13799,N_9630,N_9267);
or U13800 (N_13800,N_10110,N_11778);
nor U13801 (N_13801,N_9670,N_11304);
or U13802 (N_13802,N_9408,N_11619);
nand U13803 (N_13803,N_9300,N_11341);
nor U13804 (N_13804,N_11877,N_10641);
or U13805 (N_13805,N_10719,N_10885);
nand U13806 (N_13806,N_10454,N_11185);
or U13807 (N_13807,N_11062,N_11774);
nand U13808 (N_13808,N_11287,N_9912);
and U13809 (N_13809,N_11878,N_11128);
and U13810 (N_13810,N_9886,N_9019);
and U13811 (N_13811,N_10280,N_10170);
or U13812 (N_13812,N_10248,N_9230);
and U13813 (N_13813,N_9898,N_9332);
or U13814 (N_13814,N_11322,N_10151);
nand U13815 (N_13815,N_9657,N_9628);
and U13816 (N_13816,N_10734,N_11198);
nand U13817 (N_13817,N_9854,N_11444);
and U13818 (N_13818,N_9902,N_10381);
nor U13819 (N_13819,N_9989,N_10295);
and U13820 (N_13820,N_9591,N_9802);
or U13821 (N_13821,N_10829,N_11979);
nand U13822 (N_13822,N_9555,N_11648);
and U13823 (N_13823,N_11331,N_9495);
or U13824 (N_13824,N_11198,N_10391);
and U13825 (N_13825,N_10023,N_11832);
or U13826 (N_13826,N_9680,N_9306);
or U13827 (N_13827,N_10509,N_10662);
nor U13828 (N_13828,N_10478,N_9995);
or U13829 (N_13829,N_9128,N_9624);
and U13830 (N_13830,N_11797,N_10836);
nand U13831 (N_13831,N_9060,N_11375);
or U13832 (N_13832,N_10392,N_11038);
nand U13833 (N_13833,N_9625,N_11141);
nand U13834 (N_13834,N_9272,N_11562);
nand U13835 (N_13835,N_10344,N_11665);
and U13836 (N_13836,N_9382,N_11165);
or U13837 (N_13837,N_10398,N_10028);
nand U13838 (N_13838,N_10162,N_11213);
nor U13839 (N_13839,N_11913,N_10199);
nand U13840 (N_13840,N_11178,N_9924);
or U13841 (N_13841,N_11778,N_10618);
nor U13842 (N_13842,N_10434,N_9575);
or U13843 (N_13843,N_9734,N_11013);
nor U13844 (N_13844,N_9388,N_11636);
or U13845 (N_13845,N_10011,N_10421);
nand U13846 (N_13846,N_11664,N_11242);
nand U13847 (N_13847,N_10718,N_9936);
and U13848 (N_13848,N_10965,N_11498);
or U13849 (N_13849,N_10584,N_10361);
or U13850 (N_13850,N_9734,N_11664);
nand U13851 (N_13851,N_9506,N_10836);
nand U13852 (N_13852,N_9905,N_10585);
nor U13853 (N_13853,N_9534,N_9647);
and U13854 (N_13854,N_9931,N_10572);
nand U13855 (N_13855,N_10746,N_11223);
and U13856 (N_13856,N_11902,N_11663);
or U13857 (N_13857,N_11801,N_9984);
nand U13858 (N_13858,N_9051,N_11623);
and U13859 (N_13859,N_9506,N_10413);
nand U13860 (N_13860,N_9705,N_11911);
or U13861 (N_13861,N_9356,N_10244);
nand U13862 (N_13862,N_9137,N_10938);
nor U13863 (N_13863,N_9683,N_9917);
or U13864 (N_13864,N_9172,N_10816);
or U13865 (N_13865,N_11991,N_9480);
or U13866 (N_13866,N_9196,N_9727);
and U13867 (N_13867,N_9437,N_10679);
nand U13868 (N_13868,N_10658,N_10502);
and U13869 (N_13869,N_11158,N_9852);
or U13870 (N_13870,N_9836,N_9228);
and U13871 (N_13871,N_10334,N_11401);
or U13872 (N_13872,N_9203,N_9980);
and U13873 (N_13873,N_11560,N_9900);
and U13874 (N_13874,N_9726,N_10676);
or U13875 (N_13875,N_9677,N_9964);
nor U13876 (N_13876,N_9488,N_11104);
nand U13877 (N_13877,N_9178,N_10123);
or U13878 (N_13878,N_9884,N_10832);
and U13879 (N_13879,N_10789,N_10588);
nor U13880 (N_13880,N_11517,N_11957);
nand U13881 (N_13881,N_11819,N_9812);
or U13882 (N_13882,N_9137,N_9112);
or U13883 (N_13883,N_11516,N_10520);
or U13884 (N_13884,N_11896,N_9966);
or U13885 (N_13885,N_10256,N_11443);
nor U13886 (N_13886,N_9466,N_11003);
and U13887 (N_13887,N_9059,N_11058);
and U13888 (N_13888,N_11448,N_11190);
nor U13889 (N_13889,N_10761,N_11736);
and U13890 (N_13890,N_9024,N_9698);
and U13891 (N_13891,N_10541,N_9607);
and U13892 (N_13892,N_11822,N_11278);
nand U13893 (N_13893,N_10622,N_11063);
nand U13894 (N_13894,N_11503,N_11408);
nand U13895 (N_13895,N_10205,N_9969);
nor U13896 (N_13896,N_9175,N_10842);
nor U13897 (N_13897,N_11637,N_9793);
or U13898 (N_13898,N_9238,N_9399);
or U13899 (N_13899,N_11971,N_9512);
nor U13900 (N_13900,N_9900,N_10578);
and U13901 (N_13901,N_10267,N_9487);
or U13902 (N_13902,N_9746,N_9263);
nand U13903 (N_13903,N_11200,N_10687);
nor U13904 (N_13904,N_9714,N_9146);
or U13905 (N_13905,N_9017,N_10741);
or U13906 (N_13906,N_11787,N_10978);
nor U13907 (N_13907,N_11398,N_9034);
or U13908 (N_13908,N_10944,N_10203);
or U13909 (N_13909,N_9348,N_11988);
nand U13910 (N_13910,N_11685,N_11558);
and U13911 (N_13911,N_10261,N_11576);
nor U13912 (N_13912,N_10570,N_10113);
nor U13913 (N_13913,N_11284,N_10505);
nand U13914 (N_13914,N_9695,N_11829);
nor U13915 (N_13915,N_10744,N_9785);
and U13916 (N_13916,N_9581,N_9129);
or U13917 (N_13917,N_10868,N_10197);
nor U13918 (N_13918,N_9290,N_9867);
or U13919 (N_13919,N_11108,N_9189);
nand U13920 (N_13920,N_9490,N_10642);
or U13921 (N_13921,N_10353,N_11901);
nand U13922 (N_13922,N_9057,N_11267);
nor U13923 (N_13923,N_11050,N_9063);
or U13924 (N_13924,N_9456,N_11558);
nor U13925 (N_13925,N_9732,N_10765);
or U13926 (N_13926,N_10689,N_9712);
nor U13927 (N_13927,N_9353,N_10895);
nor U13928 (N_13928,N_11382,N_11902);
or U13929 (N_13929,N_11405,N_10290);
and U13930 (N_13930,N_11789,N_10226);
nand U13931 (N_13931,N_11924,N_10971);
nand U13932 (N_13932,N_9303,N_10981);
and U13933 (N_13933,N_11632,N_11928);
and U13934 (N_13934,N_11757,N_11509);
and U13935 (N_13935,N_10165,N_11816);
nand U13936 (N_13936,N_11992,N_10973);
nand U13937 (N_13937,N_10281,N_10440);
nor U13938 (N_13938,N_11326,N_11750);
or U13939 (N_13939,N_9279,N_9536);
nand U13940 (N_13940,N_11567,N_11634);
nand U13941 (N_13941,N_11748,N_9739);
nor U13942 (N_13942,N_9129,N_10541);
and U13943 (N_13943,N_9823,N_10919);
nand U13944 (N_13944,N_9315,N_9504);
nor U13945 (N_13945,N_10391,N_11989);
or U13946 (N_13946,N_9633,N_10673);
or U13947 (N_13947,N_9232,N_10244);
and U13948 (N_13948,N_9680,N_9749);
and U13949 (N_13949,N_9793,N_10279);
nand U13950 (N_13950,N_11394,N_9294);
and U13951 (N_13951,N_10049,N_11883);
nor U13952 (N_13952,N_11724,N_11016);
nor U13953 (N_13953,N_9626,N_10245);
and U13954 (N_13954,N_10583,N_11679);
and U13955 (N_13955,N_10143,N_11540);
and U13956 (N_13956,N_11465,N_10666);
nor U13957 (N_13957,N_9289,N_9175);
nor U13958 (N_13958,N_10681,N_11188);
nand U13959 (N_13959,N_11727,N_11480);
nor U13960 (N_13960,N_11208,N_9180);
nor U13961 (N_13961,N_10966,N_9681);
and U13962 (N_13962,N_11395,N_10046);
nor U13963 (N_13963,N_11175,N_11552);
nor U13964 (N_13964,N_9389,N_10824);
or U13965 (N_13965,N_10937,N_10802);
nor U13966 (N_13966,N_10879,N_11172);
nand U13967 (N_13967,N_10232,N_11009);
nor U13968 (N_13968,N_9657,N_11034);
or U13969 (N_13969,N_11292,N_9299);
or U13970 (N_13970,N_9795,N_10668);
nand U13971 (N_13971,N_11662,N_9438);
or U13972 (N_13972,N_9797,N_11713);
and U13973 (N_13973,N_10373,N_9945);
nand U13974 (N_13974,N_10441,N_11606);
or U13975 (N_13975,N_11855,N_10723);
nor U13976 (N_13976,N_11526,N_10095);
and U13977 (N_13977,N_9269,N_11840);
nand U13978 (N_13978,N_9259,N_10339);
and U13979 (N_13979,N_9302,N_10632);
and U13980 (N_13980,N_11081,N_11842);
nand U13981 (N_13981,N_10624,N_11018);
nor U13982 (N_13982,N_11669,N_9388);
nand U13983 (N_13983,N_9101,N_9720);
nand U13984 (N_13984,N_9422,N_11638);
nor U13985 (N_13985,N_9120,N_10159);
and U13986 (N_13986,N_11393,N_9201);
nand U13987 (N_13987,N_11670,N_11439);
or U13988 (N_13988,N_10750,N_11680);
nand U13989 (N_13989,N_9163,N_9169);
nand U13990 (N_13990,N_11559,N_11508);
nand U13991 (N_13991,N_9225,N_9019);
or U13992 (N_13992,N_9608,N_10682);
and U13993 (N_13993,N_9696,N_9630);
and U13994 (N_13994,N_10133,N_11183);
nor U13995 (N_13995,N_11980,N_11916);
nand U13996 (N_13996,N_9320,N_11306);
or U13997 (N_13997,N_9871,N_9571);
nor U13998 (N_13998,N_10033,N_11567);
and U13999 (N_13999,N_10500,N_9395);
nand U14000 (N_14000,N_9870,N_11653);
or U14001 (N_14001,N_9002,N_11463);
nand U14002 (N_14002,N_9222,N_9755);
and U14003 (N_14003,N_9594,N_10523);
and U14004 (N_14004,N_11364,N_11561);
nor U14005 (N_14005,N_9740,N_10414);
nand U14006 (N_14006,N_10362,N_10857);
nor U14007 (N_14007,N_9200,N_9662);
or U14008 (N_14008,N_9672,N_11878);
or U14009 (N_14009,N_11954,N_9764);
or U14010 (N_14010,N_11296,N_10488);
or U14011 (N_14011,N_9133,N_11031);
nor U14012 (N_14012,N_10617,N_9614);
or U14013 (N_14013,N_11151,N_11793);
and U14014 (N_14014,N_10158,N_10522);
and U14015 (N_14015,N_10872,N_11227);
and U14016 (N_14016,N_9442,N_10971);
nand U14017 (N_14017,N_11866,N_9094);
nand U14018 (N_14018,N_9655,N_9132);
and U14019 (N_14019,N_11924,N_11281);
and U14020 (N_14020,N_10690,N_11588);
and U14021 (N_14021,N_11929,N_10133);
or U14022 (N_14022,N_9490,N_11724);
nor U14023 (N_14023,N_11883,N_10925);
nand U14024 (N_14024,N_11525,N_10247);
or U14025 (N_14025,N_11668,N_11706);
or U14026 (N_14026,N_9810,N_10269);
or U14027 (N_14027,N_11413,N_9997);
nand U14028 (N_14028,N_10982,N_9559);
nand U14029 (N_14029,N_9498,N_10184);
nor U14030 (N_14030,N_11116,N_9621);
or U14031 (N_14031,N_11891,N_10905);
nand U14032 (N_14032,N_10450,N_10063);
nand U14033 (N_14033,N_9603,N_10446);
and U14034 (N_14034,N_11820,N_10501);
nand U14035 (N_14035,N_11043,N_9557);
nand U14036 (N_14036,N_11907,N_11247);
nand U14037 (N_14037,N_9595,N_9965);
nor U14038 (N_14038,N_11571,N_11916);
nand U14039 (N_14039,N_9169,N_10799);
nor U14040 (N_14040,N_11993,N_9390);
nand U14041 (N_14041,N_11818,N_11187);
nor U14042 (N_14042,N_9227,N_11404);
and U14043 (N_14043,N_11857,N_10218);
and U14044 (N_14044,N_11440,N_11350);
nor U14045 (N_14045,N_10375,N_11016);
nand U14046 (N_14046,N_9271,N_11736);
nor U14047 (N_14047,N_10495,N_11531);
nor U14048 (N_14048,N_10960,N_9229);
nor U14049 (N_14049,N_9358,N_10504);
nand U14050 (N_14050,N_9120,N_9161);
or U14051 (N_14051,N_11078,N_10838);
or U14052 (N_14052,N_9597,N_11188);
and U14053 (N_14053,N_9866,N_10095);
nor U14054 (N_14054,N_11653,N_11946);
and U14055 (N_14055,N_9684,N_11222);
nor U14056 (N_14056,N_11697,N_11885);
and U14057 (N_14057,N_11787,N_10178);
nand U14058 (N_14058,N_11695,N_9705);
and U14059 (N_14059,N_11916,N_10884);
nand U14060 (N_14060,N_9388,N_10534);
and U14061 (N_14061,N_10477,N_10335);
and U14062 (N_14062,N_11171,N_11109);
nand U14063 (N_14063,N_11743,N_11745);
nand U14064 (N_14064,N_9382,N_10471);
nand U14065 (N_14065,N_9376,N_11591);
nor U14066 (N_14066,N_9644,N_11530);
or U14067 (N_14067,N_10698,N_10634);
nor U14068 (N_14068,N_10547,N_10801);
nor U14069 (N_14069,N_11171,N_11433);
and U14070 (N_14070,N_9680,N_11172);
nand U14071 (N_14071,N_11421,N_9684);
and U14072 (N_14072,N_11994,N_10254);
nand U14073 (N_14073,N_11260,N_9719);
or U14074 (N_14074,N_11840,N_11225);
and U14075 (N_14075,N_9244,N_9905);
nand U14076 (N_14076,N_9113,N_10074);
nand U14077 (N_14077,N_9307,N_9065);
nor U14078 (N_14078,N_10465,N_9419);
or U14079 (N_14079,N_11405,N_9775);
nor U14080 (N_14080,N_10180,N_9256);
xor U14081 (N_14081,N_11180,N_9286);
or U14082 (N_14082,N_10087,N_11964);
and U14083 (N_14083,N_10589,N_11057);
and U14084 (N_14084,N_10820,N_10050);
nand U14085 (N_14085,N_9412,N_10090);
nor U14086 (N_14086,N_11661,N_9842);
and U14087 (N_14087,N_11060,N_11421);
nand U14088 (N_14088,N_11354,N_11462);
and U14089 (N_14089,N_10178,N_10591);
and U14090 (N_14090,N_9217,N_10297);
or U14091 (N_14091,N_9787,N_11170);
and U14092 (N_14092,N_11231,N_9186);
nor U14093 (N_14093,N_11824,N_9595);
nand U14094 (N_14094,N_11439,N_9419);
nand U14095 (N_14095,N_10786,N_11172);
and U14096 (N_14096,N_9564,N_10600);
and U14097 (N_14097,N_9752,N_10587);
or U14098 (N_14098,N_10876,N_11873);
and U14099 (N_14099,N_10971,N_10096);
or U14100 (N_14100,N_9874,N_11094);
or U14101 (N_14101,N_11235,N_9811);
and U14102 (N_14102,N_10341,N_9631);
nand U14103 (N_14103,N_10015,N_10037);
or U14104 (N_14104,N_11026,N_11914);
and U14105 (N_14105,N_10916,N_10048);
or U14106 (N_14106,N_9365,N_10529);
nand U14107 (N_14107,N_11474,N_9036);
nor U14108 (N_14108,N_11026,N_10188);
nand U14109 (N_14109,N_10028,N_11294);
nor U14110 (N_14110,N_10763,N_9597);
and U14111 (N_14111,N_11080,N_9818);
nand U14112 (N_14112,N_10740,N_10045);
and U14113 (N_14113,N_10153,N_10562);
and U14114 (N_14114,N_10255,N_9592);
nor U14115 (N_14115,N_10029,N_11643);
or U14116 (N_14116,N_10258,N_9388);
and U14117 (N_14117,N_11516,N_10233);
nand U14118 (N_14118,N_9838,N_10169);
nand U14119 (N_14119,N_10714,N_11163);
and U14120 (N_14120,N_11228,N_10546);
or U14121 (N_14121,N_9005,N_11237);
and U14122 (N_14122,N_10248,N_10278);
nor U14123 (N_14123,N_11209,N_9957);
nand U14124 (N_14124,N_10013,N_11284);
and U14125 (N_14125,N_11426,N_10794);
nand U14126 (N_14126,N_11857,N_9470);
nor U14127 (N_14127,N_11192,N_10538);
nor U14128 (N_14128,N_9783,N_11179);
nor U14129 (N_14129,N_10126,N_11249);
or U14130 (N_14130,N_9643,N_10981);
and U14131 (N_14131,N_10632,N_11688);
nor U14132 (N_14132,N_10706,N_11169);
nor U14133 (N_14133,N_9812,N_9379);
nand U14134 (N_14134,N_11259,N_11434);
nor U14135 (N_14135,N_11863,N_9625);
and U14136 (N_14136,N_9892,N_9067);
nand U14137 (N_14137,N_9888,N_9258);
and U14138 (N_14138,N_9969,N_10275);
or U14139 (N_14139,N_10190,N_10552);
nor U14140 (N_14140,N_9628,N_9650);
nand U14141 (N_14141,N_11973,N_10332);
nor U14142 (N_14142,N_11491,N_10845);
nor U14143 (N_14143,N_11014,N_11041);
and U14144 (N_14144,N_9330,N_11730);
nand U14145 (N_14145,N_11980,N_11534);
or U14146 (N_14146,N_9759,N_9277);
nand U14147 (N_14147,N_10071,N_9998);
and U14148 (N_14148,N_11786,N_11951);
or U14149 (N_14149,N_9593,N_11491);
nor U14150 (N_14150,N_9797,N_9193);
nand U14151 (N_14151,N_11036,N_9963);
nand U14152 (N_14152,N_11679,N_9025);
and U14153 (N_14153,N_11410,N_9656);
and U14154 (N_14154,N_11149,N_11926);
or U14155 (N_14155,N_11005,N_9696);
nor U14156 (N_14156,N_11511,N_10338);
nand U14157 (N_14157,N_9506,N_10222);
xor U14158 (N_14158,N_9296,N_11025);
nand U14159 (N_14159,N_9289,N_10784);
xnor U14160 (N_14160,N_10665,N_11287);
and U14161 (N_14161,N_10829,N_9596);
and U14162 (N_14162,N_9801,N_10212);
and U14163 (N_14163,N_11129,N_10310);
nor U14164 (N_14164,N_11556,N_10984);
nor U14165 (N_14165,N_11223,N_9340);
and U14166 (N_14166,N_11984,N_9025);
nand U14167 (N_14167,N_10783,N_10487);
nor U14168 (N_14168,N_10469,N_9677);
and U14169 (N_14169,N_10999,N_10193);
nand U14170 (N_14170,N_11423,N_11628);
nand U14171 (N_14171,N_10295,N_11381);
nand U14172 (N_14172,N_11962,N_9588);
nor U14173 (N_14173,N_9725,N_11025);
nand U14174 (N_14174,N_11856,N_9366);
and U14175 (N_14175,N_9878,N_9154);
and U14176 (N_14176,N_11686,N_10324);
and U14177 (N_14177,N_9826,N_10675);
nand U14178 (N_14178,N_9811,N_11096);
or U14179 (N_14179,N_11246,N_10846);
nand U14180 (N_14180,N_10129,N_11577);
and U14181 (N_14181,N_11306,N_11920);
and U14182 (N_14182,N_9822,N_11528);
nand U14183 (N_14183,N_9627,N_9794);
nor U14184 (N_14184,N_10258,N_9694);
nor U14185 (N_14185,N_9143,N_11903);
nand U14186 (N_14186,N_11474,N_11522);
and U14187 (N_14187,N_9771,N_10831);
nand U14188 (N_14188,N_9171,N_11396);
nand U14189 (N_14189,N_11602,N_9487);
nor U14190 (N_14190,N_11682,N_11953);
nand U14191 (N_14191,N_9826,N_11922);
and U14192 (N_14192,N_9972,N_10046);
or U14193 (N_14193,N_10632,N_10957);
nor U14194 (N_14194,N_11247,N_10259);
and U14195 (N_14195,N_9735,N_10018);
nand U14196 (N_14196,N_9737,N_9705);
nand U14197 (N_14197,N_9387,N_9620);
xnor U14198 (N_14198,N_11693,N_9552);
nor U14199 (N_14199,N_11546,N_11130);
nand U14200 (N_14200,N_9932,N_10685);
nor U14201 (N_14201,N_9133,N_10937);
and U14202 (N_14202,N_9093,N_11098);
nand U14203 (N_14203,N_11180,N_11082);
nand U14204 (N_14204,N_10474,N_9876);
and U14205 (N_14205,N_10247,N_11991);
or U14206 (N_14206,N_10197,N_9180);
nor U14207 (N_14207,N_10429,N_9932);
and U14208 (N_14208,N_9145,N_9233);
or U14209 (N_14209,N_9996,N_11205);
nand U14210 (N_14210,N_11643,N_11909);
nand U14211 (N_14211,N_11970,N_11528);
nand U14212 (N_14212,N_10979,N_11042);
nor U14213 (N_14213,N_10476,N_11441);
and U14214 (N_14214,N_9156,N_10401);
nor U14215 (N_14215,N_11899,N_10055);
nand U14216 (N_14216,N_11337,N_9077);
nor U14217 (N_14217,N_9004,N_9177);
and U14218 (N_14218,N_9344,N_11590);
or U14219 (N_14219,N_11322,N_9237);
nand U14220 (N_14220,N_10701,N_10192);
or U14221 (N_14221,N_11277,N_10218);
nor U14222 (N_14222,N_11691,N_10811);
and U14223 (N_14223,N_10659,N_10583);
nand U14224 (N_14224,N_10724,N_11081);
or U14225 (N_14225,N_11705,N_11511);
or U14226 (N_14226,N_9079,N_10084);
nor U14227 (N_14227,N_10883,N_11368);
nand U14228 (N_14228,N_9811,N_10102);
nand U14229 (N_14229,N_10592,N_9610);
nand U14230 (N_14230,N_9675,N_10128);
or U14231 (N_14231,N_9560,N_9714);
or U14232 (N_14232,N_11666,N_11562);
nor U14233 (N_14233,N_11633,N_10768);
or U14234 (N_14234,N_11241,N_10760);
nand U14235 (N_14235,N_11629,N_11030);
nand U14236 (N_14236,N_11947,N_10091);
or U14237 (N_14237,N_11340,N_11818);
nor U14238 (N_14238,N_11035,N_9198);
and U14239 (N_14239,N_10681,N_10163);
nand U14240 (N_14240,N_9425,N_10057);
nor U14241 (N_14241,N_9020,N_10882);
nand U14242 (N_14242,N_9213,N_10285);
nand U14243 (N_14243,N_11057,N_9131);
nor U14244 (N_14244,N_11366,N_11399);
and U14245 (N_14245,N_11386,N_10404);
nand U14246 (N_14246,N_10987,N_9679);
and U14247 (N_14247,N_10016,N_11459);
nand U14248 (N_14248,N_10568,N_10853);
and U14249 (N_14249,N_10234,N_9303);
nand U14250 (N_14250,N_10570,N_10596);
nor U14251 (N_14251,N_10845,N_9120);
or U14252 (N_14252,N_10785,N_10013);
nand U14253 (N_14253,N_11602,N_10417);
and U14254 (N_14254,N_11773,N_9846);
or U14255 (N_14255,N_11234,N_11874);
nand U14256 (N_14256,N_11635,N_9466);
nand U14257 (N_14257,N_9010,N_10750);
and U14258 (N_14258,N_11709,N_11663);
and U14259 (N_14259,N_11868,N_11084);
nor U14260 (N_14260,N_11167,N_11320);
nor U14261 (N_14261,N_9935,N_9746);
nand U14262 (N_14262,N_10636,N_9940);
or U14263 (N_14263,N_11882,N_10424);
nor U14264 (N_14264,N_9004,N_11695);
nor U14265 (N_14265,N_9882,N_10923);
nor U14266 (N_14266,N_11444,N_10518);
and U14267 (N_14267,N_9329,N_11503);
and U14268 (N_14268,N_10266,N_10717);
and U14269 (N_14269,N_11917,N_9127);
nor U14270 (N_14270,N_10264,N_9063);
nor U14271 (N_14271,N_10411,N_10944);
nor U14272 (N_14272,N_10285,N_10252);
nor U14273 (N_14273,N_10363,N_10833);
or U14274 (N_14274,N_11693,N_10333);
nor U14275 (N_14275,N_9103,N_11752);
and U14276 (N_14276,N_10030,N_9611);
and U14277 (N_14277,N_9215,N_10743);
nor U14278 (N_14278,N_10645,N_10376);
nor U14279 (N_14279,N_10527,N_10466);
nand U14280 (N_14280,N_9603,N_11864);
nand U14281 (N_14281,N_9345,N_10069);
or U14282 (N_14282,N_9892,N_11061);
nor U14283 (N_14283,N_9687,N_10308);
and U14284 (N_14284,N_11346,N_11964);
nand U14285 (N_14285,N_11674,N_11844);
nand U14286 (N_14286,N_11100,N_10300);
nor U14287 (N_14287,N_11212,N_11171);
nor U14288 (N_14288,N_11559,N_10447);
nand U14289 (N_14289,N_9808,N_11904);
or U14290 (N_14290,N_11994,N_9099);
nand U14291 (N_14291,N_10270,N_11173);
nor U14292 (N_14292,N_9478,N_11737);
nand U14293 (N_14293,N_10907,N_11918);
nor U14294 (N_14294,N_11915,N_10080);
nor U14295 (N_14295,N_9570,N_9870);
nand U14296 (N_14296,N_9010,N_10971);
nand U14297 (N_14297,N_9421,N_10073);
and U14298 (N_14298,N_10180,N_10781);
nand U14299 (N_14299,N_10974,N_10173);
nor U14300 (N_14300,N_11970,N_11346);
nand U14301 (N_14301,N_9431,N_10744);
nor U14302 (N_14302,N_10513,N_10917);
nand U14303 (N_14303,N_11078,N_11318);
nor U14304 (N_14304,N_11410,N_9576);
and U14305 (N_14305,N_10450,N_9441);
nor U14306 (N_14306,N_9437,N_10802);
nor U14307 (N_14307,N_9684,N_10005);
or U14308 (N_14308,N_9135,N_10491);
nand U14309 (N_14309,N_11925,N_10633);
or U14310 (N_14310,N_10338,N_11425);
nand U14311 (N_14311,N_9707,N_9813);
or U14312 (N_14312,N_11301,N_11058);
and U14313 (N_14313,N_11618,N_9973);
nand U14314 (N_14314,N_9800,N_10148);
or U14315 (N_14315,N_10483,N_10195);
xor U14316 (N_14316,N_11860,N_10532);
and U14317 (N_14317,N_10126,N_10359);
nand U14318 (N_14318,N_11887,N_9267);
nor U14319 (N_14319,N_9819,N_10386);
nor U14320 (N_14320,N_10938,N_10592);
nand U14321 (N_14321,N_11146,N_10924);
nand U14322 (N_14322,N_10786,N_10564);
and U14323 (N_14323,N_10020,N_11589);
xor U14324 (N_14324,N_11018,N_9096);
nor U14325 (N_14325,N_9156,N_11708);
nor U14326 (N_14326,N_10897,N_11306);
nor U14327 (N_14327,N_10173,N_9757);
nand U14328 (N_14328,N_9851,N_10458);
and U14329 (N_14329,N_10161,N_9937);
nor U14330 (N_14330,N_11960,N_9714);
or U14331 (N_14331,N_11927,N_11820);
nand U14332 (N_14332,N_10485,N_9279);
or U14333 (N_14333,N_9883,N_11605);
nor U14334 (N_14334,N_11771,N_10408);
nor U14335 (N_14335,N_9367,N_9196);
nor U14336 (N_14336,N_9375,N_11914);
nand U14337 (N_14337,N_10413,N_9940);
nand U14338 (N_14338,N_11138,N_10635);
or U14339 (N_14339,N_10066,N_9524);
nor U14340 (N_14340,N_9224,N_9945);
nor U14341 (N_14341,N_11610,N_11537);
or U14342 (N_14342,N_9138,N_9006);
or U14343 (N_14343,N_9495,N_9865);
nor U14344 (N_14344,N_9814,N_10130);
nor U14345 (N_14345,N_10538,N_10873);
nand U14346 (N_14346,N_10560,N_11529);
or U14347 (N_14347,N_10187,N_11394);
nor U14348 (N_14348,N_10881,N_10243);
nand U14349 (N_14349,N_11359,N_9954);
nand U14350 (N_14350,N_11904,N_11886);
or U14351 (N_14351,N_11850,N_11006);
or U14352 (N_14352,N_9537,N_10741);
nand U14353 (N_14353,N_9756,N_11030);
nand U14354 (N_14354,N_10484,N_9994);
and U14355 (N_14355,N_9196,N_10417);
or U14356 (N_14356,N_10826,N_9502);
nand U14357 (N_14357,N_9093,N_9539);
and U14358 (N_14358,N_9170,N_9967);
nand U14359 (N_14359,N_10265,N_9330);
nor U14360 (N_14360,N_9253,N_11554);
and U14361 (N_14361,N_9969,N_9324);
nand U14362 (N_14362,N_9170,N_9234);
or U14363 (N_14363,N_10872,N_11446);
nor U14364 (N_14364,N_10470,N_10722);
nand U14365 (N_14365,N_10420,N_11578);
or U14366 (N_14366,N_9969,N_11961);
nand U14367 (N_14367,N_9296,N_9090);
nand U14368 (N_14368,N_9025,N_10311);
or U14369 (N_14369,N_11946,N_11479);
or U14370 (N_14370,N_10616,N_9022);
nand U14371 (N_14371,N_11013,N_10731);
nand U14372 (N_14372,N_9767,N_11165);
or U14373 (N_14373,N_11649,N_9900);
nor U14374 (N_14374,N_11298,N_10476);
nor U14375 (N_14375,N_9152,N_10715);
nor U14376 (N_14376,N_11278,N_11588);
or U14377 (N_14377,N_9310,N_10345);
nand U14378 (N_14378,N_10274,N_10959);
and U14379 (N_14379,N_11631,N_11388);
and U14380 (N_14380,N_10044,N_9282);
and U14381 (N_14381,N_10091,N_9748);
or U14382 (N_14382,N_10883,N_9142);
nor U14383 (N_14383,N_10352,N_9635);
and U14384 (N_14384,N_9800,N_10202);
nor U14385 (N_14385,N_11805,N_9964);
nand U14386 (N_14386,N_11095,N_10765);
and U14387 (N_14387,N_10357,N_9415);
or U14388 (N_14388,N_10901,N_11669);
nand U14389 (N_14389,N_10535,N_9291);
or U14390 (N_14390,N_11717,N_11058);
nand U14391 (N_14391,N_9897,N_11585);
and U14392 (N_14392,N_10685,N_10209);
nand U14393 (N_14393,N_9228,N_11808);
nand U14394 (N_14394,N_11723,N_10358);
nor U14395 (N_14395,N_9115,N_10285);
nor U14396 (N_14396,N_10991,N_11232);
nor U14397 (N_14397,N_9875,N_10980);
nor U14398 (N_14398,N_10966,N_11729);
nor U14399 (N_14399,N_9786,N_11733);
or U14400 (N_14400,N_9880,N_9547);
nand U14401 (N_14401,N_10996,N_10940);
and U14402 (N_14402,N_11478,N_9201);
nor U14403 (N_14403,N_9221,N_11085);
nand U14404 (N_14404,N_10103,N_9460);
nand U14405 (N_14405,N_10228,N_10358);
nor U14406 (N_14406,N_10688,N_10729);
and U14407 (N_14407,N_10596,N_10389);
and U14408 (N_14408,N_9934,N_10260);
and U14409 (N_14409,N_11291,N_11660);
and U14410 (N_14410,N_10905,N_11959);
nand U14411 (N_14411,N_9453,N_11644);
nand U14412 (N_14412,N_10871,N_9190);
or U14413 (N_14413,N_11545,N_10456);
nor U14414 (N_14414,N_11309,N_10272);
nor U14415 (N_14415,N_9052,N_9508);
or U14416 (N_14416,N_10021,N_9215);
nand U14417 (N_14417,N_10403,N_11377);
nor U14418 (N_14418,N_10832,N_9601);
or U14419 (N_14419,N_11227,N_10582);
nor U14420 (N_14420,N_11004,N_9611);
nand U14421 (N_14421,N_11407,N_10086);
nor U14422 (N_14422,N_11052,N_11695);
and U14423 (N_14423,N_11940,N_10484);
nand U14424 (N_14424,N_10275,N_9963);
and U14425 (N_14425,N_11925,N_10117);
nor U14426 (N_14426,N_10640,N_9495);
or U14427 (N_14427,N_9680,N_9840);
nor U14428 (N_14428,N_9443,N_10352);
nand U14429 (N_14429,N_10181,N_11943);
or U14430 (N_14430,N_9665,N_10551);
nand U14431 (N_14431,N_9760,N_9848);
xor U14432 (N_14432,N_10924,N_10655);
nor U14433 (N_14433,N_10798,N_9023);
nand U14434 (N_14434,N_9148,N_9407);
and U14435 (N_14435,N_9391,N_11422);
and U14436 (N_14436,N_9709,N_10340);
nand U14437 (N_14437,N_10991,N_10381);
nand U14438 (N_14438,N_10324,N_10686);
nor U14439 (N_14439,N_11841,N_11948);
xnor U14440 (N_14440,N_10605,N_9193);
nand U14441 (N_14441,N_11849,N_10684);
nand U14442 (N_14442,N_9352,N_10496);
or U14443 (N_14443,N_9472,N_9088);
and U14444 (N_14444,N_11377,N_11667);
and U14445 (N_14445,N_10594,N_9147);
nor U14446 (N_14446,N_10275,N_11825);
and U14447 (N_14447,N_9145,N_11652);
nand U14448 (N_14448,N_9403,N_9408);
or U14449 (N_14449,N_11134,N_11489);
and U14450 (N_14450,N_9078,N_11590);
nor U14451 (N_14451,N_10718,N_9934);
nand U14452 (N_14452,N_11801,N_10184);
and U14453 (N_14453,N_10747,N_10848);
nor U14454 (N_14454,N_9266,N_10313);
and U14455 (N_14455,N_10167,N_10893);
nor U14456 (N_14456,N_10742,N_10384);
nand U14457 (N_14457,N_10606,N_10565);
or U14458 (N_14458,N_10927,N_11285);
nand U14459 (N_14459,N_10803,N_9395);
nor U14460 (N_14460,N_10562,N_9038);
nor U14461 (N_14461,N_10358,N_10283);
nor U14462 (N_14462,N_10904,N_11584);
nand U14463 (N_14463,N_11289,N_9478);
nand U14464 (N_14464,N_9318,N_11969);
nor U14465 (N_14465,N_11255,N_10899);
or U14466 (N_14466,N_11636,N_9163);
or U14467 (N_14467,N_11674,N_10857);
nor U14468 (N_14468,N_10381,N_11488);
nor U14469 (N_14469,N_10268,N_10971);
and U14470 (N_14470,N_9805,N_10760);
and U14471 (N_14471,N_9614,N_10290);
and U14472 (N_14472,N_11449,N_9738);
or U14473 (N_14473,N_9934,N_11481);
xor U14474 (N_14474,N_10231,N_9540);
nand U14475 (N_14475,N_9468,N_10560);
or U14476 (N_14476,N_9167,N_11552);
or U14477 (N_14477,N_11387,N_11480);
nand U14478 (N_14478,N_11667,N_11806);
nor U14479 (N_14479,N_11563,N_11968);
nand U14480 (N_14480,N_9919,N_10158);
and U14481 (N_14481,N_11614,N_11515);
or U14482 (N_14482,N_11919,N_10064);
nand U14483 (N_14483,N_9011,N_10931);
nand U14484 (N_14484,N_9525,N_11248);
nor U14485 (N_14485,N_10370,N_9338);
or U14486 (N_14486,N_10732,N_9019);
or U14487 (N_14487,N_10686,N_10365);
nor U14488 (N_14488,N_10067,N_11341);
nand U14489 (N_14489,N_11518,N_11328);
nand U14490 (N_14490,N_10611,N_9025);
nand U14491 (N_14491,N_9040,N_9749);
and U14492 (N_14492,N_10787,N_10370);
or U14493 (N_14493,N_10569,N_11921);
nor U14494 (N_14494,N_11635,N_11354);
and U14495 (N_14495,N_10837,N_10776);
nand U14496 (N_14496,N_10941,N_11073);
nor U14497 (N_14497,N_10527,N_11763);
nor U14498 (N_14498,N_10895,N_11859);
nand U14499 (N_14499,N_10309,N_9607);
nand U14500 (N_14500,N_11984,N_10333);
or U14501 (N_14501,N_10005,N_9552);
nand U14502 (N_14502,N_10675,N_9393);
nor U14503 (N_14503,N_11788,N_10758);
nand U14504 (N_14504,N_11147,N_10375);
nor U14505 (N_14505,N_9513,N_11612);
or U14506 (N_14506,N_10352,N_11655);
or U14507 (N_14507,N_11030,N_10033);
and U14508 (N_14508,N_11485,N_11997);
nand U14509 (N_14509,N_9999,N_9486);
or U14510 (N_14510,N_9532,N_9974);
nor U14511 (N_14511,N_9181,N_11687);
or U14512 (N_14512,N_10680,N_10251);
or U14513 (N_14513,N_9648,N_9677);
nor U14514 (N_14514,N_11805,N_11638);
nor U14515 (N_14515,N_11545,N_11015);
or U14516 (N_14516,N_11283,N_11119);
and U14517 (N_14517,N_10704,N_9541);
nor U14518 (N_14518,N_10743,N_10096);
nor U14519 (N_14519,N_11906,N_11777);
or U14520 (N_14520,N_11776,N_10721);
nand U14521 (N_14521,N_10106,N_10747);
nor U14522 (N_14522,N_9916,N_10095);
xor U14523 (N_14523,N_9598,N_11868);
or U14524 (N_14524,N_11389,N_10805);
and U14525 (N_14525,N_9897,N_9573);
or U14526 (N_14526,N_11738,N_9558);
or U14527 (N_14527,N_10502,N_9687);
nand U14528 (N_14528,N_11266,N_10623);
nand U14529 (N_14529,N_9836,N_11264);
or U14530 (N_14530,N_10345,N_11783);
and U14531 (N_14531,N_9656,N_10645);
and U14532 (N_14532,N_10022,N_10165);
nor U14533 (N_14533,N_9283,N_11455);
nor U14534 (N_14534,N_11862,N_11436);
or U14535 (N_14535,N_11535,N_10801);
nor U14536 (N_14536,N_11555,N_11664);
nor U14537 (N_14537,N_9380,N_10014);
nor U14538 (N_14538,N_11432,N_9235);
nand U14539 (N_14539,N_9825,N_10192);
nor U14540 (N_14540,N_11765,N_10336);
nor U14541 (N_14541,N_11431,N_9295);
or U14542 (N_14542,N_11981,N_10703);
or U14543 (N_14543,N_11006,N_9249);
and U14544 (N_14544,N_11910,N_11131);
nand U14545 (N_14545,N_10023,N_11580);
and U14546 (N_14546,N_11228,N_9997);
and U14547 (N_14547,N_9451,N_9401);
nand U14548 (N_14548,N_11830,N_9740);
nor U14549 (N_14549,N_9140,N_10951);
or U14550 (N_14550,N_11634,N_9214);
nor U14551 (N_14551,N_10556,N_10634);
nor U14552 (N_14552,N_10870,N_9361);
and U14553 (N_14553,N_11540,N_9574);
or U14554 (N_14554,N_9745,N_10666);
and U14555 (N_14555,N_9133,N_9078);
nor U14556 (N_14556,N_10195,N_10998);
and U14557 (N_14557,N_9707,N_10113);
or U14558 (N_14558,N_11796,N_9368);
and U14559 (N_14559,N_9717,N_11618);
or U14560 (N_14560,N_9786,N_9262);
nor U14561 (N_14561,N_9038,N_11479);
or U14562 (N_14562,N_10742,N_10017);
nand U14563 (N_14563,N_10618,N_11436);
and U14564 (N_14564,N_10045,N_11859);
or U14565 (N_14565,N_10040,N_9669);
nor U14566 (N_14566,N_9901,N_11361);
nand U14567 (N_14567,N_10116,N_9939);
and U14568 (N_14568,N_10927,N_9950);
or U14569 (N_14569,N_10103,N_10116);
and U14570 (N_14570,N_11885,N_11567);
and U14571 (N_14571,N_10000,N_9423);
nand U14572 (N_14572,N_10821,N_11606);
and U14573 (N_14573,N_9612,N_9062);
nand U14574 (N_14574,N_10655,N_10221);
and U14575 (N_14575,N_11388,N_11536);
or U14576 (N_14576,N_11023,N_10969);
nor U14577 (N_14577,N_11841,N_11707);
and U14578 (N_14578,N_10590,N_11815);
and U14579 (N_14579,N_9944,N_11870);
nand U14580 (N_14580,N_9580,N_9698);
nand U14581 (N_14581,N_9376,N_10760);
and U14582 (N_14582,N_9400,N_9165);
nor U14583 (N_14583,N_11991,N_9581);
nand U14584 (N_14584,N_11724,N_10679);
or U14585 (N_14585,N_9155,N_9047);
and U14586 (N_14586,N_9156,N_9926);
nor U14587 (N_14587,N_9745,N_11612);
nor U14588 (N_14588,N_9996,N_9209);
or U14589 (N_14589,N_9335,N_9543);
or U14590 (N_14590,N_11918,N_10483);
and U14591 (N_14591,N_10211,N_9289);
or U14592 (N_14592,N_10048,N_10420);
or U14593 (N_14593,N_11578,N_11025);
or U14594 (N_14594,N_11594,N_10748);
or U14595 (N_14595,N_10412,N_9819);
and U14596 (N_14596,N_9722,N_11971);
or U14597 (N_14597,N_9063,N_11547);
and U14598 (N_14598,N_10265,N_11396);
or U14599 (N_14599,N_10824,N_11500);
nand U14600 (N_14600,N_11408,N_11560);
or U14601 (N_14601,N_10898,N_11826);
nor U14602 (N_14602,N_11188,N_11306);
and U14603 (N_14603,N_11023,N_9975);
or U14604 (N_14604,N_11926,N_11404);
and U14605 (N_14605,N_11726,N_9469);
nand U14606 (N_14606,N_9642,N_9407);
and U14607 (N_14607,N_10585,N_11431);
or U14608 (N_14608,N_10681,N_9757);
nand U14609 (N_14609,N_10241,N_11384);
or U14610 (N_14610,N_9098,N_11142);
nor U14611 (N_14611,N_10639,N_11250);
or U14612 (N_14612,N_11704,N_10392);
nor U14613 (N_14613,N_9036,N_9937);
nor U14614 (N_14614,N_11365,N_11390);
nor U14615 (N_14615,N_10611,N_10901);
nand U14616 (N_14616,N_10168,N_9660);
nor U14617 (N_14617,N_11947,N_11166);
and U14618 (N_14618,N_9912,N_9337);
xor U14619 (N_14619,N_11314,N_9892);
nor U14620 (N_14620,N_10325,N_11500);
nor U14621 (N_14621,N_10280,N_11955);
nand U14622 (N_14622,N_10171,N_10691);
nor U14623 (N_14623,N_11391,N_11176);
nor U14624 (N_14624,N_10805,N_11532);
and U14625 (N_14625,N_11879,N_10974);
nand U14626 (N_14626,N_11124,N_10634);
nand U14627 (N_14627,N_10195,N_9698);
nand U14628 (N_14628,N_11061,N_10163);
nand U14629 (N_14629,N_9511,N_10926);
or U14630 (N_14630,N_10770,N_9931);
nor U14631 (N_14631,N_11842,N_9048);
nand U14632 (N_14632,N_10852,N_11066);
nand U14633 (N_14633,N_9102,N_9138);
and U14634 (N_14634,N_9560,N_11692);
or U14635 (N_14635,N_9385,N_9721);
nor U14636 (N_14636,N_10605,N_10032);
and U14637 (N_14637,N_10565,N_10566);
nor U14638 (N_14638,N_10513,N_9753);
and U14639 (N_14639,N_10699,N_11973);
or U14640 (N_14640,N_9016,N_10262);
nor U14641 (N_14641,N_11492,N_9508);
or U14642 (N_14642,N_11532,N_11381);
nand U14643 (N_14643,N_9640,N_9268);
and U14644 (N_14644,N_10398,N_11543);
or U14645 (N_14645,N_9709,N_9034);
nand U14646 (N_14646,N_9877,N_11966);
nand U14647 (N_14647,N_10861,N_11784);
and U14648 (N_14648,N_11302,N_9497);
or U14649 (N_14649,N_9703,N_9609);
nor U14650 (N_14650,N_11355,N_10583);
or U14651 (N_14651,N_9267,N_9145);
nand U14652 (N_14652,N_9021,N_9938);
nand U14653 (N_14653,N_9649,N_11811);
and U14654 (N_14654,N_11347,N_11962);
or U14655 (N_14655,N_9313,N_11388);
nor U14656 (N_14656,N_9113,N_9070);
nor U14657 (N_14657,N_9521,N_11390);
and U14658 (N_14658,N_10197,N_9333);
xnor U14659 (N_14659,N_10657,N_9769);
and U14660 (N_14660,N_11265,N_10528);
nand U14661 (N_14661,N_11509,N_11492);
nor U14662 (N_14662,N_9493,N_11142);
nor U14663 (N_14663,N_9672,N_9022);
nor U14664 (N_14664,N_9410,N_11366);
nand U14665 (N_14665,N_10119,N_10331);
nand U14666 (N_14666,N_11381,N_10013);
or U14667 (N_14667,N_11373,N_9688);
nand U14668 (N_14668,N_11458,N_9678);
and U14669 (N_14669,N_10756,N_11207);
nand U14670 (N_14670,N_11358,N_9426);
nor U14671 (N_14671,N_11866,N_9183);
and U14672 (N_14672,N_11771,N_11893);
nand U14673 (N_14673,N_9087,N_9147);
nor U14674 (N_14674,N_10032,N_11386);
or U14675 (N_14675,N_10704,N_10062);
or U14676 (N_14676,N_10254,N_10712);
nor U14677 (N_14677,N_11998,N_9632);
nor U14678 (N_14678,N_11372,N_9341);
nand U14679 (N_14679,N_10280,N_10267);
and U14680 (N_14680,N_9279,N_9228);
nor U14681 (N_14681,N_10597,N_9941);
or U14682 (N_14682,N_9072,N_10517);
nand U14683 (N_14683,N_11373,N_11520);
and U14684 (N_14684,N_9538,N_10206);
nor U14685 (N_14685,N_10507,N_11723);
nand U14686 (N_14686,N_11743,N_10500);
nor U14687 (N_14687,N_10697,N_10585);
or U14688 (N_14688,N_9641,N_11116);
nand U14689 (N_14689,N_11993,N_10749);
nand U14690 (N_14690,N_9697,N_9022);
and U14691 (N_14691,N_9772,N_9607);
nor U14692 (N_14692,N_10896,N_11699);
and U14693 (N_14693,N_11435,N_11093);
nand U14694 (N_14694,N_11745,N_9599);
nand U14695 (N_14695,N_9298,N_11716);
nand U14696 (N_14696,N_10298,N_9132);
nand U14697 (N_14697,N_10575,N_9992);
and U14698 (N_14698,N_10546,N_9222);
or U14699 (N_14699,N_9564,N_9553);
nand U14700 (N_14700,N_11479,N_10530);
nor U14701 (N_14701,N_11445,N_11381);
and U14702 (N_14702,N_11257,N_11571);
nor U14703 (N_14703,N_9157,N_11212);
nand U14704 (N_14704,N_10575,N_11988);
and U14705 (N_14705,N_10943,N_9020);
nor U14706 (N_14706,N_9552,N_10109);
nor U14707 (N_14707,N_10524,N_11050);
or U14708 (N_14708,N_11812,N_9706);
nand U14709 (N_14709,N_10663,N_9252);
nand U14710 (N_14710,N_10181,N_10089);
and U14711 (N_14711,N_10195,N_9190);
or U14712 (N_14712,N_11831,N_10861);
nor U14713 (N_14713,N_10785,N_10184);
nand U14714 (N_14714,N_11568,N_10683);
or U14715 (N_14715,N_9651,N_11626);
nand U14716 (N_14716,N_11523,N_9095);
nand U14717 (N_14717,N_9981,N_10470);
xor U14718 (N_14718,N_10345,N_11524);
nand U14719 (N_14719,N_11925,N_9123);
nor U14720 (N_14720,N_9594,N_11095);
xor U14721 (N_14721,N_9326,N_10380);
and U14722 (N_14722,N_11379,N_9880);
nand U14723 (N_14723,N_9676,N_11499);
xor U14724 (N_14724,N_10652,N_9132);
or U14725 (N_14725,N_9569,N_11129);
nand U14726 (N_14726,N_10253,N_10640);
and U14727 (N_14727,N_11693,N_9736);
and U14728 (N_14728,N_11154,N_9727);
nand U14729 (N_14729,N_10030,N_10716);
and U14730 (N_14730,N_10099,N_11237);
and U14731 (N_14731,N_9994,N_9347);
or U14732 (N_14732,N_10376,N_10518);
and U14733 (N_14733,N_10567,N_10535);
and U14734 (N_14734,N_11396,N_10373);
nand U14735 (N_14735,N_11735,N_9165);
or U14736 (N_14736,N_10434,N_9422);
and U14737 (N_14737,N_9822,N_11761);
nor U14738 (N_14738,N_11817,N_11534);
xnor U14739 (N_14739,N_9181,N_10543);
and U14740 (N_14740,N_10628,N_11841);
nand U14741 (N_14741,N_11786,N_11402);
and U14742 (N_14742,N_11384,N_9163);
and U14743 (N_14743,N_9377,N_9833);
nor U14744 (N_14744,N_10491,N_11919);
nor U14745 (N_14745,N_9294,N_10179);
nor U14746 (N_14746,N_11460,N_9387);
or U14747 (N_14747,N_11055,N_9767);
nand U14748 (N_14748,N_11197,N_10007);
or U14749 (N_14749,N_10726,N_11094);
nand U14750 (N_14750,N_11220,N_9726);
and U14751 (N_14751,N_11876,N_9300);
nor U14752 (N_14752,N_9720,N_11470);
and U14753 (N_14753,N_10179,N_11561);
and U14754 (N_14754,N_10011,N_11068);
nor U14755 (N_14755,N_10860,N_10990);
nand U14756 (N_14756,N_10879,N_10530);
or U14757 (N_14757,N_11902,N_11506);
and U14758 (N_14758,N_10910,N_10226);
nand U14759 (N_14759,N_11053,N_10019);
and U14760 (N_14760,N_9577,N_10713);
and U14761 (N_14761,N_11698,N_9499);
nand U14762 (N_14762,N_10402,N_10852);
or U14763 (N_14763,N_9110,N_10101);
nand U14764 (N_14764,N_10104,N_9570);
nor U14765 (N_14765,N_11292,N_9289);
or U14766 (N_14766,N_11374,N_9409);
and U14767 (N_14767,N_9081,N_10636);
nand U14768 (N_14768,N_10935,N_11278);
or U14769 (N_14769,N_10684,N_11003);
or U14770 (N_14770,N_10861,N_11155);
and U14771 (N_14771,N_9175,N_11844);
and U14772 (N_14772,N_11994,N_11376);
nor U14773 (N_14773,N_11996,N_9917);
or U14774 (N_14774,N_11587,N_11636);
or U14775 (N_14775,N_10323,N_10943);
nor U14776 (N_14776,N_11354,N_10517);
or U14777 (N_14777,N_11883,N_11132);
nand U14778 (N_14778,N_10203,N_10740);
or U14779 (N_14779,N_9337,N_9850);
nor U14780 (N_14780,N_11478,N_10611);
nand U14781 (N_14781,N_9985,N_10124);
or U14782 (N_14782,N_11451,N_9923);
nand U14783 (N_14783,N_10174,N_10703);
nand U14784 (N_14784,N_10206,N_9214);
nand U14785 (N_14785,N_9132,N_10782);
nor U14786 (N_14786,N_9644,N_11483);
and U14787 (N_14787,N_11267,N_9967);
and U14788 (N_14788,N_11453,N_9327);
nand U14789 (N_14789,N_11310,N_9795);
and U14790 (N_14790,N_10931,N_10727);
or U14791 (N_14791,N_11506,N_9287);
or U14792 (N_14792,N_10163,N_9188);
nand U14793 (N_14793,N_11711,N_10161);
and U14794 (N_14794,N_10698,N_9314);
nand U14795 (N_14795,N_11630,N_11888);
nand U14796 (N_14796,N_9483,N_11891);
nand U14797 (N_14797,N_11514,N_11551);
nand U14798 (N_14798,N_10943,N_11579);
nand U14799 (N_14799,N_10399,N_10415);
nand U14800 (N_14800,N_11329,N_10419);
or U14801 (N_14801,N_9587,N_11015);
nor U14802 (N_14802,N_9449,N_9980);
nor U14803 (N_14803,N_11391,N_11926);
nor U14804 (N_14804,N_10798,N_10830);
nor U14805 (N_14805,N_10764,N_11193);
nor U14806 (N_14806,N_10258,N_10637);
nor U14807 (N_14807,N_11426,N_11624);
nor U14808 (N_14808,N_9800,N_9050);
nand U14809 (N_14809,N_10931,N_10971);
and U14810 (N_14810,N_10746,N_10476);
and U14811 (N_14811,N_9508,N_10056);
nand U14812 (N_14812,N_10728,N_10181);
and U14813 (N_14813,N_10545,N_10148);
nor U14814 (N_14814,N_11804,N_11228);
or U14815 (N_14815,N_10546,N_9877);
nand U14816 (N_14816,N_11994,N_10039);
and U14817 (N_14817,N_10149,N_9007);
nor U14818 (N_14818,N_11267,N_9195);
nor U14819 (N_14819,N_9184,N_10629);
xnor U14820 (N_14820,N_11365,N_10598);
nand U14821 (N_14821,N_11604,N_9201);
nand U14822 (N_14822,N_10504,N_11958);
or U14823 (N_14823,N_9043,N_9783);
nand U14824 (N_14824,N_9236,N_9793);
xnor U14825 (N_14825,N_11239,N_10042);
or U14826 (N_14826,N_9761,N_10913);
nand U14827 (N_14827,N_10714,N_9817);
or U14828 (N_14828,N_10713,N_11903);
nand U14829 (N_14829,N_11843,N_11196);
nor U14830 (N_14830,N_11603,N_11054);
nand U14831 (N_14831,N_9149,N_11325);
nand U14832 (N_14832,N_11112,N_10041);
and U14833 (N_14833,N_10438,N_10073);
or U14834 (N_14834,N_9115,N_11922);
or U14835 (N_14835,N_11103,N_11088);
and U14836 (N_14836,N_10294,N_10594);
nor U14837 (N_14837,N_9992,N_9063);
and U14838 (N_14838,N_9380,N_11159);
and U14839 (N_14839,N_10094,N_11034);
nand U14840 (N_14840,N_10787,N_11697);
and U14841 (N_14841,N_10981,N_9526);
nor U14842 (N_14842,N_9725,N_11639);
and U14843 (N_14843,N_11894,N_10238);
or U14844 (N_14844,N_9218,N_10472);
or U14845 (N_14845,N_9194,N_10640);
nand U14846 (N_14846,N_10761,N_11615);
or U14847 (N_14847,N_10293,N_9071);
or U14848 (N_14848,N_11465,N_11716);
nor U14849 (N_14849,N_9194,N_11718);
or U14850 (N_14850,N_10400,N_11267);
and U14851 (N_14851,N_11313,N_10075);
nand U14852 (N_14852,N_9078,N_11125);
nand U14853 (N_14853,N_11772,N_10883);
nor U14854 (N_14854,N_9360,N_10694);
or U14855 (N_14855,N_9314,N_9707);
nand U14856 (N_14856,N_9236,N_9518);
and U14857 (N_14857,N_11158,N_11879);
and U14858 (N_14858,N_9347,N_10274);
and U14859 (N_14859,N_11392,N_11626);
or U14860 (N_14860,N_10038,N_10898);
or U14861 (N_14861,N_11615,N_9643);
nor U14862 (N_14862,N_9281,N_10451);
nand U14863 (N_14863,N_10449,N_11189);
and U14864 (N_14864,N_9955,N_11159);
nand U14865 (N_14865,N_11982,N_10065);
nand U14866 (N_14866,N_11611,N_10855);
nor U14867 (N_14867,N_9017,N_9841);
or U14868 (N_14868,N_11380,N_11263);
and U14869 (N_14869,N_11052,N_11820);
and U14870 (N_14870,N_11581,N_9424);
or U14871 (N_14871,N_9922,N_11512);
and U14872 (N_14872,N_9955,N_9162);
nand U14873 (N_14873,N_11587,N_11442);
and U14874 (N_14874,N_10767,N_10470);
and U14875 (N_14875,N_11065,N_11652);
nand U14876 (N_14876,N_11457,N_11797);
nand U14877 (N_14877,N_10534,N_9441);
nor U14878 (N_14878,N_11374,N_11433);
or U14879 (N_14879,N_9546,N_10814);
nor U14880 (N_14880,N_9495,N_10663);
nand U14881 (N_14881,N_11153,N_9049);
nor U14882 (N_14882,N_10846,N_9916);
nand U14883 (N_14883,N_10302,N_11916);
nand U14884 (N_14884,N_11160,N_11982);
nor U14885 (N_14885,N_10934,N_9893);
and U14886 (N_14886,N_10563,N_10395);
and U14887 (N_14887,N_10763,N_11635);
nor U14888 (N_14888,N_9586,N_11178);
nor U14889 (N_14889,N_11197,N_10809);
and U14890 (N_14890,N_11512,N_9885);
nand U14891 (N_14891,N_9991,N_10237);
and U14892 (N_14892,N_9836,N_9252);
or U14893 (N_14893,N_9917,N_10965);
or U14894 (N_14894,N_11114,N_10104);
nor U14895 (N_14895,N_11167,N_9461);
or U14896 (N_14896,N_11587,N_11444);
and U14897 (N_14897,N_9422,N_10343);
and U14898 (N_14898,N_10967,N_10798);
or U14899 (N_14899,N_9676,N_11683);
and U14900 (N_14900,N_11772,N_9860);
nand U14901 (N_14901,N_10702,N_9550);
nand U14902 (N_14902,N_11986,N_9981);
nand U14903 (N_14903,N_9949,N_10843);
or U14904 (N_14904,N_10557,N_10790);
nor U14905 (N_14905,N_10547,N_10052);
nand U14906 (N_14906,N_11724,N_10309);
or U14907 (N_14907,N_11021,N_11346);
nor U14908 (N_14908,N_9841,N_9969);
and U14909 (N_14909,N_9133,N_11068);
or U14910 (N_14910,N_11029,N_11232);
nand U14911 (N_14911,N_9973,N_10005);
or U14912 (N_14912,N_10447,N_11468);
and U14913 (N_14913,N_10385,N_9626);
or U14914 (N_14914,N_9536,N_10815);
and U14915 (N_14915,N_10388,N_10521);
and U14916 (N_14916,N_9945,N_11049);
or U14917 (N_14917,N_10325,N_9325);
and U14918 (N_14918,N_10472,N_9237);
nand U14919 (N_14919,N_11365,N_10874);
and U14920 (N_14920,N_11277,N_11595);
nand U14921 (N_14921,N_11049,N_10734);
and U14922 (N_14922,N_11826,N_9442);
nor U14923 (N_14923,N_9061,N_11891);
nand U14924 (N_14924,N_9700,N_11170);
nor U14925 (N_14925,N_9877,N_10752);
nand U14926 (N_14926,N_10264,N_9815);
or U14927 (N_14927,N_11999,N_10824);
nand U14928 (N_14928,N_9071,N_11896);
or U14929 (N_14929,N_11727,N_9678);
nand U14930 (N_14930,N_9860,N_10180);
nand U14931 (N_14931,N_11094,N_9455);
and U14932 (N_14932,N_9423,N_9921);
or U14933 (N_14933,N_10707,N_10027);
nand U14934 (N_14934,N_10078,N_11690);
xor U14935 (N_14935,N_10556,N_10443);
nand U14936 (N_14936,N_10154,N_9110);
or U14937 (N_14937,N_9246,N_11092);
and U14938 (N_14938,N_10631,N_11788);
or U14939 (N_14939,N_9478,N_9278);
or U14940 (N_14940,N_9997,N_11622);
xnor U14941 (N_14941,N_11759,N_11791);
and U14942 (N_14942,N_11295,N_9947);
nand U14943 (N_14943,N_11115,N_11613);
nor U14944 (N_14944,N_9256,N_11946);
or U14945 (N_14945,N_11697,N_10207);
or U14946 (N_14946,N_10108,N_11104);
nor U14947 (N_14947,N_11401,N_11955);
nor U14948 (N_14948,N_10708,N_11948);
nor U14949 (N_14949,N_11902,N_10092);
nor U14950 (N_14950,N_10897,N_11283);
and U14951 (N_14951,N_11557,N_9835);
nor U14952 (N_14952,N_10039,N_9134);
and U14953 (N_14953,N_10954,N_11460);
nor U14954 (N_14954,N_9794,N_11103);
nand U14955 (N_14955,N_10751,N_11893);
nand U14956 (N_14956,N_10257,N_11061);
or U14957 (N_14957,N_10357,N_11916);
and U14958 (N_14958,N_10206,N_9768);
nand U14959 (N_14959,N_11272,N_11776);
or U14960 (N_14960,N_9636,N_9899);
nand U14961 (N_14961,N_11708,N_11687);
nand U14962 (N_14962,N_10818,N_11679);
or U14963 (N_14963,N_9633,N_10783);
nor U14964 (N_14964,N_11524,N_10642);
and U14965 (N_14965,N_11203,N_9493);
and U14966 (N_14966,N_11861,N_9018);
and U14967 (N_14967,N_10122,N_10803);
nor U14968 (N_14968,N_11992,N_10438);
xor U14969 (N_14969,N_11393,N_10120);
nor U14970 (N_14970,N_9989,N_10166);
nor U14971 (N_14971,N_9457,N_10851);
and U14972 (N_14972,N_10532,N_10581);
and U14973 (N_14973,N_9258,N_9149);
nand U14974 (N_14974,N_10321,N_11845);
nand U14975 (N_14975,N_11551,N_10639);
nand U14976 (N_14976,N_10757,N_10943);
nor U14977 (N_14977,N_10949,N_9487);
nand U14978 (N_14978,N_10547,N_10930);
nor U14979 (N_14979,N_10021,N_11612);
or U14980 (N_14980,N_10574,N_11173);
or U14981 (N_14981,N_11229,N_10078);
xnor U14982 (N_14982,N_10924,N_11628);
and U14983 (N_14983,N_10458,N_9386);
or U14984 (N_14984,N_9762,N_10690);
or U14985 (N_14985,N_11211,N_9646);
and U14986 (N_14986,N_9461,N_11400);
nand U14987 (N_14987,N_10846,N_10166);
and U14988 (N_14988,N_10184,N_11514);
nand U14989 (N_14989,N_9454,N_9078);
nor U14990 (N_14990,N_9457,N_9594);
nor U14991 (N_14991,N_11902,N_9143);
or U14992 (N_14992,N_10768,N_10617);
and U14993 (N_14993,N_10282,N_11495);
and U14994 (N_14994,N_10853,N_11919);
nor U14995 (N_14995,N_10955,N_10743);
nand U14996 (N_14996,N_9018,N_10555);
and U14997 (N_14997,N_9749,N_11770);
and U14998 (N_14998,N_11955,N_11087);
and U14999 (N_14999,N_9228,N_11475);
or UO_0 (O_0,N_13015,N_14582);
nand UO_1 (O_1,N_13816,N_13175);
nand UO_2 (O_2,N_12518,N_14001);
or UO_3 (O_3,N_12483,N_12876);
nand UO_4 (O_4,N_14086,N_12355);
or UO_5 (O_5,N_14743,N_13277);
and UO_6 (O_6,N_13516,N_12607);
and UO_7 (O_7,N_12115,N_14571);
nand UO_8 (O_8,N_12639,N_13972);
nor UO_9 (O_9,N_14251,N_13592);
nor UO_10 (O_10,N_13691,N_14772);
nand UO_11 (O_11,N_13683,N_13621);
nand UO_12 (O_12,N_12753,N_12660);
and UO_13 (O_13,N_14368,N_14801);
and UO_14 (O_14,N_14745,N_12523);
or UO_15 (O_15,N_14581,N_12279);
or UO_16 (O_16,N_14053,N_13835);
and UO_17 (O_17,N_13682,N_12870);
nor UO_18 (O_18,N_14204,N_13399);
nand UO_19 (O_19,N_14671,N_13292);
nand UO_20 (O_20,N_12982,N_13892);
or UO_21 (O_21,N_14019,N_14353);
and UO_22 (O_22,N_14245,N_12033);
nand UO_23 (O_23,N_13149,N_12055);
nand UO_24 (O_24,N_12987,N_12846);
and UO_25 (O_25,N_13792,N_12818);
or UO_26 (O_26,N_13671,N_14359);
nand UO_27 (O_27,N_12413,N_14736);
or UO_28 (O_28,N_14799,N_12510);
nor UO_29 (O_29,N_12521,N_12685);
or UO_30 (O_30,N_13071,N_12623);
nand UO_31 (O_31,N_12371,N_14696);
nor UO_32 (O_32,N_13849,N_14826);
and UO_33 (O_33,N_13384,N_12156);
nor UO_34 (O_34,N_13958,N_12648);
nand UO_35 (O_35,N_14460,N_12610);
or UO_36 (O_36,N_13694,N_14013);
nand UO_37 (O_37,N_14670,N_12694);
nor UO_38 (O_38,N_12630,N_13341);
or UO_39 (O_39,N_14827,N_14751);
and UO_40 (O_40,N_14485,N_12095);
and UO_41 (O_41,N_13717,N_13209);
or UO_42 (O_42,N_13834,N_13395);
or UO_43 (O_43,N_12389,N_14823);
nor UO_44 (O_44,N_13097,N_14265);
and UO_45 (O_45,N_12892,N_14284);
nand UO_46 (O_46,N_12498,N_14159);
and UO_47 (O_47,N_13154,N_13383);
or UO_48 (O_48,N_13301,N_12627);
and UO_49 (O_49,N_12801,N_14014);
nor UO_50 (O_50,N_14203,N_13882);
nor UO_51 (O_51,N_14200,N_14329);
nor UO_52 (O_52,N_12200,N_14002);
nor UO_53 (O_53,N_14243,N_14221);
nand UO_54 (O_54,N_14762,N_14010);
nor UO_55 (O_55,N_14781,N_14474);
or UO_56 (O_56,N_12333,N_13722);
xnor UO_57 (O_57,N_12345,N_14062);
nand UO_58 (O_58,N_14985,N_12142);
nand UO_59 (O_59,N_14720,N_14958);
and UO_60 (O_60,N_12046,N_12716);
or UO_61 (O_61,N_13618,N_12168);
and UO_62 (O_62,N_12029,N_14675);
nand UO_63 (O_63,N_14924,N_12939);
nand UO_64 (O_64,N_14310,N_14396);
and UO_65 (O_65,N_14803,N_12524);
and UO_66 (O_66,N_13076,N_14822);
nor UO_67 (O_67,N_13377,N_14316);
or UO_68 (O_68,N_14000,N_14810);
nor UO_69 (O_69,N_13006,N_13656);
or UO_70 (O_70,N_13710,N_13438);
nor UO_71 (O_71,N_14256,N_14066);
or UO_72 (O_72,N_12953,N_12497);
or UO_73 (O_73,N_13235,N_12847);
and UO_74 (O_74,N_14367,N_13821);
nand UO_75 (O_75,N_14680,N_13714);
nor UO_76 (O_76,N_12773,N_13126);
or UO_77 (O_77,N_12440,N_13141);
and UO_78 (O_78,N_14858,N_14550);
or UO_79 (O_79,N_12999,N_13159);
nor UO_80 (O_80,N_14632,N_13106);
and UO_81 (O_81,N_12605,N_14651);
nand UO_82 (O_82,N_12832,N_12360);
nand UO_83 (O_83,N_14297,N_13761);
or UO_84 (O_84,N_14580,N_13394);
and UO_85 (O_85,N_14514,N_13789);
or UO_86 (O_86,N_12039,N_13840);
xor UO_87 (O_87,N_14301,N_13225);
and UO_88 (O_88,N_14929,N_12077);
or UO_89 (O_89,N_14820,N_12951);
and UO_90 (O_90,N_12928,N_12148);
and UO_91 (O_91,N_14987,N_12004);
and UO_92 (O_92,N_12394,N_13854);
and UO_93 (O_93,N_13819,N_13900);
nor UO_94 (O_94,N_13619,N_13393);
nor UO_95 (O_95,N_14092,N_14541);
and UO_96 (O_96,N_12188,N_14427);
or UO_97 (O_97,N_14175,N_12793);
or UO_98 (O_98,N_14458,N_14702);
and UO_99 (O_99,N_12068,N_14350);
and UO_100 (O_100,N_13625,N_12711);
nand UO_101 (O_101,N_13757,N_12744);
or UO_102 (O_102,N_14241,N_13226);
and UO_103 (O_103,N_14047,N_14084);
and UO_104 (O_104,N_14538,N_14943);
nor UO_105 (O_105,N_13309,N_13897);
and UO_106 (O_106,N_14761,N_14527);
nor UO_107 (O_107,N_12448,N_14999);
and UO_108 (O_108,N_14871,N_13950);
or UO_109 (O_109,N_12151,N_14641);
or UO_110 (O_110,N_13044,N_12451);
nand UO_111 (O_111,N_13969,N_14373);
or UO_112 (O_112,N_14846,N_12896);
nor UO_113 (O_113,N_13372,N_12768);
or UO_114 (O_114,N_14774,N_12102);
nor UO_115 (O_115,N_14492,N_12652);
and UO_116 (O_116,N_13063,N_12804);
and UO_117 (O_117,N_12949,N_12233);
nor UO_118 (O_118,N_12320,N_14399);
nand UO_119 (O_119,N_12754,N_12766);
nor UO_120 (O_120,N_12615,N_13780);
and UO_121 (O_121,N_12180,N_12828);
and UO_122 (O_122,N_12748,N_14837);
nand UO_123 (O_123,N_12676,N_12376);
nand UO_124 (O_124,N_12977,N_13408);
or UO_125 (O_125,N_14394,N_13296);
nand UO_126 (O_126,N_13725,N_13743);
and UO_127 (O_127,N_14590,N_12911);
nor UO_128 (O_128,N_14383,N_13651);
or UO_129 (O_129,N_13986,N_12344);
nand UO_130 (O_130,N_14401,N_13025);
nand UO_131 (O_131,N_13822,N_13387);
nor UO_132 (O_132,N_13544,N_14444);
or UO_133 (O_133,N_14973,N_14191);
and UO_134 (O_134,N_13566,N_13429);
nor UO_135 (O_135,N_14619,N_13089);
nand UO_136 (O_136,N_14638,N_14272);
or UO_137 (O_137,N_14737,N_12374);
nand UO_138 (O_138,N_13528,N_12408);
xnor UO_139 (O_139,N_12733,N_12259);
nand UO_140 (O_140,N_12063,N_13338);
nand UO_141 (O_141,N_14719,N_13649);
or UO_142 (O_142,N_14577,N_13091);
nor UO_143 (O_143,N_14250,N_14617);
nor UO_144 (O_144,N_14502,N_12570);
or UO_145 (O_145,N_12659,N_12112);
nor UO_146 (O_146,N_12737,N_13038);
and UO_147 (O_147,N_12468,N_13571);
and UO_148 (O_148,N_12281,N_12888);
or UO_149 (O_149,N_12457,N_14124);
and UO_150 (O_150,N_13692,N_13283);
nor UO_151 (O_151,N_13163,N_12508);
nor UO_152 (O_152,N_13977,N_13769);
nand UO_153 (O_153,N_12650,N_13288);
and UO_154 (O_154,N_12536,N_14239);
nand UO_155 (O_155,N_13010,N_12354);
or UO_156 (O_156,N_12092,N_12525);
nand UO_157 (O_157,N_13135,N_12635);
nand UO_158 (O_158,N_14760,N_12611);
nor UO_159 (O_159,N_14884,N_14136);
or UO_160 (O_160,N_12519,N_12075);
nand UO_161 (O_161,N_12683,N_13170);
or UO_162 (O_162,N_12455,N_12065);
or UO_163 (O_163,N_12196,N_13838);
and UO_164 (O_164,N_13872,N_12335);
nor UO_165 (O_165,N_12649,N_14295);
nor UO_166 (O_166,N_14352,N_13493);
nand UO_167 (O_167,N_13588,N_12658);
nor UO_168 (O_168,N_13947,N_14278);
nor UO_169 (O_169,N_12015,N_14102);
or UO_170 (O_170,N_12349,N_13614);
and UO_171 (O_171,N_14036,N_13253);
nor UO_172 (O_172,N_14890,N_12640);
or UO_173 (O_173,N_13564,N_13463);
and UO_174 (O_174,N_12767,N_12411);
or UO_175 (O_175,N_12989,N_14863);
nor UO_176 (O_176,N_13462,N_12171);
nor UO_177 (O_177,N_12820,N_12016);
nand UO_178 (O_178,N_14075,N_13985);
xor UO_179 (O_179,N_14174,N_12966);
nor UO_180 (O_180,N_14592,N_12032);
nand UO_181 (O_181,N_13447,N_13638);
or UO_182 (O_182,N_12019,N_12382);
nor UO_183 (O_183,N_12255,N_12158);
nand UO_184 (O_184,N_14997,N_14003);
nor UO_185 (O_185,N_12945,N_13382);
nand UO_186 (O_186,N_12388,N_14576);
and UO_187 (O_187,N_14158,N_12049);
nand UO_188 (O_188,N_12037,N_14793);
or UO_189 (O_189,N_14169,N_14875);
and UO_190 (O_190,N_13232,N_13194);
nor UO_191 (O_191,N_12079,N_14469);
and UO_192 (O_192,N_14853,N_14657);
nand UO_193 (O_193,N_14862,N_12923);
nand UO_194 (O_194,N_13634,N_12936);
nor UO_195 (O_195,N_14157,N_13844);
and UO_196 (O_196,N_14637,N_14154);
or UO_197 (O_197,N_12875,N_14931);
or UO_198 (O_198,N_12755,N_12285);
nand UO_199 (O_199,N_14497,N_14271);
nand UO_200 (O_200,N_13741,N_13965);
nand UO_201 (O_201,N_13092,N_12303);
nand UO_202 (O_202,N_14303,N_12872);
nor UO_203 (O_203,N_13502,N_12808);
nand UO_204 (O_204,N_12339,N_13559);
nor UO_205 (O_205,N_13082,N_14054);
nor UO_206 (O_206,N_12398,N_12885);
and UO_207 (O_207,N_13889,N_13146);
nand UO_208 (O_208,N_13468,N_14100);
and UO_209 (O_209,N_12211,N_14038);
and UO_210 (O_210,N_12314,N_14962);
xor UO_211 (O_211,N_13214,N_14113);
and UO_212 (O_212,N_13364,N_13654);
or UO_213 (O_213,N_13558,N_12323);
nand UO_214 (O_214,N_13160,N_14041);
and UO_215 (O_215,N_12116,N_13905);
or UO_216 (O_216,N_12183,N_14768);
or UO_217 (O_217,N_14757,N_12803);
nor UO_218 (O_218,N_12772,N_13971);
nand UO_219 (O_219,N_12462,N_12318);
and UO_220 (O_220,N_14604,N_12681);
and UO_221 (O_221,N_14838,N_12366);
nor UO_222 (O_222,N_14405,N_12535);
nor UO_223 (O_223,N_13842,N_13310);
nor UO_224 (O_224,N_14423,N_12882);
nor UO_225 (O_225,N_13650,N_12402);
or UO_226 (O_226,N_13633,N_14912);
nor UO_227 (O_227,N_14555,N_14950);
and UO_228 (O_228,N_12917,N_13198);
nor UO_229 (O_229,N_12157,N_12702);
nor UO_230 (O_230,N_14532,N_12110);
or UO_231 (O_231,N_13937,N_14107);
or UO_232 (O_232,N_14984,N_12637);
nor UO_233 (O_233,N_14536,N_14165);
or UO_234 (O_234,N_13177,N_13949);
or UO_235 (O_235,N_13832,N_13783);
nand UO_236 (O_236,N_13539,N_13648);
nor UO_237 (O_237,N_13039,N_14190);
nor UO_238 (O_238,N_12014,N_14027);
nand UO_239 (O_239,N_12194,N_12356);
or UO_240 (O_240,N_13084,N_12780);
nand UO_241 (O_241,N_14612,N_12297);
and UO_242 (O_242,N_14578,N_14094);
or UO_243 (O_243,N_14928,N_13707);
or UO_244 (O_244,N_13647,N_14800);
nor UO_245 (O_245,N_12170,N_14167);
nand UO_246 (O_246,N_12278,N_14478);
and UO_247 (O_247,N_13210,N_12909);
nor UO_248 (O_248,N_12283,N_13385);
and UO_249 (O_249,N_13998,N_14304);
nor UO_250 (O_250,N_13815,N_13906);
xnor UO_251 (O_251,N_14225,N_12262);
and UO_252 (O_252,N_13980,N_12916);
or UO_253 (O_253,N_13963,N_13280);
and UO_254 (O_254,N_13426,N_13254);
or UO_255 (O_255,N_12093,N_12573);
and UO_256 (O_256,N_14586,N_13250);
or UO_257 (O_257,N_13240,N_12581);
or UO_258 (O_258,N_14078,N_13525);
or UO_259 (O_259,N_14741,N_14982);
and UO_260 (O_260,N_12958,N_13867);
and UO_261 (O_261,N_12986,N_12691);
or UO_262 (O_262,N_13785,N_12125);
nand UO_263 (O_263,N_14818,N_13912);
nand UO_264 (O_264,N_12160,N_13435);
or UO_265 (O_265,N_12336,N_14069);
or UO_266 (O_266,N_13313,N_13579);
nand UO_267 (O_267,N_14376,N_12475);
and UO_268 (O_268,N_12133,N_12661);
and UO_269 (O_269,N_13846,N_13046);
nand UO_270 (O_270,N_13806,N_12463);
nor UO_271 (O_271,N_13970,N_13809);
nor UO_272 (O_272,N_13645,N_12493);
or UO_273 (O_273,N_12645,N_14211);
nand UO_274 (O_274,N_12239,N_13864);
nand UO_275 (O_275,N_13048,N_12131);
nand UO_276 (O_276,N_13978,N_13733);
nand UO_277 (O_277,N_12898,N_14994);
and UO_278 (O_278,N_14980,N_14883);
and UO_279 (O_279,N_14270,N_12122);
nand UO_280 (O_280,N_12775,N_13472);
or UO_281 (O_281,N_13907,N_13482);
xnor UO_282 (O_282,N_12351,N_13450);
nor UO_283 (O_283,N_12421,N_14005);
nor UO_284 (O_284,N_12657,N_13414);
or UO_285 (O_285,N_12944,N_14674);
or UO_286 (O_286,N_14517,N_13766);
and UO_287 (O_287,N_13229,N_13753);
and UO_288 (O_288,N_14626,N_13774);
xnor UO_289 (O_289,N_13400,N_14479);
and UO_290 (O_290,N_13916,N_13286);
and UO_291 (O_291,N_12861,N_13190);
nor UO_292 (O_292,N_13252,N_14499);
and UO_293 (O_293,N_13713,N_13261);
or UO_294 (O_294,N_12141,N_14573);
and UO_295 (O_295,N_12817,N_14727);
and UO_296 (O_296,N_12964,N_13933);
nor UO_297 (O_297,N_12546,N_12295);
and UO_298 (O_298,N_13077,N_13773);
nor UO_299 (O_299,N_14447,N_13183);
and UO_300 (O_300,N_13118,N_12965);
or UO_301 (O_301,N_13911,N_12363);
nor UO_302 (O_302,N_13538,N_12520);
or UO_303 (O_303,N_14711,N_12423);
or UO_304 (O_304,N_13913,N_12669);
and UO_305 (O_305,N_13522,N_13557);
nand UO_306 (O_306,N_13891,N_14850);
nand UO_307 (O_307,N_14435,N_12488);
or UO_308 (O_308,N_12175,N_12105);
nor UO_309 (O_309,N_13480,N_14686);
and UO_310 (O_310,N_14847,N_12979);
or UO_311 (O_311,N_12866,N_14120);
and UO_312 (O_312,N_12590,N_14261);
nand UO_313 (O_313,N_13058,N_12948);
nand UO_314 (O_314,N_13018,N_14417);
nand UO_315 (O_315,N_14411,N_13982);
or UO_316 (O_316,N_12526,N_12750);
nand UO_317 (O_317,N_14334,N_13192);
and UO_318 (O_318,N_14259,N_14287);
or UO_319 (O_319,N_13367,N_14426);
or UO_320 (O_320,N_12745,N_12209);
nand UO_321 (O_321,N_13088,N_13403);
nand UO_322 (O_322,N_13222,N_14722);
or UO_323 (O_323,N_13489,N_14275);
nor UO_324 (O_324,N_14237,N_14968);
nor UO_325 (O_325,N_14509,N_12073);
or UO_326 (O_326,N_13685,N_13481);
and UO_327 (O_327,N_14333,N_12862);
or UO_328 (O_328,N_12715,N_12890);
or UO_329 (O_329,N_13111,N_14083);
and UO_330 (O_330,N_14222,N_14422);
and UO_331 (O_331,N_13817,N_13431);
nand UO_332 (O_332,N_14559,N_13640);
nand UO_333 (O_333,N_12543,N_13075);
or UO_334 (O_334,N_13115,N_12061);
nand UO_335 (O_335,N_12486,N_12050);
nor UO_336 (O_336,N_13519,N_14913);
and UO_337 (O_337,N_12166,N_13790);
and UO_338 (O_338,N_14649,N_12770);
nor UO_339 (O_339,N_13184,N_13943);
and UO_340 (O_340,N_13744,N_14432);
nor UO_341 (O_341,N_14129,N_13483);
or UO_342 (O_342,N_14848,N_14959);
and UO_343 (O_343,N_14636,N_14365);
nand UO_344 (O_344,N_14519,N_14343);
nor UO_345 (O_345,N_12721,N_12026);
or UO_346 (O_346,N_13636,N_14831);
nor UO_347 (O_347,N_14842,N_13314);
nand UO_348 (O_348,N_14764,N_12460);
and UO_349 (O_349,N_12082,N_14791);
and UO_350 (O_350,N_13603,N_13424);
nand UO_351 (O_351,N_14115,N_12289);
and UO_352 (O_352,N_12057,N_13452);
nand UO_353 (O_353,N_12922,N_14391);
and UO_354 (O_354,N_14729,N_13545);
nor UO_355 (O_355,N_14055,N_13812);
nor UO_356 (O_356,N_13979,N_13706);
nor UO_357 (O_357,N_13455,N_14461);
and UO_358 (O_358,N_12176,N_12465);
and UO_359 (O_359,N_14146,N_12268);
or UO_360 (O_360,N_12980,N_12913);
or UO_361 (O_361,N_13020,N_12403);
nor UO_362 (O_362,N_12372,N_13464);
or UO_363 (O_363,N_14939,N_12001);
or UO_364 (O_364,N_14565,N_12740);
or UO_365 (O_365,N_14349,N_14882);
nor UO_366 (O_366,N_12968,N_12582);
and UO_367 (O_367,N_13151,N_13674);
nor UO_368 (O_368,N_14240,N_13787);
nand UO_369 (O_369,N_12731,N_12638);
nor UO_370 (O_370,N_13282,N_14244);
and UO_371 (O_371,N_14851,N_13487);
nand UO_372 (O_372,N_12328,N_12569);
or UO_373 (O_373,N_14067,N_14785);
nand UO_374 (O_374,N_14452,N_14624);
nand UO_375 (O_375,N_14314,N_12288);
and UO_376 (O_376,N_12636,N_13607);
and UO_377 (O_377,N_13541,N_14937);
nand UO_378 (O_378,N_12993,N_12863);
or UO_379 (O_379,N_14436,N_14537);
and UO_380 (O_380,N_12618,N_12709);
nor UO_381 (O_381,N_13735,N_12839);
and UO_382 (O_382,N_13412,N_13223);
nand UO_383 (O_383,N_14231,N_13119);
or UO_384 (O_384,N_13117,N_13373);
nor UO_385 (O_385,N_14286,N_13848);
nand UO_386 (O_386,N_12730,N_12688);
and UO_387 (O_387,N_14714,N_12656);
or UO_388 (O_388,N_12011,N_14654);
nand UO_389 (O_389,N_13410,N_13546);
and UO_390 (O_390,N_13158,N_13231);
and UO_391 (O_391,N_14560,N_12850);
nor UO_392 (O_392,N_12952,N_13078);
nand UO_393 (O_393,N_14998,N_14377);
nor UO_394 (O_394,N_12162,N_13925);
nand UO_395 (O_395,N_14777,N_12013);
or UO_396 (O_396,N_13712,N_14767);
nor UO_397 (O_397,N_14914,N_12163);
and UO_398 (O_398,N_13968,N_14776);
and UO_399 (O_399,N_14506,N_14424);
nand UO_400 (O_400,N_12806,N_14718);
and UO_401 (O_401,N_13300,N_14656);
nand UO_402 (O_402,N_12891,N_13550);
nand UO_403 (O_403,N_13698,N_13140);
and UO_404 (O_404,N_12942,N_13132);
nand UO_405 (O_405,N_12853,N_12714);
nor UO_406 (O_406,N_14336,N_12321);
nand UO_407 (O_407,N_13677,N_14212);
or UO_408 (O_408,N_12114,N_12541);
nor UO_409 (O_409,N_12879,N_14114);
or UO_410 (O_410,N_12886,N_12954);
and UO_411 (O_411,N_12734,N_12855);
or UO_412 (O_412,N_14874,N_12502);
and UO_413 (O_413,N_13771,N_12165);
or UO_414 (O_414,N_13855,N_12097);
nand UO_415 (O_415,N_12860,N_12873);
nand UO_416 (O_416,N_13054,N_13325);
and UO_417 (O_417,N_13622,N_12091);
nand UO_418 (O_418,N_14198,N_14589);
nand UO_419 (O_419,N_13055,N_12220);
nor UO_420 (O_420,N_12956,N_14712);
nand UO_421 (O_421,N_12680,N_13600);
and UO_422 (O_422,N_13779,N_13594);
and UO_423 (O_423,N_14515,N_14596);
nand UO_424 (O_424,N_14441,N_12071);
and UO_425 (O_425,N_14710,N_12791);
nor UO_426 (O_426,N_13667,N_13176);
and UO_427 (O_427,N_14684,N_13663);
nand UO_428 (O_428,N_13467,N_13257);
and UO_429 (O_429,N_14717,N_14825);
and UO_430 (O_430,N_12400,N_13643);
xnor UO_431 (O_431,N_13954,N_13556);
nor UO_432 (O_432,N_14018,N_14249);
nand UO_433 (O_433,N_12577,N_13419);
nor UO_434 (O_434,N_12111,N_12219);
and UO_435 (O_435,N_12515,N_14949);
nand UO_436 (O_436,N_14598,N_13073);
and UO_437 (O_437,N_13655,N_14451);
and UO_438 (O_438,N_13366,N_12599);
nand UO_439 (O_439,N_12858,N_14125);
nand UO_440 (O_440,N_14689,N_13488);
nor UO_441 (O_441,N_12036,N_13624);
nand UO_442 (O_442,N_14400,N_12243);
or UO_443 (O_443,N_13597,N_13868);
and UO_444 (O_444,N_13218,N_14370);
and UO_445 (O_445,N_13576,N_14993);
nand UO_446 (O_446,N_14150,N_12113);
nor UO_447 (O_447,N_12352,N_12499);
nor UO_448 (O_448,N_12369,N_12641);
nor UO_449 (O_449,N_13799,N_14983);
nor UO_450 (O_450,N_13941,N_13670);
and UO_451 (O_451,N_14260,N_12184);
or UO_452 (O_452,N_13966,N_14501);
or UO_453 (O_453,N_12434,N_12228);
nor UO_454 (O_454,N_12428,N_14236);
and UO_455 (O_455,N_12950,N_12701);
and UO_456 (O_456,N_14408,N_14317);
nand UO_457 (O_457,N_12346,N_14836);
and UO_458 (O_458,N_14516,N_13266);
or UO_459 (O_459,N_14459,N_14756);
or UO_460 (O_460,N_14881,N_13307);
and UO_461 (O_461,N_14567,N_13457);
and UO_462 (O_462,N_13895,N_14098);
and UO_463 (O_463,N_12642,N_12245);
nor UO_464 (O_464,N_12673,N_14969);
or UO_465 (O_465,N_14683,N_13860);
and UO_466 (O_466,N_12527,N_13441);
nand UO_467 (O_467,N_14111,N_13376);
nor UO_468 (O_468,N_14870,N_13794);
nor UO_469 (O_469,N_14666,N_14491);
nor UO_470 (O_470,N_14663,N_12506);
nor UO_471 (O_471,N_14557,N_12427);
or UO_472 (O_472,N_13758,N_12309);
or UO_473 (O_473,N_12576,N_12491);
nor UO_474 (O_474,N_12869,N_13927);
and UO_475 (O_475,N_12912,N_13023);
nor UO_476 (O_476,N_14542,N_12751);
nand UO_477 (O_477,N_14085,N_12560);
nand UO_478 (O_478,N_12816,N_14128);
nand UO_479 (O_479,N_12273,N_14533);
or UO_480 (O_480,N_12367,N_14979);
and UO_481 (O_481,N_14911,N_13196);
nor UO_482 (O_482,N_14963,N_12250);
and UO_483 (O_483,N_14611,N_13478);
or UO_484 (O_484,N_14347,N_14344);
nand UO_485 (O_485,N_14601,N_14210);
or UO_486 (O_486,N_12505,N_14795);
nand UO_487 (O_487,N_12189,N_12007);
nor UO_488 (O_488,N_13531,N_13616);
or UO_489 (O_489,N_14687,N_12622);
nor UO_490 (O_490,N_12210,N_12906);
nand UO_491 (O_491,N_12778,N_13595);
nor UO_492 (O_492,N_13062,N_12088);
nor UO_493 (O_493,N_12010,N_12155);
nand UO_494 (O_494,N_12988,N_13665);
nand UO_495 (O_495,N_13299,N_12823);
nand UO_496 (O_496,N_13236,N_13276);
nor UO_497 (O_497,N_13515,N_12130);
or UO_498 (O_498,N_12555,N_13258);
or UO_499 (O_499,N_12087,N_12769);
nor UO_500 (O_500,N_14690,N_13703);
and UO_501 (O_501,N_14229,N_14215);
nor UO_502 (O_502,N_14481,N_12689);
and UO_503 (O_503,N_12707,N_13620);
and UO_504 (O_504,N_14328,N_13204);
nor UO_505 (O_505,N_12054,N_12677);
or UO_506 (O_506,N_13520,N_12038);
nor UO_507 (O_507,N_13197,N_14771);
nor UO_508 (O_508,N_14902,N_12974);
nand UO_509 (O_509,N_13813,N_13275);
nand UO_510 (O_510,N_13591,N_12067);
nor UO_511 (O_511,N_12381,N_13205);
and UO_512 (O_512,N_12501,N_13763);
nor UO_513 (O_513,N_13191,N_14309);
or UO_514 (O_514,N_12103,N_12601);
xnor UO_515 (O_515,N_14425,N_14780);
and UO_516 (O_516,N_13416,N_14877);
nand UO_517 (O_517,N_13287,N_14356);
or UO_518 (O_518,N_12045,N_14170);
nand UO_519 (O_519,N_12144,N_13629);
nand UO_520 (O_520,N_12926,N_12058);
nor UO_521 (O_521,N_13021,N_12341);
or UO_522 (O_522,N_14620,N_12246);
and UO_523 (O_523,N_14942,N_12787);
nand UO_524 (O_524,N_13876,N_12881);
nor UO_525 (O_525,N_12644,N_12492);
or UO_526 (O_526,N_14247,N_13434);
nor UO_527 (O_527,N_14692,N_13173);
and UO_528 (O_528,N_13825,N_13989);
and UO_529 (O_529,N_12595,N_14856);
and UO_530 (O_530,N_12794,N_12467);
nor UO_531 (O_531,N_12761,N_14442);
and UO_532 (O_532,N_12199,N_14277);
nand UO_533 (O_533,N_13764,N_12325);
nor UO_534 (O_534,N_12654,N_13186);
nand UO_535 (O_535,N_12118,N_12729);
nor UO_536 (O_536,N_12397,N_13936);
nor UO_537 (O_537,N_14750,N_14602);
nor UO_538 (O_538,N_13042,N_14739);
or UO_539 (O_539,N_12845,N_12401);
nor UO_540 (O_540,N_12461,N_14379);
nand UO_541 (O_541,N_12710,N_13221);
and UO_542 (O_542,N_13244,N_14889);
nor UO_543 (O_543,N_14161,N_14569);
or UO_544 (O_544,N_12198,N_14915);
and UO_545 (O_545,N_14954,N_12237);
nor UO_546 (O_546,N_13931,N_13923);
and UO_547 (O_547,N_13490,N_14907);
nor UO_548 (O_548,N_12435,N_14747);
and UO_549 (O_549,N_14618,N_13788);
or UO_550 (O_550,N_13142,N_14172);
and UO_551 (O_551,N_14058,N_13930);
or UO_552 (O_552,N_14953,N_13894);
and UO_553 (O_553,N_12578,N_14733);
and UO_554 (O_554,N_13390,N_13508);
nand UO_555 (O_555,N_13919,N_14832);
or UO_556 (O_556,N_13179,N_14133);
nand UO_557 (O_557,N_13139,N_12703);
or UO_558 (O_558,N_12416,N_14936);
nand UO_559 (O_559,N_13696,N_12589);
nand UO_560 (O_560,N_13732,N_12614);
and UO_561 (O_561,N_13357,N_12101);
nand UO_562 (O_562,N_14413,N_13290);
or UO_563 (O_563,N_14591,N_13473);
or UO_564 (O_564,N_14076,N_12124);
and UO_565 (O_565,N_13368,N_12062);
and UO_566 (O_566,N_13233,N_14600);
nor UO_567 (O_567,N_12338,N_14022);
or UO_568 (O_568,N_14742,N_14224);
or UO_569 (O_569,N_12134,N_12003);
or UO_570 (O_570,N_13323,N_12963);
and UO_571 (O_571,N_12490,N_13939);
or UO_572 (O_572,N_14740,N_13755);
nor UO_573 (O_573,N_14357,N_14607);
or UO_574 (O_574,N_14269,N_12291);
nor UO_575 (O_575,N_14819,N_14678);
nor UO_576 (O_576,N_12298,N_14305);
or UO_577 (O_577,N_14951,N_14039);
nor UO_578 (O_578,N_14904,N_14143);
nand UO_579 (O_579,N_14545,N_12234);
nand UO_580 (O_580,N_14052,N_13704);
or UO_581 (O_581,N_12296,N_13355);
or UO_582 (O_582,N_13561,N_12854);
nand UO_583 (O_583,N_13530,N_12322);
nor UO_584 (O_584,N_14121,N_14787);
nand UO_585 (O_585,N_14415,N_13596);
or UO_586 (O_586,N_12624,N_13729);
nor UO_587 (O_587,N_14016,N_14547);
nor UO_588 (O_588,N_13359,N_12852);
nand UO_589 (O_589,N_14028,N_14045);
and UO_590 (O_590,N_14930,N_13418);
nor UO_591 (O_591,N_13458,N_13526);
or UO_592 (O_592,N_13474,N_12432);
nand UO_593 (O_593,N_12343,N_14910);
nand UO_594 (O_594,N_12064,N_12357);
nand UO_595 (O_595,N_14393,N_13193);
or UO_596 (O_596,N_14088,N_12182);
and UO_597 (O_597,N_14371,N_13599);
and UO_598 (O_598,N_13569,N_13259);
nor UO_599 (O_599,N_12480,N_13702);
and UO_600 (O_600,N_13182,N_13554);
nor UO_601 (O_601,N_13302,N_12606);
and UO_602 (O_602,N_13540,N_13093);
nand UO_603 (O_603,N_12782,N_12897);
or UO_604 (O_604,N_14428,N_12998);
and UO_605 (O_605,N_14669,N_12208);
or UO_606 (O_606,N_12908,N_13896);
nand UO_607 (O_607,N_13756,N_12549);
and UO_608 (O_608,N_12943,N_14414);
and UO_609 (O_609,N_13491,N_12084);
nand UO_610 (O_610,N_14653,N_13507);
or UO_611 (O_611,N_14566,N_12884);
and UO_612 (O_612,N_14570,N_13628);
and UO_613 (O_613,N_13801,N_12631);
nor UO_614 (O_614,N_14691,N_13285);
or UO_615 (O_615,N_12192,N_14730);
nor UO_616 (O_616,N_14440,N_13040);
nor UO_617 (O_617,N_13167,N_14676);
and UO_618 (O_618,N_12139,N_12018);
or UO_619 (O_619,N_12776,N_14629);
or UO_620 (O_620,N_14255,N_13884);
and UO_621 (O_621,N_13069,N_12331);
and UO_622 (O_622,N_14964,N_13778);
nand UO_623 (O_623,N_13428,N_13432);
or UO_624 (O_624,N_14978,N_12900);
nand UO_625 (O_625,N_14990,N_13272);
and UO_626 (O_626,N_12241,N_12699);
nor UO_627 (O_627,N_13249,N_12825);
nand UO_628 (O_628,N_14891,N_12020);
nand UO_629 (O_629,N_13852,N_12380);
nor UO_630 (O_630,N_12304,N_14878);
nor UO_631 (O_631,N_13866,N_13679);
or UO_632 (O_632,N_12446,N_13826);
nor UO_633 (O_633,N_14677,N_12533);
and UO_634 (O_634,N_12542,N_14164);
or UO_635 (O_635,N_13567,N_12177);
or UO_636 (O_636,N_13187,N_13731);
or UO_637 (O_637,N_14313,N_14443);
and UO_638 (O_638,N_13098,N_14346);
nor UO_639 (O_639,N_12299,N_12878);
or UO_640 (O_640,N_12668,N_12167);
nand UO_641 (O_641,N_13604,N_13331);
nand UO_642 (O_642,N_14681,N_14845);
nor UO_643 (O_643,N_12256,N_12264);
or UO_644 (O_644,N_12405,N_12274);
nor UO_645 (O_645,N_12918,N_12695);
and UO_646 (O_646,N_12666,N_12052);
nand UO_647 (O_647,N_14407,N_12620);
nor UO_648 (O_648,N_13013,N_14934);
nand UO_649 (O_649,N_14050,N_13945);
nand UO_650 (O_650,N_14382,N_12154);
nor UO_651 (O_651,N_12925,N_13066);
and UO_652 (O_652,N_14916,N_12284);
or UO_653 (O_653,N_13807,N_12662);
nor UO_654 (O_654,N_12568,N_13668);
nand UO_655 (O_655,N_13284,N_12920);
nor UO_656 (O_656,N_12072,N_12743);
nand UO_657 (O_657,N_14988,N_13208);
nor UO_658 (O_658,N_14171,N_12509);
or UO_659 (O_659,N_13380,N_13496);
and UO_660 (O_660,N_12831,N_13672);
and UO_661 (O_661,N_13877,N_13740);
and UO_662 (O_662,N_14033,N_14640);
and UO_663 (O_663,N_13751,N_14470);
and UO_664 (O_664,N_14861,N_14324);
and UO_665 (O_665,N_14679,N_14775);
nor UO_666 (O_666,N_14040,N_13716);
and UO_667 (O_667,N_14715,N_12970);
nand UO_668 (O_668,N_13765,N_14390);
or UO_669 (O_669,N_14135,N_14940);
nand UO_670 (O_670,N_14108,N_14206);
or UO_671 (O_671,N_14178,N_13984);
and UO_672 (O_672,N_12143,N_14521);
nand UO_673 (O_673,N_13157,N_13909);
or UO_674 (O_674,N_13059,N_14946);
and UO_675 (O_675,N_12080,N_12365);
and UO_676 (O_676,N_12786,N_14494);
nor UO_677 (O_677,N_14388,N_14162);
and UO_678 (O_678,N_12537,N_12790);
nor UO_679 (O_679,N_12760,N_14021);
nor UO_680 (O_680,N_14410,N_13156);
and UO_681 (O_681,N_12251,N_13995);
nand UO_682 (O_682,N_12329,N_14335);
nand UO_683 (O_683,N_13016,N_13823);
or UO_684 (O_684,N_14082,N_12311);
and UO_685 (O_685,N_14168,N_13404);
and UO_686 (O_686,N_14483,N_14864);
nor UO_687 (O_687,N_12670,N_14456);
or UO_688 (O_688,N_14996,N_12418);
nand UO_689 (O_689,N_13356,N_14412);
and UO_690 (O_690,N_14794,N_13708);
nor UO_691 (O_691,N_12871,N_12764);
nand UO_692 (O_692,N_14728,N_14700);
and UO_693 (O_693,N_14342,N_13264);
nand UO_694 (O_694,N_12571,N_14246);
or UO_695 (O_695,N_13646,N_13899);
nand UO_696 (O_696,N_12353,N_12083);
nor UO_697 (O_697,N_13676,N_13294);
and UO_698 (O_698,N_13166,N_12904);
and UO_699 (O_699,N_14397,N_13700);
nor UO_700 (O_700,N_12017,N_13334);
nor UO_701 (O_701,N_14026,N_13513);
nand UO_702 (O_702,N_14490,N_12174);
and UO_703 (O_703,N_13883,N_12302);
or UO_704 (O_704,N_12300,N_14688);
nor UO_705 (O_705,N_12552,N_12368);
nor UO_706 (O_706,N_13901,N_14790);
and UO_707 (O_707,N_14805,N_13161);
nand UO_708 (O_708,N_12370,N_12655);
and UO_709 (O_709,N_13510,N_12218);
or UO_710 (O_710,N_14263,N_12362);
or UO_711 (O_711,N_13351,N_12230);
and UO_712 (O_712,N_13199,N_12437);
nand UO_713 (O_713,N_12837,N_12708);
and UO_714 (O_714,N_13681,N_13705);
or UO_715 (O_715,N_13960,N_14181);
nand UO_716 (O_716,N_12035,N_14759);
nand UO_717 (O_717,N_13451,N_14361);
nor UO_718 (O_718,N_13255,N_12249);
or UO_719 (O_719,N_13350,N_14004);
nand UO_720 (O_720,N_13427,N_14512);
and UO_721 (O_721,N_14614,N_14531);
and UO_722 (O_722,N_12315,N_14755);
or UO_723 (O_723,N_13397,N_14369);
and UO_724 (O_724,N_13442,N_12021);
or UO_725 (O_725,N_14732,N_13471);
and UO_726 (O_726,N_12150,N_14648);
xnor UO_727 (O_727,N_12099,N_12651);
and UO_728 (O_728,N_13509,N_13856);
or UO_729 (O_729,N_13131,N_14530);
nand UO_730 (O_730,N_14043,N_12277);
or UO_731 (O_731,N_13739,N_14192);
or UO_732 (O_732,N_12895,N_14546);
nor UO_733 (O_733,N_13224,N_13371);
nand UO_734 (O_734,N_12306,N_14386);
nor UO_735 (O_735,N_13083,N_12924);
nor UO_736 (O_736,N_14661,N_13999);
nand UO_737 (O_737,N_14487,N_14326);
nand UO_738 (O_738,N_12000,N_13164);
nor UO_739 (O_739,N_13611,N_14037);
and UO_740 (O_740,N_13030,N_14685);
or UO_741 (O_741,N_12317,N_12594);
nor UO_742 (O_742,N_14392,N_12153);
nor UO_743 (O_743,N_14288,N_14202);
nor UO_744 (O_744,N_12931,N_13534);
and UO_745 (O_745,N_13737,N_13120);
or UO_746 (O_746,N_13932,N_14608);
and UO_747 (O_747,N_12551,N_14976);
or UO_748 (O_748,N_14563,N_13962);
or UO_749 (O_749,N_12937,N_13678);
or UO_750 (O_750,N_14758,N_14095);
and UO_751 (O_751,N_12819,N_14507);
or UO_752 (O_752,N_14948,N_12567);
nand UO_753 (O_753,N_13802,N_14921);
xnor UO_754 (O_754,N_12373,N_13893);
and UO_755 (O_755,N_14439,N_13695);
or UO_756 (O_756,N_13203,N_14207);
nand UO_757 (O_757,N_13928,N_14553);
nor UO_758 (O_758,N_12456,N_12994);
and UO_759 (O_759,N_12410,N_13606);
and UO_760 (O_760,N_14311,N_12385);
and UO_761 (O_761,N_14792,N_13134);
nor UO_762 (O_762,N_13590,N_12269);
or UO_763 (O_763,N_12686,N_12443);
nand UO_764 (O_764,N_14788,N_12375);
or UO_765 (O_765,N_14627,N_13498);
and UO_766 (O_766,N_12621,N_14905);
and UO_767 (O_767,N_14472,N_12991);
nor UO_768 (O_768,N_13391,N_13776);
or UO_769 (O_769,N_12056,N_12919);
nor UO_770 (O_770,N_12899,N_12173);
nand UO_771 (O_771,N_14935,N_14475);
and UO_772 (O_772,N_14524,N_13270);
nand UO_773 (O_773,N_12117,N_12212);
nor UO_774 (O_774,N_12248,N_13521);
or UO_775 (O_775,N_14103,N_14880);
and UO_776 (O_776,N_12516,N_13718);
or UO_777 (O_777,N_13251,N_12946);
and UO_778 (O_778,N_14814,N_13180);
nor UO_779 (O_779,N_13004,N_14652);
nand UO_780 (O_780,N_14032,N_12415);
nand UO_781 (O_781,N_13994,N_14378);
and UO_782 (O_782,N_12867,N_12625);
nand UO_783 (O_783,N_13219,N_12060);
and UO_784 (O_784,N_12078,N_12027);
nand UO_785 (O_785,N_13915,N_13337);
or UO_786 (O_786,N_12347,N_14079);
nand UO_787 (O_787,N_13316,N_12921);
or UO_788 (O_788,N_12634,N_13422);
nor UO_789 (O_789,N_12874,N_14738);
nand UO_790 (O_790,N_12583,N_13859);
or UO_791 (O_791,N_13565,N_12796);
nor UO_792 (O_792,N_13686,N_14960);
nor UO_793 (O_793,N_14665,N_13575);
or UO_794 (O_794,N_14060,N_13090);
nand UO_795 (O_795,N_14562,N_12824);
or UO_796 (O_796,N_12805,N_14522);
or UO_797 (O_797,N_14123,N_13612);
and UO_798 (O_798,N_14704,N_13536);
xnor UO_799 (O_799,N_13476,N_13201);
nor UO_800 (O_800,N_12700,N_14467);
nand UO_801 (O_801,N_14908,N_13991);
or UO_802 (O_802,N_13782,N_12947);
xor UO_803 (O_803,N_12140,N_14337);
nand UO_804 (O_804,N_13050,N_13697);
and UO_805 (O_805,N_12771,N_12327);
nor UO_806 (O_806,N_13109,N_13983);
nand UO_807 (O_807,N_13730,N_13415);
nand UO_808 (O_808,N_12464,N_13828);
nand UO_809 (O_809,N_13549,N_13243);
or UO_810 (O_810,N_13100,N_13318);
nor UO_811 (O_811,N_13362,N_13104);
or UO_812 (O_812,N_12450,N_14616);
nor UO_813 (O_813,N_12012,N_13171);
or UO_814 (O_814,N_13022,N_12783);
nand UO_815 (O_815,N_13110,N_13857);
and UO_816 (O_816,N_14778,N_14477);
or UO_817 (O_817,N_12364,N_12720);
xnor UO_818 (O_818,N_13661,N_13910);
nor UO_819 (O_819,N_14833,N_14748);
nand UO_820 (O_820,N_13107,N_14266);
or UO_821 (O_821,N_12253,N_12613);
and UO_822 (O_822,N_12718,N_14308);
nand UO_823 (O_823,N_13348,N_12746);
or UO_824 (O_824,N_14900,N_13644);
or UO_825 (O_825,N_13425,N_12135);
nor UO_826 (O_826,N_12697,N_14802);
nand UO_827 (O_827,N_12172,N_14145);
or UO_828 (O_828,N_14644,N_13440);
and UO_829 (O_829,N_12981,N_12675);
nand UO_830 (O_830,N_14645,N_13881);
or UO_831 (O_831,N_14089,N_13238);
or UO_832 (O_832,N_13738,N_12308);
or UO_833 (O_833,N_12992,N_14599);
and UO_834 (O_834,N_14899,N_14709);
nor UO_835 (O_835,N_12378,N_12758);
xnor UO_836 (O_836,N_14216,N_13298);
nand UO_837 (O_837,N_12564,N_14380);
and UO_838 (O_838,N_14453,N_12260);
and UO_839 (O_839,N_14753,N_14500);
nand UO_840 (O_840,N_13319,N_12827);
nand UO_841 (O_841,N_12727,N_14981);
or UO_842 (O_842,N_13870,N_14364);
nand UO_843 (O_843,N_12310,N_12407);
or UO_844 (O_844,N_14292,N_12557);
nor UO_845 (O_845,N_14584,N_14127);
or UO_846 (O_846,N_13841,N_12484);
and UO_847 (O_847,N_14199,N_14564);
nor UO_848 (O_848,N_14667,N_12213);
nor UO_849 (O_849,N_14009,N_13466);
nand UO_850 (O_850,N_13353,N_14281);
nor UO_851 (O_851,N_12217,N_12738);
nor UO_852 (O_852,N_12185,N_14438);
nand UO_853 (O_853,N_12550,N_13850);
nand UO_854 (O_854,N_14051,N_14323);
or UO_855 (O_855,N_13673,N_13843);
nand UO_856 (O_856,N_14635,N_14746);
nand UO_857 (O_857,N_12889,N_12826);
nor UO_858 (O_858,N_13370,N_12724);
and UO_859 (O_859,N_12562,N_13693);
nand UO_860 (O_860,N_12643,N_12190);
nor UO_861 (O_861,N_14134,N_14815);
and UO_862 (O_862,N_12859,N_14658);
and UO_863 (O_863,N_12433,N_13952);
or UO_864 (O_864,N_13095,N_13532);
and UO_865 (O_865,N_13724,N_14331);
and UO_866 (O_866,N_14218,N_14126);
and UO_867 (O_867,N_12361,N_13719);
and UO_868 (O_868,N_14895,N_12807);
or UO_869 (O_869,N_14077,N_12445);
nand UO_870 (O_870,N_13087,N_12337);
nand UO_871 (O_871,N_14829,N_13206);
nand UO_872 (O_872,N_12757,N_14622);
nand UO_873 (O_873,N_12044,N_12094);
nor UO_874 (O_874,N_12762,N_12313);
and UO_875 (O_875,N_13322,N_12843);
and UO_876 (O_876,N_14876,N_13155);
nor UO_877 (O_877,N_14291,N_14701);
nor UO_878 (O_878,N_14193,N_14529);
or UO_879 (O_879,N_14957,N_14320);
and UO_880 (O_880,N_14354,N_12146);
or UO_881 (O_881,N_13152,N_14844);
nand UO_882 (O_882,N_14223,N_12145);
nor UO_883 (O_883,N_14901,N_13903);
nand UO_884 (O_884,N_13829,N_12294);
and UO_885 (O_885,N_14796,N_12813);
and UO_886 (O_886,N_14523,N_12593);
nor UO_887 (O_887,N_12893,N_12193);
or UO_888 (O_888,N_12705,N_12821);
nor UO_889 (O_889,N_13981,N_14932);
xor UO_890 (O_890,N_14248,N_14012);
nand UO_891 (O_891,N_14625,N_12138);
and UO_892 (O_892,N_12602,N_14341);
nor UO_893 (O_893,N_14824,N_12085);
nor UO_894 (O_894,N_13748,N_14534);
or UO_895 (O_895,N_14307,N_12671);
nand UO_896 (O_896,N_13349,N_12472);
nand UO_897 (O_897,N_12789,N_14633);
nand UO_898 (O_898,N_14723,N_12985);
nand UO_899 (O_899,N_13306,N_13317);
or UO_900 (O_900,N_13460,N_12265);
nand UO_901 (O_901,N_13805,N_13064);
or UO_902 (O_902,N_14974,N_13747);
nand UO_903 (O_903,N_12538,N_12040);
nor UO_904 (O_904,N_12565,N_13767);
nand UO_905 (O_905,N_14322,N_13001);
nor UO_906 (O_906,N_13887,N_14185);
or UO_907 (O_907,N_14603,N_14147);
nor UO_908 (O_908,N_14015,N_14721);
nor UO_909 (O_909,N_13953,N_14437);
nand UO_910 (O_910,N_13715,N_12684);
and UO_911 (O_911,N_14042,N_14554);
or UO_912 (O_912,N_14708,N_13446);
and UO_913 (O_913,N_12290,N_13113);
and UO_914 (O_914,N_12887,N_13512);
nand UO_915 (O_915,N_12548,N_13987);
xor UO_916 (O_916,N_12591,N_14977);
nor UO_917 (O_917,N_14465,N_12814);
or UO_918 (O_918,N_14434,N_14807);
and UO_919 (O_919,N_13074,N_14482);
nand UO_920 (O_920,N_14887,N_13908);
nand UO_921 (O_921,N_13185,N_13582);
or UO_922 (O_922,N_13865,N_12191);
or UO_923 (O_923,N_12399,N_12604);
and UO_924 (O_924,N_13630,N_14840);
or UO_925 (O_925,N_12971,N_13081);
or UO_926 (O_926,N_12597,N_12042);
nor UO_927 (O_927,N_13327,N_13128);
and UO_928 (O_928,N_12732,N_12997);
and UO_929 (O_929,N_13688,N_12698);
or UO_930 (O_930,N_14897,N_14945);
or UO_931 (O_931,N_12412,N_13818);
nor UO_932 (O_932,N_14903,N_12903);
nor UO_933 (O_933,N_14262,N_14583);
or UO_934 (O_934,N_13363,N_14234);
or UO_935 (O_935,N_13666,N_12927);
nor UO_936 (O_936,N_13803,N_12513);
nor UO_937 (O_937,N_12842,N_12616);
nor UO_938 (O_938,N_14406,N_13174);
and UO_939 (O_939,N_12932,N_14070);
nand UO_940 (O_940,N_12330,N_12430);
nor UO_941 (O_941,N_14544,N_14031);
and UO_942 (O_942,N_14118,N_13626);
and UO_943 (O_943,N_13137,N_12632);
nand UO_944 (O_944,N_14065,N_13926);
or UO_945 (O_945,N_12674,N_14725);
nand UO_946 (O_946,N_12452,N_13308);
and UO_947 (O_947,N_12663,N_13375);
nand UO_948 (O_948,N_12305,N_12395);
or UO_949 (O_949,N_12287,N_14804);
nand UO_950 (O_950,N_13988,N_14011);
or UO_951 (O_951,N_12393,N_12005);
or UO_952 (O_952,N_14006,N_12186);
nor UO_953 (O_953,N_14918,N_12809);
nand UO_954 (O_954,N_13641,N_13437);
nor UO_955 (O_955,N_13990,N_12326);
and UO_956 (O_956,N_13885,N_12592);
nor UO_957 (O_957,N_14821,N_13080);
and UO_958 (O_958,N_13837,N_12678);
nand UO_959 (O_959,N_12425,N_13008);
and UO_960 (O_960,N_13632,N_14372);
nand UO_961 (O_961,N_13129,N_13269);
or UO_962 (O_962,N_12629,N_13396);
nand UO_963 (O_963,N_14034,N_12682);
or UO_964 (O_964,N_14279,N_13061);
or UO_965 (O_965,N_14920,N_14332);
nand UO_966 (O_966,N_14132,N_12471);
nor UO_967 (O_967,N_14166,N_14992);
and UO_968 (O_968,N_14232,N_13049);
nand UO_969 (O_969,N_14892,N_12002);
nor UO_970 (O_970,N_12726,N_13241);
nand UO_971 (O_971,N_12799,N_14909);
nor UO_972 (O_972,N_13609,N_13781);
and UO_973 (O_973,N_12849,N_14561);
or UO_974 (O_974,N_13475,N_13568);
nor UO_975 (O_975,N_14385,N_14090);
nor UO_976 (O_976,N_13728,N_13014);
and UO_977 (O_977,N_13922,N_12348);
and UO_978 (O_978,N_13956,N_14289);
xnor UO_979 (O_979,N_14806,N_13940);
nand UO_980 (O_980,N_14149,N_12566);
or UO_981 (O_981,N_12822,N_14068);
and UO_982 (O_982,N_13580,N_12276);
or UO_983 (O_983,N_14593,N_13007);
and UO_984 (O_984,N_12511,N_14048);
nand UO_985 (O_985,N_13045,N_14056);
nand UO_986 (O_986,N_13242,N_13027);
nor UO_987 (O_987,N_13494,N_12864);
nor UO_988 (O_988,N_12482,N_14419);
nor UO_989 (O_989,N_12696,N_13413);
nand UO_990 (O_990,N_12109,N_13863);
nand UO_991 (O_991,N_13684,N_14587);
or UO_992 (O_992,N_14366,N_13291);
and UO_993 (O_993,N_14540,N_13770);
and UO_994 (O_994,N_14639,N_14839);
or UO_995 (O_995,N_13147,N_13330);
and UO_996 (O_996,N_12836,N_13143);
or UO_997 (O_997,N_12829,N_13234);
nor UO_998 (O_998,N_13845,N_14025);
nor UO_999 (O_999,N_13517,N_12487);
nand UO_1000 (O_1000,N_14961,N_14064);
and UO_1001 (O_1001,N_14253,N_14898);
nor UO_1002 (O_1002,N_13165,N_13637);
and UO_1003 (O_1003,N_12883,N_13976);
nand UO_1004 (O_1004,N_13701,N_12967);
nand UO_1005 (O_1005,N_12429,N_14254);
or UO_1006 (O_1006,N_12585,N_13890);
or UO_1007 (O_1007,N_12008,N_14520);
nand UO_1008 (O_1008,N_13123,N_13886);
nand UO_1009 (O_1009,N_14865,N_13720);
and UO_1010 (O_1010,N_12934,N_12206);
nand UO_1011 (O_1011,N_12996,N_13858);
and UO_1012 (O_1012,N_13699,N_14293);
nand UO_1013 (O_1013,N_14119,N_14217);
or UO_1014 (O_1014,N_14956,N_12009);
nand UO_1015 (O_1015,N_12558,N_12553);
nand UO_1016 (O_1016,N_14008,N_13996);
nor UO_1017 (O_1017,N_12121,N_14450);
and UO_1018 (O_1018,N_14302,N_12031);
nor UO_1019 (O_1019,N_14360,N_14299);
and UO_1020 (O_1020,N_13037,N_13560);
or UO_1021 (O_1021,N_13938,N_13833);
or UO_1022 (O_1022,N_12706,N_14552);
and UO_1023 (O_1023,N_14613,N_12712);
and UO_1024 (O_1024,N_12136,N_14857);
nand UO_1025 (O_1025,N_12232,N_12765);
or UO_1026 (O_1026,N_13211,N_13573);
or UO_1027 (O_1027,N_14779,N_14765);
and UO_1028 (O_1028,N_13615,N_12969);
or UO_1029 (O_1029,N_14363,N_13690);
nand UO_1030 (O_1030,N_13335,N_13583);
nor UO_1031 (O_1031,N_13202,N_12128);
or UO_1032 (O_1032,N_12419,N_14059);
or UO_1033 (O_1033,N_13430,N_14511);
or UO_1034 (O_1034,N_12588,N_12784);
nand UO_1035 (O_1035,N_13034,N_12417);
and UO_1036 (O_1036,N_14242,N_12238);
or UO_1037 (O_1037,N_12123,N_13562);
or UO_1038 (O_1038,N_13324,N_14873);
or UO_1039 (O_1039,N_13381,N_14071);
or UO_1040 (O_1040,N_13918,N_12066);
nor UO_1041 (O_1041,N_13017,N_13888);
or UO_1042 (O_1042,N_14421,N_13997);
or UO_1043 (O_1043,N_13444,N_12485);
and UO_1044 (O_1044,N_12617,N_14213);
and UO_1045 (O_1045,N_14888,N_13271);
and UO_1046 (O_1046,N_12129,N_13297);
or UO_1047 (O_1047,N_14879,N_13752);
and UO_1048 (O_1048,N_12941,N_14480);
or UO_1049 (O_1049,N_12856,N_14866);
and UO_1050 (O_1050,N_12961,N_13500);
nor UO_1051 (O_1051,N_14104,N_13547);
nor UO_1052 (O_1052,N_13955,N_14744);
and UO_1053 (O_1053,N_14209,N_12090);
and UO_1054 (O_1054,N_14513,N_14828);
or UO_1055 (O_1055,N_13148,N_12529);
and UO_1056 (O_1056,N_14358,N_13181);
and UO_1057 (O_1057,N_14445,N_13329);
and UO_1058 (O_1058,N_14650,N_13070);
nand UO_1059 (O_1059,N_13332,N_12024);
nor UO_1060 (O_1060,N_14179,N_12672);
nand UO_1061 (O_1061,N_14457,N_14330);
nor UO_1062 (O_1062,N_14621,N_14518);
nand UO_1063 (O_1063,N_13114,N_14321);
nor UO_1064 (O_1064,N_14947,N_13721);
and UO_1065 (O_1065,N_13839,N_13577);
or UO_1066 (O_1066,N_14735,N_14024);
or UO_1067 (O_1067,N_13533,N_12147);
nand UO_1068 (O_1068,N_13273,N_14535);
or UO_1069 (O_1069,N_12205,N_13086);
or UO_1070 (O_1070,N_14852,N_13352);
nand UO_1071 (O_1071,N_13623,N_13005);
and UO_1072 (O_1072,N_13035,N_12976);
and UO_1073 (O_1073,N_14783,N_13032);
xnor UO_1074 (O_1074,N_14697,N_12252);
nor UO_1075 (O_1075,N_13734,N_13553);
nand UO_1076 (O_1076,N_12473,N_13026);
nand UO_1077 (O_1077,N_12907,N_14227);
and UO_1078 (O_1078,N_13116,N_12383);
nand UO_1079 (O_1079,N_13527,N_14867);
and UO_1080 (O_1080,N_12231,N_13101);
and UO_1081 (O_1081,N_14763,N_14195);
nand UO_1082 (O_1082,N_13024,N_13217);
and UO_1083 (O_1083,N_13727,N_13993);
or UO_1084 (O_1084,N_13345,N_13505);
and UO_1085 (O_1085,N_14606,N_14318);
nand UO_1086 (O_1086,N_12469,N_14398);
nand UO_1087 (O_1087,N_14187,N_14754);
or UO_1088 (O_1088,N_13246,N_13343);
or UO_1089 (O_1089,N_14579,N_14230);
nand UO_1090 (O_1090,N_14327,N_14208);
and UO_1091 (O_1091,N_13477,N_14816);
and UO_1092 (O_1092,N_12181,N_12266);
nor UO_1093 (O_1093,N_13333,N_14351);
and UO_1094 (O_1094,N_13871,N_13398);
nand UO_1095 (O_1095,N_13436,N_14811);
or UO_1096 (O_1096,N_12905,N_14646);
or UO_1097 (O_1097,N_13804,N_14110);
nor UO_1098 (O_1098,N_13320,N_14030);
or UO_1099 (O_1099,N_12324,N_13189);
or UO_1100 (O_1100,N_12575,N_12612);
and UO_1101 (O_1101,N_14152,N_12350);
nand UO_1102 (O_1102,N_13664,N_13529);
nand UO_1103 (O_1103,N_14812,N_13453);
nor UO_1104 (O_1104,N_14659,N_13499);
nand UO_1105 (O_1105,N_13935,N_13031);
nand UO_1106 (O_1106,N_12547,N_13745);
or UO_1107 (O_1107,N_12152,N_12051);
and UO_1108 (O_1108,N_13548,N_13433);
nor UO_1109 (O_1109,N_13145,N_13810);
nor UO_1110 (O_1110,N_14080,N_14160);
or UO_1111 (O_1111,N_13581,N_13542);
or UO_1112 (O_1112,N_14381,N_13336);
or UO_1113 (O_1113,N_14813,N_12938);
nor UO_1114 (O_1114,N_13003,N_13762);
nand UO_1115 (O_1115,N_14574,N_12386);
and UO_1116 (O_1116,N_14495,N_14894);
nand UO_1117 (O_1117,N_12528,N_14967);
nor UO_1118 (O_1118,N_12470,N_12119);
nor UO_1119 (O_1119,N_13178,N_14214);
or UO_1120 (O_1120,N_12242,N_12204);
and UO_1121 (O_1121,N_12739,N_14605);
and UO_1122 (O_1122,N_14252,N_14922);
nand UO_1123 (O_1123,N_12984,N_12540);
nor UO_1124 (O_1124,N_13036,N_14389);
and UO_1125 (O_1125,N_13321,N_12504);
and UO_1126 (O_1126,N_12742,N_13759);
nand UO_1127 (O_1127,N_13555,N_13880);
nand UO_1128 (O_1128,N_12935,N_14238);
nand UO_1129 (O_1129,N_13921,N_14528);
nand UO_1130 (O_1130,N_12459,N_14597);
or UO_1131 (O_1131,N_14446,N_13248);
or UO_1132 (O_1132,N_13660,N_12224);
and UO_1133 (O_1133,N_13033,N_14808);
and UO_1134 (O_1134,N_14035,N_13122);
or UO_1135 (O_1135,N_13689,N_12301);
nor UO_1136 (O_1136,N_12240,N_12137);
nor UO_1137 (O_1137,N_12723,N_14925);
and UO_1138 (O_1138,N_12161,N_14091);
or UO_1139 (O_1139,N_14233,N_13389);
nor UO_1140 (O_1140,N_14348,N_13796);
or UO_1141 (O_1141,N_13627,N_12201);
or UO_1142 (O_1142,N_13144,N_13827);
or UO_1143 (O_1143,N_13305,N_13289);
nand UO_1144 (O_1144,N_12312,N_13777);
or UO_1145 (O_1145,N_12316,N_12995);
and UO_1146 (O_1146,N_12222,N_12422);
and UO_1147 (O_1147,N_13230,N_12749);
nor UO_1148 (O_1148,N_14296,N_13002);
or UO_1149 (O_1149,N_12267,N_12584);
nor UO_1150 (O_1150,N_13365,N_13479);
or UO_1151 (O_1151,N_13130,N_13168);
nor UO_1152 (O_1152,N_13267,N_12633);
nand UO_1153 (O_1153,N_12270,N_14144);
nand UO_1154 (O_1154,N_13563,N_12481);
nor UO_1155 (O_1155,N_12391,N_13602);
nand UO_1156 (O_1156,N_13875,N_13200);
nand UO_1157 (O_1157,N_13658,N_12358);
or UO_1158 (O_1158,N_13262,N_13657);
or UO_1159 (O_1159,N_14989,N_13503);
nand UO_1160 (O_1160,N_14274,N_12159);
and UO_1161 (O_1161,N_12216,N_14660);
and UO_1162 (O_1162,N_14375,N_14893);
nand UO_1163 (O_1163,N_12258,N_13315);
or UO_1164 (O_1164,N_14623,N_13992);
nand UO_1165 (O_1165,N_12081,N_13485);
or UO_1166 (O_1166,N_12955,N_13511);
and UO_1167 (O_1167,N_14420,N_13601);
and UO_1168 (O_1168,N_12619,N_14493);
or UO_1169 (O_1169,N_14508,N_13642);
or UO_1170 (O_1170,N_12609,N_13874);
and UO_1171 (O_1171,N_12424,N_12788);
or UO_1172 (O_1172,N_14941,N_13388);
xnor UO_1173 (O_1173,N_14841,N_13497);
or UO_1174 (O_1174,N_13598,N_14300);
or UO_1175 (O_1175,N_13029,N_13736);
nand UO_1176 (O_1176,N_13245,N_14970);
nor UO_1177 (O_1177,N_12763,N_14558);
nand UO_1178 (O_1178,N_14464,N_12023);
nor UO_1179 (O_1179,N_14843,N_12495);
nor UO_1180 (O_1180,N_13456,N_13423);
and UO_1181 (O_1181,N_12126,N_14496);
or UO_1182 (O_1182,N_14294,N_14695);
xnor UO_1183 (O_1183,N_14430,N_14860);
and UO_1184 (O_1184,N_14117,N_13103);
and UO_1185 (O_1185,N_14919,N_14177);
and UO_1186 (O_1186,N_13379,N_12447);
or UO_1187 (O_1187,N_14139,N_14642);
or UO_1188 (O_1188,N_13495,N_14387);
nand UO_1189 (O_1189,N_13102,N_14610);
nand UO_1190 (O_1190,N_14896,N_13019);
nand UO_1191 (O_1191,N_12910,N_12503);
and UO_1192 (O_1192,N_14105,N_14148);
and UO_1193 (O_1193,N_12736,N_13902);
nor UO_1194 (O_1194,N_14766,N_14151);
nor UO_1195 (O_1195,N_12390,N_12086);
or UO_1196 (O_1196,N_12096,N_13518);
and UO_1197 (O_1197,N_13659,N_14319);
and UO_1198 (O_1198,N_14403,N_13405);
nor UO_1199 (O_1199,N_13263,N_14752);
nand UO_1200 (O_1200,N_12132,N_12449);
or UO_1201 (O_1201,N_13831,N_12798);
and UO_1202 (O_1202,N_13967,N_13830);
nor UO_1203 (O_1203,N_14155,N_14971);
and UO_1204 (O_1204,N_13652,N_13295);
nand UO_1205 (O_1205,N_14572,N_12841);
and UO_1206 (O_1206,N_14017,N_13946);
or UO_1207 (O_1207,N_14662,N_14374);
nand UO_1208 (O_1208,N_12179,N_12438);
nor UO_1209 (O_1209,N_12901,N_13610);
or UO_1210 (O_1210,N_14049,N_12990);
and UO_1211 (O_1211,N_14952,N_14594);
nand UO_1212 (O_1212,N_13328,N_12070);
and UO_1213 (O_1213,N_12384,N_14631);
nand UO_1214 (O_1214,N_13443,N_14835);
nand UO_1215 (O_1215,N_14101,N_14966);
or UO_1216 (O_1216,N_14306,N_13836);
nor UO_1217 (O_1217,N_13587,N_13411);
and UO_1218 (O_1218,N_12833,N_12197);
nand UO_1219 (O_1219,N_13420,N_14634);
nor UO_1220 (O_1220,N_12534,N_13772);
or UO_1221 (O_1221,N_12377,N_14917);
nand UO_1222 (O_1222,N_13504,N_14273);
nand UO_1223 (O_1223,N_13742,N_14264);
or UO_1224 (O_1224,N_14673,N_12053);
or UO_1225 (O_1225,N_14007,N_13750);
nand UO_1226 (O_1226,N_12830,N_12494);
or UO_1227 (O_1227,N_12379,N_14965);
nand UO_1228 (O_1228,N_13009,N_12409);
nor UO_1229 (O_1229,N_13053,N_14156);
and UO_1230 (O_1230,N_13929,N_13768);
nand UO_1231 (O_1231,N_14258,N_14196);
xnor UO_1232 (O_1232,N_13125,N_12725);
nand UO_1233 (O_1233,N_12420,N_13589);
xnor UO_1234 (O_1234,N_14257,N_14927);
nand UO_1235 (O_1235,N_12975,N_12756);
nand UO_1236 (O_1236,N_12530,N_14731);
nor UO_1237 (O_1237,N_12563,N_12195);
nor UO_1238 (O_1238,N_13133,N_12332);
nor UO_1239 (O_1239,N_14418,N_14433);
or UO_1240 (O_1240,N_12687,N_13484);
and UO_1241 (O_1241,N_14588,N_12444);
nor UO_1242 (O_1242,N_12580,N_14726);
nor UO_1243 (O_1243,N_12517,N_14449);
nand UO_1244 (O_1244,N_13754,N_12454);
nand UO_1245 (O_1245,N_12225,N_12202);
nor UO_1246 (O_1246,N_13639,N_14362);
nand UO_1247 (O_1247,N_13593,N_14706);
nor UO_1248 (O_1248,N_12392,N_14548);
nor UO_1249 (O_1249,N_13268,N_13537);
nand UO_1250 (O_1250,N_13265,N_12387);
nor UO_1251 (O_1251,N_14585,N_14489);
or UO_1252 (O_1252,N_14938,N_12915);
nand UO_1253 (O_1253,N_12280,N_13112);
nor UO_1254 (O_1254,N_14197,N_14575);
nor UO_1255 (O_1255,N_14830,N_12894);
nand UO_1256 (O_1256,N_13056,N_14809);
or UO_1257 (O_1257,N_14955,N_12164);
nand UO_1258 (O_1258,N_13798,N_12272);
nand UO_1259 (O_1259,N_14693,N_13094);
nor UO_1260 (O_1260,N_14184,N_14431);
and UO_1261 (O_1261,N_12025,N_12178);
or UO_1262 (O_1262,N_14734,N_13585);
and UO_1263 (O_1263,N_14609,N_13448);
or UO_1264 (O_1264,N_13068,N_12960);
and UO_1265 (O_1265,N_12215,N_14280);
nor UO_1266 (O_1266,N_12603,N_13635);
and UO_1267 (O_1267,N_12532,N_12293);
xor UO_1268 (O_1268,N_13188,N_12214);
nand UO_1269 (O_1269,N_12759,N_14355);
or UO_1270 (O_1270,N_13904,N_13814);
nand UO_1271 (O_1271,N_14205,N_12834);
and UO_1272 (O_1272,N_12275,N_14707);
nand UO_1273 (O_1273,N_14454,N_14188);
nand UO_1274 (O_1274,N_13470,N_12586);
nand UO_1275 (O_1275,N_12107,N_13551);
xnor UO_1276 (O_1276,N_14122,N_13065);
and UO_1277 (O_1277,N_13669,N_14116);
nor UO_1278 (O_1278,N_12933,N_14268);
and UO_1279 (O_1279,N_13800,N_13948);
and UO_1280 (O_1280,N_13340,N_13028);
and UO_1281 (O_1281,N_12441,N_13820);
or UO_1282 (O_1282,N_13964,N_12810);
nand UO_1283 (O_1283,N_12646,N_14628);
xor UO_1284 (O_1284,N_13797,N_13786);
nor UO_1285 (O_1285,N_12426,N_13011);
nor UO_1286 (O_1286,N_14647,N_13574);
nor UO_1287 (O_1287,N_14784,N_14180);
nand UO_1288 (O_1288,N_14448,N_12554);
nand UO_1289 (O_1289,N_12076,N_13784);
or UO_1290 (O_1290,N_13675,N_14855);
and UO_1291 (O_1291,N_14228,N_12442);
nand UO_1292 (O_1292,N_13346,N_14770);
nand UO_1293 (O_1293,N_14749,N_13354);
and UO_1294 (O_1294,N_13228,N_12006);
or UO_1295 (O_1295,N_12476,N_14926);
nor UO_1296 (O_1296,N_14539,N_13402);
and UO_1297 (O_1297,N_12261,N_13861);
or UO_1298 (O_1298,N_12539,N_13043);
or UO_1299 (O_1299,N_12857,N_12100);
or UO_1300 (O_1300,N_13369,N_13617);
or UO_1301 (O_1301,N_12692,N_14682);
or UO_1302 (O_1302,N_13072,N_12404);
nand UO_1303 (O_1303,N_13461,N_13853);
and UO_1304 (O_1304,N_14138,N_14097);
nand UO_1305 (O_1305,N_13746,N_14798);
and UO_1306 (O_1306,N_12844,N_14142);
and UO_1307 (O_1307,N_13459,N_12500);
and UO_1308 (O_1308,N_13552,N_14130);
and UO_1309 (O_1309,N_13150,N_13012);
nor UO_1310 (O_1310,N_12474,N_14986);
nor UO_1311 (O_1311,N_14338,N_13501);
nor UO_1312 (O_1312,N_14782,N_13386);
nor UO_1313 (O_1313,N_13709,N_13215);
and UO_1314 (O_1314,N_13047,N_13934);
nor UO_1315 (O_1315,N_12512,N_13445);
nand UO_1316 (O_1316,N_14789,N_14471);
or UO_1317 (O_1317,N_14283,N_13213);
or UO_1318 (O_1318,N_14201,N_14868);
and UO_1319 (O_1319,N_12034,N_13898);
nor UO_1320 (O_1320,N_12797,N_12973);
or UO_1321 (O_1321,N_12106,N_14096);
and UO_1322 (O_1322,N_12781,N_12187);
and UO_1323 (O_1323,N_13439,N_13051);
nand UO_1324 (O_1324,N_12458,N_14315);
nand UO_1325 (O_1325,N_13957,N_12647);
nor UO_1326 (O_1326,N_14194,N_14694);
nand UO_1327 (O_1327,N_12127,N_12800);
or UO_1328 (O_1328,N_12667,N_12439);
and UO_1329 (O_1329,N_14189,N_14486);
nor UO_1330 (O_1330,N_12406,N_14504);
nor UO_1331 (O_1331,N_13847,N_14859);
nor UO_1332 (O_1332,N_12340,N_13543);
nand UO_1333 (O_1333,N_14630,N_13920);
nand UO_1334 (O_1334,N_12777,N_14416);
or UO_1335 (O_1335,N_12030,N_13449);
nand UO_1336 (O_1336,N_13795,N_12203);
and UO_1337 (O_1337,N_13723,N_13347);
or UO_1338 (O_1338,N_14476,N_14044);
and UO_1339 (O_1339,N_14137,N_14468);
nor UO_1340 (O_1340,N_13524,N_13454);
nand UO_1341 (O_1341,N_14455,N_12848);
nand UO_1342 (O_1342,N_12271,N_12717);
and UO_1343 (O_1343,N_14176,N_14384);
nand UO_1344 (O_1344,N_14298,N_13293);
or UO_1345 (O_1345,N_12223,N_13279);
or UO_1346 (O_1346,N_13247,N_12972);
nand UO_1347 (O_1347,N_13862,N_13326);
nor UO_1348 (O_1348,N_12983,N_12436);
or UO_1349 (O_1349,N_14073,N_14173);
and UO_1350 (O_1350,N_14995,N_14339);
nand UO_1351 (O_1351,N_13570,N_12286);
xnor UO_1352 (O_1352,N_14724,N_14817);
nand UO_1353 (O_1353,N_14404,N_14906);
xnor UO_1354 (O_1354,N_14698,N_14713);
nor UO_1355 (O_1355,N_14466,N_14131);
nand UO_1356 (O_1356,N_12653,N_13162);
nand UO_1357 (O_1357,N_12221,N_14183);
and UO_1358 (O_1358,N_12815,N_14484);
nand UO_1359 (O_1359,N_13041,N_12069);
nor UO_1360 (O_1360,N_12959,N_13124);
and UO_1361 (O_1361,N_13407,N_12108);
nand UO_1362 (O_1362,N_13237,N_14020);
nand UO_1363 (O_1363,N_12496,N_12747);
or UO_1364 (O_1364,N_14099,N_14141);
nor UO_1365 (O_1365,N_12227,N_13811);
nor UO_1366 (O_1366,N_14526,N_12236);
and UO_1367 (O_1367,N_13195,N_14463);
nand UO_1368 (O_1368,N_12665,N_13256);
nor UO_1369 (O_1369,N_13578,N_13523);
nor UO_1370 (O_1370,N_12544,N_13760);
and UO_1371 (O_1371,N_13869,N_14703);
nor UO_1372 (O_1372,N_12207,N_12795);
and UO_1373 (O_1373,N_14163,N_12089);
nand UO_1374 (O_1374,N_13808,N_13401);
nand UO_1375 (O_1375,N_13000,N_12735);
or UO_1376 (O_1376,N_12812,N_13605);
and UO_1377 (O_1377,N_13608,N_12914);
or UO_1378 (O_1378,N_13465,N_14267);
nor UO_1379 (O_1379,N_14057,N_13914);
and UO_1380 (O_1380,N_13281,N_14106);
and UO_1381 (O_1381,N_12507,N_12596);
or UO_1382 (O_1382,N_14219,N_14220);
or UO_1383 (O_1383,N_12811,N_14834);
and UO_1384 (O_1384,N_13136,N_14551);
or UO_1385 (O_1385,N_12722,N_14872);
nand UO_1386 (O_1386,N_13060,N_12545);
nor UO_1387 (O_1387,N_14854,N_12226);
nor UO_1388 (O_1388,N_13492,N_13653);
and UO_1389 (O_1389,N_12779,N_13216);
nand UO_1390 (O_1390,N_12628,N_14186);
and UO_1391 (O_1391,N_12263,N_14429);
nor UO_1392 (O_1392,N_14074,N_13409);
and UO_1393 (O_1393,N_13220,N_14235);
nor UO_1394 (O_1394,N_14409,N_14488);
and UO_1395 (O_1395,N_13924,N_14664);
nor UO_1396 (O_1396,N_13586,N_13339);
nand UO_1397 (O_1397,N_13469,N_13121);
or UO_1398 (O_1398,N_14615,N_14975);
and UO_1399 (O_1399,N_13096,N_12104);
nor UO_1400 (O_1400,N_12522,N_13824);
or UO_1401 (O_1401,N_13879,N_14991);
nand UO_1402 (O_1402,N_12556,N_13138);
and UO_1403 (O_1403,N_13793,N_14849);
or UO_1404 (O_1404,N_13749,N_14672);
nor UO_1405 (O_1405,N_12690,N_12840);
nand UO_1406 (O_1406,N_14140,N_14543);
or UO_1407 (O_1407,N_13153,N_13358);
or UO_1408 (O_1408,N_12028,N_12047);
nand UO_1409 (O_1409,N_12396,N_13344);
nand UO_1410 (O_1410,N_13260,N_12929);
nor UO_1411 (O_1411,N_12478,N_13057);
or UO_1412 (O_1412,N_14786,N_13973);
or UO_1413 (O_1413,N_14029,N_14276);
and UO_1414 (O_1414,N_12664,N_13959);
or UO_1415 (O_1415,N_14716,N_14087);
nor UO_1416 (O_1416,N_12579,N_12307);
and UO_1417 (O_1417,N_14226,N_13942);
or UO_1418 (O_1418,N_12059,N_12957);
nor UO_1419 (O_1419,N_14081,N_12752);
xor UO_1420 (O_1420,N_13274,N_12041);
or UO_1421 (O_1421,N_12741,N_14290);
and UO_1422 (O_1422,N_14182,N_13662);
or UO_1423 (O_1423,N_12880,N_14503);
nor UO_1424 (O_1424,N_14699,N_14046);
nor UO_1425 (O_1425,N_14510,N_12940);
nor UO_1426 (O_1426,N_13514,N_14282);
nor UO_1427 (O_1427,N_13873,N_14923);
and UO_1428 (O_1428,N_14473,N_12713);
nand UO_1429 (O_1429,N_13726,N_12414);
nor UO_1430 (O_1430,N_13961,N_14869);
and UO_1431 (O_1431,N_13067,N_13105);
nor UO_1432 (O_1432,N_14312,N_12608);
or UO_1433 (O_1433,N_13239,N_12868);
nand UO_1434 (O_1434,N_12229,N_12292);
and UO_1435 (O_1435,N_13212,N_14285);
or UO_1436 (O_1436,N_12453,N_12962);
or UO_1437 (O_1437,N_12257,N_14549);
nand UO_1438 (O_1438,N_12342,N_14525);
nand UO_1439 (O_1439,N_13951,N_14595);
nand UO_1440 (O_1440,N_13207,N_13506);
nand UO_1441 (O_1441,N_13378,N_13303);
nand UO_1442 (O_1442,N_12531,N_12600);
nand UO_1443 (O_1443,N_13584,N_12693);
nor UO_1444 (O_1444,N_12359,N_13631);
nor UO_1445 (O_1445,N_12120,N_12802);
or UO_1446 (O_1446,N_13079,N_12774);
nand UO_1447 (O_1447,N_12728,N_13374);
nand UO_1448 (O_1448,N_13311,N_12559);
nand UO_1449 (O_1449,N_12598,N_12978);
nor UO_1450 (O_1450,N_12792,N_14153);
or UO_1451 (O_1451,N_13851,N_14063);
nand UO_1452 (O_1452,N_12626,N_13687);
or UO_1453 (O_1453,N_12048,N_13974);
or UO_1454 (O_1454,N_13169,N_12169);
and UO_1455 (O_1455,N_14885,N_12574);
nor UO_1456 (O_1456,N_13572,N_13878);
or UO_1457 (O_1457,N_14972,N_12043);
nand UO_1458 (O_1458,N_13278,N_12149);
and UO_1459 (O_1459,N_12877,N_13085);
nand UO_1460 (O_1460,N_14773,N_12489);
nand UO_1461 (O_1461,N_13361,N_13360);
xor UO_1462 (O_1462,N_12514,N_13127);
nand UO_1463 (O_1463,N_12479,N_13227);
nand UO_1464 (O_1464,N_12902,N_13711);
or UO_1465 (O_1465,N_14402,N_13680);
nand UO_1466 (O_1466,N_12477,N_12074);
nand UO_1467 (O_1467,N_12679,N_12254);
xnor UO_1468 (O_1468,N_13613,N_14556);
nand UO_1469 (O_1469,N_12282,N_13944);
or UO_1470 (O_1470,N_14886,N_13421);
or UO_1471 (O_1471,N_12098,N_13392);
nand UO_1472 (O_1472,N_13052,N_14395);
or UO_1473 (O_1473,N_14568,N_12431);
nor UO_1474 (O_1474,N_14944,N_14061);
nor UO_1475 (O_1475,N_13417,N_13535);
or UO_1476 (O_1476,N_14643,N_12561);
or UO_1477 (O_1477,N_12022,N_14705);
and UO_1478 (O_1478,N_13108,N_14023);
nor UO_1479 (O_1479,N_12838,N_13406);
and UO_1480 (O_1480,N_14769,N_13304);
and UO_1481 (O_1481,N_13486,N_14109);
and UO_1482 (O_1482,N_12247,N_12334);
and UO_1483 (O_1483,N_13775,N_14345);
nand UO_1484 (O_1484,N_13312,N_14933);
nand UO_1485 (O_1485,N_12235,N_12704);
and UO_1486 (O_1486,N_14340,N_14072);
or UO_1487 (O_1487,N_14498,N_14655);
and UO_1488 (O_1488,N_12719,N_14462);
or UO_1489 (O_1489,N_12851,N_12587);
and UO_1490 (O_1490,N_12785,N_12572);
nor UO_1491 (O_1491,N_12865,N_12244);
and UO_1492 (O_1492,N_13917,N_12835);
and UO_1493 (O_1493,N_14093,N_13975);
nand UO_1494 (O_1494,N_13172,N_13342);
nand UO_1495 (O_1495,N_14112,N_13099);
nor UO_1496 (O_1496,N_14325,N_12466);
and UO_1497 (O_1497,N_14505,N_14797);
and UO_1498 (O_1498,N_14668,N_13791);
nand UO_1499 (O_1499,N_12930,N_12319);
nand UO_1500 (O_1500,N_14364,N_13230);
nor UO_1501 (O_1501,N_13644,N_14723);
xnor UO_1502 (O_1502,N_12769,N_13500);
and UO_1503 (O_1503,N_12222,N_12539);
nand UO_1504 (O_1504,N_14412,N_13769);
nor UO_1505 (O_1505,N_13016,N_14654);
or UO_1506 (O_1506,N_13496,N_14143);
and UO_1507 (O_1507,N_14151,N_13051);
nand UO_1508 (O_1508,N_13168,N_14163);
nor UO_1509 (O_1509,N_12452,N_14201);
or UO_1510 (O_1510,N_13594,N_13974);
and UO_1511 (O_1511,N_14478,N_13467);
nand UO_1512 (O_1512,N_14651,N_13367);
nor UO_1513 (O_1513,N_12174,N_12403);
and UO_1514 (O_1514,N_12987,N_14425);
nand UO_1515 (O_1515,N_14270,N_14475);
nor UO_1516 (O_1516,N_12495,N_12669);
and UO_1517 (O_1517,N_13525,N_14440);
nor UO_1518 (O_1518,N_13343,N_14607);
and UO_1519 (O_1519,N_13831,N_13724);
or UO_1520 (O_1520,N_13674,N_13046);
nand UO_1521 (O_1521,N_14145,N_14518);
or UO_1522 (O_1522,N_13707,N_14493);
nand UO_1523 (O_1523,N_14983,N_14400);
nor UO_1524 (O_1524,N_14726,N_14444);
nand UO_1525 (O_1525,N_14598,N_13270);
nand UO_1526 (O_1526,N_14184,N_12878);
and UO_1527 (O_1527,N_13824,N_12464);
xor UO_1528 (O_1528,N_12890,N_14109);
and UO_1529 (O_1529,N_13445,N_14645);
nor UO_1530 (O_1530,N_12307,N_14472);
nand UO_1531 (O_1531,N_13627,N_14038);
or UO_1532 (O_1532,N_14882,N_12235);
nor UO_1533 (O_1533,N_12162,N_14697);
or UO_1534 (O_1534,N_12527,N_14711);
or UO_1535 (O_1535,N_12409,N_14883);
nor UO_1536 (O_1536,N_13805,N_14333);
nor UO_1537 (O_1537,N_14608,N_14939);
and UO_1538 (O_1538,N_14143,N_14499);
and UO_1539 (O_1539,N_12554,N_14590);
nand UO_1540 (O_1540,N_12223,N_13502);
nand UO_1541 (O_1541,N_13529,N_13982);
nor UO_1542 (O_1542,N_13330,N_12471);
nor UO_1543 (O_1543,N_12007,N_14837);
or UO_1544 (O_1544,N_14525,N_14917);
and UO_1545 (O_1545,N_14306,N_12226);
or UO_1546 (O_1546,N_14708,N_14188);
nor UO_1547 (O_1547,N_12504,N_14160);
or UO_1548 (O_1548,N_14552,N_14706);
or UO_1549 (O_1549,N_12372,N_13962);
and UO_1550 (O_1550,N_12385,N_12027);
nand UO_1551 (O_1551,N_12985,N_13151);
nand UO_1552 (O_1552,N_13559,N_12882);
nor UO_1553 (O_1553,N_12898,N_13671);
nand UO_1554 (O_1554,N_12558,N_12611);
nor UO_1555 (O_1555,N_14701,N_14693);
or UO_1556 (O_1556,N_14482,N_12760);
and UO_1557 (O_1557,N_13120,N_12148);
nor UO_1558 (O_1558,N_14649,N_14070);
nand UO_1559 (O_1559,N_12659,N_14027);
and UO_1560 (O_1560,N_13627,N_12926);
nor UO_1561 (O_1561,N_13392,N_12103);
nor UO_1562 (O_1562,N_12785,N_12876);
nand UO_1563 (O_1563,N_12703,N_12719);
nor UO_1564 (O_1564,N_14977,N_14613);
and UO_1565 (O_1565,N_14741,N_14774);
nand UO_1566 (O_1566,N_14964,N_12961);
nor UO_1567 (O_1567,N_13534,N_14480);
and UO_1568 (O_1568,N_12543,N_12716);
or UO_1569 (O_1569,N_12281,N_14900);
nand UO_1570 (O_1570,N_12955,N_14771);
nand UO_1571 (O_1571,N_12409,N_13069);
and UO_1572 (O_1572,N_13339,N_14015);
and UO_1573 (O_1573,N_13726,N_12537);
or UO_1574 (O_1574,N_14751,N_14789);
and UO_1575 (O_1575,N_13444,N_12235);
nand UO_1576 (O_1576,N_14188,N_12642);
nand UO_1577 (O_1577,N_13655,N_12913);
or UO_1578 (O_1578,N_13252,N_12934);
or UO_1579 (O_1579,N_12986,N_12819);
and UO_1580 (O_1580,N_12521,N_14501);
nor UO_1581 (O_1581,N_12478,N_14282);
nor UO_1582 (O_1582,N_12665,N_13737);
and UO_1583 (O_1583,N_13202,N_14438);
nand UO_1584 (O_1584,N_13359,N_13608);
and UO_1585 (O_1585,N_12811,N_12314);
nor UO_1586 (O_1586,N_14680,N_13960);
or UO_1587 (O_1587,N_14889,N_12481);
nand UO_1588 (O_1588,N_14232,N_12418);
and UO_1589 (O_1589,N_12177,N_13453);
nand UO_1590 (O_1590,N_13524,N_14741);
and UO_1591 (O_1591,N_14875,N_13051);
xnor UO_1592 (O_1592,N_13421,N_12896);
nor UO_1593 (O_1593,N_14022,N_14059);
or UO_1594 (O_1594,N_14158,N_14949);
or UO_1595 (O_1595,N_13611,N_12532);
nor UO_1596 (O_1596,N_13758,N_14388);
nor UO_1597 (O_1597,N_13600,N_14884);
or UO_1598 (O_1598,N_13497,N_13091);
or UO_1599 (O_1599,N_14425,N_14600);
and UO_1600 (O_1600,N_12508,N_14711);
and UO_1601 (O_1601,N_12927,N_12700);
nor UO_1602 (O_1602,N_12672,N_13113);
and UO_1603 (O_1603,N_13836,N_12939);
nand UO_1604 (O_1604,N_13438,N_13161);
or UO_1605 (O_1605,N_14790,N_14331);
nor UO_1606 (O_1606,N_14414,N_12207);
nand UO_1607 (O_1607,N_14036,N_14866);
or UO_1608 (O_1608,N_14307,N_13651);
nor UO_1609 (O_1609,N_14155,N_12711);
nand UO_1610 (O_1610,N_14113,N_13343);
or UO_1611 (O_1611,N_14177,N_13820);
or UO_1612 (O_1612,N_13490,N_13187);
nand UO_1613 (O_1613,N_14015,N_13839);
nand UO_1614 (O_1614,N_14241,N_12359);
nand UO_1615 (O_1615,N_14882,N_14450);
nand UO_1616 (O_1616,N_13372,N_14747);
nand UO_1617 (O_1617,N_12352,N_12703);
nor UO_1618 (O_1618,N_13330,N_12746);
nand UO_1619 (O_1619,N_13876,N_14977);
nor UO_1620 (O_1620,N_14258,N_14017);
or UO_1621 (O_1621,N_13480,N_12783);
nand UO_1622 (O_1622,N_14693,N_14927);
nor UO_1623 (O_1623,N_12915,N_13003);
or UO_1624 (O_1624,N_12817,N_12637);
nand UO_1625 (O_1625,N_13696,N_14391);
or UO_1626 (O_1626,N_12904,N_13690);
nand UO_1627 (O_1627,N_14796,N_13756);
and UO_1628 (O_1628,N_14794,N_13083);
or UO_1629 (O_1629,N_14133,N_13335);
nor UO_1630 (O_1630,N_14321,N_14488);
and UO_1631 (O_1631,N_14006,N_12966);
or UO_1632 (O_1632,N_13248,N_13607);
or UO_1633 (O_1633,N_14155,N_14114);
nand UO_1634 (O_1634,N_13117,N_13447);
nor UO_1635 (O_1635,N_12932,N_13649);
and UO_1636 (O_1636,N_13238,N_14308);
and UO_1637 (O_1637,N_14173,N_13126);
nand UO_1638 (O_1638,N_12381,N_12323);
or UO_1639 (O_1639,N_14454,N_13487);
nand UO_1640 (O_1640,N_14858,N_14530);
and UO_1641 (O_1641,N_13749,N_13692);
or UO_1642 (O_1642,N_14421,N_12802);
and UO_1643 (O_1643,N_14589,N_14798);
nor UO_1644 (O_1644,N_14533,N_14331);
or UO_1645 (O_1645,N_13456,N_12680);
and UO_1646 (O_1646,N_12544,N_13345);
or UO_1647 (O_1647,N_13861,N_13949);
or UO_1648 (O_1648,N_12832,N_14857);
nand UO_1649 (O_1649,N_12624,N_14288);
or UO_1650 (O_1650,N_13845,N_13676);
nand UO_1651 (O_1651,N_14013,N_14488);
nor UO_1652 (O_1652,N_13090,N_13195);
and UO_1653 (O_1653,N_14936,N_14241);
and UO_1654 (O_1654,N_14956,N_13172);
and UO_1655 (O_1655,N_12418,N_14720);
and UO_1656 (O_1656,N_14810,N_13553);
nand UO_1657 (O_1657,N_14104,N_12462);
nand UO_1658 (O_1658,N_12043,N_13452);
or UO_1659 (O_1659,N_14415,N_12855);
or UO_1660 (O_1660,N_12961,N_12296);
or UO_1661 (O_1661,N_12804,N_14210);
nand UO_1662 (O_1662,N_13022,N_13171);
nand UO_1663 (O_1663,N_13512,N_14390);
nor UO_1664 (O_1664,N_13222,N_14441);
or UO_1665 (O_1665,N_13845,N_14945);
or UO_1666 (O_1666,N_13345,N_12460);
nor UO_1667 (O_1667,N_13047,N_13101);
nand UO_1668 (O_1668,N_13872,N_14578);
nor UO_1669 (O_1669,N_12132,N_12756);
and UO_1670 (O_1670,N_12806,N_14711);
nor UO_1671 (O_1671,N_12302,N_12450);
nand UO_1672 (O_1672,N_12702,N_12084);
or UO_1673 (O_1673,N_14103,N_13324);
and UO_1674 (O_1674,N_13389,N_14310);
nand UO_1675 (O_1675,N_12963,N_12492);
nand UO_1676 (O_1676,N_14116,N_13363);
nand UO_1677 (O_1677,N_12102,N_14271);
nand UO_1678 (O_1678,N_14704,N_13592);
nand UO_1679 (O_1679,N_13488,N_14212);
xnor UO_1680 (O_1680,N_12819,N_13748);
nor UO_1681 (O_1681,N_14762,N_13534);
and UO_1682 (O_1682,N_12981,N_12531);
nor UO_1683 (O_1683,N_13690,N_14671);
nor UO_1684 (O_1684,N_14250,N_13362);
or UO_1685 (O_1685,N_12864,N_14463);
nor UO_1686 (O_1686,N_12990,N_14362);
nor UO_1687 (O_1687,N_13738,N_13191);
and UO_1688 (O_1688,N_14186,N_13879);
nand UO_1689 (O_1689,N_12206,N_13926);
xor UO_1690 (O_1690,N_14844,N_13745);
or UO_1691 (O_1691,N_13554,N_14451);
and UO_1692 (O_1692,N_12718,N_13022);
nor UO_1693 (O_1693,N_14020,N_13620);
or UO_1694 (O_1694,N_13272,N_14734);
nor UO_1695 (O_1695,N_12580,N_14781);
or UO_1696 (O_1696,N_12067,N_12273);
and UO_1697 (O_1697,N_13818,N_14936);
nor UO_1698 (O_1698,N_12153,N_12754);
and UO_1699 (O_1699,N_12366,N_12379);
and UO_1700 (O_1700,N_14604,N_12999);
nor UO_1701 (O_1701,N_14791,N_13548);
and UO_1702 (O_1702,N_14768,N_13720);
and UO_1703 (O_1703,N_13861,N_12057);
and UO_1704 (O_1704,N_13242,N_12639);
nor UO_1705 (O_1705,N_14362,N_12182);
and UO_1706 (O_1706,N_12364,N_13453);
or UO_1707 (O_1707,N_14144,N_13756);
and UO_1708 (O_1708,N_14599,N_14699);
nand UO_1709 (O_1709,N_12198,N_12642);
nor UO_1710 (O_1710,N_13269,N_13012);
nand UO_1711 (O_1711,N_14052,N_13760);
and UO_1712 (O_1712,N_13403,N_12052);
nand UO_1713 (O_1713,N_13892,N_12701);
nor UO_1714 (O_1714,N_14260,N_12453);
and UO_1715 (O_1715,N_14053,N_12491);
nor UO_1716 (O_1716,N_14925,N_12727);
nor UO_1717 (O_1717,N_14514,N_13958);
nand UO_1718 (O_1718,N_13538,N_14789);
nand UO_1719 (O_1719,N_13577,N_13087);
nor UO_1720 (O_1720,N_12913,N_14256);
nor UO_1721 (O_1721,N_13500,N_13918);
or UO_1722 (O_1722,N_13775,N_14894);
and UO_1723 (O_1723,N_12591,N_14199);
nor UO_1724 (O_1724,N_14860,N_12660);
and UO_1725 (O_1725,N_14704,N_12377);
and UO_1726 (O_1726,N_14567,N_12781);
nor UO_1727 (O_1727,N_12261,N_14520);
nor UO_1728 (O_1728,N_13796,N_13843);
and UO_1729 (O_1729,N_14859,N_13796);
nand UO_1730 (O_1730,N_14818,N_13450);
nor UO_1731 (O_1731,N_14938,N_13537);
nand UO_1732 (O_1732,N_14126,N_12627);
or UO_1733 (O_1733,N_14474,N_13932);
and UO_1734 (O_1734,N_12627,N_14052);
and UO_1735 (O_1735,N_13703,N_13793);
and UO_1736 (O_1736,N_14568,N_14910);
nor UO_1737 (O_1737,N_14100,N_14335);
nor UO_1738 (O_1738,N_14160,N_14728);
nand UO_1739 (O_1739,N_14583,N_12096);
nand UO_1740 (O_1740,N_13002,N_12166);
and UO_1741 (O_1741,N_13913,N_13818);
or UO_1742 (O_1742,N_14966,N_12467);
nor UO_1743 (O_1743,N_14541,N_14453);
xor UO_1744 (O_1744,N_12650,N_14723);
or UO_1745 (O_1745,N_14515,N_13723);
or UO_1746 (O_1746,N_12725,N_12771);
nor UO_1747 (O_1747,N_13063,N_13862);
or UO_1748 (O_1748,N_13172,N_14619);
or UO_1749 (O_1749,N_14990,N_14222);
and UO_1750 (O_1750,N_13053,N_13814);
nand UO_1751 (O_1751,N_14082,N_13001);
nand UO_1752 (O_1752,N_13447,N_14457);
nand UO_1753 (O_1753,N_13543,N_14665);
nor UO_1754 (O_1754,N_12355,N_14903);
nand UO_1755 (O_1755,N_13812,N_12849);
or UO_1756 (O_1756,N_14138,N_14679);
nand UO_1757 (O_1757,N_13714,N_14827);
nand UO_1758 (O_1758,N_13913,N_14657);
or UO_1759 (O_1759,N_13411,N_14318);
or UO_1760 (O_1760,N_13261,N_12535);
and UO_1761 (O_1761,N_14525,N_12879);
nor UO_1762 (O_1762,N_12493,N_14445);
or UO_1763 (O_1763,N_12583,N_13079);
nor UO_1764 (O_1764,N_14226,N_14767);
and UO_1765 (O_1765,N_13432,N_12643);
and UO_1766 (O_1766,N_14676,N_14261);
and UO_1767 (O_1767,N_13359,N_14454);
or UO_1768 (O_1768,N_14856,N_13964);
nand UO_1769 (O_1769,N_12049,N_14016);
nor UO_1770 (O_1770,N_14560,N_12404);
nand UO_1771 (O_1771,N_14917,N_14254);
or UO_1772 (O_1772,N_13774,N_14746);
nand UO_1773 (O_1773,N_12708,N_14397);
nor UO_1774 (O_1774,N_13829,N_12944);
nor UO_1775 (O_1775,N_14494,N_14742);
and UO_1776 (O_1776,N_12140,N_13674);
or UO_1777 (O_1777,N_12095,N_12203);
nor UO_1778 (O_1778,N_13847,N_14573);
or UO_1779 (O_1779,N_13685,N_13029);
and UO_1780 (O_1780,N_14762,N_14162);
and UO_1781 (O_1781,N_12984,N_13507);
nor UO_1782 (O_1782,N_14806,N_14062);
nor UO_1783 (O_1783,N_13475,N_13409);
nand UO_1784 (O_1784,N_12568,N_14439);
and UO_1785 (O_1785,N_13169,N_13619);
nand UO_1786 (O_1786,N_13006,N_13762);
or UO_1787 (O_1787,N_13066,N_12224);
and UO_1788 (O_1788,N_13439,N_12813);
nand UO_1789 (O_1789,N_14754,N_12710);
nand UO_1790 (O_1790,N_14774,N_12770);
or UO_1791 (O_1791,N_12435,N_12416);
and UO_1792 (O_1792,N_14238,N_14246);
and UO_1793 (O_1793,N_12454,N_12230);
and UO_1794 (O_1794,N_13850,N_13636);
nand UO_1795 (O_1795,N_13339,N_13620);
nand UO_1796 (O_1796,N_14165,N_14056);
or UO_1797 (O_1797,N_12493,N_12125);
or UO_1798 (O_1798,N_12643,N_14584);
nor UO_1799 (O_1799,N_12045,N_14601);
and UO_1800 (O_1800,N_13220,N_12081);
and UO_1801 (O_1801,N_13846,N_14167);
nor UO_1802 (O_1802,N_14472,N_13430);
nor UO_1803 (O_1803,N_13260,N_13118);
nand UO_1804 (O_1804,N_13385,N_14751);
nor UO_1805 (O_1805,N_14139,N_14941);
nor UO_1806 (O_1806,N_13948,N_12458);
or UO_1807 (O_1807,N_12117,N_13508);
nor UO_1808 (O_1808,N_13963,N_14264);
nand UO_1809 (O_1809,N_12862,N_14351);
or UO_1810 (O_1810,N_12366,N_14209);
nor UO_1811 (O_1811,N_13890,N_14682);
nand UO_1812 (O_1812,N_14573,N_13986);
and UO_1813 (O_1813,N_12945,N_14120);
or UO_1814 (O_1814,N_12435,N_13242);
nor UO_1815 (O_1815,N_13016,N_13620);
xor UO_1816 (O_1816,N_12288,N_12356);
nor UO_1817 (O_1817,N_13037,N_13243);
nor UO_1818 (O_1818,N_12443,N_12241);
or UO_1819 (O_1819,N_14473,N_13661);
nand UO_1820 (O_1820,N_13194,N_12195);
xor UO_1821 (O_1821,N_12618,N_13440);
nor UO_1822 (O_1822,N_13191,N_14932);
or UO_1823 (O_1823,N_13043,N_14350);
nor UO_1824 (O_1824,N_12734,N_14876);
nor UO_1825 (O_1825,N_14487,N_13805);
and UO_1826 (O_1826,N_12508,N_14200);
or UO_1827 (O_1827,N_14903,N_12591);
or UO_1828 (O_1828,N_14709,N_14373);
nor UO_1829 (O_1829,N_13514,N_12860);
nand UO_1830 (O_1830,N_12710,N_14450);
nand UO_1831 (O_1831,N_12074,N_12788);
and UO_1832 (O_1832,N_12782,N_12646);
and UO_1833 (O_1833,N_12066,N_12728);
or UO_1834 (O_1834,N_13586,N_12215);
and UO_1835 (O_1835,N_14133,N_14168);
and UO_1836 (O_1836,N_14573,N_13844);
and UO_1837 (O_1837,N_13257,N_12097);
or UO_1838 (O_1838,N_13388,N_12414);
nand UO_1839 (O_1839,N_12574,N_13500);
nand UO_1840 (O_1840,N_14126,N_14068);
and UO_1841 (O_1841,N_14649,N_14662);
nand UO_1842 (O_1842,N_12649,N_14749);
or UO_1843 (O_1843,N_14943,N_14203);
and UO_1844 (O_1844,N_14513,N_13315);
or UO_1845 (O_1845,N_13205,N_13177);
and UO_1846 (O_1846,N_12612,N_14830);
nor UO_1847 (O_1847,N_13725,N_12791);
and UO_1848 (O_1848,N_12781,N_12701);
nand UO_1849 (O_1849,N_12638,N_14864);
xnor UO_1850 (O_1850,N_12225,N_14510);
nand UO_1851 (O_1851,N_12863,N_13034);
nand UO_1852 (O_1852,N_13746,N_12162);
nand UO_1853 (O_1853,N_13180,N_14673);
or UO_1854 (O_1854,N_13104,N_12568);
nor UO_1855 (O_1855,N_14271,N_14240);
nor UO_1856 (O_1856,N_14204,N_14405);
nand UO_1857 (O_1857,N_12193,N_14524);
nor UO_1858 (O_1858,N_14026,N_12798);
and UO_1859 (O_1859,N_12438,N_13199);
nand UO_1860 (O_1860,N_14607,N_14006);
and UO_1861 (O_1861,N_13735,N_14754);
and UO_1862 (O_1862,N_13402,N_12781);
or UO_1863 (O_1863,N_14253,N_12672);
and UO_1864 (O_1864,N_13906,N_14894);
or UO_1865 (O_1865,N_13206,N_14097);
nor UO_1866 (O_1866,N_13820,N_14845);
nor UO_1867 (O_1867,N_14923,N_13526);
nor UO_1868 (O_1868,N_13984,N_13326);
nor UO_1869 (O_1869,N_12496,N_13524);
and UO_1870 (O_1870,N_14933,N_13132);
nor UO_1871 (O_1871,N_13632,N_13373);
nor UO_1872 (O_1872,N_12956,N_14032);
nand UO_1873 (O_1873,N_13731,N_12896);
and UO_1874 (O_1874,N_13290,N_13711);
nand UO_1875 (O_1875,N_14186,N_12830);
or UO_1876 (O_1876,N_13672,N_12257);
nor UO_1877 (O_1877,N_12933,N_14373);
or UO_1878 (O_1878,N_13326,N_14612);
nand UO_1879 (O_1879,N_13751,N_12927);
nor UO_1880 (O_1880,N_13893,N_14674);
or UO_1881 (O_1881,N_14312,N_13779);
and UO_1882 (O_1882,N_13763,N_12759);
nand UO_1883 (O_1883,N_12525,N_13437);
xor UO_1884 (O_1884,N_12607,N_13989);
nand UO_1885 (O_1885,N_12417,N_14318);
or UO_1886 (O_1886,N_14766,N_13912);
and UO_1887 (O_1887,N_12447,N_14157);
xnor UO_1888 (O_1888,N_14083,N_14214);
or UO_1889 (O_1889,N_14875,N_12011);
and UO_1890 (O_1890,N_13602,N_12845);
nor UO_1891 (O_1891,N_12871,N_14260);
or UO_1892 (O_1892,N_12958,N_14505);
nor UO_1893 (O_1893,N_12836,N_13687);
nand UO_1894 (O_1894,N_12402,N_12473);
nand UO_1895 (O_1895,N_13159,N_13953);
and UO_1896 (O_1896,N_13799,N_12776);
and UO_1897 (O_1897,N_13603,N_13119);
nand UO_1898 (O_1898,N_14625,N_12880);
nor UO_1899 (O_1899,N_14805,N_12661);
or UO_1900 (O_1900,N_13776,N_13711);
nor UO_1901 (O_1901,N_13258,N_14961);
nand UO_1902 (O_1902,N_13151,N_14062);
and UO_1903 (O_1903,N_14608,N_13067);
nor UO_1904 (O_1904,N_13878,N_14780);
or UO_1905 (O_1905,N_13729,N_14506);
and UO_1906 (O_1906,N_12658,N_13983);
nand UO_1907 (O_1907,N_13792,N_12423);
and UO_1908 (O_1908,N_14015,N_13789);
nor UO_1909 (O_1909,N_14071,N_12806);
nand UO_1910 (O_1910,N_14600,N_13909);
and UO_1911 (O_1911,N_14813,N_13161);
nor UO_1912 (O_1912,N_12629,N_12654);
or UO_1913 (O_1913,N_13098,N_12317);
and UO_1914 (O_1914,N_14622,N_12899);
or UO_1915 (O_1915,N_14378,N_14254);
nor UO_1916 (O_1916,N_14078,N_14743);
or UO_1917 (O_1917,N_12835,N_14410);
and UO_1918 (O_1918,N_13220,N_12999);
and UO_1919 (O_1919,N_12253,N_14742);
nand UO_1920 (O_1920,N_12556,N_12186);
and UO_1921 (O_1921,N_12823,N_13114);
nor UO_1922 (O_1922,N_12118,N_14042);
and UO_1923 (O_1923,N_14810,N_12673);
and UO_1924 (O_1924,N_13741,N_12042);
and UO_1925 (O_1925,N_12397,N_13906);
nor UO_1926 (O_1926,N_13006,N_14770);
nor UO_1927 (O_1927,N_12405,N_13988);
nor UO_1928 (O_1928,N_14377,N_14967);
or UO_1929 (O_1929,N_12665,N_13743);
nor UO_1930 (O_1930,N_12663,N_12588);
nor UO_1931 (O_1931,N_13767,N_14978);
or UO_1932 (O_1932,N_13786,N_12423);
and UO_1933 (O_1933,N_13648,N_14217);
or UO_1934 (O_1934,N_13550,N_14850);
nand UO_1935 (O_1935,N_14889,N_12242);
nor UO_1936 (O_1936,N_13468,N_13763);
and UO_1937 (O_1937,N_12226,N_13786);
nor UO_1938 (O_1938,N_13060,N_13904);
nand UO_1939 (O_1939,N_13718,N_12007);
and UO_1940 (O_1940,N_14306,N_14872);
and UO_1941 (O_1941,N_14733,N_13895);
nand UO_1942 (O_1942,N_13793,N_12418);
nor UO_1943 (O_1943,N_12408,N_13490);
nor UO_1944 (O_1944,N_14675,N_12253);
nand UO_1945 (O_1945,N_12024,N_13843);
nand UO_1946 (O_1946,N_12579,N_14237);
nand UO_1947 (O_1947,N_14909,N_14005);
nand UO_1948 (O_1948,N_14797,N_14265);
and UO_1949 (O_1949,N_13772,N_14658);
nand UO_1950 (O_1950,N_14070,N_14987);
nor UO_1951 (O_1951,N_12825,N_13205);
or UO_1952 (O_1952,N_13257,N_14323);
and UO_1953 (O_1953,N_14619,N_13863);
and UO_1954 (O_1954,N_14931,N_13876);
or UO_1955 (O_1955,N_13068,N_12398);
nor UO_1956 (O_1956,N_12974,N_13133);
or UO_1957 (O_1957,N_14465,N_12089);
nor UO_1958 (O_1958,N_13194,N_12069);
nand UO_1959 (O_1959,N_13658,N_14701);
and UO_1960 (O_1960,N_13565,N_14286);
nand UO_1961 (O_1961,N_14919,N_14280);
or UO_1962 (O_1962,N_12516,N_13963);
and UO_1963 (O_1963,N_12935,N_13126);
and UO_1964 (O_1964,N_12611,N_12213);
or UO_1965 (O_1965,N_14496,N_12740);
and UO_1966 (O_1966,N_13207,N_13768);
nor UO_1967 (O_1967,N_14265,N_13809);
or UO_1968 (O_1968,N_12246,N_14658);
nand UO_1969 (O_1969,N_14319,N_14658);
nor UO_1970 (O_1970,N_14409,N_12604);
and UO_1971 (O_1971,N_12285,N_13608);
nor UO_1972 (O_1972,N_13120,N_12913);
and UO_1973 (O_1973,N_13432,N_12369);
nand UO_1974 (O_1974,N_14998,N_14626);
or UO_1975 (O_1975,N_12673,N_12983);
or UO_1976 (O_1976,N_12520,N_13643);
nor UO_1977 (O_1977,N_14791,N_12764);
or UO_1978 (O_1978,N_14551,N_14628);
and UO_1979 (O_1979,N_12984,N_14716);
and UO_1980 (O_1980,N_14275,N_13602);
or UO_1981 (O_1981,N_13434,N_13911);
nand UO_1982 (O_1982,N_13552,N_13324);
nor UO_1983 (O_1983,N_14646,N_12659);
nand UO_1984 (O_1984,N_13417,N_14762);
nor UO_1985 (O_1985,N_14642,N_12561);
nor UO_1986 (O_1986,N_12240,N_13741);
nor UO_1987 (O_1987,N_12760,N_13382);
nand UO_1988 (O_1988,N_14658,N_13214);
or UO_1989 (O_1989,N_13345,N_14925);
and UO_1990 (O_1990,N_12998,N_12915);
and UO_1991 (O_1991,N_12612,N_12758);
and UO_1992 (O_1992,N_12864,N_12959);
or UO_1993 (O_1993,N_14157,N_12905);
nor UO_1994 (O_1994,N_12211,N_13599);
nand UO_1995 (O_1995,N_13651,N_14163);
and UO_1996 (O_1996,N_13074,N_13137);
nor UO_1997 (O_1997,N_14687,N_12191);
nor UO_1998 (O_1998,N_12113,N_12807);
and UO_1999 (O_1999,N_12665,N_12880);
endmodule