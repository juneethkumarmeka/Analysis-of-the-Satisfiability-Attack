module basic_2500_25000_3000_8_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1693,In_979);
xnor U1 (N_1,In_1521,In_2445);
xor U2 (N_2,In_946,In_1114);
xor U3 (N_3,In_1835,In_1143);
nand U4 (N_4,In_747,In_1604);
or U5 (N_5,In_1821,In_2408);
nand U6 (N_6,In_96,In_511);
and U7 (N_7,In_1144,In_2413);
nor U8 (N_8,In_1433,In_1776);
xnor U9 (N_9,In_1415,In_919);
nand U10 (N_10,In_1036,In_1469);
nor U11 (N_11,In_872,In_1319);
and U12 (N_12,In_1123,In_1357);
and U13 (N_13,In_421,In_150);
and U14 (N_14,In_2245,In_443);
or U15 (N_15,In_1261,In_557);
nor U16 (N_16,In_2183,In_742);
nor U17 (N_17,In_1071,In_1119);
nor U18 (N_18,In_627,In_101);
nand U19 (N_19,In_503,In_126);
nor U20 (N_20,In_1789,In_1309);
and U21 (N_21,In_2456,In_1287);
nor U22 (N_22,In_1109,In_1690);
or U23 (N_23,In_1644,In_2010);
nand U24 (N_24,In_633,In_1010);
or U25 (N_25,In_1524,In_493);
and U26 (N_26,In_2381,In_1640);
nand U27 (N_27,In_305,In_188);
xnor U28 (N_28,In_423,In_2067);
or U29 (N_29,In_482,In_894);
nand U30 (N_30,In_2475,In_1950);
nor U31 (N_31,In_2492,In_518);
and U32 (N_32,In_1273,In_2056);
xnor U33 (N_33,In_996,In_1705);
xor U34 (N_34,In_1592,In_1031);
and U35 (N_35,In_1933,In_1752);
xor U36 (N_36,In_1435,In_2231);
or U37 (N_37,In_335,In_217);
nor U38 (N_38,In_1317,In_1778);
or U39 (N_39,In_2353,In_146);
nand U40 (N_40,In_137,In_2359);
nor U41 (N_41,In_1003,In_1782);
or U42 (N_42,In_172,In_1019);
nand U43 (N_43,In_60,In_294);
nor U44 (N_44,In_2187,In_1695);
and U45 (N_45,In_981,In_1509);
xor U46 (N_46,In_958,In_1713);
and U47 (N_47,In_77,In_484);
nor U48 (N_48,In_2491,In_1994);
or U49 (N_49,In_131,In_2434);
xor U50 (N_50,In_1256,In_688);
nand U51 (N_51,In_1140,In_569);
nand U52 (N_52,In_878,In_1804);
and U53 (N_53,In_1476,In_821);
nor U54 (N_54,In_689,In_291);
nand U55 (N_55,In_1651,In_574);
or U56 (N_56,In_1955,In_247);
nand U57 (N_57,In_3,In_2029);
nor U58 (N_58,In_542,In_1969);
or U59 (N_59,In_973,In_1661);
and U60 (N_60,In_893,In_1952);
and U61 (N_61,In_1602,In_865);
or U62 (N_62,In_200,In_42);
or U63 (N_63,In_143,In_580);
nor U64 (N_64,In_1126,In_1217);
xor U65 (N_65,In_798,In_233);
nand U66 (N_66,In_2054,In_2440);
xor U67 (N_67,In_70,In_1596);
xnor U68 (N_68,In_869,In_554);
or U69 (N_69,In_1953,In_382);
or U70 (N_70,In_912,In_2454);
nand U71 (N_71,In_2298,In_1248);
or U72 (N_72,In_277,In_1872);
or U73 (N_73,In_2007,In_249);
xor U74 (N_74,In_1671,In_1079);
nor U75 (N_75,In_598,In_2487);
nand U76 (N_76,In_1424,In_1342);
and U77 (N_77,In_152,In_1910);
nand U78 (N_78,In_1384,In_750);
or U79 (N_79,In_506,In_279);
or U80 (N_80,In_221,In_161);
xnor U81 (N_81,In_1853,In_1489);
xor U82 (N_82,In_1797,In_1743);
or U83 (N_83,In_1862,In_1715);
xnor U84 (N_84,In_83,In_2105);
and U85 (N_85,In_2156,In_1701);
xnor U86 (N_86,In_134,In_2136);
or U87 (N_87,In_1292,In_193);
or U88 (N_88,In_1523,In_942);
nor U89 (N_89,In_677,In_2091);
nor U90 (N_90,In_165,In_1992);
nand U91 (N_91,In_424,In_2320);
xor U92 (N_92,In_280,In_2024);
or U93 (N_93,In_470,In_1293);
and U94 (N_94,In_2036,In_1462);
and U95 (N_95,In_2318,In_1762);
nand U96 (N_96,In_899,In_2297);
nand U97 (N_97,In_810,In_2377);
and U98 (N_98,In_1381,In_1007);
xor U99 (N_99,In_1152,In_2490);
nand U100 (N_100,In_1423,In_1628);
nand U101 (N_101,In_1400,In_100);
xnor U102 (N_102,In_2040,In_242);
and U103 (N_103,In_1444,In_1147);
xor U104 (N_104,In_517,In_1078);
xnor U105 (N_105,In_357,In_1888);
or U106 (N_106,In_1482,In_1339);
nor U107 (N_107,In_2370,In_1709);
xor U108 (N_108,In_2399,In_921);
or U109 (N_109,In_548,In_222);
and U110 (N_110,In_1497,In_2210);
nor U111 (N_111,In_1788,In_1474);
nand U112 (N_112,In_532,In_1260);
xor U113 (N_113,In_2104,In_553);
nand U114 (N_114,In_779,In_2261);
nor U115 (N_115,In_204,In_109);
and U116 (N_116,In_1304,In_863);
nand U117 (N_117,In_685,In_1407);
xor U118 (N_118,In_2484,In_130);
or U119 (N_119,In_2186,In_330);
nor U120 (N_120,In_446,In_449);
xnor U121 (N_121,In_360,In_1106);
nand U122 (N_122,In_1843,In_410);
nor U123 (N_123,In_1277,In_792);
or U124 (N_124,In_2071,In_1911);
nor U125 (N_125,In_563,In_1092);
nand U126 (N_126,In_1577,In_1494);
nand U127 (N_127,In_908,In_1070);
nand U128 (N_128,In_670,In_611);
nand U129 (N_129,In_616,In_1131);
xor U130 (N_130,In_1685,In_2066);
xnor U131 (N_131,In_412,In_1457);
nor U132 (N_132,In_1822,In_232);
nand U133 (N_133,In_1014,In_751);
and U134 (N_134,In_2425,In_1168);
or U135 (N_135,In_1421,In_2122);
xor U136 (N_136,In_2039,In_2444);
and U137 (N_137,In_2006,In_2436);
xnor U138 (N_138,In_1607,In_1894);
xor U139 (N_139,In_1191,In_2148);
nand U140 (N_140,In_195,In_832);
nor U141 (N_141,In_1166,In_2367);
or U142 (N_142,In_883,In_1241);
and U143 (N_143,In_92,In_1848);
nor U144 (N_144,In_2455,In_21);
and U145 (N_145,In_720,In_1923);
nor U146 (N_146,In_986,In_1365);
xnor U147 (N_147,In_643,In_1328);
or U148 (N_148,In_1707,In_1321);
and U149 (N_149,In_1528,In_1593);
and U150 (N_150,In_1380,In_1811);
or U151 (N_151,In_669,In_2383);
nand U152 (N_152,In_331,In_1186);
or U153 (N_153,In_80,In_884);
xnor U154 (N_154,In_464,In_2275);
xor U155 (N_155,In_2235,In_50);
and U156 (N_156,In_1032,In_2258);
nand U157 (N_157,In_61,In_966);
and U158 (N_158,In_2457,In_771);
nand U159 (N_159,In_733,In_458);
or U160 (N_160,In_2358,In_234);
xnor U161 (N_161,In_839,In_2131);
nor U162 (N_162,In_1398,In_1945);
and U163 (N_163,In_2098,In_1912);
nor U164 (N_164,In_1039,In_699);
and U165 (N_165,In_1647,In_1883);
and U166 (N_166,In_1930,In_135);
or U167 (N_167,In_2461,In_1943);
or U168 (N_168,In_45,In_584);
xor U169 (N_169,In_682,In_1845);
nor U170 (N_170,In_1688,In_1879);
nor U171 (N_171,In_708,In_1765);
and U172 (N_172,In_1857,In_793);
nor U173 (N_173,In_2124,In_620);
or U174 (N_174,In_497,In_2315);
xor U175 (N_175,In_1730,In_1868);
nor U176 (N_176,In_2017,In_229);
nor U177 (N_177,In_860,In_911);
nand U178 (N_178,In_2157,In_1597);
or U179 (N_179,In_1040,In_2253);
nand U180 (N_180,In_649,In_686);
and U181 (N_181,In_144,In_2169);
or U182 (N_182,In_1089,In_952);
and U183 (N_183,In_253,In_1138);
and U184 (N_184,In_430,In_1153);
nor U185 (N_185,In_1033,In_213);
nand U186 (N_186,In_822,In_2309);
nor U187 (N_187,In_2099,In_2155);
or U188 (N_188,In_1714,In_1649);
nor U189 (N_189,In_1145,In_466);
or U190 (N_190,In_1749,In_2119);
or U191 (N_191,In_1758,In_254);
nand U192 (N_192,In_334,In_1500);
xnor U193 (N_193,In_1043,In_1815);
or U194 (N_194,In_1030,In_1322);
nand U195 (N_195,In_93,In_235);
nor U196 (N_196,In_715,In_2174);
nor U197 (N_197,In_2372,In_1265);
xnor U198 (N_198,In_2076,In_653);
nor U199 (N_199,In_1814,In_1227);
xor U200 (N_200,In_314,In_385);
xor U201 (N_201,In_1909,In_214);
nor U202 (N_202,In_1669,In_1420);
nor U203 (N_203,In_273,In_614);
or U204 (N_204,In_1100,In_704);
xor U205 (N_205,In_1276,In_1733);
nor U206 (N_206,In_407,In_49);
nand U207 (N_207,In_1794,In_240);
or U208 (N_208,In_748,In_1545);
nand U209 (N_209,In_1860,In_887);
nor U210 (N_210,In_712,In_1452);
nor U211 (N_211,In_795,In_319);
and U212 (N_212,In_1183,In_2321);
or U213 (N_213,In_1613,In_1583);
and U214 (N_214,In_1130,In_370);
and U215 (N_215,In_898,In_376);
and U216 (N_216,In_1171,In_1581);
xor U217 (N_217,In_2121,In_72);
xor U218 (N_218,In_73,In_1691);
xnor U219 (N_219,In_393,In_2250);
xor U220 (N_220,In_586,In_1871);
or U221 (N_221,In_837,In_361);
and U222 (N_222,In_1847,In_1345);
xnor U223 (N_223,In_1696,In_1884);
and U224 (N_224,In_909,In_320);
nand U225 (N_225,In_774,In_260);
or U226 (N_226,In_1618,In_1137);
or U227 (N_227,In_626,In_64);
nor U228 (N_228,In_1591,In_1799);
xnor U229 (N_229,In_641,In_1018);
nor U230 (N_230,In_182,In_834);
nand U231 (N_231,In_198,In_2489);
nor U232 (N_232,In_2366,In_1175);
nand U233 (N_233,In_2172,In_882);
and U234 (N_234,In_787,In_1364);
and U235 (N_235,In_91,In_1989);
nand U236 (N_236,In_1934,In_2181);
xnor U237 (N_237,In_638,In_1718);
nor U238 (N_238,In_1742,In_1937);
or U239 (N_239,In_2403,In_1478);
xor U240 (N_240,In_749,In_66);
or U241 (N_241,In_270,In_731);
and U242 (N_242,In_1488,In_2483);
or U243 (N_243,In_468,In_1997);
nand U244 (N_244,In_1578,In_190);
xnor U245 (N_245,In_1247,In_230);
xnor U246 (N_246,In_125,In_2343);
nor U247 (N_247,In_1072,In_22);
nor U248 (N_248,In_426,In_1629);
or U249 (N_249,In_902,In_702);
or U250 (N_250,In_1262,In_197);
nand U251 (N_251,In_2162,In_1731);
and U252 (N_252,In_1959,In_1284);
and U253 (N_253,In_2223,In_692);
nand U254 (N_254,In_2474,In_917);
xor U255 (N_255,In_711,In_1235);
nor U256 (N_256,In_1326,In_2429);
nor U257 (N_257,In_791,In_495);
nor U258 (N_258,In_2341,In_807);
or U259 (N_259,In_414,In_889);
or U260 (N_260,In_1603,In_1267);
nand U261 (N_261,In_1812,In_2432);
nand U262 (N_262,In_1517,In_1954);
nor U263 (N_263,In_1568,In_2476);
and U264 (N_264,In_1791,In_610);
nand U265 (N_265,In_2147,In_514);
nand U266 (N_266,In_1729,In_2179);
nor U267 (N_267,In_1113,In_2171);
nand U268 (N_268,In_1639,In_2276);
and U269 (N_269,In_350,In_1826);
xor U270 (N_270,In_2000,In_1116);
xnor U271 (N_271,In_241,In_338);
xor U272 (N_272,In_2194,In_120);
nor U273 (N_273,In_2288,In_524);
and U274 (N_274,In_1162,In_647);
xnor U275 (N_275,In_238,In_2165);
xnor U276 (N_276,In_667,In_1011);
or U277 (N_277,In_1877,In_769);
xnor U278 (N_278,In_855,In_1312);
and U279 (N_279,In_1609,In_1971);
or U280 (N_280,In_2132,In_1908);
nor U281 (N_281,In_256,In_107);
xnor U282 (N_282,In_664,In_1587);
nor U283 (N_283,In_1786,In_142);
or U284 (N_284,In_2240,In_1434);
or U285 (N_285,In_830,In_1541);
xnor U286 (N_286,In_0,In_1239);
nor U287 (N_287,In_1694,In_2206);
nor U288 (N_288,In_1281,In_1915);
nor U289 (N_289,In_379,In_2146);
nor U290 (N_290,In_2488,In_29);
xor U291 (N_291,In_2266,In_383);
and U292 (N_292,In_2373,In_1684);
xnor U293 (N_293,In_1654,In_2047);
xor U294 (N_294,In_1700,In_918);
nand U295 (N_295,In_1361,In_351);
nor U296 (N_296,In_1332,In_857);
and U297 (N_297,In_781,In_417);
nand U298 (N_298,In_267,In_1856);
nand U299 (N_299,In_2219,In_2374);
and U300 (N_300,In_1250,In_459);
xor U301 (N_301,In_2224,In_2061);
and U302 (N_302,In_372,In_766);
and U303 (N_303,In_1341,In_1426);
nand U304 (N_304,In_2060,In_85);
or U305 (N_305,In_2380,In_802);
nor U306 (N_306,In_1481,In_97);
and U307 (N_307,In_2113,In_9);
nor U308 (N_308,In_833,In_2199);
nor U309 (N_309,In_46,In_419);
or U310 (N_310,In_1472,In_1851);
nand U311 (N_311,In_1254,In_1793);
nor U312 (N_312,In_1676,In_2467);
xor U313 (N_313,In_1770,In_1867);
xor U314 (N_314,In_691,In_698);
or U315 (N_315,In_2428,In_1370);
or U316 (N_316,In_1440,In_450);
or U317 (N_317,In_416,In_1672);
or U318 (N_318,In_1508,In_2233);
nor U319 (N_319,In_815,In_984);
xnor U320 (N_320,In_2072,In_307);
nand U321 (N_321,In_1211,In_1024);
nand U322 (N_322,In_177,In_356);
xnor U323 (N_323,In_2468,In_1200);
and U324 (N_324,In_48,In_1551);
nor U325 (N_325,In_1739,In_76);
nand U326 (N_326,In_1833,In_413);
or U327 (N_327,In_258,In_1150);
and U328 (N_328,In_938,In_1974);
or U329 (N_329,In_2495,In_2420);
or U330 (N_330,In_397,In_1589);
and U331 (N_331,In_1050,In_2438);
or U332 (N_332,In_2411,In_264);
and U333 (N_333,In_2202,In_1108);
nor U334 (N_334,In_1133,In_2093);
nor U335 (N_335,In_562,In_595);
and U336 (N_336,In_251,In_1846);
and U337 (N_337,In_1588,In_823);
and U338 (N_338,In_1921,In_2387);
and U339 (N_339,In_1988,In_75);
xor U340 (N_340,In_1790,In_1823);
xnor U341 (N_341,In_1366,In_601);
nor U342 (N_342,In_975,In_1062);
nor U343 (N_343,In_371,In_173);
nand U344 (N_344,In_98,In_1759);
nor U345 (N_345,In_2077,In_2482);
xnor U346 (N_346,In_651,In_299);
nand U347 (N_347,In_1456,In_2114);
or U348 (N_348,In_2059,In_223);
nand U349 (N_349,In_1330,In_1375);
and U350 (N_350,In_1471,In_395);
xor U351 (N_351,In_1720,In_1825);
nor U352 (N_352,In_1960,In_1540);
nand U353 (N_353,In_906,In_288);
and U354 (N_354,In_628,In_1525);
nor U355 (N_355,In_208,In_2479);
xor U356 (N_356,In_710,In_1664);
nor U357 (N_357,In_549,In_1772);
nor U358 (N_358,In_1001,In_951);
xor U359 (N_359,In_1643,In_454);
or U360 (N_360,In_5,In_840);
and U361 (N_361,In_63,In_1325);
nand U362 (N_362,In_1443,In_1829);
xor U363 (N_363,In_1899,In_24);
or U364 (N_364,In_491,In_879);
or U365 (N_365,In_1479,In_1327);
xor U366 (N_366,In_891,In_605);
xor U367 (N_367,In_1708,In_1864);
nor U368 (N_368,In_2433,In_1068);
nand U369 (N_369,In_1487,In_441);
or U370 (N_370,In_703,In_835);
and U371 (N_371,In_2152,In_1917);
nand U372 (N_372,In_1081,In_767);
xnor U373 (N_373,In_1827,In_2347);
or U374 (N_374,In_1129,In_1716);
nand U375 (N_375,In_2176,In_2125);
and U376 (N_376,In_545,In_31);
or U377 (N_377,In_2209,In_1228);
and U378 (N_378,In_687,In_632);
xnor U379 (N_379,In_655,In_2129);
xnor U380 (N_380,In_928,In_184);
nor U381 (N_381,In_2097,In_186);
xor U382 (N_382,In_949,In_2471);
or U383 (N_383,In_82,In_1291);
nor U384 (N_384,In_1642,In_2419);
nor U385 (N_385,In_1979,In_1965);
xnor U386 (N_386,In_683,In_1522);
and U387 (N_387,In_1165,In_1621);
nand U388 (N_388,In_1698,In_597);
and U389 (N_389,In_700,In_1873);
nor U390 (N_390,In_1041,In_1536);
or U391 (N_391,In_1249,In_355);
nor U392 (N_392,In_1185,In_585);
or U393 (N_393,In_39,In_897);
or U394 (N_394,In_2351,In_2041);
or U395 (N_395,In_2135,In_768);
xnor U396 (N_396,In_1620,In_2331);
or U397 (N_397,In_2118,In_1882);
nor U398 (N_398,In_910,In_1895);
nand U399 (N_399,In_552,In_1379);
xor U400 (N_400,In_812,In_2300);
nor U401 (N_401,In_2290,In_145);
or U402 (N_402,In_1195,In_1571);
xor U403 (N_403,In_2280,In_1492);
or U404 (N_404,In_2264,In_90);
xor U405 (N_405,In_659,In_2407);
nor U406 (N_406,In_1635,In_1725);
nand U407 (N_407,In_255,In_1294);
and U408 (N_408,In_1447,In_814);
or U409 (N_409,In_571,In_2335);
nand U410 (N_410,In_1221,In_52);
nand U411 (N_411,In_2284,In_448);
nand U412 (N_412,In_1442,In_561);
nor U413 (N_413,In_1207,In_132);
nor U414 (N_414,In_1586,In_136);
xnor U415 (N_415,In_2396,In_1454);
nand U416 (N_416,In_2355,In_1820);
and U417 (N_417,In_1561,In_1105);
xnor U418 (N_418,In_2417,In_1391);
nor U419 (N_419,In_2252,In_842);
nor U420 (N_420,In_1139,In_1362);
nand U421 (N_421,In_2262,In_353);
and U422 (N_422,In_2051,In_2191);
nand U423 (N_423,In_318,In_1021);
nand U424 (N_424,In_1060,In_104);
nand U425 (N_425,In_665,In_2352);
and U426 (N_426,In_1549,In_1615);
xor U427 (N_427,In_778,In_1617);
or U428 (N_428,In_1124,In_2295);
xnor U429 (N_429,In_1058,In_1998);
nor U430 (N_430,In_290,In_2274);
nand U431 (N_431,In_1678,In_2378);
or U432 (N_432,In_1240,In_1942);
or U433 (N_433,In_2447,In_1224);
nor U434 (N_434,In_359,In_261);
xnor U435 (N_435,In_1984,In_992);
nor U436 (N_436,In_226,In_492);
nand U437 (N_437,In_851,In_1816);
or U438 (N_438,In_87,In_2153);
xor U439 (N_439,In_2103,In_1485);
and U440 (N_440,In_971,In_993);
xnor U441 (N_441,In_2394,In_1418);
xnor U442 (N_442,In_1337,In_608);
or U443 (N_443,In_695,In_2089);
nor U444 (N_444,In_1885,In_825);
or U445 (N_445,In_1719,In_957);
and U446 (N_446,In_1412,In_576);
or U447 (N_447,In_479,In_947);
or U448 (N_448,In_35,In_818);
xnor U449 (N_449,In_1410,In_1414);
nor U450 (N_450,In_599,In_1430);
nand U451 (N_451,In_1968,In_905);
xor U452 (N_452,In_2015,In_465);
xnor U453 (N_453,In_790,In_1388);
nand U454 (N_454,In_2108,In_1244);
nor U455 (N_455,In_175,In_547);
nand U456 (N_456,In_1841,In_1726);
xor U457 (N_457,In_2271,In_2185);
and U458 (N_458,In_1194,In_1558);
or U459 (N_459,In_727,In_513);
nor U460 (N_460,In_758,In_546);
nand U461 (N_461,In_1110,In_1329);
or U462 (N_462,In_853,In_1747);
xnor U463 (N_463,In_1083,In_2239);
and U464 (N_464,In_387,In_1099);
nand U465 (N_465,In_1048,In_1289);
or U466 (N_466,In_560,In_1721);
xor U467 (N_467,In_55,In_819);
nor U468 (N_468,In_1005,In_128);
nand U469 (N_469,In_1810,In_1723);
and U470 (N_470,In_846,In_1464);
and U471 (N_471,In_1744,In_2035);
nor U472 (N_472,In_1796,In_1087);
nand U473 (N_473,In_2499,In_570);
nand U474 (N_474,In_2345,In_1034);
or U475 (N_475,In_1850,In_431);
nor U476 (N_476,In_183,In_2008);
xor U477 (N_477,In_354,In_1437);
and U478 (N_478,In_1176,In_316);
and U479 (N_479,In_1318,In_2177);
nor U480 (N_480,In_673,In_1976);
nand U481 (N_481,In_1686,In_460);
nor U482 (N_482,In_529,In_2472);
xnor U483 (N_483,In_880,In_789);
or U484 (N_484,In_964,In_2065);
nor U485 (N_485,In_94,In_2293);
nand U486 (N_486,In_1259,In_1275);
nor U487 (N_487,In_2140,In_1098);
and U488 (N_488,In_875,In_2427);
and U489 (N_489,In_1740,In_1428);
nor U490 (N_490,In_1288,In_2267);
nand U491 (N_491,In_684,In_2084);
or U492 (N_492,In_2032,In_775);
xor U493 (N_493,In_604,In_1429);
nand U494 (N_494,In_1385,In_2339);
nand U495 (N_495,In_2473,In_311);
and U496 (N_496,In_308,In_2337);
or U497 (N_497,In_617,In_1893);
nor U498 (N_498,In_2159,In_788);
nor U499 (N_499,In_1037,In_1229);
and U500 (N_500,In_1948,In_1399);
or U501 (N_501,In_138,In_1798);
and U502 (N_502,In_2312,In_20);
nor U503 (N_503,In_1122,In_1128);
xnor U504 (N_504,In_1932,In_236);
nor U505 (N_505,In_831,In_1074);
xnor U506 (N_506,In_488,In_1773);
xor U507 (N_507,In_435,In_838);
nand U508 (N_508,In_2214,In_1529);
and U509 (N_509,In_1205,In_398);
or U510 (N_510,In_1542,In_2200);
and U511 (N_511,In_1547,In_544);
xnor U512 (N_512,In_2418,In_2350);
nand U513 (N_513,In_1502,In_907);
or U514 (N_514,In_658,In_2042);
or U515 (N_515,In_127,In_1118);
or U516 (N_516,In_725,In_2395);
nand U517 (N_517,In_380,In_2069);
xnor U518 (N_518,In_476,In_1350);
and U519 (N_519,In_36,In_1962);
nand U520 (N_520,In_970,In_110);
xnor U521 (N_521,In_1225,In_1146);
nand U522 (N_522,In_119,In_2075);
xor U523 (N_523,In_1946,In_323);
nor U524 (N_524,In_2329,In_1053);
nor U525 (N_525,In_1237,In_1599);
and U526 (N_526,In_663,In_477);
and U527 (N_527,In_1750,In_2088);
or U528 (N_528,In_2415,In_939);
nor U529 (N_529,In_27,In_694);
xnor U530 (N_530,In_1483,In_1067);
nand U531 (N_531,In_661,In_988);
or U532 (N_532,In_99,In_2079);
or U533 (N_533,In_95,In_2412);
nor U534 (N_534,In_639,In_1881);
and U535 (N_535,In_642,In_2400);
nor U536 (N_536,In_1567,In_2305);
xnor U537 (N_537,In_1579,In_415);
xor U538 (N_538,In_2340,In_403);
or U539 (N_539,In_870,In_1614);
and U540 (N_540,In_1756,In_1111);
or U541 (N_541,In_1484,In_348);
and U542 (N_542,In_2178,In_1416);
and U543 (N_543,In_485,In_991);
nor U544 (N_544,In_2360,In_1148);
or U545 (N_545,In_442,In_4);
nand U546 (N_546,In_286,In_1411);
xnor U547 (N_547,In_1016,In_1652);
nand U548 (N_548,In_28,In_922);
nor U549 (N_549,In_15,In_293);
nand U550 (N_550,In_1470,In_1255);
nor U551 (N_551,In_2334,In_2441);
nor U552 (N_552,In_2189,In_1657);
and U553 (N_553,In_1344,In_346);
xor U554 (N_554,In_948,In_2126);
nand U555 (N_555,In_1734,In_1548);
or U556 (N_556,In_770,In_265);
or U557 (N_557,In_1692,In_487);
and U558 (N_558,In_1780,In_2478);
nor U559 (N_559,In_754,In_1813);
xnor U560 (N_560,In_1550,In_1073);
nor U561 (N_561,In_2435,In_1817);
or U562 (N_562,In_1272,In_199);
and U563 (N_563,In_873,In_2030);
xor U564 (N_564,In_1156,In_2406);
xor U565 (N_565,In_2278,In_2248);
xor U566 (N_566,In_1781,In_1193);
nor U567 (N_567,In_1638,In_1303);
nand U568 (N_568,In_1722,In_1238);
nand U569 (N_569,In_1570,In_2301);
xor U570 (N_570,In_2164,In_2391);
xnor U571 (N_571,In_594,In_1565);
or U572 (N_572,In_1855,In_1164);
and U573 (N_573,In_1286,In_734);
nor U574 (N_574,In_1188,In_533);
nand U575 (N_575,In_30,In_1737);
and U576 (N_576,In_2414,In_1516);
and U577 (N_577,In_954,In_480);
nor U578 (N_578,In_950,In_1646);
xnor U579 (N_579,In_1563,In_920);
nor U580 (N_580,In_637,In_1461);
nor U581 (N_581,In_1929,In_369);
or U582 (N_582,In_402,In_38);
nand U583 (N_583,In_2410,In_1012);
xnor U584 (N_584,In_746,In_266);
and U585 (N_585,In_2242,In_776);
and U586 (N_586,In_166,In_1606);
nor U587 (N_587,In_41,In_565);
nand U588 (N_588,In_390,In_530);
nand U589 (N_589,In_1585,In_1363);
nand U590 (N_590,In_1757,In_1401);
nand U591 (N_591,In_2304,In_2094);
xor U592 (N_592,In_1766,In_1880);
nand U593 (N_593,In_1920,In_1999);
nand U594 (N_594,In_2027,In_1538);
or U595 (N_595,In_352,In_526);
nand U596 (N_596,In_490,In_1904);
xor U597 (N_597,In_2203,In_457);
nor U598 (N_598,In_2204,In_115);
and U599 (N_599,In_342,In_2263);
nand U600 (N_600,In_18,In_612);
xnor U601 (N_601,In_2073,In_1179);
nand U602 (N_602,In_625,In_1069);
and U603 (N_603,In_1027,In_339);
and U604 (N_604,In_941,In_321);
nor U605 (N_605,In_40,In_7);
nand U606 (N_606,In_811,In_148);
and U607 (N_607,In_1594,In_1253);
and U608 (N_608,In_535,In_937);
and U609 (N_609,In_2449,In_1623);
or U610 (N_610,In_108,In_1167);
or U611 (N_611,In_1504,In_602);
nand U612 (N_612,In_1295,In_1512);
xnor U613 (N_613,In_1354,In_1562);
nor U614 (N_614,In_386,In_1987);
xor U615 (N_615,In_418,In_756);
and U616 (N_616,In_1966,In_174);
and U617 (N_617,In_2310,In_1712);
or U618 (N_618,In_1473,In_1828);
nor U619 (N_619,In_1091,In_1061);
nand U620 (N_620,In_538,In_1805);
and U621 (N_621,In_606,In_374);
and U622 (N_622,In_985,In_813);
xnor U623 (N_623,In_1459,In_1697);
or U624 (N_624,In_2451,In_1710);
nor U625 (N_625,In_2247,In_1458);
and U626 (N_626,In_1112,In_1449);
or U627 (N_627,In_850,In_784);
and U628 (N_628,In_434,In_33);
and U629 (N_629,In_1086,In_1054);
and U630 (N_630,In_456,In_2182);
xor U631 (N_631,In_1397,In_1981);
nand U632 (N_632,In_1333,In_1996);
nand U633 (N_633,In_219,In_592);
nand U634 (N_634,In_1097,In_1025);
nor U635 (N_635,In_2070,In_786);
and U636 (N_636,In_1299,In_933);
nor U637 (N_637,In_901,In_2459);
or U638 (N_638,In_1208,In_2038);
or U639 (N_639,In_1120,In_1906);
or U640 (N_640,In_1004,In_1637);
and U641 (N_641,In_496,In_1431);
xor U642 (N_642,In_502,In_2205);
xor U643 (N_643,In_2308,In_164);
and U644 (N_644,In_1220,In_2349);
and U645 (N_645,In_1905,In_1741);
or U646 (N_646,In_2064,In_591);
nor U647 (N_647,In_2497,In_2357);
xor U648 (N_648,In_573,In_1491);
nand U649 (N_649,In_2215,In_1600);
or U650 (N_650,In_959,In_2133);
nand U651 (N_651,In_1990,In_1395);
xor U652 (N_652,In_81,In_461);
nand U653 (N_653,In_336,In_2033);
xor U654 (N_654,In_559,In_1056);
xnor U655 (N_655,In_2333,In_729);
xnor U656 (N_656,In_540,In_874);
nor U657 (N_657,In_2127,In_567);
nand U658 (N_658,In_609,In_1002);
nor U659 (N_659,In_1633,In_2379);
or U660 (N_660,In_187,In_472);
nor U661 (N_661,In_1049,In_447);
nand U662 (N_662,In_2422,In_654);
nand U663 (N_663,In_1,In_2485);
or U664 (N_664,In_2018,In_738);
or U665 (N_665,In_1270,In_122);
and U666 (N_666,In_762,In_1065);
or U667 (N_667,In_411,In_1141);
nand U668 (N_668,In_243,In_406);
xnor U669 (N_669,In_1376,In_588);
xnor U670 (N_670,In_635,In_500);
and U671 (N_671,In_1922,In_1951);
or U672 (N_672,In_1755,In_528);
or U673 (N_673,In_1230,In_349);
or U674 (N_674,In_583,In_2238);
xor U675 (N_675,In_681,In_2037);
or U676 (N_676,In_982,In_1226);
nor U677 (N_677,In_739,In_631);
nor U678 (N_678,In_404,In_2175);
nor U679 (N_679,In_972,In_1251);
and U680 (N_680,In_391,In_1641);
and U681 (N_681,In_440,In_652);
or U682 (N_682,In_1717,In_1977);
xor U683 (N_683,In_1916,In_202);
and U684 (N_684,In_1246,In_1234);
or U685 (N_685,In_1269,In_327);
nand U686 (N_686,In_1475,In_263);
xor U687 (N_687,In_1925,In_1931);
nor U688 (N_688,In_2249,In_2);
or U689 (N_689,In_1451,In_2229);
xor U690 (N_690,In_1753,In_1212);
nand U691 (N_691,In_543,In_1085);
xor U692 (N_692,In_1135,In_2095);
nand U693 (N_693,In_1982,In_67);
and U694 (N_694,In_2082,In_1243);
or U695 (N_695,In_451,In_1889);
or U696 (N_696,In_2120,In_1689);
xor U697 (N_697,In_1679,In_1940);
or U698 (N_698,In_1764,In_1389);
nor U699 (N_699,In_252,In_844);
xor U700 (N_700,In_2058,In_111);
nand U701 (N_701,In_1409,In_147);
nand U702 (N_702,In_624,In_1610);
xor U703 (N_703,In_2074,In_1876);
and U704 (N_704,In_1566,In_2317);
xor U705 (N_705,In_437,In_206);
nand U706 (N_706,In_1338,In_1619);
or U707 (N_707,In_1297,In_618);
and U708 (N_708,In_428,In_961);
or U709 (N_709,In_1180,In_309);
xnor U710 (N_710,In_1673,In_1774);
or U711 (N_711,In_1991,In_2048);
nand U712 (N_712,In_2019,In_1575);
nor U713 (N_713,In_1674,In_304);
or U714 (N_714,In_274,In_1404);
nand U715 (N_715,In_2116,In_1665);
xnor U716 (N_716,In_520,In_276);
xnor U717 (N_717,In_196,In_2265);
xnor U718 (N_718,In_931,In_394);
nor U719 (N_719,In_1506,In_1802);
and U720 (N_720,In_827,In_1076);
or U721 (N_721,In_2004,In_2062);
and U722 (N_722,In_1616,In_764);
nor U723 (N_723,In_914,In_1849);
or U724 (N_724,In_1668,In_1495);
or U725 (N_725,In_932,In_648);
xor U726 (N_726,In_341,In_179);
nor U727 (N_727,In_888,In_2158);
nor U728 (N_728,In_796,In_510);
xor U729 (N_729,In_1543,In_2134);
nand U730 (N_730,In_763,In_1305);
or U731 (N_731,In_859,In_367);
xor U732 (N_732,In_1611,In_1983);
nand U733 (N_733,In_344,In_1169);
and U734 (N_734,In_281,In_531);
or U735 (N_735,In_2163,In_455);
and U736 (N_736,In_2212,In_2292);
nand U737 (N_737,In_2401,In_57);
or U738 (N_738,In_103,In_960);
nor U739 (N_739,In_1386,In_1505);
nand U740 (N_740,In_1973,In_1022);
nand U741 (N_741,In_1352,In_1839);
xor U742 (N_742,In_965,In_1956);
xor U743 (N_743,In_1009,In_522);
nor U744 (N_744,In_2232,In_1155);
or U745 (N_745,In_1787,In_1210);
and U746 (N_746,In_2299,In_2269);
and U747 (N_747,In_1219,In_1439);
nor U748 (N_748,In_1498,In_366);
and U749 (N_749,In_780,In_969);
nand U750 (N_750,In_1537,In_2398);
and U751 (N_751,In_1101,In_1518);
nor U752 (N_752,In_1008,In_2014);
or U753 (N_753,In_782,In_1204);
nand U754 (N_754,In_2167,In_2466);
xor U755 (N_755,In_2423,In_2306);
nor U756 (N_756,In_1631,In_1373);
xnor U757 (N_757,In_2110,In_805);
nand U758 (N_758,In_1582,In_1331);
nor U759 (N_759,In_275,In_1886);
or U760 (N_760,In_2213,In_58);
and U761 (N_761,In_1394,In_885);
nor U762 (N_762,In_1824,In_2255);
nand U763 (N_763,In_1748,In_1699);
or U764 (N_764,In_1559,In_1913);
nand U765 (N_765,In_401,In_1866);
xor U766 (N_766,In_1455,In_2043);
nor U767 (N_767,In_1675,In_1190);
xor U768 (N_768,In_1527,In_1539);
or U769 (N_769,In_1634,In_425);
or U770 (N_770,In_1367,In_1095);
or U771 (N_771,In_225,In_630);
nand U772 (N_772,In_2409,In_1136);
nand U773 (N_773,In_772,In_444);
nor U774 (N_774,In_1775,In_439);
xor U775 (N_775,In_59,In_377);
nand U776 (N_776,In_2222,In_2002);
and U777 (N_777,In_2287,In_2368);
nor U778 (N_778,In_864,In_2025);
or U779 (N_779,In_2442,In_508);
or U780 (N_780,In_736,In_445);
and U781 (N_781,In_613,In_892);
and U782 (N_782,In_1453,In_636);
or U783 (N_783,In_178,In_718);
and U784 (N_784,In_1468,In_890);
and U785 (N_785,In_1533,In_167);
nor U786 (N_786,In_714,In_1296);
and U787 (N_787,In_375,In_2439);
and U788 (N_788,In_2251,In_1222);
or U789 (N_789,In_2201,In_999);
nor U790 (N_790,In_759,In_761);
nor U791 (N_791,In_660,In_486);
or U792 (N_792,In_1035,In_1724);
or U793 (N_793,In_1532,In_2464);
xor U794 (N_794,In_32,In_995);
nand U795 (N_795,In_432,In_558);
nand U796 (N_796,In_2057,In_1274);
xor U797 (N_797,In_696,In_572);
or U798 (N_798,In_2393,In_1842);
and U799 (N_799,In_1760,In_1020);
xnor U800 (N_800,In_2376,In_2273);
nor U801 (N_801,In_2170,In_1335);
nor U802 (N_802,In_1026,In_227);
nor U803 (N_803,In_1202,In_1353);
nand U804 (N_804,In_1355,In_896);
nand U805 (N_805,In_2322,In_1159);
nand U806 (N_806,In_2256,In_396);
and U807 (N_807,In_697,In_1268);
nand U808 (N_808,In_2371,In_929);
or U809 (N_809,In_189,In_936);
nand U810 (N_810,In_1280,In_2106);
xnor U811 (N_811,In_6,In_271);
nor U812 (N_812,In_1045,In_1242);
and U813 (N_813,In_2426,In_2281);
nor U814 (N_814,In_1214,In_19);
nor U815 (N_815,In_808,In_1347);
or U816 (N_816,In_1546,In_269);
xnor U817 (N_817,In_1859,In_51);
nor U818 (N_818,In_577,In_218);
nor U819 (N_819,In_724,In_2243);
or U820 (N_820,In_2154,In_2195);
nand U821 (N_821,In_934,In_1513);
nor U822 (N_822,In_877,In_181);
nand U823 (N_823,In_1057,In_924);
nor U824 (N_824,In_1903,In_728);
and U825 (N_825,In_2081,In_755);
xnor U826 (N_826,In_1082,In_1023);
nand U827 (N_827,In_237,In_201);
nor U828 (N_828,In_332,In_930);
nand U829 (N_829,In_1157,In_358);
or U830 (N_830,In_1650,In_504);
nand U831 (N_831,In_473,In_215);
nor U832 (N_832,In_1396,In_154);
or U833 (N_833,In_2217,In_1343);
or U834 (N_834,In_706,In_1432);
or U835 (N_835,In_84,In_1387);
or U836 (N_836,In_1573,In_284);
or U837 (N_837,In_1515,In_1283);
xnor U838 (N_838,In_2404,In_155);
nand U839 (N_839,In_365,In_1324);
or U840 (N_840,In_2001,In_2141);
and U841 (N_841,In_2100,In_744);
xor U842 (N_842,In_248,In_1807);
xnor U843 (N_843,In_935,In_1093);
and U844 (N_844,In_1711,In_2244);
or U845 (N_845,In_2385,In_1656);
nor U846 (N_846,In_1944,In_112);
and U847 (N_847,In_373,In_645);
nor U848 (N_848,In_1160,In_1046);
and U849 (N_849,In_78,In_1121);
xnor U850 (N_850,In_1047,In_963);
or U851 (N_851,In_1878,In_1681);
and U852 (N_852,In_1779,In_693);
nor U853 (N_853,In_1510,In_1514);
or U854 (N_854,In_615,In_1683);
and U855 (N_855,In_1738,In_216);
and U856 (N_856,In_1154,In_1102);
xnor U857 (N_857,In_1125,In_717);
or U858 (N_858,In_1818,In_534);
nor U859 (N_859,In_1728,In_607);
xnor U860 (N_860,In_489,In_1861);
nor U861 (N_861,In_2375,In_422);
nand U862 (N_862,In_1315,In_1936);
and U863 (N_863,In_1706,In_113);
nand U864 (N_864,In_523,In_797);
and U865 (N_865,In_1422,In_1182);
or U866 (N_866,In_26,In_829);
nor U867 (N_867,In_1359,In_278);
nand U868 (N_868,In_160,In_816);
nand U869 (N_869,In_2283,In_1064);
nand U870 (N_870,In_2272,In_2384);
nand U871 (N_871,In_151,In_158);
and U872 (N_872,In_1863,In_2450);
xnor U873 (N_873,In_306,In_723);
nor U874 (N_874,In_1745,In_1213);
xor U875 (N_875,In_943,In_1466);
nor U876 (N_876,In_1519,In_521);
nand U877 (N_877,In_2448,In_2220);
xor U878 (N_878,In_1530,In_2416);
and U879 (N_879,In_2307,In_2101);
or U880 (N_880,In_2430,In_1000);
nor U881 (N_881,In_2149,In_1632);
nand U882 (N_882,In_1564,In_1052);
and U883 (N_883,In_1601,In_1203);
or U884 (N_884,In_140,In_1393);
and U885 (N_885,In_672,In_1088);
nor U886 (N_886,In_123,In_1875);
and U887 (N_887,In_2009,In_621);
and U888 (N_888,In_2003,In_2270);
or U889 (N_889,In_1995,In_1042);
nand U890 (N_890,In_1924,In_2279);
or U891 (N_891,In_662,In_121);
and U892 (N_892,In_1425,In_760);
or U893 (N_893,In_944,In_2323);
and U894 (N_894,In_2115,In_2303);
or U895 (N_895,In_980,In_2480);
or U896 (N_896,In_2234,In_2296);
or U897 (N_897,In_205,In_582);
nor U898 (N_898,In_2193,In_2382);
and U899 (N_899,In_1630,In_1792);
xnor U900 (N_900,In_399,In_721);
and U901 (N_901,In_820,In_245);
nand U902 (N_902,In_2087,In_105);
or U903 (N_903,In_537,In_2228);
xnor U904 (N_904,In_745,In_310);
and U905 (N_905,In_1446,In_363);
xor U906 (N_906,In_501,In_1096);
xor U907 (N_907,In_2139,In_551);
nor U908 (N_908,In_794,In_1170);
or U909 (N_909,In_1308,In_2184);
xor U910 (N_910,In_295,In_2302);
nor U911 (N_911,In_1560,In_713);
or U912 (N_912,In_783,In_2324);
xor U913 (N_913,In_2207,In_2236);
or U914 (N_914,In_1767,In_1844);
nand U915 (N_915,In_2465,In_854);
and U916 (N_916,In_1084,In_1531);
and U917 (N_917,In_1258,In_2470);
and U918 (N_918,In_2402,In_2463);
nand U919 (N_919,In_2111,In_876);
nor U920 (N_920,In_809,In_2123);
or U921 (N_921,In_1115,In_2130);
xor U922 (N_922,In_881,In_1993);
nand U923 (N_923,In_2053,In_1819);
nand U924 (N_924,In_1063,In_1803);
and U925 (N_925,In_1874,In_1192);
nand U926 (N_926,In_1184,In_2453);
nor U927 (N_927,In_555,In_2096);
nand U928 (N_928,In_1450,In_1413);
xnor U929 (N_929,In_1371,In_974);
or U930 (N_930,In_765,In_2364);
nand U931 (N_931,In_420,In_2260);
and U932 (N_932,In_1858,In_1612);
nand U933 (N_933,In_2392,In_841);
and U934 (N_934,In_89,In_1535);
xor U935 (N_935,In_1980,In_1939);
nor U936 (N_936,In_678,In_581);
and U937 (N_937,In_1173,In_1769);
xor U938 (N_938,In_737,In_296);
xnor U939 (N_939,In_564,In_312);
or U940 (N_940,In_56,In_824);
nand U941 (N_941,In_157,In_1534);
or U942 (N_942,In_1356,In_106);
or U943 (N_943,In_2137,In_1970);
or U944 (N_944,In_848,In_156);
nor U945 (N_945,In_220,In_62);
nor U946 (N_946,In_590,In_847);
xor U947 (N_947,In_2277,In_578);
xnor U948 (N_948,In_228,In_1900);
and U949 (N_949,In_2446,In_1314);
or U950 (N_950,In_2020,In_862);
nand U951 (N_951,In_463,In_2031);
and U952 (N_952,In_37,In_1624);
xnor U953 (N_953,In_65,In_2397);
nand U954 (N_954,In_1972,In_2336);
nor U955 (N_955,In_2462,In_803);
nand U956 (N_956,In_23,In_259);
nand U957 (N_957,In_1919,In_54);
nand U958 (N_958,In_2221,In_303);
or U959 (N_959,In_79,In_194);
nand U960 (N_960,In_707,In_2026);
nand U961 (N_961,In_977,In_800);
nand U962 (N_962,In_2055,In_2044);
and U963 (N_963,In_114,In_866);
xnor U964 (N_964,In_2190,In_298);
xor U965 (N_965,In_968,In_2338);
and U966 (N_966,In_1947,In_923);
or U967 (N_967,In_507,In_1257);
nand U968 (N_968,In_1852,In_675);
or U969 (N_969,In_953,In_705);
nor U970 (N_970,In_2045,In_1975);
and U971 (N_971,In_1831,In_1836);
or U972 (N_972,In_743,In_388);
nand U973 (N_973,In_836,In_433);
nand U974 (N_974,In_740,In_1580);
nor U975 (N_975,In_2198,In_527);
and U976 (N_976,In_1266,In_1898);
nor U977 (N_977,In_871,In_679);
nand U978 (N_978,In_452,In_1307);
xor U979 (N_979,In_550,In_1768);
xnor U980 (N_980,In_2112,In_1784);
nor U981 (N_981,In_856,In_1252);
and U982 (N_982,In_852,In_2226);
xor U983 (N_983,In_978,In_313);
nor U984 (N_984,In_34,In_1278);
xor U985 (N_985,In_1511,In_1785);
nand U986 (N_986,In_1572,In_1117);
nand U987 (N_987,In_2078,In_453);
nor U988 (N_988,In_2496,In_282);
xnor U989 (N_989,In_817,In_124);
or U990 (N_990,In_429,In_86);
xor U991 (N_991,In_2437,In_858);
or U992 (N_992,In_272,In_1206);
and U993 (N_993,In_2188,In_1015);
and U994 (N_994,In_2365,In_1406);
nor U995 (N_995,In_1104,In_1438);
nor U996 (N_996,In_752,In_690);
nand U997 (N_997,In_300,In_118);
nand U998 (N_998,In_1051,In_2166);
xnor U999 (N_999,In_895,In_1834);
nand U1000 (N_1000,In_1865,In_1687);
xor U1001 (N_1001,In_1490,In_806);
and U1002 (N_1002,In_498,In_987);
nand U1003 (N_1003,In_2012,In_1465);
and U1004 (N_1004,In_1659,In_2013);
or U1005 (N_1005,In_1436,In_735);
or U1006 (N_1006,In_368,In_799);
xor U1007 (N_1007,In_2128,In_333);
and U1008 (N_1008,In_1311,In_1625);
nand U1009 (N_1009,In_1320,In_2326);
and U1010 (N_1010,In_2327,In_1181);
nor U1011 (N_1011,In_2145,In_1149);
and U1012 (N_1012,In_163,In_1608);
nor U1013 (N_1013,In_1313,In_74);
or U1014 (N_1014,In_541,In_381);
nand U1015 (N_1015,In_1390,In_389);
xnor U1016 (N_1016,In_2151,In_2218);
nand U1017 (N_1017,In_1215,In_1187);
nor U1018 (N_1018,In_324,In_1890);
and U1019 (N_1019,In_2369,In_2405);
nor U1020 (N_1020,In_1223,In_1645);
xor U1021 (N_1021,In_2050,In_1961);
nand U1022 (N_1022,In_777,In_2291);
and U1023 (N_1023,In_1302,In_2052);
xor U1024 (N_1024,In_1151,In_927);
or U1025 (N_1025,In_1777,In_1340);
nand U1026 (N_1026,In_1006,In_68);
nand U1027 (N_1027,In_1927,In_1232);
and U1028 (N_1028,In_2268,In_16);
and U1029 (N_1029,In_141,In_1209);
or U1030 (N_1030,In_287,In_1902);
and U1031 (N_1031,In_2168,In_378);
nor U1032 (N_1032,In_1300,In_634);
and U1033 (N_1033,In_1918,In_709);
or U1034 (N_1034,In_1134,In_1897);
nand U1035 (N_1035,In_1941,In_1419);
or U1036 (N_1036,In_1198,In_2063);
and U1037 (N_1037,In_268,In_2083);
and U1038 (N_1038,In_656,In_481);
nor U1039 (N_1039,In_1427,In_2285);
or U1040 (N_1040,In_2390,In_139);
nor U1041 (N_1041,In_1349,In_427);
and U1042 (N_1042,In_1653,In_88);
nor U1043 (N_1043,In_904,In_1680);
xor U1044 (N_1044,In_845,In_2314);
and U1045 (N_1045,In_2469,In_2348);
and U1046 (N_1046,In_1736,In_1245);
and U1047 (N_1047,In_1336,In_239);
and U1048 (N_1048,In_1801,In_1928);
nand U1049 (N_1049,In_438,In_956);
xnor U1050 (N_1050,In_133,In_1298);
nor U1051 (N_1051,In_1334,In_43);
xor U1052 (N_1052,In_2192,In_207);
nand U1053 (N_1053,In_1840,In_337);
or U1054 (N_1054,In_1301,In_600);
or U1055 (N_1055,In_231,In_436);
xor U1056 (N_1056,In_1236,In_257);
nor U1057 (N_1057,In_843,In_1094);
xnor U1058 (N_1058,In_1378,In_1595);
nand U1059 (N_1059,In_2173,In_1914);
nor U1060 (N_1060,In_191,In_159);
nand U1061 (N_1061,In_1441,In_471);
nand U1062 (N_1062,In_2011,In_1556);
nor U1063 (N_1063,In_1554,In_1735);
or U1064 (N_1064,In_210,In_1754);
nor U1065 (N_1065,In_1503,In_1590);
and U1066 (N_1066,In_1044,In_1935);
or U1067 (N_1067,In_2117,In_1477);
or U1068 (N_1068,In_329,In_405);
nand U1069 (N_1069,In_1795,In_469);
xor U1070 (N_1070,In_69,In_2227);
nand U1071 (N_1071,In_701,In_483);
or U1072 (N_1072,In_325,In_593);
nand U1073 (N_1073,In_1201,In_1369);
nand U1074 (N_1074,In_1132,In_1196);
and U1075 (N_1075,In_657,In_1907);
or U1076 (N_1076,In_1177,In_2005);
nand U1077 (N_1077,In_1127,In_1964);
nand U1078 (N_1078,In_1727,In_1526);
nand U1079 (N_1079,In_176,In_467);
and U1080 (N_1080,In_2028,In_2486);
and U1081 (N_1081,In_250,In_849);
nor U1082 (N_1082,In_976,In_1763);
xnor U1083 (N_1083,In_224,In_1783);
xor U1084 (N_1084,In_1501,In_1448);
nand U1085 (N_1085,In_2289,In_1271);
nand U1086 (N_1086,In_2142,In_512);
nand U1087 (N_1087,In_1463,In_1926);
or U1088 (N_1088,In_2138,In_1028);
and U1089 (N_1089,In_2196,In_1499);
or U1090 (N_1090,In_1626,In_1677);
or U1091 (N_1091,In_297,In_170);
or U1092 (N_1092,In_2388,In_328);
xor U1093 (N_1093,In_1574,In_867);
xor U1094 (N_1094,In_1891,In_915);
xor U1095 (N_1095,In_1392,In_2021);
nor U1096 (N_1096,In_2016,In_2328);
and U1097 (N_1097,In_1938,In_556);
nor U1098 (N_1098,In_2356,In_2498);
xor U1099 (N_1099,In_1417,In_1013);
and U1100 (N_1100,In_302,In_2046);
or U1101 (N_1101,In_1838,In_861);
or U1102 (N_1102,In_994,In_680);
nand U1103 (N_1103,In_1158,In_1544);
or U1104 (N_1104,In_180,In_668);
and U1105 (N_1105,In_1648,In_116);
nand U1106 (N_1106,In_2319,In_1103);
nor U1107 (N_1107,In_153,In_989);
and U1108 (N_1108,In_539,In_1372);
or U1109 (N_1109,In_925,In_2246);
nor U1110 (N_1110,In_25,In_285);
or U1111 (N_1111,In_1080,In_1075);
xor U1112 (N_1112,In_801,In_2068);
and U1113 (N_1113,In_1598,In_1704);
xnor U1114 (N_1114,In_1066,In_185);
and U1115 (N_1115,In_11,In_262);
and U1116 (N_1116,In_826,In_1869);
and U1117 (N_1117,In_340,In_2493);
nand U1118 (N_1118,In_53,In_1460);
or U1119 (N_1119,In_192,In_603);
nand U1120 (N_1120,In_1809,In_1077);
xnor U1121 (N_1121,In_102,In_10);
xor U1122 (N_1122,In_998,In_400);
nor U1123 (N_1123,In_650,In_566);
and U1124 (N_1124,In_1507,In_1408);
or U1125 (N_1125,In_525,In_1285);
and U1126 (N_1126,In_1557,In_1142);
and U1127 (N_1127,In_828,In_1374);
and U1128 (N_1128,In_2311,In_983);
or U1129 (N_1129,In_1360,In_1306);
and U1130 (N_1130,In_347,In_44);
or U1131 (N_1131,In_47,In_623);
xor U1132 (N_1132,In_1553,In_474);
and U1133 (N_1133,In_2144,In_2431);
or U1134 (N_1134,In_644,In_945);
nand U1135 (N_1135,In_1189,In_886);
nor U1136 (N_1136,In_536,In_1161);
or U1137 (N_1137,In_2460,In_716);
or U1138 (N_1138,In_1830,In_2034);
nor U1139 (N_1139,In_384,In_1216);
xnor U1140 (N_1140,In_1218,In_2085);
and U1141 (N_1141,In_203,In_1520);
nor U1142 (N_1142,In_1486,In_2230);
or U1143 (N_1143,In_913,In_1958);
nand U1144 (N_1144,In_940,In_12);
nor U1145 (N_1145,In_162,In_2208);
and U1146 (N_1146,In_2086,In_1771);
nand U1147 (N_1147,In_1351,In_2225);
nor U1148 (N_1148,In_71,In_2237);
and U1149 (N_1149,In_409,In_1382);
and U1150 (N_1150,In_967,In_343);
nor U1151 (N_1151,In_1800,In_17);
xnor U1152 (N_1152,In_1667,In_868);
and U1153 (N_1153,In_1901,In_283);
xor U1154 (N_1154,In_990,In_2458);
nand U1155 (N_1155,In_246,In_1854);
xnor U1156 (N_1156,In_1163,In_129);
or U1157 (N_1157,In_646,In_1746);
nand U1158 (N_1158,In_1493,In_2346);
and U1159 (N_1159,In_2362,In_1808);
nand U1160 (N_1160,In_2294,In_515);
and U1161 (N_1161,In_244,In_364);
nor U1162 (N_1162,In_1978,In_212);
or U1163 (N_1163,In_345,In_1832);
nor U1164 (N_1164,In_1172,In_640);
nor U1165 (N_1165,In_619,In_462);
xnor U1166 (N_1166,In_362,In_1670);
nand U1167 (N_1167,In_2344,In_1887);
and U1168 (N_1168,In_516,In_1584);
or U1169 (N_1169,In_1663,In_209);
or U1170 (N_1170,In_719,In_997);
and U1171 (N_1171,In_1178,In_1233);
and U1172 (N_1172,In_13,In_1368);
xnor U1173 (N_1173,In_1038,In_757);
nor U1174 (N_1174,In_666,In_2023);
and U1175 (N_1175,In_2080,In_1107);
nand U1176 (N_1176,In_1290,In_2354);
xnor U1177 (N_1177,In_2424,In_1480);
or U1178 (N_1178,In_326,In_1358);
or U1179 (N_1179,In_2421,In_730);
xor U1180 (N_1180,In_2452,In_408);
and U1181 (N_1181,In_1282,In_596);
or U1182 (N_1182,In_2443,In_509);
and U1183 (N_1183,In_317,In_962);
nand U1184 (N_1184,In_1576,In_475);
nor U1185 (N_1185,In_1445,In_1896);
or U1186 (N_1186,In_2342,In_1985);
nand U1187 (N_1187,In_1666,In_1627);
xnor U1188 (N_1188,In_2092,In_1197);
nand U1189 (N_1189,In_1231,In_671);
xnor U1190 (N_1190,In_2313,In_1605);
or U1191 (N_1191,In_1806,In_2282);
and U1192 (N_1192,In_1348,In_292);
nor U1193 (N_1193,In_1264,In_773);
nand U1194 (N_1194,In_1703,In_169);
and U1195 (N_1195,In_2363,In_322);
nand U1196 (N_1196,In_2494,In_2259);
and U1197 (N_1197,In_1662,In_1090);
and U1198 (N_1198,In_1316,In_519);
or U1199 (N_1199,In_1383,In_726);
and U1200 (N_1200,In_1279,In_1986);
xor U1201 (N_1201,In_1658,In_1029);
nor U1202 (N_1202,In_392,In_926);
xnor U1203 (N_1203,In_8,In_900);
nor U1204 (N_1204,In_2090,In_1837);
or U1205 (N_1205,In_1732,In_2211);
xor U1206 (N_1206,In_1622,In_587);
nor U1207 (N_1207,In_2022,In_2481);
and U1208 (N_1208,In_2150,In_1949);
nor U1209 (N_1209,In_494,In_2332);
or U1210 (N_1210,In_589,In_301);
nor U1211 (N_1211,In_1377,In_804);
xor U1212 (N_1212,In_1751,In_1263);
or U1213 (N_1213,In_2241,In_14);
nand U1214 (N_1214,In_2160,In_722);
nand U1215 (N_1215,In_753,In_505);
and U1216 (N_1216,In_2330,In_1870);
xor U1217 (N_1217,In_785,In_955);
and U1218 (N_1218,In_1963,In_289);
and U1219 (N_1219,In_732,In_149);
xor U1220 (N_1220,In_1761,In_1346);
or U1221 (N_1221,In_1017,In_1660);
or U1222 (N_1222,In_2389,In_1467);
nand U1223 (N_1223,In_2049,In_1636);
and U1224 (N_1224,In_1957,In_579);
nor U1225 (N_1225,In_903,In_1323);
nor U1226 (N_1226,In_2286,In_1496);
or U1227 (N_1227,In_1702,In_2161);
and U1228 (N_1228,In_2180,In_674);
nor U1229 (N_1229,In_2197,In_2477);
nand U1230 (N_1230,In_1569,In_622);
or U1231 (N_1231,In_1967,In_499);
or U1232 (N_1232,In_168,In_2109);
and U1233 (N_1233,In_629,In_1402);
nor U1234 (N_1234,In_741,In_568);
nor U1235 (N_1235,In_2316,In_916);
and U1236 (N_1236,In_1892,In_2325);
nand U1237 (N_1237,In_211,In_1310);
or U1238 (N_1238,In_1199,In_2143);
nand U1239 (N_1239,In_2254,In_1682);
and U1240 (N_1240,In_2257,In_676);
nor U1241 (N_1241,In_1655,In_2216);
and U1242 (N_1242,In_1059,In_2361);
nand U1243 (N_1243,In_171,In_1555);
and U1244 (N_1244,In_2386,In_117);
xnor U1245 (N_1245,In_1055,In_1174);
xnor U1246 (N_1246,In_478,In_575);
nor U1247 (N_1247,In_1403,In_2107);
xor U1248 (N_1248,In_1552,In_2102);
or U1249 (N_1249,In_1405,In_315);
and U1250 (N_1250,In_491,In_150);
nor U1251 (N_1251,In_1298,In_2122);
xnor U1252 (N_1252,In_1632,In_1728);
nand U1253 (N_1253,In_1494,In_1469);
and U1254 (N_1254,In_525,In_137);
and U1255 (N_1255,In_1014,In_150);
xnor U1256 (N_1256,In_554,In_1022);
nand U1257 (N_1257,In_908,In_274);
xor U1258 (N_1258,In_100,In_679);
or U1259 (N_1259,In_1538,In_1161);
nand U1260 (N_1260,In_165,In_1793);
or U1261 (N_1261,In_753,In_599);
nand U1262 (N_1262,In_2392,In_1627);
xnor U1263 (N_1263,In_2146,In_1339);
nor U1264 (N_1264,In_1743,In_1759);
xnor U1265 (N_1265,In_1196,In_468);
xor U1266 (N_1266,In_1146,In_1256);
and U1267 (N_1267,In_683,In_2497);
nor U1268 (N_1268,In_1125,In_1755);
or U1269 (N_1269,In_912,In_451);
nor U1270 (N_1270,In_2120,In_1792);
nand U1271 (N_1271,In_941,In_1465);
nor U1272 (N_1272,In_1090,In_1844);
nor U1273 (N_1273,In_1573,In_945);
nor U1274 (N_1274,In_184,In_1321);
xnor U1275 (N_1275,In_1752,In_1772);
and U1276 (N_1276,In_436,In_925);
and U1277 (N_1277,In_499,In_1425);
or U1278 (N_1278,In_638,In_299);
nor U1279 (N_1279,In_2125,In_99);
or U1280 (N_1280,In_637,In_2208);
or U1281 (N_1281,In_217,In_694);
and U1282 (N_1282,In_250,In_1148);
nand U1283 (N_1283,In_13,In_1707);
and U1284 (N_1284,In_354,In_937);
nor U1285 (N_1285,In_63,In_1153);
xor U1286 (N_1286,In_1761,In_568);
nor U1287 (N_1287,In_1038,In_1636);
nor U1288 (N_1288,In_1727,In_1268);
nand U1289 (N_1289,In_858,In_956);
nand U1290 (N_1290,In_1749,In_543);
xnor U1291 (N_1291,In_354,In_2238);
or U1292 (N_1292,In_2256,In_448);
xnor U1293 (N_1293,In_1211,In_2005);
nand U1294 (N_1294,In_2107,In_1975);
or U1295 (N_1295,In_2387,In_1411);
or U1296 (N_1296,In_1257,In_2336);
nand U1297 (N_1297,In_892,In_516);
nor U1298 (N_1298,In_1460,In_1662);
nand U1299 (N_1299,In_319,In_877);
or U1300 (N_1300,In_1600,In_2226);
nand U1301 (N_1301,In_897,In_384);
xor U1302 (N_1302,In_496,In_1720);
or U1303 (N_1303,In_187,In_1149);
nor U1304 (N_1304,In_1634,In_173);
and U1305 (N_1305,In_2374,In_201);
nand U1306 (N_1306,In_1592,In_1446);
nand U1307 (N_1307,In_2328,In_354);
xor U1308 (N_1308,In_855,In_1197);
nor U1309 (N_1309,In_1916,In_1627);
and U1310 (N_1310,In_1964,In_381);
and U1311 (N_1311,In_58,In_409);
nor U1312 (N_1312,In_2029,In_110);
nor U1313 (N_1313,In_1712,In_2359);
nor U1314 (N_1314,In_1058,In_132);
nand U1315 (N_1315,In_1356,In_345);
or U1316 (N_1316,In_1253,In_212);
or U1317 (N_1317,In_261,In_986);
nor U1318 (N_1318,In_2319,In_1949);
xor U1319 (N_1319,In_2060,In_2241);
xnor U1320 (N_1320,In_1364,In_938);
nand U1321 (N_1321,In_1580,In_1876);
nand U1322 (N_1322,In_727,In_448);
nor U1323 (N_1323,In_367,In_2214);
nor U1324 (N_1324,In_2388,In_2212);
xnor U1325 (N_1325,In_1922,In_1646);
nand U1326 (N_1326,In_1180,In_2324);
nand U1327 (N_1327,In_1942,In_2037);
nand U1328 (N_1328,In_2057,In_776);
nor U1329 (N_1329,In_1214,In_1876);
and U1330 (N_1330,In_1698,In_934);
nor U1331 (N_1331,In_1201,In_74);
nand U1332 (N_1332,In_1070,In_834);
and U1333 (N_1333,In_237,In_1932);
nand U1334 (N_1334,In_273,In_1906);
xor U1335 (N_1335,In_1823,In_1031);
xnor U1336 (N_1336,In_1109,In_2418);
and U1337 (N_1337,In_1629,In_503);
xnor U1338 (N_1338,In_391,In_2219);
and U1339 (N_1339,In_53,In_1560);
nand U1340 (N_1340,In_1696,In_1786);
xor U1341 (N_1341,In_1256,In_843);
and U1342 (N_1342,In_1672,In_962);
nand U1343 (N_1343,In_501,In_316);
nor U1344 (N_1344,In_781,In_1768);
nand U1345 (N_1345,In_1827,In_1759);
nand U1346 (N_1346,In_794,In_801);
xor U1347 (N_1347,In_778,In_1814);
nor U1348 (N_1348,In_1571,In_2009);
or U1349 (N_1349,In_303,In_1644);
nor U1350 (N_1350,In_1803,In_1797);
xnor U1351 (N_1351,In_2363,In_1402);
xor U1352 (N_1352,In_2303,In_2018);
xor U1353 (N_1353,In_1098,In_1382);
nand U1354 (N_1354,In_113,In_2268);
xor U1355 (N_1355,In_118,In_1779);
nor U1356 (N_1356,In_2068,In_766);
xor U1357 (N_1357,In_2300,In_1774);
xnor U1358 (N_1358,In_2101,In_682);
xor U1359 (N_1359,In_1976,In_2230);
and U1360 (N_1360,In_942,In_1893);
nor U1361 (N_1361,In_1638,In_11);
or U1362 (N_1362,In_87,In_977);
nor U1363 (N_1363,In_291,In_1216);
nor U1364 (N_1364,In_1878,In_382);
and U1365 (N_1365,In_2189,In_2187);
nand U1366 (N_1366,In_265,In_64);
nor U1367 (N_1367,In_1178,In_299);
nor U1368 (N_1368,In_980,In_2322);
or U1369 (N_1369,In_496,In_1430);
or U1370 (N_1370,In_725,In_749);
xor U1371 (N_1371,In_47,In_1447);
nor U1372 (N_1372,In_1847,In_76);
xnor U1373 (N_1373,In_1383,In_133);
nand U1374 (N_1374,In_1038,In_1779);
and U1375 (N_1375,In_806,In_557);
nand U1376 (N_1376,In_1953,In_631);
or U1377 (N_1377,In_2037,In_1114);
or U1378 (N_1378,In_196,In_1079);
or U1379 (N_1379,In_1792,In_723);
and U1380 (N_1380,In_649,In_2438);
and U1381 (N_1381,In_647,In_814);
xor U1382 (N_1382,In_2136,In_910);
nand U1383 (N_1383,In_665,In_826);
nand U1384 (N_1384,In_1277,In_898);
nor U1385 (N_1385,In_37,In_1424);
nand U1386 (N_1386,In_1583,In_1116);
or U1387 (N_1387,In_1285,In_285);
or U1388 (N_1388,In_1437,In_2441);
and U1389 (N_1389,In_2286,In_144);
and U1390 (N_1390,In_1052,In_387);
xnor U1391 (N_1391,In_342,In_547);
or U1392 (N_1392,In_673,In_133);
xor U1393 (N_1393,In_1614,In_1895);
nand U1394 (N_1394,In_745,In_1289);
and U1395 (N_1395,In_1843,In_301);
xnor U1396 (N_1396,In_2115,In_599);
xnor U1397 (N_1397,In_1394,In_1268);
or U1398 (N_1398,In_179,In_107);
and U1399 (N_1399,In_498,In_619);
nor U1400 (N_1400,In_1502,In_1467);
xor U1401 (N_1401,In_281,In_2045);
and U1402 (N_1402,In_2452,In_961);
xnor U1403 (N_1403,In_2473,In_855);
and U1404 (N_1404,In_2397,In_2272);
xor U1405 (N_1405,In_1323,In_1826);
xor U1406 (N_1406,In_2292,In_655);
and U1407 (N_1407,In_316,In_1422);
xnor U1408 (N_1408,In_1824,In_1787);
nor U1409 (N_1409,In_1619,In_662);
or U1410 (N_1410,In_1510,In_1588);
xor U1411 (N_1411,In_1067,In_428);
and U1412 (N_1412,In_2359,In_184);
nor U1413 (N_1413,In_724,In_2394);
nand U1414 (N_1414,In_1607,In_2068);
xnor U1415 (N_1415,In_279,In_681);
and U1416 (N_1416,In_2348,In_1803);
nor U1417 (N_1417,In_1581,In_1447);
nand U1418 (N_1418,In_383,In_1301);
xor U1419 (N_1419,In_1523,In_865);
nor U1420 (N_1420,In_1672,In_309);
xnor U1421 (N_1421,In_885,In_1325);
or U1422 (N_1422,In_1008,In_786);
nand U1423 (N_1423,In_2138,In_1992);
and U1424 (N_1424,In_1782,In_2095);
nor U1425 (N_1425,In_2189,In_1642);
or U1426 (N_1426,In_1254,In_1604);
xnor U1427 (N_1427,In_486,In_631);
nor U1428 (N_1428,In_1524,In_1876);
nand U1429 (N_1429,In_1114,In_342);
and U1430 (N_1430,In_1396,In_541);
xor U1431 (N_1431,In_1340,In_1471);
nand U1432 (N_1432,In_1292,In_2152);
xor U1433 (N_1433,In_318,In_1136);
nand U1434 (N_1434,In_1019,In_539);
nand U1435 (N_1435,In_1476,In_410);
xnor U1436 (N_1436,In_2356,In_1369);
or U1437 (N_1437,In_958,In_1116);
and U1438 (N_1438,In_483,In_1199);
nand U1439 (N_1439,In_1425,In_1398);
nand U1440 (N_1440,In_2113,In_714);
nor U1441 (N_1441,In_1257,In_425);
and U1442 (N_1442,In_2137,In_1531);
xnor U1443 (N_1443,In_55,In_1078);
or U1444 (N_1444,In_740,In_848);
and U1445 (N_1445,In_2367,In_1030);
or U1446 (N_1446,In_83,In_1662);
xnor U1447 (N_1447,In_613,In_376);
nor U1448 (N_1448,In_179,In_2207);
nor U1449 (N_1449,In_1053,In_2166);
nor U1450 (N_1450,In_1391,In_113);
and U1451 (N_1451,In_2135,In_1725);
or U1452 (N_1452,In_977,In_837);
or U1453 (N_1453,In_2057,In_773);
or U1454 (N_1454,In_2304,In_996);
nand U1455 (N_1455,In_2191,In_1485);
nor U1456 (N_1456,In_2309,In_1981);
nand U1457 (N_1457,In_2061,In_1774);
or U1458 (N_1458,In_1705,In_1207);
xnor U1459 (N_1459,In_983,In_950);
nand U1460 (N_1460,In_1294,In_1850);
or U1461 (N_1461,In_1138,In_2291);
or U1462 (N_1462,In_2192,In_507);
or U1463 (N_1463,In_2491,In_926);
nand U1464 (N_1464,In_2094,In_1796);
xnor U1465 (N_1465,In_895,In_1518);
and U1466 (N_1466,In_2052,In_886);
and U1467 (N_1467,In_1665,In_2362);
nand U1468 (N_1468,In_1037,In_1067);
or U1469 (N_1469,In_1263,In_2352);
xnor U1470 (N_1470,In_498,In_676);
or U1471 (N_1471,In_922,In_146);
and U1472 (N_1472,In_2059,In_266);
xnor U1473 (N_1473,In_310,In_2280);
and U1474 (N_1474,In_1390,In_885);
xor U1475 (N_1475,In_1215,In_2088);
xnor U1476 (N_1476,In_1106,In_474);
xor U1477 (N_1477,In_1571,In_2345);
nand U1478 (N_1478,In_1893,In_1890);
or U1479 (N_1479,In_2180,In_601);
nor U1480 (N_1480,In_681,In_457);
xnor U1481 (N_1481,In_103,In_757);
and U1482 (N_1482,In_1827,In_694);
nor U1483 (N_1483,In_792,In_1553);
or U1484 (N_1484,In_1551,In_2327);
nand U1485 (N_1485,In_2399,In_2029);
nand U1486 (N_1486,In_1990,In_2083);
xnor U1487 (N_1487,In_1354,In_1149);
xor U1488 (N_1488,In_1286,In_910);
xor U1489 (N_1489,In_1786,In_1244);
and U1490 (N_1490,In_615,In_592);
and U1491 (N_1491,In_1181,In_1457);
nand U1492 (N_1492,In_1302,In_998);
xnor U1493 (N_1493,In_832,In_190);
nor U1494 (N_1494,In_452,In_1507);
nor U1495 (N_1495,In_2096,In_739);
or U1496 (N_1496,In_532,In_1702);
xnor U1497 (N_1497,In_1253,In_150);
or U1498 (N_1498,In_1483,In_1883);
or U1499 (N_1499,In_2274,In_636);
nand U1500 (N_1500,In_571,In_2241);
nor U1501 (N_1501,In_1909,In_1771);
or U1502 (N_1502,In_1465,In_2350);
and U1503 (N_1503,In_21,In_1123);
nand U1504 (N_1504,In_2345,In_1629);
or U1505 (N_1505,In_2142,In_1166);
nand U1506 (N_1506,In_1760,In_1715);
and U1507 (N_1507,In_2262,In_2178);
and U1508 (N_1508,In_2121,In_571);
or U1509 (N_1509,In_1839,In_1058);
or U1510 (N_1510,In_887,In_519);
nor U1511 (N_1511,In_706,In_1667);
and U1512 (N_1512,In_6,In_1206);
and U1513 (N_1513,In_1255,In_978);
or U1514 (N_1514,In_299,In_2410);
nor U1515 (N_1515,In_732,In_1570);
xor U1516 (N_1516,In_1453,In_1060);
or U1517 (N_1517,In_470,In_1457);
or U1518 (N_1518,In_2301,In_768);
nand U1519 (N_1519,In_1074,In_936);
and U1520 (N_1520,In_572,In_417);
or U1521 (N_1521,In_1851,In_1440);
nand U1522 (N_1522,In_991,In_607);
nor U1523 (N_1523,In_1825,In_1808);
xnor U1524 (N_1524,In_2226,In_936);
nand U1525 (N_1525,In_450,In_2376);
xnor U1526 (N_1526,In_59,In_309);
and U1527 (N_1527,In_846,In_1732);
xor U1528 (N_1528,In_692,In_1343);
and U1529 (N_1529,In_1152,In_247);
nand U1530 (N_1530,In_655,In_1654);
or U1531 (N_1531,In_588,In_1115);
nand U1532 (N_1532,In_925,In_667);
nor U1533 (N_1533,In_508,In_1194);
nor U1534 (N_1534,In_906,In_1672);
and U1535 (N_1535,In_867,In_1779);
nand U1536 (N_1536,In_574,In_1384);
nor U1537 (N_1537,In_1591,In_219);
nand U1538 (N_1538,In_512,In_1025);
nand U1539 (N_1539,In_1068,In_1186);
nand U1540 (N_1540,In_861,In_303);
or U1541 (N_1541,In_1104,In_2319);
nand U1542 (N_1542,In_2082,In_749);
and U1543 (N_1543,In_2120,In_1698);
nor U1544 (N_1544,In_897,In_448);
and U1545 (N_1545,In_1519,In_193);
nor U1546 (N_1546,In_414,In_1536);
or U1547 (N_1547,In_2166,In_1220);
xnor U1548 (N_1548,In_471,In_846);
nand U1549 (N_1549,In_57,In_1548);
nand U1550 (N_1550,In_1773,In_1722);
xor U1551 (N_1551,In_2433,In_2156);
xor U1552 (N_1552,In_1074,In_165);
xor U1553 (N_1553,In_1121,In_2454);
nor U1554 (N_1554,In_829,In_2268);
or U1555 (N_1555,In_291,In_132);
and U1556 (N_1556,In_1528,In_1666);
nand U1557 (N_1557,In_575,In_2072);
and U1558 (N_1558,In_624,In_2414);
or U1559 (N_1559,In_2397,In_995);
or U1560 (N_1560,In_963,In_810);
or U1561 (N_1561,In_1179,In_1161);
or U1562 (N_1562,In_686,In_2241);
and U1563 (N_1563,In_2498,In_1233);
xor U1564 (N_1564,In_977,In_1515);
nor U1565 (N_1565,In_501,In_1207);
and U1566 (N_1566,In_1661,In_780);
nor U1567 (N_1567,In_2329,In_1805);
or U1568 (N_1568,In_870,In_530);
xnor U1569 (N_1569,In_276,In_2418);
or U1570 (N_1570,In_419,In_1);
or U1571 (N_1571,In_5,In_571);
xor U1572 (N_1572,In_240,In_168);
nand U1573 (N_1573,In_2113,In_2140);
xnor U1574 (N_1574,In_703,In_722);
or U1575 (N_1575,In_2323,In_1511);
nand U1576 (N_1576,In_2227,In_763);
nor U1577 (N_1577,In_1932,In_550);
nor U1578 (N_1578,In_1043,In_78);
or U1579 (N_1579,In_597,In_520);
xnor U1580 (N_1580,In_1688,In_1164);
nand U1581 (N_1581,In_1172,In_1229);
and U1582 (N_1582,In_1285,In_1207);
nor U1583 (N_1583,In_938,In_784);
and U1584 (N_1584,In_186,In_1811);
nand U1585 (N_1585,In_402,In_1638);
or U1586 (N_1586,In_308,In_118);
nor U1587 (N_1587,In_1282,In_383);
or U1588 (N_1588,In_1121,In_1681);
xnor U1589 (N_1589,In_2181,In_749);
and U1590 (N_1590,In_1844,In_1002);
xor U1591 (N_1591,In_2310,In_1070);
or U1592 (N_1592,In_2413,In_302);
and U1593 (N_1593,In_1418,In_1884);
xnor U1594 (N_1594,In_707,In_2457);
nor U1595 (N_1595,In_887,In_2056);
xnor U1596 (N_1596,In_1476,In_1827);
xnor U1597 (N_1597,In_2121,In_472);
nand U1598 (N_1598,In_1939,In_225);
xor U1599 (N_1599,In_32,In_1660);
xnor U1600 (N_1600,In_465,In_1323);
and U1601 (N_1601,In_1951,In_662);
nor U1602 (N_1602,In_59,In_268);
and U1603 (N_1603,In_371,In_2458);
xor U1604 (N_1604,In_2443,In_2094);
nor U1605 (N_1605,In_1487,In_1151);
or U1606 (N_1606,In_472,In_956);
nand U1607 (N_1607,In_767,In_282);
or U1608 (N_1608,In_578,In_824);
or U1609 (N_1609,In_2273,In_2090);
xor U1610 (N_1610,In_828,In_52);
nor U1611 (N_1611,In_1668,In_1907);
or U1612 (N_1612,In_798,In_1740);
xor U1613 (N_1613,In_627,In_1856);
nor U1614 (N_1614,In_1103,In_1976);
nor U1615 (N_1615,In_2287,In_1800);
and U1616 (N_1616,In_663,In_409);
nand U1617 (N_1617,In_1554,In_788);
nand U1618 (N_1618,In_780,In_1677);
or U1619 (N_1619,In_1173,In_2317);
or U1620 (N_1620,In_1313,In_2429);
nor U1621 (N_1621,In_917,In_1716);
nor U1622 (N_1622,In_1484,In_1121);
and U1623 (N_1623,In_2419,In_2404);
or U1624 (N_1624,In_696,In_121);
nor U1625 (N_1625,In_1941,In_80);
xor U1626 (N_1626,In_1078,In_755);
or U1627 (N_1627,In_956,In_1821);
xor U1628 (N_1628,In_163,In_313);
nand U1629 (N_1629,In_336,In_898);
xor U1630 (N_1630,In_786,In_2453);
nand U1631 (N_1631,In_1682,In_451);
or U1632 (N_1632,In_1229,In_730);
nand U1633 (N_1633,In_495,In_1199);
and U1634 (N_1634,In_1894,In_1191);
nor U1635 (N_1635,In_512,In_486);
nor U1636 (N_1636,In_1711,In_1026);
and U1637 (N_1637,In_1747,In_66);
or U1638 (N_1638,In_62,In_861);
or U1639 (N_1639,In_792,In_19);
nor U1640 (N_1640,In_722,In_1878);
or U1641 (N_1641,In_2053,In_1406);
and U1642 (N_1642,In_1450,In_2229);
nor U1643 (N_1643,In_475,In_1340);
nand U1644 (N_1644,In_2399,In_1852);
and U1645 (N_1645,In_1577,In_1599);
nor U1646 (N_1646,In_2035,In_220);
xor U1647 (N_1647,In_764,In_397);
xor U1648 (N_1648,In_2057,In_1153);
and U1649 (N_1649,In_1936,In_239);
nand U1650 (N_1650,In_990,In_35);
nand U1651 (N_1651,In_265,In_1406);
xor U1652 (N_1652,In_386,In_766);
nand U1653 (N_1653,In_2087,In_1957);
or U1654 (N_1654,In_47,In_1562);
nor U1655 (N_1655,In_810,In_1184);
or U1656 (N_1656,In_1126,In_1387);
xnor U1657 (N_1657,In_624,In_2254);
xor U1658 (N_1658,In_881,In_38);
nor U1659 (N_1659,In_332,In_1086);
or U1660 (N_1660,In_1592,In_1273);
nor U1661 (N_1661,In_2217,In_1517);
xnor U1662 (N_1662,In_1356,In_80);
or U1663 (N_1663,In_1972,In_2152);
nand U1664 (N_1664,In_27,In_410);
xor U1665 (N_1665,In_395,In_285);
xnor U1666 (N_1666,In_2332,In_2083);
nor U1667 (N_1667,In_1538,In_112);
xnor U1668 (N_1668,In_123,In_601);
nor U1669 (N_1669,In_321,In_2007);
or U1670 (N_1670,In_2499,In_1523);
and U1671 (N_1671,In_2418,In_831);
and U1672 (N_1672,In_877,In_1232);
and U1673 (N_1673,In_1271,In_677);
and U1674 (N_1674,In_1601,In_2411);
xor U1675 (N_1675,In_1933,In_2094);
or U1676 (N_1676,In_1210,In_1077);
nor U1677 (N_1677,In_2231,In_1663);
and U1678 (N_1678,In_1138,In_2044);
and U1679 (N_1679,In_42,In_2299);
nand U1680 (N_1680,In_944,In_1376);
or U1681 (N_1681,In_2054,In_2243);
or U1682 (N_1682,In_736,In_290);
xor U1683 (N_1683,In_2286,In_542);
or U1684 (N_1684,In_955,In_535);
nor U1685 (N_1685,In_1782,In_637);
and U1686 (N_1686,In_376,In_944);
nor U1687 (N_1687,In_149,In_701);
nor U1688 (N_1688,In_1370,In_1340);
and U1689 (N_1689,In_716,In_1313);
or U1690 (N_1690,In_1861,In_797);
xor U1691 (N_1691,In_2013,In_2000);
xnor U1692 (N_1692,In_1236,In_1943);
nand U1693 (N_1693,In_75,In_1931);
nand U1694 (N_1694,In_2203,In_2273);
or U1695 (N_1695,In_347,In_1872);
nor U1696 (N_1696,In_493,In_1034);
nor U1697 (N_1697,In_949,In_2090);
nand U1698 (N_1698,In_1433,In_2399);
nor U1699 (N_1699,In_1043,In_2056);
nand U1700 (N_1700,In_524,In_1078);
nor U1701 (N_1701,In_121,In_671);
nand U1702 (N_1702,In_374,In_1059);
nand U1703 (N_1703,In_1580,In_1888);
and U1704 (N_1704,In_1108,In_588);
xor U1705 (N_1705,In_1461,In_1034);
or U1706 (N_1706,In_1623,In_1549);
nor U1707 (N_1707,In_1349,In_1828);
or U1708 (N_1708,In_2399,In_1506);
xnor U1709 (N_1709,In_2267,In_1253);
xor U1710 (N_1710,In_1018,In_1233);
nand U1711 (N_1711,In_2198,In_364);
and U1712 (N_1712,In_431,In_1505);
nor U1713 (N_1713,In_1848,In_2404);
nor U1714 (N_1714,In_1088,In_428);
nor U1715 (N_1715,In_1485,In_198);
and U1716 (N_1716,In_1051,In_972);
and U1717 (N_1717,In_355,In_535);
and U1718 (N_1718,In_1531,In_1611);
xor U1719 (N_1719,In_1127,In_380);
or U1720 (N_1720,In_594,In_605);
or U1721 (N_1721,In_461,In_2067);
and U1722 (N_1722,In_475,In_1362);
and U1723 (N_1723,In_2457,In_353);
or U1724 (N_1724,In_1402,In_19);
nand U1725 (N_1725,In_1998,In_984);
and U1726 (N_1726,In_1189,In_1852);
or U1727 (N_1727,In_558,In_256);
and U1728 (N_1728,In_2101,In_627);
xor U1729 (N_1729,In_602,In_1317);
xnor U1730 (N_1730,In_1891,In_958);
and U1731 (N_1731,In_1799,In_1938);
nand U1732 (N_1732,In_976,In_567);
or U1733 (N_1733,In_1136,In_1810);
nand U1734 (N_1734,In_941,In_1329);
xor U1735 (N_1735,In_121,In_629);
or U1736 (N_1736,In_550,In_433);
or U1737 (N_1737,In_1300,In_178);
nor U1738 (N_1738,In_2283,In_910);
or U1739 (N_1739,In_476,In_1754);
or U1740 (N_1740,In_1852,In_988);
nor U1741 (N_1741,In_2200,In_503);
nor U1742 (N_1742,In_1563,In_1870);
and U1743 (N_1743,In_2186,In_1848);
xor U1744 (N_1744,In_1608,In_2003);
or U1745 (N_1745,In_1462,In_1190);
xor U1746 (N_1746,In_2493,In_121);
or U1747 (N_1747,In_2246,In_842);
or U1748 (N_1748,In_1428,In_2288);
or U1749 (N_1749,In_1688,In_1307);
and U1750 (N_1750,In_1532,In_2414);
nor U1751 (N_1751,In_546,In_763);
or U1752 (N_1752,In_1919,In_1891);
nand U1753 (N_1753,In_2111,In_1999);
xor U1754 (N_1754,In_2198,In_987);
nand U1755 (N_1755,In_803,In_579);
nor U1756 (N_1756,In_1100,In_1524);
and U1757 (N_1757,In_871,In_250);
xor U1758 (N_1758,In_634,In_1533);
or U1759 (N_1759,In_259,In_1324);
nand U1760 (N_1760,In_1837,In_2464);
and U1761 (N_1761,In_161,In_2174);
xnor U1762 (N_1762,In_908,In_2463);
nand U1763 (N_1763,In_1519,In_1537);
nand U1764 (N_1764,In_1768,In_1514);
or U1765 (N_1765,In_906,In_1566);
nand U1766 (N_1766,In_2175,In_1911);
or U1767 (N_1767,In_1823,In_636);
nand U1768 (N_1768,In_498,In_353);
xnor U1769 (N_1769,In_1716,In_219);
or U1770 (N_1770,In_2126,In_779);
or U1771 (N_1771,In_1040,In_838);
and U1772 (N_1772,In_2225,In_84);
and U1773 (N_1773,In_669,In_2430);
nor U1774 (N_1774,In_1596,In_1703);
nor U1775 (N_1775,In_424,In_523);
xor U1776 (N_1776,In_2021,In_1042);
and U1777 (N_1777,In_2204,In_986);
nand U1778 (N_1778,In_1865,In_1601);
xor U1779 (N_1779,In_1017,In_34);
or U1780 (N_1780,In_868,In_2464);
nor U1781 (N_1781,In_1451,In_1185);
and U1782 (N_1782,In_2364,In_308);
xor U1783 (N_1783,In_1416,In_2143);
and U1784 (N_1784,In_336,In_758);
nor U1785 (N_1785,In_935,In_67);
nand U1786 (N_1786,In_2116,In_860);
nor U1787 (N_1787,In_1598,In_64);
xnor U1788 (N_1788,In_1626,In_2163);
nor U1789 (N_1789,In_2414,In_2290);
or U1790 (N_1790,In_369,In_267);
xor U1791 (N_1791,In_197,In_1645);
or U1792 (N_1792,In_736,In_1247);
nor U1793 (N_1793,In_1632,In_2192);
xor U1794 (N_1794,In_533,In_1834);
xnor U1795 (N_1795,In_907,In_2468);
nand U1796 (N_1796,In_981,In_2426);
nand U1797 (N_1797,In_1876,In_1671);
nand U1798 (N_1798,In_1839,In_354);
or U1799 (N_1799,In_1414,In_423);
nor U1800 (N_1800,In_1662,In_1615);
or U1801 (N_1801,In_1653,In_1901);
nand U1802 (N_1802,In_146,In_1446);
nor U1803 (N_1803,In_2319,In_2481);
and U1804 (N_1804,In_86,In_2323);
xor U1805 (N_1805,In_216,In_2243);
or U1806 (N_1806,In_2103,In_1128);
and U1807 (N_1807,In_650,In_1593);
xnor U1808 (N_1808,In_554,In_1459);
nand U1809 (N_1809,In_469,In_1195);
and U1810 (N_1810,In_86,In_736);
xor U1811 (N_1811,In_1750,In_1764);
nor U1812 (N_1812,In_2482,In_1354);
and U1813 (N_1813,In_19,In_1114);
or U1814 (N_1814,In_775,In_1454);
nand U1815 (N_1815,In_1744,In_2201);
nor U1816 (N_1816,In_1807,In_1178);
xor U1817 (N_1817,In_322,In_2097);
and U1818 (N_1818,In_210,In_1816);
and U1819 (N_1819,In_999,In_1088);
and U1820 (N_1820,In_1959,In_963);
nand U1821 (N_1821,In_73,In_1948);
or U1822 (N_1822,In_2032,In_556);
and U1823 (N_1823,In_104,In_311);
xnor U1824 (N_1824,In_704,In_2357);
and U1825 (N_1825,In_456,In_1635);
or U1826 (N_1826,In_1318,In_1436);
nor U1827 (N_1827,In_1081,In_2165);
or U1828 (N_1828,In_749,In_948);
nand U1829 (N_1829,In_1448,In_1413);
xnor U1830 (N_1830,In_612,In_213);
and U1831 (N_1831,In_418,In_366);
and U1832 (N_1832,In_943,In_208);
or U1833 (N_1833,In_1147,In_952);
nor U1834 (N_1834,In_505,In_1398);
or U1835 (N_1835,In_2287,In_986);
and U1836 (N_1836,In_578,In_138);
and U1837 (N_1837,In_23,In_1273);
nor U1838 (N_1838,In_20,In_768);
and U1839 (N_1839,In_952,In_2109);
and U1840 (N_1840,In_1096,In_155);
or U1841 (N_1841,In_463,In_2413);
nand U1842 (N_1842,In_1874,In_1484);
and U1843 (N_1843,In_2317,In_612);
or U1844 (N_1844,In_1425,In_1181);
and U1845 (N_1845,In_2455,In_2063);
xor U1846 (N_1846,In_1040,In_2397);
nor U1847 (N_1847,In_1805,In_924);
nor U1848 (N_1848,In_2365,In_356);
nor U1849 (N_1849,In_1541,In_1274);
nand U1850 (N_1850,In_893,In_326);
or U1851 (N_1851,In_2451,In_2410);
nand U1852 (N_1852,In_1875,In_147);
or U1853 (N_1853,In_1647,In_121);
nand U1854 (N_1854,In_53,In_475);
and U1855 (N_1855,In_1192,In_321);
xor U1856 (N_1856,In_1373,In_1673);
xnor U1857 (N_1857,In_653,In_2026);
nor U1858 (N_1858,In_1157,In_2216);
nand U1859 (N_1859,In_2332,In_629);
or U1860 (N_1860,In_630,In_632);
xnor U1861 (N_1861,In_1449,In_548);
nand U1862 (N_1862,In_1522,In_1485);
nor U1863 (N_1863,In_1954,In_317);
xor U1864 (N_1864,In_1684,In_1588);
nor U1865 (N_1865,In_2009,In_688);
xor U1866 (N_1866,In_71,In_1849);
nand U1867 (N_1867,In_376,In_1434);
nand U1868 (N_1868,In_776,In_1205);
and U1869 (N_1869,In_2035,In_1150);
xor U1870 (N_1870,In_1439,In_155);
nor U1871 (N_1871,In_1962,In_1792);
nand U1872 (N_1872,In_655,In_2126);
xor U1873 (N_1873,In_1836,In_2224);
nand U1874 (N_1874,In_1134,In_2378);
xor U1875 (N_1875,In_1938,In_730);
or U1876 (N_1876,In_2421,In_1422);
or U1877 (N_1877,In_395,In_1592);
xnor U1878 (N_1878,In_2435,In_1286);
and U1879 (N_1879,In_861,In_840);
and U1880 (N_1880,In_363,In_707);
nor U1881 (N_1881,In_551,In_1959);
nor U1882 (N_1882,In_1891,In_2205);
and U1883 (N_1883,In_642,In_837);
nor U1884 (N_1884,In_1053,In_2025);
or U1885 (N_1885,In_1924,In_103);
nor U1886 (N_1886,In_2466,In_315);
xor U1887 (N_1887,In_2492,In_1870);
xnor U1888 (N_1888,In_1279,In_43);
and U1889 (N_1889,In_1393,In_1010);
nor U1890 (N_1890,In_1092,In_1758);
nand U1891 (N_1891,In_1475,In_1109);
nand U1892 (N_1892,In_1003,In_2315);
xor U1893 (N_1893,In_1670,In_1262);
or U1894 (N_1894,In_101,In_765);
or U1895 (N_1895,In_512,In_1106);
nor U1896 (N_1896,In_2130,In_1918);
or U1897 (N_1897,In_723,In_237);
nand U1898 (N_1898,In_806,In_1904);
or U1899 (N_1899,In_2469,In_954);
and U1900 (N_1900,In_1223,In_1911);
and U1901 (N_1901,In_1786,In_292);
nand U1902 (N_1902,In_3,In_2356);
xor U1903 (N_1903,In_1298,In_1170);
xnor U1904 (N_1904,In_348,In_84);
nand U1905 (N_1905,In_19,In_2235);
or U1906 (N_1906,In_1834,In_1128);
and U1907 (N_1907,In_1272,In_465);
nor U1908 (N_1908,In_208,In_50);
xor U1909 (N_1909,In_699,In_296);
xnor U1910 (N_1910,In_295,In_949);
nand U1911 (N_1911,In_2309,In_917);
xor U1912 (N_1912,In_2209,In_823);
nor U1913 (N_1913,In_1467,In_2317);
nand U1914 (N_1914,In_602,In_194);
nand U1915 (N_1915,In_2128,In_35);
nor U1916 (N_1916,In_176,In_1180);
xnor U1917 (N_1917,In_1632,In_2485);
nor U1918 (N_1918,In_888,In_1176);
nand U1919 (N_1919,In_1701,In_2162);
or U1920 (N_1920,In_1163,In_2041);
and U1921 (N_1921,In_2465,In_2031);
and U1922 (N_1922,In_877,In_1025);
nand U1923 (N_1923,In_1439,In_2083);
or U1924 (N_1924,In_949,In_2042);
or U1925 (N_1925,In_1854,In_1750);
and U1926 (N_1926,In_1335,In_2011);
and U1927 (N_1927,In_720,In_1089);
or U1928 (N_1928,In_2098,In_398);
xnor U1929 (N_1929,In_1940,In_439);
or U1930 (N_1930,In_1984,In_1059);
and U1931 (N_1931,In_52,In_816);
nand U1932 (N_1932,In_201,In_2244);
and U1933 (N_1933,In_1656,In_989);
or U1934 (N_1934,In_1670,In_1855);
or U1935 (N_1935,In_1609,In_1176);
nand U1936 (N_1936,In_27,In_429);
and U1937 (N_1937,In_564,In_709);
xnor U1938 (N_1938,In_1573,In_1529);
nor U1939 (N_1939,In_1562,In_1305);
and U1940 (N_1940,In_149,In_94);
or U1941 (N_1941,In_1872,In_2412);
and U1942 (N_1942,In_132,In_883);
nand U1943 (N_1943,In_1691,In_2306);
xor U1944 (N_1944,In_60,In_467);
xnor U1945 (N_1945,In_1724,In_943);
and U1946 (N_1946,In_2069,In_244);
or U1947 (N_1947,In_415,In_1246);
xnor U1948 (N_1948,In_1891,In_859);
xnor U1949 (N_1949,In_344,In_1494);
xnor U1950 (N_1950,In_2143,In_486);
xor U1951 (N_1951,In_922,In_980);
and U1952 (N_1952,In_2276,In_164);
or U1953 (N_1953,In_2146,In_1411);
and U1954 (N_1954,In_1768,In_1115);
xnor U1955 (N_1955,In_1758,In_381);
and U1956 (N_1956,In_2253,In_2076);
or U1957 (N_1957,In_865,In_1748);
nor U1958 (N_1958,In_1437,In_2337);
nand U1959 (N_1959,In_1370,In_763);
nand U1960 (N_1960,In_393,In_841);
nor U1961 (N_1961,In_1426,In_1699);
nand U1962 (N_1962,In_2070,In_626);
or U1963 (N_1963,In_2085,In_1323);
or U1964 (N_1964,In_93,In_503);
nor U1965 (N_1965,In_2279,In_271);
xnor U1966 (N_1966,In_1647,In_694);
xnor U1967 (N_1967,In_757,In_921);
or U1968 (N_1968,In_1394,In_1987);
or U1969 (N_1969,In_2238,In_1196);
xor U1970 (N_1970,In_1341,In_2037);
xor U1971 (N_1971,In_260,In_2365);
nor U1972 (N_1972,In_1664,In_1943);
or U1973 (N_1973,In_1135,In_1260);
xor U1974 (N_1974,In_2403,In_655);
xnor U1975 (N_1975,In_231,In_1127);
nand U1976 (N_1976,In_1810,In_1080);
and U1977 (N_1977,In_2361,In_1490);
or U1978 (N_1978,In_347,In_895);
or U1979 (N_1979,In_687,In_321);
nor U1980 (N_1980,In_844,In_318);
xor U1981 (N_1981,In_674,In_610);
and U1982 (N_1982,In_507,In_1720);
xnor U1983 (N_1983,In_1159,In_422);
nor U1984 (N_1984,In_828,In_604);
and U1985 (N_1985,In_2365,In_776);
nor U1986 (N_1986,In_927,In_975);
and U1987 (N_1987,In_1351,In_1381);
or U1988 (N_1988,In_1822,In_1742);
and U1989 (N_1989,In_682,In_166);
and U1990 (N_1990,In_1182,In_1862);
nand U1991 (N_1991,In_2364,In_800);
nand U1992 (N_1992,In_2101,In_1735);
and U1993 (N_1993,In_1724,In_246);
and U1994 (N_1994,In_2263,In_1847);
nand U1995 (N_1995,In_989,In_1810);
nand U1996 (N_1996,In_972,In_210);
nand U1997 (N_1997,In_1119,In_2027);
nand U1998 (N_1998,In_2246,In_1286);
xnor U1999 (N_1999,In_946,In_1073);
xor U2000 (N_2000,In_1353,In_1456);
or U2001 (N_2001,In_135,In_328);
xor U2002 (N_2002,In_208,In_1981);
nand U2003 (N_2003,In_2363,In_1006);
and U2004 (N_2004,In_936,In_90);
and U2005 (N_2005,In_1208,In_2131);
and U2006 (N_2006,In_264,In_495);
or U2007 (N_2007,In_1505,In_2270);
nand U2008 (N_2008,In_2001,In_786);
and U2009 (N_2009,In_143,In_2358);
nor U2010 (N_2010,In_784,In_2493);
or U2011 (N_2011,In_1178,In_1527);
or U2012 (N_2012,In_1079,In_2093);
nand U2013 (N_2013,In_663,In_1056);
nand U2014 (N_2014,In_983,In_1076);
nor U2015 (N_2015,In_2350,In_1885);
xnor U2016 (N_2016,In_767,In_1831);
nor U2017 (N_2017,In_2161,In_484);
and U2018 (N_2018,In_376,In_1225);
and U2019 (N_2019,In_285,In_1164);
nand U2020 (N_2020,In_940,In_766);
nor U2021 (N_2021,In_2119,In_322);
nor U2022 (N_2022,In_243,In_301);
nand U2023 (N_2023,In_1654,In_52);
and U2024 (N_2024,In_875,In_785);
or U2025 (N_2025,In_1024,In_1795);
and U2026 (N_2026,In_768,In_2136);
nand U2027 (N_2027,In_2133,In_1209);
or U2028 (N_2028,In_452,In_1962);
xor U2029 (N_2029,In_635,In_2036);
or U2030 (N_2030,In_1990,In_1618);
and U2031 (N_2031,In_1995,In_851);
nor U2032 (N_2032,In_534,In_1015);
nand U2033 (N_2033,In_8,In_1298);
nor U2034 (N_2034,In_546,In_794);
and U2035 (N_2035,In_2095,In_817);
nor U2036 (N_2036,In_574,In_981);
xor U2037 (N_2037,In_2310,In_1864);
nor U2038 (N_2038,In_1229,In_934);
nand U2039 (N_2039,In_1260,In_431);
and U2040 (N_2040,In_309,In_368);
or U2041 (N_2041,In_580,In_444);
xor U2042 (N_2042,In_75,In_2437);
xnor U2043 (N_2043,In_32,In_1107);
nor U2044 (N_2044,In_416,In_2429);
or U2045 (N_2045,In_613,In_329);
and U2046 (N_2046,In_419,In_1033);
and U2047 (N_2047,In_413,In_2482);
nand U2048 (N_2048,In_1839,In_1385);
nor U2049 (N_2049,In_1332,In_886);
xor U2050 (N_2050,In_2374,In_1318);
nand U2051 (N_2051,In_2156,In_1393);
and U2052 (N_2052,In_1068,In_1602);
nand U2053 (N_2053,In_1400,In_894);
xor U2054 (N_2054,In_2127,In_184);
or U2055 (N_2055,In_1051,In_2221);
and U2056 (N_2056,In_306,In_939);
or U2057 (N_2057,In_1217,In_1060);
nor U2058 (N_2058,In_1689,In_574);
or U2059 (N_2059,In_1341,In_858);
and U2060 (N_2060,In_477,In_975);
or U2061 (N_2061,In_1501,In_1076);
and U2062 (N_2062,In_453,In_1933);
nor U2063 (N_2063,In_2217,In_641);
nand U2064 (N_2064,In_1325,In_1272);
nand U2065 (N_2065,In_618,In_1288);
xnor U2066 (N_2066,In_1036,In_1506);
or U2067 (N_2067,In_2364,In_535);
nand U2068 (N_2068,In_1606,In_2306);
nor U2069 (N_2069,In_610,In_1836);
xnor U2070 (N_2070,In_1118,In_1447);
nand U2071 (N_2071,In_2186,In_1266);
nand U2072 (N_2072,In_1221,In_724);
and U2073 (N_2073,In_1840,In_894);
nand U2074 (N_2074,In_2291,In_765);
and U2075 (N_2075,In_2313,In_931);
and U2076 (N_2076,In_1450,In_1072);
nand U2077 (N_2077,In_1507,In_2496);
nand U2078 (N_2078,In_829,In_1467);
nand U2079 (N_2079,In_254,In_1002);
nor U2080 (N_2080,In_1569,In_1526);
and U2081 (N_2081,In_1012,In_2386);
nand U2082 (N_2082,In_654,In_625);
nand U2083 (N_2083,In_1200,In_192);
or U2084 (N_2084,In_651,In_948);
and U2085 (N_2085,In_1601,In_2103);
and U2086 (N_2086,In_1577,In_2196);
and U2087 (N_2087,In_38,In_417);
xor U2088 (N_2088,In_1454,In_2438);
nand U2089 (N_2089,In_1895,In_373);
and U2090 (N_2090,In_997,In_1748);
or U2091 (N_2091,In_1616,In_1800);
nor U2092 (N_2092,In_1946,In_509);
nor U2093 (N_2093,In_2185,In_1808);
nor U2094 (N_2094,In_1089,In_485);
nor U2095 (N_2095,In_403,In_602);
nor U2096 (N_2096,In_2044,In_1997);
and U2097 (N_2097,In_2013,In_327);
nor U2098 (N_2098,In_929,In_1359);
and U2099 (N_2099,In_1556,In_2288);
nand U2100 (N_2100,In_516,In_1998);
and U2101 (N_2101,In_1074,In_533);
xor U2102 (N_2102,In_2252,In_2498);
xor U2103 (N_2103,In_2311,In_2226);
or U2104 (N_2104,In_1660,In_733);
and U2105 (N_2105,In_710,In_2196);
nor U2106 (N_2106,In_271,In_640);
and U2107 (N_2107,In_783,In_1655);
or U2108 (N_2108,In_110,In_1816);
nor U2109 (N_2109,In_357,In_1662);
or U2110 (N_2110,In_2351,In_1908);
and U2111 (N_2111,In_1286,In_1304);
and U2112 (N_2112,In_729,In_577);
and U2113 (N_2113,In_1622,In_621);
or U2114 (N_2114,In_974,In_449);
xnor U2115 (N_2115,In_1202,In_1901);
xor U2116 (N_2116,In_1380,In_180);
and U2117 (N_2117,In_1922,In_591);
xor U2118 (N_2118,In_459,In_213);
nor U2119 (N_2119,In_407,In_1655);
nor U2120 (N_2120,In_109,In_1423);
xnor U2121 (N_2121,In_37,In_1861);
and U2122 (N_2122,In_684,In_2019);
nor U2123 (N_2123,In_333,In_1630);
nor U2124 (N_2124,In_1664,In_1179);
and U2125 (N_2125,In_402,In_1397);
nor U2126 (N_2126,In_1954,In_1188);
nand U2127 (N_2127,In_1057,In_1980);
or U2128 (N_2128,In_2312,In_2294);
or U2129 (N_2129,In_2018,In_223);
xnor U2130 (N_2130,In_2150,In_1130);
nor U2131 (N_2131,In_128,In_330);
xor U2132 (N_2132,In_1575,In_1930);
nand U2133 (N_2133,In_2204,In_513);
nor U2134 (N_2134,In_1945,In_1837);
and U2135 (N_2135,In_2044,In_1493);
and U2136 (N_2136,In_962,In_1722);
and U2137 (N_2137,In_1234,In_940);
xor U2138 (N_2138,In_1076,In_1761);
and U2139 (N_2139,In_2338,In_672);
nor U2140 (N_2140,In_1163,In_1301);
nand U2141 (N_2141,In_1782,In_2123);
or U2142 (N_2142,In_2459,In_2492);
nand U2143 (N_2143,In_646,In_1790);
nor U2144 (N_2144,In_2216,In_728);
nand U2145 (N_2145,In_1625,In_1880);
xnor U2146 (N_2146,In_1862,In_1334);
nor U2147 (N_2147,In_310,In_1569);
or U2148 (N_2148,In_197,In_941);
xnor U2149 (N_2149,In_2352,In_1818);
or U2150 (N_2150,In_915,In_825);
nor U2151 (N_2151,In_320,In_520);
and U2152 (N_2152,In_1904,In_2432);
nand U2153 (N_2153,In_1980,In_2125);
nor U2154 (N_2154,In_703,In_0);
xnor U2155 (N_2155,In_1563,In_230);
nand U2156 (N_2156,In_1592,In_422);
xnor U2157 (N_2157,In_1895,In_1069);
nor U2158 (N_2158,In_103,In_90);
xnor U2159 (N_2159,In_2122,In_533);
and U2160 (N_2160,In_2175,In_1047);
nand U2161 (N_2161,In_73,In_1080);
nor U2162 (N_2162,In_1490,In_850);
xor U2163 (N_2163,In_2391,In_858);
xnor U2164 (N_2164,In_558,In_1027);
or U2165 (N_2165,In_2024,In_636);
nand U2166 (N_2166,In_1595,In_969);
xnor U2167 (N_2167,In_1224,In_2424);
nand U2168 (N_2168,In_4,In_340);
nand U2169 (N_2169,In_1080,In_290);
nand U2170 (N_2170,In_1580,In_1132);
xor U2171 (N_2171,In_773,In_620);
nand U2172 (N_2172,In_1351,In_51);
or U2173 (N_2173,In_1868,In_1300);
nand U2174 (N_2174,In_1309,In_1184);
nor U2175 (N_2175,In_633,In_235);
nand U2176 (N_2176,In_2046,In_757);
or U2177 (N_2177,In_1604,In_1527);
and U2178 (N_2178,In_674,In_284);
nand U2179 (N_2179,In_2284,In_1132);
and U2180 (N_2180,In_1601,In_1676);
and U2181 (N_2181,In_201,In_1093);
nor U2182 (N_2182,In_2083,In_2328);
and U2183 (N_2183,In_525,In_2069);
xnor U2184 (N_2184,In_1834,In_2194);
or U2185 (N_2185,In_1529,In_740);
nor U2186 (N_2186,In_2191,In_1769);
nor U2187 (N_2187,In_1748,In_1591);
xnor U2188 (N_2188,In_526,In_634);
and U2189 (N_2189,In_198,In_2019);
and U2190 (N_2190,In_2472,In_1046);
xor U2191 (N_2191,In_2375,In_1912);
or U2192 (N_2192,In_1773,In_2114);
nand U2193 (N_2193,In_1576,In_697);
nor U2194 (N_2194,In_1208,In_1780);
xor U2195 (N_2195,In_784,In_2107);
xnor U2196 (N_2196,In_819,In_2138);
xor U2197 (N_2197,In_533,In_406);
nor U2198 (N_2198,In_1277,In_1710);
nand U2199 (N_2199,In_2182,In_1174);
or U2200 (N_2200,In_2240,In_708);
nor U2201 (N_2201,In_1574,In_1225);
or U2202 (N_2202,In_519,In_1143);
xor U2203 (N_2203,In_2216,In_586);
and U2204 (N_2204,In_719,In_1642);
or U2205 (N_2205,In_1168,In_1288);
or U2206 (N_2206,In_2092,In_2160);
and U2207 (N_2207,In_675,In_1395);
nand U2208 (N_2208,In_1661,In_359);
or U2209 (N_2209,In_1645,In_1902);
nor U2210 (N_2210,In_933,In_131);
and U2211 (N_2211,In_103,In_1953);
or U2212 (N_2212,In_1215,In_115);
nand U2213 (N_2213,In_1162,In_1943);
xor U2214 (N_2214,In_1558,In_1184);
nor U2215 (N_2215,In_1743,In_1575);
or U2216 (N_2216,In_1996,In_1076);
or U2217 (N_2217,In_1451,In_398);
xor U2218 (N_2218,In_1017,In_556);
nand U2219 (N_2219,In_520,In_395);
xor U2220 (N_2220,In_2390,In_1951);
xor U2221 (N_2221,In_728,In_1405);
nor U2222 (N_2222,In_1149,In_951);
and U2223 (N_2223,In_609,In_500);
and U2224 (N_2224,In_263,In_2088);
nor U2225 (N_2225,In_175,In_1688);
nand U2226 (N_2226,In_299,In_117);
and U2227 (N_2227,In_558,In_2121);
nand U2228 (N_2228,In_606,In_2386);
nand U2229 (N_2229,In_1549,In_1095);
or U2230 (N_2230,In_1592,In_491);
xor U2231 (N_2231,In_1524,In_1587);
nand U2232 (N_2232,In_1990,In_230);
xnor U2233 (N_2233,In_2290,In_136);
or U2234 (N_2234,In_1573,In_2125);
nor U2235 (N_2235,In_2054,In_1727);
and U2236 (N_2236,In_2368,In_2398);
nand U2237 (N_2237,In_540,In_2249);
nor U2238 (N_2238,In_1187,In_1318);
xnor U2239 (N_2239,In_868,In_915);
xor U2240 (N_2240,In_1296,In_2067);
and U2241 (N_2241,In_2459,In_1334);
nor U2242 (N_2242,In_1251,In_498);
nand U2243 (N_2243,In_2079,In_234);
xor U2244 (N_2244,In_1615,In_1369);
nand U2245 (N_2245,In_1964,In_834);
and U2246 (N_2246,In_1734,In_1160);
or U2247 (N_2247,In_1383,In_1609);
nand U2248 (N_2248,In_1056,In_2337);
or U2249 (N_2249,In_1797,In_2339);
or U2250 (N_2250,In_2475,In_785);
nor U2251 (N_2251,In_227,In_2351);
or U2252 (N_2252,In_193,In_1937);
xor U2253 (N_2253,In_426,In_2375);
and U2254 (N_2254,In_949,In_447);
nand U2255 (N_2255,In_1712,In_731);
xor U2256 (N_2256,In_1163,In_2369);
xnor U2257 (N_2257,In_182,In_2463);
and U2258 (N_2258,In_615,In_635);
or U2259 (N_2259,In_1148,In_1926);
nor U2260 (N_2260,In_2238,In_730);
nand U2261 (N_2261,In_278,In_2349);
xor U2262 (N_2262,In_2346,In_151);
nor U2263 (N_2263,In_1667,In_492);
or U2264 (N_2264,In_1974,In_1741);
or U2265 (N_2265,In_1872,In_90);
nor U2266 (N_2266,In_493,In_119);
nor U2267 (N_2267,In_1530,In_426);
xor U2268 (N_2268,In_1670,In_2192);
xnor U2269 (N_2269,In_133,In_507);
nor U2270 (N_2270,In_2184,In_874);
nor U2271 (N_2271,In_1321,In_1481);
and U2272 (N_2272,In_1655,In_1856);
or U2273 (N_2273,In_553,In_2180);
xnor U2274 (N_2274,In_1451,In_7);
and U2275 (N_2275,In_1439,In_1034);
or U2276 (N_2276,In_936,In_900);
nand U2277 (N_2277,In_1070,In_2488);
nand U2278 (N_2278,In_2287,In_258);
xnor U2279 (N_2279,In_2042,In_2470);
nor U2280 (N_2280,In_1077,In_736);
nor U2281 (N_2281,In_1399,In_425);
and U2282 (N_2282,In_1655,In_535);
nor U2283 (N_2283,In_1054,In_1485);
nand U2284 (N_2284,In_1807,In_1768);
nor U2285 (N_2285,In_116,In_1158);
and U2286 (N_2286,In_1944,In_2391);
xnor U2287 (N_2287,In_717,In_1954);
nor U2288 (N_2288,In_433,In_1970);
or U2289 (N_2289,In_2307,In_1914);
or U2290 (N_2290,In_1913,In_2282);
nor U2291 (N_2291,In_2341,In_582);
and U2292 (N_2292,In_878,In_1476);
nand U2293 (N_2293,In_1942,In_1540);
nor U2294 (N_2294,In_2219,In_466);
or U2295 (N_2295,In_272,In_195);
or U2296 (N_2296,In_621,In_2455);
or U2297 (N_2297,In_2445,In_1622);
and U2298 (N_2298,In_2189,In_1856);
xnor U2299 (N_2299,In_1839,In_355);
or U2300 (N_2300,In_44,In_882);
and U2301 (N_2301,In_2312,In_327);
or U2302 (N_2302,In_1539,In_1925);
xor U2303 (N_2303,In_1052,In_953);
nand U2304 (N_2304,In_251,In_2398);
nand U2305 (N_2305,In_2080,In_1685);
nor U2306 (N_2306,In_2343,In_1129);
or U2307 (N_2307,In_1179,In_412);
nor U2308 (N_2308,In_2016,In_772);
and U2309 (N_2309,In_510,In_1785);
nor U2310 (N_2310,In_1507,In_248);
xor U2311 (N_2311,In_1238,In_815);
and U2312 (N_2312,In_1321,In_2037);
or U2313 (N_2313,In_1428,In_740);
nand U2314 (N_2314,In_2025,In_2099);
xnor U2315 (N_2315,In_1440,In_1503);
xnor U2316 (N_2316,In_1075,In_516);
nor U2317 (N_2317,In_1691,In_1198);
and U2318 (N_2318,In_2144,In_1867);
xnor U2319 (N_2319,In_32,In_840);
or U2320 (N_2320,In_2395,In_329);
or U2321 (N_2321,In_288,In_1469);
and U2322 (N_2322,In_744,In_1498);
nand U2323 (N_2323,In_1477,In_249);
nor U2324 (N_2324,In_2444,In_2204);
xnor U2325 (N_2325,In_2071,In_2187);
nand U2326 (N_2326,In_1262,In_2168);
xor U2327 (N_2327,In_2447,In_1280);
or U2328 (N_2328,In_2048,In_1560);
xor U2329 (N_2329,In_1767,In_2466);
and U2330 (N_2330,In_594,In_475);
or U2331 (N_2331,In_1610,In_1086);
nor U2332 (N_2332,In_1515,In_1960);
xor U2333 (N_2333,In_1606,In_1087);
nand U2334 (N_2334,In_370,In_915);
or U2335 (N_2335,In_1262,In_379);
xor U2336 (N_2336,In_102,In_1747);
nand U2337 (N_2337,In_1120,In_988);
and U2338 (N_2338,In_2419,In_1700);
xor U2339 (N_2339,In_2185,In_67);
nand U2340 (N_2340,In_442,In_2270);
and U2341 (N_2341,In_404,In_1570);
or U2342 (N_2342,In_589,In_2000);
or U2343 (N_2343,In_965,In_2127);
nand U2344 (N_2344,In_1075,In_2481);
nand U2345 (N_2345,In_1538,In_1402);
or U2346 (N_2346,In_493,In_355);
nand U2347 (N_2347,In_382,In_651);
and U2348 (N_2348,In_1351,In_30);
nand U2349 (N_2349,In_2134,In_365);
nor U2350 (N_2350,In_3,In_305);
nand U2351 (N_2351,In_1576,In_508);
xor U2352 (N_2352,In_2398,In_1920);
nor U2353 (N_2353,In_783,In_2181);
nand U2354 (N_2354,In_1073,In_1901);
xnor U2355 (N_2355,In_1963,In_1940);
and U2356 (N_2356,In_1240,In_1383);
and U2357 (N_2357,In_1102,In_2467);
xor U2358 (N_2358,In_93,In_313);
xor U2359 (N_2359,In_2385,In_1371);
or U2360 (N_2360,In_1156,In_2460);
and U2361 (N_2361,In_2356,In_1331);
or U2362 (N_2362,In_1915,In_54);
or U2363 (N_2363,In_956,In_411);
or U2364 (N_2364,In_134,In_110);
nand U2365 (N_2365,In_206,In_2351);
nor U2366 (N_2366,In_1200,In_867);
nor U2367 (N_2367,In_2284,In_2019);
nor U2368 (N_2368,In_2448,In_477);
and U2369 (N_2369,In_1033,In_44);
xnor U2370 (N_2370,In_1400,In_1940);
nand U2371 (N_2371,In_2107,In_1519);
or U2372 (N_2372,In_2315,In_288);
nand U2373 (N_2373,In_1052,In_1030);
nand U2374 (N_2374,In_2174,In_1378);
xor U2375 (N_2375,In_1771,In_1982);
nor U2376 (N_2376,In_2207,In_782);
nand U2377 (N_2377,In_1060,In_721);
nor U2378 (N_2378,In_1318,In_516);
and U2379 (N_2379,In_1054,In_646);
nor U2380 (N_2380,In_1861,In_1112);
nand U2381 (N_2381,In_560,In_1805);
nand U2382 (N_2382,In_2252,In_1361);
xnor U2383 (N_2383,In_224,In_694);
or U2384 (N_2384,In_2285,In_2498);
and U2385 (N_2385,In_1340,In_1469);
xnor U2386 (N_2386,In_1055,In_2137);
nand U2387 (N_2387,In_1749,In_526);
nand U2388 (N_2388,In_1919,In_1437);
and U2389 (N_2389,In_1531,In_774);
and U2390 (N_2390,In_2358,In_1956);
nand U2391 (N_2391,In_1049,In_2022);
nor U2392 (N_2392,In_1251,In_843);
nor U2393 (N_2393,In_2230,In_1382);
nand U2394 (N_2394,In_317,In_511);
and U2395 (N_2395,In_2067,In_572);
and U2396 (N_2396,In_1252,In_362);
and U2397 (N_2397,In_1969,In_1190);
nor U2398 (N_2398,In_2438,In_2216);
nor U2399 (N_2399,In_1416,In_1689);
nor U2400 (N_2400,In_2277,In_1327);
or U2401 (N_2401,In_46,In_772);
and U2402 (N_2402,In_1836,In_319);
nand U2403 (N_2403,In_279,In_771);
nand U2404 (N_2404,In_209,In_169);
or U2405 (N_2405,In_1711,In_2368);
or U2406 (N_2406,In_2092,In_550);
or U2407 (N_2407,In_1527,In_1997);
and U2408 (N_2408,In_1871,In_234);
nand U2409 (N_2409,In_1947,In_242);
and U2410 (N_2410,In_115,In_896);
nand U2411 (N_2411,In_2027,In_1765);
nand U2412 (N_2412,In_310,In_2295);
nand U2413 (N_2413,In_2260,In_1817);
xnor U2414 (N_2414,In_1725,In_2340);
nor U2415 (N_2415,In_822,In_2141);
and U2416 (N_2416,In_1697,In_2405);
nand U2417 (N_2417,In_792,In_1579);
nand U2418 (N_2418,In_1327,In_1445);
nand U2419 (N_2419,In_2085,In_373);
xor U2420 (N_2420,In_804,In_1335);
or U2421 (N_2421,In_929,In_761);
xor U2422 (N_2422,In_516,In_1171);
nand U2423 (N_2423,In_116,In_407);
nand U2424 (N_2424,In_792,In_311);
or U2425 (N_2425,In_637,In_502);
and U2426 (N_2426,In_1674,In_1144);
nor U2427 (N_2427,In_844,In_631);
nor U2428 (N_2428,In_101,In_2297);
nor U2429 (N_2429,In_837,In_1670);
xnor U2430 (N_2430,In_657,In_973);
nor U2431 (N_2431,In_1464,In_1316);
nand U2432 (N_2432,In_671,In_1477);
and U2433 (N_2433,In_2292,In_1184);
nand U2434 (N_2434,In_271,In_2388);
xor U2435 (N_2435,In_1686,In_2422);
xor U2436 (N_2436,In_1903,In_1);
nand U2437 (N_2437,In_1952,In_903);
nand U2438 (N_2438,In_475,In_1132);
and U2439 (N_2439,In_920,In_940);
xnor U2440 (N_2440,In_224,In_2402);
and U2441 (N_2441,In_928,In_1958);
xnor U2442 (N_2442,In_1237,In_1451);
xor U2443 (N_2443,In_2189,In_367);
and U2444 (N_2444,In_2476,In_1651);
or U2445 (N_2445,In_962,In_468);
and U2446 (N_2446,In_425,In_1214);
xnor U2447 (N_2447,In_1808,In_580);
xnor U2448 (N_2448,In_1901,In_1077);
xnor U2449 (N_2449,In_2250,In_1451);
nor U2450 (N_2450,In_763,In_419);
nand U2451 (N_2451,In_900,In_613);
and U2452 (N_2452,In_2443,In_2226);
nor U2453 (N_2453,In_1355,In_121);
nand U2454 (N_2454,In_1773,In_233);
nor U2455 (N_2455,In_218,In_692);
or U2456 (N_2456,In_877,In_292);
nand U2457 (N_2457,In_93,In_1607);
and U2458 (N_2458,In_1119,In_409);
nor U2459 (N_2459,In_381,In_1667);
nand U2460 (N_2460,In_2298,In_818);
or U2461 (N_2461,In_922,In_208);
nor U2462 (N_2462,In_1948,In_731);
nor U2463 (N_2463,In_1457,In_186);
xor U2464 (N_2464,In_1718,In_23);
nor U2465 (N_2465,In_854,In_1626);
and U2466 (N_2466,In_1645,In_322);
xor U2467 (N_2467,In_1399,In_1111);
and U2468 (N_2468,In_2412,In_1997);
and U2469 (N_2469,In_785,In_2494);
xor U2470 (N_2470,In_1041,In_1596);
or U2471 (N_2471,In_179,In_256);
or U2472 (N_2472,In_1630,In_1205);
nor U2473 (N_2473,In_167,In_181);
nand U2474 (N_2474,In_589,In_890);
or U2475 (N_2475,In_1859,In_1601);
nor U2476 (N_2476,In_2415,In_1951);
nor U2477 (N_2477,In_1723,In_1171);
nor U2478 (N_2478,In_991,In_1317);
nor U2479 (N_2479,In_2430,In_1315);
or U2480 (N_2480,In_1420,In_1389);
or U2481 (N_2481,In_1474,In_150);
or U2482 (N_2482,In_2192,In_1769);
nor U2483 (N_2483,In_1821,In_2465);
nand U2484 (N_2484,In_2421,In_1951);
nor U2485 (N_2485,In_252,In_2082);
nor U2486 (N_2486,In_2267,In_694);
xor U2487 (N_2487,In_192,In_347);
nor U2488 (N_2488,In_114,In_1354);
nor U2489 (N_2489,In_131,In_316);
nor U2490 (N_2490,In_1202,In_1499);
xor U2491 (N_2491,In_2498,In_193);
xor U2492 (N_2492,In_2227,In_502);
xnor U2493 (N_2493,In_172,In_2275);
nor U2494 (N_2494,In_1816,In_417);
nand U2495 (N_2495,In_1973,In_1238);
nor U2496 (N_2496,In_2259,In_394);
xor U2497 (N_2497,In_749,In_1980);
nand U2498 (N_2498,In_1986,In_734);
and U2499 (N_2499,In_2004,In_2452);
xnor U2500 (N_2500,In_15,In_946);
nor U2501 (N_2501,In_790,In_717);
xnor U2502 (N_2502,In_2060,In_1010);
nor U2503 (N_2503,In_495,In_398);
nand U2504 (N_2504,In_2352,In_1230);
and U2505 (N_2505,In_1298,In_49);
nor U2506 (N_2506,In_642,In_1601);
xor U2507 (N_2507,In_1388,In_630);
and U2508 (N_2508,In_2006,In_954);
nor U2509 (N_2509,In_1033,In_1423);
and U2510 (N_2510,In_1678,In_1613);
nor U2511 (N_2511,In_2290,In_1217);
and U2512 (N_2512,In_519,In_1346);
and U2513 (N_2513,In_2130,In_29);
and U2514 (N_2514,In_1314,In_1682);
xnor U2515 (N_2515,In_1831,In_479);
nand U2516 (N_2516,In_1138,In_2055);
nand U2517 (N_2517,In_2087,In_81);
nor U2518 (N_2518,In_547,In_1343);
nand U2519 (N_2519,In_1488,In_2326);
and U2520 (N_2520,In_2483,In_607);
and U2521 (N_2521,In_1210,In_1458);
and U2522 (N_2522,In_2277,In_2255);
nor U2523 (N_2523,In_605,In_1971);
xor U2524 (N_2524,In_2021,In_1072);
nand U2525 (N_2525,In_435,In_1093);
xor U2526 (N_2526,In_326,In_1055);
and U2527 (N_2527,In_2096,In_448);
and U2528 (N_2528,In_1264,In_2289);
nor U2529 (N_2529,In_1762,In_2296);
and U2530 (N_2530,In_978,In_991);
xnor U2531 (N_2531,In_539,In_1024);
and U2532 (N_2532,In_867,In_327);
nand U2533 (N_2533,In_2094,In_1297);
and U2534 (N_2534,In_1814,In_2452);
and U2535 (N_2535,In_528,In_179);
or U2536 (N_2536,In_1416,In_489);
nand U2537 (N_2537,In_2147,In_554);
xor U2538 (N_2538,In_535,In_800);
and U2539 (N_2539,In_1815,In_1258);
and U2540 (N_2540,In_1898,In_2447);
nor U2541 (N_2541,In_1936,In_894);
nor U2542 (N_2542,In_602,In_1526);
nor U2543 (N_2543,In_1343,In_1666);
and U2544 (N_2544,In_104,In_1798);
nand U2545 (N_2545,In_109,In_118);
nor U2546 (N_2546,In_643,In_85);
nand U2547 (N_2547,In_1963,In_1034);
and U2548 (N_2548,In_1862,In_2092);
xnor U2549 (N_2549,In_1811,In_719);
or U2550 (N_2550,In_2495,In_445);
and U2551 (N_2551,In_2211,In_86);
nand U2552 (N_2552,In_2172,In_497);
nand U2553 (N_2553,In_274,In_242);
nor U2554 (N_2554,In_734,In_311);
or U2555 (N_2555,In_1767,In_2014);
nor U2556 (N_2556,In_183,In_798);
xor U2557 (N_2557,In_1909,In_2041);
nor U2558 (N_2558,In_1576,In_673);
nor U2559 (N_2559,In_1480,In_900);
nand U2560 (N_2560,In_1498,In_84);
nor U2561 (N_2561,In_914,In_1130);
and U2562 (N_2562,In_1092,In_2082);
xnor U2563 (N_2563,In_2232,In_63);
xnor U2564 (N_2564,In_1534,In_948);
nand U2565 (N_2565,In_1832,In_1441);
and U2566 (N_2566,In_1548,In_2204);
and U2567 (N_2567,In_2174,In_2160);
and U2568 (N_2568,In_601,In_1979);
xnor U2569 (N_2569,In_1388,In_1118);
nand U2570 (N_2570,In_1308,In_725);
and U2571 (N_2571,In_1934,In_814);
or U2572 (N_2572,In_1185,In_2143);
nand U2573 (N_2573,In_1484,In_669);
nand U2574 (N_2574,In_255,In_2456);
xnor U2575 (N_2575,In_944,In_1009);
nor U2576 (N_2576,In_962,In_730);
and U2577 (N_2577,In_1467,In_1510);
nor U2578 (N_2578,In_2193,In_768);
nor U2579 (N_2579,In_2258,In_933);
nor U2580 (N_2580,In_1775,In_1713);
or U2581 (N_2581,In_419,In_1025);
nor U2582 (N_2582,In_1118,In_1068);
nor U2583 (N_2583,In_1894,In_329);
or U2584 (N_2584,In_446,In_931);
or U2585 (N_2585,In_1783,In_244);
nor U2586 (N_2586,In_1373,In_173);
and U2587 (N_2587,In_280,In_1357);
or U2588 (N_2588,In_2093,In_1443);
nor U2589 (N_2589,In_394,In_1271);
xor U2590 (N_2590,In_802,In_693);
and U2591 (N_2591,In_135,In_406);
and U2592 (N_2592,In_2305,In_1272);
or U2593 (N_2593,In_1593,In_1301);
and U2594 (N_2594,In_2206,In_1328);
nand U2595 (N_2595,In_109,In_1750);
or U2596 (N_2596,In_656,In_1326);
and U2597 (N_2597,In_1449,In_2094);
nand U2598 (N_2598,In_1073,In_1898);
and U2599 (N_2599,In_1440,In_509);
xor U2600 (N_2600,In_1878,In_2348);
or U2601 (N_2601,In_1372,In_1848);
nand U2602 (N_2602,In_63,In_1810);
or U2603 (N_2603,In_364,In_948);
xnor U2604 (N_2604,In_1810,In_325);
nand U2605 (N_2605,In_383,In_69);
or U2606 (N_2606,In_879,In_1480);
nor U2607 (N_2607,In_2239,In_2178);
or U2608 (N_2608,In_1777,In_1342);
and U2609 (N_2609,In_190,In_205);
or U2610 (N_2610,In_2096,In_1951);
or U2611 (N_2611,In_1078,In_727);
nand U2612 (N_2612,In_1561,In_1330);
nand U2613 (N_2613,In_2463,In_1025);
and U2614 (N_2614,In_1033,In_179);
nor U2615 (N_2615,In_1059,In_1760);
and U2616 (N_2616,In_585,In_1009);
and U2617 (N_2617,In_2426,In_1474);
and U2618 (N_2618,In_886,In_1248);
and U2619 (N_2619,In_291,In_428);
nand U2620 (N_2620,In_1358,In_1830);
xor U2621 (N_2621,In_2495,In_2478);
nand U2622 (N_2622,In_1008,In_1129);
xor U2623 (N_2623,In_249,In_1461);
xnor U2624 (N_2624,In_552,In_1350);
xor U2625 (N_2625,In_1129,In_2268);
nand U2626 (N_2626,In_831,In_2305);
and U2627 (N_2627,In_2496,In_1378);
xnor U2628 (N_2628,In_854,In_58);
xnor U2629 (N_2629,In_2334,In_1474);
and U2630 (N_2630,In_2290,In_1150);
xor U2631 (N_2631,In_2289,In_824);
or U2632 (N_2632,In_77,In_2336);
nor U2633 (N_2633,In_501,In_1722);
nand U2634 (N_2634,In_1222,In_1351);
and U2635 (N_2635,In_43,In_2371);
xnor U2636 (N_2636,In_25,In_661);
nor U2637 (N_2637,In_1418,In_320);
and U2638 (N_2638,In_1988,In_885);
or U2639 (N_2639,In_2345,In_1462);
and U2640 (N_2640,In_2310,In_275);
nand U2641 (N_2641,In_1295,In_1071);
nor U2642 (N_2642,In_1029,In_2000);
and U2643 (N_2643,In_1702,In_1847);
xnor U2644 (N_2644,In_1304,In_1266);
or U2645 (N_2645,In_968,In_914);
and U2646 (N_2646,In_301,In_2043);
xor U2647 (N_2647,In_2329,In_1551);
xor U2648 (N_2648,In_1403,In_1068);
and U2649 (N_2649,In_1239,In_904);
or U2650 (N_2650,In_958,In_1535);
nor U2651 (N_2651,In_2252,In_2045);
xnor U2652 (N_2652,In_784,In_84);
nand U2653 (N_2653,In_362,In_705);
and U2654 (N_2654,In_794,In_131);
nor U2655 (N_2655,In_1559,In_667);
and U2656 (N_2656,In_2356,In_849);
xor U2657 (N_2657,In_2183,In_884);
nor U2658 (N_2658,In_2223,In_2218);
nand U2659 (N_2659,In_614,In_2019);
nand U2660 (N_2660,In_108,In_2201);
and U2661 (N_2661,In_1706,In_2383);
nand U2662 (N_2662,In_1081,In_1118);
or U2663 (N_2663,In_634,In_2107);
and U2664 (N_2664,In_1500,In_259);
nor U2665 (N_2665,In_2268,In_1139);
xor U2666 (N_2666,In_955,In_2143);
and U2667 (N_2667,In_665,In_818);
or U2668 (N_2668,In_894,In_1366);
xor U2669 (N_2669,In_478,In_2241);
or U2670 (N_2670,In_257,In_738);
nand U2671 (N_2671,In_623,In_1828);
nand U2672 (N_2672,In_1438,In_2469);
or U2673 (N_2673,In_1531,In_1977);
xor U2674 (N_2674,In_467,In_199);
and U2675 (N_2675,In_1417,In_1900);
or U2676 (N_2676,In_1354,In_1205);
xnor U2677 (N_2677,In_287,In_1464);
xnor U2678 (N_2678,In_481,In_541);
or U2679 (N_2679,In_379,In_1877);
and U2680 (N_2680,In_421,In_488);
nor U2681 (N_2681,In_644,In_552);
nor U2682 (N_2682,In_1291,In_1278);
and U2683 (N_2683,In_88,In_2361);
or U2684 (N_2684,In_1694,In_998);
or U2685 (N_2685,In_305,In_1641);
and U2686 (N_2686,In_221,In_467);
xor U2687 (N_2687,In_1854,In_707);
or U2688 (N_2688,In_1216,In_1246);
and U2689 (N_2689,In_1517,In_1893);
nand U2690 (N_2690,In_499,In_985);
nor U2691 (N_2691,In_1903,In_1637);
and U2692 (N_2692,In_2340,In_490);
nand U2693 (N_2693,In_2295,In_1753);
xnor U2694 (N_2694,In_1925,In_265);
and U2695 (N_2695,In_577,In_2200);
and U2696 (N_2696,In_1870,In_211);
and U2697 (N_2697,In_1780,In_2324);
nand U2698 (N_2698,In_1822,In_1468);
and U2699 (N_2699,In_1844,In_380);
nor U2700 (N_2700,In_137,In_925);
nor U2701 (N_2701,In_2032,In_32);
or U2702 (N_2702,In_1569,In_1427);
or U2703 (N_2703,In_283,In_413);
xor U2704 (N_2704,In_339,In_1713);
and U2705 (N_2705,In_2083,In_1708);
xor U2706 (N_2706,In_559,In_1563);
and U2707 (N_2707,In_745,In_1604);
or U2708 (N_2708,In_1248,In_1351);
nor U2709 (N_2709,In_2012,In_1999);
and U2710 (N_2710,In_32,In_912);
nor U2711 (N_2711,In_2420,In_76);
and U2712 (N_2712,In_2143,In_1609);
nor U2713 (N_2713,In_2097,In_466);
or U2714 (N_2714,In_1501,In_1227);
or U2715 (N_2715,In_1152,In_2274);
and U2716 (N_2716,In_1558,In_957);
xnor U2717 (N_2717,In_2324,In_1568);
and U2718 (N_2718,In_2436,In_1755);
or U2719 (N_2719,In_1104,In_776);
and U2720 (N_2720,In_1552,In_41);
or U2721 (N_2721,In_367,In_1265);
and U2722 (N_2722,In_1326,In_55);
nand U2723 (N_2723,In_1221,In_167);
and U2724 (N_2724,In_1199,In_1942);
and U2725 (N_2725,In_985,In_163);
and U2726 (N_2726,In_1024,In_1764);
nor U2727 (N_2727,In_1897,In_1277);
nand U2728 (N_2728,In_1114,In_55);
nor U2729 (N_2729,In_347,In_2475);
xor U2730 (N_2730,In_1487,In_1284);
nand U2731 (N_2731,In_1511,In_1456);
and U2732 (N_2732,In_1604,In_2067);
xnor U2733 (N_2733,In_786,In_1772);
xor U2734 (N_2734,In_787,In_1941);
and U2735 (N_2735,In_848,In_739);
and U2736 (N_2736,In_1345,In_1324);
nor U2737 (N_2737,In_656,In_1039);
nor U2738 (N_2738,In_2453,In_784);
nor U2739 (N_2739,In_1321,In_2133);
and U2740 (N_2740,In_921,In_196);
and U2741 (N_2741,In_2224,In_1667);
nor U2742 (N_2742,In_1423,In_1536);
nand U2743 (N_2743,In_1703,In_1445);
nand U2744 (N_2744,In_1831,In_2288);
xnor U2745 (N_2745,In_877,In_40);
or U2746 (N_2746,In_1953,In_2316);
nor U2747 (N_2747,In_2251,In_1566);
nand U2748 (N_2748,In_1605,In_2151);
nand U2749 (N_2749,In_2226,In_305);
xor U2750 (N_2750,In_2391,In_783);
and U2751 (N_2751,In_173,In_866);
xor U2752 (N_2752,In_1984,In_648);
xnor U2753 (N_2753,In_2163,In_1329);
and U2754 (N_2754,In_1809,In_1720);
xnor U2755 (N_2755,In_2118,In_2343);
and U2756 (N_2756,In_398,In_833);
nand U2757 (N_2757,In_2376,In_1671);
and U2758 (N_2758,In_2376,In_1827);
nor U2759 (N_2759,In_2490,In_1109);
nand U2760 (N_2760,In_322,In_1723);
or U2761 (N_2761,In_2306,In_2313);
or U2762 (N_2762,In_579,In_2141);
and U2763 (N_2763,In_2284,In_1890);
or U2764 (N_2764,In_1508,In_35);
or U2765 (N_2765,In_912,In_1238);
or U2766 (N_2766,In_1817,In_2417);
and U2767 (N_2767,In_432,In_1734);
nand U2768 (N_2768,In_0,In_1053);
or U2769 (N_2769,In_2331,In_762);
xnor U2770 (N_2770,In_2390,In_168);
xnor U2771 (N_2771,In_295,In_1471);
or U2772 (N_2772,In_1677,In_945);
nand U2773 (N_2773,In_513,In_223);
nor U2774 (N_2774,In_113,In_2048);
nor U2775 (N_2775,In_2156,In_471);
and U2776 (N_2776,In_1839,In_712);
and U2777 (N_2777,In_253,In_279);
nor U2778 (N_2778,In_600,In_297);
and U2779 (N_2779,In_2022,In_1341);
and U2780 (N_2780,In_2307,In_1545);
xor U2781 (N_2781,In_1446,In_2098);
nor U2782 (N_2782,In_1977,In_209);
nand U2783 (N_2783,In_1121,In_1722);
nand U2784 (N_2784,In_732,In_1757);
nor U2785 (N_2785,In_2332,In_1330);
nor U2786 (N_2786,In_2115,In_742);
or U2787 (N_2787,In_2008,In_1115);
nor U2788 (N_2788,In_1184,In_1488);
and U2789 (N_2789,In_1563,In_1702);
and U2790 (N_2790,In_241,In_449);
nor U2791 (N_2791,In_1021,In_353);
or U2792 (N_2792,In_2346,In_2480);
nand U2793 (N_2793,In_1674,In_42);
or U2794 (N_2794,In_1961,In_694);
nor U2795 (N_2795,In_28,In_1582);
and U2796 (N_2796,In_278,In_1234);
or U2797 (N_2797,In_1086,In_929);
nand U2798 (N_2798,In_330,In_1256);
xor U2799 (N_2799,In_229,In_209);
nand U2800 (N_2800,In_510,In_372);
xnor U2801 (N_2801,In_1913,In_2475);
xor U2802 (N_2802,In_858,In_9);
or U2803 (N_2803,In_93,In_307);
xnor U2804 (N_2804,In_435,In_42);
or U2805 (N_2805,In_545,In_62);
xnor U2806 (N_2806,In_140,In_1156);
nor U2807 (N_2807,In_866,In_308);
or U2808 (N_2808,In_1407,In_2492);
nor U2809 (N_2809,In_1668,In_1710);
nor U2810 (N_2810,In_1419,In_1059);
xnor U2811 (N_2811,In_18,In_393);
and U2812 (N_2812,In_97,In_1649);
nor U2813 (N_2813,In_1267,In_2203);
or U2814 (N_2814,In_1300,In_790);
or U2815 (N_2815,In_463,In_1009);
nand U2816 (N_2816,In_803,In_357);
and U2817 (N_2817,In_2230,In_549);
or U2818 (N_2818,In_2427,In_2104);
and U2819 (N_2819,In_361,In_281);
nand U2820 (N_2820,In_1591,In_33);
nor U2821 (N_2821,In_1216,In_54);
and U2822 (N_2822,In_1285,In_2154);
xor U2823 (N_2823,In_1800,In_814);
nor U2824 (N_2824,In_1362,In_459);
xnor U2825 (N_2825,In_508,In_349);
nor U2826 (N_2826,In_2146,In_1366);
xnor U2827 (N_2827,In_2026,In_1469);
and U2828 (N_2828,In_2348,In_1849);
nand U2829 (N_2829,In_1989,In_1104);
nand U2830 (N_2830,In_1546,In_86);
and U2831 (N_2831,In_1469,In_1121);
nand U2832 (N_2832,In_2315,In_1044);
xor U2833 (N_2833,In_2040,In_1454);
nor U2834 (N_2834,In_2243,In_203);
and U2835 (N_2835,In_826,In_548);
nand U2836 (N_2836,In_1344,In_1216);
nor U2837 (N_2837,In_778,In_745);
and U2838 (N_2838,In_252,In_57);
nand U2839 (N_2839,In_1657,In_1313);
nor U2840 (N_2840,In_262,In_2082);
or U2841 (N_2841,In_1641,In_565);
nand U2842 (N_2842,In_1790,In_1138);
nor U2843 (N_2843,In_2076,In_2059);
and U2844 (N_2844,In_1445,In_417);
and U2845 (N_2845,In_527,In_824);
xor U2846 (N_2846,In_1996,In_217);
nor U2847 (N_2847,In_1575,In_2436);
or U2848 (N_2848,In_2204,In_2360);
xnor U2849 (N_2849,In_2068,In_1471);
and U2850 (N_2850,In_1771,In_749);
nor U2851 (N_2851,In_2451,In_718);
nor U2852 (N_2852,In_517,In_1296);
nand U2853 (N_2853,In_386,In_208);
nand U2854 (N_2854,In_1651,In_748);
xnor U2855 (N_2855,In_306,In_1394);
nor U2856 (N_2856,In_753,In_2306);
xor U2857 (N_2857,In_1710,In_1442);
or U2858 (N_2858,In_1057,In_2151);
and U2859 (N_2859,In_1525,In_76);
nand U2860 (N_2860,In_1256,In_1433);
nand U2861 (N_2861,In_1146,In_906);
or U2862 (N_2862,In_2237,In_708);
nor U2863 (N_2863,In_1833,In_2496);
or U2864 (N_2864,In_1680,In_1751);
and U2865 (N_2865,In_2149,In_180);
nor U2866 (N_2866,In_1788,In_1065);
xor U2867 (N_2867,In_1879,In_124);
nor U2868 (N_2868,In_355,In_1613);
xnor U2869 (N_2869,In_828,In_1192);
or U2870 (N_2870,In_1397,In_985);
nor U2871 (N_2871,In_1891,In_208);
nand U2872 (N_2872,In_1897,In_1630);
nor U2873 (N_2873,In_298,In_1910);
nand U2874 (N_2874,In_1438,In_2131);
or U2875 (N_2875,In_328,In_1593);
xor U2876 (N_2876,In_1511,In_1240);
and U2877 (N_2877,In_218,In_232);
or U2878 (N_2878,In_289,In_1859);
nor U2879 (N_2879,In_1290,In_174);
xor U2880 (N_2880,In_29,In_1652);
nand U2881 (N_2881,In_941,In_354);
nand U2882 (N_2882,In_2241,In_162);
xor U2883 (N_2883,In_2423,In_1257);
and U2884 (N_2884,In_1898,In_558);
or U2885 (N_2885,In_1545,In_1559);
xnor U2886 (N_2886,In_1514,In_1478);
xnor U2887 (N_2887,In_528,In_1437);
nor U2888 (N_2888,In_1587,In_2225);
or U2889 (N_2889,In_1776,In_292);
and U2890 (N_2890,In_890,In_1084);
and U2891 (N_2891,In_2213,In_226);
xnor U2892 (N_2892,In_669,In_2278);
xnor U2893 (N_2893,In_2471,In_1948);
and U2894 (N_2894,In_1519,In_203);
nand U2895 (N_2895,In_1527,In_379);
nand U2896 (N_2896,In_32,In_2369);
or U2897 (N_2897,In_1123,In_1366);
nor U2898 (N_2898,In_1745,In_2377);
nand U2899 (N_2899,In_1464,In_1492);
nand U2900 (N_2900,In_1042,In_111);
and U2901 (N_2901,In_557,In_1305);
nor U2902 (N_2902,In_2469,In_2209);
nand U2903 (N_2903,In_1501,In_1780);
or U2904 (N_2904,In_562,In_2388);
xor U2905 (N_2905,In_603,In_2299);
nand U2906 (N_2906,In_1340,In_1804);
or U2907 (N_2907,In_1281,In_1241);
or U2908 (N_2908,In_2051,In_384);
nor U2909 (N_2909,In_1682,In_2125);
or U2910 (N_2910,In_2014,In_1193);
or U2911 (N_2911,In_948,In_2442);
or U2912 (N_2912,In_1333,In_253);
and U2913 (N_2913,In_1843,In_240);
nor U2914 (N_2914,In_1512,In_2150);
nand U2915 (N_2915,In_2134,In_1011);
nor U2916 (N_2916,In_2101,In_1645);
and U2917 (N_2917,In_2449,In_249);
nor U2918 (N_2918,In_524,In_781);
and U2919 (N_2919,In_723,In_483);
nand U2920 (N_2920,In_2413,In_969);
nand U2921 (N_2921,In_1016,In_2440);
nor U2922 (N_2922,In_1119,In_1223);
nand U2923 (N_2923,In_2039,In_1548);
nand U2924 (N_2924,In_1411,In_547);
nand U2925 (N_2925,In_1115,In_2421);
nor U2926 (N_2926,In_1443,In_381);
xnor U2927 (N_2927,In_992,In_517);
and U2928 (N_2928,In_2085,In_1981);
xor U2929 (N_2929,In_1671,In_250);
xor U2930 (N_2930,In_1241,In_1909);
xor U2931 (N_2931,In_336,In_1821);
nor U2932 (N_2932,In_751,In_618);
or U2933 (N_2933,In_678,In_2066);
and U2934 (N_2934,In_1747,In_2087);
or U2935 (N_2935,In_1865,In_1323);
xnor U2936 (N_2936,In_110,In_430);
nor U2937 (N_2937,In_791,In_1191);
xor U2938 (N_2938,In_1350,In_2445);
and U2939 (N_2939,In_2270,In_177);
nand U2940 (N_2940,In_767,In_1503);
xnor U2941 (N_2941,In_2170,In_744);
and U2942 (N_2942,In_193,In_931);
xnor U2943 (N_2943,In_1319,In_1565);
xor U2944 (N_2944,In_2084,In_1553);
xor U2945 (N_2945,In_1010,In_533);
or U2946 (N_2946,In_1686,In_753);
xor U2947 (N_2947,In_1718,In_2310);
nand U2948 (N_2948,In_1214,In_1946);
xnor U2949 (N_2949,In_1889,In_906);
or U2950 (N_2950,In_89,In_932);
and U2951 (N_2951,In_1917,In_1309);
or U2952 (N_2952,In_2200,In_90);
xor U2953 (N_2953,In_2131,In_1528);
and U2954 (N_2954,In_653,In_295);
and U2955 (N_2955,In_1786,In_65);
or U2956 (N_2956,In_1090,In_2162);
or U2957 (N_2957,In_653,In_1287);
nand U2958 (N_2958,In_223,In_1035);
nand U2959 (N_2959,In_305,In_550);
and U2960 (N_2960,In_1325,In_1985);
nor U2961 (N_2961,In_1710,In_291);
nor U2962 (N_2962,In_1269,In_2041);
or U2963 (N_2963,In_1861,In_2421);
nor U2964 (N_2964,In_2373,In_361);
xor U2965 (N_2965,In_950,In_1577);
nand U2966 (N_2966,In_101,In_1178);
and U2967 (N_2967,In_1884,In_1206);
or U2968 (N_2968,In_2351,In_1847);
nand U2969 (N_2969,In_712,In_1740);
nor U2970 (N_2970,In_2255,In_616);
or U2971 (N_2971,In_1233,In_262);
and U2972 (N_2972,In_2057,In_1727);
and U2973 (N_2973,In_350,In_136);
or U2974 (N_2974,In_160,In_763);
nand U2975 (N_2975,In_916,In_475);
or U2976 (N_2976,In_146,In_2052);
or U2977 (N_2977,In_2410,In_2480);
xor U2978 (N_2978,In_1643,In_808);
nor U2979 (N_2979,In_263,In_816);
or U2980 (N_2980,In_465,In_383);
or U2981 (N_2981,In_1834,In_966);
and U2982 (N_2982,In_766,In_633);
nor U2983 (N_2983,In_1061,In_179);
nor U2984 (N_2984,In_612,In_1035);
and U2985 (N_2985,In_1146,In_1151);
nand U2986 (N_2986,In_872,In_2080);
xnor U2987 (N_2987,In_251,In_1274);
nor U2988 (N_2988,In_1349,In_1979);
nand U2989 (N_2989,In_1693,In_412);
xor U2990 (N_2990,In_526,In_1700);
xnor U2991 (N_2991,In_2112,In_1352);
nand U2992 (N_2992,In_427,In_1866);
nor U2993 (N_2993,In_1997,In_106);
nor U2994 (N_2994,In_219,In_989);
nor U2995 (N_2995,In_1644,In_1918);
nand U2996 (N_2996,In_1789,In_695);
and U2997 (N_2997,In_1226,In_2434);
nand U2998 (N_2998,In_2002,In_1729);
nand U2999 (N_2999,In_267,In_1492);
xor U3000 (N_3000,In_115,In_2218);
nor U3001 (N_3001,In_1059,In_2497);
xor U3002 (N_3002,In_470,In_1475);
nand U3003 (N_3003,In_1434,In_1370);
xor U3004 (N_3004,In_1519,In_1742);
xor U3005 (N_3005,In_972,In_78);
xnor U3006 (N_3006,In_936,In_2249);
and U3007 (N_3007,In_756,In_1605);
nor U3008 (N_3008,In_1697,In_845);
and U3009 (N_3009,In_2464,In_1748);
and U3010 (N_3010,In_2315,In_2147);
and U3011 (N_3011,In_503,In_1024);
or U3012 (N_3012,In_893,In_2062);
nor U3013 (N_3013,In_963,In_1986);
or U3014 (N_3014,In_1011,In_906);
xor U3015 (N_3015,In_829,In_2125);
nand U3016 (N_3016,In_2170,In_602);
or U3017 (N_3017,In_2208,In_181);
and U3018 (N_3018,In_2256,In_122);
and U3019 (N_3019,In_1966,In_1874);
nor U3020 (N_3020,In_1326,In_289);
or U3021 (N_3021,In_382,In_2174);
nand U3022 (N_3022,In_634,In_1269);
or U3023 (N_3023,In_1405,In_859);
and U3024 (N_3024,In_1913,In_1843);
or U3025 (N_3025,In_1208,In_8);
nor U3026 (N_3026,In_2376,In_41);
xor U3027 (N_3027,In_99,In_44);
nor U3028 (N_3028,In_1539,In_2377);
nor U3029 (N_3029,In_336,In_127);
and U3030 (N_3030,In_518,In_438);
xnor U3031 (N_3031,In_2240,In_849);
xor U3032 (N_3032,In_718,In_887);
or U3033 (N_3033,In_1131,In_2393);
xor U3034 (N_3034,In_1330,In_65);
and U3035 (N_3035,In_307,In_860);
and U3036 (N_3036,In_1995,In_762);
nand U3037 (N_3037,In_105,In_1927);
xnor U3038 (N_3038,In_2279,In_2200);
and U3039 (N_3039,In_1902,In_2120);
nor U3040 (N_3040,In_764,In_1296);
or U3041 (N_3041,In_1552,In_352);
and U3042 (N_3042,In_1653,In_1843);
and U3043 (N_3043,In_187,In_1007);
xor U3044 (N_3044,In_1507,In_1739);
and U3045 (N_3045,In_317,In_786);
nand U3046 (N_3046,In_1423,In_2476);
or U3047 (N_3047,In_773,In_1917);
nand U3048 (N_3048,In_1263,In_2082);
xor U3049 (N_3049,In_442,In_423);
and U3050 (N_3050,In_1688,In_1618);
nor U3051 (N_3051,In_941,In_1199);
xor U3052 (N_3052,In_233,In_1734);
or U3053 (N_3053,In_1773,In_1532);
nor U3054 (N_3054,In_279,In_1076);
nor U3055 (N_3055,In_1609,In_1979);
and U3056 (N_3056,In_1753,In_824);
nand U3057 (N_3057,In_1665,In_1599);
xor U3058 (N_3058,In_859,In_1707);
nor U3059 (N_3059,In_1986,In_495);
xnor U3060 (N_3060,In_1639,In_2054);
nand U3061 (N_3061,In_659,In_1174);
and U3062 (N_3062,In_2261,In_142);
xor U3063 (N_3063,In_663,In_1652);
nor U3064 (N_3064,In_2073,In_1225);
xor U3065 (N_3065,In_2366,In_623);
or U3066 (N_3066,In_928,In_1072);
nor U3067 (N_3067,In_68,In_1448);
xnor U3068 (N_3068,In_202,In_1295);
nand U3069 (N_3069,In_176,In_180);
and U3070 (N_3070,In_168,In_1495);
nand U3071 (N_3071,In_1981,In_975);
xnor U3072 (N_3072,In_947,In_913);
nor U3073 (N_3073,In_271,In_1327);
xnor U3074 (N_3074,In_1980,In_2160);
and U3075 (N_3075,In_275,In_284);
or U3076 (N_3076,In_1920,In_36);
and U3077 (N_3077,In_922,In_1737);
xor U3078 (N_3078,In_265,In_26);
or U3079 (N_3079,In_724,In_323);
nor U3080 (N_3080,In_2334,In_839);
or U3081 (N_3081,In_1811,In_1283);
xor U3082 (N_3082,In_2453,In_1225);
nor U3083 (N_3083,In_70,In_400);
nand U3084 (N_3084,In_289,In_1033);
and U3085 (N_3085,In_980,In_2323);
or U3086 (N_3086,In_1344,In_1927);
and U3087 (N_3087,In_1101,In_515);
or U3088 (N_3088,In_661,In_2132);
and U3089 (N_3089,In_1333,In_2018);
and U3090 (N_3090,In_1638,In_2369);
or U3091 (N_3091,In_2177,In_1250);
and U3092 (N_3092,In_42,In_1998);
and U3093 (N_3093,In_403,In_225);
or U3094 (N_3094,In_1263,In_100);
nor U3095 (N_3095,In_115,In_641);
nand U3096 (N_3096,In_1892,In_252);
nand U3097 (N_3097,In_1482,In_417);
and U3098 (N_3098,In_1539,In_1551);
nand U3099 (N_3099,In_1278,In_1427);
xnor U3100 (N_3100,In_1715,In_1701);
nand U3101 (N_3101,In_2373,In_1812);
and U3102 (N_3102,In_899,In_1874);
nor U3103 (N_3103,In_1807,In_1642);
and U3104 (N_3104,In_300,In_990);
and U3105 (N_3105,In_1290,In_906);
nor U3106 (N_3106,In_914,In_25);
xor U3107 (N_3107,In_2152,In_978);
or U3108 (N_3108,In_1355,In_22);
nand U3109 (N_3109,In_820,In_2047);
xnor U3110 (N_3110,In_2237,In_924);
or U3111 (N_3111,In_1249,In_2228);
nand U3112 (N_3112,In_342,In_220);
or U3113 (N_3113,In_1552,In_1885);
nor U3114 (N_3114,In_1846,In_2463);
or U3115 (N_3115,In_2182,In_1384);
nor U3116 (N_3116,In_1152,In_2460);
nor U3117 (N_3117,In_1999,In_1555);
xnor U3118 (N_3118,In_1396,In_1355);
and U3119 (N_3119,In_735,In_272);
nor U3120 (N_3120,In_2051,In_1195);
nand U3121 (N_3121,In_813,In_318);
and U3122 (N_3122,In_2472,In_1836);
nor U3123 (N_3123,In_425,In_899);
nand U3124 (N_3124,In_2307,In_1164);
or U3125 (N_3125,N_515,N_1420);
nand U3126 (N_3126,N_1213,N_872);
and U3127 (N_3127,N_3027,N_1330);
xnor U3128 (N_3128,N_558,N_2917);
nor U3129 (N_3129,N_1345,N_2958);
xnor U3130 (N_3130,N_2526,N_917);
xor U3131 (N_3131,N_1349,N_103);
xor U3132 (N_3132,N_822,N_812);
or U3133 (N_3133,N_2372,N_2508);
and U3134 (N_3134,N_2159,N_2876);
and U3135 (N_3135,N_2607,N_2498);
or U3136 (N_3136,N_221,N_1685);
xor U3137 (N_3137,N_1613,N_147);
and U3138 (N_3138,N_2129,N_2535);
or U3139 (N_3139,N_215,N_1909);
or U3140 (N_3140,N_849,N_119);
nor U3141 (N_3141,N_413,N_2707);
nand U3142 (N_3142,N_1552,N_2527);
nor U3143 (N_3143,N_288,N_130);
nand U3144 (N_3144,N_1939,N_611);
nand U3145 (N_3145,N_654,N_1236);
or U3146 (N_3146,N_132,N_2888);
or U3147 (N_3147,N_1474,N_2740);
or U3148 (N_3148,N_1350,N_1805);
xor U3149 (N_3149,N_2761,N_428);
nand U3150 (N_3150,N_2257,N_908);
nand U3151 (N_3151,N_225,N_1186);
xnor U3152 (N_3152,N_635,N_2260);
nand U3153 (N_3153,N_861,N_2478);
or U3154 (N_3154,N_844,N_1392);
and U3155 (N_3155,N_1734,N_869);
nand U3156 (N_3156,N_1256,N_757);
and U3157 (N_3157,N_1468,N_2911);
and U3158 (N_3158,N_2020,N_1817);
xor U3159 (N_3159,N_2988,N_1949);
nand U3160 (N_3160,N_456,N_169);
or U3161 (N_3161,N_1629,N_2142);
and U3162 (N_3162,N_67,N_3079);
xnor U3163 (N_3163,N_2060,N_2480);
nor U3164 (N_3164,N_1559,N_213);
or U3165 (N_3165,N_1176,N_2834);
or U3166 (N_3166,N_2269,N_475);
nand U3167 (N_3167,N_1381,N_3054);
xor U3168 (N_3168,N_2727,N_2419);
or U3169 (N_3169,N_1369,N_2791);
and U3170 (N_3170,N_2253,N_749);
xor U3171 (N_3171,N_1780,N_1918);
xnor U3172 (N_3172,N_203,N_426);
or U3173 (N_3173,N_2246,N_887);
nand U3174 (N_3174,N_2795,N_1996);
nor U3175 (N_3175,N_2453,N_2733);
xor U3176 (N_3176,N_1466,N_634);
or U3177 (N_3177,N_1793,N_149);
xor U3178 (N_3178,N_2803,N_264);
xor U3179 (N_3179,N_1305,N_1973);
and U3180 (N_3180,N_2821,N_2776);
nor U3181 (N_3181,N_1153,N_365);
xor U3182 (N_3182,N_2034,N_1658);
nand U3183 (N_3183,N_702,N_695);
nand U3184 (N_3184,N_1818,N_1244);
nand U3185 (N_3185,N_853,N_2642);
and U3186 (N_3186,N_2348,N_404);
nor U3187 (N_3187,N_446,N_1219);
xnor U3188 (N_3188,N_2681,N_1616);
or U3189 (N_3189,N_1344,N_2062);
or U3190 (N_3190,N_1763,N_1985);
nor U3191 (N_3191,N_2657,N_1907);
nand U3192 (N_3192,N_907,N_1239);
nand U3193 (N_3193,N_1592,N_2202);
or U3194 (N_3194,N_1881,N_2183);
or U3195 (N_3195,N_2154,N_470);
or U3196 (N_3196,N_2933,N_370);
nand U3197 (N_3197,N_2583,N_1892);
or U3198 (N_3198,N_246,N_98);
and U3199 (N_3199,N_2742,N_1396);
nand U3200 (N_3200,N_2076,N_2381);
or U3201 (N_3201,N_922,N_1462);
xor U3202 (N_3202,N_2061,N_81);
and U3203 (N_3203,N_2237,N_2843);
xnor U3204 (N_3204,N_619,N_2333);
or U3205 (N_3205,N_2838,N_2551);
nor U3206 (N_3206,N_776,N_1777);
xnor U3207 (N_3207,N_1540,N_701);
and U3208 (N_3208,N_273,N_1773);
and U3209 (N_3209,N_728,N_2284);
and U3210 (N_3210,N_2053,N_2601);
xnor U3211 (N_3211,N_1944,N_2920);
nand U3212 (N_3212,N_1150,N_1578);
nor U3213 (N_3213,N_958,N_2177);
xor U3214 (N_3214,N_735,N_2712);
or U3215 (N_3215,N_2358,N_1648);
nor U3216 (N_3216,N_1485,N_1687);
and U3217 (N_3217,N_1946,N_2107);
xnor U3218 (N_3218,N_2702,N_1260);
nor U3219 (N_3219,N_1122,N_2529);
or U3220 (N_3220,N_1107,N_2957);
nand U3221 (N_3221,N_2695,N_129);
nor U3222 (N_3222,N_1285,N_1174);
nand U3223 (N_3223,N_2282,N_3006);
xnor U3224 (N_3224,N_2645,N_3001);
or U3225 (N_3225,N_1776,N_206);
nand U3226 (N_3226,N_1187,N_915);
and U3227 (N_3227,N_2597,N_2747);
or U3228 (N_3228,N_1661,N_2998);
and U3229 (N_3229,N_583,N_2229);
or U3230 (N_3230,N_272,N_2932);
nor U3231 (N_3231,N_545,N_1560);
and U3232 (N_3232,N_926,N_218);
and U3233 (N_3233,N_598,N_3121);
and U3234 (N_3234,N_1994,N_2627);
or U3235 (N_3235,N_2739,N_948);
xnor U3236 (N_3236,N_2696,N_2287);
nand U3237 (N_3237,N_2418,N_1097);
xor U3238 (N_3238,N_1880,N_592);
and U3239 (N_3239,N_651,N_2305);
xnor U3240 (N_3240,N_464,N_1503);
nand U3241 (N_3241,N_1408,N_1163);
and U3242 (N_3242,N_2522,N_1223);
and U3243 (N_3243,N_2134,N_1445);
and U3244 (N_3244,N_667,N_1741);
and U3245 (N_3245,N_860,N_2209);
nor U3246 (N_3246,N_1078,N_1536);
xor U3247 (N_3247,N_2798,N_612);
nor U3248 (N_3248,N_2839,N_2077);
nor U3249 (N_3249,N_2547,N_700);
xnor U3250 (N_3250,N_2891,N_383);
xnor U3251 (N_3251,N_307,N_1940);
xnor U3252 (N_3252,N_2617,N_1338);
and U3253 (N_3253,N_3111,N_521);
nand U3254 (N_3254,N_1724,N_568);
or U3255 (N_3255,N_940,N_1073);
nor U3256 (N_3256,N_769,N_1572);
xnor U3257 (N_3257,N_2560,N_2506);
xor U3258 (N_3258,N_2511,N_1189);
nand U3259 (N_3259,N_109,N_1768);
nand U3260 (N_3260,N_376,N_2599);
xor U3261 (N_3261,N_1027,N_3117);
nand U3262 (N_3262,N_1309,N_152);
nor U3263 (N_3263,N_1827,N_1436);
and U3264 (N_3264,N_1937,N_11);
xor U3265 (N_3265,N_54,N_1293);
or U3266 (N_3266,N_2173,N_3094);
and U3267 (N_3267,N_236,N_3123);
nor U3268 (N_3268,N_854,N_280);
nand U3269 (N_3269,N_688,N_153);
nand U3270 (N_3270,N_2189,N_1790);
and U3271 (N_3271,N_2774,N_2910);
nor U3272 (N_3272,N_2996,N_1282);
nand U3273 (N_3273,N_1885,N_1422);
and U3274 (N_3274,N_1393,N_1755);
nor U3275 (N_3275,N_2896,N_2240);
and U3276 (N_3276,N_481,N_431);
or U3277 (N_3277,N_179,N_1705);
and U3278 (N_3278,N_2937,N_2572);
and U3279 (N_3279,N_577,N_1821);
xor U3280 (N_3280,N_2647,N_1888);
nand U3281 (N_3281,N_1489,N_2847);
or U3282 (N_3282,N_1575,N_39);
xor U3283 (N_3283,N_2852,N_214);
or U3284 (N_3284,N_3069,N_3098);
xor U3285 (N_3285,N_704,N_834);
xor U3286 (N_3286,N_2280,N_1923);
nand U3287 (N_3287,N_227,N_1134);
xnor U3288 (N_3288,N_2631,N_2801);
nand U3289 (N_3289,N_393,N_151);
xnor U3290 (N_3290,N_1523,N_1448);
nand U3291 (N_3291,N_2045,N_259);
or U3292 (N_3292,N_348,N_689);
xnor U3293 (N_3293,N_2255,N_48);
and U3294 (N_3294,N_2448,N_355);
nand U3295 (N_3295,N_380,N_2353);
xnor U3296 (N_3296,N_1605,N_2944);
or U3297 (N_3297,N_111,N_1972);
nand U3298 (N_3298,N_2454,N_3025);
and U3299 (N_3299,N_867,N_989);
and U3300 (N_3300,N_707,N_2168);
nor U3301 (N_3301,N_3071,N_2576);
nor U3302 (N_3302,N_1838,N_2513);
xor U3303 (N_3303,N_596,N_2635);
nand U3304 (N_3304,N_2703,N_184);
or U3305 (N_3305,N_358,N_1142);
xor U3306 (N_3306,N_293,N_1371);
and U3307 (N_3307,N_3101,N_1263);
nor U3308 (N_3308,N_1669,N_1841);
nand U3309 (N_3309,N_966,N_138);
nand U3310 (N_3310,N_2789,N_2351);
nand U3311 (N_3311,N_507,N_30);
xor U3312 (N_3312,N_1671,N_874);
or U3313 (N_3313,N_2857,N_2660);
or U3314 (N_3314,N_2016,N_1759);
xor U3315 (N_3315,N_2644,N_1662);
nand U3316 (N_3316,N_2244,N_1678);
nand U3317 (N_3317,N_1866,N_1303);
xnor U3318 (N_3318,N_99,N_2011);
nand U3319 (N_3319,N_1382,N_212);
or U3320 (N_3320,N_2462,N_552);
nand U3321 (N_3321,N_2380,N_2063);
or U3322 (N_3322,N_1155,N_1585);
nor U3323 (N_3323,N_2230,N_2374);
nor U3324 (N_3324,N_3011,N_1357);
and U3325 (N_3325,N_2112,N_27);
nand U3326 (N_3326,N_1913,N_2503);
nand U3327 (N_3327,N_3085,N_2434);
or U3328 (N_3328,N_12,N_1103);
and U3329 (N_3329,N_462,N_378);
xnor U3330 (N_3330,N_1049,N_604);
nand U3331 (N_3331,N_2971,N_2516);
nor U3332 (N_3332,N_2466,N_122);
xor U3333 (N_3333,N_782,N_1947);
or U3334 (N_3334,N_1315,N_1091);
and U3335 (N_3335,N_2952,N_3099);
or U3336 (N_3336,N_1221,N_713);
nand U3337 (N_3337,N_2141,N_2231);
and U3338 (N_3338,N_1370,N_2771);
or U3339 (N_3339,N_2805,N_1201);
or U3340 (N_3340,N_2867,N_2864);
xnor U3341 (N_3341,N_2036,N_1031);
nor U3342 (N_3342,N_1518,N_2766);
nand U3343 (N_3343,N_1531,N_1300);
nor U3344 (N_3344,N_1602,N_1264);
nor U3345 (N_3345,N_9,N_3093);
xnor U3346 (N_3346,N_180,N_1086);
nand U3347 (N_3347,N_1415,N_2356);
nand U3348 (N_3348,N_59,N_2127);
and U3349 (N_3349,N_925,N_2382);
and U3350 (N_3350,N_2406,N_235);
xor U3351 (N_3351,N_315,N_1989);
xnor U3352 (N_3352,N_255,N_1197);
nand U3353 (N_3353,N_1891,N_994);
nand U3354 (N_3354,N_680,N_912);
xnor U3355 (N_3355,N_395,N_1438);
and U3356 (N_3356,N_1116,N_2714);
xor U3357 (N_3357,N_1495,N_2677);
xor U3358 (N_3358,N_2171,N_2428);
nor U3359 (N_3359,N_501,N_675);
or U3360 (N_3360,N_2442,N_1214);
xnor U3361 (N_3361,N_2967,N_2978);
or U3362 (N_3362,N_194,N_2916);
or U3363 (N_3363,N_1261,N_250);
xnor U3364 (N_3364,N_1803,N_1360);
nor U3365 (N_3365,N_311,N_3089);
or U3366 (N_3366,N_1191,N_1576);
and U3367 (N_3367,N_3051,N_2038);
nor U3368 (N_3368,N_2737,N_1886);
nor U3369 (N_3369,N_461,N_553);
or U3370 (N_3370,N_1463,N_208);
xor U3371 (N_3371,N_1290,N_1809);
nand U3372 (N_3372,N_114,N_1858);
or U3373 (N_3373,N_1204,N_2412);
nand U3374 (N_3374,N_1610,N_2043);
xor U3375 (N_3375,N_2689,N_1520);
and U3376 (N_3376,N_1980,N_1646);
or U3377 (N_3377,N_674,N_626);
xor U3378 (N_3378,N_1123,N_1500);
and U3379 (N_3379,N_237,N_488);
nand U3380 (N_3380,N_2673,N_2410);
xnor U3381 (N_3381,N_2544,N_1513);
nand U3382 (N_3382,N_1063,N_2698);
xnor U3383 (N_3383,N_3070,N_2268);
and U3384 (N_3384,N_2056,N_1852);
or U3385 (N_3385,N_2012,N_2717);
or U3386 (N_3386,N_136,N_1159);
xnor U3387 (N_3387,N_121,N_1043);
nor U3388 (N_3388,N_2040,N_1988);
nor U3389 (N_3389,N_1728,N_594);
nor U3390 (N_3390,N_262,N_597);
nand U3391 (N_3391,N_2423,N_2709);
and U3392 (N_3392,N_344,N_1541);
or U3393 (N_3393,N_2598,N_1215);
xnor U3394 (N_3394,N_2652,N_2494);
nand U3395 (N_3395,N_832,N_1826);
nor U3396 (N_3396,N_2935,N_1016);
nor U3397 (N_3397,N_714,N_284);
or U3398 (N_3398,N_772,N_679);
nor U3399 (N_3399,N_2854,N_1553);
and U3400 (N_3400,N_1179,N_229);
xnor U3401 (N_3401,N_2403,N_2985);
or U3402 (N_3402,N_1795,N_791);
nor U3403 (N_3403,N_2666,N_1033);
nor U3404 (N_3404,N_1726,N_1651);
xnor U3405 (N_3405,N_327,N_1090);
nor U3406 (N_3406,N_471,N_2161);
nand U3407 (N_3407,N_833,N_1053);
xnor U3408 (N_3408,N_2340,N_1311);
and U3409 (N_3409,N_1475,N_2745);
and U3410 (N_3410,N_2267,N_736);
xnor U3411 (N_3411,N_2215,N_2893);
and U3412 (N_3412,N_2605,N_1919);
or U3413 (N_3413,N_440,N_652);
nand U3414 (N_3414,N_2172,N_74);
nor U3415 (N_3415,N_982,N_1524);
nand U3416 (N_3416,N_172,N_1681);
or U3417 (N_3417,N_325,N_985);
and U3418 (N_3418,N_949,N_1618);
nand U3419 (N_3419,N_1932,N_1854);
nand U3420 (N_3420,N_1899,N_1253);
or U3421 (N_3421,N_2882,N_23);
and U3422 (N_3422,N_2117,N_992);
nand U3423 (N_3423,N_2819,N_2729);
or U3424 (N_3424,N_2730,N_1908);
nor U3425 (N_3425,N_450,N_1138);
xor U3426 (N_3426,N_2554,N_1125);
and U3427 (N_3427,N_2977,N_331);
xor U3428 (N_3428,N_300,N_2279);
xnor U3429 (N_3429,N_805,N_1226);
or U3430 (N_3430,N_686,N_2178);
and U3431 (N_3431,N_1268,N_3034);
or U3432 (N_3432,N_645,N_1292);
xnor U3433 (N_3433,N_2700,N_3072);
nand U3434 (N_3434,N_2311,N_2349);
nor U3435 (N_3435,N_517,N_1644);
xnor U3436 (N_3436,N_173,N_1164);
and U3437 (N_3437,N_2846,N_2797);
xor U3438 (N_3438,N_2997,N_2271);
xnor U3439 (N_3439,N_1067,N_1959);
nor U3440 (N_3440,N_973,N_2759);
nand U3441 (N_3441,N_1596,N_1433);
or U3442 (N_3442,N_160,N_34);
nor U3443 (N_3443,N_2900,N_1504);
nand U3444 (N_3444,N_2118,N_1787);
xnor U3445 (N_3445,N_807,N_1151);
nor U3446 (N_3446,N_2779,N_362);
xor U3447 (N_3447,N_1346,N_540);
nand U3448 (N_3448,N_1961,N_1248);
xnor U3449 (N_3449,N_3108,N_199);
nand U3450 (N_3450,N_3060,N_238);
xor U3451 (N_3451,N_936,N_3017);
nor U3452 (N_3452,N_2580,N_1570);
and U3453 (N_3453,N_2197,N_677);
nor U3454 (N_3454,N_274,N_2122);
and U3455 (N_3455,N_1427,N_2947);
or U3456 (N_3456,N_555,N_459);
nand U3457 (N_3457,N_1341,N_1836);
nor U3458 (N_3458,N_251,N_896);
or U3459 (N_3459,N_1626,N_734);
and U3460 (N_3460,N_2969,N_1377);
xnor U3461 (N_3461,N_1353,N_68);
nand U3462 (N_3462,N_2102,N_163);
and U3463 (N_3463,N_2426,N_216);
and U3464 (N_3464,N_2938,N_722);
xnor U3465 (N_3465,N_1431,N_1679);
xnor U3466 (N_3466,N_2042,N_2588);
nand U3467 (N_3467,N_1343,N_512);
xor U3468 (N_3468,N_1326,N_942);
or U3469 (N_3469,N_2457,N_1563);
or U3470 (N_3470,N_1272,N_2567);
xnor U3471 (N_3471,N_929,N_1404);
xnor U3472 (N_3472,N_1794,N_2549);
nor U3473 (N_3473,N_2181,N_490);
xnor U3474 (N_3474,N_1745,N_790);
and U3475 (N_3475,N_1772,N_340);
nor U3476 (N_3476,N_220,N_3106);
nand U3477 (N_3477,N_1102,N_58);
xnor U3478 (N_3478,N_2310,N_2460);
nor U3479 (N_3479,N_642,N_1006);
nor U3480 (N_3480,N_1896,N_1428);
or U3481 (N_3481,N_276,N_1586);
nor U3482 (N_3482,N_1539,N_36);
xnor U3483 (N_3483,N_1365,N_1479);
xnor U3484 (N_3484,N_1339,N_1842);
nor U3485 (N_3485,N_513,N_2908);
nand U3486 (N_3486,N_601,N_2905);
nor U3487 (N_3487,N_143,N_1169);
and U3488 (N_3488,N_2366,N_715);
or U3489 (N_3489,N_1133,N_1258);
and U3490 (N_3490,N_2636,N_1275);
nor U3491 (N_3491,N_1635,N_2481);
and U3492 (N_3492,N_2497,N_1684);
nor U3493 (N_3493,N_1440,N_1753);
nor U3494 (N_3494,N_2620,N_2565);
and U3495 (N_3495,N_2357,N_224);
nor U3496 (N_3496,N_338,N_1711);
and U3497 (N_3497,N_2166,N_1906);
and U3498 (N_3498,N_2536,N_2039);
xnor U3499 (N_3499,N_1421,N_2022);
and U3500 (N_3500,N_2800,N_1259);
or U3501 (N_3501,N_2590,N_2989);
nor U3502 (N_3502,N_2048,N_110);
xnor U3503 (N_3503,N_2639,N_1653);
xnor U3504 (N_3504,N_267,N_719);
xor U3505 (N_3505,N_2085,N_1655);
or U3506 (N_3506,N_885,N_1200);
xnor U3507 (N_3507,N_100,N_1114);
nand U3508 (N_3508,N_275,N_2436);
nand U3509 (N_3509,N_1783,N_209);
xnor U3510 (N_3510,N_1266,N_2806);
and U3511 (N_3511,N_2135,N_2548);
and U3512 (N_3512,N_2114,N_2818);
or U3513 (N_3513,N_2788,N_1281);
and U3514 (N_3514,N_2973,N_802);
and U3515 (N_3515,N_1695,N_484);
xnor U3516 (N_3516,N_1098,N_361);
nor U3517 (N_3517,N_312,N_967);
nor U3518 (N_3518,N_207,N_3020);
xor U3519 (N_3519,N_3107,N_2324);
and U3520 (N_3520,N_460,N_1639);
nand U3521 (N_3521,N_299,N_2467);
nand U3522 (N_3522,N_2828,N_70);
nor U3523 (N_3523,N_632,N_1957);
and U3524 (N_3524,N_899,N_2608);
xor U3525 (N_3525,N_1108,N_831);
and U3526 (N_3526,N_981,N_472);
or U3527 (N_3527,N_166,N_1530);
and U3528 (N_3528,N_1921,N_774);
or U3529 (N_3529,N_876,N_1686);
and U3530 (N_3530,N_1625,N_1855);
or U3531 (N_3531,N_1879,N_2325);
xor U3532 (N_3532,N_2878,N_711);
or U3533 (N_3533,N_2004,N_3084);
xor U3534 (N_3534,N_3086,N_581);
xor U3535 (N_3535,N_465,N_1407);
nor U3536 (N_3536,N_2869,N_1725);
or U3537 (N_3537,N_3103,N_656);
or U3538 (N_3538,N_2850,N_396);
nor U3539 (N_3539,N_2691,N_2261);
nor U3540 (N_3540,N_2139,N_1432);
or U3541 (N_3541,N_525,N_1434);
nand U3542 (N_3542,N_741,N_2276);
nand U3543 (N_3543,N_964,N_432);
or U3544 (N_3544,N_1136,N_478);
nor U3545 (N_3545,N_3065,N_1351);
nand U3546 (N_3546,N_1757,N_1514);
xor U3547 (N_3547,N_1731,N_1727);
nand U3548 (N_3548,N_1140,N_2868);
or U3549 (N_3549,N_600,N_1864);
xor U3550 (N_3550,N_1549,N_2272);
and U3551 (N_3551,N_780,N_51);
or U3552 (N_3552,N_1829,N_1770);
or U3553 (N_3553,N_988,N_932);
and U3554 (N_3554,N_535,N_2365);
or U3555 (N_3555,N_532,N_2743);
nor U3556 (N_3556,N_2624,N_1109);
nor U3557 (N_3557,N_1743,N_2095);
xor U3558 (N_3558,N_603,N_1166);
xor U3559 (N_3559,N_156,N_2507);
nor U3560 (N_3560,N_1619,N_1287);
xor U3561 (N_3561,N_2972,N_590);
or U3562 (N_3562,N_2519,N_1419);
and U3563 (N_3563,N_1167,N_3083);
xnor U3564 (N_3564,N_894,N_1627);
nand U3565 (N_3565,N_838,N_2811);
or U3566 (N_3566,N_1609,N_1249);
nand U3567 (N_3567,N_2674,N_2283);
nor U3568 (N_3568,N_2451,N_1364);
nor U3569 (N_3569,N_1218,N_1933);
or U3570 (N_3570,N_2784,N_2780);
nor U3571 (N_3571,N_738,N_2749);
nand U3572 (N_3572,N_848,N_493);
and U3573 (N_3573,N_2254,N_2955);
xor U3574 (N_3574,N_352,N_2465);
nand U3575 (N_3575,N_3050,N_2658);
xnor U3576 (N_3576,N_2438,N_1331);
or U3577 (N_3577,N_2662,N_2236);
nand U3578 (N_3578,N_2315,N_624);
nand U3579 (N_3579,N_1708,N_2754);
nand U3580 (N_3580,N_2592,N_923);
nand U3581 (N_3581,N_2185,N_2678);
nand U3582 (N_3582,N_1308,N_3021);
and U3583 (N_3583,N_947,N_1235);
nand U3584 (N_3584,N_1981,N_2706);
and U3585 (N_3585,N_1938,N_2377);
xor U3586 (N_3586,N_247,N_2224);
and U3587 (N_3587,N_2025,N_1190);
nand U3588 (N_3588,N_3053,N_2940);
or U3589 (N_3589,N_1205,N_1461);
or U3590 (N_3590,N_319,N_2918);
or U3591 (N_3591,N_2295,N_2245);
nor U3592 (N_3592,N_1958,N_566);
xnor U3593 (N_3593,N_1825,N_1361);
and U3594 (N_3594,N_2387,N_1914);
xor U3595 (N_3595,N_761,N_93);
xnor U3596 (N_3596,N_2833,N_1188);
nand U3597 (N_3597,N_1397,N_888);
nand U3598 (N_3598,N_368,N_1367);
nand U3599 (N_3599,N_1130,N_2830);
xnor U3600 (N_3600,N_1784,N_2094);
and U3601 (N_3601,N_31,N_2802);
nor U3602 (N_3602,N_494,N_1245);
or U3603 (N_3603,N_1736,N_723);
nor U3604 (N_3604,N_2625,N_2354);
or U3605 (N_3605,N_1974,N_938);
or U3606 (N_3606,N_1323,N_332);
or U3607 (N_3607,N_2075,N_476);
or U3608 (N_3608,N_1481,N_1577);
nand U3609 (N_3609,N_2078,N_2408);
and U3610 (N_3610,N_526,N_2005);
nor U3611 (N_3611,N_633,N_980);
nand U3612 (N_3612,N_2555,N_2923);
nor U3613 (N_3613,N_328,N_1079);
nand U3614 (N_3614,N_984,N_2182);
or U3615 (N_3615,N_2212,N_659);
nand U3616 (N_3616,N_181,N_1508);
or U3617 (N_3617,N_1358,N_1143);
and U3618 (N_3618,N_913,N_2247);
nor U3619 (N_3619,N_105,N_1088);
xnor U3620 (N_3620,N_278,N_509);
nand U3621 (N_3621,N_2961,N_1267);
or U3622 (N_3622,N_3029,N_1294);
and U3623 (N_3623,N_1556,N_669);
and U3624 (N_3624,N_1922,N_1769);
or U3625 (N_3625,N_2655,N_1161);
nor U3626 (N_3626,N_1643,N_1291);
and U3627 (N_3627,N_2836,N_930);
and U3628 (N_3628,N_1680,N_1929);
xor U3629 (N_3629,N_2734,N_1041);
or U3630 (N_3630,N_3024,N_2711);
nand U3631 (N_3631,N_1177,N_2108);
and U3632 (N_3632,N_268,N_3014);
nand U3633 (N_3633,N_2347,N_2007);
nand U3634 (N_3634,N_1354,N_754);
nand U3635 (N_3635,N_1488,N_2088);
xnor U3636 (N_3636,N_480,N_1173);
and U3637 (N_3637,N_297,N_131);
or U3638 (N_3638,N_400,N_745);
or U3639 (N_3639,N_2928,N_1149);
or U3640 (N_3640,N_2898,N_241);
xor U3641 (N_3641,N_3008,N_2637);
or U3642 (N_3642,N_1774,N_2621);
xnor U3643 (N_3643,N_1699,N_359);
nor U3644 (N_3644,N_1657,N_2775);
nand U3645 (N_3645,N_2006,N_1312);
or U3646 (N_3646,N_2772,N_260);
nand U3647 (N_3647,N_1286,N_1252);
or U3648 (N_3648,N_1857,N_2610);
and U3649 (N_3649,N_3082,N_1663);
or U3650 (N_3650,N_1322,N_1232);
nor U3651 (N_3651,N_1546,N_200);
xor U3652 (N_3652,N_2687,N_2630);
or U3653 (N_3653,N_1324,N_219);
or U3654 (N_3654,N_2456,N_1194);
nand U3655 (N_3655,N_2713,N_2299);
nor U3656 (N_3656,N_2326,N_112);
xnor U3657 (N_3657,N_2603,N_2623);
nand U3658 (N_3658,N_349,N_1320);
or U3659 (N_3659,N_306,N_1614);
nand U3660 (N_3660,N_1273,N_2962);
or U3661 (N_3661,N_1995,N_2037);
nor U3662 (N_3662,N_2330,N_2907);
and U3663 (N_3663,N_574,N_803);
and U3664 (N_3664,N_824,N_1172);
or U3665 (N_3665,N_1652,N_217);
nor U3666 (N_3666,N_998,N_1051);
xnor U3667 (N_3667,N_623,N_2849);
xor U3668 (N_3668,N_1758,N_1111);
nor U3669 (N_3669,N_2521,N_582);
or U3670 (N_3670,N_613,N_1059);
xnor U3671 (N_3671,N_858,N_2723);
and U3672 (N_3672,N_430,N_2760);
nor U3673 (N_3673,N_2770,N_2979);
and U3674 (N_3674,N_901,N_2401);
nand U3675 (N_3675,N_1387,N_2106);
and U3676 (N_3676,N_1670,N_1442);
or U3677 (N_3677,N_97,N_2787);
xor U3678 (N_3678,N_1454,N_808);
nand U3679 (N_3679,N_3000,N_324);
xor U3680 (N_3680,N_1470,N_2407);
nand U3681 (N_3681,N_1534,N_573);
and U3682 (N_3682,N_763,N_2219);
or U3683 (N_3683,N_1963,N_845);
nand U3684 (N_3684,N_1782,N_2110);
xnor U3685 (N_3685,N_3032,N_350);
xor U3686 (N_3686,N_2708,N_2697);
and U3687 (N_3687,N_2067,N_382);
or U3688 (N_3688,N_2518,N_1129);
xor U3689 (N_3689,N_2029,N_1976);
xnor U3690 (N_3690,N_2336,N_2028);
nor U3691 (N_3691,N_115,N_232);
nand U3692 (N_3692,N_157,N_2501);
nor U3693 (N_3693,N_2143,N_534);
and U3694 (N_3694,N_1469,N_171);
nor U3695 (N_3695,N_1110,N_730);
nor U3696 (N_3696,N_1982,N_2594);
or U3697 (N_3697,N_2479,N_847);
nor U3698 (N_3698,N_2119,N_2649);
nor U3699 (N_3699,N_733,N_289);
nor U3700 (N_3700,N_1316,N_1017);
nor U3701 (N_3701,N_1117,N_1271);
and U3702 (N_3702,N_871,N_2715);
nand U3703 (N_3703,N_1391,N_294);
nor U3704 (N_3704,N_257,N_2781);
nand U3705 (N_3705,N_1398,N_1579);
xnor U3706 (N_3706,N_1449,N_2825);
and U3707 (N_3707,N_2184,N_2589);
or U3708 (N_3708,N_502,N_458);
or U3709 (N_3709,N_1065,N_1760);
xor U3710 (N_3710,N_148,N_2384);
nor U3711 (N_3711,N_2096,N_423);
and U3712 (N_3712,N_1617,N_1732);
or U3713 (N_3713,N_2885,N_1688);
nor U3714 (N_3714,N_580,N_1990);
nand U3715 (N_3715,N_630,N_21);
and U3716 (N_3716,N_1486,N_1762);
and U3717 (N_3717,N_2470,N_823);
and U3718 (N_3718,N_387,N_2402);
nand U3719 (N_3719,N_2090,N_690);
xor U3720 (N_3720,N_1081,N_2364);
nand U3721 (N_3721,N_2203,N_718);
or U3722 (N_3722,N_1713,N_843);
xnor U3723 (N_3723,N_2121,N_302);
and U3724 (N_3724,N_561,N_1222);
nand U3725 (N_3725,N_969,N_3031);
nor U3726 (N_3726,N_2871,N_1395);
and U3727 (N_3727,N_1069,N_1505);
xor U3728 (N_3728,N_2158,N_617);
nor U3729 (N_3729,N_2704,N_2449);
and U3730 (N_3730,N_2270,N_2277);
nor U3731 (N_3731,N_408,N_2131);
nand U3732 (N_3732,N_295,N_2919);
nand U3733 (N_3733,N_3066,N_189);
nand U3734 (N_3734,N_2101,N_2359);
xnor U3735 (N_3735,N_2853,N_1359);
or U3736 (N_3736,N_1650,N_1941);
xor U3737 (N_3737,N_1372,N_231);
xnor U3738 (N_3738,N_2650,N_137);
and U3739 (N_3739,N_1837,N_1876);
xnor U3740 (N_3740,N_602,N_2595);
xnor U3741 (N_3741,N_1180,N_2870);
and U3742 (N_3742,N_155,N_84);
or U3743 (N_3743,N_510,N_664);
nand U3744 (N_3744,N_1574,N_1093);
or U3745 (N_3745,N_2072,N_2093);
nand U3746 (N_3746,N_1230,N_1830);
or U3747 (N_3747,N_2782,N_2485);
nor U3748 (N_3748,N_2640,N_33);
nor U3749 (N_3749,N_2323,N_125);
xor U3750 (N_3750,N_2217,N_3105);
nand U3751 (N_3751,N_233,N_2570);
or U3752 (N_3752,N_2653,N_1611);
or U3753 (N_3753,N_2471,N_2822);
and U3754 (N_3754,N_740,N_756);
nand U3755 (N_3755,N_2213,N_2345);
or U3756 (N_3756,N_2533,N_1057);
nor U3757 (N_3757,N_1867,N_618);
or U3758 (N_3758,N_1924,N_1135);
nor U3759 (N_3759,N_2027,N_1856);
and U3760 (N_3760,N_437,N_856);
or U3761 (N_3761,N_2433,N_1642);
or U3762 (N_3762,N_1493,N_1127);
xnor U3763 (N_3763,N_198,N_2091);
or U3764 (N_3764,N_2050,N_2568);
and U3765 (N_3765,N_2285,N_1243);
or U3766 (N_3766,N_705,N_1738);
xnor U3767 (N_3767,N_641,N_2472);
and U3768 (N_3768,N_2648,N_1411);
nand U3769 (N_3769,N_990,N_3049);
and U3770 (N_3770,N_1714,N_37);
or U3771 (N_3771,N_2814,N_2807);
and U3772 (N_3772,N_2206,N_2622);
or U3773 (N_3773,N_1340,N_902);
xnor U3774 (N_3774,N_1878,N_2953);
and U3775 (N_3775,N_2738,N_2400);
xnor U3776 (N_3776,N_2899,N_1791);
nand U3777 (N_3777,N_1729,N_2582);
or U3778 (N_3778,N_1105,N_1517);
nor U3779 (N_3779,N_1280,N_644);
and U3780 (N_3780,N_1979,N_2409);
nand U3781 (N_3781,N_778,N_411);
nor U3782 (N_3782,N_2473,N_2338);
and U3783 (N_3783,N_3112,N_2201);
xnor U3784 (N_3784,N_316,N_2534);
or U3785 (N_3785,N_742,N_692);
nor U3786 (N_3786,N_489,N_2395);
xor U3787 (N_3787,N_2492,N_385);
or U3788 (N_3788,N_1378,N_1698);
nand U3789 (N_3789,N_1401,N_92);
nor U3790 (N_3790,N_2634,N_193);
nand U3791 (N_3791,N_1023,N_341);
nand U3792 (N_3792,N_1636,N_83);
nand U3793 (N_3793,N_1975,N_2227);
and U3794 (N_3794,N_556,N_1615);
or U3795 (N_3795,N_770,N_2191);
nand U3796 (N_3796,N_1147,N_3119);
nor U3797 (N_3797,N_3087,N_2126);
nand U3798 (N_3798,N_1342,N_296);
xor U3799 (N_3799,N_1935,N_1945);
nor U3800 (N_3800,N_1526,N_2424);
and U3801 (N_3801,N_572,N_1094);
xnor U3802 (N_3802,N_1998,N_205);
and U3803 (N_3803,N_2301,N_451);
nand U3804 (N_3804,N_2092,N_2413);
and U3805 (N_3805,N_1347,N_1840);
or U3806 (N_3806,N_3002,N_3064);
and U3807 (N_3807,N_1953,N_1689);
nor U3808 (N_3808,N_2505,N_1363);
nand U3809 (N_3809,N_851,N_85);
nor U3810 (N_3810,N_606,N_2222);
or U3811 (N_3811,N_2017,N_45);
nand U3812 (N_3812,N_977,N_2884);
nor U3813 (N_3813,N_1209,N_2469);
nor U3814 (N_3814,N_1955,N_2569);
and U3815 (N_3815,N_2872,N_1074);
and U3816 (N_3816,N_374,N_1668);
xnor U3817 (N_3817,N_1238,N_89);
or U3818 (N_3818,N_1018,N_2186);
or U3819 (N_3819,N_14,N_2320);
or U3820 (N_3820,N_1740,N_1457);
nor U3821 (N_3821,N_55,N_71);
and U3822 (N_3822,N_2959,N_1744);
nand U3823 (N_3823,N_2930,N_775);
nor U3824 (N_3824,N_239,N_2499);
nor U3825 (N_3825,N_1608,N_2286);
nand U3826 (N_3826,N_781,N_177);
nor U3827 (N_3827,N_62,N_321);
and U3828 (N_3828,N_2651,N_784);
or U3829 (N_3829,N_1024,N_3055);
nor U3830 (N_3830,N_3015,N_684);
nand U3831 (N_3831,N_2581,N_1336);
and U3832 (N_3832,N_1936,N_787);
nand U3833 (N_3833,N_3036,N_1203);
xor U3834 (N_3834,N_2982,N_1237);
xnor U3835 (N_3835,N_1516,N_308);
nand U3836 (N_3836,N_1597,N_815);
xnor U3837 (N_3837,N_2252,N_2238);
nand U3838 (N_3838,N_279,N_483);
nand U3839 (N_3839,N_2970,N_2394);
or U3840 (N_3840,N_96,N_2273);
nand U3841 (N_3841,N_204,N_107);
or U3842 (N_3842,N_2146,N_1555);
and U3843 (N_3843,N_2099,N_375);
xnor U3844 (N_3844,N_126,N_1765);
nand U3845 (N_3845,N_1843,N_2951);
nor U3846 (N_3846,N_2912,N_2373);
or U3847 (N_3847,N_1895,N_113);
xor U3848 (N_3848,N_1198,N_2720);
and U3849 (N_3849,N_1785,N_2437);
nor U3850 (N_3850,N_1441,N_1716);
and U3851 (N_3851,N_889,N_41);
and U3852 (N_3852,N_2509,N_859);
xor U3853 (N_3853,N_3073,N_1633);
xnor U3854 (N_3854,N_142,N_1160);
and U3855 (N_3855,N_2542,N_457);
or U3856 (N_3856,N_1484,N_2162);
or U3857 (N_3857,N_1849,N_139);
nor U3858 (N_3858,N_2491,N_2378);
nand U3859 (N_3859,N_1390,N_1719);
nand U3860 (N_3860,N_1499,N_1003);
or U3861 (N_3861,N_1375,N_2541);
or U3862 (N_3862,N_317,N_1634);
xnor U3863 (N_3863,N_1321,N_2223);
xor U3864 (N_3864,N_1423,N_2266);
nor U3865 (N_3865,N_1224,N_2724);
xnor U3866 (N_3866,N_2915,N_3028);
and U3867 (N_3867,N_1460,N_643);
xnor U3868 (N_3868,N_760,N_971);
or U3869 (N_3869,N_2894,N_1565);
xnor U3870 (N_3870,N_962,N_1195);
nand U3871 (N_3871,N_244,N_591);
nor U3872 (N_3872,N_1413,N_1584);
xnor U3873 (N_3873,N_230,N_1580);
xor U3874 (N_3874,N_1385,N_895);
xor U3875 (N_3875,N_1380,N_384);
or U3876 (N_3876,N_32,N_970);
xor U3877 (N_3877,N_2435,N_1631);
xor U3878 (N_3878,N_564,N_1970);
and U3879 (N_3879,N_1862,N_3);
nand U3880 (N_3880,N_3059,N_1096);
xnor U3881 (N_3881,N_2752,N_2105);
nand U3882 (N_3882,N_1869,N_2071);
nor U3883 (N_3883,N_3113,N_369);
and U3884 (N_3884,N_2816,N_2086);
nand U3885 (N_3885,N_1178,N_846);
or U3886 (N_3886,N_1811,N_291);
nand U3887 (N_3887,N_82,N_2104);
or U3888 (N_3888,N_2153,N_2024);
or U3889 (N_3889,N_266,N_176);
nand U3890 (N_3890,N_19,N_398);
nor U3891 (N_3891,N_403,N_1416);
nor U3892 (N_3892,N_621,N_3039);
and U3893 (N_3893,N_1877,N_2753);
nor U3894 (N_3894,N_419,N_1522);
xnor U3895 (N_3895,N_2573,N_167);
and U3896 (N_3896,N_1106,N_7);
xor U3897 (N_3897,N_1250,N_1806);
or U3898 (N_3898,N_2431,N_2342);
nor U3899 (N_3899,N_820,N_202);
and U3900 (N_3900,N_60,N_2524);
and U3901 (N_3901,N_2054,N_1477);
nand U3902 (N_3902,N_2559,N_2389);
nand U3903 (N_3903,N_696,N_63);
nor U3904 (N_3904,N_422,N_1046);
xor U3905 (N_3905,N_1464,N_671);
nand U3906 (N_3906,N_2577,N_263);
nand U3907 (N_3907,N_2441,N_3077);
nand U3908 (N_3908,N_2537,N_35);
nand U3909 (N_3909,N_1848,N_439);
nand U3910 (N_3910,N_2602,N_960);
or U3911 (N_3911,N_201,N_1182);
nor U3912 (N_3912,N_2773,N_1170);
nor U3913 (N_3913,N_1384,N_648);
or U3914 (N_3914,N_1751,N_2525);
and U3915 (N_3915,N_1601,N_38);
nor U3916 (N_3916,N_1590,N_2539);
xnor U3917 (N_3917,N_1394,N_371);
nor U3918 (N_3918,N_1020,N_1604);
nor U3919 (N_3919,N_1026,N_636);
xnor U3920 (N_3920,N_2615,N_1999);
xnor U3921 (N_3921,N_2019,N_318);
nor U3922 (N_3922,N_2137,N_1873);
nor U3923 (N_3923,N_2232,N_2379);
xnor U3924 (N_3924,N_2490,N_2921);
nor U3925 (N_3925,N_2880,N_1217);
xnor U3926 (N_3926,N_1567,N_2512);
and U3927 (N_3927,N_453,N_245);
or U3928 (N_3928,N_442,N_2484);
xnor U3929 (N_3929,N_762,N_2123);
and U3930 (N_3930,N_2587,N_1764);
or U3931 (N_3931,N_1456,N_2082);
and U3932 (N_3932,N_2632,N_1084);
nor U3933 (N_3933,N_427,N_2686);
nand U3934 (N_3934,N_1747,N_717);
xor U3935 (N_3935,N_282,N_2561);
nor U3936 (N_3936,N_1297,N_495);
nor U3937 (N_3937,N_1298,N_599);
nand U3938 (N_3938,N_2297,N_1894);
xor U3939 (N_3939,N_785,N_3067);
and U3940 (N_3940,N_409,N_305);
and U3941 (N_3941,N_197,N_2721);
nor U3942 (N_3942,N_283,N_2532);
nand U3943 (N_3943,N_28,N_3076);
nand U3944 (N_3944,N_2163,N_976);
and U3945 (N_3945,N_2155,N_554);
or U3946 (N_3946,N_865,N_1589);
xnor U3947 (N_3947,N_1694,N_2430);
xor U3948 (N_3948,N_254,N_2487);
xnor U3949 (N_3949,N_124,N_628);
nand U3950 (N_3950,N_2152,N_134);
xor U3951 (N_3951,N_265,N_694);
nand U3952 (N_3952,N_499,N_2445);
and U3953 (N_3953,N_2823,N_1443);
xnor U3954 (N_3954,N_1011,N_2432);
xnor U3955 (N_3955,N_2820,N_1196);
or U3956 (N_3956,N_228,N_405);
nor U3957 (N_3957,N_1682,N_607);
or U3958 (N_3958,N_133,N_892);
nand U3959 (N_3959,N_1497,N_893);
and U3960 (N_3960,N_1956,N_390);
xnor U3961 (N_3961,N_354,N_1969);
or U3962 (N_3962,N_1255,N_367);
or U3963 (N_3963,N_2170,N_2187);
xnor U3964 (N_3964,N_520,N_2069);
nand U3965 (N_3965,N_1859,N_1872);
nor U3966 (N_3966,N_2455,N_3019);
or U3967 (N_3967,N_190,N_3046);
or U3968 (N_3968,N_945,N_2370);
xnor U3969 (N_3969,N_2300,N_864);
nor U3970 (N_3970,N_1622,N_3100);
and U3971 (N_3971,N_1403,N_1893);
nor U3972 (N_3972,N_1376,N_588);
or U3973 (N_3973,N_1156,N_2986);
xor U3974 (N_3974,N_2726,N_813);
or U3975 (N_3975,N_2926,N_516);
xnor U3976 (N_3976,N_2386,N_531);
xor U3977 (N_3977,N_905,N_1807);
nor U3978 (N_3978,N_953,N_933);
nor U3979 (N_3979,N_301,N_1402);
xnor U3980 (N_3980,N_3038,N_937);
nand U3981 (N_3981,N_1863,N_2009);
xor U3982 (N_3982,N_794,N_3115);
nor U3983 (N_3983,N_1414,N_979);
or U3984 (N_3984,N_1916,N_928);
or U3985 (N_3985,N_2474,N_753);
xnor U3986 (N_3986,N_2304,N_2860);
nor U3987 (N_3987,N_1032,N_1943);
xnor U3988 (N_3988,N_1379,N_2502);
or U3989 (N_3989,N_2327,N_1928);
or U3990 (N_3990,N_2874,N_3078);
or U3991 (N_3991,N_2844,N_2855);
or U3992 (N_3992,N_2664,N_187);
xnor U3993 (N_3993,N_1834,N_2768);
and U3994 (N_3994,N_377,N_1965);
nor U3995 (N_3995,N_2486,N_1665);
nor U3996 (N_3996,N_2316,N_1950);
or U3997 (N_3997,N_2515,N_2198);
xor U3998 (N_3998,N_1833,N_2109);
xor U3999 (N_3999,N_1529,N_1257);
and U4000 (N_4000,N_178,N_898);
nor U4001 (N_4001,N_2892,N_2942);
xnor U4002 (N_4002,N_2530,N_287);
and U4003 (N_4003,N_1702,N_466);
nand U4004 (N_4004,N_2165,N_2321);
and U4005 (N_4005,N_2783,N_1571);
or U4006 (N_4006,N_1192,N_668);
nor U4007 (N_4007,N_1798,N_1673);
and U4008 (N_4008,N_1072,N_40);
nor U4009 (N_4009,N_758,N_941);
xnor U4010 (N_4010,N_2682,N_435);
or U4011 (N_4011,N_1676,N_346);
or U4012 (N_4012,N_708,N_2661);
or U4013 (N_4013,N_2196,N_1749);
nand U4014 (N_4014,N_2906,N_578);
nand U4015 (N_4015,N_1846,N_3109);
xnor U4016 (N_4016,N_1816,N_1019);
nand U4017 (N_4017,N_2879,N_1366);
xnor U4018 (N_4018,N_2427,N_829);
nand U4019 (N_4019,N_421,N_2463);
nor U4020 (N_4020,N_1987,N_2993);
or U4021 (N_4021,N_1701,N_830);
nand U4022 (N_4022,N_13,N_1451);
and U4023 (N_4023,N_1591,N_347);
nor U4024 (N_4024,N_356,N_529);
and U4025 (N_4025,N_2992,N_486);
nand U4026 (N_4026,N_2157,N_1796);
nand U4027 (N_4027,N_2190,N_2690);
xor U4028 (N_4028,N_691,N_1832);
or U4029 (N_4029,N_2719,N_943);
nor U4030 (N_4030,N_269,N_2444);
xnor U4031 (N_4031,N_1240,N_818);
nor U4032 (N_4032,N_1897,N_2176);
or U4033 (N_4033,N_2446,N_1779);
nor U4034 (N_4034,N_2361,N_827);
nand U4035 (N_4035,N_2762,N_1700);
and U4036 (N_4036,N_1502,N_783);
nand U4037 (N_4037,N_118,N_721);
nor U4038 (N_4038,N_570,N_18);
nor U4039 (N_4039,N_2520,N_1284);
nand U4040 (N_4040,N_102,N_3118);
or U4041 (N_4041,N_309,N_2945);
xnor U4042 (N_4042,N_956,N_1720);
xor U4043 (N_4043,N_2543,N_505);
or U4044 (N_4044,N_547,N_2523);
and U4045 (N_4045,N_1389,N_72);
nand U4046 (N_4046,N_1012,N_2575);
xnor U4047 (N_4047,N_2517,N_1501);
xor U4048 (N_4048,N_290,N_750);
and U4049 (N_4049,N_2001,N_2566);
or U4050 (N_4050,N_2552,N_2769);
nor U4051 (N_4051,N_2943,N_1145);
nand U4052 (N_4052,N_1001,N_2999);
xor U4053 (N_4053,N_2068,N_2332);
or U4054 (N_4054,N_3114,N_2929);
and U4055 (N_4055,N_2675,N_2968);
and U4056 (N_4056,N_2015,N_1115);
or U4057 (N_4057,N_685,N_391);
xnor U4058 (N_4058,N_1158,N_434);
and U4059 (N_4059,N_1690,N_1767);
or U4060 (N_4060,N_1064,N_2116);
nand U4061 (N_4061,N_2574,N_3095);
nor U4062 (N_4062,N_1455,N_660);
or U4063 (N_4063,N_786,N_1047);
xnor U4064 (N_4064,N_1822,N_145);
xnor U4065 (N_4065,N_66,N_357);
or U4066 (N_4066,N_1313,N_571);
nand U4067 (N_4067,N_539,N_866);
nor U4068 (N_4068,N_270,N_890);
nand U4069 (N_4069,N_2670,N_836);
or U4070 (N_4070,N_3004,N_2241);
xnor U4071 (N_4071,N_1234,N_445);
and U4072 (N_4072,N_2464,N_1332);
and U4073 (N_4073,N_1100,N_372);
nor U4074 (N_4074,N_1472,N_2578);
nand U4075 (N_4075,N_2368,N_154);
xor U4076 (N_4076,N_1638,N_868);
and U4077 (N_4077,N_2540,N_2562);
or U4078 (N_4078,N_855,N_1562);
nor U4079 (N_4079,N_1055,N_2841);
xnor U4080 (N_4080,N_1124,N_1473);
nand U4081 (N_4081,N_2718,N_1126);
xnor U4082 (N_4082,N_2861,N_1692);
and U4083 (N_4083,N_1528,N_1162);
nor U4084 (N_4084,N_3052,N_2618);
and U4085 (N_4085,N_3016,N_1992);
nor U4086 (N_4086,N_1659,N_454);
xor U4087 (N_4087,N_755,N_2393);
nand U4088 (N_4088,N_1588,N_2180);
or U4089 (N_4089,N_709,N_1550);
xor U4090 (N_4090,N_168,N_2831);
nor U4091 (N_4091,N_1551,N_682);
nand U4092 (N_4092,N_1672,N_165);
and U4093 (N_4093,N_50,N_2294);
and U4094 (N_4094,N_1507,N_765);
nand U4095 (N_4095,N_986,N_389);
nand U4096 (N_4096,N_595,N_2981);
or U4097 (N_4097,N_2987,N_2777);
xnor U4098 (N_4098,N_339,N_101);
or U4099 (N_4099,N_1865,N_252);
xnor U4100 (N_4100,N_1737,N_2440);
nor U4101 (N_4101,N_954,N_2475);
and U4102 (N_4102,N_1104,N_463);
nor U4103 (N_4103,N_1868,N_759);
and U4104 (N_4104,N_2679,N_2205);
xnor U4105 (N_4105,N_1071,N_816);
or U4106 (N_4106,N_342,N_2767);
or U4107 (N_4107,N_1693,N_968);
nand U4108 (N_4108,N_2044,N_549);
or U4109 (N_4109,N_2417,N_3035);
nand U4110 (N_4110,N_353,N_1722);
xor U4111 (N_4111,N_518,N_1733);
nand U4112 (N_4112,N_1247,N_397);
nor U4113 (N_4113,N_2046,N_2302);
xor U4114 (N_4114,N_2021,N_3096);
nand U4115 (N_4115,N_2643,N_1131);
xor U4116 (N_4116,N_2790,N_629);
or U4117 (N_4117,N_2826,N_286);
nor U4118 (N_4118,N_1060,N_1476);
nor U4119 (N_4119,N_2376,N_2756);
xnor U4120 (N_4120,N_2793,N_1492);
nor U4121 (N_4121,N_127,N_2221);
nor U4122 (N_4122,N_681,N_983);
and U4123 (N_4123,N_3062,N_394);
nor U4124 (N_4124,N_2000,N_1035);
xnor U4125 (N_4125,N_1742,N_665);
nand U4126 (N_4126,N_2318,N_2732);
nor U4127 (N_4127,N_77,N_1675);
nand U4128 (N_4128,N_2030,N_1004);
or U4129 (N_4129,N_2329,N_2363);
nor U4130 (N_4130,N_479,N_2751);
or U4131 (N_4131,N_2367,N_1335);
nand U4132 (N_4132,N_1383,N_1593);
and U4133 (N_4133,N_996,N_1527);
or U4134 (N_4134,N_94,N_1844);
nor U4135 (N_4135,N_1612,N_563);
xor U4136 (N_4136,N_410,N_2994);
xor U4137 (N_4137,N_916,N_3081);
and U4138 (N_4138,N_3061,N_1487);
xor U4139 (N_4139,N_839,N_914);
nor U4140 (N_4140,N_2659,N_1144);
xnor U4141 (N_4141,N_2335,N_1212);
and U4142 (N_4142,N_1882,N_1748);
nand U4143 (N_4143,N_746,N_1242);
or U4144 (N_4144,N_2482,N_258);
xnor U4145 (N_4145,N_2488,N_2120);
or U4146 (N_4146,N_2948,N_1799);
nor U4147 (N_4147,N_2669,N_814);
nor U4148 (N_4148,N_90,N_386);
or U4149 (N_4149,N_5,N_1075);
or U4150 (N_4150,N_1184,N_2242);
nand U4151 (N_4151,N_2125,N_196);
and U4152 (N_4152,N_2676,N_2397);
or U4153 (N_4153,N_64,N_993);
and U4154 (N_4154,N_2328,N_3026);
xor U4155 (N_4155,N_1883,N_1547);
nand U4156 (N_4156,N_1712,N_322);
nand U4157 (N_4157,N_1412,N_1446);
xnor U4158 (N_4158,N_333,N_957);
or U4159 (N_4159,N_182,N_1934);
xor U4160 (N_4160,N_2405,N_1545);
nor U4161 (N_4161,N_1621,N_3092);
nor U4162 (N_4162,N_447,N_873);
and U4163 (N_4163,N_417,N_1034);
or U4164 (N_4164,N_1120,N_1010);
nand U4165 (N_4165,N_2748,N_2832);
nand U4166 (N_4166,N_2538,N_1569);
nor U4167 (N_4167,N_1519,N_95);
nand U4168 (N_4168,N_314,N_2792);
or U4169 (N_4169,N_75,N_3010);
xnor U4170 (N_4170,N_1645,N_584);
nor U4171 (N_4171,N_364,N_2633);
xnor U4172 (N_4172,N_2274,N_2736);
nand U4173 (N_4173,N_1623,N_751);
nor U4174 (N_4174,N_1310,N_589);
and U4175 (N_4175,N_2974,N_927);
xor U4176 (N_4176,N_2145,N_2827);
nor U4177 (N_4177,N_841,N_2495);
nor U4178 (N_4178,N_764,N_1426);
xor U4179 (N_4179,N_1101,N_699);
xor U4180 (N_4180,N_2901,N_825);
nor U4181 (N_4181,N_381,N_2388);
or U4182 (N_4182,N_3033,N_1603);
nand U4183 (N_4183,N_2375,N_3009);
and U4184 (N_4184,N_2809,N_725);
or U4185 (N_4185,N_2411,N_49);
nor U4186 (N_4186,N_1754,N_2404);
or U4187 (N_4187,N_429,N_672);
xor U4188 (N_4188,N_3057,N_2313);
nor U4189 (N_4189,N_3056,N_141);
and U4190 (N_4190,N_2584,N_650);
xnor U4191 (N_4191,N_1600,N_2052);
nand U4192 (N_4192,N_6,N_304);
and U4193 (N_4193,N_1241,N_2817);
nand U4194 (N_4194,N_2100,N_880);
xnor U4195 (N_4195,N_801,N_811);
nor U4196 (N_4196,N_1089,N_2208);
nand U4197 (N_4197,N_1056,N_2468);
nand U4198 (N_4198,N_2235,N_2);
xnor U4199 (N_4199,N_2646,N_2895);
nand U4200 (N_4200,N_185,N_1014);
nand U4201 (N_4201,N_57,N_3013);
nand U4202 (N_4202,N_2684,N_1008);
nand U4203 (N_4203,N_1917,N_2701);
nand U4204 (N_4204,N_2609,N_3075);
and U4205 (N_4205,N_2192,N_1815);
or U4206 (N_4206,N_2080,N_2964);
nand U4207 (N_4207,N_797,N_1641);
or U4208 (N_4208,N_1930,N_1048);
nand U4209 (N_4209,N_1948,N_1068);
nor U4210 (N_4210,N_543,N_1542);
nor U4211 (N_4211,N_1983,N_1573);
or U4212 (N_4212,N_622,N_1993);
nand U4213 (N_4213,N_877,N_2604);
nand U4214 (N_4214,N_2344,N_1039);
or U4215 (N_4215,N_2991,N_1664);
and U4216 (N_4216,N_1278,N_1325);
nand U4217 (N_4217,N_3097,N_26);
and U4218 (N_4218,N_2835,N_87);
or U4219 (N_4219,N_1092,N_3124);
and U4220 (N_4220,N_2983,N_1061);
nor U4221 (N_4221,N_2322,N_657);
or U4222 (N_4222,N_2392,N_1009);
xnor U4223 (N_4223,N_2167,N_2925);
xnor U4224 (N_4224,N_826,N_1042);
and U4225 (N_4225,N_2638,N_2735);
nor U4226 (N_4226,N_2258,N_646);
nand U4227 (N_4227,N_2616,N_655);
nor U4228 (N_4228,N_1374,N_777);
and U4229 (N_4229,N_1515,N_2256);
or U4230 (N_4230,N_1802,N_909);
nor U4231 (N_4231,N_2909,N_1410);
and U4232 (N_4232,N_44,N_670);
xnor U4233 (N_4233,N_2859,N_2963);
and U4234 (N_4234,N_326,N_1801);
xnor U4235 (N_4235,N_2263,N_792);
and U4236 (N_4236,N_2954,N_2023);
xnor U4237 (N_4237,N_351,N_2233);
xnor U4238 (N_4238,N_2965,N_2824);
nand U4239 (N_4239,N_449,N_2188);
nand U4240 (N_4240,N_747,N_2611);
xor U4241 (N_4241,N_2799,N_373);
nor U4242 (N_4242,N_1207,N_452);
nor U4243 (N_4243,N_1337,N_934);
and U4244 (N_4244,N_2579,N_2103);
or U4245 (N_4245,N_1220,N_997);
xor U4246 (N_4246,N_732,N_2026);
and U4247 (N_4247,N_804,N_2966);
nor U4248 (N_4248,N_2725,N_562);
and U4249 (N_4249,N_1211,N_56);
xor U4250 (N_4250,N_1640,N_2563);
nor U4251 (N_4251,N_1400,N_2308);
nor U4252 (N_4252,N_2493,N_1710);
and U4253 (N_4253,N_586,N_2425);
nand U4254 (N_4254,N_2150,N_536);
or U4255 (N_4255,N_10,N_3090);
or U4256 (N_4256,N_1185,N_653);
or U4257 (N_4257,N_1450,N_1007);
or U4258 (N_4258,N_211,N_2319);
nor U4259 (N_4259,N_2946,N_1289);
and U4260 (N_4260,N_1628,N_503);
or U4261 (N_4261,N_1544,N_527);
or U4262 (N_4262,N_1952,N_1168);
xnor U4263 (N_4263,N_1058,N_729);
xnor U4264 (N_4264,N_1707,N_533);
or U4265 (N_4265,N_1991,N_2136);
and U4266 (N_4266,N_2851,N_1181);
and U4267 (N_4267,N_47,N_292);
xor U4268 (N_4268,N_455,N_1792);
xnor U4269 (N_4269,N_878,N_2049);
or U4270 (N_4270,N_2556,N_2098);
nand U4271 (N_4271,N_3022,N_2606);
nand U4272 (N_4272,N_1183,N_1839);
or U4273 (N_4273,N_1632,N_1691);
xor U4274 (N_4274,N_519,N_1637);
nor U4275 (N_4275,N_2641,N_2902);
and U4276 (N_4276,N_1262,N_128);
nand U4277 (N_4277,N_1202,N_303);
xnor U4278 (N_4278,N_2169,N_1750);
and U4279 (N_4279,N_2360,N_438);
and U4280 (N_4280,N_638,N_2528);
nand U4281 (N_4281,N_1082,N_1954);
and U4282 (N_4282,N_0,N_120);
nand U4283 (N_4283,N_806,N_2003);
nor U4284 (N_4284,N_1927,N_80);
and U4285 (N_4285,N_3030,N_2975);
nand U4286 (N_4286,N_1482,N_587);
nand U4287 (N_4287,N_1478,N_1789);
xnor U4288 (N_4288,N_1583,N_1333);
or U4289 (N_4289,N_2084,N_2693);
or U4290 (N_4290,N_2504,N_506);
xor U4291 (N_4291,N_951,N_1813);
or U4292 (N_4292,N_2292,N_281);
xor U4293 (N_4293,N_65,N_538);
nor U4294 (N_4294,N_1797,N_2097);
nor U4295 (N_4295,N_1911,N_1874);
nand U4296 (N_4296,N_1037,N_2210);
nor U4297 (N_4297,N_1022,N_24);
xor U4298 (N_4298,N_2710,N_676);
nand U4299 (N_4299,N_1417,N_20);
nor U4300 (N_4300,N_1971,N_2980);
xor U4301 (N_4301,N_2211,N_2138);
nor U4302 (N_4302,N_2371,N_243);
xnor U4303 (N_4303,N_1775,N_183);
nand U4304 (N_4304,N_2443,N_1295);
nor U4305 (N_4305,N_1860,N_2346);
or U4306 (N_4306,N_1931,N_3116);
nand U4307 (N_4307,N_162,N_1132);
nor U4308 (N_4308,N_1568,N_1459);
xnor U4309 (N_4309,N_1532,N_2922);
nand U4310 (N_4310,N_575,N_2362);
nor U4311 (N_4311,N_2309,N_2794);
nor U4312 (N_4312,N_3063,N_2585);
xnor U4313 (N_4313,N_1274,N_2663);
or U4314 (N_4314,N_1141,N_1444);
nor U4315 (N_4315,N_2293,N_1228);
and U4316 (N_4316,N_3005,N_2035);
nor U4317 (N_4317,N_559,N_334);
and U4318 (N_4318,N_1430,N_1352);
nand U4319 (N_4319,N_1070,N_1746);
nand U4320 (N_4320,N_1861,N_444);
xor U4321 (N_4321,N_2476,N_2510);
nand U4322 (N_4322,N_661,N_2600);
and U4323 (N_4323,N_2941,N_1566);
nor U4324 (N_4324,N_2553,N_810);
and U4325 (N_4325,N_248,N_2214);
xnor U4326 (N_4326,N_329,N_1962);
or U4327 (N_4327,N_1052,N_76);
nor U4328 (N_4328,N_2033,N_2842);
xnor U4329 (N_4329,N_2939,N_2164);
and U4330 (N_4330,N_1066,N_330);
and U4331 (N_4331,N_766,N_1208);
or U4332 (N_4332,N_53,N_1887);
and U4333 (N_4333,N_2949,N_1823);
and U4334 (N_4334,N_974,N_919);
xnor U4335 (N_4335,N_2074,N_1083);
and U4336 (N_4336,N_2728,N_1915);
or U4337 (N_4337,N_817,N_2204);
xor U4338 (N_4338,N_2369,N_2699);
and U4339 (N_4339,N_104,N_593);
nand U4340 (N_4340,N_2564,N_420);
and U4341 (N_4341,N_2667,N_1697);
nor U4342 (N_4342,N_1660,N_195);
nand U4343 (N_4343,N_2385,N_425);
or U4344 (N_4344,N_2398,N_2070);
nor U4345 (N_4345,N_1870,N_2193);
nand U4346 (N_4346,N_491,N_2778);
or U4347 (N_4347,N_2422,N_1044);
nand U4348 (N_4348,N_1647,N_2133);
or U4349 (N_4349,N_150,N_1667);
nor U4350 (N_4350,N_2924,N_1128);
xnor U4351 (N_4351,N_17,N_2848);
or U4352 (N_4352,N_1171,N_1677);
nor U4353 (N_4353,N_2059,N_363);
and U4354 (N_4354,N_2031,N_900);
or U4355 (N_4355,N_2160,N_1276);
and U4356 (N_4356,N_2877,N_1319);
or U4357 (N_4357,N_1512,N_498);
nand U4358 (N_4358,N_253,N_337);
or U4359 (N_4359,N_2694,N_857);
nor U4360 (N_4360,N_2862,N_658);
and U4361 (N_4361,N_2950,N_298);
and U4362 (N_4362,N_924,N_2010);
or U4363 (N_4363,N_1761,N_1002);
nand U4364 (N_4364,N_414,N_412);
and U4365 (N_4365,N_2722,N_1439);
and U4366 (N_4366,N_3018,N_2840);
nor U4367 (N_4367,N_2990,N_443);
and U4368 (N_4368,N_2500,N_3003);
and U4369 (N_4369,N_2705,N_551);
xor U4370 (N_4370,N_2249,N_366);
nor U4371 (N_4371,N_91,N_1654);
and U4372 (N_4372,N_2995,N_796);
nand U4373 (N_4373,N_2414,N_1146);
nor U4374 (N_4374,N_1062,N_1025);
or U4375 (N_4375,N_987,N_852);
and U4376 (N_4376,N_1175,N_3045);
xnor U4377 (N_4377,N_3080,N_2680);
nor U4378 (N_4378,N_2303,N_3042);
nor U4379 (N_4379,N_1535,N_2612);
or U4380 (N_4380,N_1087,N_1595);
nor U4381 (N_4381,N_1013,N_2248);
or U4382 (N_4382,N_2113,N_2875);
nor U4383 (N_4383,N_1582,N_399);
and U4384 (N_4384,N_1452,N_921);
xnor U4385 (N_4385,N_2956,N_2264);
xnor U4386 (N_4386,N_2883,N_2195);
or U4387 (N_4387,N_2275,N_2066);
or U4388 (N_4388,N_1509,N_3012);
or U4389 (N_4389,N_879,N_2858);
xnor U4390 (N_4390,N_1808,N_2334);
xnor U4391 (N_4391,N_1334,N_1040);
xnor U4392 (N_4392,N_1498,N_482);
and U4393 (N_4393,N_662,N_1328);
and U4394 (N_4394,N_2786,N_1521);
or U4395 (N_4395,N_123,N_1080);
nand U4396 (N_4396,N_2626,N_1875);
nand U4397 (N_4397,N_487,N_3041);
and U4398 (N_4398,N_88,N_379);
xnor U4399 (N_4399,N_1227,N_249);
nand U4400 (N_4400,N_767,N_616);
xor U4401 (N_4401,N_1606,N_1752);
and U4402 (N_4402,N_146,N_2081);
nor U4403 (N_4403,N_1756,N_697);
nor U4404 (N_4404,N_862,N_1630);
nor U4405 (N_4405,N_2447,N_609);
nor U4406 (N_4406,N_1471,N_911);
nand U4407 (N_4407,N_1301,N_946);
nor U4408 (N_4408,N_2808,N_904);
nor U4409 (N_4409,N_978,N_918);
nand U4410 (N_4410,N_508,N_2804);
xor U4411 (N_4411,N_1302,N_3102);
and U4412 (N_4412,N_1704,N_2278);
nor U4413 (N_4413,N_2396,N_546);
and U4414 (N_4414,N_175,N_2934);
xor U4415 (N_4415,N_2337,N_550);
xor U4416 (N_4416,N_1960,N_1118);
xnor U4417 (N_4417,N_1021,N_2459);
nor U4418 (N_4418,N_1265,N_1373);
nor U4419 (N_4419,N_1543,N_2421);
or U4420 (N_4420,N_1409,N_1910);
and U4421 (N_4421,N_2262,N_2115);
or U4422 (N_4422,N_360,N_1157);
nand U4423 (N_4423,N_703,N_548);
or U4424 (N_4424,N_952,N_712);
xnor U4425 (N_4425,N_1314,N_3104);
or U4426 (N_4426,N_789,N_310);
nor U4427 (N_4427,N_140,N_511);
nand U4428 (N_4428,N_1491,N_2341);
and U4429 (N_4429,N_407,N_875);
and U4430 (N_4430,N_1119,N_2557);
or U4431 (N_4431,N_544,N_313);
nand U4432 (N_4432,N_1327,N_2936);
and U4433 (N_4433,N_1453,N_1307);
or U4434 (N_4434,N_727,N_1113);
xor U4435 (N_4435,N_1231,N_52);
xnor U4436 (N_4436,N_1810,N_1210);
nand U4437 (N_4437,N_1229,N_418);
and U4438 (N_4438,N_3091,N_234);
nand U4439 (N_4439,N_1005,N_726);
nor U4440 (N_4440,N_2913,N_1406);
nand U4441 (N_4441,N_1649,N_1299);
nor U4442 (N_4442,N_2429,N_1269);
or U4443 (N_4443,N_2619,N_835);
nand U4444 (N_4444,N_710,N_637);
and U4445 (N_4445,N_891,N_2124);
or U4446 (N_4446,N_240,N_608);
nor U4447 (N_4447,N_2812,N_625);
and U4448 (N_4448,N_1318,N_567);
nand U4449 (N_4449,N_388,N_2550);
or U4450 (N_4450,N_886,N_1997);
xnor U4451 (N_4451,N_2383,N_724);
nor U4452 (N_4452,N_1425,N_2243);
xor U4453 (N_4453,N_2018,N_2614);
and U4454 (N_4454,N_1554,N_605);
xor U4455 (N_4455,N_2665,N_29);
and U4456 (N_4456,N_2757,N_1028);
or U4457 (N_4457,N_473,N_1465);
xnor U4458 (N_4458,N_2654,N_1050);
or U4459 (N_4459,N_3074,N_2586);
nor U4460 (N_4460,N_743,N_336);
xnor U4461 (N_4461,N_639,N_1820);
or U4462 (N_4462,N_15,N_2306);
nor U4463 (N_4463,N_1418,N_2483);
and U4464 (N_4464,N_752,N_2343);
nor U4465 (N_4465,N_86,N_117);
or U4466 (N_4466,N_819,N_1283);
nor U4467 (N_4467,N_2489,N_2914);
xnor U4468 (N_4468,N_2355,N_1786);
or U4469 (N_4469,N_2194,N_935);
nand U4470 (N_4470,N_1348,N_565);
and U4471 (N_4471,N_1429,N_2148);
or U4472 (N_4472,N_1853,N_2047);
and U4473 (N_4473,N_1986,N_1045);
nand U4474 (N_4474,N_3037,N_647);
nor U4475 (N_4475,N_1399,N_2350);
and U4476 (N_4476,N_910,N_2289);
nor U4477 (N_4477,N_773,N_436);
and U4478 (N_4478,N_1557,N_1905);
nor U4479 (N_4479,N_882,N_1831);
and U4480 (N_4480,N_795,N_1766);
or U4481 (N_4481,N_106,N_2314);
xnor U4482 (N_4482,N_392,N_2927);
or U4483 (N_4483,N_620,N_2416);
or U4484 (N_4484,N_3043,N_2886);
nor U4485 (N_4485,N_1015,N_2265);
nor U4486 (N_4486,N_2591,N_2458);
nand U4487 (N_4487,N_1148,N_1828);
nand U4488 (N_4488,N_108,N_116);
nor U4489 (N_4489,N_944,N_2755);
xnor U4490 (N_4490,N_837,N_2281);
or U4491 (N_4491,N_1926,N_2593);
or U4492 (N_4492,N_2668,N_828);
and U4493 (N_4493,N_939,N_406);
and U4494 (N_4494,N_1920,N_1494);
or U4495 (N_4495,N_991,N_144);
xnor U4496 (N_4496,N_1706,N_2140);
xnor U4497 (N_4497,N_698,N_706);
nand U4498 (N_4498,N_1814,N_1904);
or U4499 (N_4499,N_4,N_1715);
or U4500 (N_4500,N_2220,N_1721);
or U4501 (N_4501,N_1884,N_2496);
nand U4502 (N_4502,N_474,N_2087);
nor U4503 (N_4503,N_2041,N_779);
xnor U4504 (N_4504,N_716,N_1942);
xor U4505 (N_4505,N_2064,N_192);
xnor U4506 (N_4506,N_1900,N_2758);
xor U4507 (N_4507,N_975,N_1951);
or U4508 (N_4508,N_1000,N_1656);
xnor U4509 (N_4509,N_1054,N_1388);
and U4510 (N_4510,N_2629,N_2741);
nor U4511 (N_4511,N_995,N_345);
nand U4512 (N_4512,N_768,N_541);
or U4513 (N_4513,N_1447,N_2179);
nor U4514 (N_4514,N_2312,N_416);
nor U4515 (N_4515,N_1788,N_1279);
and U4516 (N_4516,N_277,N_485);
nand U4517 (N_4517,N_1077,N_1835);
and U4518 (N_4518,N_2317,N_1723);
and U4519 (N_4519,N_161,N_2290);
or U4520 (N_4520,N_530,N_2251);
xnor U4521 (N_4521,N_2288,N_2002);
nand U4522 (N_4522,N_1537,N_2339);
and U4523 (N_4523,N_2452,N_2796);
or U4524 (N_4524,N_1386,N_2765);
or U4525 (N_4525,N_1296,N_800);
nor U4526 (N_4526,N_1800,N_1558);
nor U4527 (N_4527,N_448,N_1480);
and U4528 (N_4528,N_223,N_640);
nand U4529 (N_4529,N_164,N_2234);
nor U4530 (N_4530,N_2889,N_2683);
or U4531 (N_4531,N_693,N_2815);
or U4532 (N_4532,N_2250,N_3023);
nor U4533 (N_4533,N_2079,N_1030);
xor U4534 (N_4534,N_1076,N_2259);
nor U4535 (N_4535,N_3110,N_1139);
nor U4536 (N_4536,N_1778,N_2866);
nor U4537 (N_4537,N_576,N_771);
xor U4538 (N_4538,N_610,N_191);
nor U4539 (N_4539,N_1912,N_2558);
or U4540 (N_4540,N_1564,N_2785);
or U4541 (N_4541,N_2130,N_3120);
and U4542 (N_4542,N_528,N_2731);
nor U4543 (N_4543,N_1718,N_2596);
nand U4544 (N_4544,N_2055,N_2656);
xnor U4545 (N_4545,N_25,N_186);
or U4546 (N_4546,N_2763,N_1288);
and U4547 (N_4547,N_1871,N_1329);
and U4548 (N_4548,N_1525,N_2688);
nor U4549 (N_4549,N_950,N_731);
and U4550 (N_4550,N_2764,N_1599);
nand U4551 (N_4551,N_1355,N_2174);
nand U4552 (N_4552,N_883,N_1405);
and U4553 (N_4553,N_226,N_1902);
and U4554 (N_4554,N_174,N_69);
nor U4555 (N_4555,N_1966,N_965);
and U4556 (N_4556,N_903,N_1812);
nor U4557 (N_4557,N_931,N_1099);
nand U4558 (N_4558,N_2228,N_863);
nand U4559 (N_4559,N_920,N_2671);
nor U4560 (N_4560,N_2352,N_1851);
nor U4561 (N_4561,N_1968,N_43);
nand U4562 (N_4562,N_2439,N_2065);
and U4563 (N_4563,N_1901,N_1121);
and U4564 (N_4564,N_1624,N_1548);
xor U4565 (N_4565,N_2420,N_1964);
and U4566 (N_4566,N_2225,N_3068);
or U4567 (N_4567,N_2175,N_2477);
nand U4568 (N_4568,N_1511,N_678);
nand U4569 (N_4569,N_1977,N_1);
nand U4570 (N_4570,N_2147,N_744);
nand U4571 (N_4571,N_788,N_2083);
nand U4572 (N_4572,N_8,N_1437);
and U4573 (N_4573,N_2746,N_1251);
nand U4574 (N_4574,N_1095,N_2813);
xor U4575 (N_4575,N_271,N_2207);
xor U4576 (N_4576,N_809,N_673);
nor U4577 (N_4577,N_222,N_2829);
nand U4578 (N_4578,N_1984,N_2128);
or U4579 (N_4579,N_2013,N_1771);
xnor U4580 (N_4580,N_1368,N_1362);
and U4581 (N_4581,N_1233,N_1967);
or U4582 (N_4582,N_1824,N_1903);
and U4583 (N_4583,N_504,N_1847);
xor U4584 (N_4584,N_2897,N_2628);
or U4585 (N_4585,N_2390,N_467);
or U4586 (N_4586,N_22,N_2399);
nor U4587 (N_4587,N_2331,N_1561);
xor U4588 (N_4588,N_2514,N_468);
nor U4589 (N_4589,N_585,N_2298);
xnor U4590 (N_4590,N_3048,N_793);
or U4591 (N_4591,N_1850,N_881);
and U4592 (N_4592,N_2008,N_3058);
xnor U4593 (N_4593,N_2051,N_2199);
and U4594 (N_4594,N_614,N_2296);
nand U4595 (N_4595,N_537,N_3047);
and U4596 (N_4596,N_188,N_799);
or U4597 (N_4597,N_1165,N_2837);
nor U4598 (N_4598,N_955,N_2545);
nor U4599 (N_4599,N_1199,N_492);
and U4600 (N_4600,N_242,N_1717);
nor U4601 (N_4601,N_798,N_850);
nand U4602 (N_4602,N_2685,N_2032);
xnor U4603 (N_4603,N_524,N_1137);
xor U4604 (N_4604,N_2291,N_1898);
or U4605 (N_4605,N_2672,N_500);
nand U4606 (N_4606,N_842,N_2960);
and U4607 (N_4607,N_2149,N_424);
nor U4608 (N_4608,N_73,N_158);
nor U4609 (N_4609,N_739,N_210);
nand U4610 (N_4610,N_42,N_79);
or U4611 (N_4611,N_1029,N_159);
nand U4612 (N_4612,N_256,N_3044);
xnor U4613 (N_4613,N_2744,N_2014);
nor U4614 (N_4614,N_1317,N_2571);
or U4615 (N_4615,N_1581,N_1510);
nand U4616 (N_4616,N_496,N_2546);
or U4617 (N_4617,N_343,N_285);
or U4618 (N_4618,N_1038,N_78);
nor U4619 (N_4619,N_2156,N_1206);
and U4620 (N_4620,N_261,N_720);
or U4621 (N_4621,N_1735,N_1304);
nor U4622 (N_4622,N_2111,N_1216);
nand U4623 (N_4623,N_2057,N_1496);
nor U4624 (N_4624,N_1152,N_2531);
or U4625 (N_4625,N_1533,N_569);
nand U4626 (N_4626,N_1246,N_46);
and U4627 (N_4627,N_1819,N_402);
or U4628 (N_4628,N_2904,N_1607);
xor U4629 (N_4629,N_972,N_2200);
and U4630 (N_4630,N_821,N_1112);
xor U4631 (N_4631,N_2750,N_2218);
xor U4632 (N_4632,N_3040,N_3007);
nand U4633 (N_4633,N_2845,N_557);
or U4634 (N_4634,N_2450,N_2810);
and U4635 (N_4635,N_469,N_1666);
or U4636 (N_4636,N_1978,N_2716);
nor U4637 (N_4637,N_1506,N_649);
nor U4638 (N_4638,N_441,N_2058);
and U4639 (N_4639,N_2226,N_1483);
xnor U4640 (N_4640,N_3122,N_542);
xor U4641 (N_4641,N_523,N_1085);
xnor U4642 (N_4642,N_2613,N_627);
nor U4643 (N_4643,N_2863,N_2151);
xor U4644 (N_4644,N_1490,N_2239);
xor U4645 (N_4645,N_61,N_477);
or U4646 (N_4646,N_2887,N_906);
nor U4647 (N_4647,N_1703,N_737);
xnor U4648 (N_4648,N_1270,N_1154);
xor U4649 (N_4649,N_1424,N_1709);
nor U4650 (N_4650,N_3088,N_415);
nand U4651 (N_4651,N_687,N_1696);
nand U4652 (N_4652,N_1781,N_1845);
nand U4653 (N_4653,N_323,N_1594);
xnor U4654 (N_4654,N_1467,N_897);
xor U4655 (N_4655,N_1804,N_663);
or U4656 (N_4656,N_2391,N_2984);
and U4657 (N_4657,N_1598,N_1620);
nand U4658 (N_4658,N_1254,N_2856);
nand U4659 (N_4659,N_2881,N_2865);
nor U4660 (N_4660,N_1890,N_1925);
and U4661 (N_4661,N_579,N_2307);
xnor U4662 (N_4662,N_514,N_666);
and U4663 (N_4663,N_748,N_2890);
xnor U4664 (N_4664,N_961,N_1277);
or U4665 (N_4665,N_1674,N_1889);
or U4666 (N_4666,N_2461,N_2415);
nand U4667 (N_4667,N_840,N_522);
nand U4668 (N_4668,N_1587,N_683);
nand U4669 (N_4669,N_1739,N_2089);
xnor U4670 (N_4670,N_335,N_631);
and U4671 (N_4671,N_2903,N_401);
nand U4672 (N_4672,N_959,N_2073);
or U4673 (N_4673,N_170,N_1306);
nor U4674 (N_4674,N_2144,N_2692);
nor U4675 (N_4675,N_1458,N_870);
nor U4676 (N_4676,N_2873,N_16);
or U4677 (N_4677,N_615,N_497);
or U4678 (N_4678,N_2976,N_1435);
nand U4679 (N_4679,N_2931,N_1356);
nor U4680 (N_4680,N_1683,N_1730);
xnor U4681 (N_4681,N_560,N_1538);
xnor U4682 (N_4682,N_2132,N_1036);
nor U4683 (N_4683,N_963,N_433);
nor U4684 (N_4684,N_320,N_2216);
xor U4685 (N_4685,N_135,N_1225);
xor U4686 (N_4686,N_1193,N_884);
nor U4687 (N_4687,N_999,N_2733);
and U4688 (N_4688,N_2349,N_2003);
nand U4689 (N_4689,N_854,N_3081);
and U4690 (N_4690,N_258,N_565);
xnor U4691 (N_4691,N_2218,N_1236);
nor U4692 (N_4692,N_1440,N_3101);
or U4693 (N_4693,N_1037,N_2802);
nand U4694 (N_4694,N_2599,N_126);
or U4695 (N_4695,N_2497,N_1734);
nand U4696 (N_4696,N_1775,N_873);
xnor U4697 (N_4697,N_1755,N_2266);
nor U4698 (N_4698,N_473,N_1185);
nor U4699 (N_4699,N_3023,N_1853);
xnor U4700 (N_4700,N_2060,N_2007);
xor U4701 (N_4701,N_1070,N_664);
or U4702 (N_4702,N_1847,N_2119);
and U4703 (N_4703,N_2673,N_1873);
nor U4704 (N_4704,N_680,N_1733);
nand U4705 (N_4705,N_2432,N_470);
nor U4706 (N_4706,N_2342,N_914);
or U4707 (N_4707,N_1544,N_1880);
nand U4708 (N_4708,N_1603,N_2427);
xnor U4709 (N_4709,N_62,N_982);
or U4710 (N_4710,N_1403,N_473);
and U4711 (N_4711,N_1111,N_2687);
or U4712 (N_4712,N_1579,N_2960);
xnor U4713 (N_4713,N_2063,N_1164);
xnor U4714 (N_4714,N_2346,N_1485);
nor U4715 (N_4715,N_2718,N_863);
nor U4716 (N_4716,N_1479,N_1856);
nor U4717 (N_4717,N_3020,N_2922);
xor U4718 (N_4718,N_1111,N_2458);
nor U4719 (N_4719,N_368,N_184);
and U4720 (N_4720,N_1318,N_1492);
and U4721 (N_4721,N_639,N_2624);
or U4722 (N_4722,N_1270,N_707);
or U4723 (N_4723,N_173,N_977);
xnor U4724 (N_4724,N_1127,N_1153);
nand U4725 (N_4725,N_2273,N_2556);
and U4726 (N_4726,N_350,N_1855);
xnor U4727 (N_4727,N_2767,N_616);
or U4728 (N_4728,N_1625,N_1673);
or U4729 (N_4729,N_632,N_2625);
and U4730 (N_4730,N_632,N_2037);
or U4731 (N_4731,N_2713,N_549);
and U4732 (N_4732,N_2961,N_2520);
and U4733 (N_4733,N_599,N_2310);
nor U4734 (N_4734,N_2086,N_173);
and U4735 (N_4735,N_3072,N_2665);
or U4736 (N_4736,N_1628,N_543);
and U4737 (N_4737,N_743,N_658);
nor U4738 (N_4738,N_508,N_2014);
or U4739 (N_4739,N_1849,N_947);
nand U4740 (N_4740,N_1156,N_62);
or U4741 (N_4741,N_1723,N_498);
xor U4742 (N_4742,N_1840,N_573);
xnor U4743 (N_4743,N_1212,N_2185);
or U4744 (N_4744,N_1423,N_608);
nand U4745 (N_4745,N_2438,N_2437);
and U4746 (N_4746,N_424,N_1153);
and U4747 (N_4747,N_1318,N_793);
xnor U4748 (N_4748,N_2785,N_1596);
xor U4749 (N_4749,N_503,N_355);
and U4750 (N_4750,N_626,N_637);
nand U4751 (N_4751,N_1566,N_3106);
nand U4752 (N_4752,N_2704,N_3047);
and U4753 (N_4753,N_501,N_805);
or U4754 (N_4754,N_1641,N_1342);
nor U4755 (N_4755,N_2706,N_2790);
nand U4756 (N_4756,N_2886,N_1505);
xor U4757 (N_4757,N_3057,N_2207);
xnor U4758 (N_4758,N_3040,N_662);
xor U4759 (N_4759,N_747,N_2700);
or U4760 (N_4760,N_2957,N_979);
or U4761 (N_4761,N_1159,N_1496);
and U4762 (N_4762,N_2954,N_1529);
nand U4763 (N_4763,N_825,N_3048);
nand U4764 (N_4764,N_786,N_1278);
nand U4765 (N_4765,N_256,N_426);
and U4766 (N_4766,N_1667,N_2154);
and U4767 (N_4767,N_1518,N_3061);
and U4768 (N_4768,N_1201,N_418);
and U4769 (N_4769,N_713,N_636);
xor U4770 (N_4770,N_552,N_970);
nor U4771 (N_4771,N_1278,N_219);
and U4772 (N_4772,N_2933,N_2104);
nor U4773 (N_4773,N_1647,N_783);
or U4774 (N_4774,N_679,N_1664);
xor U4775 (N_4775,N_715,N_782);
nand U4776 (N_4776,N_1099,N_3042);
or U4777 (N_4777,N_677,N_1351);
nor U4778 (N_4778,N_1061,N_1650);
nor U4779 (N_4779,N_114,N_2455);
xnor U4780 (N_4780,N_1186,N_916);
nand U4781 (N_4781,N_833,N_2224);
or U4782 (N_4782,N_1317,N_279);
and U4783 (N_4783,N_606,N_2631);
xor U4784 (N_4784,N_1916,N_1182);
or U4785 (N_4785,N_1130,N_2405);
nor U4786 (N_4786,N_603,N_3037);
nor U4787 (N_4787,N_1262,N_1581);
and U4788 (N_4788,N_907,N_1134);
or U4789 (N_4789,N_2353,N_1678);
nand U4790 (N_4790,N_1427,N_651);
and U4791 (N_4791,N_2126,N_1240);
and U4792 (N_4792,N_1182,N_2019);
and U4793 (N_4793,N_789,N_805);
xor U4794 (N_4794,N_123,N_657);
nor U4795 (N_4795,N_45,N_1191);
or U4796 (N_4796,N_1968,N_1434);
or U4797 (N_4797,N_19,N_1025);
and U4798 (N_4798,N_2980,N_2411);
xor U4799 (N_4799,N_911,N_1327);
nor U4800 (N_4800,N_2462,N_793);
xor U4801 (N_4801,N_2591,N_1368);
and U4802 (N_4802,N_1803,N_1539);
nand U4803 (N_4803,N_1508,N_1815);
nand U4804 (N_4804,N_665,N_740);
and U4805 (N_4805,N_1880,N_606);
and U4806 (N_4806,N_1655,N_789);
nor U4807 (N_4807,N_1510,N_157);
or U4808 (N_4808,N_2533,N_2434);
and U4809 (N_4809,N_2153,N_1133);
and U4810 (N_4810,N_478,N_2912);
xnor U4811 (N_4811,N_1035,N_2674);
nand U4812 (N_4812,N_717,N_2129);
nor U4813 (N_4813,N_2188,N_2703);
and U4814 (N_4814,N_590,N_1002);
and U4815 (N_4815,N_2307,N_572);
or U4816 (N_4816,N_880,N_294);
nor U4817 (N_4817,N_2016,N_1946);
nor U4818 (N_4818,N_3010,N_2751);
nor U4819 (N_4819,N_2658,N_141);
xor U4820 (N_4820,N_41,N_1280);
or U4821 (N_4821,N_3065,N_3087);
or U4822 (N_4822,N_462,N_188);
nor U4823 (N_4823,N_246,N_2031);
nor U4824 (N_4824,N_1722,N_2295);
and U4825 (N_4825,N_2917,N_966);
nor U4826 (N_4826,N_1114,N_760);
and U4827 (N_4827,N_1874,N_181);
xor U4828 (N_4828,N_967,N_998);
and U4829 (N_4829,N_2369,N_622);
or U4830 (N_4830,N_1946,N_2348);
and U4831 (N_4831,N_2283,N_98);
or U4832 (N_4832,N_3008,N_2726);
nor U4833 (N_4833,N_496,N_504);
xor U4834 (N_4834,N_44,N_269);
or U4835 (N_4835,N_861,N_1);
xnor U4836 (N_4836,N_2763,N_2031);
and U4837 (N_4837,N_485,N_2108);
xor U4838 (N_4838,N_2185,N_1509);
or U4839 (N_4839,N_946,N_240);
and U4840 (N_4840,N_986,N_1840);
nor U4841 (N_4841,N_325,N_1562);
xnor U4842 (N_4842,N_2970,N_1315);
nor U4843 (N_4843,N_1579,N_60);
and U4844 (N_4844,N_1763,N_2625);
nand U4845 (N_4845,N_2721,N_1152);
nand U4846 (N_4846,N_329,N_1054);
or U4847 (N_4847,N_3109,N_272);
or U4848 (N_4848,N_1266,N_771);
nand U4849 (N_4849,N_144,N_2207);
or U4850 (N_4850,N_2136,N_568);
xor U4851 (N_4851,N_627,N_1744);
and U4852 (N_4852,N_3027,N_520);
nand U4853 (N_4853,N_2940,N_1319);
nand U4854 (N_4854,N_2874,N_1227);
nor U4855 (N_4855,N_1150,N_2036);
xor U4856 (N_4856,N_2296,N_1304);
nand U4857 (N_4857,N_1287,N_640);
nor U4858 (N_4858,N_1676,N_1987);
xor U4859 (N_4859,N_364,N_455);
nor U4860 (N_4860,N_388,N_1469);
nor U4861 (N_4861,N_462,N_897);
xnor U4862 (N_4862,N_2733,N_714);
nand U4863 (N_4863,N_106,N_1917);
and U4864 (N_4864,N_678,N_1429);
nand U4865 (N_4865,N_2421,N_249);
nor U4866 (N_4866,N_1185,N_301);
and U4867 (N_4867,N_42,N_593);
or U4868 (N_4868,N_2491,N_2725);
xor U4869 (N_4869,N_302,N_1610);
and U4870 (N_4870,N_475,N_1838);
and U4871 (N_4871,N_1838,N_751);
or U4872 (N_4872,N_1254,N_1502);
or U4873 (N_4873,N_2437,N_81);
nor U4874 (N_4874,N_2246,N_1120);
or U4875 (N_4875,N_2417,N_1424);
nand U4876 (N_4876,N_1044,N_1495);
nand U4877 (N_4877,N_2787,N_2586);
and U4878 (N_4878,N_2041,N_2473);
or U4879 (N_4879,N_1482,N_158);
nand U4880 (N_4880,N_1954,N_2460);
nand U4881 (N_4881,N_1732,N_413);
nor U4882 (N_4882,N_2484,N_2146);
nand U4883 (N_4883,N_2076,N_2760);
or U4884 (N_4884,N_270,N_330);
nand U4885 (N_4885,N_2475,N_2470);
xor U4886 (N_4886,N_2857,N_2836);
and U4887 (N_4887,N_2479,N_460);
or U4888 (N_4888,N_2279,N_2153);
xor U4889 (N_4889,N_655,N_1676);
xnor U4890 (N_4890,N_1744,N_1441);
nor U4891 (N_4891,N_1139,N_2796);
nor U4892 (N_4892,N_1150,N_163);
or U4893 (N_4893,N_2471,N_1231);
or U4894 (N_4894,N_3004,N_2113);
nor U4895 (N_4895,N_1690,N_956);
nor U4896 (N_4896,N_1080,N_1450);
or U4897 (N_4897,N_25,N_977);
nand U4898 (N_4898,N_2940,N_1751);
or U4899 (N_4899,N_2048,N_2378);
or U4900 (N_4900,N_1967,N_177);
xnor U4901 (N_4901,N_1868,N_1803);
nor U4902 (N_4902,N_1180,N_703);
nand U4903 (N_4903,N_1839,N_669);
or U4904 (N_4904,N_1915,N_889);
and U4905 (N_4905,N_1341,N_2431);
and U4906 (N_4906,N_898,N_1074);
nor U4907 (N_4907,N_2777,N_688);
and U4908 (N_4908,N_793,N_902);
and U4909 (N_4909,N_402,N_458);
xnor U4910 (N_4910,N_458,N_650);
or U4911 (N_4911,N_1411,N_138);
or U4912 (N_4912,N_1707,N_3035);
and U4913 (N_4913,N_2566,N_275);
xnor U4914 (N_4914,N_1517,N_2664);
xnor U4915 (N_4915,N_699,N_1057);
or U4916 (N_4916,N_2235,N_2012);
nor U4917 (N_4917,N_701,N_1457);
nand U4918 (N_4918,N_524,N_1767);
or U4919 (N_4919,N_2546,N_991);
nand U4920 (N_4920,N_2254,N_355);
and U4921 (N_4921,N_210,N_1598);
xor U4922 (N_4922,N_2542,N_2105);
nor U4923 (N_4923,N_1227,N_984);
xor U4924 (N_4924,N_2445,N_352);
nand U4925 (N_4925,N_2219,N_2222);
xor U4926 (N_4926,N_2665,N_954);
nor U4927 (N_4927,N_1308,N_2157);
xor U4928 (N_4928,N_789,N_1538);
and U4929 (N_4929,N_1961,N_1318);
xnor U4930 (N_4930,N_2377,N_877);
xnor U4931 (N_4931,N_1402,N_2742);
and U4932 (N_4932,N_124,N_1625);
nand U4933 (N_4933,N_674,N_3082);
and U4934 (N_4934,N_2815,N_2559);
xor U4935 (N_4935,N_986,N_3077);
nor U4936 (N_4936,N_1824,N_104);
or U4937 (N_4937,N_2600,N_2616);
and U4938 (N_4938,N_685,N_1793);
nor U4939 (N_4939,N_2716,N_2678);
nand U4940 (N_4940,N_908,N_171);
xor U4941 (N_4941,N_3051,N_998);
xnor U4942 (N_4942,N_351,N_1690);
or U4943 (N_4943,N_1872,N_3050);
nand U4944 (N_4944,N_689,N_266);
xnor U4945 (N_4945,N_1583,N_1426);
nor U4946 (N_4946,N_2683,N_3036);
nand U4947 (N_4947,N_1268,N_1991);
xnor U4948 (N_4948,N_2618,N_252);
and U4949 (N_4949,N_1403,N_2179);
and U4950 (N_4950,N_2169,N_1909);
and U4951 (N_4951,N_1118,N_556);
and U4952 (N_4952,N_1793,N_467);
xor U4953 (N_4953,N_1756,N_1472);
or U4954 (N_4954,N_1750,N_1519);
xor U4955 (N_4955,N_2828,N_2086);
or U4956 (N_4956,N_2366,N_1754);
and U4957 (N_4957,N_2455,N_2582);
and U4958 (N_4958,N_3004,N_1078);
nor U4959 (N_4959,N_564,N_2911);
xnor U4960 (N_4960,N_2338,N_1653);
nand U4961 (N_4961,N_916,N_221);
xnor U4962 (N_4962,N_2193,N_685);
nor U4963 (N_4963,N_2889,N_2163);
and U4964 (N_4964,N_1792,N_3120);
xnor U4965 (N_4965,N_2113,N_2247);
nand U4966 (N_4966,N_2265,N_357);
or U4967 (N_4967,N_2493,N_1134);
nor U4968 (N_4968,N_2189,N_2895);
xnor U4969 (N_4969,N_2627,N_1641);
nor U4970 (N_4970,N_2688,N_2155);
nand U4971 (N_4971,N_541,N_2960);
nand U4972 (N_4972,N_1669,N_52);
nor U4973 (N_4973,N_36,N_1735);
or U4974 (N_4974,N_2707,N_460);
or U4975 (N_4975,N_2840,N_767);
or U4976 (N_4976,N_713,N_2686);
xnor U4977 (N_4977,N_1403,N_1006);
and U4978 (N_4978,N_1011,N_1058);
nand U4979 (N_4979,N_2927,N_735);
nand U4980 (N_4980,N_2288,N_1682);
nor U4981 (N_4981,N_1809,N_529);
or U4982 (N_4982,N_2352,N_394);
xor U4983 (N_4983,N_252,N_238);
nand U4984 (N_4984,N_1830,N_1859);
nor U4985 (N_4985,N_1829,N_1968);
or U4986 (N_4986,N_743,N_2603);
or U4987 (N_4987,N_970,N_191);
xor U4988 (N_4988,N_2412,N_465);
xor U4989 (N_4989,N_2418,N_901);
or U4990 (N_4990,N_1898,N_2474);
and U4991 (N_4991,N_2937,N_1659);
nand U4992 (N_4992,N_3118,N_4);
xor U4993 (N_4993,N_2070,N_1865);
nor U4994 (N_4994,N_1456,N_1520);
nor U4995 (N_4995,N_1376,N_1438);
xor U4996 (N_4996,N_368,N_1139);
and U4997 (N_4997,N_123,N_3055);
xnor U4998 (N_4998,N_1419,N_1690);
or U4999 (N_4999,N_1576,N_2886);
xor U5000 (N_5000,N_2068,N_2409);
and U5001 (N_5001,N_2010,N_59);
and U5002 (N_5002,N_2955,N_549);
nor U5003 (N_5003,N_836,N_438);
nand U5004 (N_5004,N_2011,N_1363);
nand U5005 (N_5005,N_1191,N_1581);
xnor U5006 (N_5006,N_2946,N_422);
nand U5007 (N_5007,N_526,N_1904);
xor U5008 (N_5008,N_1333,N_2873);
and U5009 (N_5009,N_805,N_2815);
xor U5010 (N_5010,N_421,N_2105);
nand U5011 (N_5011,N_2122,N_2180);
nand U5012 (N_5012,N_754,N_2933);
or U5013 (N_5013,N_2263,N_3016);
and U5014 (N_5014,N_2769,N_883);
xnor U5015 (N_5015,N_1003,N_1107);
or U5016 (N_5016,N_914,N_940);
nand U5017 (N_5017,N_1354,N_146);
and U5018 (N_5018,N_1231,N_1558);
nor U5019 (N_5019,N_2562,N_322);
and U5020 (N_5020,N_1539,N_570);
and U5021 (N_5021,N_2806,N_2690);
nor U5022 (N_5022,N_42,N_1257);
or U5023 (N_5023,N_1123,N_49);
or U5024 (N_5024,N_1097,N_169);
xor U5025 (N_5025,N_1313,N_80);
xnor U5026 (N_5026,N_1932,N_642);
or U5027 (N_5027,N_2393,N_59);
nand U5028 (N_5028,N_629,N_1236);
xor U5029 (N_5029,N_3084,N_1906);
nand U5030 (N_5030,N_1115,N_1068);
nor U5031 (N_5031,N_1714,N_2950);
or U5032 (N_5032,N_978,N_1317);
nor U5033 (N_5033,N_533,N_899);
nor U5034 (N_5034,N_1467,N_1695);
or U5035 (N_5035,N_632,N_1687);
and U5036 (N_5036,N_2854,N_2506);
nand U5037 (N_5037,N_801,N_1184);
xnor U5038 (N_5038,N_675,N_887);
nand U5039 (N_5039,N_1206,N_574);
xnor U5040 (N_5040,N_1328,N_2782);
or U5041 (N_5041,N_2297,N_1538);
and U5042 (N_5042,N_129,N_2595);
nand U5043 (N_5043,N_1610,N_141);
or U5044 (N_5044,N_2379,N_1224);
nand U5045 (N_5045,N_694,N_1220);
and U5046 (N_5046,N_91,N_2429);
and U5047 (N_5047,N_1590,N_2880);
xor U5048 (N_5048,N_597,N_1057);
xnor U5049 (N_5049,N_2422,N_1327);
xor U5050 (N_5050,N_2783,N_2255);
and U5051 (N_5051,N_2060,N_702);
and U5052 (N_5052,N_485,N_1972);
nor U5053 (N_5053,N_1255,N_1240);
or U5054 (N_5054,N_227,N_647);
nand U5055 (N_5055,N_601,N_2359);
xnor U5056 (N_5056,N_1890,N_277);
xnor U5057 (N_5057,N_849,N_1723);
xnor U5058 (N_5058,N_1757,N_2978);
nand U5059 (N_5059,N_2097,N_2121);
and U5060 (N_5060,N_665,N_1824);
or U5061 (N_5061,N_2070,N_1981);
and U5062 (N_5062,N_362,N_1091);
nor U5063 (N_5063,N_1378,N_943);
xnor U5064 (N_5064,N_1045,N_2463);
nor U5065 (N_5065,N_150,N_140);
and U5066 (N_5066,N_922,N_46);
or U5067 (N_5067,N_2312,N_242);
nor U5068 (N_5068,N_165,N_2035);
nor U5069 (N_5069,N_731,N_2685);
and U5070 (N_5070,N_2646,N_2772);
and U5071 (N_5071,N_1707,N_1276);
and U5072 (N_5072,N_2027,N_2180);
or U5073 (N_5073,N_2960,N_3105);
and U5074 (N_5074,N_271,N_499);
and U5075 (N_5075,N_2047,N_1832);
xor U5076 (N_5076,N_2459,N_1895);
and U5077 (N_5077,N_1189,N_1889);
nor U5078 (N_5078,N_24,N_1635);
nand U5079 (N_5079,N_1304,N_2565);
and U5080 (N_5080,N_794,N_1894);
or U5081 (N_5081,N_1587,N_760);
and U5082 (N_5082,N_2305,N_2556);
or U5083 (N_5083,N_2274,N_827);
or U5084 (N_5084,N_367,N_2710);
xnor U5085 (N_5085,N_2158,N_3062);
xnor U5086 (N_5086,N_1835,N_907);
nand U5087 (N_5087,N_1917,N_2171);
and U5088 (N_5088,N_2249,N_337);
and U5089 (N_5089,N_1313,N_3048);
xnor U5090 (N_5090,N_1709,N_575);
and U5091 (N_5091,N_259,N_1251);
or U5092 (N_5092,N_2034,N_1852);
xnor U5093 (N_5093,N_818,N_2008);
and U5094 (N_5094,N_3009,N_489);
nand U5095 (N_5095,N_229,N_1840);
xor U5096 (N_5096,N_2524,N_447);
xnor U5097 (N_5097,N_1265,N_682);
nand U5098 (N_5098,N_1498,N_35);
xnor U5099 (N_5099,N_699,N_1842);
and U5100 (N_5100,N_2648,N_99);
nor U5101 (N_5101,N_1561,N_1369);
and U5102 (N_5102,N_2235,N_2735);
nand U5103 (N_5103,N_1633,N_2940);
or U5104 (N_5104,N_631,N_464);
or U5105 (N_5105,N_141,N_973);
or U5106 (N_5106,N_2386,N_2165);
nor U5107 (N_5107,N_1859,N_120);
and U5108 (N_5108,N_203,N_2509);
and U5109 (N_5109,N_198,N_1653);
nor U5110 (N_5110,N_1899,N_2944);
xnor U5111 (N_5111,N_3121,N_1997);
nand U5112 (N_5112,N_2205,N_1652);
nand U5113 (N_5113,N_2752,N_227);
and U5114 (N_5114,N_1938,N_837);
xnor U5115 (N_5115,N_455,N_2929);
or U5116 (N_5116,N_798,N_858);
nand U5117 (N_5117,N_1930,N_1309);
and U5118 (N_5118,N_2943,N_2801);
xor U5119 (N_5119,N_1020,N_3115);
nand U5120 (N_5120,N_2763,N_303);
and U5121 (N_5121,N_2886,N_1688);
nor U5122 (N_5122,N_1500,N_919);
nor U5123 (N_5123,N_1154,N_131);
nand U5124 (N_5124,N_2252,N_3036);
and U5125 (N_5125,N_792,N_1111);
xor U5126 (N_5126,N_2159,N_2553);
nand U5127 (N_5127,N_1616,N_553);
nand U5128 (N_5128,N_6,N_930);
or U5129 (N_5129,N_1296,N_160);
nand U5130 (N_5130,N_1969,N_968);
xor U5131 (N_5131,N_977,N_1396);
nand U5132 (N_5132,N_3100,N_666);
or U5133 (N_5133,N_1131,N_2313);
xnor U5134 (N_5134,N_2691,N_2056);
or U5135 (N_5135,N_1745,N_2427);
nor U5136 (N_5136,N_1181,N_1125);
and U5137 (N_5137,N_532,N_2575);
and U5138 (N_5138,N_1439,N_2919);
or U5139 (N_5139,N_734,N_1970);
xor U5140 (N_5140,N_150,N_1895);
or U5141 (N_5141,N_2130,N_471);
xor U5142 (N_5142,N_711,N_726);
xor U5143 (N_5143,N_766,N_777);
xor U5144 (N_5144,N_1622,N_3034);
xnor U5145 (N_5145,N_436,N_1681);
xor U5146 (N_5146,N_3021,N_163);
and U5147 (N_5147,N_913,N_2360);
and U5148 (N_5148,N_1628,N_1633);
nand U5149 (N_5149,N_2528,N_2706);
nand U5150 (N_5150,N_2246,N_2223);
nand U5151 (N_5151,N_1685,N_1001);
and U5152 (N_5152,N_2948,N_2196);
nor U5153 (N_5153,N_2933,N_2232);
or U5154 (N_5154,N_1649,N_1316);
and U5155 (N_5155,N_2552,N_1523);
or U5156 (N_5156,N_722,N_2803);
or U5157 (N_5157,N_2315,N_532);
xor U5158 (N_5158,N_2966,N_602);
xor U5159 (N_5159,N_2792,N_498);
nand U5160 (N_5160,N_1517,N_999);
or U5161 (N_5161,N_2639,N_950);
xnor U5162 (N_5162,N_1024,N_2986);
xor U5163 (N_5163,N_21,N_1570);
xnor U5164 (N_5164,N_579,N_1487);
xor U5165 (N_5165,N_474,N_2486);
nand U5166 (N_5166,N_139,N_1522);
xnor U5167 (N_5167,N_2147,N_1298);
nand U5168 (N_5168,N_2416,N_392);
or U5169 (N_5169,N_1714,N_2072);
nand U5170 (N_5170,N_2556,N_2825);
or U5171 (N_5171,N_2019,N_1947);
xnor U5172 (N_5172,N_334,N_1185);
nand U5173 (N_5173,N_2967,N_1840);
nand U5174 (N_5174,N_1102,N_827);
xnor U5175 (N_5175,N_679,N_2722);
nand U5176 (N_5176,N_1924,N_2099);
xnor U5177 (N_5177,N_2439,N_340);
or U5178 (N_5178,N_1429,N_2154);
and U5179 (N_5179,N_2727,N_1927);
nor U5180 (N_5180,N_2928,N_2217);
nor U5181 (N_5181,N_164,N_565);
nor U5182 (N_5182,N_1597,N_1631);
and U5183 (N_5183,N_1797,N_3099);
and U5184 (N_5184,N_1792,N_93);
and U5185 (N_5185,N_3101,N_278);
xnor U5186 (N_5186,N_514,N_2668);
xnor U5187 (N_5187,N_2686,N_273);
xnor U5188 (N_5188,N_658,N_1854);
or U5189 (N_5189,N_2485,N_703);
xor U5190 (N_5190,N_2312,N_327);
nand U5191 (N_5191,N_3064,N_1260);
and U5192 (N_5192,N_2154,N_452);
nand U5193 (N_5193,N_1019,N_2285);
nand U5194 (N_5194,N_2849,N_34);
or U5195 (N_5195,N_2792,N_1893);
or U5196 (N_5196,N_2088,N_2202);
nor U5197 (N_5197,N_581,N_34);
or U5198 (N_5198,N_1817,N_1864);
nor U5199 (N_5199,N_1623,N_571);
nor U5200 (N_5200,N_685,N_2941);
nand U5201 (N_5201,N_609,N_1516);
nand U5202 (N_5202,N_2377,N_742);
nand U5203 (N_5203,N_1088,N_1603);
nor U5204 (N_5204,N_2245,N_2519);
nor U5205 (N_5205,N_916,N_1897);
or U5206 (N_5206,N_1130,N_1068);
or U5207 (N_5207,N_2621,N_1253);
or U5208 (N_5208,N_879,N_2349);
and U5209 (N_5209,N_1779,N_2503);
nand U5210 (N_5210,N_1987,N_2846);
and U5211 (N_5211,N_1207,N_2716);
nor U5212 (N_5212,N_2759,N_1808);
nor U5213 (N_5213,N_3053,N_2339);
nand U5214 (N_5214,N_589,N_1541);
xor U5215 (N_5215,N_645,N_1907);
xnor U5216 (N_5216,N_3029,N_394);
xor U5217 (N_5217,N_762,N_2036);
xor U5218 (N_5218,N_533,N_2306);
nor U5219 (N_5219,N_1024,N_378);
nor U5220 (N_5220,N_466,N_1611);
nand U5221 (N_5221,N_2503,N_3002);
and U5222 (N_5222,N_212,N_956);
or U5223 (N_5223,N_759,N_2748);
xor U5224 (N_5224,N_1640,N_1756);
or U5225 (N_5225,N_545,N_2338);
and U5226 (N_5226,N_222,N_742);
or U5227 (N_5227,N_2142,N_1584);
and U5228 (N_5228,N_8,N_2151);
and U5229 (N_5229,N_1594,N_908);
nand U5230 (N_5230,N_2619,N_885);
nand U5231 (N_5231,N_913,N_997);
nor U5232 (N_5232,N_2564,N_1076);
and U5233 (N_5233,N_2243,N_486);
nor U5234 (N_5234,N_800,N_1300);
and U5235 (N_5235,N_1099,N_2262);
and U5236 (N_5236,N_2952,N_1115);
and U5237 (N_5237,N_839,N_2001);
or U5238 (N_5238,N_127,N_1947);
xor U5239 (N_5239,N_116,N_61);
xor U5240 (N_5240,N_1485,N_641);
nand U5241 (N_5241,N_985,N_764);
xnor U5242 (N_5242,N_2068,N_3078);
nand U5243 (N_5243,N_786,N_545);
nor U5244 (N_5244,N_2540,N_239);
nor U5245 (N_5245,N_2740,N_249);
nor U5246 (N_5246,N_703,N_2340);
nand U5247 (N_5247,N_2237,N_2673);
xor U5248 (N_5248,N_2537,N_2422);
xnor U5249 (N_5249,N_921,N_3041);
xnor U5250 (N_5250,N_250,N_1255);
xnor U5251 (N_5251,N_2406,N_444);
nand U5252 (N_5252,N_2761,N_1152);
or U5253 (N_5253,N_2914,N_544);
nand U5254 (N_5254,N_285,N_2271);
or U5255 (N_5255,N_1525,N_3105);
nor U5256 (N_5256,N_1295,N_2690);
nand U5257 (N_5257,N_2753,N_2938);
xor U5258 (N_5258,N_2502,N_1378);
nand U5259 (N_5259,N_404,N_2113);
or U5260 (N_5260,N_2410,N_2858);
xnor U5261 (N_5261,N_390,N_617);
or U5262 (N_5262,N_483,N_486);
or U5263 (N_5263,N_364,N_1629);
nor U5264 (N_5264,N_111,N_2065);
and U5265 (N_5265,N_1092,N_2002);
nor U5266 (N_5266,N_1515,N_2215);
xor U5267 (N_5267,N_548,N_678);
nor U5268 (N_5268,N_1982,N_1644);
and U5269 (N_5269,N_2468,N_2940);
nor U5270 (N_5270,N_1076,N_2640);
nand U5271 (N_5271,N_2921,N_742);
nand U5272 (N_5272,N_2758,N_2081);
or U5273 (N_5273,N_1023,N_1584);
or U5274 (N_5274,N_1189,N_685);
xor U5275 (N_5275,N_1744,N_2056);
and U5276 (N_5276,N_84,N_2789);
nor U5277 (N_5277,N_2790,N_2980);
or U5278 (N_5278,N_601,N_276);
nor U5279 (N_5279,N_2183,N_139);
nor U5280 (N_5280,N_277,N_1281);
and U5281 (N_5281,N_2646,N_1482);
nand U5282 (N_5282,N_2411,N_1316);
and U5283 (N_5283,N_2400,N_3021);
and U5284 (N_5284,N_340,N_432);
nor U5285 (N_5285,N_1689,N_2209);
or U5286 (N_5286,N_264,N_775);
xnor U5287 (N_5287,N_2749,N_1174);
xor U5288 (N_5288,N_1724,N_1928);
and U5289 (N_5289,N_2409,N_18);
xor U5290 (N_5290,N_194,N_15);
nand U5291 (N_5291,N_1566,N_844);
xor U5292 (N_5292,N_226,N_719);
and U5293 (N_5293,N_668,N_1096);
and U5294 (N_5294,N_1428,N_1885);
or U5295 (N_5295,N_1947,N_162);
xnor U5296 (N_5296,N_1197,N_1476);
xnor U5297 (N_5297,N_2846,N_2826);
or U5298 (N_5298,N_927,N_717);
or U5299 (N_5299,N_2242,N_1813);
and U5300 (N_5300,N_2323,N_2929);
and U5301 (N_5301,N_1428,N_270);
nand U5302 (N_5302,N_924,N_1993);
nand U5303 (N_5303,N_139,N_2961);
or U5304 (N_5304,N_30,N_2732);
and U5305 (N_5305,N_1356,N_1174);
nand U5306 (N_5306,N_987,N_896);
nor U5307 (N_5307,N_2401,N_1660);
and U5308 (N_5308,N_1178,N_2404);
nor U5309 (N_5309,N_415,N_2490);
nor U5310 (N_5310,N_2860,N_344);
or U5311 (N_5311,N_1377,N_247);
or U5312 (N_5312,N_1356,N_3004);
or U5313 (N_5313,N_1777,N_2971);
or U5314 (N_5314,N_38,N_1633);
nand U5315 (N_5315,N_3098,N_3004);
xnor U5316 (N_5316,N_1045,N_96);
and U5317 (N_5317,N_1047,N_1867);
nor U5318 (N_5318,N_551,N_1652);
or U5319 (N_5319,N_2047,N_402);
nor U5320 (N_5320,N_1012,N_1933);
and U5321 (N_5321,N_2941,N_1608);
and U5322 (N_5322,N_860,N_3124);
or U5323 (N_5323,N_116,N_1609);
nor U5324 (N_5324,N_1245,N_1017);
and U5325 (N_5325,N_959,N_777);
xnor U5326 (N_5326,N_2535,N_2549);
nand U5327 (N_5327,N_2766,N_468);
nor U5328 (N_5328,N_2658,N_2758);
nand U5329 (N_5329,N_2531,N_256);
nand U5330 (N_5330,N_178,N_2594);
and U5331 (N_5331,N_2520,N_1524);
or U5332 (N_5332,N_2330,N_160);
xnor U5333 (N_5333,N_386,N_2353);
or U5334 (N_5334,N_1143,N_1282);
nor U5335 (N_5335,N_369,N_455);
or U5336 (N_5336,N_2019,N_2394);
nor U5337 (N_5337,N_1357,N_2182);
nand U5338 (N_5338,N_1185,N_2700);
and U5339 (N_5339,N_728,N_1482);
xnor U5340 (N_5340,N_1741,N_72);
nand U5341 (N_5341,N_1145,N_656);
nand U5342 (N_5342,N_953,N_239);
and U5343 (N_5343,N_2625,N_222);
nand U5344 (N_5344,N_1966,N_2009);
nor U5345 (N_5345,N_2038,N_541);
xor U5346 (N_5346,N_119,N_1464);
xor U5347 (N_5347,N_315,N_481);
nor U5348 (N_5348,N_2354,N_2025);
xor U5349 (N_5349,N_16,N_1938);
or U5350 (N_5350,N_2240,N_439);
or U5351 (N_5351,N_2365,N_2358);
xor U5352 (N_5352,N_41,N_439);
and U5353 (N_5353,N_388,N_2367);
nor U5354 (N_5354,N_232,N_1980);
nor U5355 (N_5355,N_2364,N_1500);
nand U5356 (N_5356,N_1964,N_1321);
or U5357 (N_5357,N_119,N_2901);
or U5358 (N_5358,N_524,N_2876);
and U5359 (N_5359,N_100,N_2783);
xnor U5360 (N_5360,N_1644,N_1377);
nor U5361 (N_5361,N_15,N_2661);
nor U5362 (N_5362,N_1489,N_2500);
or U5363 (N_5363,N_314,N_1556);
and U5364 (N_5364,N_2644,N_2980);
and U5365 (N_5365,N_2204,N_1188);
and U5366 (N_5366,N_904,N_2246);
xor U5367 (N_5367,N_320,N_2398);
or U5368 (N_5368,N_2250,N_2464);
nand U5369 (N_5369,N_374,N_856);
nor U5370 (N_5370,N_1810,N_367);
and U5371 (N_5371,N_528,N_774);
or U5372 (N_5372,N_2789,N_2927);
nand U5373 (N_5373,N_53,N_491);
xnor U5374 (N_5374,N_514,N_384);
or U5375 (N_5375,N_1665,N_2396);
nor U5376 (N_5376,N_2785,N_2434);
nand U5377 (N_5377,N_48,N_1200);
xor U5378 (N_5378,N_687,N_2358);
xnor U5379 (N_5379,N_59,N_1535);
and U5380 (N_5380,N_192,N_1611);
nor U5381 (N_5381,N_1,N_527);
and U5382 (N_5382,N_2398,N_368);
and U5383 (N_5383,N_1354,N_139);
and U5384 (N_5384,N_1596,N_669);
nor U5385 (N_5385,N_966,N_1117);
and U5386 (N_5386,N_258,N_439);
xnor U5387 (N_5387,N_1658,N_2274);
nor U5388 (N_5388,N_593,N_3063);
and U5389 (N_5389,N_2250,N_464);
xnor U5390 (N_5390,N_1479,N_132);
nand U5391 (N_5391,N_2395,N_47);
or U5392 (N_5392,N_2887,N_2613);
and U5393 (N_5393,N_1095,N_859);
nor U5394 (N_5394,N_2806,N_2246);
and U5395 (N_5395,N_2307,N_295);
xnor U5396 (N_5396,N_93,N_1610);
nor U5397 (N_5397,N_2633,N_246);
nor U5398 (N_5398,N_1896,N_153);
nand U5399 (N_5399,N_1551,N_1423);
xnor U5400 (N_5400,N_604,N_526);
xnor U5401 (N_5401,N_1223,N_3037);
or U5402 (N_5402,N_1984,N_2862);
and U5403 (N_5403,N_979,N_2816);
and U5404 (N_5404,N_333,N_980);
nand U5405 (N_5405,N_2585,N_225);
nor U5406 (N_5406,N_2344,N_691);
or U5407 (N_5407,N_1905,N_2999);
nor U5408 (N_5408,N_1095,N_1211);
nand U5409 (N_5409,N_735,N_1167);
or U5410 (N_5410,N_2134,N_1832);
xor U5411 (N_5411,N_38,N_651);
xor U5412 (N_5412,N_671,N_2766);
nand U5413 (N_5413,N_2429,N_630);
or U5414 (N_5414,N_2802,N_2913);
and U5415 (N_5415,N_2481,N_197);
nand U5416 (N_5416,N_1400,N_1620);
nand U5417 (N_5417,N_529,N_2281);
nor U5418 (N_5418,N_2339,N_98);
or U5419 (N_5419,N_2781,N_2001);
xnor U5420 (N_5420,N_763,N_2059);
nor U5421 (N_5421,N_679,N_2744);
or U5422 (N_5422,N_137,N_2506);
nand U5423 (N_5423,N_1218,N_1210);
nor U5424 (N_5424,N_2516,N_1356);
xnor U5425 (N_5425,N_308,N_106);
xor U5426 (N_5426,N_2940,N_2989);
or U5427 (N_5427,N_2466,N_1688);
nor U5428 (N_5428,N_1807,N_1656);
or U5429 (N_5429,N_2945,N_1637);
nand U5430 (N_5430,N_702,N_529);
xnor U5431 (N_5431,N_777,N_327);
nand U5432 (N_5432,N_2520,N_153);
nor U5433 (N_5433,N_1526,N_2335);
or U5434 (N_5434,N_774,N_472);
nand U5435 (N_5435,N_1814,N_2133);
nor U5436 (N_5436,N_1525,N_1964);
xnor U5437 (N_5437,N_2784,N_1144);
nand U5438 (N_5438,N_1230,N_1724);
xnor U5439 (N_5439,N_1831,N_1545);
nand U5440 (N_5440,N_2355,N_256);
or U5441 (N_5441,N_1924,N_2288);
nor U5442 (N_5442,N_2287,N_1751);
nand U5443 (N_5443,N_3044,N_3078);
nand U5444 (N_5444,N_320,N_1788);
nand U5445 (N_5445,N_3060,N_1181);
nand U5446 (N_5446,N_2725,N_281);
and U5447 (N_5447,N_217,N_218);
xor U5448 (N_5448,N_1878,N_428);
xor U5449 (N_5449,N_2389,N_729);
nor U5450 (N_5450,N_60,N_3059);
and U5451 (N_5451,N_2428,N_2878);
nand U5452 (N_5452,N_713,N_1897);
or U5453 (N_5453,N_372,N_1106);
or U5454 (N_5454,N_2801,N_163);
or U5455 (N_5455,N_1079,N_2780);
nand U5456 (N_5456,N_1803,N_2893);
or U5457 (N_5457,N_2916,N_2311);
xnor U5458 (N_5458,N_1409,N_2833);
nor U5459 (N_5459,N_2148,N_129);
and U5460 (N_5460,N_225,N_3023);
nand U5461 (N_5461,N_1233,N_1365);
or U5462 (N_5462,N_758,N_2622);
nand U5463 (N_5463,N_1234,N_1533);
nor U5464 (N_5464,N_596,N_1340);
or U5465 (N_5465,N_2480,N_149);
or U5466 (N_5466,N_863,N_1261);
xnor U5467 (N_5467,N_2380,N_2675);
or U5468 (N_5468,N_1256,N_2418);
nor U5469 (N_5469,N_500,N_594);
nor U5470 (N_5470,N_728,N_2627);
nand U5471 (N_5471,N_2870,N_676);
nor U5472 (N_5472,N_842,N_2023);
or U5473 (N_5473,N_470,N_2049);
xnor U5474 (N_5474,N_771,N_1474);
nor U5475 (N_5475,N_1586,N_703);
nand U5476 (N_5476,N_357,N_399);
nand U5477 (N_5477,N_1249,N_1424);
nand U5478 (N_5478,N_7,N_1240);
or U5479 (N_5479,N_1700,N_555);
xor U5480 (N_5480,N_491,N_1262);
or U5481 (N_5481,N_993,N_1864);
and U5482 (N_5482,N_991,N_1965);
and U5483 (N_5483,N_342,N_2846);
xor U5484 (N_5484,N_1901,N_2730);
nand U5485 (N_5485,N_1784,N_2080);
and U5486 (N_5486,N_1312,N_2561);
xor U5487 (N_5487,N_2502,N_2673);
and U5488 (N_5488,N_3033,N_1643);
and U5489 (N_5489,N_1338,N_612);
xor U5490 (N_5490,N_2967,N_2175);
or U5491 (N_5491,N_1195,N_3122);
nand U5492 (N_5492,N_1793,N_2697);
xor U5493 (N_5493,N_2417,N_106);
and U5494 (N_5494,N_1233,N_2355);
nand U5495 (N_5495,N_2075,N_2013);
and U5496 (N_5496,N_143,N_469);
and U5497 (N_5497,N_2392,N_845);
and U5498 (N_5498,N_697,N_2873);
or U5499 (N_5499,N_2580,N_2126);
xor U5500 (N_5500,N_2955,N_2616);
nor U5501 (N_5501,N_2063,N_2309);
xnor U5502 (N_5502,N_1175,N_1635);
nand U5503 (N_5503,N_1140,N_1170);
nor U5504 (N_5504,N_464,N_2362);
and U5505 (N_5505,N_658,N_1692);
xor U5506 (N_5506,N_3078,N_1189);
nor U5507 (N_5507,N_3008,N_2225);
or U5508 (N_5508,N_1304,N_2102);
nand U5509 (N_5509,N_1891,N_2555);
nand U5510 (N_5510,N_925,N_210);
or U5511 (N_5511,N_2302,N_1153);
or U5512 (N_5512,N_2165,N_288);
nor U5513 (N_5513,N_1165,N_1879);
xnor U5514 (N_5514,N_2331,N_747);
nand U5515 (N_5515,N_1751,N_2782);
xor U5516 (N_5516,N_1561,N_229);
or U5517 (N_5517,N_764,N_2955);
or U5518 (N_5518,N_1181,N_1803);
nand U5519 (N_5519,N_3020,N_2333);
nor U5520 (N_5520,N_2016,N_2785);
xnor U5521 (N_5521,N_2464,N_651);
or U5522 (N_5522,N_2842,N_1740);
and U5523 (N_5523,N_2883,N_37);
or U5524 (N_5524,N_128,N_148);
nand U5525 (N_5525,N_208,N_1181);
or U5526 (N_5526,N_1855,N_735);
or U5527 (N_5527,N_2546,N_48);
or U5528 (N_5528,N_1945,N_2682);
nor U5529 (N_5529,N_2964,N_243);
nor U5530 (N_5530,N_2357,N_1186);
and U5531 (N_5531,N_1480,N_2491);
xor U5532 (N_5532,N_2586,N_2700);
xnor U5533 (N_5533,N_1983,N_1587);
or U5534 (N_5534,N_1018,N_496);
and U5535 (N_5535,N_911,N_1429);
nand U5536 (N_5536,N_2771,N_2441);
nand U5537 (N_5537,N_2959,N_1810);
nor U5538 (N_5538,N_2793,N_2335);
or U5539 (N_5539,N_1449,N_3012);
nand U5540 (N_5540,N_691,N_2475);
xnor U5541 (N_5541,N_347,N_1700);
nand U5542 (N_5542,N_1468,N_733);
xnor U5543 (N_5543,N_2232,N_1931);
nand U5544 (N_5544,N_2733,N_2572);
xor U5545 (N_5545,N_1202,N_2702);
xnor U5546 (N_5546,N_2859,N_92);
or U5547 (N_5547,N_490,N_410);
nor U5548 (N_5548,N_1421,N_800);
or U5549 (N_5549,N_1259,N_1988);
nor U5550 (N_5550,N_1642,N_325);
nand U5551 (N_5551,N_1801,N_2915);
and U5552 (N_5552,N_757,N_617);
xor U5553 (N_5553,N_517,N_2403);
nor U5554 (N_5554,N_2485,N_1989);
nor U5555 (N_5555,N_915,N_3116);
and U5556 (N_5556,N_5,N_373);
nor U5557 (N_5557,N_448,N_1018);
xor U5558 (N_5558,N_1711,N_1797);
and U5559 (N_5559,N_2684,N_2785);
xnor U5560 (N_5560,N_3061,N_217);
nor U5561 (N_5561,N_2428,N_1081);
xor U5562 (N_5562,N_160,N_699);
nand U5563 (N_5563,N_214,N_987);
and U5564 (N_5564,N_847,N_362);
and U5565 (N_5565,N_2509,N_1579);
nand U5566 (N_5566,N_1299,N_2617);
nand U5567 (N_5567,N_609,N_530);
nor U5568 (N_5568,N_1887,N_2445);
or U5569 (N_5569,N_441,N_2744);
xor U5570 (N_5570,N_86,N_925);
nand U5571 (N_5571,N_1508,N_89);
or U5572 (N_5572,N_703,N_2433);
and U5573 (N_5573,N_2519,N_2150);
nand U5574 (N_5574,N_865,N_1874);
or U5575 (N_5575,N_1604,N_1909);
or U5576 (N_5576,N_974,N_2897);
nand U5577 (N_5577,N_2696,N_1113);
nor U5578 (N_5578,N_2086,N_2035);
or U5579 (N_5579,N_744,N_741);
nand U5580 (N_5580,N_1006,N_373);
and U5581 (N_5581,N_1,N_1428);
and U5582 (N_5582,N_244,N_149);
nor U5583 (N_5583,N_309,N_1499);
nor U5584 (N_5584,N_1766,N_3077);
or U5585 (N_5585,N_2574,N_3072);
xnor U5586 (N_5586,N_305,N_1029);
nand U5587 (N_5587,N_1329,N_161);
xnor U5588 (N_5588,N_47,N_295);
xor U5589 (N_5589,N_228,N_58);
nor U5590 (N_5590,N_2419,N_3004);
nand U5591 (N_5591,N_2824,N_1124);
xnor U5592 (N_5592,N_644,N_472);
nand U5593 (N_5593,N_2079,N_1487);
and U5594 (N_5594,N_2873,N_898);
or U5595 (N_5595,N_1212,N_2569);
nand U5596 (N_5596,N_526,N_2634);
or U5597 (N_5597,N_1737,N_1391);
xor U5598 (N_5598,N_216,N_2497);
nor U5599 (N_5599,N_1897,N_2160);
nand U5600 (N_5600,N_999,N_1544);
xor U5601 (N_5601,N_2610,N_946);
xnor U5602 (N_5602,N_75,N_1632);
and U5603 (N_5603,N_580,N_2565);
or U5604 (N_5604,N_686,N_195);
nor U5605 (N_5605,N_2956,N_1267);
and U5606 (N_5606,N_1513,N_456);
and U5607 (N_5607,N_1973,N_1445);
and U5608 (N_5608,N_1454,N_300);
nor U5609 (N_5609,N_1482,N_311);
xnor U5610 (N_5610,N_1274,N_877);
or U5611 (N_5611,N_1474,N_880);
or U5612 (N_5612,N_657,N_1511);
nand U5613 (N_5613,N_1892,N_686);
or U5614 (N_5614,N_2152,N_2768);
and U5615 (N_5615,N_484,N_1766);
and U5616 (N_5616,N_1462,N_260);
or U5617 (N_5617,N_973,N_3071);
and U5618 (N_5618,N_654,N_555);
xor U5619 (N_5619,N_1975,N_3063);
xnor U5620 (N_5620,N_1806,N_2705);
and U5621 (N_5621,N_1316,N_34);
xnor U5622 (N_5622,N_2939,N_2907);
nand U5623 (N_5623,N_1434,N_458);
nor U5624 (N_5624,N_562,N_1779);
nand U5625 (N_5625,N_994,N_1344);
nand U5626 (N_5626,N_1046,N_1466);
nand U5627 (N_5627,N_903,N_743);
nor U5628 (N_5628,N_2022,N_375);
nor U5629 (N_5629,N_2554,N_2547);
nand U5630 (N_5630,N_1941,N_530);
or U5631 (N_5631,N_652,N_1657);
and U5632 (N_5632,N_1759,N_2513);
or U5633 (N_5633,N_2315,N_714);
nor U5634 (N_5634,N_2817,N_1454);
nor U5635 (N_5635,N_350,N_2976);
and U5636 (N_5636,N_2243,N_177);
nand U5637 (N_5637,N_2112,N_1783);
and U5638 (N_5638,N_3051,N_610);
nor U5639 (N_5639,N_1886,N_1474);
xor U5640 (N_5640,N_432,N_2368);
or U5641 (N_5641,N_2660,N_514);
xor U5642 (N_5642,N_1233,N_2512);
nand U5643 (N_5643,N_1336,N_787);
and U5644 (N_5644,N_1100,N_2667);
xnor U5645 (N_5645,N_2034,N_1521);
or U5646 (N_5646,N_1802,N_1781);
or U5647 (N_5647,N_1799,N_493);
or U5648 (N_5648,N_3017,N_2036);
nor U5649 (N_5649,N_2632,N_628);
nand U5650 (N_5650,N_128,N_2314);
nor U5651 (N_5651,N_1012,N_99);
or U5652 (N_5652,N_919,N_2574);
xor U5653 (N_5653,N_1183,N_54);
nor U5654 (N_5654,N_1622,N_185);
nor U5655 (N_5655,N_2683,N_1731);
xor U5656 (N_5656,N_815,N_1174);
nor U5657 (N_5657,N_1858,N_2797);
or U5658 (N_5658,N_1512,N_2107);
or U5659 (N_5659,N_2408,N_543);
nor U5660 (N_5660,N_2357,N_397);
or U5661 (N_5661,N_2887,N_2922);
and U5662 (N_5662,N_501,N_450);
or U5663 (N_5663,N_572,N_1326);
nand U5664 (N_5664,N_1342,N_2042);
and U5665 (N_5665,N_2728,N_2199);
nand U5666 (N_5666,N_717,N_2227);
xnor U5667 (N_5667,N_868,N_2417);
xnor U5668 (N_5668,N_1326,N_975);
or U5669 (N_5669,N_2224,N_2099);
and U5670 (N_5670,N_1653,N_1723);
nor U5671 (N_5671,N_2820,N_2391);
and U5672 (N_5672,N_2468,N_943);
nor U5673 (N_5673,N_2614,N_2607);
or U5674 (N_5674,N_1808,N_1150);
and U5675 (N_5675,N_2521,N_889);
nor U5676 (N_5676,N_197,N_1141);
or U5677 (N_5677,N_2878,N_1607);
nor U5678 (N_5678,N_1957,N_1701);
xor U5679 (N_5679,N_670,N_297);
nand U5680 (N_5680,N_1608,N_2033);
nor U5681 (N_5681,N_2261,N_1131);
nor U5682 (N_5682,N_2641,N_624);
xnor U5683 (N_5683,N_1687,N_729);
nand U5684 (N_5684,N_2328,N_2365);
nor U5685 (N_5685,N_2658,N_2467);
or U5686 (N_5686,N_1345,N_592);
and U5687 (N_5687,N_2123,N_1980);
nor U5688 (N_5688,N_821,N_2674);
nand U5689 (N_5689,N_2600,N_728);
and U5690 (N_5690,N_2680,N_747);
and U5691 (N_5691,N_123,N_1113);
nand U5692 (N_5692,N_2908,N_2373);
nand U5693 (N_5693,N_1912,N_2453);
nand U5694 (N_5694,N_190,N_3121);
xnor U5695 (N_5695,N_2160,N_1308);
xnor U5696 (N_5696,N_974,N_1870);
xnor U5697 (N_5697,N_544,N_2973);
xnor U5698 (N_5698,N_2535,N_95);
nand U5699 (N_5699,N_340,N_2901);
or U5700 (N_5700,N_1026,N_1394);
nand U5701 (N_5701,N_900,N_455);
or U5702 (N_5702,N_1244,N_185);
and U5703 (N_5703,N_747,N_2214);
xnor U5704 (N_5704,N_2474,N_542);
nor U5705 (N_5705,N_2436,N_2201);
nor U5706 (N_5706,N_1322,N_285);
or U5707 (N_5707,N_2452,N_937);
nand U5708 (N_5708,N_115,N_1087);
or U5709 (N_5709,N_874,N_1652);
and U5710 (N_5710,N_1918,N_1450);
and U5711 (N_5711,N_2849,N_1079);
or U5712 (N_5712,N_2604,N_1321);
or U5713 (N_5713,N_2075,N_260);
nand U5714 (N_5714,N_2067,N_1963);
nand U5715 (N_5715,N_106,N_1957);
or U5716 (N_5716,N_1008,N_1724);
nand U5717 (N_5717,N_531,N_88);
nand U5718 (N_5718,N_2862,N_384);
and U5719 (N_5719,N_2579,N_2277);
and U5720 (N_5720,N_1741,N_2299);
xor U5721 (N_5721,N_2872,N_2752);
or U5722 (N_5722,N_2264,N_323);
nor U5723 (N_5723,N_520,N_135);
nor U5724 (N_5724,N_2872,N_2136);
and U5725 (N_5725,N_2816,N_1314);
nand U5726 (N_5726,N_2990,N_1167);
xnor U5727 (N_5727,N_868,N_2828);
xor U5728 (N_5728,N_2226,N_755);
or U5729 (N_5729,N_2418,N_1874);
and U5730 (N_5730,N_15,N_2871);
nor U5731 (N_5731,N_1507,N_1832);
and U5732 (N_5732,N_56,N_1048);
nor U5733 (N_5733,N_1474,N_851);
or U5734 (N_5734,N_1005,N_1143);
xor U5735 (N_5735,N_1113,N_1328);
nor U5736 (N_5736,N_48,N_781);
nand U5737 (N_5737,N_361,N_54);
nor U5738 (N_5738,N_1709,N_2621);
nand U5739 (N_5739,N_2012,N_2219);
and U5740 (N_5740,N_2431,N_1633);
xor U5741 (N_5741,N_1082,N_734);
nor U5742 (N_5742,N_2884,N_737);
and U5743 (N_5743,N_2926,N_2488);
and U5744 (N_5744,N_721,N_1566);
nand U5745 (N_5745,N_1412,N_3060);
or U5746 (N_5746,N_1509,N_2444);
or U5747 (N_5747,N_1852,N_1785);
or U5748 (N_5748,N_2406,N_2077);
and U5749 (N_5749,N_1458,N_1161);
nor U5750 (N_5750,N_2769,N_553);
and U5751 (N_5751,N_2885,N_2974);
nor U5752 (N_5752,N_1716,N_2286);
and U5753 (N_5753,N_156,N_2464);
nand U5754 (N_5754,N_1268,N_1361);
or U5755 (N_5755,N_2429,N_3024);
or U5756 (N_5756,N_1278,N_2668);
nand U5757 (N_5757,N_764,N_54);
and U5758 (N_5758,N_2767,N_216);
nand U5759 (N_5759,N_2574,N_1152);
and U5760 (N_5760,N_2520,N_2946);
nand U5761 (N_5761,N_3002,N_323);
xor U5762 (N_5762,N_1096,N_1573);
or U5763 (N_5763,N_644,N_2603);
xor U5764 (N_5764,N_2904,N_1893);
or U5765 (N_5765,N_2995,N_2950);
nor U5766 (N_5766,N_2480,N_1915);
nand U5767 (N_5767,N_2026,N_306);
nor U5768 (N_5768,N_2095,N_2221);
and U5769 (N_5769,N_1140,N_2367);
and U5770 (N_5770,N_80,N_1078);
and U5771 (N_5771,N_174,N_875);
nor U5772 (N_5772,N_2194,N_2899);
and U5773 (N_5773,N_906,N_2530);
or U5774 (N_5774,N_1538,N_2072);
and U5775 (N_5775,N_2205,N_1611);
and U5776 (N_5776,N_169,N_1234);
nand U5777 (N_5777,N_2662,N_939);
or U5778 (N_5778,N_136,N_1060);
and U5779 (N_5779,N_2045,N_576);
xor U5780 (N_5780,N_520,N_2265);
xor U5781 (N_5781,N_863,N_2765);
and U5782 (N_5782,N_198,N_692);
xnor U5783 (N_5783,N_2760,N_1883);
or U5784 (N_5784,N_1269,N_2164);
nand U5785 (N_5785,N_1300,N_628);
nand U5786 (N_5786,N_556,N_468);
or U5787 (N_5787,N_1208,N_520);
nand U5788 (N_5788,N_1260,N_351);
nor U5789 (N_5789,N_1856,N_1093);
and U5790 (N_5790,N_2294,N_494);
or U5791 (N_5791,N_36,N_118);
nor U5792 (N_5792,N_684,N_768);
and U5793 (N_5793,N_1551,N_2637);
nand U5794 (N_5794,N_1024,N_2972);
and U5795 (N_5795,N_1832,N_2664);
nand U5796 (N_5796,N_1919,N_2565);
nor U5797 (N_5797,N_2455,N_1001);
nor U5798 (N_5798,N_757,N_1828);
and U5799 (N_5799,N_445,N_1617);
and U5800 (N_5800,N_748,N_199);
xor U5801 (N_5801,N_1890,N_2249);
nand U5802 (N_5802,N_1884,N_2708);
or U5803 (N_5803,N_807,N_1943);
or U5804 (N_5804,N_3046,N_2350);
nand U5805 (N_5805,N_433,N_1507);
xnor U5806 (N_5806,N_1787,N_624);
xor U5807 (N_5807,N_1481,N_2279);
nand U5808 (N_5808,N_2404,N_1882);
nand U5809 (N_5809,N_1150,N_2832);
and U5810 (N_5810,N_1960,N_1476);
nor U5811 (N_5811,N_155,N_681);
nand U5812 (N_5812,N_1524,N_2361);
nor U5813 (N_5813,N_2407,N_2527);
xnor U5814 (N_5814,N_1165,N_1017);
nand U5815 (N_5815,N_322,N_97);
nor U5816 (N_5816,N_1472,N_1949);
nor U5817 (N_5817,N_962,N_1701);
or U5818 (N_5818,N_1766,N_1612);
nor U5819 (N_5819,N_817,N_1209);
nor U5820 (N_5820,N_2219,N_865);
nor U5821 (N_5821,N_1945,N_1508);
nor U5822 (N_5822,N_2301,N_1326);
and U5823 (N_5823,N_1974,N_2466);
or U5824 (N_5824,N_644,N_141);
or U5825 (N_5825,N_320,N_2099);
and U5826 (N_5826,N_2949,N_120);
nand U5827 (N_5827,N_95,N_611);
or U5828 (N_5828,N_2969,N_837);
and U5829 (N_5829,N_616,N_1577);
and U5830 (N_5830,N_1476,N_1582);
or U5831 (N_5831,N_2464,N_3100);
nor U5832 (N_5832,N_2320,N_1694);
nor U5833 (N_5833,N_2819,N_431);
or U5834 (N_5834,N_1420,N_1815);
nor U5835 (N_5835,N_702,N_2863);
nand U5836 (N_5836,N_914,N_1707);
xor U5837 (N_5837,N_2027,N_2379);
and U5838 (N_5838,N_2288,N_2484);
nor U5839 (N_5839,N_685,N_1625);
nand U5840 (N_5840,N_735,N_1371);
nand U5841 (N_5841,N_210,N_2592);
xnor U5842 (N_5842,N_549,N_716);
or U5843 (N_5843,N_2165,N_134);
and U5844 (N_5844,N_1997,N_1026);
nand U5845 (N_5845,N_869,N_1470);
or U5846 (N_5846,N_650,N_402);
or U5847 (N_5847,N_1171,N_264);
or U5848 (N_5848,N_1872,N_1032);
or U5849 (N_5849,N_2821,N_2726);
nor U5850 (N_5850,N_1586,N_65);
nor U5851 (N_5851,N_2673,N_2762);
or U5852 (N_5852,N_131,N_1802);
or U5853 (N_5853,N_1177,N_2654);
nor U5854 (N_5854,N_3052,N_842);
nor U5855 (N_5855,N_1806,N_68);
xor U5856 (N_5856,N_2076,N_2984);
xnor U5857 (N_5857,N_1098,N_2149);
nor U5858 (N_5858,N_941,N_1342);
nor U5859 (N_5859,N_1100,N_3082);
nand U5860 (N_5860,N_2348,N_839);
xnor U5861 (N_5861,N_1698,N_1119);
or U5862 (N_5862,N_2446,N_2355);
or U5863 (N_5863,N_548,N_1339);
nor U5864 (N_5864,N_1338,N_368);
nand U5865 (N_5865,N_694,N_698);
nor U5866 (N_5866,N_2035,N_1264);
nand U5867 (N_5867,N_1009,N_2872);
xor U5868 (N_5868,N_2336,N_2537);
xnor U5869 (N_5869,N_556,N_516);
or U5870 (N_5870,N_1037,N_998);
or U5871 (N_5871,N_1207,N_1501);
and U5872 (N_5872,N_1546,N_1010);
and U5873 (N_5873,N_2410,N_2448);
and U5874 (N_5874,N_2310,N_2731);
nand U5875 (N_5875,N_1552,N_2712);
nor U5876 (N_5876,N_224,N_2503);
nor U5877 (N_5877,N_613,N_697);
or U5878 (N_5878,N_818,N_1640);
nand U5879 (N_5879,N_308,N_1344);
and U5880 (N_5880,N_2361,N_330);
nand U5881 (N_5881,N_711,N_2549);
and U5882 (N_5882,N_1761,N_1715);
nor U5883 (N_5883,N_1184,N_2247);
nand U5884 (N_5884,N_1693,N_1424);
or U5885 (N_5885,N_284,N_842);
nor U5886 (N_5886,N_431,N_607);
nor U5887 (N_5887,N_577,N_941);
and U5888 (N_5888,N_1788,N_1785);
and U5889 (N_5889,N_1089,N_1411);
nand U5890 (N_5890,N_2169,N_954);
and U5891 (N_5891,N_2112,N_1938);
xor U5892 (N_5892,N_2447,N_3052);
and U5893 (N_5893,N_1320,N_2956);
xor U5894 (N_5894,N_1674,N_377);
nor U5895 (N_5895,N_2440,N_756);
xnor U5896 (N_5896,N_1461,N_1297);
and U5897 (N_5897,N_1382,N_196);
xor U5898 (N_5898,N_138,N_1384);
and U5899 (N_5899,N_2478,N_912);
or U5900 (N_5900,N_1972,N_1358);
nand U5901 (N_5901,N_2667,N_2250);
nor U5902 (N_5902,N_929,N_1383);
or U5903 (N_5903,N_2103,N_2844);
xnor U5904 (N_5904,N_1157,N_2539);
nand U5905 (N_5905,N_2467,N_833);
nor U5906 (N_5906,N_3100,N_1545);
xor U5907 (N_5907,N_478,N_2711);
nand U5908 (N_5908,N_1170,N_1189);
and U5909 (N_5909,N_2591,N_1350);
xnor U5910 (N_5910,N_1374,N_2656);
and U5911 (N_5911,N_3090,N_1877);
xnor U5912 (N_5912,N_1996,N_2825);
or U5913 (N_5913,N_1589,N_1991);
or U5914 (N_5914,N_1520,N_1025);
or U5915 (N_5915,N_1648,N_1370);
or U5916 (N_5916,N_719,N_626);
and U5917 (N_5917,N_1310,N_1833);
or U5918 (N_5918,N_1032,N_2190);
nand U5919 (N_5919,N_2764,N_1821);
xor U5920 (N_5920,N_1714,N_2472);
xor U5921 (N_5921,N_512,N_976);
nor U5922 (N_5922,N_759,N_1890);
nor U5923 (N_5923,N_438,N_1983);
and U5924 (N_5924,N_2510,N_2243);
nor U5925 (N_5925,N_1616,N_306);
or U5926 (N_5926,N_2484,N_280);
xnor U5927 (N_5927,N_2354,N_1276);
or U5928 (N_5928,N_13,N_348);
nand U5929 (N_5929,N_2302,N_1776);
and U5930 (N_5930,N_2176,N_1717);
nor U5931 (N_5931,N_1865,N_2427);
xnor U5932 (N_5932,N_2998,N_2527);
xor U5933 (N_5933,N_2429,N_3090);
nand U5934 (N_5934,N_3041,N_960);
xor U5935 (N_5935,N_2618,N_2921);
or U5936 (N_5936,N_1387,N_909);
nor U5937 (N_5937,N_1324,N_168);
nor U5938 (N_5938,N_2181,N_303);
xnor U5939 (N_5939,N_2549,N_342);
xor U5940 (N_5940,N_2275,N_618);
xnor U5941 (N_5941,N_963,N_878);
and U5942 (N_5942,N_1028,N_2636);
nor U5943 (N_5943,N_2542,N_3089);
nor U5944 (N_5944,N_2818,N_1817);
and U5945 (N_5945,N_1991,N_1578);
nor U5946 (N_5946,N_735,N_1357);
xnor U5947 (N_5947,N_214,N_1516);
and U5948 (N_5948,N_742,N_765);
xor U5949 (N_5949,N_1978,N_2164);
or U5950 (N_5950,N_1968,N_2949);
nor U5951 (N_5951,N_878,N_2979);
and U5952 (N_5952,N_2722,N_1828);
nand U5953 (N_5953,N_808,N_1649);
xnor U5954 (N_5954,N_2070,N_433);
nor U5955 (N_5955,N_222,N_1271);
or U5956 (N_5956,N_999,N_2675);
nor U5957 (N_5957,N_2053,N_2307);
and U5958 (N_5958,N_2474,N_1895);
and U5959 (N_5959,N_232,N_118);
nor U5960 (N_5960,N_2234,N_2974);
xnor U5961 (N_5961,N_1945,N_3046);
and U5962 (N_5962,N_2191,N_2329);
and U5963 (N_5963,N_1039,N_1485);
xor U5964 (N_5964,N_281,N_369);
or U5965 (N_5965,N_2708,N_2688);
nor U5966 (N_5966,N_2031,N_690);
xnor U5967 (N_5967,N_3098,N_116);
xnor U5968 (N_5968,N_1120,N_1246);
nor U5969 (N_5969,N_2759,N_2395);
xor U5970 (N_5970,N_2042,N_2655);
nor U5971 (N_5971,N_2192,N_825);
nor U5972 (N_5972,N_497,N_1550);
xor U5973 (N_5973,N_2193,N_2862);
nor U5974 (N_5974,N_2919,N_1519);
xor U5975 (N_5975,N_2176,N_2445);
or U5976 (N_5976,N_1994,N_1133);
nand U5977 (N_5977,N_2447,N_563);
nand U5978 (N_5978,N_2277,N_1521);
and U5979 (N_5979,N_433,N_2111);
nand U5980 (N_5980,N_2606,N_335);
nor U5981 (N_5981,N_1103,N_803);
nor U5982 (N_5982,N_1255,N_2942);
xor U5983 (N_5983,N_2968,N_2580);
or U5984 (N_5984,N_993,N_344);
nor U5985 (N_5985,N_1301,N_1564);
nand U5986 (N_5986,N_1307,N_935);
and U5987 (N_5987,N_2606,N_840);
nor U5988 (N_5988,N_2126,N_69);
nor U5989 (N_5989,N_2359,N_568);
nand U5990 (N_5990,N_2067,N_2821);
and U5991 (N_5991,N_2985,N_2732);
and U5992 (N_5992,N_2837,N_1857);
nand U5993 (N_5993,N_1249,N_1348);
xnor U5994 (N_5994,N_620,N_1667);
nor U5995 (N_5995,N_2594,N_2734);
xor U5996 (N_5996,N_2088,N_3109);
or U5997 (N_5997,N_1577,N_1028);
nor U5998 (N_5998,N_298,N_2661);
xor U5999 (N_5999,N_2971,N_1074);
nor U6000 (N_6000,N_1409,N_2637);
nand U6001 (N_6001,N_2333,N_1056);
nor U6002 (N_6002,N_2653,N_2202);
xor U6003 (N_6003,N_2271,N_739);
or U6004 (N_6004,N_2674,N_1642);
or U6005 (N_6005,N_1415,N_1101);
or U6006 (N_6006,N_2257,N_1264);
and U6007 (N_6007,N_2601,N_2959);
or U6008 (N_6008,N_2324,N_186);
xor U6009 (N_6009,N_473,N_1576);
and U6010 (N_6010,N_2443,N_506);
nor U6011 (N_6011,N_529,N_1783);
nor U6012 (N_6012,N_2816,N_2720);
nand U6013 (N_6013,N_1952,N_1013);
and U6014 (N_6014,N_2448,N_125);
and U6015 (N_6015,N_1111,N_321);
nand U6016 (N_6016,N_686,N_483);
nor U6017 (N_6017,N_1132,N_3077);
xor U6018 (N_6018,N_420,N_251);
nand U6019 (N_6019,N_2108,N_2393);
xnor U6020 (N_6020,N_1331,N_1582);
xor U6021 (N_6021,N_2164,N_1000);
xor U6022 (N_6022,N_325,N_2664);
nor U6023 (N_6023,N_2418,N_2816);
nand U6024 (N_6024,N_1549,N_1633);
nor U6025 (N_6025,N_762,N_371);
and U6026 (N_6026,N_706,N_2527);
or U6027 (N_6027,N_2707,N_720);
and U6028 (N_6028,N_553,N_2938);
and U6029 (N_6029,N_565,N_3085);
nand U6030 (N_6030,N_1144,N_2725);
nor U6031 (N_6031,N_812,N_844);
nor U6032 (N_6032,N_2483,N_453);
xor U6033 (N_6033,N_2739,N_1716);
xnor U6034 (N_6034,N_2893,N_180);
and U6035 (N_6035,N_2634,N_380);
or U6036 (N_6036,N_43,N_2796);
and U6037 (N_6037,N_1191,N_2243);
nor U6038 (N_6038,N_1328,N_2611);
nand U6039 (N_6039,N_2775,N_1104);
and U6040 (N_6040,N_2984,N_700);
nand U6041 (N_6041,N_2055,N_3053);
nand U6042 (N_6042,N_418,N_342);
nor U6043 (N_6043,N_1617,N_2037);
or U6044 (N_6044,N_2428,N_2643);
or U6045 (N_6045,N_2690,N_64);
and U6046 (N_6046,N_1269,N_947);
and U6047 (N_6047,N_1096,N_728);
nand U6048 (N_6048,N_3097,N_71);
nor U6049 (N_6049,N_3104,N_2906);
or U6050 (N_6050,N_1465,N_3029);
xnor U6051 (N_6051,N_2929,N_1726);
xor U6052 (N_6052,N_1411,N_242);
or U6053 (N_6053,N_454,N_2042);
xor U6054 (N_6054,N_3066,N_1679);
nor U6055 (N_6055,N_71,N_865);
nand U6056 (N_6056,N_2509,N_2828);
and U6057 (N_6057,N_1455,N_303);
and U6058 (N_6058,N_2664,N_339);
nor U6059 (N_6059,N_316,N_77);
nand U6060 (N_6060,N_1339,N_554);
xor U6061 (N_6061,N_1366,N_891);
nand U6062 (N_6062,N_532,N_1257);
nand U6063 (N_6063,N_979,N_621);
xor U6064 (N_6064,N_1059,N_1529);
and U6065 (N_6065,N_3076,N_2448);
and U6066 (N_6066,N_1590,N_1347);
nor U6067 (N_6067,N_2233,N_2361);
nand U6068 (N_6068,N_585,N_2471);
or U6069 (N_6069,N_2403,N_817);
and U6070 (N_6070,N_545,N_1868);
and U6071 (N_6071,N_2858,N_3090);
or U6072 (N_6072,N_263,N_1811);
and U6073 (N_6073,N_3106,N_61);
nor U6074 (N_6074,N_2649,N_1925);
nand U6075 (N_6075,N_3111,N_1260);
xor U6076 (N_6076,N_1173,N_2923);
nor U6077 (N_6077,N_759,N_2226);
and U6078 (N_6078,N_1486,N_1342);
and U6079 (N_6079,N_1166,N_1096);
nor U6080 (N_6080,N_1310,N_1832);
xor U6081 (N_6081,N_408,N_445);
nor U6082 (N_6082,N_2113,N_804);
xor U6083 (N_6083,N_274,N_2805);
xor U6084 (N_6084,N_1952,N_2354);
and U6085 (N_6085,N_948,N_2270);
and U6086 (N_6086,N_2672,N_2113);
nand U6087 (N_6087,N_2408,N_1756);
or U6088 (N_6088,N_2931,N_2731);
nor U6089 (N_6089,N_603,N_360);
nor U6090 (N_6090,N_1755,N_1860);
nand U6091 (N_6091,N_2512,N_226);
xor U6092 (N_6092,N_1801,N_1182);
nand U6093 (N_6093,N_610,N_461);
xnor U6094 (N_6094,N_1044,N_1145);
nand U6095 (N_6095,N_1615,N_1833);
nand U6096 (N_6096,N_49,N_811);
nand U6097 (N_6097,N_636,N_97);
and U6098 (N_6098,N_2112,N_2352);
and U6099 (N_6099,N_2266,N_1666);
or U6100 (N_6100,N_386,N_570);
or U6101 (N_6101,N_2973,N_2765);
and U6102 (N_6102,N_209,N_602);
nor U6103 (N_6103,N_1176,N_2870);
or U6104 (N_6104,N_690,N_2270);
nand U6105 (N_6105,N_2506,N_186);
nand U6106 (N_6106,N_2189,N_700);
or U6107 (N_6107,N_1017,N_1548);
and U6108 (N_6108,N_720,N_134);
or U6109 (N_6109,N_1574,N_1616);
xor U6110 (N_6110,N_49,N_766);
xnor U6111 (N_6111,N_1737,N_1209);
nor U6112 (N_6112,N_1258,N_1644);
xor U6113 (N_6113,N_583,N_161);
nand U6114 (N_6114,N_1280,N_2031);
nor U6115 (N_6115,N_3035,N_497);
and U6116 (N_6116,N_2265,N_1644);
nor U6117 (N_6117,N_2044,N_1999);
nand U6118 (N_6118,N_18,N_1664);
nand U6119 (N_6119,N_931,N_1216);
and U6120 (N_6120,N_968,N_2181);
xor U6121 (N_6121,N_1259,N_50);
nor U6122 (N_6122,N_361,N_533);
and U6123 (N_6123,N_2222,N_0);
xnor U6124 (N_6124,N_2570,N_1538);
nor U6125 (N_6125,N_2059,N_3123);
or U6126 (N_6126,N_2009,N_740);
xor U6127 (N_6127,N_1752,N_2111);
or U6128 (N_6128,N_1976,N_3043);
nor U6129 (N_6129,N_2396,N_505);
and U6130 (N_6130,N_2105,N_2457);
nor U6131 (N_6131,N_3064,N_1361);
and U6132 (N_6132,N_1287,N_2382);
nor U6133 (N_6133,N_33,N_691);
nor U6134 (N_6134,N_455,N_1006);
nand U6135 (N_6135,N_3052,N_1171);
xor U6136 (N_6136,N_1692,N_99);
nand U6137 (N_6137,N_2557,N_2803);
and U6138 (N_6138,N_2979,N_842);
or U6139 (N_6139,N_321,N_2230);
nor U6140 (N_6140,N_114,N_2158);
xor U6141 (N_6141,N_2658,N_2859);
nor U6142 (N_6142,N_2437,N_1419);
nor U6143 (N_6143,N_202,N_598);
nand U6144 (N_6144,N_1360,N_3001);
nor U6145 (N_6145,N_564,N_2662);
and U6146 (N_6146,N_2557,N_1762);
and U6147 (N_6147,N_1454,N_1267);
and U6148 (N_6148,N_466,N_2164);
or U6149 (N_6149,N_343,N_576);
or U6150 (N_6150,N_678,N_1573);
and U6151 (N_6151,N_2337,N_895);
or U6152 (N_6152,N_737,N_1789);
or U6153 (N_6153,N_2365,N_2305);
nor U6154 (N_6154,N_1719,N_986);
nand U6155 (N_6155,N_1724,N_1424);
and U6156 (N_6156,N_2441,N_813);
nor U6157 (N_6157,N_1829,N_1396);
nand U6158 (N_6158,N_1805,N_2477);
nor U6159 (N_6159,N_1187,N_1456);
xor U6160 (N_6160,N_2589,N_22);
xor U6161 (N_6161,N_1724,N_356);
nor U6162 (N_6162,N_1636,N_1148);
and U6163 (N_6163,N_1618,N_2899);
and U6164 (N_6164,N_1346,N_869);
nand U6165 (N_6165,N_2076,N_2557);
and U6166 (N_6166,N_1709,N_1096);
xor U6167 (N_6167,N_2198,N_148);
nand U6168 (N_6168,N_113,N_2230);
xor U6169 (N_6169,N_19,N_1559);
or U6170 (N_6170,N_848,N_2094);
nand U6171 (N_6171,N_2233,N_1214);
and U6172 (N_6172,N_2430,N_2915);
or U6173 (N_6173,N_1290,N_2281);
xor U6174 (N_6174,N_986,N_2072);
or U6175 (N_6175,N_2379,N_1454);
or U6176 (N_6176,N_1355,N_1730);
nand U6177 (N_6177,N_2424,N_573);
nand U6178 (N_6178,N_340,N_2736);
or U6179 (N_6179,N_417,N_1725);
nand U6180 (N_6180,N_1939,N_2903);
nor U6181 (N_6181,N_1881,N_1427);
or U6182 (N_6182,N_2244,N_1361);
xnor U6183 (N_6183,N_2582,N_1875);
nor U6184 (N_6184,N_1976,N_1159);
and U6185 (N_6185,N_2851,N_952);
nor U6186 (N_6186,N_1937,N_1228);
or U6187 (N_6187,N_1914,N_2836);
xor U6188 (N_6188,N_1994,N_1471);
nor U6189 (N_6189,N_388,N_862);
and U6190 (N_6190,N_391,N_2031);
xnor U6191 (N_6191,N_1576,N_1446);
nor U6192 (N_6192,N_1294,N_1370);
nor U6193 (N_6193,N_2853,N_1858);
or U6194 (N_6194,N_4,N_3112);
nor U6195 (N_6195,N_1096,N_1615);
nor U6196 (N_6196,N_805,N_1784);
xnor U6197 (N_6197,N_2069,N_671);
nor U6198 (N_6198,N_1627,N_840);
nor U6199 (N_6199,N_2235,N_2560);
nor U6200 (N_6200,N_2498,N_376);
or U6201 (N_6201,N_2429,N_2193);
or U6202 (N_6202,N_3052,N_2146);
nor U6203 (N_6203,N_1917,N_1773);
xor U6204 (N_6204,N_847,N_2799);
nand U6205 (N_6205,N_2923,N_150);
xor U6206 (N_6206,N_1524,N_237);
and U6207 (N_6207,N_1612,N_1669);
or U6208 (N_6208,N_3048,N_231);
xnor U6209 (N_6209,N_1076,N_1499);
xor U6210 (N_6210,N_423,N_1526);
or U6211 (N_6211,N_2990,N_999);
nand U6212 (N_6212,N_456,N_183);
xnor U6213 (N_6213,N_2213,N_2879);
or U6214 (N_6214,N_2758,N_60);
and U6215 (N_6215,N_2455,N_1460);
and U6216 (N_6216,N_1702,N_2268);
nand U6217 (N_6217,N_1443,N_2251);
or U6218 (N_6218,N_2641,N_80);
nand U6219 (N_6219,N_2782,N_1010);
or U6220 (N_6220,N_408,N_760);
nor U6221 (N_6221,N_1423,N_3055);
nand U6222 (N_6222,N_1281,N_2535);
xnor U6223 (N_6223,N_2793,N_797);
xnor U6224 (N_6224,N_560,N_2029);
xnor U6225 (N_6225,N_1752,N_1808);
xor U6226 (N_6226,N_2981,N_1599);
nand U6227 (N_6227,N_1701,N_73);
nor U6228 (N_6228,N_114,N_217);
and U6229 (N_6229,N_178,N_1185);
or U6230 (N_6230,N_984,N_636);
or U6231 (N_6231,N_1991,N_1728);
nand U6232 (N_6232,N_1066,N_1341);
nand U6233 (N_6233,N_1962,N_2413);
nand U6234 (N_6234,N_2871,N_1119);
xnor U6235 (N_6235,N_1750,N_2826);
or U6236 (N_6236,N_961,N_360);
xnor U6237 (N_6237,N_804,N_859);
and U6238 (N_6238,N_1876,N_319);
and U6239 (N_6239,N_1318,N_1640);
and U6240 (N_6240,N_2750,N_1658);
and U6241 (N_6241,N_2527,N_636);
or U6242 (N_6242,N_1553,N_1684);
nand U6243 (N_6243,N_101,N_3098);
nor U6244 (N_6244,N_2678,N_827);
or U6245 (N_6245,N_2551,N_2594);
nand U6246 (N_6246,N_1722,N_2168);
and U6247 (N_6247,N_3121,N_3026);
or U6248 (N_6248,N_2686,N_518);
nor U6249 (N_6249,N_73,N_3112);
nand U6250 (N_6250,N_4680,N_4971);
or U6251 (N_6251,N_4667,N_6086);
xor U6252 (N_6252,N_3920,N_5490);
and U6253 (N_6253,N_4157,N_4583);
xor U6254 (N_6254,N_3463,N_5095);
or U6255 (N_6255,N_5661,N_5254);
nor U6256 (N_6256,N_4325,N_4316);
or U6257 (N_6257,N_5064,N_4982);
nand U6258 (N_6258,N_5894,N_4349);
xor U6259 (N_6259,N_4653,N_4106);
nand U6260 (N_6260,N_5308,N_3706);
nand U6261 (N_6261,N_3255,N_4202);
and U6262 (N_6262,N_3814,N_5132);
and U6263 (N_6263,N_4035,N_3905);
nand U6264 (N_6264,N_3574,N_5443);
nand U6265 (N_6265,N_5334,N_4968);
and U6266 (N_6266,N_5524,N_5702);
xnor U6267 (N_6267,N_5548,N_5795);
xnor U6268 (N_6268,N_5311,N_5775);
nor U6269 (N_6269,N_4016,N_5142);
nor U6270 (N_6270,N_4387,N_5350);
and U6271 (N_6271,N_3151,N_3800);
nor U6272 (N_6272,N_4203,N_5750);
or U6273 (N_6273,N_4489,N_5836);
nand U6274 (N_6274,N_4439,N_5258);
nand U6275 (N_6275,N_5442,N_5186);
and U6276 (N_6276,N_4189,N_4878);
or U6277 (N_6277,N_6197,N_5358);
xor U6278 (N_6278,N_4624,N_3392);
and U6279 (N_6279,N_4223,N_5454);
xnor U6280 (N_6280,N_4039,N_4314);
xor U6281 (N_6281,N_6191,N_3939);
or U6282 (N_6282,N_6174,N_3628);
nor U6283 (N_6283,N_4412,N_4527);
nand U6284 (N_6284,N_3139,N_4509);
xnor U6285 (N_6285,N_3481,N_4603);
xnor U6286 (N_6286,N_4111,N_3619);
nand U6287 (N_6287,N_3368,N_5204);
or U6288 (N_6288,N_5387,N_3684);
xor U6289 (N_6289,N_4083,N_6007);
or U6290 (N_6290,N_5944,N_5847);
nor U6291 (N_6291,N_4249,N_5874);
nor U6292 (N_6292,N_3710,N_3325);
and U6293 (N_6293,N_3835,N_3329);
xor U6294 (N_6294,N_3885,N_5299);
or U6295 (N_6295,N_5042,N_4540);
or U6296 (N_6296,N_4415,N_5351);
nor U6297 (N_6297,N_3522,N_4569);
nor U6298 (N_6298,N_5079,N_4827);
nor U6299 (N_6299,N_3896,N_3491);
xnor U6300 (N_6300,N_5901,N_5316);
and U6301 (N_6301,N_3848,N_3185);
or U6302 (N_6302,N_4721,N_4462);
xnor U6303 (N_6303,N_3761,N_4405);
nand U6304 (N_6304,N_3886,N_4816);
nor U6305 (N_6305,N_3948,N_5958);
nor U6306 (N_6306,N_5029,N_4551);
xnor U6307 (N_6307,N_4262,N_5163);
nor U6308 (N_6308,N_4863,N_4438);
nand U6309 (N_6309,N_6018,N_4440);
or U6310 (N_6310,N_5943,N_4549);
nand U6311 (N_6311,N_3488,N_3916);
xor U6312 (N_6312,N_6024,N_3533);
nor U6313 (N_6313,N_5536,N_3798);
or U6314 (N_6314,N_4781,N_4080);
or U6315 (N_6315,N_4972,N_4825);
nand U6316 (N_6316,N_4801,N_5066);
nand U6317 (N_6317,N_3371,N_3564);
nor U6318 (N_6318,N_3213,N_3793);
and U6319 (N_6319,N_4796,N_5229);
and U6320 (N_6320,N_4174,N_3446);
nor U6321 (N_6321,N_3892,N_4764);
and U6322 (N_6322,N_3356,N_4402);
nor U6323 (N_6323,N_6234,N_4390);
and U6324 (N_6324,N_3223,N_6222);
nand U6325 (N_6325,N_6240,N_4485);
nor U6326 (N_6326,N_4498,N_4430);
nand U6327 (N_6327,N_3526,N_5113);
nor U6328 (N_6328,N_4678,N_4280);
and U6329 (N_6329,N_4924,N_4885);
nand U6330 (N_6330,N_4564,N_4115);
and U6331 (N_6331,N_5125,N_3869);
xnor U6332 (N_6332,N_3182,N_5551);
nor U6333 (N_6333,N_3958,N_5920);
or U6334 (N_6334,N_4619,N_4759);
and U6335 (N_6335,N_5354,N_5276);
nor U6336 (N_6336,N_3842,N_6134);
nand U6337 (N_6337,N_5057,N_4058);
xnor U6338 (N_6338,N_5124,N_5205);
and U6339 (N_6339,N_3521,N_3246);
nor U6340 (N_6340,N_5019,N_4938);
or U6341 (N_6341,N_5882,N_4481);
or U6342 (N_6342,N_4589,N_4451);
xor U6343 (N_6343,N_4196,N_3999);
nand U6344 (N_6344,N_5723,N_5245);
xor U6345 (N_6345,N_3895,N_4735);
and U6346 (N_6346,N_4985,N_6047);
or U6347 (N_6347,N_3668,N_4154);
and U6348 (N_6348,N_5459,N_3728);
xnor U6349 (N_6349,N_5889,N_4719);
nor U6350 (N_6350,N_3161,N_3423);
xnor U6351 (N_6351,N_5456,N_4151);
nand U6352 (N_6352,N_4118,N_4399);
nand U6353 (N_6353,N_3499,N_4018);
or U6354 (N_6354,N_5198,N_5671);
nor U6355 (N_6355,N_4236,N_3157);
xnor U6356 (N_6356,N_4665,N_5699);
xor U6357 (N_6357,N_4534,N_3769);
nor U6358 (N_6358,N_3860,N_4024);
and U6359 (N_6359,N_3959,N_3303);
and U6360 (N_6360,N_3688,N_5626);
or U6361 (N_6361,N_6224,N_5462);
or U6362 (N_6362,N_3301,N_3504);
or U6363 (N_6363,N_4817,N_3682);
or U6364 (N_6364,N_4561,N_3782);
nand U6365 (N_6365,N_6182,N_4255);
nor U6366 (N_6366,N_5323,N_5252);
xnor U6367 (N_6367,N_6011,N_4932);
and U6368 (N_6368,N_5578,N_3722);
xor U6369 (N_6369,N_4260,N_6040);
and U6370 (N_6370,N_3954,N_4282);
nand U6371 (N_6371,N_4826,N_5213);
nand U6372 (N_6372,N_5261,N_5195);
xor U6373 (N_6373,N_4431,N_3679);
nor U6374 (N_6374,N_5729,N_5785);
and U6375 (N_6375,N_4297,N_6218);
or U6376 (N_6376,N_3426,N_5914);
and U6377 (N_6377,N_4342,N_3808);
xnor U6378 (N_6378,N_3512,N_4284);
nor U6379 (N_6379,N_6150,N_5864);
nand U6380 (N_6380,N_4334,N_5848);
or U6381 (N_6381,N_4171,N_3334);
nor U6382 (N_6382,N_6121,N_5881);
nand U6383 (N_6383,N_3134,N_3695);
nand U6384 (N_6384,N_5869,N_5022);
xor U6385 (N_6385,N_3340,N_3984);
and U6386 (N_6386,N_5556,N_5405);
and U6387 (N_6387,N_4013,N_5660);
or U6388 (N_6388,N_3534,N_3353);
or U6389 (N_6389,N_3751,N_4285);
or U6390 (N_6390,N_5087,N_5784);
or U6391 (N_6391,N_3432,N_4696);
or U6392 (N_6392,N_3511,N_4020);
and U6393 (N_6393,N_6177,N_4537);
and U6394 (N_6394,N_5497,N_3830);
xnor U6395 (N_6395,N_5840,N_4898);
or U6396 (N_6396,N_5967,N_3925);
or U6397 (N_6397,N_3600,N_5709);
nor U6398 (N_6398,N_3639,N_5046);
or U6399 (N_6399,N_5054,N_3897);
and U6400 (N_6400,N_3322,N_5665);
xor U6401 (N_6401,N_4046,N_5515);
nand U6402 (N_6402,N_4882,N_5475);
and U6403 (N_6403,N_5724,N_6242);
nand U6404 (N_6404,N_4650,N_3545);
nor U6405 (N_6405,N_5557,N_3215);
xor U6406 (N_6406,N_6032,N_5169);
xnor U6407 (N_6407,N_5071,N_4194);
xor U6408 (N_6408,N_3713,N_4628);
nor U6409 (N_6409,N_3376,N_5588);
and U6410 (N_6410,N_5994,N_4277);
nand U6411 (N_6411,N_3396,N_4948);
or U6412 (N_6412,N_3256,N_6084);
nor U6413 (N_6413,N_3456,N_3549);
or U6414 (N_6414,N_5838,N_4598);
and U6415 (N_6415,N_4553,N_5814);
nor U6416 (N_6416,N_6217,N_5867);
nor U6417 (N_6417,N_3765,N_4069);
nor U6418 (N_6418,N_5675,N_3351);
nor U6419 (N_6419,N_3384,N_5008);
nand U6420 (N_6420,N_3703,N_6168);
xor U6421 (N_6421,N_4208,N_6066);
and U6422 (N_6422,N_3757,N_5689);
nand U6423 (N_6423,N_5286,N_5324);
nand U6424 (N_6424,N_5432,N_3516);
or U6425 (N_6425,N_4011,N_3982);
xor U6426 (N_6426,N_5266,N_4158);
or U6427 (N_6427,N_6090,N_5826);
nor U6428 (N_6428,N_5230,N_5346);
and U6429 (N_6429,N_3324,N_5649);
nand U6430 (N_6430,N_5232,N_4471);
and U6431 (N_6431,N_3160,N_4045);
and U6432 (N_6432,N_5484,N_4067);
or U6433 (N_6433,N_4579,N_5282);
and U6434 (N_6434,N_6227,N_3261);
xor U6435 (N_6435,N_4596,N_5651);
nor U6436 (N_6436,N_4983,N_4450);
and U6437 (N_6437,N_5612,N_5220);
nand U6438 (N_6438,N_4261,N_5973);
or U6439 (N_6439,N_5221,N_3854);
and U6440 (N_6440,N_5818,N_5005);
xnor U6441 (N_6441,N_3727,N_4522);
or U6442 (N_6442,N_3667,N_5604);
and U6443 (N_6443,N_5440,N_3462);
nand U6444 (N_6444,N_5104,N_5697);
and U6445 (N_6445,N_3152,N_4986);
xor U6446 (N_6446,N_5883,N_4144);
nand U6447 (N_6447,N_4312,N_3572);
xor U6448 (N_6448,N_4946,N_5152);
or U6449 (N_6449,N_4516,N_5381);
and U6450 (N_6450,N_3225,N_4818);
nor U6451 (N_6451,N_5957,N_3956);
and U6452 (N_6452,N_4183,N_4793);
or U6453 (N_6453,N_4164,N_5806);
xor U6454 (N_6454,N_3767,N_4857);
nor U6455 (N_6455,N_5929,N_6035);
nand U6456 (N_6456,N_5561,N_5128);
xnor U6457 (N_6457,N_3887,N_5614);
and U6458 (N_6458,N_5802,N_4404);
and U6459 (N_6459,N_5747,N_5117);
xnor U6460 (N_6460,N_4211,N_6152);
nor U6461 (N_6461,N_5295,N_4259);
and U6462 (N_6462,N_3654,N_4695);
nand U6463 (N_6463,N_4469,N_3269);
xor U6464 (N_6464,N_5518,N_3715);
xnor U6465 (N_6465,N_6194,N_5068);
nand U6466 (N_6466,N_5255,N_5341);
nand U6467 (N_6467,N_5584,N_4022);
nor U6468 (N_6468,N_3657,N_3699);
nand U6469 (N_6469,N_5954,N_5373);
nand U6470 (N_6470,N_3485,N_4820);
nor U6471 (N_6471,N_6235,N_3228);
xor U6472 (N_6472,N_5922,N_5568);
xor U6473 (N_6473,N_5242,N_6188);
xor U6474 (N_6474,N_4251,N_5167);
and U6475 (N_6475,N_4877,N_6204);
and U6476 (N_6476,N_6102,N_6119);
xnor U6477 (N_6477,N_3541,N_6097);
xor U6478 (N_6478,N_5344,N_5051);
or U6479 (N_6479,N_5892,N_5099);
or U6480 (N_6480,N_3853,N_4136);
nand U6481 (N_6481,N_5366,N_4830);
nor U6482 (N_6482,N_3764,N_3788);
or U6483 (N_6483,N_3821,N_5809);
and U6484 (N_6484,N_5160,N_3841);
nor U6485 (N_6485,N_3746,N_3467);
nor U6486 (N_6486,N_3955,N_4162);
or U6487 (N_6487,N_5940,N_4293);
and U6488 (N_6488,N_4751,N_4071);
xor U6489 (N_6489,N_3405,N_4864);
nor U6490 (N_6490,N_5240,N_4905);
and U6491 (N_6491,N_5203,N_3586);
xnor U6492 (N_6492,N_3929,N_4874);
nand U6493 (N_6493,N_3671,N_3336);
and U6494 (N_6494,N_3778,N_4386);
or U6495 (N_6495,N_3608,N_6172);
or U6496 (N_6496,N_5370,N_5359);
or U6497 (N_6497,N_6198,N_3293);
or U6498 (N_6498,N_4239,N_3655);
xor U6499 (N_6499,N_4178,N_6108);
xnor U6500 (N_6500,N_5445,N_3242);
and U6501 (N_6501,N_3431,N_3866);
or U6502 (N_6502,N_5131,N_6214);
nand U6503 (N_6503,N_5530,N_4831);
nor U6504 (N_6504,N_4021,N_5762);
or U6505 (N_6505,N_5768,N_3359);
nor U6506 (N_6506,N_6075,N_4576);
or U6507 (N_6507,N_3846,N_5942);
or U6508 (N_6508,N_5212,N_5711);
nor U6509 (N_6509,N_4992,N_6044);
or U6510 (N_6510,N_5457,N_5815);
nor U6511 (N_6511,N_4886,N_4682);
nor U6512 (N_6512,N_4423,N_3993);
nor U6513 (N_6513,N_4951,N_4879);
nand U6514 (N_6514,N_3579,N_3622);
xnor U6515 (N_6515,N_5663,N_4359);
or U6516 (N_6516,N_5368,N_5062);
nand U6517 (N_6517,N_3878,N_5494);
and U6518 (N_6518,N_5392,N_5021);
xor U6519 (N_6519,N_3643,N_5035);
and U6520 (N_6520,N_5790,N_6176);
xnor U6521 (N_6521,N_5791,N_6233);
or U6522 (N_6522,N_4833,N_3427);
nand U6523 (N_6523,N_5734,N_5356);
xor U6524 (N_6524,N_4432,N_5899);
nand U6525 (N_6525,N_4233,N_4687);
nor U6526 (N_6526,N_4466,N_5759);
or U6527 (N_6527,N_3128,N_3805);
xnor U6528 (N_6528,N_5946,N_5849);
xor U6529 (N_6529,N_5102,N_3683);
and U6530 (N_6530,N_4729,N_4588);
nand U6531 (N_6531,N_3637,N_5783);
xnor U6532 (N_6532,N_3973,N_5673);
nor U6533 (N_6533,N_3820,N_4281);
nor U6534 (N_6534,N_5306,N_3365);
and U6535 (N_6535,N_4774,N_6170);
or U6536 (N_6536,N_4899,N_5859);
nand U6537 (N_6537,N_5645,N_4704);
or U6538 (N_6538,N_4943,N_4843);
nand U6539 (N_6539,N_6023,N_4936);
nand U6540 (N_6540,N_6115,N_3164);
or U6541 (N_6541,N_4231,N_4274);
nor U6542 (N_6542,N_5602,N_5371);
xor U6543 (N_6543,N_5813,N_5285);
xor U6544 (N_6544,N_5406,N_3882);
nor U6545 (N_6545,N_6117,N_3864);
xnor U6546 (N_6546,N_5315,N_5260);
xnor U6547 (N_6547,N_3720,N_5599);
nor U6548 (N_6548,N_4889,N_5119);
xnor U6549 (N_6549,N_5329,N_4602);
and U6550 (N_6550,N_4959,N_4135);
and U6551 (N_6551,N_3749,N_3131);
nand U6552 (N_6552,N_4934,N_4989);
or U6553 (N_6553,N_5837,N_4548);
nand U6554 (N_6554,N_4963,N_5722);
or U6555 (N_6555,N_5577,N_5177);
nand U6556 (N_6556,N_5357,N_5969);
nand U6557 (N_6557,N_4378,N_3346);
and U6558 (N_6558,N_5644,N_4822);
nand U6559 (N_6559,N_4718,N_5992);
or U6560 (N_6560,N_3216,N_6226);
and U6561 (N_6561,N_3861,N_5120);
or U6562 (N_6562,N_5915,N_3507);
nor U6563 (N_6563,N_4110,N_5735);
nor U6564 (N_6564,N_5547,N_5294);
nor U6565 (N_6565,N_5433,N_4813);
nand U6566 (N_6566,N_4909,N_5179);
and U6567 (N_6567,N_5631,N_5707);
xnor U6568 (N_6568,N_4993,N_4988);
and U6569 (N_6569,N_5025,N_4317);
or U6570 (N_6570,N_6037,N_4321);
and U6571 (N_6571,N_4256,N_4949);
and U6572 (N_6572,N_5235,N_5620);
xnor U6573 (N_6573,N_3226,N_3287);
and U6574 (N_6574,N_6199,N_3898);
nor U6575 (N_6575,N_4790,N_3919);
and U6576 (N_6576,N_4383,N_5115);
or U6577 (N_6577,N_5118,N_3957);
nor U6578 (N_6578,N_6207,N_3232);
nand U6579 (N_6579,N_3424,N_4419);
xnor U6580 (N_6580,N_5710,N_4077);
or U6581 (N_6581,N_5372,N_5652);
nor U6582 (N_6582,N_6058,N_3294);
or U6583 (N_6583,N_4304,N_4368);
and U6584 (N_6584,N_5465,N_3525);
nand U6585 (N_6585,N_4005,N_3341);
or U6586 (N_6586,N_3941,N_4300);
nor U6587 (N_6587,N_6073,N_4829);
xnor U6588 (N_6588,N_3125,N_6062);
and U6589 (N_6589,N_3694,N_5540);
and U6590 (N_6590,N_3809,N_4453);
nor U6591 (N_6591,N_5581,N_5900);
nand U6592 (N_6592,N_3357,N_3961);
and U6593 (N_6593,N_3707,N_4320);
nand U6594 (N_6594,N_5844,N_6074);
nor U6595 (N_6595,N_3771,N_5478);
nor U6596 (N_6596,N_4961,N_3557);
and U6597 (N_6597,N_4927,N_5367);
or U6598 (N_6598,N_5448,N_3280);
nand U6599 (N_6599,N_3690,N_5298);
xor U6600 (N_6600,N_3460,N_5403);
nand U6601 (N_6601,N_6034,N_4814);
or U6602 (N_6602,N_4147,N_5793);
nor U6603 (N_6603,N_4313,N_6083);
nand U6604 (N_6604,N_5075,N_4710);
or U6605 (N_6605,N_6051,N_3502);
nor U6606 (N_6606,N_5634,N_3971);
nor U6607 (N_6607,N_3986,N_3593);
xor U6608 (N_6608,N_4715,N_4187);
nor U6609 (N_6609,N_3388,N_4240);
xnor U6610 (N_6610,N_5196,N_5538);
and U6611 (N_6611,N_4608,N_5932);
and U6612 (N_6612,N_5880,N_6022);
or U6613 (N_6613,N_5312,N_4273);
and U6614 (N_6614,N_5953,N_5017);
and U6615 (N_6615,N_6243,N_4858);
and U6616 (N_6616,N_3438,N_4031);
nand U6617 (N_6617,N_5126,N_3385);
and U6618 (N_6618,N_4488,N_4631);
nor U6619 (N_6619,N_4640,N_5045);
and U6620 (N_6620,N_3308,N_4424);
nor U6621 (N_6621,N_5617,N_4056);
nand U6622 (N_6622,N_3748,N_4875);
nand U6623 (N_6623,N_4844,N_3291);
and U6624 (N_6624,N_4230,N_3678);
and U6625 (N_6625,N_5486,N_3621);
nor U6626 (N_6626,N_5474,N_4351);
xor U6627 (N_6627,N_5917,N_3307);
or U6628 (N_6628,N_4605,N_6027);
and U6629 (N_6629,N_5730,N_5871);
and U6630 (N_6630,N_4305,N_5677);
xor U6631 (N_6631,N_5236,N_5326);
xnor U6632 (N_6632,N_5265,N_5646);
nor U6633 (N_6633,N_4894,N_6196);
nand U6634 (N_6634,N_4308,N_4769);
nand U6635 (N_6635,N_4819,N_4686);
nand U6636 (N_6636,N_4152,N_3791);
xor U6637 (N_6637,N_3740,N_4614);
nor U6638 (N_6638,N_5907,N_3188);
nand U6639 (N_6639,N_4703,N_3561);
and U6640 (N_6640,N_6205,N_3449);
and U6641 (N_6641,N_3802,N_3270);
nor U6642 (N_6642,N_4955,N_4768);
nand U6643 (N_6643,N_4684,N_3960);
xnor U6644 (N_6644,N_4384,N_4190);
nand U6645 (N_6645,N_3172,N_5077);
nand U6646 (N_6646,N_4445,N_6057);
nand U6647 (N_6647,N_4900,N_3349);
nor U6648 (N_6648,N_5292,N_5909);
and U6649 (N_6649,N_3949,N_4268);
nor U6650 (N_6650,N_3493,N_4647);
nand U6651 (N_6651,N_3163,N_5253);
nand U6652 (N_6652,N_5480,N_6000);
nor U6653 (N_6653,N_5704,N_3144);
nor U6654 (N_6654,N_4966,N_5185);
or U6655 (N_6655,N_5267,N_3487);
xnor U6656 (N_6656,N_5239,N_3738);
nor U6657 (N_6657,N_3320,N_4141);
xnor U6658 (N_6658,N_4129,N_5580);
xnor U6659 (N_6659,N_5703,N_3286);
or U6660 (N_6660,N_5855,N_4165);
and U6661 (N_6661,N_5216,N_5168);
xnor U6662 (N_6662,N_3165,N_4573);
and U6663 (N_6663,N_5964,N_5352);
xor U6664 (N_6664,N_5107,N_6021);
and U6665 (N_6665,N_5879,N_3935);
xor U6666 (N_6666,N_5514,N_6089);
or U6667 (N_6667,N_5569,N_3482);
or U6668 (N_6668,N_3147,N_4860);
and U6669 (N_6669,N_4738,N_4693);
and U6670 (N_6670,N_4287,N_3855);
nor U6671 (N_6671,N_6165,N_5829);
xnor U6672 (N_6672,N_4101,N_3776);
xnor U6673 (N_6673,N_3563,N_6181);
and U6674 (N_6674,N_3209,N_5091);
nor U6675 (N_6675,N_4117,N_4558);
nor U6676 (N_6676,N_3410,N_4258);
and U6677 (N_6677,N_3863,N_3772);
nand U6678 (N_6678,N_5165,N_3338);
xnor U6679 (N_6679,N_4195,N_3317);
and U6680 (N_6680,N_3179,N_3374);
or U6681 (N_6681,N_4995,N_3360);
nor U6682 (N_6682,N_3766,N_6179);
nand U6683 (N_6683,N_5476,N_4969);
nand U6684 (N_6684,N_5544,N_5714);
and U6685 (N_6685,N_4883,N_3989);
and U6686 (N_6686,N_5090,N_3590);
nand U6687 (N_6687,N_5106,N_4267);
nor U6688 (N_6688,N_3250,N_5184);
nand U6689 (N_6689,N_3180,N_3302);
and U6690 (N_6690,N_4395,N_4524);
xor U6691 (N_6691,N_5805,N_4168);
nand U6692 (N_6692,N_5803,N_3795);
nand U6693 (N_6693,N_5755,N_3605);
or U6694 (N_6694,N_4847,N_4007);
nand U6695 (N_6695,N_5846,N_4263);
xor U6696 (N_6696,N_5197,N_3581);
xor U6697 (N_6697,N_5629,N_4737);
nor U6698 (N_6698,N_3737,N_3646);
and U6699 (N_6699,N_4520,N_5962);
nand U6700 (N_6700,N_5789,N_5891);
nor U6701 (N_6701,N_4355,N_5166);
nor U6702 (N_6702,N_5310,N_3127);
nor U6703 (N_6703,N_4252,N_3260);
nand U6704 (N_6704,N_3430,N_6136);
nor U6705 (N_6705,N_3422,N_5794);
nand U6706 (N_6706,N_3344,N_5435);
nor U6707 (N_6707,N_3921,N_5419);
xnor U6708 (N_6708,N_4902,N_4322);
and U6709 (N_6709,N_5369,N_4473);
or U6710 (N_6710,N_3677,N_4023);
or U6711 (N_6711,N_4458,N_4414);
nor U6712 (N_6712,N_3570,N_5636);
xnor U6713 (N_6713,N_4926,N_5233);
or U6714 (N_6714,N_3254,N_3972);
nand U6715 (N_6715,N_5209,N_5136);
nand U6716 (N_6716,N_4246,N_5738);
xor U6717 (N_6717,N_4786,N_4149);
xor U6718 (N_6718,N_4627,N_4166);
and U6719 (N_6719,N_4798,N_5579);
nand U6720 (N_6720,N_6206,N_5774);
and U6721 (N_6721,N_4805,N_3580);
or U6722 (N_6722,N_3618,N_3296);
nor U6723 (N_6723,N_3816,N_5641);
and U6724 (N_6724,N_5741,N_5437);
and U6725 (N_6725,N_3859,N_6158);
nand U6726 (N_6726,N_5609,N_4760);
nor U6727 (N_6727,N_5420,N_5439);
xor U6728 (N_6728,N_4155,N_5458);
and U6729 (N_6729,N_4610,N_5016);
and U6730 (N_6730,N_3753,N_5975);
nand U6731 (N_6731,N_3942,N_4339);
and U6732 (N_6732,N_3790,N_3888);
xor U6733 (N_6733,N_3631,N_5746);
and U6734 (N_6734,N_3328,N_3966);
or U6735 (N_6735,N_6033,N_5244);
nor U6736 (N_6736,N_6178,N_5553);
or U6737 (N_6737,N_3355,N_3244);
nand U6738 (N_6738,N_4787,N_4783);
and U6739 (N_6739,N_4919,N_4767);
xor U6740 (N_6740,N_4213,N_3873);
nand U6741 (N_6741,N_4958,N_5309);
or U6742 (N_6742,N_5274,N_3691);
nand U6743 (N_6743,N_4538,N_5382);
nand U6744 (N_6744,N_3718,N_3400);
nor U6745 (N_6745,N_3797,N_3983);
nor U6746 (N_6746,N_5332,N_3364);
or U6747 (N_6747,N_6050,N_3506);
xor U6748 (N_6748,N_6146,N_5876);
nand U6749 (N_6749,N_3466,N_4269);
xnor U6750 (N_6750,N_5215,N_3568);
or U6751 (N_6751,N_5401,N_5006);
or U6752 (N_6752,N_5955,N_3451);
and U6753 (N_6753,N_5526,N_5903);
and U6754 (N_6754,N_4075,N_4091);
and U6755 (N_6755,N_6085,N_4750);
or U6756 (N_6756,N_3285,N_4517);
xnor U6757 (N_6757,N_3497,N_3810);
nand U6758 (N_6758,N_4933,N_5549);
nand U6759 (N_6759,N_4884,N_3652);
xor U6760 (N_6760,N_4761,N_3343);
or U6761 (N_6761,N_4657,N_5831);
or U6762 (N_6762,N_5491,N_5362);
nor U6763 (N_6763,N_5187,N_3265);
and U6764 (N_6764,N_4109,N_4809);
nor U6765 (N_6765,N_5788,N_6025);
nand U6766 (N_6766,N_5503,N_3465);
and U6767 (N_6767,N_3697,N_5009);
xnor U6768 (N_6768,N_3141,N_4662);
nor U6769 (N_6769,N_3730,N_5269);
xor U6770 (N_6770,N_3704,N_3434);
nand U6771 (N_6771,N_3890,N_4341);
or U6772 (N_6772,N_3535,N_5182);
nor U6773 (N_6773,N_3552,N_5007);
nor U6774 (N_6774,N_4594,N_4116);
nand U6775 (N_6775,N_3378,N_3923);
and U6776 (N_6776,N_3596,N_6093);
nor U6777 (N_6777,N_5289,N_3756);
or U6778 (N_6778,N_4965,N_3907);
or U6779 (N_6779,N_5725,N_3473);
and U6780 (N_6780,N_6041,N_3803);
xor U6781 (N_6781,N_5947,N_3943);
xnor U6782 (N_6782,N_4570,N_4775);
nand U6783 (N_6783,N_5749,N_4294);
or U6784 (N_6784,N_3539,N_4229);
nand U6785 (N_6785,N_5015,N_5317);
xnor U6786 (N_6786,N_5905,N_3967);
or U6787 (N_6787,N_6052,N_3509);
xor U6788 (N_6788,N_3616,N_3201);
nand U6789 (N_6789,N_5180,N_5687);
or U6790 (N_6790,N_4501,N_5110);
nor U6791 (N_6791,N_4301,N_6038);
xnor U6792 (N_6792,N_6163,N_4379);
nand U6793 (N_6793,N_4890,N_6127);
and U6794 (N_6794,N_4177,N_3833);
xor U6795 (N_6795,N_5679,N_5094);
or U6796 (N_6796,N_5979,N_3229);
nor U6797 (N_6797,N_5098,N_5500);
nand U6798 (N_6798,N_6036,N_3447);
and U6799 (N_6799,N_5558,N_4601);
nand U6800 (N_6800,N_5823,N_5694);
xor U6801 (N_6801,N_5069,N_5933);
nor U6802 (N_6802,N_3649,N_3632);
or U6803 (N_6803,N_5930,N_4915);
nand U6804 (N_6804,N_3700,N_4757);
or U6805 (N_6805,N_3382,N_5380);
or U6806 (N_6806,N_5632,N_4571);
nand U6807 (N_6807,N_6118,N_4871);
nand U6808 (N_6808,N_4743,N_6123);
or U6809 (N_6809,N_3458,N_6081);
xnor U6810 (N_6810,N_4398,N_3146);
and U6811 (N_6811,N_4523,N_4426);
or U6812 (N_6812,N_4868,N_5997);
nand U6813 (N_6813,N_3309,N_5504);
nor U6814 (N_6814,N_5527,N_5379);
xnor U6815 (N_6815,N_3316,N_5429);
xor U6816 (N_6816,N_4870,N_5345);
nor U6817 (N_6817,N_5686,N_3498);
nor U6818 (N_6818,N_4169,N_5934);
and U6819 (N_6819,N_6210,N_5134);
or U6820 (N_6820,N_3834,N_5228);
and U6821 (N_6821,N_5541,N_5586);
and U6822 (N_6822,N_4480,N_4047);
and U6823 (N_6823,N_3183,N_3236);
and U6824 (N_6824,N_5231,N_3413);
nand U6825 (N_6825,N_5479,N_3996);
and U6826 (N_6826,N_3598,N_4791);
nand U6827 (N_6827,N_4367,N_5904);
nor U6828 (N_6828,N_4725,N_6185);
or U6829 (N_6829,N_4505,N_3175);
or U6830 (N_6830,N_5400,N_3965);
or U6831 (N_6831,N_3673,N_5191);
xor U6832 (N_6832,N_5928,N_5175);
or U6833 (N_6833,N_5648,N_5246);
nor U6834 (N_6834,N_4150,N_4974);
nor U6835 (N_6835,N_4228,N_3962);
or U6836 (N_6836,N_5241,N_5885);
and U6837 (N_6837,N_3674,N_4407);
xnor U6838 (N_6838,N_5960,N_5669);
xor U6839 (N_6839,N_6230,N_4952);
nand U6840 (N_6840,N_5890,N_3726);
nor U6841 (N_6841,N_5845,N_5833);
or U6842 (N_6842,N_3947,N_3208);
xor U6843 (N_6843,N_5452,N_4089);
xnor U6844 (N_6844,N_4265,N_3398);
nor U6845 (N_6845,N_4506,N_5726);
and U6846 (N_6846,N_4173,N_4145);
nand U6847 (N_6847,N_3559,N_3288);
xor U6848 (N_6848,N_5112,N_5966);
nor U6849 (N_6849,N_4586,N_5081);
xnor U6850 (N_6850,N_4618,N_4338);
nor U6851 (N_6851,N_3658,N_3211);
nand U6852 (N_6852,N_3744,N_4357);
nand U6853 (N_6853,N_3856,N_5576);
and U6854 (N_6854,N_6125,N_3192);
or U6855 (N_6855,N_5083,N_4073);
nand U6856 (N_6856,N_4418,N_6048);
xor U6857 (N_6857,N_5528,N_5884);
nand U6858 (N_6858,N_5619,N_6190);
nand U6859 (N_6859,N_4036,N_4731);
nor U6860 (N_6860,N_5451,N_4954);
or U6861 (N_6861,N_4241,N_3997);
or U6862 (N_6862,N_3537,N_4253);
nand U6863 (N_6863,N_5060,N_4510);
nand U6864 (N_6864,N_3573,N_4507);
nand U6865 (N_6865,N_4937,N_4944);
xnor U6866 (N_6866,N_4443,N_5206);
nor U6867 (N_6867,N_4138,N_4595);
nand U6868 (N_6868,N_3492,N_4872);
and U6869 (N_6869,N_4747,N_3200);
nor U6870 (N_6870,N_4771,N_3445);
or U6871 (N_6871,N_5571,N_4499);
and U6872 (N_6872,N_5361,N_4609);
nor U6873 (N_6873,N_5301,N_4393);
or U6874 (N_6874,N_3259,N_5630);
and U6875 (N_6875,N_3661,N_5529);
nand U6876 (N_6876,N_3436,N_3263);
nor U6877 (N_6877,N_5193,N_5348);
or U6878 (N_6878,N_3138,N_5798);
or U6879 (N_6879,N_5611,N_3304);
xor U6880 (N_6880,N_3524,N_3331);
xnor U6881 (N_6881,N_4120,N_4072);
xnor U6882 (N_6882,N_3785,N_3932);
nand U6883 (N_6883,N_4513,N_5485);
nor U6884 (N_6884,N_3926,N_4690);
and U6885 (N_6885,N_6137,N_5516);
or U6886 (N_6886,N_5383,N_5866);
nand U6887 (N_6887,N_3305,N_5336);
or U6888 (N_6888,N_4708,N_5302);
nor U6889 (N_6889,N_4235,N_5386);
and U6890 (N_6890,N_5583,N_5053);
nor U6891 (N_6891,N_3470,N_5293);
xor U6892 (N_6892,N_4688,N_3807);
and U6893 (N_6893,N_3312,N_3237);
nor U6894 (N_6894,N_4654,N_5415);
nand U6895 (N_6895,N_3933,N_5657);
xor U6896 (N_6896,N_3289,N_3532);
xnor U6897 (N_6897,N_5183,N_5926);
nor U6898 (N_6898,N_3571,N_3686);
nor U6899 (N_6899,N_3610,N_5918);
nor U6900 (N_6900,N_4176,N_3333);
nand U6901 (N_6901,N_4720,N_3725);
and U6902 (N_6902,N_6079,N_5375);
nand U6903 (N_6903,N_6076,N_3931);
or U6904 (N_6904,N_3543,N_5510);
nand U6905 (N_6905,N_5225,N_5002);
nand U6906 (N_6906,N_5978,N_4292);
xnor U6907 (N_6907,N_4180,N_5519);
xnor U6908 (N_6908,N_4699,N_3137);
xnor U6909 (N_6909,N_5539,N_4185);
xor U6910 (N_6910,N_3985,N_3173);
and U6911 (N_6911,N_3290,N_4560);
nor U6912 (N_6912,N_5248,N_4925);
or U6913 (N_6913,N_5720,N_4566);
or U6914 (N_6914,N_5407,N_4330);
or U6915 (N_6915,N_5404,N_3197);
xor U6916 (N_6916,N_5176,N_5273);
or U6917 (N_6917,N_4722,N_3812);
or U6918 (N_6918,N_3702,N_3372);
nor U6919 (N_6919,N_4343,N_6215);
or U6920 (N_6920,N_4795,N_3184);
nor U6921 (N_6921,N_4163,N_5399);
and U6922 (N_6922,N_6175,N_5048);
nor U6923 (N_6923,N_3397,N_3310);
xnor U6924 (N_6924,N_4289,N_4681);
nor U6925 (N_6925,N_5434,N_5656);
nor U6926 (N_6926,N_6148,N_5925);
nand U6927 (N_6927,N_5825,N_5270);
xor U6928 (N_6928,N_5692,N_4172);
nor U6929 (N_6929,N_4861,N_5897);
or U6930 (N_6930,N_5961,N_3421);
nand U6931 (N_6931,N_5014,N_5421);
or U6932 (N_6932,N_4403,N_3406);
xnor U6933 (N_6933,N_3448,N_3402);
or U6934 (N_6934,N_4859,N_3267);
and U6935 (N_6935,N_3453,N_3844);
and U6936 (N_6936,N_3441,N_3930);
nand U6937 (N_6937,N_4362,N_5446);
xor U6938 (N_6938,N_5719,N_5817);
and U6939 (N_6939,N_4051,N_4193);
xor U6940 (N_6940,N_3547,N_3851);
nand U6941 (N_6941,N_5397,N_4673);
nor U6942 (N_6942,N_4794,N_3528);
xnor U6943 (N_6943,N_6059,N_4804);
xor U6944 (N_6944,N_5149,N_4496);
xor U6945 (N_6945,N_6114,N_6193);
or U6946 (N_6946,N_4726,N_4901);
or U6947 (N_6947,N_5765,N_3205);
nand U6948 (N_6948,N_5314,N_3550);
or U6949 (N_6949,N_3784,N_4550);
nor U6950 (N_6950,N_4019,N_4494);
xor U6951 (N_6951,N_4380,N_4643);
xnor U6952 (N_6952,N_4264,N_4064);
nor U6953 (N_6953,N_5633,N_4812);
and U6954 (N_6954,N_3804,N_5893);
or U6955 (N_6955,N_3754,N_5695);
nor U6956 (N_6956,N_3604,N_3486);
and U6957 (N_6957,N_4048,N_4832);
or U6958 (N_6958,N_5171,N_3531);
nand U6959 (N_6959,N_4060,N_5467);
nand U6960 (N_6960,N_5347,N_5853);
nor U6961 (N_6961,N_5607,N_3934);
xor U6962 (N_6962,N_3159,N_5505);
and U6963 (N_6963,N_5562,N_5279);
nand U6964 (N_6964,N_4545,N_5986);
xnor U6965 (N_6965,N_4562,N_6220);
or U6966 (N_6966,N_4008,N_5878);
or U6967 (N_6967,N_4492,N_4401);
xnor U6968 (N_6968,N_4327,N_6019);
and U6969 (N_6969,N_5792,N_4087);
or U6970 (N_6970,N_5086,N_3944);
or U6971 (N_6971,N_3578,N_4978);
and U6972 (N_6972,N_5658,N_6238);
and U6973 (N_6973,N_5919,N_3544);
xor U6974 (N_6974,N_5650,N_4685);
xnor U6975 (N_6975,N_5003,N_5856);
and U6976 (N_6976,N_5801,N_3554);
nand U6977 (N_6977,N_3464,N_3420);
and U6978 (N_6978,N_3723,N_4433);
and U6979 (N_6979,N_3154,N_5659);
xnor U6980 (N_6980,N_5756,N_5464);
and U6981 (N_6981,N_6232,N_3249);
nand U6982 (N_6982,N_5628,N_3224);
nand U6983 (N_6983,N_3817,N_4392);
and U6984 (N_6984,N_3763,N_3373);
or U6985 (N_6985,N_5908,N_6147);
or U6986 (N_6986,N_5174,N_5036);
nand U6987 (N_6987,N_3323,N_4286);
xor U6988 (N_6988,N_3811,N_6078);
nor U6989 (N_6989,N_4838,N_4599);
nand U6990 (N_6990,N_5394,N_5249);
nand U6991 (N_6991,N_5761,N_4114);
and U6992 (N_6992,N_5574,N_3362);
nand U6993 (N_6993,N_5304,N_5477);
nor U6994 (N_6994,N_6069,N_3515);
nor U6995 (N_6995,N_5772,N_4425);
nor U6996 (N_6996,N_5374,N_4408);
xor U6997 (N_6997,N_5408,N_5565);
xor U6998 (N_6998,N_4706,N_3520);
nand U6999 (N_6999,N_3472,N_5453);
nand U7000 (N_7000,N_4616,N_5854);
xnor U7001 (N_7001,N_3783,N_5340);
xnor U7002 (N_7002,N_3476,N_5780);
and U7003 (N_7003,N_5898,N_4092);
xnor U7004 (N_7004,N_5088,N_5977);
xnor U7005 (N_7005,N_4808,N_5263);
nor U7006 (N_7006,N_5396,N_5776);
xor U7007 (N_7007,N_4869,N_6239);
nand U7008 (N_7008,N_3681,N_3626);
and U7009 (N_7009,N_5593,N_3850);
nor U7010 (N_7010,N_5868,N_3251);
nor U7011 (N_7011,N_6106,N_4800);
xor U7012 (N_7012,N_5506,N_3174);
and U7013 (N_7013,N_5012,N_5339);
xnor U7014 (N_7014,N_5281,N_5771);
nor U7015 (N_7015,N_5821,N_5618);
nor U7016 (N_7016,N_5861,N_4337);
nor U7017 (N_7017,N_5684,N_5123);
nand U7018 (N_7018,N_4906,N_4372);
or U7019 (N_7019,N_4724,N_5028);
and U7020 (N_7020,N_4454,N_4385);
or U7021 (N_7021,N_5201,N_4348);
nor U7022 (N_7022,N_3339,N_4784);
xnor U7023 (N_7023,N_4600,N_4962);
or U7024 (N_7024,N_4088,N_5389);
or U7025 (N_7025,N_3990,N_3221);
nor U7026 (N_7026,N_4474,N_3332);
nor U7027 (N_7027,N_3911,N_5038);
nor U7028 (N_7028,N_3428,N_5596);
and U7029 (N_7029,N_4345,N_3452);
nand U7030 (N_7030,N_4642,N_3739);
nor U7031 (N_7031,N_5272,N_5655);
nor U7032 (N_7032,N_5065,N_5981);
nor U7033 (N_7033,N_6216,N_4984);
xor U7034 (N_7034,N_3217,N_3130);
and U7035 (N_7035,N_5402,N_4170);
and U7036 (N_7036,N_4855,N_6096);
or U7037 (N_7037,N_3634,N_4788);
nand U7038 (N_7038,N_4659,N_5935);
nor U7039 (N_7039,N_3826,N_4713);
nor U7040 (N_7040,N_5804,N_5237);
xor U7041 (N_7041,N_5959,N_6248);
nand U7042 (N_7042,N_4973,N_4000);
or U7043 (N_7043,N_4104,N_4119);
and U7044 (N_7044,N_4622,N_5546);
xnor U7045 (N_7045,N_4333,N_4059);
nor U7046 (N_7046,N_4375,N_6124);
nand U7047 (N_7047,N_3779,N_3149);
nand U7048 (N_7048,N_4590,N_4668);
nand U7049 (N_7049,N_5325,N_5585);
nor U7050 (N_7050,N_4302,N_3393);
xnor U7051 (N_7051,N_4908,N_5319);
nor U7052 (N_7052,N_5024,N_4503);
nand U7053 (N_7053,N_4621,N_5690);
nor U7054 (N_7054,N_5461,N_3514);
nor U7055 (N_7055,N_4137,N_4346);
or U7056 (N_7056,N_5140,N_3822);
or U7057 (N_7057,N_3276,N_5084);
or U7058 (N_7058,N_5812,N_5983);
xnor U7059 (N_7059,N_5096,N_5322);
nand U7060 (N_7060,N_3978,N_3662);
xnor U7061 (N_7061,N_3140,N_4483);
or U7062 (N_7062,N_6002,N_4998);
xnor U7063 (N_7063,N_4428,N_6109);
nand U7064 (N_7064,N_5116,N_3190);
nor U7065 (N_7065,N_4002,N_5985);
xor U7066 (N_7066,N_3369,N_4126);
xnor U7067 (N_7067,N_4382,N_4782);
nand U7068 (N_7068,N_4777,N_5070);
and U7069 (N_7069,N_3577,N_4467);
xor U7070 (N_7070,N_4250,N_4922);
nand U7071 (N_7071,N_5318,N_5101);
and U7072 (N_7072,N_5906,N_6009);
xnor U7073 (N_7073,N_4648,N_4098);
xnor U7074 (N_7074,N_4295,N_4449);
and U7075 (N_7075,N_6043,N_5698);
and U7076 (N_7076,N_4465,N_3951);
xnor U7077 (N_7077,N_4409,N_4911);
xnor U7078 (N_7078,N_4096,N_4730);
nor U7079 (N_7079,N_5450,N_3459);
and U7080 (N_7080,N_5605,N_4736);
or U7081 (N_7081,N_4082,N_5037);
nand U7082 (N_7082,N_4037,N_5590);
xor U7083 (N_7083,N_5680,N_4361);
or U7084 (N_7084,N_4099,N_3976);
nand U7085 (N_7085,N_4369,N_4744);
or U7086 (N_7086,N_3773,N_3243);
nand U7087 (N_7087,N_5337,N_3644);
nand U7088 (N_7088,N_3529,N_4133);
or U7089 (N_7089,N_5639,N_5828);
xor U7090 (N_7090,N_4876,N_4139);
xor U7091 (N_7091,N_5135,N_5447);
xnor U7092 (N_7092,N_5436,N_5666);
nand U7093 (N_7093,N_5888,N_5059);
or U7094 (N_7094,N_5150,N_5748);
and U7095 (N_7095,N_4447,N_4207);
and U7096 (N_7096,N_4977,N_4531);
or U7097 (N_7097,N_4063,N_3629);
or U7098 (N_7098,N_3780,N_4856);
nand U7099 (N_7099,N_4200,N_4987);
or U7100 (N_7100,N_3852,N_3587);
nor U7101 (N_7101,N_4756,N_5208);
xor U7102 (N_7102,N_4698,N_6167);
nand U7103 (N_7103,N_3937,N_3927);
nand U7104 (N_7104,N_5970,N_4604);
nor U7105 (N_7105,N_4733,N_3158);
nand U7106 (N_7106,N_4270,N_5105);
or U7107 (N_7107,N_4417,N_5664);
nor U7108 (N_7108,N_3518,N_4004);
nor U7109 (N_7109,N_3602,N_5509);
nor U7110 (N_7110,N_5563,N_3991);
or U7111 (N_7111,N_4477,N_4778);
and U7112 (N_7112,N_5030,N_3177);
or U7113 (N_7113,N_6145,N_4543);
and U7114 (N_7114,N_5156,N_3567);
xnor U7115 (N_7115,N_4947,N_4518);
nand U7116 (N_7116,N_3575,N_3836);
or U7117 (N_7117,N_4220,N_3613);
nor U7118 (N_7118,N_4146,N_4991);
or U7119 (N_7119,N_3248,N_4219);
nand U7120 (N_7120,N_4705,N_5378);
and U7121 (N_7121,N_4606,N_3870);
and U7122 (N_7122,N_4310,N_3418);
or U7123 (N_7123,N_4460,N_4288);
nand U7124 (N_7124,N_5582,N_3714);
nand U7125 (N_7125,N_3204,N_3366);
nand U7126 (N_7126,N_6133,N_6042);
nand U7127 (N_7127,N_5441,N_5424);
xnor U7128 (N_7128,N_5567,N_5839);
or U7129 (N_7129,N_5870,N_3635);
xor U7130 (N_7130,N_5830,N_3741);
xor U7131 (N_7131,N_5533,N_4572);
or U7132 (N_7132,N_3900,N_5573);
xnor U7133 (N_7133,N_3214,N_5887);
and U7134 (N_7134,N_6173,N_6156);
xnor U7135 (N_7135,N_4749,N_3268);
and U7136 (N_7136,N_6180,N_5594);
and U7137 (N_7137,N_3663,N_5601);
and U7138 (N_7138,N_5770,N_5409);
xor U7139 (N_7139,N_4070,N_3721);
or U7140 (N_7140,N_4865,N_5753);
nor U7141 (N_7141,N_4429,N_3454);
nand U7142 (N_7142,N_5542,N_4085);
or U7143 (N_7143,N_5471,N_3945);
or U7144 (N_7144,N_5760,N_3917);
nand U7145 (N_7145,N_3136,N_6055);
and U7146 (N_7146,N_3517,N_4365);
nor U7147 (N_7147,N_3245,N_5395);
and U7148 (N_7148,N_6135,N_3712);
nand U7149 (N_7149,N_4084,N_4641);
xor U7150 (N_7150,N_5916,N_3789);
nor U7151 (N_7151,N_5027,N_5712);
nor U7152 (N_7152,N_4556,N_3212);
xnor U7153 (N_7153,N_4683,N_4873);
and U7154 (N_7154,N_3994,N_4806);
xnor U7155 (N_7155,N_5353,N_6151);
xor U7156 (N_7156,N_4611,N_4497);
or U7157 (N_7157,N_4309,N_5923);
nand U7158 (N_7158,N_4222,N_4242);
and U7159 (N_7159,N_4994,N_3591);
and U7160 (N_7160,N_6053,N_4612);
xnor U7161 (N_7161,N_5757,N_4842);
xor U7162 (N_7162,N_4525,N_4416);
xor U7163 (N_7163,N_4672,N_4635);
nor U7164 (N_7164,N_5218,N_5033);
xor U7165 (N_7165,N_4487,N_3735);
and U7166 (N_7166,N_4702,N_4095);
nor U7167 (N_7167,N_3500,N_3416);
or U7168 (N_7168,N_6183,N_4980);
or U7169 (N_7169,N_4532,N_3282);
or U7170 (N_7170,N_3505,N_6110);
xnor U7171 (N_7171,N_5559,N_3231);
nand U7172 (N_7172,N_3314,N_6064);
nor U7173 (N_7173,N_3443,N_5200);
nor U7174 (N_7174,N_5653,N_4040);
xor U7175 (N_7175,N_5535,N_4533);
nand U7176 (N_7176,N_5277,N_4329);
nor U7177 (N_7177,N_4676,N_4464);
nor U7178 (N_7178,N_3227,N_5532);
nor U7179 (N_7179,N_5262,N_4912);
nand U7180 (N_7180,N_4862,N_6101);
nand U7181 (N_7181,N_5835,N_4353);
nand U7182 (N_7182,N_3411,N_3395);
and U7183 (N_7183,N_5688,N_5886);
xnor U7184 (N_7184,N_4577,N_4043);
nand U7185 (N_7185,N_5146,N_3195);
and U7186 (N_7186,N_6091,N_4188);
or U7187 (N_7187,N_6184,N_4664);
xnor U7188 (N_7188,N_4807,N_5921);
xor U7189 (N_7189,N_5164,N_3648);
and U7190 (N_7190,N_4448,N_6098);
xor U7191 (N_7191,N_5534,N_4148);
and U7192 (N_7192,N_6122,N_5335);
or U7193 (N_7193,N_4354,N_4519);
nand U7194 (N_7194,N_5388,N_3377);
or U7195 (N_7195,N_3903,N_3620);
or U7196 (N_7196,N_5018,N_3548);
xnor U7197 (N_7197,N_4701,N_5740);
nor U7198 (N_7198,N_5819,N_3698);
or U7199 (N_7199,N_5020,N_5108);
and U7200 (N_7200,N_6157,N_4254);
nor U7201 (N_7201,N_3562,N_5924);
and U7202 (N_7202,N_5043,N_5268);
xor U7203 (N_7203,N_3233,N_4159);
xnor U7204 (N_7204,N_3647,N_5974);
or U7205 (N_7205,N_3689,N_3240);
xnor U7206 (N_7206,N_6003,N_4128);
nand U7207 (N_7207,N_3513,N_4742);
and U7208 (N_7208,N_4575,N_4153);
or U7209 (N_7209,N_5615,N_4526);
and U7210 (N_7210,N_3489,N_6070);
or U7211 (N_7211,N_4475,N_3582);
or U7212 (N_7212,N_6192,N_4340);
nand U7213 (N_7213,N_3519,N_4468);
nor U7214 (N_7214,N_3238,N_4739);
nor U7215 (N_7215,N_3968,N_3440);
nand U7216 (N_7216,N_6161,N_3638);
and U7217 (N_7217,N_5564,N_4567);
nand U7218 (N_7218,N_3603,N_4344);
and U7219 (N_7219,N_3189,N_4366);
nand U7220 (N_7220,N_5470,N_3666);
or U7221 (N_7221,N_3148,N_5416);
xnor U7222 (N_7222,N_5004,N_4298);
or U7223 (N_7223,N_4065,N_5627);
nand U7224 (N_7224,N_5455,N_3444);
nand U7225 (N_7225,N_5623,N_5133);
nor U7226 (N_7226,N_3350,N_5560);
nor U7227 (N_7227,N_5226,N_4296);
and U7228 (N_7228,N_3363,N_5449);
xnor U7229 (N_7229,N_4132,N_4651);
xnor U7230 (N_7230,N_5365,N_3565);
xnor U7231 (N_7231,N_4754,N_5330);
xor U7232 (N_7232,N_4175,N_4057);
and U7233 (N_7233,N_6131,N_5520);
and U7234 (N_7234,N_5188,N_5693);
nor U7235 (N_7235,N_4247,N_5550);
nand U7236 (N_7236,N_5877,N_3928);
xnor U7237 (N_7237,N_5857,N_4849);
xnor U7238 (N_7238,N_5010,N_4062);
nor U7239 (N_7239,N_5718,N_3871);
nand U7240 (N_7240,N_5824,N_5787);
nand U7241 (N_7241,N_4544,N_5154);
xor U7242 (N_7242,N_3258,N_3595);
xor U7243 (N_7243,N_3969,N_4904);
nand U7244 (N_7244,N_4597,N_5144);
or U7245 (N_7245,N_5080,N_5852);
nor U7246 (N_7246,N_3247,N_4086);
and U7247 (N_7247,N_5089,N_4852);
xor U7248 (N_7248,N_5157,N_5498);
nor U7249 (N_7249,N_6082,N_4941);
and U7250 (N_7250,N_5937,N_4076);
or U7251 (N_7251,N_3153,N_3806);
or U7252 (N_7252,N_3370,N_5287);
xor U7253 (N_7253,N_4753,N_5811);
or U7254 (N_7254,N_5779,N_4555);
or U7255 (N_7255,N_6087,N_5100);
or U7256 (N_7256,N_4956,N_5320);
xor U7257 (N_7257,N_3193,N_6231);
xor U7258 (N_7258,N_4484,N_4283);
xor U7259 (N_7259,N_5616,N_6006);
nand U7260 (N_7260,N_5951,N_5363);
nor U7261 (N_7261,N_6209,N_4032);
and U7262 (N_7262,N_5192,N_3938);
nor U7263 (N_7263,N_4266,N_3902);
xnor U7264 (N_7264,N_3477,N_3615);
nand U7265 (N_7265,N_3899,N_3987);
nor U7266 (N_7266,N_5224,N_4243);
and U7267 (N_7267,N_6088,N_5682);
nor U7268 (N_7268,N_3693,N_4113);
and U7269 (N_7269,N_4463,N_4130);
nor U7270 (N_7270,N_6056,N_4935);
nand U7271 (N_7271,N_5219,N_5222);
xor U7272 (N_7272,N_3755,N_4903);
or U7273 (N_7273,N_3656,N_4030);
and U7274 (N_7274,N_3275,N_4388);
nor U7275 (N_7275,N_6046,N_5816);
nand U7276 (N_7276,N_5716,N_3199);
xnor U7277 (N_7277,N_4529,N_4557);
xnor U7278 (N_7278,N_5786,N_4061);
and U7279 (N_7279,N_5902,N_3904);
nand U7280 (N_7280,N_3828,N_3429);
and U7281 (N_7281,N_6228,N_5214);
nor U7282 (N_7282,N_5278,N_3150);
nor U7283 (N_7283,N_4967,N_5678);
or U7284 (N_7284,N_4565,N_4041);
xnor U7285 (N_7285,N_4824,N_3202);
nor U7286 (N_7286,N_5654,N_5778);
nor U7287 (N_7287,N_5050,N_4815);
nand U7288 (N_7288,N_4850,N_3566);
or U7289 (N_7289,N_3455,N_5000);
and U7290 (N_7290,N_5511,N_3381);
nor U7291 (N_7291,N_5047,N_5610);
nor U7292 (N_7292,N_6159,N_3641);
xor U7293 (N_7293,N_6001,N_4881);
and U7294 (N_7294,N_5555,N_3633);
and U7295 (N_7295,N_5624,N_5468);
nor U7296 (N_7296,N_5976,N_4181);
nor U7297 (N_7297,N_4891,N_4323);
xor U7298 (N_7298,N_5744,N_3589);
nand U7299 (N_7299,N_3433,N_6014);
and U7300 (N_7300,N_4186,N_5732);
or U7301 (N_7301,N_3880,N_4632);
or U7302 (N_7302,N_5280,N_5913);
xor U7303 (N_7303,N_5049,N_4848);
xor U7304 (N_7304,N_3560,N_4275);
nand U7305 (N_7305,N_5492,N_6142);
nor U7306 (N_7306,N_4182,N_5438);
nor U7307 (N_7307,N_3998,N_3551);
and U7308 (N_7308,N_3218,N_5247);
and U7309 (N_7309,N_6104,N_5872);
nor U7310 (N_7310,N_3361,N_4237);
nand U7311 (N_7311,N_5114,N_4400);
or U7312 (N_7312,N_5938,N_3330);
nand U7313 (N_7313,N_4762,N_5499);
nand U7314 (N_7314,N_6187,N_4257);
nor U7315 (N_7315,N_4493,N_4939);
and U7316 (N_7316,N_5283,N_5328);
nor U7317 (N_7317,N_3471,N_4613);
and U7318 (N_7318,N_4221,N_5109);
or U7319 (N_7319,N_5860,N_5622);
xnor U7320 (N_7320,N_4326,N_5463);
nor U7321 (N_7321,N_4913,N_5858);
nor U7322 (N_7322,N_5841,N_3168);
nor U7323 (N_7323,N_3914,N_4964);
nand U7324 (N_7324,N_4996,N_3665);
xor U7325 (N_7325,N_3404,N_5194);
or U7326 (N_7326,N_4055,N_4479);
or U7327 (N_7327,N_3352,N_5321);
nand U7328 (N_7328,N_3910,N_4364);
or U7329 (N_7329,N_5121,N_3838);
nor U7330 (N_7330,N_3394,N_4649);
and U7331 (N_7331,N_4502,N_6016);
nand U7332 (N_7332,N_5143,N_4666);
and U7333 (N_7333,N_6203,N_3558);
xor U7334 (N_7334,N_3599,N_6202);
nand U7335 (N_7335,N_4957,N_3419);
nor U7336 (N_7336,N_3768,N_3716);
nor U7337 (N_7337,N_4160,N_4225);
and U7338 (N_7338,N_4887,N_5338);
or U7339 (N_7339,N_4434,N_3813);
and U7340 (N_7340,N_4476,N_4198);
xor U7341 (N_7341,N_5572,N_5950);
or U7342 (N_7342,N_6095,N_3298);
xnor U7343 (N_7343,N_4238,N_4636);
xnor U7344 (N_7344,N_4105,N_5766);
nand U7345 (N_7345,N_3386,N_3536);
nand U7346 (N_7346,N_3415,N_5148);
nor U7347 (N_7347,N_3274,N_4358);
nor U7348 (N_7348,N_4625,N_5288);
and U7349 (N_7349,N_4012,N_6237);
xnor U7350 (N_7350,N_3264,N_4929);
xnor U7351 (N_7351,N_4478,N_3770);
nor U7352 (N_7352,N_5376,N_5412);
nor U7353 (N_7353,N_4315,N_5987);
nand U7354 (N_7354,N_3345,N_4711);
xnor U7355 (N_7355,N_3414,N_4435);
xor U7356 (N_7356,N_5972,N_5799);
nor U7357 (N_7357,N_5482,N_3819);
nand U7358 (N_7358,N_5078,N_4244);
or U7359 (N_7359,N_4671,N_4717);
xnor U7360 (N_7360,N_4920,N_4331);
nand U7361 (N_7361,N_3759,N_4552);
nand U7362 (N_7362,N_5493,N_5426);
nor U7363 (N_7363,N_5948,N_4585);
or U7364 (N_7364,N_5127,N_5001);
nand U7365 (N_7365,N_3818,N_4054);
or U7366 (N_7366,N_5863,N_3733);
nor U7367 (N_7367,N_3257,N_4940);
or U7368 (N_7368,N_5625,N_4779);
nor U7369 (N_7369,N_5072,N_4845);
or U7370 (N_7370,N_4212,N_6054);
and U7371 (N_7371,N_3709,N_3437);
nor U7372 (N_7372,N_3876,N_3435);
nand U7373 (N_7373,N_4834,N_6200);
and U7374 (N_7374,N_5398,N_4078);
or U7375 (N_7375,N_5642,N_4319);
nor U7376 (N_7376,N_3169,N_5111);
xor U7377 (N_7377,N_5313,N_6211);
nand U7378 (N_7378,N_3210,N_3747);
xnor U7379 (N_7379,N_5752,N_6149);
or U7380 (N_7380,N_4811,N_3319);
nor U7381 (N_7381,N_4363,N_5264);
xnor U7382 (N_7382,N_6030,N_4707);
xor U7383 (N_7383,N_4712,N_4131);
nor U7384 (N_7384,N_4074,N_3196);
or U7385 (N_7385,N_5391,N_5769);
xor U7386 (N_7386,N_3760,N_4124);
and U7387 (N_7387,N_4197,N_3630);
nand U7388 (N_7388,N_4248,N_4638);
xnor U7389 (N_7389,N_4215,N_3617);
nand U7390 (N_7390,N_6201,N_5256);
and U7391 (N_7391,N_4490,N_3736);
nor U7392 (N_7392,N_4942,N_3321);
and U7393 (N_7393,N_4746,N_3827);
xnor U7394 (N_7394,N_3865,N_3901);
and U7395 (N_7395,N_4541,N_5589);
and U7396 (N_7396,N_5044,N_4279);
nor U7397 (N_7397,N_4615,N_4457);
and U7398 (N_7398,N_3743,N_3203);
nand U7399 (N_7399,N_4508,N_4629);
xnor U7400 (N_7400,N_3335,N_4107);
or U7401 (N_7401,N_5843,N_5199);
xor U7402 (N_7402,N_4732,N_3417);
nand U7403 (N_7403,N_5250,N_5425);
xnor U7404 (N_7404,N_5137,N_4581);
or U7405 (N_7405,N_5608,N_3295);
nor U7406 (N_7406,N_4437,N_5800);
nor U7407 (N_7407,N_4634,N_3266);
nor U7408 (N_7408,N_6068,N_3909);
nor U7409 (N_7409,N_4979,N_3717);
or U7410 (N_7410,N_3597,N_3891);
nand U7411 (N_7411,N_5427,N_4970);
xnor U7412 (N_7412,N_4655,N_3311);
xnor U7413 (N_7413,N_5384,N_3915);
nand U7414 (N_7414,N_4918,N_5207);
nand U7415 (N_7415,N_4134,N_5965);
xnor U7416 (N_7416,N_5414,N_5989);
and U7417 (N_7417,N_5181,N_5980);
nand U7418 (N_7418,N_3680,N_6100);
xnor U7419 (N_7419,N_3843,N_4491);
nand U7420 (N_7420,N_6219,N_4360);
or U7421 (N_7421,N_3234,N_5773);
or U7422 (N_7422,N_3981,N_4376);
nor U7423 (N_7423,N_3979,N_3170);
or U7424 (N_7424,N_3992,N_4892);
or U7425 (N_7425,N_4097,N_4675);
nand U7426 (N_7426,N_4637,N_3840);
nor U7427 (N_7427,N_3407,N_4079);
and U7428 (N_7428,N_3829,N_6008);
and U7429 (N_7429,N_3468,N_6020);
nand U7430 (N_7430,N_3676,N_3946);
nor U7431 (N_7431,N_5234,N_5613);
or U7432 (N_7432,N_3687,N_5728);
xor U7433 (N_7433,N_3913,N_4542);
nor U7434 (N_7434,N_3391,N_3609);
and U7435 (N_7435,N_6246,N_5349);
and U7436 (N_7436,N_5418,N_3664);
nor U7437 (N_7437,N_3696,N_4436);
xnor U7438 (N_7438,N_5993,N_5417);
nand U7439 (N_7439,N_5377,N_5097);
or U7440 (N_7440,N_4318,N_3889);
xor U7441 (N_7441,N_4975,N_6017);
and U7442 (N_7442,N_3669,N_4559);
and U7443 (N_7443,N_4931,N_5063);
or U7444 (N_7444,N_5190,N_6077);
and U7445 (N_7445,N_4514,N_6208);
nand U7446 (N_7446,N_5290,N_4607);
nand U7447 (N_7447,N_4851,N_5570);
nor U7448 (N_7448,N_6010,N_3594);
or U7449 (N_7449,N_5502,N_4332);
nand U7450 (N_7450,N_3542,N_3457);
nor U7451 (N_7451,N_4728,N_5092);
nor U7452 (N_7452,N_3879,N_6031);
nor U7453 (N_7453,N_4006,N_3734);
nor U7454 (N_7454,N_6154,N_3490);
or U7455 (N_7455,N_5522,N_3781);
or U7456 (N_7456,N_4276,N_4123);
and U7457 (N_7457,N_3186,N_5466);
and U7458 (N_7458,N_5743,N_3166);
and U7459 (N_7459,N_4504,N_4692);
and U7460 (N_7460,N_6099,N_3940);
nor U7461 (N_7461,N_6060,N_4748);
or U7462 (N_7462,N_4652,N_5731);
nor U7463 (N_7463,N_5676,N_3412);
or U7464 (N_7464,N_6113,N_3752);
or U7465 (N_7465,N_5764,N_4206);
xnor U7466 (N_7466,N_4381,N_3636);
xor U7467 (N_7467,N_4772,N_4745);
nor U7468 (N_7468,N_4580,N_6012);
nand U7469 (N_7469,N_3847,N_5865);
or U7470 (N_7470,N_6103,N_5158);
and U7471 (N_7471,N_5284,N_5850);
and U7472 (N_7472,N_3953,N_3347);
nand U7473 (N_7473,N_5672,N_3884);
or U7474 (N_7474,N_4444,N_5512);
xor U7475 (N_7475,N_5061,N_5172);
or U7476 (N_7476,N_4455,N_6092);
nor U7477 (N_7477,N_4568,N_6140);
and U7478 (N_7478,N_4950,N_6105);
nand U7479 (N_7479,N_6225,N_3272);
nand U7480 (N_7480,N_6162,N_3645);
nand U7481 (N_7481,N_4199,N_4500);
or U7482 (N_7482,N_4880,N_3750);
and U7483 (N_7483,N_3796,N_5227);
or U7484 (N_7484,N_5223,N_3450);
or U7485 (N_7485,N_4535,N_3906);
nor U7486 (N_7486,N_5170,N_3874);
nor U7487 (N_7487,N_5495,N_4821);
and U7488 (N_7488,N_5963,N_4734);
and U7489 (N_7489,N_4916,N_3823);
nor U7490 (N_7490,N_4910,N_5034);
nor U7491 (N_7491,N_5355,N_4773);
nand U7492 (N_7492,N_3777,N_3877);
and U7493 (N_7493,N_4917,N_5307);
or U7494 (N_7494,N_6126,N_5713);
or U7495 (N_7495,N_6186,N_6015);
nor U7496 (N_7496,N_3672,N_4578);
or U7497 (N_7497,N_6171,N_6236);
or U7498 (N_7498,N_4373,N_5911);
and U7499 (N_7499,N_5305,N_5595);
nor U7500 (N_7500,N_4156,N_3762);
nor U7501 (N_7501,N_3837,N_4161);
nor U7502 (N_7502,N_5483,N_5685);
xnor U7503 (N_7503,N_4752,N_5945);
and U7504 (N_7504,N_5895,N_6005);
and U7505 (N_7505,N_4026,N_3478);
nor U7506 (N_7506,N_6155,N_5056);
nand U7507 (N_7507,N_4352,N_5173);
or U7508 (N_7508,N_3640,N_5489);
and U7509 (N_7509,N_3623,N_5552);
or U7510 (N_7510,N_5727,N_3569);
nor U7511 (N_7511,N_4945,N_5635);
nand U7512 (N_7512,N_4617,N_4226);
xor U7513 (N_7513,N_3742,N_5822);
nor U7514 (N_7514,N_5566,N_4841);
and U7515 (N_7515,N_5257,N_5827);
xor U7516 (N_7516,N_5032,N_4727);
or U7517 (N_7517,N_5982,N_5130);
nor U7518 (N_7518,N_3262,N_4646);
and U7519 (N_7519,N_3230,N_4823);
xnor U7520 (N_7520,N_5862,N_3625);
nor U7521 (N_7521,N_5668,N_6039);
nor U7522 (N_7522,N_4981,N_5472);
or U7523 (N_7523,N_4232,N_4554);
or U7524 (N_7524,N_5670,N_3387);
xnor U7525 (N_7525,N_3277,N_3300);
xnor U7526 (N_7526,N_4205,N_5621);
nor U7527 (N_7527,N_3936,N_3495);
nand U7528 (N_7528,N_4674,N_4953);
nand U7529 (N_7529,N_3474,N_3912);
and U7530 (N_7530,N_5139,N_6169);
nand U7531 (N_7531,N_4741,N_4397);
nand U7532 (N_7532,N_3318,N_5159);
nor U7533 (N_7533,N_4486,N_5782);
xnor U7534 (N_7534,N_4461,N_4291);
nor U7535 (N_7535,N_4515,N_3556);
or U7536 (N_7536,N_4630,N_3786);
xnor U7537 (N_7537,N_3538,N_6229);
nand U7538 (N_7538,N_4694,N_5910);
or U7539 (N_7539,N_4740,N_4660);
and U7540 (N_7540,N_5390,N_3857);
nor U7541 (N_7541,N_6072,N_3142);
nor U7542 (N_7542,N_6241,N_4028);
xnor U7543 (N_7543,N_3132,N_4810);
nor U7544 (N_7544,N_4593,N_5781);
nand U7545 (N_7545,N_5151,N_5984);
nand U7546 (N_7546,N_5896,N_3719);
nand U7547 (N_7547,N_6120,N_5074);
and U7548 (N_7548,N_5543,N_4914);
xnor U7549 (N_7549,N_3187,N_5501);
and U7550 (N_7550,N_4411,N_4015);
xor U7551 (N_7551,N_3974,N_4797);
and U7552 (N_7552,N_4976,N_4201);
nand U7553 (N_7553,N_4038,N_3881);
nand U7554 (N_7554,N_6045,N_5956);
or U7555 (N_7555,N_3975,N_3181);
and U7556 (N_7556,N_6013,N_5041);
and U7557 (N_7557,N_4785,N_4033);
xnor U7558 (N_7558,N_4081,N_3614);
xnor U7559 (N_7559,N_4644,N_5705);
and U7560 (N_7560,N_5851,N_4658);
nand U7561 (N_7561,N_5742,N_4780);
and U7562 (N_7562,N_6223,N_3523);
and U7563 (N_7563,N_5597,N_4027);
or U7564 (N_7564,N_5291,N_3483);
or U7565 (N_7565,N_4521,N_6244);
and U7566 (N_7566,N_3675,N_4209);
xnor U7567 (N_7567,N_4427,N_4299);
or U7568 (N_7568,N_3692,N_4770);
nand U7569 (N_7569,N_4691,N_3642);
nand U7570 (N_7570,N_4528,N_4482);
nor U7571 (N_7571,N_5603,N_4066);
nand U7572 (N_7572,N_3584,N_4799);
nor U7573 (N_7573,N_4001,N_5696);
xnor U7574 (N_7574,N_5912,N_5739);
xnor U7575 (N_7575,N_5430,N_3794);
nor U7576 (N_7576,N_4034,N_3601);
nor U7577 (N_7577,N_6141,N_3327);
xnor U7578 (N_7578,N_4546,N_5717);
nor U7579 (N_7579,N_4716,N_3883);
nand U7580 (N_7580,N_3194,N_3708);
xnor U7581 (N_7581,N_4846,N_4420);
and U7582 (N_7582,N_3607,N_4895);
xor U7583 (N_7583,N_3546,N_3867);
or U7584 (N_7584,N_4563,N_3252);
and U7585 (N_7585,N_3401,N_3283);
nor U7586 (N_7586,N_5385,N_5271);
and U7587 (N_7587,N_3297,N_6067);
or U7588 (N_7588,N_3815,N_4125);
nand U7589 (N_7589,N_4866,N_4452);
nand U7590 (N_7590,N_4389,N_5939);
or U7591 (N_7591,N_4587,N_5076);
and U7592 (N_7592,N_3281,N_3253);
or U7593 (N_7593,N_5217,N_3849);
and U7594 (N_7594,N_6065,N_5055);
or U7595 (N_7595,N_5129,N_4789);
or U7596 (N_7596,N_4574,N_3143);
nor U7597 (N_7597,N_5155,N_5708);
xnor U7598 (N_7598,N_6112,N_4495);
or U7599 (N_7599,N_4142,N_3496);
or U7600 (N_7600,N_4620,N_4290);
or U7601 (N_7601,N_3375,N_4422);
or U7602 (N_7602,N_3950,N_3745);
or U7603 (N_7603,N_5591,N_5138);
or U7604 (N_7604,N_5999,N_6153);
nand U7605 (N_7605,N_5763,N_3831);
or U7606 (N_7606,N_4669,N_4143);
nand U7607 (N_7607,N_5473,N_5093);
nand U7608 (N_7608,N_5667,N_4536);
and U7609 (N_7609,N_5342,N_3342);
nor U7610 (N_7610,N_5481,N_3479);
nor U7611 (N_7611,N_3279,N_4582);
and U7612 (N_7612,N_5701,N_4052);
xor U7613 (N_7613,N_4307,N_5927);
or U7614 (N_7614,N_4472,N_6213);
nand U7615 (N_7615,N_3724,N_4167);
and U7616 (N_7616,N_6028,N_5810);
xor U7617 (N_7617,N_4446,N_4394);
xor U7618 (N_7618,N_3271,N_3701);
nand U7619 (N_7619,N_5875,N_6094);
nor U7620 (N_7620,N_6249,N_3135);
nand U7621 (N_7621,N_3868,N_4689);
xnor U7622 (N_7622,N_4700,N_4723);
nor U7623 (N_7623,N_3354,N_3711);
or U7624 (N_7624,N_4714,N_4893);
xor U7625 (N_7625,N_4396,N_4100);
nor U7626 (N_7626,N_5211,N_3832);
xnor U7627 (N_7627,N_4413,N_3299);
and U7628 (N_7628,N_4639,N_4214);
and U7629 (N_7629,N_5243,N_3403);
nor U7630 (N_7630,N_3178,N_3670);
nor U7631 (N_7631,N_3408,N_6166);
and U7632 (N_7632,N_5428,N_3553);
and U7633 (N_7633,N_3176,N_5751);
nand U7634 (N_7634,N_5842,N_3758);
nand U7635 (N_7635,N_5998,N_4324);
or U7636 (N_7636,N_3845,N_3390);
or U7637 (N_7637,N_4763,N_5715);
nor U7638 (N_7638,N_5706,N_3729);
or U7639 (N_7639,N_5990,N_5259);
xor U7640 (N_7640,N_4356,N_5327);
and U7641 (N_7641,N_6128,N_5331);
xnor U7642 (N_7642,N_4335,N_3306);
xor U7643 (N_7643,N_3379,N_5643);
and U7644 (N_7644,N_5600,N_4184);
nor U7645 (N_7645,N_3908,N_3659);
or U7646 (N_7646,N_6144,N_3611);
nor U7647 (N_7647,N_3155,N_3315);
nand U7648 (N_7648,N_4347,N_4839);
nand U7649 (N_7649,N_5052,N_4512);
nor U7650 (N_7650,N_3380,N_5554);
xnor U7651 (N_7651,N_6212,N_3731);
xnor U7652 (N_7652,N_4923,N_4670);
and U7653 (N_7653,N_3461,N_6130);
xor U7654 (N_7654,N_5085,N_3167);
and U7655 (N_7655,N_3126,N_5162);
and U7656 (N_7656,N_4679,N_6189);
nand U7657 (N_7657,N_4539,N_5733);
xor U7658 (N_7658,N_3425,N_4306);
or U7659 (N_7659,N_5777,N_6004);
xnor U7660 (N_7660,N_3222,N_3963);
or U7661 (N_7661,N_4350,N_4053);
nor U7662 (N_7662,N_4930,N_4547);
nor U7663 (N_7663,N_3273,N_5410);
and U7664 (N_7664,N_5640,N_5251);
or U7665 (N_7665,N_5189,N_4192);
and U7666 (N_7666,N_4792,N_6195);
xnor U7667 (N_7667,N_4234,N_3508);
xnor U7668 (N_7668,N_3774,N_6111);
xor U7669 (N_7669,N_4093,N_4271);
or U7670 (N_7670,N_5296,N_3358);
and U7671 (N_7671,N_4303,N_6116);
xor U7672 (N_7672,N_5161,N_3585);
nand U7673 (N_7673,N_3555,N_4272);
and U7674 (N_7674,N_5073,N_4836);
or U7675 (N_7675,N_5598,N_5508);
nor U7676 (N_7676,N_4837,N_3313);
or U7677 (N_7677,N_4108,N_4371);
and U7678 (N_7678,N_3510,N_4907);
and U7679 (N_7679,N_5995,N_5745);
or U7680 (N_7680,N_4278,N_5587);
and U7681 (N_7681,N_4888,N_6245);
and U7682 (N_7682,N_6061,N_5531);
or U7683 (N_7683,N_3922,N_4867);
and U7684 (N_7684,N_3156,N_3799);
nor U7685 (N_7685,N_4050,N_5991);
nand U7686 (N_7686,N_5638,N_5873);
or U7687 (N_7687,N_3980,N_3162);
nor U7688 (N_7688,N_6164,N_3651);
or U7689 (N_7689,N_3970,N_4328);
nor U7690 (N_7690,N_5721,N_3145);
or U7691 (N_7691,N_4311,N_6138);
and U7692 (N_7692,N_5647,N_5988);
or U7693 (N_7693,N_5525,N_3627);
xor U7694 (N_7694,N_3540,N_3475);
or U7695 (N_7695,N_5507,N_3530);
or U7696 (N_7696,N_5360,N_3995);
nand U7697 (N_7697,N_3650,N_6221);
nand U7698 (N_7698,N_4470,N_3893);
nor U7699 (N_7699,N_3348,N_3501);
and U7700 (N_7700,N_5202,N_4840);
xnor U7701 (N_7701,N_5011,N_5941);
nand U7702 (N_7702,N_4224,N_4191);
and U7703 (N_7703,N_4218,N_5662);
and U7704 (N_7704,N_5058,N_3326);
and U7705 (N_7705,N_4204,N_3624);
nor U7706 (N_7706,N_5082,N_3787);
or U7707 (N_7707,N_5968,N_3824);
xnor U7708 (N_7708,N_4042,N_4370);
xnor U7709 (N_7709,N_6247,N_5039);
nor U7710 (N_7710,N_5423,N_6107);
nor U7711 (N_7711,N_3894,N_4025);
and U7712 (N_7712,N_4921,N_3977);
or U7713 (N_7713,N_3409,N_4591);
xnor U7714 (N_7714,N_5496,N_5996);
or U7715 (N_7715,N_4127,N_5691);
nor U7716 (N_7716,N_5297,N_5931);
nand U7717 (N_7717,N_5949,N_5808);
or U7718 (N_7718,N_5592,N_3875);
nand U7719 (N_7719,N_5469,N_4336);
nor U7720 (N_7720,N_6063,N_5210);
xnor U7721 (N_7721,N_3278,N_3592);
nand U7722 (N_7722,N_3284,N_5537);
and U7723 (N_7723,N_5521,N_4661);
and U7724 (N_7724,N_4990,N_4928);
and U7725 (N_7725,N_3732,N_5683);
xnor U7726 (N_7726,N_3612,N_3653);
nor U7727 (N_7727,N_3191,N_5488);
xor U7728 (N_7728,N_5147,N_5737);
nand U7729 (N_7729,N_4626,N_3576);
or U7730 (N_7730,N_4960,N_5971);
xor U7731 (N_7731,N_3292,N_4459);
xor U7732 (N_7732,N_5431,N_3399);
and U7733 (N_7733,N_5606,N_3337);
nor U7734 (N_7734,N_4102,N_4584);
nor U7735 (N_7735,N_6029,N_4103);
xor U7736 (N_7736,N_3480,N_5487);
nand U7737 (N_7737,N_4697,N_4997);
and U7738 (N_7738,N_5681,N_5460);
or U7739 (N_7739,N_3133,N_3588);
and U7740 (N_7740,N_4828,N_5300);
nor U7741 (N_7741,N_5513,N_3801);
and U7742 (N_7742,N_4530,N_4755);
or U7743 (N_7743,N_5026,N_4003);
xor U7744 (N_7744,N_4663,N_4623);
and U7745 (N_7745,N_6132,N_4374);
or U7746 (N_7746,N_4758,N_4441);
or U7747 (N_7747,N_5674,N_3964);
and U7748 (N_7748,N_6071,N_3239);
or U7749 (N_7749,N_5145,N_3792);
xnor U7750 (N_7750,N_5343,N_5023);
nand U7751 (N_7751,N_4896,N_5754);
nor U7752 (N_7752,N_4245,N_3606);
nand U7753 (N_7753,N_3918,N_5422);
nand U7754 (N_7754,N_3952,N_3839);
nand U7755 (N_7755,N_4009,N_4456);
or U7756 (N_7756,N_5067,N_3862);
or U7757 (N_7757,N_4999,N_3367);
or U7758 (N_7758,N_5275,N_3685);
or U7759 (N_7759,N_5141,N_5238);
nand U7760 (N_7760,N_6143,N_4897);
nand U7761 (N_7761,N_3469,N_5393);
and U7762 (N_7762,N_5758,N_5040);
nor U7763 (N_7763,N_4179,N_3503);
nand U7764 (N_7764,N_4709,N_4227);
nor U7765 (N_7765,N_4511,N_4014);
or U7766 (N_7766,N_4802,N_3583);
nand U7767 (N_7767,N_4633,N_5178);
nor U7768 (N_7768,N_3219,N_5444);
and U7769 (N_7769,N_5736,N_3206);
and U7770 (N_7770,N_3705,N_4017);
xnor U7771 (N_7771,N_3484,N_4049);
or U7772 (N_7772,N_4854,N_3241);
nand U7773 (N_7773,N_5122,N_4391);
xor U7774 (N_7774,N_5832,N_5364);
nand U7775 (N_7775,N_5031,N_3389);
and U7776 (N_7776,N_5796,N_4765);
or U7777 (N_7777,N_4122,N_4216);
nor U7778 (N_7778,N_4645,N_5637);
or U7779 (N_7779,N_4406,N_3220);
nor U7780 (N_7780,N_5807,N_4210);
or U7781 (N_7781,N_3872,N_3494);
nand U7782 (N_7782,N_3439,N_5333);
and U7783 (N_7783,N_6129,N_5013);
or U7784 (N_7784,N_4090,N_3660);
or U7785 (N_7785,N_5411,N_6026);
nor U7786 (N_7786,N_6160,N_4068);
and U7787 (N_7787,N_5103,N_5820);
nor U7788 (N_7788,N_5523,N_5936);
or U7789 (N_7789,N_5575,N_4766);
or U7790 (N_7790,N_3235,N_3775);
nor U7791 (N_7791,N_5545,N_4410);
nand U7792 (N_7792,N_5303,N_4029);
and U7793 (N_7793,N_6080,N_3383);
nor U7794 (N_7794,N_3527,N_5952);
nor U7795 (N_7795,N_4592,N_3924);
nand U7796 (N_7796,N_4853,N_4803);
nand U7797 (N_7797,N_3171,N_3207);
or U7798 (N_7798,N_4140,N_4656);
nor U7799 (N_7799,N_5153,N_3442);
xor U7800 (N_7800,N_6139,N_5700);
nand U7801 (N_7801,N_5797,N_3858);
nor U7802 (N_7802,N_4776,N_3129);
or U7803 (N_7803,N_4112,N_5413);
xnor U7804 (N_7804,N_4044,N_4442);
or U7805 (N_7805,N_5517,N_4677);
nor U7806 (N_7806,N_4377,N_4094);
nor U7807 (N_7807,N_4121,N_4010);
xnor U7808 (N_7808,N_5834,N_6049);
and U7809 (N_7809,N_5767,N_3825);
xnor U7810 (N_7810,N_4835,N_4421);
xnor U7811 (N_7811,N_3988,N_4217);
nor U7812 (N_7812,N_3198,N_3760);
xor U7813 (N_7813,N_3816,N_4117);
nand U7814 (N_7814,N_3949,N_4425);
nor U7815 (N_7815,N_3355,N_5302);
xor U7816 (N_7816,N_3169,N_3507);
or U7817 (N_7817,N_5875,N_3467);
or U7818 (N_7818,N_4406,N_5088);
xnor U7819 (N_7819,N_4128,N_6186);
and U7820 (N_7820,N_3809,N_3436);
nor U7821 (N_7821,N_5714,N_4872);
and U7822 (N_7822,N_5707,N_3636);
or U7823 (N_7823,N_4966,N_3417);
or U7824 (N_7824,N_3818,N_3676);
or U7825 (N_7825,N_5285,N_5008);
nand U7826 (N_7826,N_3484,N_5917);
nor U7827 (N_7827,N_3412,N_5773);
nor U7828 (N_7828,N_5993,N_6125);
xor U7829 (N_7829,N_3398,N_4302);
xnor U7830 (N_7830,N_5448,N_3917);
xnor U7831 (N_7831,N_5688,N_6147);
or U7832 (N_7832,N_3225,N_4140);
nand U7833 (N_7833,N_5666,N_4133);
nand U7834 (N_7834,N_5912,N_4995);
xnor U7835 (N_7835,N_4970,N_5619);
nand U7836 (N_7836,N_5743,N_3474);
or U7837 (N_7837,N_6142,N_3301);
and U7838 (N_7838,N_3826,N_5446);
nand U7839 (N_7839,N_4822,N_3343);
xor U7840 (N_7840,N_5818,N_4074);
nor U7841 (N_7841,N_5646,N_4512);
and U7842 (N_7842,N_5428,N_5290);
and U7843 (N_7843,N_4858,N_3722);
nand U7844 (N_7844,N_4431,N_5975);
nor U7845 (N_7845,N_5521,N_4209);
or U7846 (N_7846,N_5649,N_5578);
or U7847 (N_7847,N_4588,N_5204);
nand U7848 (N_7848,N_5104,N_5106);
or U7849 (N_7849,N_4915,N_4236);
nand U7850 (N_7850,N_4354,N_3176);
xor U7851 (N_7851,N_3733,N_4987);
nand U7852 (N_7852,N_4568,N_3605);
and U7853 (N_7853,N_5442,N_5356);
xnor U7854 (N_7854,N_5494,N_5121);
nand U7855 (N_7855,N_5735,N_5315);
and U7856 (N_7856,N_5480,N_3658);
and U7857 (N_7857,N_5547,N_5014);
nor U7858 (N_7858,N_4933,N_3827);
or U7859 (N_7859,N_3837,N_5285);
nand U7860 (N_7860,N_3871,N_5824);
xor U7861 (N_7861,N_5798,N_3676);
or U7862 (N_7862,N_5048,N_5829);
and U7863 (N_7863,N_6001,N_3694);
and U7864 (N_7864,N_3558,N_4796);
xor U7865 (N_7865,N_5382,N_5941);
nor U7866 (N_7866,N_5864,N_5059);
and U7867 (N_7867,N_3294,N_4422);
or U7868 (N_7868,N_5841,N_6216);
xor U7869 (N_7869,N_5892,N_5063);
xor U7870 (N_7870,N_3378,N_6106);
nand U7871 (N_7871,N_5365,N_3787);
xnor U7872 (N_7872,N_3334,N_5516);
xor U7873 (N_7873,N_4635,N_3638);
or U7874 (N_7874,N_3654,N_5981);
nand U7875 (N_7875,N_6054,N_5682);
xor U7876 (N_7876,N_4435,N_6035);
nand U7877 (N_7877,N_6224,N_4741);
nand U7878 (N_7878,N_4504,N_4695);
nor U7879 (N_7879,N_5129,N_5363);
xor U7880 (N_7880,N_6074,N_3943);
xnor U7881 (N_7881,N_4583,N_3620);
nand U7882 (N_7882,N_5834,N_5801);
and U7883 (N_7883,N_6054,N_4298);
nand U7884 (N_7884,N_5882,N_4043);
or U7885 (N_7885,N_3623,N_3771);
xor U7886 (N_7886,N_6073,N_6032);
nand U7887 (N_7887,N_4206,N_5219);
xor U7888 (N_7888,N_5049,N_6136);
nor U7889 (N_7889,N_6093,N_4016);
nand U7890 (N_7890,N_3161,N_6194);
xor U7891 (N_7891,N_4048,N_5610);
xnor U7892 (N_7892,N_3410,N_4166);
nand U7893 (N_7893,N_4934,N_4957);
xnor U7894 (N_7894,N_3895,N_5500);
and U7895 (N_7895,N_5219,N_4583);
and U7896 (N_7896,N_4943,N_5026);
xnor U7897 (N_7897,N_3759,N_3264);
nor U7898 (N_7898,N_5660,N_6046);
nor U7899 (N_7899,N_3358,N_5624);
nor U7900 (N_7900,N_6182,N_4741);
xor U7901 (N_7901,N_5777,N_5146);
or U7902 (N_7902,N_5845,N_6243);
nor U7903 (N_7903,N_4291,N_4568);
or U7904 (N_7904,N_5577,N_3753);
or U7905 (N_7905,N_3160,N_4495);
nor U7906 (N_7906,N_3960,N_3151);
xnor U7907 (N_7907,N_4357,N_5025);
and U7908 (N_7908,N_4159,N_4742);
or U7909 (N_7909,N_3327,N_4909);
and U7910 (N_7910,N_5254,N_3394);
or U7911 (N_7911,N_3343,N_5073);
or U7912 (N_7912,N_5035,N_4617);
xor U7913 (N_7913,N_5760,N_3367);
and U7914 (N_7914,N_5676,N_6076);
nand U7915 (N_7915,N_3930,N_4137);
nor U7916 (N_7916,N_3217,N_3574);
or U7917 (N_7917,N_4352,N_5880);
nand U7918 (N_7918,N_4694,N_4398);
nor U7919 (N_7919,N_3744,N_3914);
and U7920 (N_7920,N_4194,N_4227);
xor U7921 (N_7921,N_3823,N_5260);
xnor U7922 (N_7922,N_5113,N_3419);
nand U7923 (N_7923,N_3830,N_4367);
xnor U7924 (N_7924,N_5488,N_3632);
nand U7925 (N_7925,N_4852,N_4596);
or U7926 (N_7926,N_3631,N_3826);
nand U7927 (N_7927,N_5283,N_3971);
or U7928 (N_7928,N_3486,N_3758);
nand U7929 (N_7929,N_6111,N_3895);
or U7930 (N_7930,N_3363,N_3636);
xor U7931 (N_7931,N_4021,N_3277);
and U7932 (N_7932,N_3682,N_3613);
and U7933 (N_7933,N_3777,N_5683);
or U7934 (N_7934,N_5121,N_5390);
or U7935 (N_7935,N_5814,N_4020);
xor U7936 (N_7936,N_4600,N_3623);
and U7937 (N_7937,N_3649,N_5915);
nand U7938 (N_7938,N_5666,N_5029);
xnor U7939 (N_7939,N_3316,N_3383);
and U7940 (N_7940,N_3806,N_5244);
or U7941 (N_7941,N_4628,N_6063);
and U7942 (N_7942,N_4473,N_4638);
or U7943 (N_7943,N_5983,N_4471);
and U7944 (N_7944,N_5111,N_4419);
xnor U7945 (N_7945,N_5348,N_4150);
and U7946 (N_7946,N_6061,N_5955);
or U7947 (N_7947,N_4639,N_5869);
nand U7948 (N_7948,N_3448,N_3730);
and U7949 (N_7949,N_3136,N_4984);
nor U7950 (N_7950,N_5545,N_5964);
xnor U7951 (N_7951,N_4835,N_5811);
xor U7952 (N_7952,N_5728,N_5618);
nor U7953 (N_7953,N_4046,N_4206);
or U7954 (N_7954,N_4746,N_3808);
xor U7955 (N_7955,N_5608,N_5755);
nor U7956 (N_7956,N_3371,N_5665);
nor U7957 (N_7957,N_5511,N_5060);
and U7958 (N_7958,N_3399,N_4880);
nor U7959 (N_7959,N_5384,N_5617);
and U7960 (N_7960,N_4245,N_3995);
nor U7961 (N_7961,N_5555,N_4861);
nor U7962 (N_7962,N_4577,N_3195);
nand U7963 (N_7963,N_5677,N_4257);
or U7964 (N_7964,N_3982,N_4275);
nand U7965 (N_7965,N_3816,N_4417);
nand U7966 (N_7966,N_3513,N_4391);
nand U7967 (N_7967,N_5561,N_5061);
nor U7968 (N_7968,N_4245,N_5606);
nand U7969 (N_7969,N_4924,N_4339);
nand U7970 (N_7970,N_3196,N_3615);
nor U7971 (N_7971,N_4101,N_5656);
xnor U7972 (N_7972,N_5821,N_5472);
nand U7973 (N_7973,N_5491,N_4205);
nand U7974 (N_7974,N_3331,N_4947);
or U7975 (N_7975,N_4661,N_5482);
or U7976 (N_7976,N_4237,N_5944);
or U7977 (N_7977,N_4979,N_4150);
nand U7978 (N_7978,N_5791,N_5407);
nand U7979 (N_7979,N_4890,N_3503);
xnor U7980 (N_7980,N_4039,N_4547);
and U7981 (N_7981,N_4434,N_4336);
nand U7982 (N_7982,N_4368,N_3583);
xnor U7983 (N_7983,N_5275,N_5539);
or U7984 (N_7984,N_5096,N_6019);
and U7985 (N_7985,N_4308,N_4893);
nor U7986 (N_7986,N_3398,N_4228);
or U7987 (N_7987,N_6067,N_5905);
or U7988 (N_7988,N_4066,N_5151);
nor U7989 (N_7989,N_4086,N_5766);
or U7990 (N_7990,N_4388,N_4259);
nand U7991 (N_7991,N_5400,N_3921);
xor U7992 (N_7992,N_5935,N_5595);
nor U7993 (N_7993,N_5488,N_5839);
xor U7994 (N_7994,N_3574,N_3478);
and U7995 (N_7995,N_5213,N_3948);
xnor U7996 (N_7996,N_5625,N_5939);
xnor U7997 (N_7997,N_6011,N_4182);
or U7998 (N_7998,N_5731,N_4339);
and U7999 (N_7999,N_3862,N_4949);
and U8000 (N_8000,N_5514,N_3163);
nor U8001 (N_8001,N_5699,N_4086);
and U8002 (N_8002,N_4796,N_4470);
nor U8003 (N_8003,N_5181,N_5818);
nor U8004 (N_8004,N_3234,N_4238);
xnor U8005 (N_8005,N_4972,N_4446);
or U8006 (N_8006,N_5315,N_6048);
or U8007 (N_8007,N_5278,N_5122);
xor U8008 (N_8008,N_4180,N_3163);
or U8009 (N_8009,N_3645,N_3689);
and U8010 (N_8010,N_4887,N_3485);
xnor U8011 (N_8011,N_4192,N_3210);
nor U8012 (N_8012,N_3617,N_3559);
xor U8013 (N_8013,N_4532,N_4383);
nor U8014 (N_8014,N_3956,N_4339);
or U8015 (N_8015,N_3192,N_4898);
nor U8016 (N_8016,N_3396,N_3297);
nand U8017 (N_8017,N_3914,N_5871);
or U8018 (N_8018,N_3280,N_5944);
nand U8019 (N_8019,N_4367,N_4430);
and U8020 (N_8020,N_3927,N_4512);
xor U8021 (N_8021,N_5741,N_5201);
nor U8022 (N_8022,N_5280,N_5909);
or U8023 (N_8023,N_3905,N_3353);
nand U8024 (N_8024,N_3651,N_3723);
nor U8025 (N_8025,N_3659,N_3743);
or U8026 (N_8026,N_5141,N_3345);
nor U8027 (N_8027,N_4923,N_3683);
and U8028 (N_8028,N_4891,N_3180);
nand U8029 (N_8029,N_4795,N_3843);
nor U8030 (N_8030,N_5967,N_3978);
nor U8031 (N_8031,N_5808,N_5057);
nor U8032 (N_8032,N_3544,N_4571);
and U8033 (N_8033,N_3459,N_3375);
and U8034 (N_8034,N_5257,N_3518);
or U8035 (N_8035,N_5521,N_5650);
nand U8036 (N_8036,N_4383,N_4174);
and U8037 (N_8037,N_4922,N_3378);
nand U8038 (N_8038,N_5657,N_3602);
nor U8039 (N_8039,N_3660,N_6045);
nor U8040 (N_8040,N_3435,N_5989);
or U8041 (N_8041,N_3968,N_5037);
xnor U8042 (N_8042,N_3882,N_4074);
nor U8043 (N_8043,N_5806,N_4933);
xor U8044 (N_8044,N_3511,N_3598);
or U8045 (N_8045,N_3290,N_4218);
and U8046 (N_8046,N_4257,N_5085);
and U8047 (N_8047,N_5061,N_4843);
nor U8048 (N_8048,N_3413,N_4875);
or U8049 (N_8049,N_3187,N_3758);
or U8050 (N_8050,N_4744,N_4609);
and U8051 (N_8051,N_4545,N_3908);
nand U8052 (N_8052,N_4270,N_5715);
nor U8053 (N_8053,N_5032,N_3246);
or U8054 (N_8054,N_4228,N_4329);
and U8055 (N_8055,N_4504,N_5851);
or U8056 (N_8056,N_5969,N_4066);
nor U8057 (N_8057,N_5415,N_4181);
and U8058 (N_8058,N_3335,N_4553);
nand U8059 (N_8059,N_3446,N_4308);
nor U8060 (N_8060,N_3912,N_4797);
and U8061 (N_8061,N_3193,N_6081);
nor U8062 (N_8062,N_3848,N_5948);
nor U8063 (N_8063,N_6029,N_5213);
xnor U8064 (N_8064,N_5581,N_5172);
nand U8065 (N_8065,N_4330,N_5470);
xnor U8066 (N_8066,N_3566,N_3785);
xnor U8067 (N_8067,N_4441,N_4785);
nand U8068 (N_8068,N_5061,N_4310);
nor U8069 (N_8069,N_4897,N_5635);
and U8070 (N_8070,N_3483,N_5602);
or U8071 (N_8071,N_4188,N_3279);
nor U8072 (N_8072,N_4652,N_5295);
and U8073 (N_8073,N_5103,N_6050);
and U8074 (N_8074,N_6189,N_5390);
and U8075 (N_8075,N_4136,N_3159);
nand U8076 (N_8076,N_5365,N_3961);
xor U8077 (N_8077,N_3845,N_3333);
or U8078 (N_8078,N_4694,N_3271);
and U8079 (N_8079,N_4826,N_6017);
nor U8080 (N_8080,N_5934,N_4206);
nand U8081 (N_8081,N_5470,N_4161);
and U8082 (N_8082,N_3695,N_4171);
xor U8083 (N_8083,N_4218,N_5516);
and U8084 (N_8084,N_5587,N_4990);
nor U8085 (N_8085,N_5207,N_5887);
and U8086 (N_8086,N_5012,N_3456);
nand U8087 (N_8087,N_4791,N_5109);
nor U8088 (N_8088,N_4932,N_5488);
or U8089 (N_8089,N_3953,N_5754);
xor U8090 (N_8090,N_5161,N_5081);
xnor U8091 (N_8091,N_3545,N_3153);
nor U8092 (N_8092,N_5707,N_6051);
nand U8093 (N_8093,N_5027,N_5896);
xnor U8094 (N_8094,N_3296,N_3780);
xor U8095 (N_8095,N_3579,N_5311);
xor U8096 (N_8096,N_3770,N_3448);
and U8097 (N_8097,N_3753,N_5622);
nor U8098 (N_8098,N_4713,N_4080);
and U8099 (N_8099,N_6059,N_3610);
nand U8100 (N_8100,N_5713,N_4754);
nor U8101 (N_8101,N_4545,N_5446);
nor U8102 (N_8102,N_3131,N_5415);
and U8103 (N_8103,N_4484,N_6159);
nor U8104 (N_8104,N_4834,N_4282);
or U8105 (N_8105,N_5248,N_5522);
xnor U8106 (N_8106,N_4403,N_4005);
and U8107 (N_8107,N_5440,N_4624);
or U8108 (N_8108,N_3269,N_4992);
nand U8109 (N_8109,N_3954,N_5127);
xnor U8110 (N_8110,N_5829,N_4750);
and U8111 (N_8111,N_4435,N_4956);
nand U8112 (N_8112,N_5689,N_4131);
or U8113 (N_8113,N_4918,N_3306);
nor U8114 (N_8114,N_4666,N_4436);
xor U8115 (N_8115,N_4478,N_4982);
nand U8116 (N_8116,N_4838,N_4065);
nor U8117 (N_8117,N_3279,N_5355);
nand U8118 (N_8118,N_5210,N_5542);
and U8119 (N_8119,N_6030,N_5590);
or U8120 (N_8120,N_5171,N_3720);
or U8121 (N_8121,N_4674,N_5657);
nor U8122 (N_8122,N_5364,N_5100);
or U8123 (N_8123,N_3958,N_3852);
xnor U8124 (N_8124,N_5355,N_5974);
or U8125 (N_8125,N_5888,N_3425);
nor U8126 (N_8126,N_4149,N_6186);
and U8127 (N_8127,N_3386,N_5642);
xor U8128 (N_8128,N_3373,N_5523);
and U8129 (N_8129,N_5257,N_4293);
or U8130 (N_8130,N_3598,N_4990);
xnor U8131 (N_8131,N_3153,N_4223);
nor U8132 (N_8132,N_5356,N_4056);
and U8133 (N_8133,N_3212,N_5903);
nand U8134 (N_8134,N_5120,N_5524);
or U8135 (N_8135,N_5448,N_5351);
and U8136 (N_8136,N_5039,N_4560);
and U8137 (N_8137,N_4257,N_4948);
or U8138 (N_8138,N_4458,N_5891);
or U8139 (N_8139,N_4856,N_3238);
xnor U8140 (N_8140,N_3611,N_3357);
nor U8141 (N_8141,N_5451,N_4208);
or U8142 (N_8142,N_3821,N_6224);
or U8143 (N_8143,N_3540,N_3978);
nand U8144 (N_8144,N_4518,N_3737);
nor U8145 (N_8145,N_5239,N_3687);
xor U8146 (N_8146,N_4136,N_3432);
nand U8147 (N_8147,N_3958,N_6111);
nor U8148 (N_8148,N_4044,N_4770);
and U8149 (N_8149,N_5743,N_3955);
or U8150 (N_8150,N_5911,N_5200);
or U8151 (N_8151,N_5984,N_5082);
nand U8152 (N_8152,N_4272,N_3215);
xor U8153 (N_8153,N_3514,N_3139);
xor U8154 (N_8154,N_5532,N_5199);
nand U8155 (N_8155,N_6041,N_6227);
nand U8156 (N_8156,N_5930,N_6008);
or U8157 (N_8157,N_5842,N_4504);
nor U8158 (N_8158,N_3506,N_4536);
and U8159 (N_8159,N_5573,N_5000);
nand U8160 (N_8160,N_4462,N_5217);
and U8161 (N_8161,N_3248,N_5248);
and U8162 (N_8162,N_3464,N_3914);
nor U8163 (N_8163,N_5941,N_4339);
nand U8164 (N_8164,N_5471,N_5719);
and U8165 (N_8165,N_6135,N_5676);
and U8166 (N_8166,N_5528,N_3973);
nor U8167 (N_8167,N_3538,N_5552);
or U8168 (N_8168,N_4554,N_4833);
and U8169 (N_8169,N_6196,N_3922);
or U8170 (N_8170,N_5762,N_5047);
nand U8171 (N_8171,N_4735,N_5770);
or U8172 (N_8172,N_3141,N_6244);
nor U8173 (N_8173,N_4937,N_3541);
nand U8174 (N_8174,N_3281,N_5234);
or U8175 (N_8175,N_5324,N_5185);
or U8176 (N_8176,N_3322,N_4354);
xor U8177 (N_8177,N_4533,N_5848);
or U8178 (N_8178,N_5677,N_3650);
nor U8179 (N_8179,N_3241,N_6124);
xnor U8180 (N_8180,N_4654,N_3308);
xor U8181 (N_8181,N_6084,N_4392);
or U8182 (N_8182,N_5405,N_5517);
and U8183 (N_8183,N_5396,N_6069);
xnor U8184 (N_8184,N_6120,N_6148);
or U8185 (N_8185,N_4905,N_3504);
or U8186 (N_8186,N_3746,N_4621);
nor U8187 (N_8187,N_5883,N_5846);
or U8188 (N_8188,N_3551,N_4998);
nor U8189 (N_8189,N_5398,N_5891);
and U8190 (N_8190,N_4667,N_5219);
and U8191 (N_8191,N_6038,N_5851);
nor U8192 (N_8192,N_5402,N_4948);
xnor U8193 (N_8193,N_5084,N_5484);
nand U8194 (N_8194,N_4181,N_5502);
or U8195 (N_8195,N_5520,N_3631);
nand U8196 (N_8196,N_5210,N_5832);
and U8197 (N_8197,N_3768,N_4632);
xor U8198 (N_8198,N_6084,N_5181);
nor U8199 (N_8199,N_5301,N_6176);
or U8200 (N_8200,N_4475,N_5568);
xor U8201 (N_8201,N_3471,N_3578);
nand U8202 (N_8202,N_4569,N_5247);
xnor U8203 (N_8203,N_4512,N_4535);
or U8204 (N_8204,N_5693,N_4596);
nor U8205 (N_8205,N_5091,N_6104);
nor U8206 (N_8206,N_5731,N_5059);
and U8207 (N_8207,N_4334,N_3554);
nand U8208 (N_8208,N_3408,N_3670);
and U8209 (N_8209,N_4869,N_5447);
or U8210 (N_8210,N_4167,N_4993);
nand U8211 (N_8211,N_4532,N_5743);
nor U8212 (N_8212,N_6068,N_4824);
nand U8213 (N_8213,N_5931,N_4443);
nand U8214 (N_8214,N_4710,N_5631);
nand U8215 (N_8215,N_3336,N_3319);
and U8216 (N_8216,N_5535,N_3232);
and U8217 (N_8217,N_3651,N_3541);
nor U8218 (N_8218,N_5154,N_3806);
or U8219 (N_8219,N_5910,N_4080);
xor U8220 (N_8220,N_6103,N_4564);
xor U8221 (N_8221,N_6206,N_5946);
and U8222 (N_8222,N_5729,N_4282);
and U8223 (N_8223,N_3840,N_3971);
xnor U8224 (N_8224,N_4248,N_3490);
and U8225 (N_8225,N_3926,N_5020);
and U8226 (N_8226,N_3364,N_5596);
xnor U8227 (N_8227,N_3724,N_3540);
and U8228 (N_8228,N_5634,N_3906);
nand U8229 (N_8229,N_3377,N_5751);
and U8230 (N_8230,N_5449,N_3573);
or U8231 (N_8231,N_4051,N_4300);
and U8232 (N_8232,N_6155,N_3494);
xor U8233 (N_8233,N_4869,N_3877);
or U8234 (N_8234,N_6222,N_5753);
nand U8235 (N_8235,N_5485,N_6184);
xor U8236 (N_8236,N_5225,N_5017);
or U8237 (N_8237,N_5898,N_5897);
nand U8238 (N_8238,N_4661,N_4213);
and U8239 (N_8239,N_3662,N_4330);
and U8240 (N_8240,N_4151,N_5235);
and U8241 (N_8241,N_4944,N_5653);
nor U8242 (N_8242,N_3420,N_5759);
or U8243 (N_8243,N_5090,N_6069);
or U8244 (N_8244,N_3747,N_4182);
nor U8245 (N_8245,N_4414,N_4877);
nor U8246 (N_8246,N_5061,N_6126);
nor U8247 (N_8247,N_5626,N_3445);
and U8248 (N_8248,N_3811,N_6181);
and U8249 (N_8249,N_3250,N_5527);
or U8250 (N_8250,N_4260,N_3908);
nor U8251 (N_8251,N_3371,N_5816);
nor U8252 (N_8252,N_3634,N_5032);
or U8253 (N_8253,N_3953,N_4034);
xor U8254 (N_8254,N_4355,N_5963);
nor U8255 (N_8255,N_6104,N_3486);
xor U8256 (N_8256,N_3787,N_4308);
nand U8257 (N_8257,N_6206,N_5832);
xor U8258 (N_8258,N_6201,N_5695);
nand U8259 (N_8259,N_5821,N_5494);
or U8260 (N_8260,N_6062,N_3784);
nor U8261 (N_8261,N_4406,N_4345);
xor U8262 (N_8262,N_4664,N_3493);
nand U8263 (N_8263,N_4827,N_3211);
or U8264 (N_8264,N_4490,N_3712);
and U8265 (N_8265,N_5060,N_4701);
nor U8266 (N_8266,N_3629,N_5534);
nor U8267 (N_8267,N_3777,N_3137);
nor U8268 (N_8268,N_4790,N_4744);
and U8269 (N_8269,N_3786,N_4509);
nand U8270 (N_8270,N_3783,N_5389);
nand U8271 (N_8271,N_3719,N_4707);
and U8272 (N_8272,N_3438,N_4382);
and U8273 (N_8273,N_3510,N_5214);
xnor U8274 (N_8274,N_4062,N_3834);
nand U8275 (N_8275,N_3937,N_4349);
nand U8276 (N_8276,N_5694,N_3779);
nor U8277 (N_8277,N_6209,N_4945);
xnor U8278 (N_8278,N_5719,N_3410);
and U8279 (N_8279,N_6237,N_4179);
nor U8280 (N_8280,N_5775,N_3755);
or U8281 (N_8281,N_3812,N_5820);
xor U8282 (N_8282,N_3821,N_3928);
or U8283 (N_8283,N_3765,N_3635);
or U8284 (N_8284,N_4617,N_4300);
and U8285 (N_8285,N_4253,N_6097);
nand U8286 (N_8286,N_5453,N_5108);
or U8287 (N_8287,N_3806,N_4989);
nor U8288 (N_8288,N_6178,N_3158);
or U8289 (N_8289,N_4785,N_3786);
nand U8290 (N_8290,N_3413,N_4461);
and U8291 (N_8291,N_5722,N_3235);
nand U8292 (N_8292,N_3895,N_3436);
or U8293 (N_8293,N_4091,N_3195);
nand U8294 (N_8294,N_3544,N_5074);
nor U8295 (N_8295,N_4574,N_4582);
or U8296 (N_8296,N_6044,N_5456);
and U8297 (N_8297,N_4602,N_3926);
xnor U8298 (N_8298,N_3987,N_4475);
and U8299 (N_8299,N_6026,N_6113);
nor U8300 (N_8300,N_4900,N_4917);
and U8301 (N_8301,N_4200,N_5253);
xor U8302 (N_8302,N_6010,N_4810);
xor U8303 (N_8303,N_6146,N_5364);
and U8304 (N_8304,N_3973,N_5065);
xnor U8305 (N_8305,N_3181,N_3456);
nor U8306 (N_8306,N_3644,N_4342);
or U8307 (N_8307,N_5342,N_6005);
and U8308 (N_8308,N_5910,N_4730);
nand U8309 (N_8309,N_5907,N_3583);
xnor U8310 (N_8310,N_3275,N_3371);
xor U8311 (N_8311,N_4741,N_5175);
nand U8312 (N_8312,N_5020,N_3997);
and U8313 (N_8313,N_4753,N_4536);
nor U8314 (N_8314,N_3582,N_5679);
nand U8315 (N_8315,N_3508,N_5546);
nand U8316 (N_8316,N_4902,N_5722);
and U8317 (N_8317,N_3379,N_5917);
and U8318 (N_8318,N_4509,N_5832);
nor U8319 (N_8319,N_4819,N_3178);
nand U8320 (N_8320,N_4429,N_4577);
nand U8321 (N_8321,N_3942,N_5241);
nand U8322 (N_8322,N_3403,N_3248);
nor U8323 (N_8323,N_4040,N_4536);
xnor U8324 (N_8324,N_5758,N_3807);
and U8325 (N_8325,N_5389,N_3309);
nor U8326 (N_8326,N_3159,N_4183);
or U8327 (N_8327,N_4089,N_3401);
xnor U8328 (N_8328,N_3181,N_5108);
xor U8329 (N_8329,N_5917,N_3446);
xnor U8330 (N_8330,N_4434,N_4771);
and U8331 (N_8331,N_3920,N_5861);
nand U8332 (N_8332,N_3316,N_5759);
and U8333 (N_8333,N_3895,N_3373);
and U8334 (N_8334,N_5973,N_3679);
or U8335 (N_8335,N_5155,N_5658);
and U8336 (N_8336,N_4512,N_4996);
nor U8337 (N_8337,N_4126,N_4252);
nand U8338 (N_8338,N_6231,N_4327);
and U8339 (N_8339,N_5473,N_3322);
xor U8340 (N_8340,N_6190,N_4346);
nor U8341 (N_8341,N_5185,N_4328);
xor U8342 (N_8342,N_3979,N_4572);
nor U8343 (N_8343,N_3840,N_5343);
and U8344 (N_8344,N_3605,N_4428);
or U8345 (N_8345,N_3283,N_3880);
and U8346 (N_8346,N_3795,N_3592);
or U8347 (N_8347,N_4174,N_5161);
nand U8348 (N_8348,N_5815,N_3322);
and U8349 (N_8349,N_5619,N_4969);
nand U8350 (N_8350,N_4404,N_3851);
or U8351 (N_8351,N_4246,N_5969);
or U8352 (N_8352,N_5336,N_5746);
nor U8353 (N_8353,N_5925,N_4612);
or U8354 (N_8354,N_5898,N_5421);
nor U8355 (N_8355,N_4969,N_3186);
and U8356 (N_8356,N_3138,N_3520);
xor U8357 (N_8357,N_3876,N_4057);
nor U8358 (N_8358,N_4131,N_4358);
nor U8359 (N_8359,N_4766,N_3667);
xnor U8360 (N_8360,N_4612,N_5868);
xor U8361 (N_8361,N_3682,N_5734);
and U8362 (N_8362,N_4921,N_5610);
nand U8363 (N_8363,N_3976,N_3461);
nor U8364 (N_8364,N_3406,N_6100);
nor U8365 (N_8365,N_5513,N_3443);
nor U8366 (N_8366,N_5123,N_4115);
nor U8367 (N_8367,N_3707,N_6126);
xor U8368 (N_8368,N_3222,N_5523);
nor U8369 (N_8369,N_3462,N_5952);
nand U8370 (N_8370,N_4805,N_4453);
nor U8371 (N_8371,N_3544,N_4994);
xor U8372 (N_8372,N_4088,N_5936);
xor U8373 (N_8373,N_5092,N_3382);
and U8374 (N_8374,N_6165,N_3701);
and U8375 (N_8375,N_4428,N_4062);
xor U8376 (N_8376,N_6081,N_3597);
and U8377 (N_8377,N_4747,N_3271);
and U8378 (N_8378,N_5533,N_4267);
and U8379 (N_8379,N_4853,N_4688);
xor U8380 (N_8380,N_3850,N_3635);
nor U8381 (N_8381,N_5978,N_5362);
or U8382 (N_8382,N_3829,N_5343);
nand U8383 (N_8383,N_6028,N_5152);
nand U8384 (N_8384,N_5719,N_5007);
xor U8385 (N_8385,N_4408,N_3386);
nor U8386 (N_8386,N_5827,N_5717);
and U8387 (N_8387,N_4275,N_5914);
xnor U8388 (N_8388,N_4935,N_4011);
nand U8389 (N_8389,N_6196,N_5325);
or U8390 (N_8390,N_6177,N_5105);
xnor U8391 (N_8391,N_4209,N_3485);
nor U8392 (N_8392,N_3676,N_5193);
and U8393 (N_8393,N_4488,N_6186);
or U8394 (N_8394,N_5798,N_4694);
xnor U8395 (N_8395,N_4460,N_4356);
nand U8396 (N_8396,N_5197,N_6242);
xor U8397 (N_8397,N_5351,N_6039);
or U8398 (N_8398,N_5145,N_4586);
xnor U8399 (N_8399,N_4473,N_4678);
and U8400 (N_8400,N_4230,N_6025);
or U8401 (N_8401,N_5650,N_3215);
or U8402 (N_8402,N_4738,N_5448);
nand U8403 (N_8403,N_6100,N_4756);
nand U8404 (N_8404,N_5499,N_5176);
nand U8405 (N_8405,N_5399,N_3193);
or U8406 (N_8406,N_5672,N_5662);
and U8407 (N_8407,N_4421,N_3910);
xor U8408 (N_8408,N_4362,N_4438);
nor U8409 (N_8409,N_4462,N_6021);
or U8410 (N_8410,N_4107,N_5679);
or U8411 (N_8411,N_3150,N_5520);
or U8412 (N_8412,N_5326,N_5153);
xor U8413 (N_8413,N_5723,N_4618);
nand U8414 (N_8414,N_3498,N_3919);
and U8415 (N_8415,N_5524,N_5707);
xor U8416 (N_8416,N_3732,N_6241);
and U8417 (N_8417,N_4240,N_4696);
xnor U8418 (N_8418,N_5998,N_5280);
and U8419 (N_8419,N_4677,N_4252);
and U8420 (N_8420,N_5656,N_3645);
xnor U8421 (N_8421,N_5072,N_5732);
nor U8422 (N_8422,N_3914,N_4112);
nand U8423 (N_8423,N_5039,N_3883);
and U8424 (N_8424,N_4096,N_4029);
nor U8425 (N_8425,N_4249,N_5166);
nor U8426 (N_8426,N_5659,N_4643);
xor U8427 (N_8427,N_6069,N_3630);
and U8428 (N_8428,N_3645,N_5561);
and U8429 (N_8429,N_5802,N_4887);
nand U8430 (N_8430,N_3827,N_4326);
nand U8431 (N_8431,N_3130,N_3398);
or U8432 (N_8432,N_4928,N_4624);
or U8433 (N_8433,N_5640,N_3494);
xnor U8434 (N_8434,N_3421,N_5634);
and U8435 (N_8435,N_4507,N_5159);
or U8436 (N_8436,N_5021,N_4487);
nand U8437 (N_8437,N_5524,N_3821);
or U8438 (N_8438,N_5343,N_3498);
or U8439 (N_8439,N_6031,N_4555);
nor U8440 (N_8440,N_3741,N_4929);
xnor U8441 (N_8441,N_3487,N_5610);
nor U8442 (N_8442,N_5474,N_3344);
or U8443 (N_8443,N_6005,N_3183);
xor U8444 (N_8444,N_5206,N_4145);
nor U8445 (N_8445,N_3652,N_5520);
nor U8446 (N_8446,N_5540,N_5024);
xor U8447 (N_8447,N_5762,N_4301);
or U8448 (N_8448,N_3471,N_4647);
or U8449 (N_8449,N_3809,N_3942);
nor U8450 (N_8450,N_4738,N_3598);
and U8451 (N_8451,N_4647,N_5014);
nor U8452 (N_8452,N_3627,N_6053);
or U8453 (N_8453,N_6042,N_4596);
nand U8454 (N_8454,N_5843,N_3255);
nand U8455 (N_8455,N_3775,N_5537);
nand U8456 (N_8456,N_4862,N_3541);
nor U8457 (N_8457,N_3996,N_5592);
xnor U8458 (N_8458,N_5163,N_5071);
or U8459 (N_8459,N_4023,N_5052);
or U8460 (N_8460,N_4472,N_4633);
and U8461 (N_8461,N_4645,N_5194);
or U8462 (N_8462,N_3157,N_3994);
or U8463 (N_8463,N_5981,N_6168);
nor U8464 (N_8464,N_5433,N_4607);
nand U8465 (N_8465,N_5022,N_5660);
nand U8466 (N_8466,N_5095,N_6112);
or U8467 (N_8467,N_5498,N_4192);
xor U8468 (N_8468,N_5279,N_5355);
or U8469 (N_8469,N_3514,N_5481);
xnor U8470 (N_8470,N_6173,N_5503);
nand U8471 (N_8471,N_5063,N_3887);
xor U8472 (N_8472,N_5122,N_4790);
or U8473 (N_8473,N_5503,N_4401);
and U8474 (N_8474,N_3391,N_3959);
xnor U8475 (N_8475,N_3759,N_5177);
nor U8476 (N_8476,N_5964,N_3383);
or U8477 (N_8477,N_3140,N_4514);
nand U8478 (N_8478,N_4328,N_3686);
and U8479 (N_8479,N_3938,N_5278);
and U8480 (N_8480,N_5839,N_4131);
and U8481 (N_8481,N_4790,N_3597);
or U8482 (N_8482,N_4532,N_3259);
or U8483 (N_8483,N_6059,N_4926);
nand U8484 (N_8484,N_4017,N_3275);
or U8485 (N_8485,N_4544,N_6013);
or U8486 (N_8486,N_3375,N_3491);
and U8487 (N_8487,N_4817,N_5016);
nand U8488 (N_8488,N_3315,N_6162);
or U8489 (N_8489,N_5464,N_4637);
or U8490 (N_8490,N_5147,N_6122);
nor U8491 (N_8491,N_5525,N_3601);
nor U8492 (N_8492,N_6170,N_5098);
nand U8493 (N_8493,N_5183,N_5371);
xor U8494 (N_8494,N_3513,N_5140);
or U8495 (N_8495,N_3572,N_4280);
nand U8496 (N_8496,N_3460,N_6163);
xnor U8497 (N_8497,N_4436,N_4854);
xnor U8498 (N_8498,N_5732,N_4554);
nand U8499 (N_8499,N_4097,N_3601);
xor U8500 (N_8500,N_5472,N_4756);
nand U8501 (N_8501,N_3294,N_4918);
xnor U8502 (N_8502,N_5233,N_5898);
and U8503 (N_8503,N_3487,N_5577);
or U8504 (N_8504,N_4104,N_4755);
and U8505 (N_8505,N_4145,N_4261);
and U8506 (N_8506,N_5204,N_3821);
nor U8507 (N_8507,N_4966,N_4131);
or U8508 (N_8508,N_5813,N_3286);
or U8509 (N_8509,N_5431,N_4248);
or U8510 (N_8510,N_5534,N_4895);
nor U8511 (N_8511,N_5868,N_4528);
or U8512 (N_8512,N_3332,N_5827);
or U8513 (N_8513,N_5871,N_4747);
and U8514 (N_8514,N_5781,N_3913);
or U8515 (N_8515,N_4676,N_4947);
nor U8516 (N_8516,N_3752,N_6198);
or U8517 (N_8517,N_4423,N_3544);
nor U8518 (N_8518,N_4956,N_3484);
or U8519 (N_8519,N_5918,N_5464);
xor U8520 (N_8520,N_6164,N_5691);
nand U8521 (N_8521,N_5828,N_3355);
or U8522 (N_8522,N_6068,N_5217);
xor U8523 (N_8523,N_5599,N_6132);
or U8524 (N_8524,N_5214,N_6054);
nor U8525 (N_8525,N_3558,N_5122);
and U8526 (N_8526,N_3219,N_4678);
nor U8527 (N_8527,N_5973,N_4780);
nor U8528 (N_8528,N_3156,N_4526);
nand U8529 (N_8529,N_5991,N_3406);
and U8530 (N_8530,N_6170,N_6122);
nand U8531 (N_8531,N_5984,N_6009);
and U8532 (N_8532,N_6199,N_5196);
and U8533 (N_8533,N_6057,N_5890);
or U8534 (N_8534,N_3965,N_4185);
nor U8535 (N_8535,N_6067,N_5743);
or U8536 (N_8536,N_5929,N_3516);
or U8537 (N_8537,N_4787,N_4984);
and U8538 (N_8538,N_3782,N_4784);
or U8539 (N_8539,N_3938,N_5677);
xor U8540 (N_8540,N_4646,N_5748);
or U8541 (N_8541,N_3178,N_4642);
or U8542 (N_8542,N_3334,N_4925);
nor U8543 (N_8543,N_5019,N_5855);
and U8544 (N_8544,N_6043,N_5274);
or U8545 (N_8545,N_3571,N_5670);
and U8546 (N_8546,N_5196,N_4090);
or U8547 (N_8547,N_4690,N_6105);
xnor U8548 (N_8548,N_3157,N_5885);
and U8549 (N_8549,N_4136,N_5106);
nand U8550 (N_8550,N_5091,N_5006);
nor U8551 (N_8551,N_5657,N_6205);
nor U8552 (N_8552,N_5542,N_3729);
xor U8553 (N_8553,N_5814,N_5735);
or U8554 (N_8554,N_5721,N_5294);
nor U8555 (N_8555,N_4601,N_3449);
nand U8556 (N_8556,N_4014,N_5840);
nand U8557 (N_8557,N_5034,N_5627);
or U8558 (N_8558,N_4664,N_3719);
nand U8559 (N_8559,N_5082,N_3324);
nand U8560 (N_8560,N_4316,N_6184);
or U8561 (N_8561,N_5745,N_5302);
or U8562 (N_8562,N_5317,N_3768);
nand U8563 (N_8563,N_5835,N_5159);
nor U8564 (N_8564,N_4275,N_5359);
xor U8565 (N_8565,N_4466,N_4839);
nand U8566 (N_8566,N_3472,N_4383);
nor U8567 (N_8567,N_3172,N_5009);
nand U8568 (N_8568,N_3243,N_5853);
nand U8569 (N_8569,N_3639,N_4113);
nand U8570 (N_8570,N_5085,N_4682);
and U8571 (N_8571,N_3225,N_3298);
xor U8572 (N_8572,N_5223,N_3994);
xor U8573 (N_8573,N_5329,N_4443);
xnor U8574 (N_8574,N_4503,N_3909);
nand U8575 (N_8575,N_4511,N_4069);
or U8576 (N_8576,N_5578,N_4396);
or U8577 (N_8577,N_3325,N_4831);
xnor U8578 (N_8578,N_5212,N_4035);
nand U8579 (N_8579,N_3134,N_5137);
or U8580 (N_8580,N_5520,N_4624);
nor U8581 (N_8581,N_4007,N_3986);
and U8582 (N_8582,N_5324,N_6094);
and U8583 (N_8583,N_3508,N_3669);
xnor U8584 (N_8584,N_3581,N_3909);
nand U8585 (N_8585,N_4114,N_5854);
xor U8586 (N_8586,N_4549,N_3141);
nor U8587 (N_8587,N_3263,N_4678);
nand U8588 (N_8588,N_3680,N_3298);
xor U8589 (N_8589,N_4136,N_4507);
or U8590 (N_8590,N_4073,N_6020);
xnor U8591 (N_8591,N_5759,N_6213);
nor U8592 (N_8592,N_4409,N_6192);
xor U8593 (N_8593,N_4527,N_3822);
and U8594 (N_8594,N_3355,N_4084);
or U8595 (N_8595,N_6138,N_4748);
or U8596 (N_8596,N_3884,N_5559);
nand U8597 (N_8597,N_4618,N_4744);
or U8598 (N_8598,N_5590,N_4202);
nand U8599 (N_8599,N_4466,N_5682);
or U8600 (N_8600,N_5880,N_5726);
nor U8601 (N_8601,N_6017,N_4677);
and U8602 (N_8602,N_4957,N_3584);
or U8603 (N_8603,N_3942,N_3965);
nand U8604 (N_8604,N_4527,N_3171);
and U8605 (N_8605,N_4595,N_3868);
and U8606 (N_8606,N_5324,N_6143);
xnor U8607 (N_8607,N_6116,N_5474);
and U8608 (N_8608,N_6131,N_4268);
and U8609 (N_8609,N_6004,N_5855);
and U8610 (N_8610,N_5029,N_5345);
and U8611 (N_8611,N_5039,N_5086);
nor U8612 (N_8612,N_3771,N_5720);
xnor U8613 (N_8613,N_3738,N_4127);
and U8614 (N_8614,N_4369,N_3569);
nor U8615 (N_8615,N_4631,N_3909);
nor U8616 (N_8616,N_6236,N_3444);
and U8617 (N_8617,N_4704,N_3131);
or U8618 (N_8618,N_5681,N_4563);
or U8619 (N_8619,N_4826,N_5512);
and U8620 (N_8620,N_3441,N_4947);
xor U8621 (N_8621,N_3691,N_5204);
nor U8622 (N_8622,N_3781,N_4731);
xor U8623 (N_8623,N_4143,N_3842);
or U8624 (N_8624,N_3870,N_3362);
and U8625 (N_8625,N_4110,N_5160);
nor U8626 (N_8626,N_4884,N_3355);
nor U8627 (N_8627,N_6085,N_3439);
and U8628 (N_8628,N_3235,N_5314);
or U8629 (N_8629,N_6052,N_3611);
nor U8630 (N_8630,N_4243,N_6100);
xnor U8631 (N_8631,N_3662,N_6214);
and U8632 (N_8632,N_5053,N_4928);
xnor U8633 (N_8633,N_4409,N_3382);
and U8634 (N_8634,N_4308,N_5019);
nor U8635 (N_8635,N_5797,N_3464);
nand U8636 (N_8636,N_4806,N_3460);
or U8637 (N_8637,N_6068,N_5091);
nor U8638 (N_8638,N_5999,N_3487);
nor U8639 (N_8639,N_5834,N_3873);
nor U8640 (N_8640,N_5702,N_5098);
nor U8641 (N_8641,N_4801,N_3858);
nand U8642 (N_8642,N_5791,N_3682);
xor U8643 (N_8643,N_3755,N_3718);
nand U8644 (N_8644,N_4050,N_4844);
xor U8645 (N_8645,N_5299,N_3738);
or U8646 (N_8646,N_3473,N_5772);
nor U8647 (N_8647,N_3645,N_5196);
xnor U8648 (N_8648,N_5205,N_4359);
nand U8649 (N_8649,N_5451,N_3205);
nand U8650 (N_8650,N_4641,N_6056);
nor U8651 (N_8651,N_4490,N_5410);
or U8652 (N_8652,N_4433,N_5869);
nand U8653 (N_8653,N_4545,N_4135);
and U8654 (N_8654,N_3365,N_5625);
or U8655 (N_8655,N_4932,N_5904);
xor U8656 (N_8656,N_3127,N_3866);
nand U8657 (N_8657,N_4377,N_4301);
xnor U8658 (N_8658,N_4292,N_4697);
or U8659 (N_8659,N_6169,N_6170);
nand U8660 (N_8660,N_3999,N_3419);
and U8661 (N_8661,N_5619,N_5103);
xnor U8662 (N_8662,N_4460,N_4863);
xnor U8663 (N_8663,N_5551,N_6020);
nand U8664 (N_8664,N_3755,N_3789);
and U8665 (N_8665,N_5564,N_5668);
nor U8666 (N_8666,N_4134,N_3449);
nand U8667 (N_8667,N_4005,N_4247);
nor U8668 (N_8668,N_3372,N_6122);
and U8669 (N_8669,N_5893,N_5608);
nor U8670 (N_8670,N_5909,N_5532);
or U8671 (N_8671,N_6103,N_6030);
nor U8672 (N_8672,N_5699,N_4311);
or U8673 (N_8673,N_4338,N_3317);
xor U8674 (N_8674,N_4531,N_5644);
or U8675 (N_8675,N_5144,N_5608);
nor U8676 (N_8676,N_6133,N_4855);
nand U8677 (N_8677,N_4125,N_5774);
and U8678 (N_8678,N_4132,N_6071);
xor U8679 (N_8679,N_4541,N_4323);
nor U8680 (N_8680,N_5815,N_4845);
or U8681 (N_8681,N_3591,N_4584);
or U8682 (N_8682,N_3220,N_3515);
nand U8683 (N_8683,N_4541,N_5134);
xor U8684 (N_8684,N_5911,N_5184);
xor U8685 (N_8685,N_3714,N_5158);
xor U8686 (N_8686,N_5065,N_4381);
and U8687 (N_8687,N_5040,N_3652);
or U8688 (N_8688,N_3386,N_5963);
and U8689 (N_8689,N_4516,N_6199);
nand U8690 (N_8690,N_4136,N_3729);
or U8691 (N_8691,N_4542,N_3996);
xor U8692 (N_8692,N_3266,N_5944);
or U8693 (N_8693,N_5908,N_3397);
and U8694 (N_8694,N_3533,N_3356);
xor U8695 (N_8695,N_4347,N_4638);
and U8696 (N_8696,N_5083,N_3867);
xor U8697 (N_8697,N_3458,N_6066);
nand U8698 (N_8698,N_4466,N_4621);
and U8699 (N_8699,N_4648,N_4788);
xor U8700 (N_8700,N_3577,N_3677);
or U8701 (N_8701,N_4403,N_4841);
nor U8702 (N_8702,N_3768,N_4282);
and U8703 (N_8703,N_4588,N_5385);
nor U8704 (N_8704,N_5096,N_4851);
or U8705 (N_8705,N_4397,N_4930);
nor U8706 (N_8706,N_4541,N_5023);
nand U8707 (N_8707,N_5657,N_3360);
or U8708 (N_8708,N_3546,N_3911);
nor U8709 (N_8709,N_4614,N_3930);
nor U8710 (N_8710,N_4192,N_5033);
nand U8711 (N_8711,N_3949,N_5727);
xnor U8712 (N_8712,N_4173,N_4048);
nor U8713 (N_8713,N_4587,N_5197);
xor U8714 (N_8714,N_3726,N_3492);
or U8715 (N_8715,N_5410,N_5890);
nor U8716 (N_8716,N_4757,N_4285);
or U8717 (N_8717,N_3979,N_4582);
and U8718 (N_8718,N_5433,N_6221);
and U8719 (N_8719,N_4172,N_4411);
nand U8720 (N_8720,N_5366,N_3864);
or U8721 (N_8721,N_4129,N_6117);
nor U8722 (N_8722,N_5256,N_4564);
nand U8723 (N_8723,N_3848,N_4665);
or U8724 (N_8724,N_3791,N_5501);
xnor U8725 (N_8725,N_4559,N_4986);
nor U8726 (N_8726,N_4649,N_4425);
xor U8727 (N_8727,N_5794,N_4523);
xnor U8728 (N_8728,N_4580,N_5190);
nand U8729 (N_8729,N_3251,N_5217);
and U8730 (N_8730,N_6024,N_4175);
or U8731 (N_8731,N_5211,N_3702);
nand U8732 (N_8732,N_5167,N_5917);
and U8733 (N_8733,N_5462,N_6188);
and U8734 (N_8734,N_5566,N_4963);
nor U8735 (N_8735,N_5196,N_3141);
and U8736 (N_8736,N_6177,N_3492);
and U8737 (N_8737,N_4693,N_3241);
nand U8738 (N_8738,N_4407,N_4092);
and U8739 (N_8739,N_5594,N_3423);
nand U8740 (N_8740,N_3804,N_3151);
nor U8741 (N_8741,N_3244,N_3549);
or U8742 (N_8742,N_4511,N_4446);
or U8743 (N_8743,N_3582,N_5435);
or U8744 (N_8744,N_4438,N_5589);
or U8745 (N_8745,N_5792,N_3574);
and U8746 (N_8746,N_3314,N_3923);
nor U8747 (N_8747,N_3533,N_3861);
xor U8748 (N_8748,N_6172,N_3530);
and U8749 (N_8749,N_6054,N_4497);
and U8750 (N_8750,N_6133,N_4079);
nand U8751 (N_8751,N_3852,N_5546);
xnor U8752 (N_8752,N_6068,N_3967);
and U8753 (N_8753,N_5186,N_4894);
nand U8754 (N_8754,N_4040,N_3576);
xor U8755 (N_8755,N_4415,N_5159);
nor U8756 (N_8756,N_4102,N_4212);
nor U8757 (N_8757,N_4343,N_5993);
xnor U8758 (N_8758,N_3349,N_5853);
or U8759 (N_8759,N_3996,N_3185);
or U8760 (N_8760,N_3556,N_4586);
and U8761 (N_8761,N_4458,N_4829);
nand U8762 (N_8762,N_5195,N_4420);
and U8763 (N_8763,N_5759,N_5003);
nor U8764 (N_8764,N_4720,N_3895);
nand U8765 (N_8765,N_5646,N_3329);
and U8766 (N_8766,N_3139,N_5714);
xnor U8767 (N_8767,N_5469,N_4681);
and U8768 (N_8768,N_4168,N_3862);
xnor U8769 (N_8769,N_4316,N_3278);
or U8770 (N_8770,N_4617,N_5795);
and U8771 (N_8771,N_3848,N_5772);
nand U8772 (N_8772,N_5417,N_5424);
nor U8773 (N_8773,N_5891,N_4739);
nor U8774 (N_8774,N_3801,N_4010);
nand U8775 (N_8775,N_5337,N_5155);
nand U8776 (N_8776,N_6103,N_4358);
or U8777 (N_8777,N_5040,N_5176);
or U8778 (N_8778,N_4206,N_5088);
nand U8779 (N_8779,N_3716,N_5351);
xnor U8780 (N_8780,N_6186,N_5360);
and U8781 (N_8781,N_4282,N_3370);
or U8782 (N_8782,N_4068,N_5565);
nand U8783 (N_8783,N_3367,N_3757);
nor U8784 (N_8784,N_3935,N_5703);
or U8785 (N_8785,N_5614,N_4190);
nand U8786 (N_8786,N_3620,N_4611);
and U8787 (N_8787,N_3133,N_6193);
nand U8788 (N_8788,N_5023,N_4666);
or U8789 (N_8789,N_5427,N_6248);
nor U8790 (N_8790,N_4103,N_3133);
nand U8791 (N_8791,N_3450,N_4735);
nor U8792 (N_8792,N_5545,N_5314);
or U8793 (N_8793,N_3210,N_4773);
and U8794 (N_8794,N_5382,N_3414);
or U8795 (N_8795,N_6134,N_5032);
xnor U8796 (N_8796,N_5673,N_5819);
nand U8797 (N_8797,N_3165,N_4378);
or U8798 (N_8798,N_5581,N_5074);
or U8799 (N_8799,N_4924,N_4272);
nand U8800 (N_8800,N_5367,N_3545);
or U8801 (N_8801,N_4356,N_4110);
or U8802 (N_8802,N_5833,N_3536);
and U8803 (N_8803,N_5941,N_3764);
xnor U8804 (N_8804,N_5894,N_5853);
or U8805 (N_8805,N_4029,N_5747);
nor U8806 (N_8806,N_5911,N_3591);
nand U8807 (N_8807,N_5904,N_4194);
and U8808 (N_8808,N_5328,N_5082);
or U8809 (N_8809,N_5545,N_3667);
nor U8810 (N_8810,N_4166,N_3508);
nor U8811 (N_8811,N_3435,N_5464);
xnor U8812 (N_8812,N_5810,N_3459);
nor U8813 (N_8813,N_4961,N_3906);
and U8814 (N_8814,N_4492,N_3177);
and U8815 (N_8815,N_3468,N_5311);
nand U8816 (N_8816,N_5514,N_5708);
or U8817 (N_8817,N_4276,N_5068);
and U8818 (N_8818,N_4288,N_4680);
nor U8819 (N_8819,N_4927,N_4651);
nor U8820 (N_8820,N_5978,N_4499);
xor U8821 (N_8821,N_4377,N_4484);
xnor U8822 (N_8822,N_5205,N_6035);
and U8823 (N_8823,N_5390,N_5042);
xor U8824 (N_8824,N_3398,N_4547);
nand U8825 (N_8825,N_6221,N_4761);
and U8826 (N_8826,N_3803,N_5643);
xor U8827 (N_8827,N_5435,N_4604);
nand U8828 (N_8828,N_3365,N_5759);
or U8829 (N_8829,N_3931,N_4471);
nor U8830 (N_8830,N_4666,N_3775);
or U8831 (N_8831,N_5220,N_4861);
or U8832 (N_8832,N_4466,N_3885);
and U8833 (N_8833,N_5288,N_5166);
nor U8834 (N_8834,N_4147,N_3657);
or U8835 (N_8835,N_3760,N_4555);
or U8836 (N_8836,N_4484,N_5416);
xor U8837 (N_8837,N_3642,N_4958);
and U8838 (N_8838,N_6022,N_6058);
nor U8839 (N_8839,N_4829,N_5557);
nand U8840 (N_8840,N_4391,N_5487);
xor U8841 (N_8841,N_6026,N_4584);
and U8842 (N_8842,N_5563,N_4660);
xor U8843 (N_8843,N_3227,N_4865);
nor U8844 (N_8844,N_4845,N_5202);
or U8845 (N_8845,N_5821,N_6119);
nand U8846 (N_8846,N_5942,N_3996);
nand U8847 (N_8847,N_5318,N_4320);
xnor U8848 (N_8848,N_5077,N_4519);
or U8849 (N_8849,N_5992,N_4557);
nand U8850 (N_8850,N_5307,N_6143);
nor U8851 (N_8851,N_6017,N_4337);
and U8852 (N_8852,N_5117,N_4349);
or U8853 (N_8853,N_3622,N_4095);
nor U8854 (N_8854,N_3441,N_4937);
and U8855 (N_8855,N_3912,N_5413);
nand U8856 (N_8856,N_4964,N_4932);
nor U8857 (N_8857,N_5041,N_3591);
nor U8858 (N_8858,N_5592,N_4639);
nand U8859 (N_8859,N_5747,N_5566);
and U8860 (N_8860,N_4914,N_4409);
or U8861 (N_8861,N_4718,N_5158);
nand U8862 (N_8862,N_4077,N_5740);
and U8863 (N_8863,N_3989,N_4458);
and U8864 (N_8864,N_3130,N_5562);
nor U8865 (N_8865,N_5285,N_4657);
or U8866 (N_8866,N_5815,N_6179);
nand U8867 (N_8867,N_3863,N_5906);
or U8868 (N_8868,N_5713,N_5493);
xor U8869 (N_8869,N_5209,N_6168);
or U8870 (N_8870,N_6143,N_5694);
and U8871 (N_8871,N_4662,N_5704);
nor U8872 (N_8872,N_4086,N_3504);
xor U8873 (N_8873,N_6090,N_4536);
and U8874 (N_8874,N_5594,N_4604);
xor U8875 (N_8875,N_5562,N_6050);
nand U8876 (N_8876,N_3405,N_3263);
and U8877 (N_8877,N_3935,N_4793);
and U8878 (N_8878,N_4537,N_3350);
or U8879 (N_8879,N_5080,N_4328);
and U8880 (N_8880,N_4302,N_4566);
nor U8881 (N_8881,N_4944,N_5590);
or U8882 (N_8882,N_3720,N_4231);
xor U8883 (N_8883,N_5722,N_3429);
or U8884 (N_8884,N_4507,N_3226);
nor U8885 (N_8885,N_3344,N_4601);
or U8886 (N_8886,N_5428,N_3626);
nand U8887 (N_8887,N_4570,N_5846);
xor U8888 (N_8888,N_5959,N_3389);
nor U8889 (N_8889,N_3832,N_4280);
nand U8890 (N_8890,N_3592,N_3863);
or U8891 (N_8891,N_5462,N_3389);
nor U8892 (N_8892,N_4687,N_3974);
or U8893 (N_8893,N_4645,N_5868);
xnor U8894 (N_8894,N_4989,N_5265);
or U8895 (N_8895,N_3434,N_6188);
nor U8896 (N_8896,N_5196,N_4039);
nand U8897 (N_8897,N_3441,N_5182);
nor U8898 (N_8898,N_3527,N_3683);
nor U8899 (N_8899,N_3519,N_5244);
xnor U8900 (N_8900,N_5899,N_3367);
nand U8901 (N_8901,N_4398,N_5178);
xor U8902 (N_8902,N_4369,N_3408);
and U8903 (N_8903,N_4372,N_3300);
or U8904 (N_8904,N_4506,N_4337);
xnor U8905 (N_8905,N_3547,N_3607);
nor U8906 (N_8906,N_4009,N_4474);
nand U8907 (N_8907,N_4656,N_5276);
and U8908 (N_8908,N_6206,N_5089);
xor U8909 (N_8909,N_6086,N_4253);
nor U8910 (N_8910,N_3212,N_5786);
xor U8911 (N_8911,N_5256,N_4658);
or U8912 (N_8912,N_6163,N_3448);
or U8913 (N_8913,N_3539,N_3675);
nor U8914 (N_8914,N_3215,N_3768);
nand U8915 (N_8915,N_4328,N_6152);
and U8916 (N_8916,N_5421,N_3229);
or U8917 (N_8917,N_5284,N_4512);
nand U8918 (N_8918,N_4774,N_5572);
nand U8919 (N_8919,N_6030,N_5069);
xor U8920 (N_8920,N_5089,N_5257);
and U8921 (N_8921,N_5969,N_4266);
xnor U8922 (N_8922,N_3484,N_4977);
and U8923 (N_8923,N_4428,N_4504);
nand U8924 (N_8924,N_4383,N_5193);
and U8925 (N_8925,N_4257,N_4996);
xnor U8926 (N_8926,N_4678,N_4821);
xnor U8927 (N_8927,N_5465,N_5517);
nor U8928 (N_8928,N_5639,N_4336);
nand U8929 (N_8929,N_4994,N_3690);
nand U8930 (N_8930,N_3419,N_4974);
or U8931 (N_8931,N_3172,N_4183);
or U8932 (N_8932,N_3355,N_3526);
and U8933 (N_8933,N_3855,N_4150);
nand U8934 (N_8934,N_5574,N_5572);
nand U8935 (N_8935,N_3464,N_4701);
xnor U8936 (N_8936,N_5654,N_3558);
nand U8937 (N_8937,N_6222,N_3473);
xor U8938 (N_8938,N_4720,N_5820);
nor U8939 (N_8939,N_4685,N_5303);
or U8940 (N_8940,N_4746,N_3298);
nand U8941 (N_8941,N_3393,N_5438);
and U8942 (N_8942,N_5539,N_5257);
nor U8943 (N_8943,N_4610,N_5098);
and U8944 (N_8944,N_5025,N_4554);
nor U8945 (N_8945,N_6016,N_5384);
nor U8946 (N_8946,N_5412,N_4016);
and U8947 (N_8947,N_5984,N_5993);
or U8948 (N_8948,N_4488,N_6076);
nor U8949 (N_8949,N_3129,N_4333);
nand U8950 (N_8950,N_5672,N_4676);
xnor U8951 (N_8951,N_6188,N_4051);
and U8952 (N_8952,N_3969,N_3717);
xor U8953 (N_8953,N_4479,N_5155);
or U8954 (N_8954,N_5358,N_3540);
nor U8955 (N_8955,N_3772,N_4610);
nor U8956 (N_8956,N_3725,N_3175);
or U8957 (N_8957,N_3529,N_4093);
and U8958 (N_8958,N_5095,N_3881);
or U8959 (N_8959,N_4940,N_6146);
or U8960 (N_8960,N_3344,N_5074);
nor U8961 (N_8961,N_6106,N_4435);
nand U8962 (N_8962,N_4860,N_3606);
nor U8963 (N_8963,N_3448,N_4029);
and U8964 (N_8964,N_4831,N_5804);
or U8965 (N_8965,N_5941,N_5380);
xor U8966 (N_8966,N_4067,N_5947);
or U8967 (N_8967,N_4478,N_4566);
nor U8968 (N_8968,N_3931,N_3642);
nand U8969 (N_8969,N_4919,N_4072);
nand U8970 (N_8970,N_4256,N_4741);
and U8971 (N_8971,N_5953,N_4499);
nor U8972 (N_8972,N_6075,N_3238);
or U8973 (N_8973,N_3824,N_3815);
xor U8974 (N_8974,N_3203,N_4367);
and U8975 (N_8975,N_5376,N_4517);
nor U8976 (N_8976,N_5467,N_4257);
and U8977 (N_8977,N_5213,N_4149);
nor U8978 (N_8978,N_4537,N_6063);
or U8979 (N_8979,N_3522,N_3892);
nor U8980 (N_8980,N_4701,N_6147);
nor U8981 (N_8981,N_3415,N_5104);
or U8982 (N_8982,N_4942,N_3595);
and U8983 (N_8983,N_4325,N_4815);
nor U8984 (N_8984,N_3838,N_4547);
nor U8985 (N_8985,N_6102,N_3319);
and U8986 (N_8986,N_6185,N_5798);
nand U8987 (N_8987,N_5078,N_4312);
nand U8988 (N_8988,N_3976,N_4951);
nand U8989 (N_8989,N_4093,N_3769);
and U8990 (N_8990,N_5338,N_5942);
nand U8991 (N_8991,N_4583,N_5842);
xor U8992 (N_8992,N_5012,N_5616);
and U8993 (N_8993,N_4609,N_3669);
or U8994 (N_8994,N_5634,N_3136);
nor U8995 (N_8995,N_6216,N_6018);
and U8996 (N_8996,N_3869,N_4163);
nor U8997 (N_8997,N_3551,N_3926);
and U8998 (N_8998,N_4157,N_3200);
xnor U8999 (N_8999,N_4310,N_5582);
nor U9000 (N_9000,N_4220,N_3180);
or U9001 (N_9001,N_3395,N_3991);
or U9002 (N_9002,N_6085,N_6078);
nand U9003 (N_9003,N_3836,N_5584);
nand U9004 (N_9004,N_4299,N_4923);
or U9005 (N_9005,N_5869,N_5700);
xnor U9006 (N_9006,N_4559,N_5907);
or U9007 (N_9007,N_5421,N_3633);
or U9008 (N_9008,N_4133,N_5290);
and U9009 (N_9009,N_6204,N_5364);
nand U9010 (N_9010,N_4512,N_3837);
nor U9011 (N_9011,N_3296,N_3439);
xnor U9012 (N_9012,N_3559,N_3760);
nor U9013 (N_9013,N_5455,N_5262);
nor U9014 (N_9014,N_3746,N_4256);
or U9015 (N_9015,N_5350,N_4831);
and U9016 (N_9016,N_5787,N_5947);
nand U9017 (N_9017,N_5568,N_5680);
nor U9018 (N_9018,N_4340,N_3418);
nand U9019 (N_9019,N_5271,N_4696);
xor U9020 (N_9020,N_3640,N_5414);
nand U9021 (N_9021,N_5154,N_4972);
xor U9022 (N_9022,N_3774,N_5756);
nor U9023 (N_9023,N_5094,N_5610);
nand U9024 (N_9024,N_3848,N_5728);
and U9025 (N_9025,N_3620,N_5494);
nor U9026 (N_9026,N_5992,N_6248);
and U9027 (N_9027,N_3522,N_5118);
nor U9028 (N_9028,N_3332,N_3156);
xnor U9029 (N_9029,N_4541,N_3906);
nor U9030 (N_9030,N_5203,N_4681);
and U9031 (N_9031,N_3541,N_5669);
xnor U9032 (N_9032,N_4153,N_3753);
or U9033 (N_9033,N_4381,N_5558);
nand U9034 (N_9034,N_6248,N_5126);
xor U9035 (N_9035,N_4927,N_3235);
and U9036 (N_9036,N_6228,N_4290);
nor U9037 (N_9037,N_4937,N_5784);
or U9038 (N_9038,N_5395,N_5727);
or U9039 (N_9039,N_5103,N_4330);
nand U9040 (N_9040,N_3792,N_5262);
and U9041 (N_9041,N_5092,N_4172);
and U9042 (N_9042,N_5210,N_4582);
xor U9043 (N_9043,N_4577,N_4124);
xor U9044 (N_9044,N_6074,N_4316);
xnor U9045 (N_9045,N_3600,N_3175);
nor U9046 (N_9046,N_4251,N_4445);
nor U9047 (N_9047,N_5869,N_4512);
and U9048 (N_9048,N_4805,N_6237);
xor U9049 (N_9049,N_4134,N_4171);
nor U9050 (N_9050,N_5832,N_3446);
nand U9051 (N_9051,N_3539,N_5195);
nand U9052 (N_9052,N_4430,N_5768);
nor U9053 (N_9053,N_3575,N_5772);
or U9054 (N_9054,N_3508,N_5214);
and U9055 (N_9055,N_3350,N_5538);
or U9056 (N_9056,N_4213,N_5969);
nor U9057 (N_9057,N_3813,N_3363);
and U9058 (N_9058,N_6231,N_4206);
xnor U9059 (N_9059,N_3271,N_3786);
nor U9060 (N_9060,N_5035,N_5759);
xnor U9061 (N_9061,N_5909,N_5938);
or U9062 (N_9062,N_4267,N_3385);
xor U9063 (N_9063,N_3659,N_6180);
and U9064 (N_9064,N_5626,N_5167);
nor U9065 (N_9065,N_3829,N_6227);
xnor U9066 (N_9066,N_4490,N_5753);
nand U9067 (N_9067,N_5830,N_4254);
nor U9068 (N_9068,N_4311,N_4887);
or U9069 (N_9069,N_5403,N_5217);
xor U9070 (N_9070,N_5311,N_4332);
nand U9071 (N_9071,N_5116,N_3867);
nand U9072 (N_9072,N_4640,N_5795);
and U9073 (N_9073,N_5787,N_4898);
xor U9074 (N_9074,N_5310,N_6009);
xnor U9075 (N_9075,N_5424,N_5321);
xor U9076 (N_9076,N_5633,N_5742);
and U9077 (N_9077,N_3575,N_3564);
xor U9078 (N_9078,N_4966,N_5380);
or U9079 (N_9079,N_5168,N_5526);
xor U9080 (N_9080,N_4824,N_4112);
nor U9081 (N_9081,N_5840,N_3556);
or U9082 (N_9082,N_3486,N_4791);
nor U9083 (N_9083,N_4693,N_4999);
and U9084 (N_9084,N_5786,N_3996);
and U9085 (N_9085,N_5341,N_5122);
or U9086 (N_9086,N_4278,N_4702);
xnor U9087 (N_9087,N_6099,N_4149);
or U9088 (N_9088,N_4832,N_5469);
nor U9089 (N_9089,N_3488,N_4984);
nor U9090 (N_9090,N_3382,N_4538);
nand U9091 (N_9091,N_4764,N_4491);
or U9092 (N_9092,N_4452,N_6026);
xor U9093 (N_9093,N_3653,N_4243);
and U9094 (N_9094,N_5806,N_3492);
nor U9095 (N_9095,N_3781,N_3772);
and U9096 (N_9096,N_5842,N_3974);
and U9097 (N_9097,N_4591,N_5623);
and U9098 (N_9098,N_3978,N_3776);
nand U9099 (N_9099,N_5419,N_4178);
or U9100 (N_9100,N_6093,N_5102);
nor U9101 (N_9101,N_4650,N_3743);
nor U9102 (N_9102,N_5927,N_3900);
or U9103 (N_9103,N_5562,N_3527);
and U9104 (N_9104,N_5614,N_4330);
nor U9105 (N_9105,N_5128,N_3755);
xor U9106 (N_9106,N_5946,N_3724);
xor U9107 (N_9107,N_3486,N_4140);
and U9108 (N_9108,N_5635,N_5904);
or U9109 (N_9109,N_6011,N_3368);
nand U9110 (N_9110,N_3313,N_5357);
nand U9111 (N_9111,N_4316,N_5851);
xnor U9112 (N_9112,N_5527,N_3496);
nand U9113 (N_9113,N_3761,N_4258);
nor U9114 (N_9114,N_5568,N_5455);
xor U9115 (N_9115,N_3769,N_6041);
or U9116 (N_9116,N_3590,N_4620);
nand U9117 (N_9117,N_4009,N_4957);
nand U9118 (N_9118,N_4515,N_3692);
and U9119 (N_9119,N_5869,N_4735);
xnor U9120 (N_9120,N_5798,N_4194);
nand U9121 (N_9121,N_4822,N_4675);
nor U9122 (N_9122,N_6211,N_4046);
nand U9123 (N_9123,N_4559,N_4130);
and U9124 (N_9124,N_4897,N_5340);
nand U9125 (N_9125,N_4632,N_5353);
nor U9126 (N_9126,N_3663,N_5373);
xor U9127 (N_9127,N_3768,N_5047);
nand U9128 (N_9128,N_5278,N_4626);
xor U9129 (N_9129,N_5287,N_3275);
xnor U9130 (N_9130,N_5944,N_6126);
nor U9131 (N_9131,N_3429,N_4271);
and U9132 (N_9132,N_4641,N_4986);
nor U9133 (N_9133,N_5931,N_5669);
or U9134 (N_9134,N_5859,N_5922);
nor U9135 (N_9135,N_3396,N_3989);
nand U9136 (N_9136,N_3223,N_4698);
nand U9137 (N_9137,N_4163,N_5877);
and U9138 (N_9138,N_5808,N_3786);
nand U9139 (N_9139,N_4576,N_3217);
or U9140 (N_9140,N_3528,N_4868);
and U9141 (N_9141,N_4497,N_6139);
xor U9142 (N_9142,N_5322,N_5761);
nand U9143 (N_9143,N_3235,N_5120);
or U9144 (N_9144,N_5943,N_5102);
nor U9145 (N_9145,N_5308,N_3713);
and U9146 (N_9146,N_6167,N_4358);
and U9147 (N_9147,N_5332,N_4584);
nand U9148 (N_9148,N_5258,N_5175);
nand U9149 (N_9149,N_4586,N_6198);
or U9150 (N_9150,N_5302,N_5210);
or U9151 (N_9151,N_6183,N_5609);
nor U9152 (N_9152,N_5850,N_5427);
nor U9153 (N_9153,N_6190,N_5497);
and U9154 (N_9154,N_3848,N_6017);
xor U9155 (N_9155,N_3687,N_5162);
or U9156 (N_9156,N_3561,N_3327);
xnor U9157 (N_9157,N_4803,N_5250);
or U9158 (N_9158,N_3427,N_3932);
and U9159 (N_9159,N_5204,N_3885);
nor U9160 (N_9160,N_3695,N_4080);
xnor U9161 (N_9161,N_3549,N_4263);
xor U9162 (N_9162,N_5409,N_4599);
or U9163 (N_9163,N_5719,N_3471);
nand U9164 (N_9164,N_5903,N_5832);
xor U9165 (N_9165,N_4831,N_5724);
or U9166 (N_9166,N_4844,N_3680);
nor U9167 (N_9167,N_4616,N_6068);
or U9168 (N_9168,N_5722,N_4905);
nand U9169 (N_9169,N_3537,N_3714);
nand U9170 (N_9170,N_3682,N_3339);
xnor U9171 (N_9171,N_3437,N_4473);
and U9172 (N_9172,N_3781,N_5300);
or U9173 (N_9173,N_5406,N_5396);
nor U9174 (N_9174,N_3767,N_6058);
nor U9175 (N_9175,N_6198,N_5536);
xnor U9176 (N_9176,N_6030,N_4321);
nand U9177 (N_9177,N_4705,N_3430);
or U9178 (N_9178,N_5337,N_5453);
xor U9179 (N_9179,N_4947,N_3180);
nand U9180 (N_9180,N_6135,N_4974);
xor U9181 (N_9181,N_5576,N_5298);
nand U9182 (N_9182,N_6173,N_4368);
xor U9183 (N_9183,N_5504,N_5626);
and U9184 (N_9184,N_4095,N_3196);
nand U9185 (N_9185,N_4865,N_4273);
or U9186 (N_9186,N_4621,N_4898);
nor U9187 (N_9187,N_5817,N_4923);
xor U9188 (N_9188,N_4098,N_5472);
and U9189 (N_9189,N_3610,N_3377);
xnor U9190 (N_9190,N_4306,N_5705);
xnor U9191 (N_9191,N_4247,N_4312);
nor U9192 (N_9192,N_5755,N_6052);
or U9193 (N_9193,N_6199,N_4174);
nor U9194 (N_9194,N_6024,N_5778);
and U9195 (N_9195,N_3988,N_5745);
xor U9196 (N_9196,N_5445,N_4356);
and U9197 (N_9197,N_3374,N_4444);
xnor U9198 (N_9198,N_4635,N_5980);
and U9199 (N_9199,N_5401,N_4901);
nor U9200 (N_9200,N_3190,N_4389);
xor U9201 (N_9201,N_5423,N_3445);
xor U9202 (N_9202,N_4993,N_4407);
or U9203 (N_9203,N_5406,N_3557);
nand U9204 (N_9204,N_5652,N_5463);
or U9205 (N_9205,N_4389,N_5691);
or U9206 (N_9206,N_5765,N_5501);
and U9207 (N_9207,N_3293,N_5427);
and U9208 (N_9208,N_3929,N_5010);
nor U9209 (N_9209,N_5914,N_4746);
nor U9210 (N_9210,N_4858,N_5950);
xnor U9211 (N_9211,N_3881,N_5464);
nor U9212 (N_9212,N_5421,N_4371);
and U9213 (N_9213,N_5282,N_4986);
nand U9214 (N_9214,N_5526,N_4154);
nor U9215 (N_9215,N_6228,N_3307);
or U9216 (N_9216,N_5878,N_5733);
or U9217 (N_9217,N_5813,N_4108);
nand U9218 (N_9218,N_5659,N_3892);
and U9219 (N_9219,N_4555,N_4269);
or U9220 (N_9220,N_6157,N_4693);
xor U9221 (N_9221,N_3356,N_5127);
xnor U9222 (N_9222,N_5847,N_3529);
nand U9223 (N_9223,N_4572,N_4238);
xor U9224 (N_9224,N_3321,N_6218);
and U9225 (N_9225,N_5065,N_5709);
nand U9226 (N_9226,N_5008,N_6106);
xnor U9227 (N_9227,N_4116,N_3637);
nor U9228 (N_9228,N_3257,N_3217);
or U9229 (N_9229,N_3485,N_3566);
xor U9230 (N_9230,N_4516,N_4013);
nand U9231 (N_9231,N_4261,N_5531);
nand U9232 (N_9232,N_4762,N_3906);
and U9233 (N_9233,N_3429,N_3458);
nor U9234 (N_9234,N_4097,N_5459);
and U9235 (N_9235,N_5502,N_4062);
nand U9236 (N_9236,N_4378,N_5298);
nand U9237 (N_9237,N_3832,N_5933);
nand U9238 (N_9238,N_3791,N_5524);
xor U9239 (N_9239,N_3819,N_3228);
nand U9240 (N_9240,N_4173,N_5978);
nor U9241 (N_9241,N_3195,N_3260);
and U9242 (N_9242,N_5974,N_5679);
and U9243 (N_9243,N_5187,N_6087);
xnor U9244 (N_9244,N_4072,N_5850);
nor U9245 (N_9245,N_4810,N_5582);
and U9246 (N_9246,N_4499,N_4680);
or U9247 (N_9247,N_6196,N_5977);
and U9248 (N_9248,N_3374,N_3355);
nand U9249 (N_9249,N_5679,N_6192);
and U9250 (N_9250,N_4087,N_3708);
xor U9251 (N_9251,N_3694,N_6025);
or U9252 (N_9252,N_3719,N_4127);
xor U9253 (N_9253,N_5705,N_3881);
nand U9254 (N_9254,N_5551,N_3544);
and U9255 (N_9255,N_3167,N_5077);
or U9256 (N_9256,N_4617,N_4761);
nor U9257 (N_9257,N_3627,N_3282);
and U9258 (N_9258,N_5118,N_5325);
nor U9259 (N_9259,N_4126,N_3997);
xnor U9260 (N_9260,N_4324,N_4820);
or U9261 (N_9261,N_3578,N_4147);
xor U9262 (N_9262,N_4956,N_5758);
or U9263 (N_9263,N_5642,N_5996);
xnor U9264 (N_9264,N_4898,N_5535);
xnor U9265 (N_9265,N_4048,N_6094);
xnor U9266 (N_9266,N_3302,N_4891);
and U9267 (N_9267,N_5983,N_4280);
and U9268 (N_9268,N_5693,N_4956);
nor U9269 (N_9269,N_3263,N_3657);
or U9270 (N_9270,N_4285,N_4956);
and U9271 (N_9271,N_3707,N_5413);
nand U9272 (N_9272,N_3424,N_4120);
xnor U9273 (N_9273,N_5986,N_3636);
or U9274 (N_9274,N_3133,N_4858);
nand U9275 (N_9275,N_3373,N_4332);
and U9276 (N_9276,N_5252,N_3400);
or U9277 (N_9277,N_5505,N_4394);
xnor U9278 (N_9278,N_4522,N_4520);
and U9279 (N_9279,N_3278,N_4112);
xnor U9280 (N_9280,N_3565,N_3344);
xnor U9281 (N_9281,N_4913,N_3957);
nand U9282 (N_9282,N_6176,N_5467);
or U9283 (N_9283,N_3560,N_3818);
xor U9284 (N_9284,N_4451,N_4906);
or U9285 (N_9285,N_3362,N_5248);
xnor U9286 (N_9286,N_6132,N_4453);
nand U9287 (N_9287,N_4380,N_4210);
and U9288 (N_9288,N_4941,N_3462);
nor U9289 (N_9289,N_4446,N_4748);
nor U9290 (N_9290,N_5603,N_5412);
xor U9291 (N_9291,N_3703,N_5122);
nand U9292 (N_9292,N_4955,N_3478);
or U9293 (N_9293,N_4053,N_5863);
or U9294 (N_9294,N_5745,N_3252);
nor U9295 (N_9295,N_4659,N_5447);
and U9296 (N_9296,N_6236,N_4473);
or U9297 (N_9297,N_5081,N_6031);
or U9298 (N_9298,N_5909,N_4214);
or U9299 (N_9299,N_6000,N_4032);
and U9300 (N_9300,N_5268,N_3531);
nor U9301 (N_9301,N_5738,N_3459);
nand U9302 (N_9302,N_4207,N_6006);
xnor U9303 (N_9303,N_5694,N_4993);
nand U9304 (N_9304,N_5838,N_5409);
or U9305 (N_9305,N_5478,N_4704);
nand U9306 (N_9306,N_4492,N_5611);
nand U9307 (N_9307,N_3343,N_4359);
or U9308 (N_9308,N_6132,N_3186);
or U9309 (N_9309,N_4767,N_6088);
xnor U9310 (N_9310,N_6058,N_3463);
xor U9311 (N_9311,N_5186,N_4815);
or U9312 (N_9312,N_5976,N_3209);
xnor U9313 (N_9313,N_3983,N_4629);
and U9314 (N_9314,N_5201,N_5570);
and U9315 (N_9315,N_5119,N_6190);
and U9316 (N_9316,N_4880,N_5608);
and U9317 (N_9317,N_3984,N_4520);
xnor U9318 (N_9318,N_5999,N_5258);
nor U9319 (N_9319,N_6230,N_3475);
and U9320 (N_9320,N_4848,N_3787);
nor U9321 (N_9321,N_4015,N_4368);
or U9322 (N_9322,N_3684,N_6231);
xnor U9323 (N_9323,N_4395,N_4257);
and U9324 (N_9324,N_6064,N_4080);
nand U9325 (N_9325,N_6008,N_5961);
or U9326 (N_9326,N_4826,N_3879);
xnor U9327 (N_9327,N_4343,N_5512);
nor U9328 (N_9328,N_5567,N_5327);
nand U9329 (N_9329,N_4212,N_5778);
or U9330 (N_9330,N_4198,N_4571);
and U9331 (N_9331,N_3812,N_3698);
or U9332 (N_9332,N_4748,N_6140);
nand U9333 (N_9333,N_3310,N_4770);
and U9334 (N_9334,N_5482,N_5607);
nor U9335 (N_9335,N_4305,N_3251);
or U9336 (N_9336,N_6133,N_4155);
nor U9337 (N_9337,N_3186,N_4291);
and U9338 (N_9338,N_4695,N_5234);
nand U9339 (N_9339,N_5604,N_4209);
nor U9340 (N_9340,N_4269,N_4609);
nor U9341 (N_9341,N_3253,N_3516);
xnor U9342 (N_9342,N_3538,N_5318);
nor U9343 (N_9343,N_3566,N_5006);
and U9344 (N_9344,N_5279,N_3694);
or U9345 (N_9345,N_4243,N_3174);
xnor U9346 (N_9346,N_3327,N_3798);
nor U9347 (N_9347,N_4497,N_3772);
and U9348 (N_9348,N_4425,N_6077);
and U9349 (N_9349,N_6155,N_3608);
or U9350 (N_9350,N_4663,N_4617);
xnor U9351 (N_9351,N_5806,N_6076);
nor U9352 (N_9352,N_3175,N_5852);
xor U9353 (N_9353,N_5193,N_4187);
xnor U9354 (N_9354,N_5490,N_5608);
xor U9355 (N_9355,N_5793,N_3417);
and U9356 (N_9356,N_4266,N_3348);
xnor U9357 (N_9357,N_3361,N_5633);
nand U9358 (N_9358,N_3410,N_6036);
and U9359 (N_9359,N_5138,N_5952);
nor U9360 (N_9360,N_6042,N_5421);
nor U9361 (N_9361,N_5153,N_3348);
or U9362 (N_9362,N_5729,N_5161);
and U9363 (N_9363,N_4794,N_4850);
or U9364 (N_9364,N_5626,N_4229);
and U9365 (N_9365,N_4884,N_4983);
or U9366 (N_9366,N_3459,N_3138);
and U9367 (N_9367,N_5760,N_5906);
xnor U9368 (N_9368,N_4531,N_6193);
or U9369 (N_9369,N_3881,N_3555);
xnor U9370 (N_9370,N_5221,N_4186);
and U9371 (N_9371,N_4538,N_3349);
or U9372 (N_9372,N_4222,N_3148);
nand U9373 (N_9373,N_5845,N_5670);
and U9374 (N_9374,N_3910,N_5488);
nor U9375 (N_9375,N_8937,N_7848);
nand U9376 (N_9376,N_9121,N_6853);
nor U9377 (N_9377,N_6384,N_6928);
nor U9378 (N_9378,N_8274,N_6849);
and U9379 (N_9379,N_8970,N_8050);
or U9380 (N_9380,N_7884,N_7595);
and U9381 (N_9381,N_6885,N_8989);
nand U9382 (N_9382,N_8422,N_8960);
nand U9383 (N_9383,N_6336,N_7210);
and U9384 (N_9384,N_6924,N_8961);
or U9385 (N_9385,N_8327,N_7394);
xor U9386 (N_9386,N_8882,N_8218);
or U9387 (N_9387,N_7347,N_6338);
nor U9388 (N_9388,N_8753,N_7203);
xor U9389 (N_9389,N_9160,N_7546);
nand U9390 (N_9390,N_8527,N_8235);
nand U9391 (N_9391,N_7915,N_6567);
or U9392 (N_9392,N_7752,N_8959);
and U9393 (N_9393,N_6960,N_7312);
xor U9394 (N_9394,N_8483,N_7531);
nand U9395 (N_9395,N_6882,N_8906);
nor U9396 (N_9396,N_7651,N_7891);
or U9397 (N_9397,N_6592,N_8522);
nand U9398 (N_9398,N_8369,N_7042);
xor U9399 (N_9399,N_6827,N_9130);
nor U9400 (N_9400,N_8407,N_8975);
and U9401 (N_9401,N_8087,N_6536);
or U9402 (N_9402,N_6324,N_6902);
nor U9403 (N_9403,N_6999,N_9374);
and U9404 (N_9404,N_7188,N_6441);
nand U9405 (N_9405,N_8197,N_6252);
or U9406 (N_9406,N_8063,N_9247);
nor U9407 (N_9407,N_8652,N_8557);
nor U9408 (N_9408,N_7068,N_6780);
or U9409 (N_9409,N_7348,N_6971);
xor U9410 (N_9410,N_6843,N_7942);
xnor U9411 (N_9411,N_6740,N_8449);
or U9412 (N_9412,N_7716,N_6758);
or U9413 (N_9413,N_6713,N_7467);
xnor U9414 (N_9414,N_8699,N_6491);
nor U9415 (N_9415,N_7742,N_9353);
and U9416 (N_9416,N_8356,N_8328);
nor U9417 (N_9417,N_6301,N_6719);
nand U9418 (N_9418,N_8592,N_7382);
nand U9419 (N_9419,N_8284,N_8894);
and U9420 (N_9420,N_8568,N_9307);
nor U9421 (N_9421,N_7237,N_7196);
nand U9422 (N_9422,N_8459,N_6275);
nand U9423 (N_9423,N_8291,N_7634);
nor U9424 (N_9424,N_9313,N_6907);
or U9425 (N_9425,N_8554,N_7044);
and U9426 (N_9426,N_6285,N_9032);
and U9427 (N_9427,N_9324,N_9286);
and U9428 (N_9428,N_7316,N_9285);
or U9429 (N_9429,N_7500,N_8084);
or U9430 (N_9430,N_7153,N_7739);
or U9431 (N_9431,N_9170,N_7217);
and U9432 (N_9432,N_9188,N_9345);
nor U9433 (N_9433,N_7853,N_9097);
and U9434 (N_9434,N_7714,N_8768);
xnor U9435 (N_9435,N_6998,N_7048);
or U9436 (N_9436,N_7779,N_7307);
nor U9437 (N_9437,N_7137,N_8175);
xor U9438 (N_9438,N_8412,N_8021);
nand U9439 (N_9439,N_9262,N_6559);
or U9440 (N_9440,N_7588,N_9323);
and U9441 (N_9441,N_7116,N_7402);
nand U9442 (N_9442,N_7285,N_7940);
nand U9443 (N_9443,N_7232,N_8132);
and U9444 (N_9444,N_7579,N_8386);
nand U9445 (N_9445,N_8897,N_7882);
nand U9446 (N_9446,N_9151,N_7009);
xnor U9447 (N_9447,N_8129,N_7379);
nor U9448 (N_9448,N_6817,N_8671);
and U9449 (N_9449,N_7252,N_7168);
or U9450 (N_9450,N_8865,N_7087);
or U9451 (N_9451,N_6577,N_7273);
xor U9452 (N_9452,N_8102,N_8619);
or U9453 (N_9453,N_6271,N_6553);
nor U9454 (N_9454,N_9108,N_6564);
xnor U9455 (N_9455,N_8280,N_7064);
nand U9456 (N_9456,N_6445,N_8228);
nand U9457 (N_9457,N_6506,N_8501);
or U9458 (N_9458,N_8822,N_6593);
nand U9459 (N_9459,N_8012,N_6693);
or U9460 (N_9460,N_8874,N_7350);
or U9461 (N_9461,N_6478,N_6305);
xnor U9462 (N_9462,N_6905,N_6258);
and U9463 (N_9463,N_7002,N_7615);
nor U9464 (N_9464,N_7099,N_8016);
and U9465 (N_9465,N_6594,N_9265);
or U9466 (N_9466,N_8342,N_7338);
and U9467 (N_9467,N_8775,N_6666);
nor U9468 (N_9468,N_9341,N_9318);
xnor U9469 (N_9469,N_8672,N_7280);
nor U9470 (N_9470,N_8635,N_7695);
xnor U9471 (N_9471,N_8582,N_8643);
nor U9472 (N_9472,N_7559,N_9009);
or U9473 (N_9473,N_7731,N_8073);
nand U9474 (N_9474,N_8831,N_6661);
nand U9475 (N_9475,N_8437,N_8622);
nand U9476 (N_9476,N_8337,N_6634);
or U9477 (N_9477,N_8921,N_9225);
nor U9478 (N_9478,N_8811,N_8880);
or U9479 (N_9479,N_7664,N_8944);
nor U9480 (N_9480,N_7767,N_7907);
xor U9481 (N_9481,N_7992,N_9146);
xnor U9482 (N_9482,N_7981,N_7341);
or U9483 (N_9483,N_6379,N_8697);
and U9484 (N_9484,N_6997,N_6936);
and U9485 (N_9485,N_8787,N_9276);
nor U9486 (N_9486,N_8268,N_7233);
or U9487 (N_9487,N_6408,N_6763);
or U9488 (N_9488,N_8227,N_6462);
nand U9489 (N_9489,N_8067,N_8427);
and U9490 (N_9490,N_6565,N_7735);
xor U9491 (N_9491,N_7246,N_7673);
nand U9492 (N_9492,N_7791,N_7620);
nor U9493 (N_9493,N_8154,N_7671);
xor U9494 (N_9494,N_7386,N_6818);
nor U9495 (N_9495,N_7310,N_7287);
nor U9496 (N_9496,N_9366,N_9205);
and U9497 (N_9497,N_7163,N_8692);
or U9498 (N_9498,N_8322,N_7461);
or U9499 (N_9499,N_7425,N_9252);
xor U9500 (N_9500,N_7961,N_6814);
nor U9501 (N_9501,N_7570,N_6720);
xor U9502 (N_9502,N_7100,N_8372);
nor U9503 (N_9503,N_7846,N_9005);
and U9504 (N_9504,N_7096,N_7337);
nand U9505 (N_9505,N_6953,N_9199);
nand U9506 (N_9506,N_7950,N_6291);
and U9507 (N_9507,N_6544,N_8763);
nand U9508 (N_9508,N_9254,N_8898);
xnor U9509 (N_9509,N_6304,N_9042);
xnor U9510 (N_9510,N_9350,N_8296);
nor U9511 (N_9511,N_6516,N_8998);
nand U9512 (N_9512,N_7880,N_6345);
xnor U9513 (N_9513,N_9292,N_8347);
nor U9514 (N_9514,N_8077,N_9166);
nand U9515 (N_9515,N_8172,N_7229);
nor U9516 (N_9516,N_6606,N_7085);
nor U9517 (N_9517,N_9371,N_7383);
nand U9518 (N_9518,N_8444,N_8247);
xnor U9519 (N_9519,N_6829,N_6947);
and U9520 (N_9520,N_6630,N_8840);
or U9521 (N_9521,N_8443,N_9145);
and U9522 (N_9522,N_7244,N_8148);
xnor U9523 (N_9523,N_8118,N_7655);
nand U9524 (N_9524,N_8758,N_8955);
xor U9525 (N_9525,N_8976,N_9361);
nor U9526 (N_9526,N_8595,N_6812);
or U9527 (N_9527,N_8720,N_8552);
xor U9528 (N_9528,N_8942,N_7984);
nor U9529 (N_9529,N_6357,N_6628);
nand U9530 (N_9530,N_8425,N_7335);
xor U9531 (N_9531,N_6671,N_8694);
nor U9532 (N_9532,N_6958,N_9331);
or U9533 (N_9533,N_8168,N_9141);
xnor U9534 (N_9534,N_6311,N_9217);
or U9535 (N_9535,N_6471,N_9048);
or U9536 (N_9536,N_8515,N_8233);
and U9537 (N_9537,N_6522,N_8415);
or U9538 (N_9538,N_8001,N_7737);
and U9539 (N_9539,N_6648,N_7759);
or U9540 (N_9540,N_6312,N_9024);
nand U9541 (N_9541,N_7859,N_8588);
nand U9542 (N_9542,N_9260,N_6844);
and U9543 (N_9543,N_7231,N_9190);
xor U9544 (N_9544,N_6281,N_7870);
nor U9545 (N_9545,N_6932,N_8778);
xor U9546 (N_9546,N_6691,N_6868);
nand U9547 (N_9547,N_6317,N_6543);
nor U9548 (N_9548,N_6860,N_6439);
xnor U9549 (N_9549,N_7303,N_8690);
nand U9550 (N_9550,N_7200,N_7052);
and U9551 (N_9551,N_7705,N_6508);
nor U9552 (N_9552,N_8941,N_8518);
nand U9553 (N_9553,N_9177,N_7957);
or U9554 (N_9554,N_9129,N_6857);
or U9555 (N_9555,N_6854,N_7076);
nor U9556 (N_9556,N_9301,N_9279);
nor U9557 (N_9557,N_6485,N_7575);
and U9558 (N_9558,N_9251,N_8452);
nand U9559 (N_9559,N_6383,N_8004);
or U9560 (N_9560,N_7165,N_6802);
and U9561 (N_9561,N_8508,N_9191);
or U9562 (N_9562,N_7783,N_7998);
and U9563 (N_9563,N_6475,N_9155);
xor U9564 (N_9564,N_7612,N_7888);
xor U9565 (N_9565,N_8761,N_6764);
nand U9566 (N_9566,N_6529,N_6514);
nor U9567 (N_9567,N_7840,N_7360);
nor U9568 (N_9568,N_9359,N_9369);
nor U9569 (N_9569,N_6406,N_8473);
or U9570 (N_9570,N_6526,N_7352);
nand U9571 (N_9571,N_7486,N_6443);
or U9572 (N_9572,N_6956,N_7972);
xnor U9573 (N_9573,N_9072,N_8752);
or U9574 (N_9574,N_9302,N_6315);
and U9575 (N_9575,N_7283,N_9104);
nand U9576 (N_9576,N_6783,N_7452);
or U9577 (N_9577,N_6959,N_6675);
or U9578 (N_9578,N_8948,N_8082);
nor U9579 (N_9579,N_8376,N_7922);
nand U9580 (N_9580,N_8361,N_6869);
or U9581 (N_9581,N_8613,N_7679);
and U9582 (N_9582,N_7920,N_6512);
xnor U9583 (N_9583,N_7806,N_7581);
and U9584 (N_9584,N_8185,N_7154);
nor U9585 (N_9585,N_9028,N_6663);
xor U9586 (N_9586,N_9185,N_6389);
xnor U9587 (N_9587,N_8278,N_7496);
nand U9588 (N_9588,N_7063,N_8302);
nand U9589 (N_9589,N_8064,N_9117);
or U9590 (N_9590,N_7158,N_7953);
xor U9591 (N_9591,N_7417,N_8032);
xor U9592 (N_9592,N_6294,N_8236);
xnor U9593 (N_9593,N_9106,N_7462);
nor U9594 (N_9594,N_7430,N_7230);
and U9595 (N_9595,N_6979,N_7123);
or U9596 (N_9596,N_7276,N_9221);
or U9597 (N_9597,N_8325,N_7794);
xor U9598 (N_9598,N_7369,N_8266);
nor U9599 (N_9599,N_8027,N_7666);
or U9600 (N_9600,N_6468,N_7808);
nand U9601 (N_9601,N_6912,N_7811);
xor U9602 (N_9602,N_8769,N_9314);
nand U9603 (N_9603,N_7120,N_7242);
nand U9604 (N_9604,N_7647,N_8928);
nand U9605 (N_9605,N_8782,N_8277);
and U9606 (N_9606,N_7008,N_6296);
nor U9607 (N_9607,N_7440,N_7975);
and U9608 (N_9608,N_6450,N_8366);
nor U9609 (N_9609,N_6431,N_7195);
nor U9610 (N_9610,N_7562,N_7066);
or U9611 (N_9611,N_8910,N_7224);
nor U9612 (N_9612,N_8226,N_7684);
nand U9613 (N_9613,N_6641,N_6741);
and U9614 (N_9614,N_7499,N_7091);
xor U9615 (N_9615,N_6795,N_8124);
or U9616 (N_9616,N_8585,N_8204);
xor U9617 (N_9617,N_7751,N_7807);
xnor U9618 (N_9618,N_6569,N_6284);
xor U9619 (N_9619,N_8086,N_8377);
nor U9620 (N_9620,N_8355,N_6974);
xnor U9621 (N_9621,N_6388,N_7512);
and U9622 (N_9622,N_8661,N_8640);
xnor U9623 (N_9623,N_7162,N_9256);
nand U9624 (N_9624,N_8137,N_6801);
nand U9625 (N_9625,N_6323,N_8288);
nor U9626 (N_9626,N_9334,N_6303);
or U9627 (N_9627,N_7175,N_8162);
nor U9628 (N_9628,N_6415,N_7646);
xnor U9629 (N_9629,N_6405,N_6267);
nand U9630 (N_9630,N_6697,N_8287);
xnor U9631 (N_9631,N_8112,N_7326);
nand U9632 (N_9632,N_6263,N_8789);
nand U9633 (N_9633,N_9149,N_7243);
and U9634 (N_9634,N_7334,N_8859);
and U9635 (N_9635,N_9243,N_9278);
and U9636 (N_9636,N_6841,N_6626);
xnor U9637 (N_9637,N_7970,N_6609);
nor U9638 (N_9638,N_8191,N_7994);
nand U9639 (N_9639,N_9362,N_7182);
nand U9640 (N_9640,N_6807,N_6957);
xor U9641 (N_9641,N_7962,N_6743);
xor U9642 (N_9642,N_8974,N_8923);
nand U9643 (N_9643,N_8825,N_9241);
nand U9644 (N_9644,N_8035,N_6699);
nand U9645 (N_9645,N_9158,N_8860);
or U9646 (N_9646,N_7327,N_8591);
nand U9647 (N_9647,N_7368,N_8007);
and U9648 (N_9648,N_7543,N_8349);
or U9649 (N_9649,N_7306,N_8419);
or U9650 (N_9650,N_7223,N_6799);
and U9651 (N_9651,N_7995,N_8780);
nand U9652 (N_9652,N_8766,N_8359);
nor U9653 (N_9653,N_8065,N_8094);
nand U9654 (N_9654,N_8621,N_7477);
nand U9655 (N_9655,N_8754,N_6550);
nand U9656 (N_9656,N_8712,N_9264);
nor U9657 (N_9657,N_9257,N_8649);
and U9658 (N_9658,N_9337,N_8790);
nor U9659 (N_9659,N_8156,N_8547);
and U9660 (N_9660,N_6989,N_6749);
nor U9661 (N_9661,N_8890,N_8827);
xor U9662 (N_9662,N_7221,N_9330);
xor U9663 (N_9663,N_8237,N_6916);
xnor U9664 (N_9664,N_8187,N_8584);
nand U9665 (N_9665,N_8441,N_9184);
and U9666 (N_9666,N_8866,N_7411);
nor U9667 (N_9667,N_9290,N_7112);
nand U9668 (N_9668,N_6386,N_7340);
nand U9669 (N_9669,N_7007,N_8549);
nor U9670 (N_9670,N_8949,N_8689);
xnor U9671 (N_9671,N_7429,N_7713);
and U9672 (N_9672,N_8988,N_8855);
or U9673 (N_9673,N_7375,N_6921);
nand U9674 (N_9674,N_6861,N_6422);
xnor U9675 (N_9675,N_9201,N_6488);
nor U9676 (N_9676,N_6880,N_6419);
nand U9677 (N_9677,N_6694,N_8160);
nor U9678 (N_9678,N_7792,N_7226);
xnor U9679 (N_9679,N_8996,N_9136);
xnor U9680 (N_9680,N_7032,N_9019);
nor U9681 (N_9681,N_7171,N_9275);
nor U9682 (N_9682,N_6401,N_8310);
or U9683 (N_9683,N_7687,N_7463);
nand U9684 (N_9684,N_6341,N_9312);
or U9685 (N_9685,N_8269,N_6629);
xnor U9686 (N_9686,N_8543,N_7480);
and U9687 (N_9687,N_6253,N_7979);
nor U9688 (N_9688,N_6310,N_7895);
or U9689 (N_9689,N_8106,N_9063);
nor U9690 (N_9690,N_8755,N_8646);
nand U9691 (N_9691,N_7639,N_6403);
and U9692 (N_9692,N_7189,N_9043);
and U9693 (N_9693,N_7835,N_7427);
or U9694 (N_9694,N_7134,N_8757);
or U9695 (N_9695,N_6446,N_6931);
nand U9696 (N_9696,N_8911,N_8678);
or U9697 (N_9697,N_8668,N_8290);
nand U9698 (N_9698,N_6266,N_8696);
nor U9699 (N_9699,N_8079,N_8177);
nand U9700 (N_9700,N_8215,N_7321);
nand U9701 (N_9701,N_7997,N_7569);
or U9702 (N_9702,N_6993,N_7143);
nand U9703 (N_9703,N_6600,N_7865);
nor U9704 (N_9704,N_6494,N_7589);
nand U9705 (N_9705,N_7667,N_8326);
and U9706 (N_9706,N_6788,N_7260);
or U9707 (N_9707,N_7024,N_7636);
and U9708 (N_9708,N_8194,N_8428);
nand U9709 (N_9709,N_6973,N_7017);
or U9710 (N_9710,N_6917,N_8273);
and U9711 (N_9711,N_7552,N_6346);
xor U9712 (N_9712,N_8492,N_7109);
or U9713 (N_9713,N_7057,N_8511);
or U9714 (N_9714,N_8371,N_7625);
nand U9715 (N_9715,N_8963,N_8465);
nor U9716 (N_9716,N_6988,N_7917);
or U9717 (N_9717,N_6903,N_8301);
and U9718 (N_9718,N_8935,N_7385);
xnor U9719 (N_9719,N_8157,N_8275);
and U9720 (N_9720,N_6487,N_7353);
or U9721 (N_9721,N_6887,N_6520);
nor U9722 (N_9722,N_8623,N_8135);
and U9723 (N_9723,N_8940,N_7799);
nor U9724 (N_9724,N_9046,N_8122);
nor U9725 (N_9725,N_7263,N_7339);
or U9726 (N_9726,N_7180,N_8479);
and U9727 (N_9727,N_7088,N_7094);
or U9728 (N_9728,N_9053,N_8489);
nor U9729 (N_9729,N_7645,N_9013);
xor U9730 (N_9730,N_6654,N_8389);
and U9731 (N_9731,N_8017,N_7756);
and U9732 (N_9732,N_7851,N_6704);
nand U9733 (N_9733,N_7305,N_7935);
nor U9734 (N_9734,N_7839,N_7689);
nor U9735 (N_9735,N_8872,N_8715);
or U9736 (N_9736,N_9189,N_8971);
xnor U9737 (N_9737,N_8926,N_6748);
and U9738 (N_9738,N_7003,N_9029);
or U9739 (N_9739,N_7373,N_8048);
nand U9740 (N_9740,N_8219,N_8812);
nand U9741 (N_9741,N_7801,N_6963);
nand U9742 (N_9742,N_6874,N_7278);
xor U9743 (N_9743,N_7971,N_8297);
xnor U9744 (N_9744,N_8128,N_7358);
or U9745 (N_9745,N_6863,N_6413);
xor U9746 (N_9746,N_9233,N_6725);
xnor U9747 (N_9747,N_7660,N_7146);
nor U9748 (N_9748,N_8282,N_8517);
nor U9749 (N_9749,N_9325,N_6679);
nor U9750 (N_9750,N_8009,N_7771);
nor U9751 (N_9751,N_7184,N_6709);
nand U9752 (N_9752,N_6798,N_7604);
nand U9753 (N_9753,N_7758,N_9015);
and U9754 (N_9754,N_6562,N_6673);
or U9755 (N_9755,N_7897,N_8136);
and U9756 (N_9756,N_9351,N_7185);
and U9757 (N_9757,N_7055,N_6632);
xor U9758 (N_9758,N_8630,N_9213);
nor U9759 (N_9759,N_8446,N_8388);
and U9760 (N_9760,N_8817,N_6615);
nand U9761 (N_9761,N_8184,N_6394);
or U9762 (N_9762,N_6968,N_9234);
or U9763 (N_9763,N_8411,N_7867);
nor U9764 (N_9764,N_6940,N_7471);
or U9765 (N_9765,N_8597,N_8615);
or U9766 (N_9766,N_8934,N_8662);
or U9767 (N_9767,N_6273,N_6366);
xnor U9768 (N_9768,N_6608,N_7495);
nor U9769 (N_9769,N_7700,N_8829);
nand U9770 (N_9770,N_8406,N_7843);
and U9771 (N_9771,N_7147,N_6333);
or U9772 (N_9772,N_7124,N_7565);
nand U9773 (N_9773,N_8564,N_7852);
nand U9774 (N_9774,N_8113,N_6256);
or U9775 (N_9775,N_6762,N_8313);
nor U9776 (N_9776,N_7643,N_9332);
nor U9777 (N_9777,N_7138,N_7072);
xor U9778 (N_9778,N_8555,N_8445);
and U9779 (N_9779,N_7193,N_7857);
xnor U9780 (N_9780,N_7026,N_8498);
and U9781 (N_9781,N_9085,N_7789);
or U9782 (N_9782,N_9127,N_6352);
nand U9783 (N_9783,N_6436,N_9171);
and U9784 (N_9784,N_6250,N_7458);
nor U9785 (N_9785,N_8503,N_6635);
or U9786 (N_9786,N_6778,N_6847);
or U9787 (N_9787,N_8793,N_8464);
and U9788 (N_9788,N_7381,N_8059);
or U9789 (N_9789,N_6686,N_9088);
and U9790 (N_9790,N_9195,N_8045);
or U9791 (N_9791,N_8861,N_7431);
and U9792 (N_9792,N_8138,N_8056);
and U9793 (N_9793,N_8131,N_9220);
and U9794 (N_9794,N_6942,N_8693);
and U9795 (N_9795,N_8442,N_8058);
and U9796 (N_9796,N_8206,N_9354);
nor U9797 (N_9797,N_8466,N_8256);
nor U9798 (N_9798,N_8022,N_6604);
xnor U9799 (N_9799,N_7564,N_7762);
or U9800 (N_9800,N_6913,N_7934);
or U9801 (N_9801,N_6325,N_8270);
and U9802 (N_9802,N_6919,N_9102);
and U9803 (N_9803,N_6385,N_8783);
xnor U9804 (N_9804,N_7568,N_8691);
and U9805 (N_9805,N_7628,N_7019);
nor U9806 (N_9806,N_7421,N_7412);
or U9807 (N_9807,N_8913,N_9211);
xor U9808 (N_9808,N_7904,N_7557);
or U9809 (N_9809,N_7028,N_8977);
nor U9810 (N_9810,N_8494,N_6850);
xnor U9811 (N_9811,N_8669,N_8516);
xnor U9812 (N_9812,N_8026,N_8309);
and U9813 (N_9813,N_8216,N_6257);
nor U9814 (N_9814,N_7982,N_6918);
or U9815 (N_9815,N_8895,N_9197);
and U9816 (N_9816,N_9230,N_8777);
or U9817 (N_9817,N_6486,N_7038);
nand U9818 (N_9818,N_7308,N_7874);
nand U9819 (N_9819,N_6546,N_8809);
and U9820 (N_9820,N_6731,N_8920);
xnor U9821 (N_9821,N_8900,N_6994);
nor U9822 (N_9822,N_6915,N_7111);
nand U9823 (N_9823,N_8545,N_8510);
and U9824 (N_9824,N_6347,N_6852);
and U9825 (N_9825,N_7602,N_7558);
xor U9826 (N_9826,N_6750,N_8736);
nor U9827 (N_9827,N_8765,N_7067);
xor U9828 (N_9828,N_8011,N_8727);
xnor U9829 (N_9829,N_7649,N_6706);
nor U9830 (N_9830,N_8409,N_8606);
nor U9831 (N_9831,N_8565,N_9316);
or U9832 (N_9832,N_7130,N_7034);
xor U9833 (N_9833,N_7551,N_6888);
or U9834 (N_9834,N_7760,N_7618);
nand U9835 (N_9835,N_6734,N_7344);
and U9836 (N_9836,N_8468,N_7419);
or U9837 (N_9837,N_6356,N_6566);
nand U9838 (N_9838,N_7355,N_8467);
nand U9839 (N_9839,N_7033,N_6644);
nor U9840 (N_9840,N_6779,N_8375);
xnor U9841 (N_9841,N_6484,N_8097);
nor U9842 (N_9842,N_6745,N_7816);
nand U9843 (N_9843,N_8312,N_7489);
or U9844 (N_9844,N_7747,N_9250);
and U9845 (N_9845,N_7483,N_7030);
nor U9846 (N_9846,N_8719,N_8364);
nor U9847 (N_9847,N_8474,N_9087);
or U9848 (N_9848,N_6705,N_7626);
nor U9849 (N_9849,N_7723,N_7554);
xor U9850 (N_9850,N_6738,N_9216);
or U9851 (N_9851,N_8810,N_8524);
nor U9852 (N_9852,N_8458,N_7613);
xnor U9853 (N_9853,N_8749,N_8987);
or U9854 (N_9854,N_8487,N_8253);
and U9855 (N_9855,N_7528,N_7459);
or U9856 (N_9856,N_6752,N_8519);
xnor U9857 (N_9857,N_7608,N_7715);
nand U9858 (N_9858,N_8319,N_8573);
and U9859 (N_9859,N_7240,N_6714);
nand U9860 (N_9860,N_8805,N_8847);
and U9861 (N_9861,N_8907,N_8330);
nor U9862 (N_9862,N_7600,N_7491);
or U9863 (N_9863,N_8841,N_8682);
xor U9864 (N_9864,N_7782,N_7829);
xnor U9865 (N_9865,N_6339,N_7343);
or U9866 (N_9866,N_8701,N_8387);
nor U9867 (N_9867,N_8786,N_9299);
xnor U9868 (N_9868,N_8808,N_8535);
nand U9869 (N_9869,N_6667,N_6344);
nor U9870 (N_9870,N_7014,N_7466);
or U9871 (N_9871,N_6668,N_8737);
nor U9872 (N_9872,N_7474,N_8260);
xnor U9873 (N_9873,N_9114,N_7775);
and U9874 (N_9874,N_8311,N_8929);
or U9875 (N_9875,N_7652,N_9266);
and U9876 (N_9876,N_8374,N_9288);
nor U9877 (N_9877,N_8222,N_7875);
or U9878 (N_9878,N_8587,N_6515);
nand U9879 (N_9879,N_7468,N_8257);
xor U9880 (N_9880,N_6261,N_9271);
and U9881 (N_9881,N_8031,N_8202);
xnor U9882 (N_9882,N_7586,N_7482);
or U9883 (N_9883,N_6502,N_8542);
nand U9884 (N_9884,N_7623,N_7728);
or U9885 (N_9885,N_8676,N_6283);
nand U9886 (N_9886,N_8835,N_6677);
xnor U9887 (N_9887,N_7409,N_7694);
or U9888 (N_9888,N_8698,N_9041);
nor U9889 (N_9889,N_8149,N_7621);
and U9890 (N_9890,N_8603,N_8248);
and U9891 (N_9891,N_8687,N_6776);
xnor U9892 (N_9892,N_6302,N_8391);
and U9893 (N_9893,N_8601,N_6922);
and U9894 (N_9894,N_6967,N_9289);
or U9895 (N_9895,N_7454,N_7749);
xnor U9896 (N_9896,N_8345,N_8071);
and U9897 (N_9897,N_7314,N_6981);
nor U9898 (N_9898,N_7380,N_8540);
xor U9899 (N_9899,N_8803,N_7131);
or U9900 (N_9900,N_6378,N_7703);
or U9901 (N_9901,N_8040,N_9124);
nor U9902 (N_9902,N_8674,N_8881);
and U9903 (N_9903,N_8807,N_9293);
nand U9904 (N_9904,N_7768,N_6627);
or U9905 (N_9905,N_8702,N_7271);
nand U9906 (N_9906,N_7476,N_6897);
xor U9907 (N_9907,N_6448,N_7896);
xor U9908 (N_9908,N_9335,N_8069);
xor U9909 (N_9909,N_7854,N_7989);
and U9910 (N_9910,N_7932,N_9020);
or U9911 (N_9911,N_7401,N_8085);
and U9912 (N_9912,N_8667,N_8343);
xor U9913 (N_9913,N_7773,N_8858);
or U9914 (N_9914,N_8706,N_8735);
nor U9915 (N_9915,N_8478,N_7186);
and U9916 (N_9916,N_6334,N_9210);
and U9917 (N_9917,N_6893,N_6987);
xor U9918 (N_9918,N_9273,N_9356);
or U9919 (N_9919,N_7079,N_7718);
and U9920 (N_9920,N_8878,N_6838);
xor U9921 (N_9921,N_6949,N_8605);
nor U9922 (N_9922,N_8480,N_6370);
nand U9923 (N_9923,N_7785,N_9056);
nand U9924 (N_9924,N_7365,N_8324);
nor U9925 (N_9925,N_8558,N_8196);
or U9926 (N_9926,N_7886,N_7879);
nand U9927 (N_9927,N_7199,N_6355);
nand U9928 (N_9928,N_6265,N_8908);
xnor U9929 (N_9929,N_8728,N_7885);
nand U9930 (N_9930,N_6495,N_8481);
and U9931 (N_9931,N_6376,N_8648);
nand U9932 (N_9932,N_7822,N_7809);
or U9933 (N_9933,N_8747,N_6730);
xor U9934 (N_9934,N_8450,N_7503);
xnor U9935 (N_9935,N_8150,N_7227);
and U9936 (N_9936,N_7844,N_7659);
xnor U9937 (N_9937,N_7540,N_7672);
and U9938 (N_9938,N_9207,N_7553);
nor U9939 (N_9939,N_6449,N_6782);
nor U9940 (N_9940,N_6617,N_6765);
or U9941 (N_9941,N_8639,N_6984);
xnor U9942 (N_9942,N_7336,N_6652);
xnor U9943 (N_9943,N_8143,N_7911);
and U9944 (N_9944,N_8212,N_7733);
and U9945 (N_9945,N_7289,N_6396);
or U9946 (N_9946,N_7023,N_8875);
xnor U9947 (N_9947,N_9125,N_6687);
or U9948 (N_9948,N_8457,N_8852);
or U9949 (N_9949,N_9159,N_6262);
xnor U9950 (N_9950,N_7062,N_8018);
nor U9951 (N_9951,N_7893,N_8813);
nor U9952 (N_9952,N_7319,N_9100);
nand U9953 (N_9953,N_6803,N_8801);
and U9954 (N_9954,N_7389,N_7204);
nand U9955 (N_9955,N_9202,N_7113);
or U9956 (N_9956,N_9086,N_9135);
and U9957 (N_9957,N_6417,N_7601);
nor U9958 (N_9958,N_7555,N_7370);
nand U9959 (N_9959,N_7658,N_7787);
nor U9960 (N_9960,N_7800,N_8146);
nand U9961 (N_9961,N_7545,N_7926);
nor U9962 (N_9962,N_8850,N_9030);
and U9963 (N_9963,N_8657,N_8883);
nor U9964 (N_9964,N_8658,N_8307);
nand U9965 (N_9965,N_7590,N_7029);
xnor U9966 (N_9966,N_6466,N_9038);
and U9967 (N_9967,N_7945,N_9223);
nand U9968 (N_9968,N_7209,N_7083);
and U9969 (N_9969,N_6532,N_7295);
nand U9970 (N_9970,N_7630,N_7219);
xor U9971 (N_9971,N_9245,N_6678);
and U9972 (N_9972,N_8417,N_8338);
nand U9973 (N_9973,N_9258,N_7257);
and U9974 (N_9974,N_8695,N_8551);
nor U9975 (N_9975,N_7596,N_7465);
nand U9976 (N_9976,N_7141,N_8198);
or U9977 (N_9977,N_9248,N_6811);
nand U9978 (N_9978,N_8958,N_8109);
nand U9979 (N_9979,N_6461,N_8802);
nor U9980 (N_9980,N_7245,N_8774);
nor U9981 (N_9981,N_7294,N_7675);
xor U9982 (N_9982,N_7092,N_8434);
and U9983 (N_9983,N_8263,N_7399);
xor U9984 (N_9984,N_9154,N_8500);
nor U9985 (N_9985,N_6923,N_7374);
xnor U9986 (N_9986,N_8344,N_7918);
nand U9987 (N_9987,N_6631,N_9113);
xnor U9988 (N_9988,N_8981,N_9070);
xnor U9989 (N_9989,N_6969,N_8153);
xor U9990 (N_9990,N_7721,N_7754);
or U9991 (N_9991,N_6605,N_7247);
nand U9992 (N_9992,N_6753,N_7858);
nor U9993 (N_9993,N_6380,N_6268);
nand U9994 (N_9994,N_6768,N_8532);
or U9995 (N_9995,N_7969,N_7678);
and U9996 (N_9996,N_7603,N_8486);
nor U9997 (N_9997,N_8339,N_8098);
and U9998 (N_9998,N_9014,N_7827);
and U9999 (N_9999,N_8750,N_6517);
and U10000 (N_10000,N_7508,N_8488);
or U10001 (N_10001,N_8870,N_6911);
nor U10002 (N_10002,N_7354,N_6427);
or U10003 (N_10003,N_8392,N_7272);
xnor U10004 (N_10004,N_8628,N_7148);
and U10005 (N_10005,N_8904,N_9016);
nand U10006 (N_10006,N_7881,N_7892);
xnor U10007 (N_10007,N_6733,N_9208);
or U10008 (N_10008,N_7396,N_8167);
nor U10009 (N_10009,N_7160,N_6597);
or U10010 (N_10010,N_8068,N_6761);
nand U10011 (N_10011,N_7925,N_6826);
nand U10012 (N_10012,N_9196,N_7764);
nand U10013 (N_10013,N_9007,N_6790);
and U10014 (N_10014,N_6497,N_8709);
nor U10015 (N_10015,N_7817,N_7016);
xnor U10016 (N_10016,N_8722,N_7699);
nand U10017 (N_10017,N_8484,N_6322);
nor U10018 (N_10018,N_7490,N_6400);
nor U10019 (N_10019,N_8626,N_7298);
nand U10020 (N_10020,N_8556,N_7951);
xor U10021 (N_10021,N_8916,N_8529);
nand U10022 (N_10022,N_9284,N_8461);
or U10023 (N_10023,N_7547,N_6642);
nand U10024 (N_10024,N_8675,N_9176);
and U10025 (N_10025,N_7597,N_6585);
nor U10026 (N_10026,N_8523,N_8688);
and U10027 (N_10027,N_8966,N_7309);
and U10028 (N_10028,N_6476,N_8834);
and U10029 (N_10029,N_8379,N_7202);
nand U10030 (N_10030,N_9182,N_8182);
xnor U10031 (N_10031,N_7363,N_6664);
nor U10032 (N_10032,N_6759,N_6821);
nand U10033 (N_10033,N_8088,N_6650);
nor U10034 (N_10034,N_8477,N_6382);
or U10035 (N_10035,N_8785,N_7592);
and U10036 (N_10036,N_8740,N_7930);
or U10037 (N_10037,N_6343,N_7662);
nand U10038 (N_10038,N_7318,N_6321);
and U10039 (N_10039,N_6521,N_8612);
xor U10040 (N_10040,N_7583,N_6744);
xor U10041 (N_10041,N_6499,N_6548);
nor U10042 (N_10042,N_8436,N_7937);
nor U10043 (N_10043,N_7929,N_9180);
nor U10044 (N_10044,N_8276,N_7438);
and U10045 (N_10045,N_7433,N_7212);
nor U10046 (N_10046,N_7403,N_8956);
and U10047 (N_10047,N_8429,N_8395);
xnor U10048 (N_10048,N_7191,N_6460);
nor U10049 (N_10049,N_7624,N_6426);
and U10050 (N_10050,N_7797,N_7426);
xor U10051 (N_10051,N_8072,N_6552);
xnor U10052 (N_10052,N_7906,N_7697);
xnor U10053 (N_10053,N_7021,N_6950);
and U10054 (N_10054,N_8654,N_6819);
and U10055 (N_10055,N_7407,N_6368);
nand U10056 (N_10056,N_6480,N_7416);
nand U10057 (N_10057,N_9281,N_6469);
nor U10058 (N_10058,N_6681,N_8115);
nor U10059 (N_10059,N_9066,N_8561);
and U10060 (N_10060,N_7708,N_9122);
nand U10061 (N_10061,N_7549,N_9112);
xor U10062 (N_10062,N_8243,N_8193);
xnor U10063 (N_10063,N_6830,N_8285);
xor U10064 (N_10064,N_8854,N_6329);
or U10065 (N_10065,N_6732,N_9120);
xor U10066 (N_10066,N_8061,N_7157);
nor U10067 (N_10067,N_7506,N_7434);
nor U10068 (N_10068,N_7702,N_8317);
nand U10069 (N_10069,N_9000,N_8036);
and U10070 (N_10070,N_8250,N_7686);
and U10071 (N_10071,N_6920,N_8303);
or U10072 (N_10072,N_8821,N_8943);
and U10073 (N_10073,N_7734,N_6598);
or U10074 (N_10074,N_8502,N_7404);
nand U10075 (N_10075,N_6409,N_7712);
or U10076 (N_10076,N_8081,N_6781);
xor U10077 (N_10077,N_8864,N_8567);
nor U10078 (N_10078,N_8103,N_8856);
nor U10079 (N_10079,N_8938,N_6473);
xnor U10080 (N_10080,N_8015,N_7359);
or U10081 (N_10081,N_6474,N_7627);
nor U10082 (N_10082,N_8410,N_7324);
nor U10083 (N_10083,N_6530,N_8924);
nand U10084 (N_10084,N_8070,N_8060);
or U10085 (N_10085,N_8370,N_9057);
nand U10086 (N_10086,N_8224,N_8828);
xnor U10087 (N_10087,N_9274,N_7328);
nand U10088 (N_10088,N_7949,N_8209);
and U10089 (N_10089,N_6537,N_7027);
nor U10090 (N_10090,N_8188,N_8659);
or U10091 (N_10091,N_9297,N_8548);
nor U10092 (N_10092,N_9272,N_6454);
and U10093 (N_10093,N_6437,N_6278);
xnor U10094 (N_10094,N_6685,N_6784);
nand U10095 (N_10095,N_7074,N_8490);
or U10096 (N_10096,N_9139,N_7248);
and U10097 (N_10097,N_8525,N_8795);
nand U10098 (N_10098,N_7190,N_7692);
or U10099 (N_10099,N_6856,N_9075);
and U10100 (N_10100,N_7075,N_7296);
or U10101 (N_10101,N_7005,N_7236);
nor U10102 (N_10102,N_6943,N_6331);
nor U10103 (N_10103,N_6910,N_8586);
nand U10104 (N_10104,N_7776,N_9179);
nand U10105 (N_10105,N_6944,N_7082);
nor U10106 (N_10106,N_6490,N_7078);
or U10107 (N_10107,N_6452,N_9143);
nor U10108 (N_10108,N_8936,N_7680);
xnor U10109 (N_10109,N_8869,N_6282);
or U10110 (N_10110,N_8433,N_7650);
nand U10111 (N_10111,N_7206,N_6712);
xnor U10112 (N_10112,N_8931,N_7436);
or U10113 (N_10113,N_7484,N_7432);
or U10114 (N_10114,N_8889,N_8289);
and U10115 (N_10115,N_8884,N_7900);
nor U10116 (N_10116,N_7566,N_6618);
nor U10117 (N_10117,N_8631,N_9222);
xnor U10118 (N_10118,N_8726,N_9173);
xnor U10119 (N_10119,N_7923,N_8251);
or U10120 (N_10120,N_9193,N_8868);
nor U10121 (N_10121,N_7442,N_8363);
and U10122 (N_10122,N_9123,N_6961);
nand U10123 (N_10123,N_7821,N_6767);
and U10124 (N_10124,N_6833,N_7047);
or U10125 (N_10125,N_7297,N_9333);
or U10126 (N_10126,N_6806,N_8451);
and U10127 (N_10127,N_7323,N_8730);
xor U10128 (N_10128,N_8843,N_6501);
nor U10129 (N_10129,N_6272,N_8531);
or U10130 (N_10130,N_8141,N_6711);
or U10131 (N_10131,N_9282,N_8155);
and U10132 (N_10132,N_9103,N_7053);
and U10133 (N_10133,N_8946,N_7863);
nor U10134 (N_10134,N_9227,N_6264);
nor U10135 (N_10135,N_8578,N_6815);
xor U10136 (N_10136,N_8333,N_6739);
xnor U10137 (N_10137,N_7862,N_9023);
xor U10138 (N_10138,N_9107,N_7039);
and U10139 (N_10139,N_7395,N_7525);
and U10140 (N_10140,N_7960,N_7963);
and U10141 (N_10141,N_7423,N_8348);
or U10142 (N_10142,N_7522,N_9174);
nand U10143 (N_10143,N_8354,N_7761);
nand U10144 (N_10144,N_6337,N_8380);
and U10145 (N_10145,N_6723,N_6978);
or U10146 (N_10146,N_8598,N_7267);
and U10147 (N_10147,N_7656,N_7599);
or U10148 (N_10148,N_8718,N_7266);
or U10149 (N_10149,N_7333,N_9261);
and U10150 (N_10150,N_6404,N_8930);
nand U10151 (N_10151,N_8849,N_6930);
nand U10152 (N_10152,N_7473,N_8426);
and U10153 (N_10153,N_7560,N_6507);
nand U10154 (N_10154,N_7107,N_6787);
and U10155 (N_10155,N_7833,N_7576);
and U10156 (N_10156,N_6805,N_7170);
and U10157 (N_10157,N_9172,N_8491);
and U10158 (N_10158,N_6875,N_7115);
nor U10159 (N_10159,N_8965,N_8005);
nor U10160 (N_10160,N_7125,N_8533);
nor U10161 (N_10161,N_8408,N_7080);
nor U10162 (N_10162,N_8779,N_8095);
xnor U10163 (N_10163,N_8378,N_7707);
xor U10164 (N_10164,N_7346,N_9105);
or U10165 (N_10165,N_6307,N_9340);
nand U10166 (N_10166,N_7861,N_9206);
nand U10167 (N_10167,N_6619,N_6260);
or U10168 (N_10168,N_8100,N_7460);
or U10169 (N_10169,N_6858,N_8358);
and U10170 (N_10170,N_6390,N_7890);
nor U10171 (N_10171,N_6540,N_8539);
nand U10172 (N_10172,N_8254,N_7530);
or U10173 (N_10173,N_8402,N_8315);
and U10174 (N_10174,N_7282,N_7043);
or U10175 (N_10175,N_8192,N_8321);
nand U10176 (N_10176,N_8221,N_6946);
and U10177 (N_10177,N_7018,N_8123);
and U10178 (N_10178,N_7174,N_6718);
xnor U10179 (N_10179,N_6688,N_7020);
nand U10180 (N_10180,N_9110,N_8704);
nand U10181 (N_10181,N_8589,N_6983);
xor U10182 (N_10182,N_8089,N_8632);
nor U10183 (N_10183,N_7156,N_8006);
and U10184 (N_10184,N_7629,N_7855);
xnor U10185 (N_10185,N_7691,N_9054);
or U10186 (N_10186,N_8482,N_8190);
nor U10187 (N_10187,N_6290,N_8838);
and U10188 (N_10188,N_6926,N_8074);
and U10189 (N_10189,N_7898,N_6879);
nand U10190 (N_10190,N_8851,N_7813);
and U10191 (N_10191,N_8255,N_7081);
nand U10192 (N_10192,N_7172,N_8314);
and U10193 (N_10193,N_7674,N_8199);
xnor U10194 (N_10194,N_7805,N_6612);
or U10195 (N_10195,N_8756,N_7927);
or U10196 (N_10196,N_8888,N_7919);
xnor U10197 (N_10197,N_8609,N_7578);
or U10198 (N_10198,N_9153,N_7520);
or U10199 (N_10199,N_9084,N_8161);
nor U10200 (N_10200,N_8528,N_9012);
xor U10201 (N_10201,N_9026,N_6834);
and U10202 (N_10202,N_8700,N_8717);
xnor U10203 (N_10203,N_6736,N_6500);
or U10204 (N_10204,N_6775,N_8246);
nor U10205 (N_10205,N_8341,N_8863);
nor U10206 (N_10206,N_6896,N_8723);
xor U10207 (N_10207,N_7591,N_9059);
xnor U10208 (N_10208,N_7445,N_9090);
xnor U10209 (N_10209,N_9320,N_7611);
xnor U10210 (N_10210,N_7408,N_7086);
or U10211 (N_10211,N_9060,N_8013);
nor U10212 (N_10212,N_9101,N_7012);
and U10213 (N_10213,N_6938,N_7978);
nor U10214 (N_10214,N_8041,N_6373);
and U10215 (N_10215,N_8267,N_6318);
xnor U10216 (N_10216,N_8600,N_6493);
and U10217 (N_10217,N_7952,N_8220);
nor U10218 (N_10218,N_7139,N_8980);
and U10219 (N_10219,N_8716,N_7103);
and U10220 (N_10220,N_7571,N_9296);
or U10221 (N_10221,N_8876,N_9004);
nand U10222 (N_10222,N_8617,N_6866);
xor U10223 (N_10223,N_8304,N_8877);
or U10224 (N_10224,N_7241,N_7574);
or U10225 (N_10225,N_7993,N_8384);
and U10226 (N_10226,N_8857,N_8159);
nor U10227 (N_10227,N_6898,N_9076);
nand U10228 (N_10228,N_8424,N_8833);
nor U10229 (N_10229,N_6794,N_6483);
xnor U10230 (N_10230,N_8305,N_7104);
and U10231 (N_10231,N_7941,N_8207);
nor U10232 (N_10232,N_8447,N_7538);
nand U10233 (N_10233,N_7831,N_7819);
or U10234 (N_10234,N_6276,N_7069);
nor U10235 (N_10235,N_8331,N_8830);
or U10236 (N_10236,N_8295,N_8166);
nand U10237 (N_10237,N_8028,N_8902);
nor U10238 (N_10238,N_7834,N_6398);
nor U10239 (N_10239,N_9242,N_6259);
xnor U10240 (N_10240,N_8526,N_7367);
nand U10241 (N_10241,N_6581,N_8962);
nand U10242 (N_10242,N_6574,N_8707);
and U10243 (N_10243,N_6397,N_7356);
nand U10244 (N_10244,N_7780,N_7725);
xnor U10245 (N_10245,N_8550,N_8788);
nand U10246 (N_10246,N_6717,N_9167);
nand U10247 (N_10247,N_9355,N_7584);
or U10248 (N_10248,N_8679,N_9071);
xnor U10249 (N_10249,N_8413,N_8078);
nor U10250 (N_10250,N_8634,N_6570);
nand U10251 (N_10251,N_8431,N_8351);
xor U10252 (N_10252,N_9349,N_9039);
nand U10253 (N_10253,N_9240,N_7536);
nor U10254 (N_10254,N_6726,N_6822);
and U10255 (N_10255,N_8281,N_7743);
nor U10256 (N_10256,N_8705,N_8799);
or U10257 (N_10257,N_9329,N_8738);
or U10258 (N_10258,N_6651,N_8213);
or U10259 (N_10259,N_9315,N_8832);
and U10260 (N_10260,N_8912,N_8915);
nor U10261 (N_10261,N_7931,N_7428);
xnor U10262 (N_10262,N_7959,N_7514);
and U10263 (N_10263,N_6870,N_7820);
xnor U10264 (N_10264,N_6412,N_7825);
or U10265 (N_10265,N_8044,N_6287);
nand U10266 (N_10266,N_8057,N_9078);
nand U10267 (N_10267,N_8683,N_7740);
and U10268 (N_10268,N_8108,N_6899);
nand U10269 (N_10269,N_9126,N_7669);
nor U10270 (N_10270,N_8504,N_8435);
and U10271 (N_10271,N_7877,N_8229);
xor U10272 (N_10272,N_6985,N_8183);
and U10273 (N_10273,N_6377,N_9095);
nor U10274 (N_10274,N_7145,N_6735);
and U10275 (N_10275,N_9270,N_6937);
nand U10276 (N_10276,N_7259,N_7207);
nor U10277 (N_10277,N_8781,N_8887);
nor U10278 (N_10278,N_8127,N_7046);
xor U10279 (N_10279,N_7676,N_7330);
or U10280 (N_10280,N_6865,N_8563);
xor U10281 (N_10281,N_6308,N_6751);
or U10282 (N_10282,N_8165,N_8186);
and U10283 (N_10283,N_8404,N_7290);
xnor U10284 (N_10284,N_6653,N_7084);
or U10285 (N_10285,N_7256,N_7261);
nor U10286 (N_10286,N_9231,N_7331);
nor U10287 (N_10287,N_7539,N_8945);
and U10288 (N_10288,N_7117,N_6482);
and U10289 (N_10289,N_9094,N_6724);
nor U10290 (N_10290,N_9169,N_6533);
nor U10291 (N_10291,N_7455,N_6340);
xnor U10292 (N_10292,N_8453,N_7698);
or U10293 (N_10293,N_8771,N_7372);
nor U10294 (N_10294,N_7633,N_7441);
xnor U10295 (N_10295,N_9049,N_8939);
xnor U10296 (N_10296,N_6848,N_6579);
or U10297 (N_10297,N_7616,N_6746);
or U10298 (N_10298,N_8403,N_8579);
nand U10299 (N_10299,N_7128,N_7924);
xor U10300 (N_10300,N_8265,N_7325);
or U10301 (N_10301,N_7869,N_8670);
or U10302 (N_10302,N_8052,N_8990);
or U10303 (N_10303,N_7910,N_6561);
xor U10304 (N_10304,N_8475,N_7093);
and U10305 (N_10305,N_6492,N_8729);
xnor U10306 (N_10306,N_7663,N_8497);
and U10307 (N_10307,N_7249,N_8393);
or U10308 (N_10308,N_6465,N_8918);
nor U10309 (N_10309,N_9317,N_6438);
xor U10310 (N_10310,N_7685,N_6335);
nand U10311 (N_10311,N_6447,N_8093);
xor U10312 (N_10312,N_7198,N_6568);
or U10313 (N_10313,N_7849,N_6756);
and U10314 (N_10314,N_9244,N_8842);
nand U10315 (N_10315,N_6927,N_8982);
and U10316 (N_10316,N_6289,N_9215);
xor U10317 (N_10317,N_6659,N_7173);
nor U10318 (N_10318,N_8681,N_8000);
xor U10319 (N_10319,N_6472,N_9119);
nand U10320 (N_10320,N_9268,N_8636);
nand U10321 (N_10321,N_7954,N_8614);
and U10322 (N_10322,N_6809,N_6769);
and U10323 (N_10323,N_7635,N_8179);
nand U10324 (N_10324,N_9259,N_8680);
nor U10325 (N_10325,N_7976,N_8530);
xnor U10326 (N_10326,N_6364,N_7098);
xnor U10327 (N_10327,N_8460,N_9306);
and U10328 (N_10328,N_9069,N_8003);
nand U10329 (N_10329,N_6908,N_9357);
nand U10330 (N_10330,N_7215,N_7770);
and U10331 (N_10331,N_9156,N_6645);
and U10332 (N_10332,N_7351,N_8439);
nor U10333 (N_10333,N_7619,N_7121);
nor U10334 (N_10334,N_6410,N_6358);
and U10335 (N_10335,N_7845,N_6872);
nor U10336 (N_10336,N_8163,N_7580);
and U10337 (N_10337,N_6372,N_8576);
nor U10338 (N_10338,N_6434,N_9368);
or U10339 (N_10339,N_8332,N_7523);
and U10340 (N_10340,N_6622,N_7938);
and U10341 (N_10341,N_8538,N_6578);
nor U10342 (N_10342,N_7449,N_7238);
or U10343 (N_10343,N_8047,N_6539);
or U10344 (N_10344,N_8432,N_8507);
xnor U10345 (N_10345,N_9336,N_6479);
or U10346 (N_10346,N_7812,N_8002);
and U10347 (N_10347,N_6672,N_8189);
nor U10348 (N_10348,N_7453,N_6549);
xor U10349 (N_10349,N_6951,N_6391);
or U10350 (N_10350,N_7118,N_7814);
xor U10351 (N_10351,N_7510,N_6877);
xnor U10352 (N_10352,N_7059,N_8748);
nor U10353 (N_10353,N_7255,N_8583);
or U10354 (N_10354,N_6513,N_8140);
and U10355 (N_10355,N_8145,N_6255);
xor U10356 (N_10356,N_9037,N_6700);
and U10357 (N_10357,N_9062,N_8663);
nor U10358 (N_10358,N_7035,N_8566);
or U10359 (N_10359,N_8957,N_6760);
or U10360 (N_10360,N_6547,N_7661);
and U10361 (N_10361,N_8396,N_7050);
nand U10362 (N_10362,N_8845,N_6607);
and U10363 (N_10363,N_8650,N_6962);
and U10364 (N_10364,N_8463,N_9181);
and U10365 (N_10365,N_6873,N_7977);
xnor U10366 (N_10366,N_7720,N_8365);
nand U10367 (N_10367,N_8454,N_9157);
nand U10368 (N_10368,N_8329,N_8784);
nand U10369 (N_10369,N_6871,N_8819);
or U10370 (N_10370,N_8947,N_6891);
or U10371 (N_10371,N_8455,N_6414);
and U10372 (N_10372,N_6295,N_8147);
nor U10373 (N_10373,N_6728,N_6657);
and U10374 (N_10374,N_6286,N_8995);
and U10375 (N_10375,N_6941,N_8505);
nor U10376 (N_10376,N_7786,N_6563);
nand U10377 (N_10377,N_9347,N_8390);
or U10378 (N_10378,N_7302,N_7097);
and U10379 (N_10379,N_6862,N_8292);
nor U10380 (N_10380,N_7987,N_8741);
and U10381 (N_10381,N_8899,N_8685);
nor U10382 (N_10382,N_8979,N_7345);
or U10383 (N_10383,N_7968,N_8927);
or U10384 (N_10384,N_7967,N_7903);
nand U10385 (N_10385,N_9200,N_9232);
and U10386 (N_10386,N_7349,N_8211);
nor U10387 (N_10387,N_7983,N_7013);
xnor U10388 (N_10388,N_9142,N_7299);
nor U10389 (N_10389,N_6707,N_8972);
xnor U10390 (N_10390,N_7110,N_8397);
or U10391 (N_10391,N_8170,N_8495);
and U10392 (N_10392,N_7795,N_6399);
nand U10393 (N_10393,N_7509,N_9035);
or U10394 (N_10394,N_9079,N_7504);
nand U10395 (N_10395,N_8038,N_8773);
xnor U10396 (N_10396,N_6625,N_7777);
and U10397 (N_10397,N_9081,N_6939);
nand U10398 (N_10398,N_7136,N_8398);
xnor U10399 (N_10399,N_7485,N_7548);
or U10400 (N_10400,N_7727,N_7573);
or U10401 (N_10401,N_8896,N_8120);
and U10402 (N_10402,N_7251,N_6935);
nor U10403 (N_10403,N_7435,N_7996);
xor U10404 (N_10404,N_7830,N_7515);
nand U10405 (N_10405,N_8151,N_8745);
or U10406 (N_10406,N_8575,N_9148);
nand U10407 (N_10407,N_6800,N_8111);
and U10408 (N_10408,N_6892,N_7524);
nand U10409 (N_10409,N_7179,N_7609);
or U10410 (N_10410,N_6326,N_7868);
nand U10411 (N_10411,N_6572,N_9140);
and U10412 (N_10412,N_8107,N_8953);
nand U10413 (N_10413,N_7481,N_7511);
or U10414 (N_10414,N_9065,N_9226);
nor U10415 (N_10415,N_7837,N_7479);
xnor U10416 (N_10416,N_6375,N_7832);
xor U10417 (N_10417,N_7757,N_8967);
nand U10418 (N_10418,N_7332,N_7724);
nor U10419 (N_10419,N_7980,N_6674);
nor U10420 (N_10420,N_9194,N_8399);
nand U10421 (N_10421,N_7322,N_7745);
nand U10422 (N_10422,N_8653,N_7550);
nand U10423 (N_10423,N_6793,N_6692);
xor U10424 (N_10424,N_6433,N_6786);
or U10425 (N_10425,N_7513,N_8373);
or U10426 (N_10426,N_9373,N_6933);
nor U10427 (N_10427,N_8867,N_9161);
xor U10428 (N_10428,N_6481,N_7642);
nor U10429 (N_10429,N_7956,N_8034);
and U10430 (N_10430,N_8666,N_7748);
nand U10431 (N_10431,N_9040,N_7598);
xor U10432 (N_10432,N_8080,N_8133);
nand U10433 (N_10433,N_9092,N_8512);
and U10434 (N_10434,N_7443,N_6867);
or U10435 (N_10435,N_8950,N_6402);
xor U10436 (N_10436,N_6591,N_7284);
nand U10437 (N_10437,N_8053,N_8994);
or U10438 (N_10438,N_7281,N_7293);
or U10439 (N_10439,N_8110,N_7753);
nand U10440 (N_10440,N_8993,N_9022);
and U10441 (N_10441,N_7638,N_7631);
xor U10442 (N_10442,N_7225,N_7133);
xor U10443 (N_10443,N_6986,N_8010);
and U10444 (N_10444,N_9358,N_7400);
xor U10445 (N_10445,N_7211,N_9138);
nand U10446 (N_10446,N_7011,N_8837);
xnor U10447 (N_10447,N_6429,N_7944);
nand U10448 (N_10448,N_6698,N_6771);
nor U10449 (N_10449,N_8520,N_6970);
nand U10450 (N_10450,N_8534,N_6837);
nor U10451 (N_10451,N_8200,N_8180);
and U10452 (N_10452,N_8234,N_6727);
nand U10453 (N_10453,N_6430,N_8008);
nand U10454 (N_10454,N_7641,N_9219);
or U10455 (N_10455,N_6766,N_8580);
nand U10456 (N_10456,N_8879,N_7250);
or U10457 (N_10457,N_6509,N_7690);
and U10458 (N_10458,N_8797,N_7222);
nand U10459 (N_10459,N_7451,N_9360);
xnor U10460 (N_10460,N_7873,N_9163);
and U10461 (N_10461,N_6791,N_6573);
or U10462 (N_10462,N_6977,N_7682);
or U10463 (N_10463,N_6589,N_6407);
or U10464 (N_10464,N_8909,N_7384);
xnor U10465 (N_10465,N_7887,N_7717);
nor U10466 (N_10466,N_8471,N_8121);
or U10467 (N_10467,N_6254,N_7850);
and U10468 (N_10468,N_6639,N_6270);
or U10469 (N_10469,N_9168,N_7693);
xnor U10470 (N_10470,N_6442,N_6842);
nand U10471 (N_10471,N_7220,N_7593);
nand U10472 (N_10472,N_7527,N_8381);
or U10473 (N_10473,N_6280,N_8299);
xnor U10474 (N_10474,N_6316,N_7472);
xnor U10475 (N_10475,N_8335,N_9235);
xor U10476 (N_10476,N_7140,N_6348);
nand U10477 (N_10477,N_8271,N_6676);
or U10478 (N_10478,N_7286,N_9017);
xnor U10479 (N_10479,N_6505,N_6583);
xor U10480 (N_10480,N_7535,N_7572);
xnor U10481 (N_10481,N_6489,N_6524);
xnor U10482 (N_10482,N_8438,N_8569);
nand U10483 (N_10483,N_6670,N_7406);
xnor U10484 (N_10484,N_7135,N_7914);
and U10485 (N_10485,N_7774,N_8416);
and U10486 (N_10486,N_8096,N_8772);
nor U10487 (N_10487,N_9212,N_7329);
xnor U10488 (N_10488,N_7711,N_6655);
or U10489 (N_10489,N_6996,N_8286);
nand U10490 (N_10490,N_7045,N_8798);
nand U10491 (N_10491,N_7958,N_7908);
nor U10492 (N_10492,N_9025,N_7398);
and U10493 (N_10493,N_7793,N_6351);
nor U10494 (N_10494,N_7493,N_7706);
xor U10495 (N_10495,N_7939,N_8973);
xnor U10496 (N_10496,N_8724,N_7688);
nand U10497 (N_10497,N_7022,N_8721);
and U10498 (N_10498,N_7010,N_9067);
nand U10499 (N_10499,N_6392,N_9363);
xnor U10500 (N_10500,N_7313,N_8252);
nand U10501 (N_10501,N_8130,N_6929);
xor U10502 (N_10502,N_7405,N_7371);
or U10503 (N_10503,N_8318,N_8677);
nor U10504 (N_10504,N_8051,N_8242);
nand U10505 (N_10505,N_8240,N_9093);
or U10506 (N_10506,N_7205,N_8647);
nand U10507 (N_10507,N_9277,N_8405);
nor U10508 (N_10508,N_7004,N_9064);
and U10509 (N_10509,N_8020,N_9061);
nand U10510 (N_10510,N_8114,N_7391);
xor U10511 (N_10511,N_8792,N_8201);
xnor U10512 (N_10512,N_8101,N_8298);
or U10513 (N_10513,N_7056,N_7828);
and U10514 (N_10514,N_8346,N_7364);
xnor U10515 (N_10515,N_7563,N_8572);
nand U10516 (N_10516,N_8824,N_8323);
or U10517 (N_10517,N_6640,N_7640);
nor U10518 (N_10518,N_8823,N_9280);
or U10519 (N_10519,N_9144,N_7444);
nor U10520 (N_10520,N_6901,N_6878);
nor U10521 (N_10521,N_7447,N_8744);
or U10522 (N_10522,N_7475,N_8300);
nor U10523 (N_10523,N_8514,N_6754);
or U10524 (N_10524,N_7183,N_9098);
nor U10525 (N_10525,N_7913,N_6682);
nor U10526 (N_10526,N_6722,N_7264);
xnor U10527 (N_10527,N_9192,N_6538);
and U10528 (N_10528,N_7006,N_9115);
and U10529 (N_10529,N_8742,N_7317);
nor U10530 (N_10530,N_8029,N_6658);
nand U10531 (N_10531,N_6274,N_6535);
nor U10532 (N_10532,N_8932,N_6596);
xor U10533 (N_10533,N_9291,N_9036);
xor U10534 (N_10534,N_7095,N_8594);
nand U10535 (N_10535,N_9343,N_8751);
nand U10536 (N_10536,N_7274,N_9294);
nor U10537 (N_10537,N_6846,N_8686);
or U10538 (N_10538,N_8456,N_9096);
nor U10539 (N_10539,N_6601,N_8951);
or U10540 (N_10540,N_6428,N_7637);
nor U10541 (N_10541,N_6435,N_8306);
nor U10542 (N_10542,N_6855,N_7040);
nor U10543 (N_10543,N_6319,N_7114);
nor U10544 (N_10544,N_8039,N_6808);
and U10545 (N_10545,N_8571,N_7410);
xnor U10546 (N_10546,N_7418,N_7025);
and U10547 (N_10547,N_9300,N_6851);
nand U10548 (N_10548,N_8144,N_6525);
or U10549 (N_10549,N_6541,N_8090);
nor U10550 (N_10550,N_9308,N_7726);
nor U10551 (N_10551,N_6715,N_8049);
nand U10552 (N_10552,N_6649,N_9338);
and U10553 (N_10553,N_8862,N_7065);
nand U10554 (N_10554,N_6595,N_8205);
and U10555 (N_10555,N_7561,N_7089);
nand U10556 (N_10556,N_6836,N_8925);
xor U10557 (N_10557,N_9175,N_6721);
nor U10558 (N_10558,N_7653,N_6785);
xnor U10559 (N_10559,N_9283,N_8249);
nand U10560 (N_10560,N_6555,N_7413);
nand U10561 (N_10561,N_8826,N_8019);
or U10562 (N_10562,N_8616,N_9287);
nor U10563 (N_10563,N_7772,N_7320);
and U10564 (N_10564,N_7741,N_6588);
xor U10565 (N_10565,N_9295,N_6934);
xnor U10566 (N_10566,N_9111,N_8570);
nand U10567 (N_10567,N_9305,N_9089);
or U10568 (N_10568,N_9326,N_6528);
xnor U10569 (N_10569,N_7105,N_7736);
xor U10570 (N_10570,N_6584,N_6418);
and U10571 (N_10571,N_7037,N_6299);
or U10572 (N_10572,N_7750,N_9237);
nand U10573 (N_10573,N_7778,N_8762);
and U10574 (N_10574,N_9021,N_8791);
xor U10575 (N_10575,N_8362,N_7965);
or U10576 (N_10576,N_8746,N_7054);
nor U10577 (N_10577,N_9050,N_9178);
or U10578 (N_10578,N_8844,N_6456);
xor U10579 (N_10579,N_7070,N_9162);
and U10580 (N_10580,N_6883,N_7446);
or U10581 (N_10581,N_7730,N_7342);
nor U10582 (N_10582,N_7860,N_7871);
nand U10583 (N_10583,N_6656,N_8978);
xnor U10584 (N_10584,N_6554,N_7798);
or U10585 (N_10585,N_8033,N_6365);
and U10586 (N_10586,N_8476,N_7802);
and U10587 (N_10587,N_7108,N_7804);
nand U10588 (N_10588,N_6895,N_7614);
xor U10589 (N_10589,N_6695,N_8030);
nand U10590 (N_10590,N_8440,N_7526);
xnor U10591 (N_10591,N_7390,N_8985);
and U10592 (N_10592,N_6810,N_8760);
nor U10593 (N_10593,N_7818,N_9165);
nand U10594 (N_10594,N_6496,N_7487);
nor U10595 (N_10595,N_8673,N_6884);
or U10596 (N_10596,N_6534,N_7159);
or U10597 (N_10597,N_8024,N_9203);
or U10598 (N_10598,N_8394,N_6511);
xor U10599 (N_10599,N_7889,N_7178);
nor U10600 (N_10600,N_7765,N_8816);
nor U10601 (N_10601,N_8593,N_7270);
and U10602 (N_10602,N_8385,N_6510);
nor U10603 (N_10603,N_7529,N_8092);
or U10604 (N_10604,N_6458,N_9027);
or U10605 (N_10605,N_7732,N_8602);
nor U10606 (N_10606,N_7061,N_8176);
and U10607 (N_10607,N_7155,N_6327);
or U10608 (N_10608,N_6354,N_8546);
or U10609 (N_10609,N_6952,N_6464);
xor U10610 (N_10610,N_7905,N_8553);
nor U10611 (N_10611,N_9311,N_8917);
xnor U10612 (N_10612,N_7494,N_9218);
nand U10613 (N_10613,N_6909,N_6804);
and U10614 (N_10614,N_6470,N_8214);
nor U10615 (N_10615,N_7738,N_8025);
xnor U10616 (N_10616,N_7311,N_9328);
and U10617 (N_10617,N_7388,N_6503);
nor U10618 (N_10618,N_7909,N_8983);
xor U10619 (N_10619,N_6369,N_8382);
xnor U10620 (N_10620,N_6620,N_6966);
nor U10621 (N_10621,N_8217,N_9010);
nor U10622 (N_10622,N_7719,N_7387);
and U10623 (N_10623,N_6906,N_9310);
xor U10624 (N_10624,N_7644,N_7464);
or U10625 (N_10625,N_7999,N_6914);
or U10626 (N_10626,N_8914,N_8258);
nand U10627 (N_10627,N_8656,N_9134);
nand U10628 (N_10628,N_8562,N_8627);
xnor U10629 (N_10629,N_8559,N_8637);
nor U10630 (N_10630,N_6519,N_6297);
and U10631 (N_10631,N_8764,N_8984);
xor U10632 (N_10632,N_6689,N_7051);
nor U10633 (N_10633,N_6954,N_6602);
nor U10634 (N_10634,N_6633,N_8767);
or U10635 (N_10635,N_7254,N_7823);
xnor U10636 (N_10636,N_6531,N_9083);
nor U10637 (N_10637,N_7985,N_8091);
nor U10638 (N_10638,N_6742,N_9080);
or U10639 (N_10639,N_7213,N_6948);
nor U10640 (N_10640,N_7166,N_6662);
nor U10641 (N_10641,N_7151,N_8919);
or U10642 (N_10642,N_8590,N_9133);
or U10643 (N_10643,N_6309,N_8645);
or U10644 (N_10644,N_6975,N_7049);
nor U10645 (N_10645,N_7164,N_7605);
and U10646 (N_10646,N_7492,N_6498);
or U10647 (N_10647,N_8903,N_6982);
xnor U10648 (N_10648,N_8066,N_9011);
nor U10649 (N_10649,N_7677,N_7946);
nor U10650 (N_10650,N_8577,N_6342);
and U10651 (N_10651,N_8173,N_7606);
nor U10652 (N_10652,N_7582,N_6360);
xnor U10653 (N_10653,N_9339,N_8743);
nand U10654 (N_10654,N_6457,N_9372);
and U10655 (N_10655,N_8836,N_7439);
xnor U10656 (N_10656,N_7916,N_7142);
nand U10657 (N_10657,N_8999,N_7000);
or U10658 (N_10658,N_8873,N_7991);
and U10659 (N_10659,N_7275,N_8541);
nor U10660 (N_10660,N_6774,N_8839);
xor U10661 (N_10661,N_6359,N_7132);
and U10662 (N_10662,N_9074,N_8933);
xor U10663 (N_10663,N_8283,N_9077);
xor U10664 (N_10664,N_7755,N_8076);
nand U10665 (N_10665,N_8272,N_6773);
xor U10666 (N_10666,N_8664,N_8770);
or U10667 (N_10667,N_6859,N_8794);
nand U10668 (N_10668,N_8624,N_7187);
nand U10669 (N_10669,N_8493,N_6716);
or U10670 (N_10670,N_9352,N_6876);
and U10671 (N_10671,N_7534,N_7060);
nor U10672 (N_10672,N_6825,N_7448);
and U10673 (N_10673,N_8336,N_6864);
nand U10674 (N_10674,N_8629,N_7665);
or U10675 (N_10675,N_9116,N_7228);
nand U10676 (N_10676,N_6611,N_7933);
and U10677 (N_10677,N_8203,N_7567);
nand U10678 (N_10678,N_7670,N_8997);
nand U10679 (N_10679,N_8367,N_8261);
and U10680 (N_10680,N_6955,N_7488);
xor U10681 (N_10681,N_9186,N_8633);
nand U10682 (N_10682,N_8075,N_7815);
or U10683 (N_10683,N_7696,N_8116);
or U10684 (N_10684,N_8181,N_7810);
and U10685 (N_10685,N_7701,N_7258);
nor U10686 (N_10686,N_7169,N_8368);
or U10687 (N_10687,N_6886,N_8905);
nor U10688 (N_10688,N_9348,N_7362);
nor U10689 (N_10689,N_8814,N_6831);
xnor U10690 (N_10690,N_6616,N_8733);
or U10691 (N_10691,N_6425,N_7763);
nand U10692 (N_10692,N_8901,N_9214);
nand U10693 (N_10693,N_7533,N_6976);
or U10694 (N_10694,N_8713,N_6638);
nand U10695 (N_10695,N_9137,N_8174);
nor U10696 (N_10696,N_8644,N_6575);
or U10697 (N_10697,N_7766,N_6381);
and U10698 (N_10698,N_8641,N_8400);
nand U10699 (N_10699,N_7216,N_6816);
nand U10700 (N_10700,N_6703,N_8684);
and U10701 (N_10701,N_8796,N_9344);
or U10702 (N_10702,N_7262,N_7974);
xor U10703 (N_10703,N_6796,N_9051);
nand U10704 (N_10704,N_6965,N_7150);
nor U10705 (N_10705,N_6835,N_8776);
and U10706 (N_10706,N_7177,N_6990);
nor U10707 (N_10707,N_8800,N_7990);
nor U10708 (N_10708,N_8308,N_8506);
xor U10709 (N_10709,N_6251,N_8964);
or U10710 (N_10710,N_7424,N_7936);
nor U10711 (N_10711,N_6440,N_7239);
and U10712 (N_10712,N_8642,N_7912);
or U10713 (N_10713,N_6696,N_8886);
nand U10714 (N_10714,N_6964,N_7126);
xor U10715 (N_10715,N_8223,N_6665);
nand U10716 (N_10716,N_7015,N_7966);
xor U10717 (N_10717,N_9045,N_8350);
xnor U10718 (N_10718,N_6710,N_6374);
nor U10719 (N_10719,N_7781,N_8158);
and U10720 (N_10720,N_7277,N_7361);
and U10721 (N_10721,N_7607,N_8334);
nand U10722 (N_10722,N_7101,N_8152);
nand U10723 (N_10723,N_6680,N_7144);
nand U10724 (N_10724,N_8142,N_6328);
or U10725 (N_10725,N_7681,N_6832);
or U10726 (N_10726,N_7516,N_6904);
xnor U10727 (N_10727,N_7149,N_7841);
nand U10728 (N_10728,N_8340,N_6306);
nand U10729 (N_10729,N_8430,N_7478);
or U10730 (N_10730,N_8245,N_7106);
xor U10731 (N_10731,N_8208,N_7234);
or U10732 (N_10732,N_6277,N_7668);
xor U10733 (N_10733,N_8625,N_7377);
or U10734 (N_10734,N_9298,N_7197);
nor U10735 (N_10735,N_8893,N_6279);
and U10736 (N_10736,N_7986,N_8448);
and U10737 (N_10737,N_8560,N_6518);
nor U10738 (N_10738,N_8231,N_6839);
or U10739 (N_10739,N_8139,N_7501);
nand U10740 (N_10740,N_6757,N_8871);
or U10741 (N_10741,N_9058,N_7803);
xnor U10742 (N_10742,N_7058,N_8262);
nand U10743 (N_10743,N_6362,N_7710);
xor U10744 (N_10744,N_6980,N_6701);
xor U10745 (N_10745,N_8725,N_8259);
nor U10746 (N_10746,N_8848,N_8046);
nor U10747 (N_10747,N_9109,N_6416);
nor U10748 (N_10748,N_7842,N_7235);
or U10749 (N_10749,N_8225,N_7292);
nor U10750 (N_10750,N_9008,N_7654);
and U10751 (N_10751,N_6314,N_7899);
and U10752 (N_10752,N_7378,N_8470);
xor U10753 (N_10753,N_7102,N_6647);
nor U10754 (N_10754,N_7683,N_7796);
and U10755 (N_10755,N_8171,N_7948);
and U10756 (N_10756,N_8353,N_6580);
and U10757 (N_10757,N_7883,N_8496);
or U10758 (N_10758,N_7521,N_7878);
nor U10759 (N_10759,N_8420,N_6636);
nor U10760 (N_10760,N_8521,N_6770);
xnor U10761 (N_10761,N_6894,N_7279);
xor U10762 (N_10762,N_7208,N_8608);
xnor U10763 (N_10763,N_8604,N_8195);
xnor U10764 (N_10764,N_6945,N_8952);
or U10765 (N_10765,N_6363,N_8232);
and U10766 (N_10766,N_9152,N_7657);
and U10767 (N_10767,N_6823,N_7176);
and U10768 (N_10768,N_8230,N_7541);
or U10769 (N_10769,N_7746,N_7366);
or U10770 (N_10770,N_8134,N_6395);
nand U10771 (N_10771,N_9018,N_8055);
and U10772 (N_10772,N_8986,N_6925);
nand U10773 (N_10773,N_9239,N_6298);
and U10774 (N_10774,N_6542,N_7826);
or U10775 (N_10775,N_7648,N_7866);
and U10776 (N_10776,N_7201,N_7194);
or U10777 (N_10777,N_6293,N_7422);
nor U10778 (N_10778,N_6599,N_7090);
or U10779 (N_10779,N_8037,N_7632);
nand U10780 (N_10780,N_8210,N_8014);
or U10781 (N_10781,N_8731,N_8509);
or U10782 (N_10782,N_8418,N_7585);
and U10783 (N_10783,N_8119,N_6523);
xor U10784 (N_10784,N_7788,N_6313);
nor U10785 (N_10785,N_7397,N_7988);
and U10786 (N_10786,N_6556,N_8991);
xor U10787 (N_10787,N_8804,N_6972);
and U10788 (N_10788,N_6551,N_7457);
and U10789 (N_10789,N_8099,N_7617);
nand U10790 (N_10790,N_6330,N_8759);
nor U10791 (N_10791,N_8885,N_8818);
or U10792 (N_10792,N_6840,N_7357);
or U10793 (N_10793,N_7192,N_6683);
and U10794 (N_10794,N_9055,N_8610);
or U10795 (N_10795,N_7838,N_8665);
nand U10796 (N_10796,N_6320,N_6453);
nor U10797 (N_10797,N_8423,N_9187);
xnor U10798 (N_10798,N_7577,N_7376);
xor U10799 (N_10799,N_8638,N_7393);
nand U10800 (N_10800,N_8846,N_6504);
and U10801 (N_10801,N_6571,N_7450);
or U10802 (N_10802,N_8599,N_9002);
nand U10803 (N_10803,N_9236,N_9342);
xnor U10804 (N_10804,N_9367,N_8401);
nand U10805 (N_10805,N_8620,N_8414);
and U10806 (N_10806,N_6747,N_8294);
nor U10807 (N_10807,N_6424,N_6755);
and U10808 (N_10808,N_7542,N_8853);
and U10809 (N_10809,N_8739,N_9228);
xnor U10810 (N_10810,N_7469,N_6797);
or U10811 (N_10811,N_6845,N_6421);
or U10812 (N_10812,N_6560,N_7836);
xnor U10813 (N_10813,N_6557,N_9034);
xor U10814 (N_10814,N_7291,N_8574);
xnor U10815 (N_10815,N_7532,N_6637);
nand U10816 (N_10816,N_7594,N_8054);
and U10817 (N_10817,N_6603,N_6269);
nand U10818 (N_10818,N_8581,N_6992);
or U10819 (N_10819,N_8169,N_7928);
xnor U10820 (N_10820,N_8513,N_6991);
xor U10821 (N_10821,N_6828,N_6455);
nor U10822 (N_10822,N_7790,N_7587);
xnor U10823 (N_10823,N_6288,N_8655);
nor U10824 (N_10824,N_7744,N_8732);
nand U10825 (N_10825,N_6367,N_8244);
and U10826 (N_10826,N_7704,N_9303);
or U10827 (N_10827,N_6463,N_9052);
and U10828 (N_10828,N_7077,N_7901);
or U10829 (N_10829,N_7784,N_6387);
nor U10830 (N_10830,N_9132,N_7824);
and U10831 (N_10831,N_6881,N_6824);
and U10832 (N_10832,N_8316,N_8499);
nand U10833 (N_10833,N_6361,N_8238);
nor U10834 (N_10834,N_8992,N_7181);
or U10835 (N_10835,N_8485,N_9364);
nor U10836 (N_10836,N_6820,N_7218);
xor U10837 (N_10837,N_9118,N_7973);
or U10838 (N_10838,N_8820,N_8462);
nor U10839 (N_10839,N_6576,N_9003);
and U10840 (N_10840,N_7921,N_6613);
nor U10841 (N_10841,N_7268,N_6545);
nand U10842 (N_10842,N_8293,N_7300);
or U10843 (N_10843,N_8611,N_7847);
and U10844 (N_10844,N_7519,N_9073);
xor U10845 (N_10845,N_9304,N_6300);
or U10846 (N_10846,N_8279,N_6420);
and U10847 (N_10847,N_8607,N_6423);
nand U10848 (N_10848,N_7073,N_8596);
and U10849 (N_10849,N_7265,N_9365);
nand U10850 (N_10850,N_6621,N_8544);
nor U10851 (N_10851,N_8714,N_6995);
and U10852 (N_10852,N_8472,N_6332);
xnor U10853 (N_10853,N_7031,N_7518);
or U10854 (N_10854,N_6350,N_7456);
and U10855 (N_10855,N_9249,N_6590);
and U10856 (N_10856,N_8922,N_9229);
or U10857 (N_10857,N_6813,N_6527);
nand U10858 (N_10858,N_9319,N_8469);
xnor U10859 (N_10859,N_8708,N_7537);
or U10860 (N_10860,N_7214,N_7036);
and U10861 (N_10861,N_7269,N_8383);
xnor U10862 (N_10862,N_7288,N_7392);
nand U10863 (N_10863,N_9001,N_7304);
xor U10864 (N_10864,N_8239,N_9044);
or U10865 (N_10865,N_7729,N_9183);
or U10866 (N_10866,N_7556,N_7856);
and U10867 (N_10867,N_8164,N_6459);
nand U10868 (N_10868,N_9309,N_7610);
xor U10869 (N_10869,N_7071,N_8891);
and U10870 (N_10870,N_9370,N_9091);
nand U10871 (N_10871,N_6789,N_8360);
nor U10872 (N_10872,N_9006,N_6777);
and U10873 (N_10873,N_8703,N_8083);
nand U10874 (N_10874,N_9164,N_7622);
and U10875 (N_10875,N_8618,N_8660);
and U10876 (N_10876,N_6702,N_6729);
nand U10877 (N_10877,N_7420,N_7769);
or U10878 (N_10878,N_7502,N_8023);
nand U10879 (N_10879,N_9255,N_7864);
or U10880 (N_10880,N_7415,N_7152);
or U10881 (N_10881,N_9209,N_9099);
xor U10882 (N_10882,N_9246,N_7709);
xnor U10883 (N_10883,N_6772,N_7507);
nand U10884 (N_10884,N_6371,N_9131);
xnor U10885 (N_10885,N_8320,N_9082);
nor U10886 (N_10886,N_9269,N_9128);
nand U10887 (N_10887,N_8043,N_8734);
or U10888 (N_10888,N_8954,N_8117);
or U10889 (N_10889,N_9238,N_6467);
nand U10890 (N_10890,N_9346,N_6586);
or U10891 (N_10891,N_7498,N_7127);
or U10892 (N_10892,N_7122,N_8264);
xor U10893 (N_10893,N_7876,N_7414);
or U10894 (N_10894,N_6349,N_8651);
xor U10895 (N_10895,N_7943,N_7505);
nor U10896 (N_10896,N_6292,N_9224);
xor U10897 (N_10897,N_8126,N_9150);
nor U10898 (N_10898,N_6684,N_7517);
xnor U10899 (N_10899,N_6708,N_8352);
nor U10900 (N_10900,N_8892,N_8421);
xor U10901 (N_10901,N_9267,N_6587);
or U10902 (N_10902,N_9033,N_7315);
nor U10903 (N_10903,N_9322,N_6558);
nor U10904 (N_10904,N_9327,N_7964);
nand U10905 (N_10905,N_9263,N_6432);
nand U10906 (N_10906,N_8710,N_6477);
and U10907 (N_10907,N_6393,N_7001);
nand U10908 (N_10908,N_8105,N_9147);
and U10909 (N_10909,N_9321,N_7167);
xnor U10910 (N_10910,N_7722,N_6353);
or U10911 (N_10911,N_8178,N_7497);
nor U10912 (N_10912,N_8969,N_7301);
nand U10913 (N_10913,N_9068,N_8062);
and U10914 (N_10914,N_6582,N_6646);
xnor U10915 (N_10915,N_8241,N_7041);
nor U10916 (N_10916,N_6624,N_6643);
nand U10917 (N_10917,N_8537,N_7470);
xnor U10918 (N_10918,N_8104,N_7544);
and U10919 (N_10919,N_7947,N_9031);
or U10920 (N_10920,N_9253,N_7894);
nor U10921 (N_10921,N_6623,N_6451);
and U10922 (N_10922,N_8042,N_6610);
nand U10923 (N_10923,N_7119,N_7437);
or U10924 (N_10924,N_7129,N_8357);
and U10925 (N_10925,N_8536,N_7902);
xnor U10926 (N_10926,N_6889,N_6614);
nor U10927 (N_10927,N_6444,N_6737);
nand U10928 (N_10928,N_8125,N_8968);
nor U10929 (N_10929,N_7253,N_6411);
and U10930 (N_10930,N_6660,N_7872);
or U10931 (N_10931,N_7955,N_8711);
or U10932 (N_10932,N_8815,N_9198);
nor U10933 (N_10933,N_8806,N_6792);
xor U10934 (N_10934,N_6900,N_6890);
nor U10935 (N_10935,N_9204,N_7161);
nand U10936 (N_10936,N_9047,N_6669);
or U10937 (N_10937,N_6690,N_8634);
and U10938 (N_10938,N_9318,N_6354);
nand U10939 (N_10939,N_8893,N_8017);
and U10940 (N_10940,N_8122,N_6600);
or U10941 (N_10941,N_8370,N_7957);
nand U10942 (N_10942,N_6315,N_6703);
and U10943 (N_10943,N_7987,N_8330);
nor U10944 (N_10944,N_7651,N_8489);
nand U10945 (N_10945,N_8165,N_7436);
nand U10946 (N_10946,N_7273,N_7240);
and U10947 (N_10947,N_8062,N_9271);
or U10948 (N_10948,N_7673,N_8671);
nor U10949 (N_10949,N_9330,N_8397);
nor U10950 (N_10950,N_6849,N_6465);
and U10951 (N_10951,N_6865,N_9233);
and U10952 (N_10952,N_8128,N_9030);
nor U10953 (N_10953,N_8658,N_7258);
xnor U10954 (N_10954,N_7022,N_8488);
nand U10955 (N_10955,N_6925,N_8238);
xor U10956 (N_10956,N_7047,N_7181);
xnor U10957 (N_10957,N_9339,N_8541);
nand U10958 (N_10958,N_6359,N_8897);
or U10959 (N_10959,N_7810,N_8289);
nor U10960 (N_10960,N_8036,N_8891);
or U10961 (N_10961,N_9026,N_7575);
and U10962 (N_10962,N_7109,N_8735);
nand U10963 (N_10963,N_7078,N_7579);
or U10964 (N_10964,N_6804,N_7391);
nor U10965 (N_10965,N_9327,N_8127);
xnor U10966 (N_10966,N_7684,N_8929);
and U10967 (N_10967,N_6496,N_7436);
nor U10968 (N_10968,N_6686,N_6792);
nor U10969 (N_10969,N_8542,N_7693);
nand U10970 (N_10970,N_8386,N_7518);
nand U10971 (N_10971,N_7637,N_8677);
nand U10972 (N_10972,N_6473,N_7636);
xor U10973 (N_10973,N_7769,N_8993);
and U10974 (N_10974,N_7839,N_8121);
xor U10975 (N_10975,N_7508,N_6762);
nand U10976 (N_10976,N_7420,N_9355);
xor U10977 (N_10977,N_7602,N_7054);
nand U10978 (N_10978,N_8366,N_6401);
nor U10979 (N_10979,N_6578,N_6929);
xnor U10980 (N_10980,N_8758,N_8518);
nor U10981 (N_10981,N_7456,N_8718);
or U10982 (N_10982,N_8145,N_6856);
nand U10983 (N_10983,N_6756,N_7371);
and U10984 (N_10984,N_8183,N_6699);
nand U10985 (N_10985,N_7557,N_8046);
nor U10986 (N_10986,N_9133,N_8686);
or U10987 (N_10987,N_6569,N_6829);
nand U10988 (N_10988,N_7328,N_8588);
nand U10989 (N_10989,N_6899,N_7985);
nand U10990 (N_10990,N_9317,N_8886);
nor U10991 (N_10991,N_7582,N_6302);
or U10992 (N_10992,N_7296,N_8049);
xor U10993 (N_10993,N_8332,N_8633);
nand U10994 (N_10994,N_8415,N_9365);
and U10995 (N_10995,N_8693,N_8914);
or U10996 (N_10996,N_8682,N_7669);
nor U10997 (N_10997,N_9106,N_8247);
or U10998 (N_10998,N_9274,N_9333);
nor U10999 (N_10999,N_7530,N_6745);
nor U11000 (N_11000,N_8903,N_7005);
and U11001 (N_11001,N_7864,N_7172);
or U11002 (N_11002,N_7607,N_7972);
and U11003 (N_11003,N_6579,N_8854);
or U11004 (N_11004,N_8986,N_7857);
nand U11005 (N_11005,N_8849,N_8084);
nor U11006 (N_11006,N_7167,N_8367);
nand U11007 (N_11007,N_8416,N_8005);
and U11008 (N_11008,N_8161,N_6609);
xnor U11009 (N_11009,N_7507,N_6577);
nor U11010 (N_11010,N_7190,N_7277);
nor U11011 (N_11011,N_7328,N_7841);
xor U11012 (N_11012,N_9202,N_7987);
xnor U11013 (N_11013,N_9272,N_7916);
nor U11014 (N_11014,N_7737,N_8217);
and U11015 (N_11015,N_9133,N_6825);
or U11016 (N_11016,N_6663,N_6930);
or U11017 (N_11017,N_6926,N_8029);
nand U11018 (N_11018,N_8103,N_8427);
nand U11019 (N_11019,N_6493,N_7138);
nand U11020 (N_11020,N_9160,N_7697);
nor U11021 (N_11021,N_8936,N_9217);
xnor U11022 (N_11022,N_8878,N_8999);
or U11023 (N_11023,N_6569,N_8079);
nand U11024 (N_11024,N_6773,N_8318);
nand U11025 (N_11025,N_7137,N_8795);
xor U11026 (N_11026,N_9030,N_6497);
nand U11027 (N_11027,N_7370,N_8662);
and U11028 (N_11028,N_7996,N_9108);
or U11029 (N_11029,N_6990,N_8657);
nand U11030 (N_11030,N_9289,N_6724);
nor U11031 (N_11031,N_6763,N_8139);
xor U11032 (N_11032,N_9302,N_8086);
and U11033 (N_11033,N_6906,N_8166);
nand U11034 (N_11034,N_8859,N_6969);
nand U11035 (N_11035,N_9077,N_7851);
nor U11036 (N_11036,N_8507,N_8031);
and U11037 (N_11037,N_7514,N_7391);
nand U11038 (N_11038,N_8725,N_9359);
and U11039 (N_11039,N_8072,N_7791);
or U11040 (N_11040,N_8612,N_9247);
xor U11041 (N_11041,N_6725,N_6799);
nand U11042 (N_11042,N_8581,N_7052);
nand U11043 (N_11043,N_8810,N_7558);
xor U11044 (N_11044,N_7989,N_8444);
and U11045 (N_11045,N_9114,N_8450);
xor U11046 (N_11046,N_7437,N_8989);
and U11047 (N_11047,N_9101,N_6715);
nand U11048 (N_11048,N_8086,N_7893);
nand U11049 (N_11049,N_8046,N_8025);
or U11050 (N_11050,N_8442,N_6994);
nor U11051 (N_11051,N_7832,N_7021);
nor U11052 (N_11052,N_8246,N_8861);
and U11053 (N_11053,N_7290,N_8405);
xnor U11054 (N_11054,N_7225,N_8960);
and U11055 (N_11055,N_8758,N_8024);
xor U11056 (N_11056,N_8810,N_7246);
nand U11057 (N_11057,N_9154,N_7784);
nand U11058 (N_11058,N_8854,N_8364);
nor U11059 (N_11059,N_7043,N_9045);
and U11060 (N_11060,N_9198,N_8046);
nand U11061 (N_11061,N_8934,N_7096);
and U11062 (N_11062,N_7802,N_9216);
or U11063 (N_11063,N_8577,N_7852);
nor U11064 (N_11064,N_7016,N_6284);
xnor U11065 (N_11065,N_8898,N_7147);
or U11066 (N_11066,N_8805,N_9317);
nor U11067 (N_11067,N_9071,N_6431);
and U11068 (N_11068,N_8485,N_6431);
and U11069 (N_11069,N_8414,N_6691);
and U11070 (N_11070,N_8698,N_8915);
or U11071 (N_11071,N_7194,N_6787);
nor U11072 (N_11072,N_7809,N_8421);
and U11073 (N_11073,N_8332,N_8523);
or U11074 (N_11074,N_6820,N_8411);
nor U11075 (N_11075,N_8190,N_7251);
nand U11076 (N_11076,N_7732,N_7834);
and U11077 (N_11077,N_6650,N_6404);
nand U11078 (N_11078,N_8140,N_7378);
nor U11079 (N_11079,N_8227,N_7756);
xnor U11080 (N_11080,N_9045,N_8897);
and U11081 (N_11081,N_6462,N_6349);
or U11082 (N_11082,N_7344,N_7226);
nor U11083 (N_11083,N_6438,N_7660);
or U11084 (N_11084,N_6254,N_7090);
nor U11085 (N_11085,N_7750,N_8885);
nor U11086 (N_11086,N_7319,N_8012);
nand U11087 (N_11087,N_7535,N_8495);
xnor U11088 (N_11088,N_8946,N_9102);
nand U11089 (N_11089,N_8865,N_8741);
or U11090 (N_11090,N_6762,N_8163);
and U11091 (N_11091,N_6812,N_8381);
xor U11092 (N_11092,N_6321,N_9205);
or U11093 (N_11093,N_8364,N_9228);
nor U11094 (N_11094,N_9078,N_6384);
nor U11095 (N_11095,N_8893,N_7250);
and U11096 (N_11096,N_9200,N_6312);
and U11097 (N_11097,N_7306,N_6486);
xnor U11098 (N_11098,N_8438,N_7792);
or U11099 (N_11099,N_7737,N_9136);
nand U11100 (N_11100,N_9032,N_8771);
nor U11101 (N_11101,N_9336,N_7311);
xor U11102 (N_11102,N_7354,N_6361);
nor U11103 (N_11103,N_7797,N_8058);
xnor U11104 (N_11104,N_8968,N_8929);
xnor U11105 (N_11105,N_7059,N_8360);
or U11106 (N_11106,N_8672,N_7078);
nand U11107 (N_11107,N_8453,N_9324);
xnor U11108 (N_11108,N_9158,N_9293);
nor U11109 (N_11109,N_6854,N_7152);
and U11110 (N_11110,N_8526,N_6526);
xor U11111 (N_11111,N_7219,N_9028);
xor U11112 (N_11112,N_6753,N_9351);
and U11113 (N_11113,N_7333,N_6979);
xnor U11114 (N_11114,N_6949,N_6666);
nand U11115 (N_11115,N_7282,N_7099);
nor U11116 (N_11116,N_6812,N_6843);
and U11117 (N_11117,N_7325,N_6517);
and U11118 (N_11118,N_7017,N_6955);
xor U11119 (N_11119,N_7472,N_6597);
nor U11120 (N_11120,N_6786,N_8385);
nor U11121 (N_11121,N_7439,N_6851);
nand U11122 (N_11122,N_6281,N_6962);
and U11123 (N_11123,N_7847,N_8941);
and U11124 (N_11124,N_8651,N_8356);
and U11125 (N_11125,N_6567,N_8940);
or U11126 (N_11126,N_6358,N_7951);
xor U11127 (N_11127,N_9336,N_7569);
nand U11128 (N_11128,N_6608,N_7303);
xor U11129 (N_11129,N_6285,N_7235);
and U11130 (N_11130,N_7481,N_8028);
nor U11131 (N_11131,N_8230,N_9317);
nand U11132 (N_11132,N_8979,N_8070);
nor U11133 (N_11133,N_8731,N_6754);
nand U11134 (N_11134,N_9315,N_9187);
xor U11135 (N_11135,N_7863,N_8226);
or U11136 (N_11136,N_7773,N_8802);
or U11137 (N_11137,N_6987,N_8170);
nor U11138 (N_11138,N_7620,N_7161);
nor U11139 (N_11139,N_6408,N_7205);
xor U11140 (N_11140,N_7110,N_7892);
xor U11141 (N_11141,N_7489,N_8455);
nor U11142 (N_11142,N_7238,N_9054);
xor U11143 (N_11143,N_8139,N_6814);
xnor U11144 (N_11144,N_7590,N_7611);
and U11145 (N_11145,N_7120,N_9014);
nor U11146 (N_11146,N_7913,N_7020);
nand U11147 (N_11147,N_9050,N_8016);
nand U11148 (N_11148,N_8126,N_8799);
and U11149 (N_11149,N_7142,N_8375);
and U11150 (N_11150,N_8450,N_7137);
or U11151 (N_11151,N_6970,N_6817);
and U11152 (N_11152,N_9314,N_9122);
nor U11153 (N_11153,N_7818,N_7301);
nand U11154 (N_11154,N_6785,N_7219);
xor U11155 (N_11155,N_7029,N_9086);
xor U11156 (N_11156,N_8746,N_6552);
nand U11157 (N_11157,N_7556,N_6309);
xor U11158 (N_11158,N_8111,N_8253);
xnor U11159 (N_11159,N_6650,N_9276);
or U11160 (N_11160,N_8751,N_8827);
nand U11161 (N_11161,N_7230,N_7724);
or U11162 (N_11162,N_8905,N_7910);
and U11163 (N_11163,N_9154,N_6501);
nand U11164 (N_11164,N_8766,N_7882);
and U11165 (N_11165,N_8886,N_7988);
or U11166 (N_11166,N_7967,N_6600);
nor U11167 (N_11167,N_8253,N_9226);
xnor U11168 (N_11168,N_6838,N_8367);
nor U11169 (N_11169,N_7989,N_6327);
xor U11170 (N_11170,N_9325,N_9302);
nor U11171 (N_11171,N_8065,N_8424);
nand U11172 (N_11172,N_6320,N_7443);
or U11173 (N_11173,N_7935,N_9035);
or U11174 (N_11174,N_8779,N_6854);
nor U11175 (N_11175,N_8467,N_6785);
nor U11176 (N_11176,N_6298,N_7100);
or U11177 (N_11177,N_9370,N_8310);
nand U11178 (N_11178,N_7301,N_7243);
and U11179 (N_11179,N_6761,N_6441);
nand U11180 (N_11180,N_7907,N_7786);
or U11181 (N_11181,N_7538,N_7569);
and U11182 (N_11182,N_7791,N_8672);
xnor U11183 (N_11183,N_6981,N_6833);
nand U11184 (N_11184,N_6585,N_9185);
nand U11185 (N_11185,N_8617,N_6986);
nor U11186 (N_11186,N_9091,N_6387);
xnor U11187 (N_11187,N_8429,N_8908);
xor U11188 (N_11188,N_6305,N_7771);
nand U11189 (N_11189,N_7770,N_6932);
nand U11190 (N_11190,N_7710,N_6932);
nor U11191 (N_11191,N_8062,N_8298);
or U11192 (N_11192,N_6963,N_7416);
or U11193 (N_11193,N_7235,N_7382);
or U11194 (N_11194,N_8103,N_7741);
or U11195 (N_11195,N_8703,N_7515);
nor U11196 (N_11196,N_8399,N_6905);
and U11197 (N_11197,N_9040,N_9116);
or U11198 (N_11198,N_7621,N_8137);
xnor U11199 (N_11199,N_6795,N_7888);
nor U11200 (N_11200,N_7198,N_9078);
and U11201 (N_11201,N_6655,N_9224);
or U11202 (N_11202,N_6788,N_6611);
and U11203 (N_11203,N_8078,N_8152);
or U11204 (N_11204,N_9210,N_6822);
and U11205 (N_11205,N_7234,N_6665);
nand U11206 (N_11206,N_6269,N_7615);
nor U11207 (N_11207,N_6634,N_9158);
or U11208 (N_11208,N_7779,N_7069);
xor U11209 (N_11209,N_8090,N_9034);
and U11210 (N_11210,N_7217,N_8863);
nor U11211 (N_11211,N_8359,N_7173);
nand U11212 (N_11212,N_7587,N_8201);
and U11213 (N_11213,N_6516,N_6854);
nand U11214 (N_11214,N_7696,N_6990);
and U11215 (N_11215,N_7619,N_8831);
or U11216 (N_11216,N_9367,N_7538);
nand U11217 (N_11217,N_8472,N_6775);
xnor U11218 (N_11218,N_8492,N_8032);
xor U11219 (N_11219,N_7114,N_8909);
xnor U11220 (N_11220,N_6501,N_6743);
xor U11221 (N_11221,N_7051,N_9154);
xor U11222 (N_11222,N_8523,N_8963);
and U11223 (N_11223,N_9131,N_9001);
xor U11224 (N_11224,N_7298,N_8531);
or U11225 (N_11225,N_7766,N_6896);
nand U11226 (N_11226,N_6781,N_6510);
nand U11227 (N_11227,N_7332,N_6609);
and U11228 (N_11228,N_6548,N_7777);
or U11229 (N_11229,N_7741,N_6943);
nand U11230 (N_11230,N_8424,N_6591);
or U11231 (N_11231,N_8539,N_6888);
and U11232 (N_11232,N_8375,N_8590);
xor U11233 (N_11233,N_7817,N_8451);
and U11234 (N_11234,N_6264,N_7599);
nor U11235 (N_11235,N_8413,N_8957);
xor U11236 (N_11236,N_8564,N_8659);
and U11237 (N_11237,N_8764,N_9203);
nand U11238 (N_11238,N_8773,N_8639);
and U11239 (N_11239,N_7470,N_9141);
or U11240 (N_11240,N_6900,N_7660);
or U11241 (N_11241,N_8843,N_6667);
and U11242 (N_11242,N_7043,N_8954);
nor U11243 (N_11243,N_6534,N_7611);
and U11244 (N_11244,N_6928,N_8871);
xor U11245 (N_11245,N_6911,N_7620);
nor U11246 (N_11246,N_8515,N_7792);
and U11247 (N_11247,N_9023,N_9036);
xor U11248 (N_11248,N_7183,N_6908);
nor U11249 (N_11249,N_6363,N_6724);
xor U11250 (N_11250,N_9225,N_6710);
nand U11251 (N_11251,N_7638,N_8559);
nand U11252 (N_11252,N_7161,N_7936);
and U11253 (N_11253,N_6729,N_8073);
nor U11254 (N_11254,N_8917,N_6642);
xnor U11255 (N_11255,N_7734,N_9312);
and U11256 (N_11256,N_7383,N_7597);
nor U11257 (N_11257,N_6841,N_6335);
xor U11258 (N_11258,N_8406,N_7256);
nor U11259 (N_11259,N_7852,N_8916);
xor U11260 (N_11260,N_6968,N_7959);
xor U11261 (N_11261,N_7646,N_6338);
and U11262 (N_11262,N_7008,N_7081);
or U11263 (N_11263,N_9252,N_8553);
nand U11264 (N_11264,N_8405,N_7718);
or U11265 (N_11265,N_7524,N_9350);
or U11266 (N_11266,N_7288,N_7581);
nand U11267 (N_11267,N_6386,N_7116);
xor U11268 (N_11268,N_6594,N_6932);
xnor U11269 (N_11269,N_9275,N_8356);
nand U11270 (N_11270,N_7039,N_7718);
and U11271 (N_11271,N_8534,N_8005);
nor U11272 (N_11272,N_6722,N_6276);
or U11273 (N_11273,N_9189,N_7484);
and U11274 (N_11274,N_8810,N_6949);
or U11275 (N_11275,N_8502,N_8169);
or U11276 (N_11276,N_8884,N_8054);
nand U11277 (N_11277,N_6477,N_7483);
xor U11278 (N_11278,N_7184,N_7611);
xnor U11279 (N_11279,N_6390,N_8545);
and U11280 (N_11280,N_6320,N_6606);
xor U11281 (N_11281,N_8374,N_8419);
or U11282 (N_11282,N_7462,N_6793);
nor U11283 (N_11283,N_7275,N_6648);
xnor U11284 (N_11284,N_8959,N_8732);
nand U11285 (N_11285,N_6979,N_7403);
nor U11286 (N_11286,N_6287,N_7755);
nor U11287 (N_11287,N_9282,N_6753);
nand U11288 (N_11288,N_8547,N_8499);
nand U11289 (N_11289,N_9272,N_6456);
or U11290 (N_11290,N_7508,N_8437);
nand U11291 (N_11291,N_8945,N_9225);
or U11292 (N_11292,N_8942,N_7211);
and U11293 (N_11293,N_7136,N_8575);
or U11294 (N_11294,N_7116,N_7997);
nor U11295 (N_11295,N_7125,N_8696);
xnor U11296 (N_11296,N_8740,N_7601);
or U11297 (N_11297,N_8781,N_7370);
nor U11298 (N_11298,N_8711,N_7611);
or U11299 (N_11299,N_7192,N_7368);
xor U11300 (N_11300,N_8044,N_7316);
and U11301 (N_11301,N_7694,N_8355);
or U11302 (N_11302,N_6804,N_8942);
or U11303 (N_11303,N_7869,N_8296);
or U11304 (N_11304,N_8430,N_7296);
nor U11305 (N_11305,N_9108,N_6782);
and U11306 (N_11306,N_8758,N_8366);
nand U11307 (N_11307,N_7279,N_9051);
xor U11308 (N_11308,N_7733,N_6421);
nand U11309 (N_11309,N_8542,N_7604);
nor U11310 (N_11310,N_7074,N_7640);
and U11311 (N_11311,N_9096,N_8461);
nand U11312 (N_11312,N_6953,N_6994);
xnor U11313 (N_11313,N_8985,N_8874);
or U11314 (N_11314,N_6387,N_6980);
nor U11315 (N_11315,N_7275,N_7541);
and U11316 (N_11316,N_6493,N_7752);
nand U11317 (N_11317,N_7037,N_6510);
xnor U11318 (N_11318,N_7849,N_7394);
or U11319 (N_11319,N_6668,N_6906);
nand U11320 (N_11320,N_7890,N_8777);
and U11321 (N_11321,N_7998,N_8854);
or U11322 (N_11322,N_6345,N_9309);
or U11323 (N_11323,N_7113,N_8607);
or U11324 (N_11324,N_8113,N_6480);
nor U11325 (N_11325,N_6849,N_8424);
nand U11326 (N_11326,N_8164,N_8435);
nand U11327 (N_11327,N_6667,N_6871);
nor U11328 (N_11328,N_8477,N_8645);
nor U11329 (N_11329,N_6792,N_7757);
nor U11330 (N_11330,N_7236,N_6599);
xnor U11331 (N_11331,N_8050,N_9049);
and U11332 (N_11332,N_7499,N_7457);
nor U11333 (N_11333,N_7488,N_8747);
xnor U11334 (N_11334,N_8031,N_7191);
nor U11335 (N_11335,N_6747,N_9327);
nand U11336 (N_11336,N_7973,N_6417);
nor U11337 (N_11337,N_7945,N_6861);
and U11338 (N_11338,N_8101,N_8370);
nand U11339 (N_11339,N_7010,N_7160);
or U11340 (N_11340,N_6919,N_6432);
and U11341 (N_11341,N_9165,N_7571);
and U11342 (N_11342,N_7464,N_8303);
xnor U11343 (N_11343,N_6969,N_7526);
or U11344 (N_11344,N_7831,N_6674);
nand U11345 (N_11345,N_8398,N_8778);
and U11346 (N_11346,N_8354,N_6730);
and U11347 (N_11347,N_7603,N_6911);
and U11348 (N_11348,N_6370,N_6412);
nand U11349 (N_11349,N_9020,N_6667);
xor U11350 (N_11350,N_9332,N_6436);
nand U11351 (N_11351,N_8795,N_8113);
or U11352 (N_11352,N_8823,N_7640);
or U11353 (N_11353,N_7532,N_8445);
and U11354 (N_11354,N_6324,N_6819);
and U11355 (N_11355,N_7633,N_7065);
nor U11356 (N_11356,N_6989,N_6471);
nand U11357 (N_11357,N_7521,N_8499);
xnor U11358 (N_11358,N_7942,N_8835);
nor U11359 (N_11359,N_7364,N_8177);
nand U11360 (N_11360,N_6618,N_6665);
nor U11361 (N_11361,N_9352,N_8155);
xnor U11362 (N_11362,N_7586,N_9183);
or U11363 (N_11363,N_8090,N_7051);
xnor U11364 (N_11364,N_6967,N_7982);
xor U11365 (N_11365,N_7089,N_7587);
xnor U11366 (N_11366,N_8648,N_7390);
nand U11367 (N_11367,N_7160,N_8699);
xor U11368 (N_11368,N_9216,N_7480);
nand U11369 (N_11369,N_8012,N_6425);
or U11370 (N_11370,N_7392,N_8788);
nand U11371 (N_11371,N_7272,N_6263);
and U11372 (N_11372,N_8539,N_7942);
nor U11373 (N_11373,N_7507,N_6538);
or U11374 (N_11374,N_7746,N_6375);
nor U11375 (N_11375,N_8829,N_7568);
or U11376 (N_11376,N_7312,N_7302);
xnor U11377 (N_11377,N_8987,N_7939);
nor U11378 (N_11378,N_8728,N_8694);
xor U11379 (N_11379,N_9214,N_9374);
or U11380 (N_11380,N_7911,N_6688);
nor U11381 (N_11381,N_6674,N_9128);
and U11382 (N_11382,N_6925,N_7798);
or U11383 (N_11383,N_9097,N_7705);
nor U11384 (N_11384,N_6631,N_6765);
or U11385 (N_11385,N_7931,N_6370);
xor U11386 (N_11386,N_7045,N_7528);
xor U11387 (N_11387,N_8769,N_9270);
nor U11388 (N_11388,N_6492,N_8292);
and U11389 (N_11389,N_7204,N_7487);
xor U11390 (N_11390,N_6675,N_9115);
xnor U11391 (N_11391,N_6368,N_6329);
xnor U11392 (N_11392,N_9106,N_8569);
and U11393 (N_11393,N_7764,N_6758);
nor U11394 (N_11394,N_7688,N_6827);
and U11395 (N_11395,N_7595,N_7573);
and U11396 (N_11396,N_7994,N_8558);
or U11397 (N_11397,N_8550,N_7535);
nor U11398 (N_11398,N_6839,N_7921);
or U11399 (N_11399,N_8498,N_6417);
xor U11400 (N_11400,N_7889,N_8274);
and U11401 (N_11401,N_9321,N_6313);
xnor U11402 (N_11402,N_6527,N_7248);
nand U11403 (N_11403,N_8977,N_7970);
nand U11404 (N_11404,N_7493,N_8203);
or U11405 (N_11405,N_9228,N_8422);
xor U11406 (N_11406,N_6697,N_8329);
nor U11407 (N_11407,N_8064,N_7171);
xnor U11408 (N_11408,N_8371,N_7393);
xor U11409 (N_11409,N_9088,N_9344);
or U11410 (N_11410,N_7260,N_7860);
nand U11411 (N_11411,N_8930,N_8320);
or U11412 (N_11412,N_7324,N_8335);
or U11413 (N_11413,N_7717,N_6607);
nand U11414 (N_11414,N_8036,N_7392);
nand U11415 (N_11415,N_6787,N_8900);
xnor U11416 (N_11416,N_7089,N_8592);
nor U11417 (N_11417,N_7483,N_7472);
nor U11418 (N_11418,N_8951,N_7704);
nor U11419 (N_11419,N_8407,N_8708);
or U11420 (N_11420,N_7563,N_7140);
xor U11421 (N_11421,N_7087,N_7888);
nor U11422 (N_11422,N_7573,N_9015);
and U11423 (N_11423,N_7265,N_6822);
xnor U11424 (N_11424,N_6583,N_7736);
and U11425 (N_11425,N_7185,N_7323);
or U11426 (N_11426,N_6264,N_9335);
xor U11427 (N_11427,N_8538,N_8996);
xor U11428 (N_11428,N_7295,N_6875);
and U11429 (N_11429,N_8849,N_7386);
nor U11430 (N_11430,N_8023,N_6381);
nor U11431 (N_11431,N_6485,N_7753);
or U11432 (N_11432,N_8173,N_7744);
or U11433 (N_11433,N_8264,N_6340);
nand U11434 (N_11434,N_8780,N_7758);
or U11435 (N_11435,N_6807,N_7066);
or U11436 (N_11436,N_8414,N_7899);
xor U11437 (N_11437,N_9060,N_6608);
or U11438 (N_11438,N_6826,N_8676);
or U11439 (N_11439,N_6767,N_8922);
nor U11440 (N_11440,N_8174,N_7794);
xor U11441 (N_11441,N_9082,N_6380);
and U11442 (N_11442,N_7255,N_6946);
nor U11443 (N_11443,N_6334,N_6552);
or U11444 (N_11444,N_7636,N_6501);
and U11445 (N_11445,N_8880,N_7801);
and U11446 (N_11446,N_6536,N_8215);
nand U11447 (N_11447,N_9077,N_8705);
xnor U11448 (N_11448,N_8157,N_6604);
and U11449 (N_11449,N_8267,N_7613);
nor U11450 (N_11450,N_8165,N_9170);
and U11451 (N_11451,N_7945,N_7089);
xnor U11452 (N_11452,N_7708,N_6610);
and U11453 (N_11453,N_7947,N_7261);
xnor U11454 (N_11454,N_7272,N_8665);
or U11455 (N_11455,N_6711,N_7830);
nand U11456 (N_11456,N_6592,N_6253);
or U11457 (N_11457,N_9047,N_7217);
or U11458 (N_11458,N_8981,N_6652);
xor U11459 (N_11459,N_9102,N_9030);
and U11460 (N_11460,N_6339,N_7749);
nor U11461 (N_11461,N_7827,N_8488);
or U11462 (N_11462,N_7839,N_6271);
and U11463 (N_11463,N_8457,N_8461);
or U11464 (N_11464,N_8334,N_8756);
and U11465 (N_11465,N_7889,N_7616);
and U11466 (N_11466,N_8938,N_9079);
nand U11467 (N_11467,N_6557,N_9015);
nor U11468 (N_11468,N_7528,N_6450);
xnor U11469 (N_11469,N_7440,N_7922);
and U11470 (N_11470,N_6985,N_7304);
xnor U11471 (N_11471,N_6679,N_7242);
nor U11472 (N_11472,N_8930,N_9102);
nand U11473 (N_11473,N_9081,N_6328);
and U11474 (N_11474,N_9111,N_7957);
nand U11475 (N_11475,N_6342,N_7333);
and U11476 (N_11476,N_9179,N_9030);
xnor U11477 (N_11477,N_7223,N_9285);
and U11478 (N_11478,N_6545,N_8136);
or U11479 (N_11479,N_7537,N_8933);
xor U11480 (N_11480,N_7383,N_7192);
nand U11481 (N_11481,N_8602,N_6938);
xor U11482 (N_11482,N_8159,N_6554);
and U11483 (N_11483,N_9077,N_9192);
nand U11484 (N_11484,N_8227,N_6544);
nand U11485 (N_11485,N_6988,N_7499);
nand U11486 (N_11486,N_8577,N_6861);
xnor U11487 (N_11487,N_8969,N_7695);
or U11488 (N_11488,N_8528,N_8939);
nor U11489 (N_11489,N_7537,N_8031);
xnor U11490 (N_11490,N_8569,N_7176);
nand U11491 (N_11491,N_9011,N_7972);
and U11492 (N_11492,N_8125,N_7091);
and U11493 (N_11493,N_9112,N_9222);
nor U11494 (N_11494,N_6353,N_6848);
nor U11495 (N_11495,N_8596,N_8090);
and U11496 (N_11496,N_7798,N_8721);
or U11497 (N_11497,N_8311,N_8843);
nor U11498 (N_11498,N_9146,N_7356);
nor U11499 (N_11499,N_8027,N_6989);
or U11500 (N_11500,N_6701,N_9304);
nand U11501 (N_11501,N_6376,N_8484);
and U11502 (N_11502,N_9101,N_7962);
and U11503 (N_11503,N_9135,N_8713);
and U11504 (N_11504,N_9046,N_6888);
and U11505 (N_11505,N_6730,N_8292);
and U11506 (N_11506,N_7311,N_6698);
nand U11507 (N_11507,N_6282,N_7816);
xor U11508 (N_11508,N_7007,N_7544);
and U11509 (N_11509,N_9060,N_8758);
and U11510 (N_11510,N_9340,N_8180);
or U11511 (N_11511,N_8884,N_7463);
xor U11512 (N_11512,N_8483,N_8230);
nand U11513 (N_11513,N_6830,N_8367);
and U11514 (N_11514,N_6741,N_9189);
nand U11515 (N_11515,N_6557,N_6611);
nor U11516 (N_11516,N_7413,N_7177);
or U11517 (N_11517,N_8463,N_7755);
nand U11518 (N_11518,N_6462,N_7866);
or U11519 (N_11519,N_7098,N_8377);
nor U11520 (N_11520,N_6876,N_8425);
or U11521 (N_11521,N_7537,N_7489);
xnor U11522 (N_11522,N_9152,N_8565);
xnor U11523 (N_11523,N_7652,N_6808);
or U11524 (N_11524,N_7312,N_8642);
and U11525 (N_11525,N_9115,N_7119);
xnor U11526 (N_11526,N_6646,N_8853);
and U11527 (N_11527,N_6984,N_7318);
nand U11528 (N_11528,N_7799,N_8095);
xor U11529 (N_11529,N_7773,N_6307);
or U11530 (N_11530,N_8355,N_7661);
or U11531 (N_11531,N_8076,N_7283);
nand U11532 (N_11532,N_8059,N_9336);
and U11533 (N_11533,N_8887,N_9294);
nor U11534 (N_11534,N_7333,N_8256);
nand U11535 (N_11535,N_8648,N_6529);
and U11536 (N_11536,N_8324,N_7628);
or U11537 (N_11537,N_8540,N_8287);
or U11538 (N_11538,N_8091,N_7684);
nor U11539 (N_11539,N_7144,N_7468);
nand U11540 (N_11540,N_6459,N_7547);
or U11541 (N_11541,N_6892,N_8516);
nor U11542 (N_11542,N_8910,N_8473);
nand U11543 (N_11543,N_6599,N_8329);
xnor U11544 (N_11544,N_7590,N_6301);
nor U11545 (N_11545,N_7666,N_7022);
or U11546 (N_11546,N_9256,N_8873);
or U11547 (N_11547,N_8765,N_8386);
and U11548 (N_11548,N_8823,N_9040);
and U11549 (N_11549,N_8381,N_7480);
nor U11550 (N_11550,N_7286,N_7545);
xor U11551 (N_11551,N_8155,N_7727);
nor U11552 (N_11552,N_7117,N_6578);
and U11553 (N_11553,N_6790,N_7481);
nor U11554 (N_11554,N_7157,N_7230);
or U11555 (N_11555,N_8388,N_7283);
and U11556 (N_11556,N_6669,N_6763);
nor U11557 (N_11557,N_7895,N_8109);
nor U11558 (N_11558,N_7282,N_8224);
or U11559 (N_11559,N_9280,N_6372);
or U11560 (N_11560,N_7796,N_7914);
xor U11561 (N_11561,N_8114,N_7339);
nand U11562 (N_11562,N_8156,N_9049);
and U11563 (N_11563,N_8885,N_7642);
nand U11564 (N_11564,N_8633,N_8571);
nand U11565 (N_11565,N_8229,N_9141);
nor U11566 (N_11566,N_8530,N_8966);
and U11567 (N_11567,N_7496,N_7796);
nand U11568 (N_11568,N_6793,N_7974);
xor U11569 (N_11569,N_8405,N_7604);
xnor U11570 (N_11570,N_8131,N_8741);
and U11571 (N_11571,N_6947,N_8955);
and U11572 (N_11572,N_8874,N_8590);
nand U11573 (N_11573,N_8772,N_7719);
xnor U11574 (N_11574,N_7501,N_8845);
and U11575 (N_11575,N_6832,N_6720);
and U11576 (N_11576,N_9231,N_8455);
or U11577 (N_11577,N_8963,N_7422);
xor U11578 (N_11578,N_7035,N_8601);
or U11579 (N_11579,N_7197,N_7255);
xor U11580 (N_11580,N_8663,N_8641);
nor U11581 (N_11581,N_9193,N_6287);
or U11582 (N_11582,N_7212,N_7069);
nor U11583 (N_11583,N_8092,N_7701);
xnor U11584 (N_11584,N_6754,N_7069);
nor U11585 (N_11585,N_8551,N_7115);
or U11586 (N_11586,N_7738,N_7323);
or U11587 (N_11587,N_7588,N_8222);
and U11588 (N_11588,N_7725,N_6455);
xnor U11589 (N_11589,N_6263,N_9184);
nor U11590 (N_11590,N_8691,N_7078);
xnor U11591 (N_11591,N_9172,N_7260);
nand U11592 (N_11592,N_6987,N_9338);
nand U11593 (N_11593,N_6699,N_7710);
and U11594 (N_11594,N_6904,N_8240);
or U11595 (N_11595,N_9052,N_7583);
nor U11596 (N_11596,N_6728,N_9260);
xnor U11597 (N_11597,N_8286,N_6366);
or U11598 (N_11598,N_7324,N_7978);
xor U11599 (N_11599,N_8346,N_7715);
nor U11600 (N_11600,N_7667,N_8854);
nand U11601 (N_11601,N_6285,N_8449);
nor U11602 (N_11602,N_6384,N_8195);
nor U11603 (N_11603,N_9107,N_7726);
nand U11604 (N_11604,N_7781,N_8560);
xnor U11605 (N_11605,N_7186,N_8651);
or U11606 (N_11606,N_7233,N_8633);
nor U11607 (N_11607,N_7780,N_8781);
nor U11608 (N_11608,N_6626,N_7032);
nand U11609 (N_11609,N_8443,N_6310);
or U11610 (N_11610,N_7404,N_8394);
and U11611 (N_11611,N_6457,N_7163);
or U11612 (N_11612,N_9259,N_8587);
and U11613 (N_11613,N_8772,N_7472);
nand U11614 (N_11614,N_8655,N_8323);
or U11615 (N_11615,N_8008,N_7904);
xor U11616 (N_11616,N_8153,N_6570);
nor U11617 (N_11617,N_7307,N_7837);
or U11618 (N_11618,N_9204,N_9066);
nor U11619 (N_11619,N_8236,N_7685);
nand U11620 (N_11620,N_6785,N_7423);
nand U11621 (N_11621,N_7703,N_8244);
nor U11622 (N_11622,N_7979,N_8438);
nor U11623 (N_11623,N_6950,N_8446);
and U11624 (N_11624,N_6826,N_6815);
xnor U11625 (N_11625,N_6664,N_7488);
and U11626 (N_11626,N_8376,N_8194);
nand U11627 (N_11627,N_6707,N_7784);
and U11628 (N_11628,N_7636,N_6848);
nor U11629 (N_11629,N_8672,N_9155);
nand U11630 (N_11630,N_6738,N_7789);
nor U11631 (N_11631,N_8348,N_7879);
and U11632 (N_11632,N_8713,N_7675);
nand U11633 (N_11633,N_6481,N_7854);
or U11634 (N_11634,N_7507,N_7920);
nand U11635 (N_11635,N_6549,N_6772);
xor U11636 (N_11636,N_8275,N_7058);
and U11637 (N_11637,N_9229,N_8291);
xor U11638 (N_11638,N_6791,N_9139);
nor U11639 (N_11639,N_9349,N_8498);
nor U11640 (N_11640,N_7635,N_7184);
nand U11641 (N_11641,N_8305,N_8044);
nand U11642 (N_11642,N_7137,N_7925);
xnor U11643 (N_11643,N_8794,N_8134);
and U11644 (N_11644,N_8338,N_7247);
and U11645 (N_11645,N_6743,N_8370);
or U11646 (N_11646,N_8936,N_9286);
nor U11647 (N_11647,N_8092,N_9291);
nor U11648 (N_11648,N_8467,N_9077);
nor U11649 (N_11649,N_6422,N_9335);
xor U11650 (N_11650,N_6984,N_8439);
and U11651 (N_11651,N_8580,N_7340);
xor U11652 (N_11652,N_8552,N_7122);
xnor U11653 (N_11653,N_6603,N_8211);
xnor U11654 (N_11654,N_8197,N_7702);
nand U11655 (N_11655,N_8779,N_7811);
nand U11656 (N_11656,N_8439,N_7944);
nand U11657 (N_11657,N_8441,N_8966);
or U11658 (N_11658,N_6668,N_6749);
nand U11659 (N_11659,N_8399,N_8319);
or U11660 (N_11660,N_6694,N_7912);
nor U11661 (N_11661,N_7141,N_8846);
nand U11662 (N_11662,N_6661,N_8735);
or U11663 (N_11663,N_7237,N_6705);
xnor U11664 (N_11664,N_6886,N_6448);
nor U11665 (N_11665,N_8299,N_6741);
and U11666 (N_11666,N_7072,N_6745);
and U11667 (N_11667,N_7768,N_6796);
xnor U11668 (N_11668,N_7117,N_6841);
nor U11669 (N_11669,N_7725,N_7578);
xor U11670 (N_11670,N_7833,N_7715);
nand U11671 (N_11671,N_6645,N_6561);
nor U11672 (N_11672,N_7937,N_7047);
and U11673 (N_11673,N_6503,N_7668);
nor U11674 (N_11674,N_8144,N_6474);
or U11675 (N_11675,N_7771,N_8464);
or U11676 (N_11676,N_6522,N_6555);
xnor U11677 (N_11677,N_8685,N_7585);
nor U11678 (N_11678,N_7397,N_9093);
xnor U11679 (N_11679,N_6599,N_9097);
nand U11680 (N_11680,N_7445,N_7410);
and U11681 (N_11681,N_8396,N_6623);
or U11682 (N_11682,N_8059,N_8693);
xnor U11683 (N_11683,N_8037,N_7016);
or U11684 (N_11684,N_6837,N_7494);
nor U11685 (N_11685,N_8806,N_8134);
nor U11686 (N_11686,N_8613,N_8427);
nor U11687 (N_11687,N_8260,N_7444);
nand U11688 (N_11688,N_7246,N_7501);
or U11689 (N_11689,N_6427,N_7177);
and U11690 (N_11690,N_7660,N_8905);
nor U11691 (N_11691,N_8934,N_8027);
nor U11692 (N_11692,N_9027,N_6773);
nor U11693 (N_11693,N_8448,N_9251);
nand U11694 (N_11694,N_7009,N_8302);
nand U11695 (N_11695,N_7205,N_8929);
or U11696 (N_11696,N_7141,N_8491);
nand U11697 (N_11697,N_8049,N_6944);
and U11698 (N_11698,N_8860,N_8106);
nor U11699 (N_11699,N_9100,N_7057);
xor U11700 (N_11700,N_7532,N_6384);
nand U11701 (N_11701,N_7003,N_6895);
xnor U11702 (N_11702,N_6480,N_8853);
nand U11703 (N_11703,N_9128,N_8068);
nor U11704 (N_11704,N_8138,N_9152);
xnor U11705 (N_11705,N_7826,N_8309);
xor U11706 (N_11706,N_6911,N_8527);
nand U11707 (N_11707,N_7748,N_7671);
nand U11708 (N_11708,N_7084,N_8295);
nand U11709 (N_11709,N_8650,N_9188);
or U11710 (N_11710,N_7582,N_8488);
and U11711 (N_11711,N_8651,N_8894);
xnor U11712 (N_11712,N_7409,N_8463);
and U11713 (N_11713,N_8503,N_6672);
xnor U11714 (N_11714,N_8894,N_7468);
nand U11715 (N_11715,N_7728,N_7838);
nor U11716 (N_11716,N_8564,N_8286);
or U11717 (N_11717,N_7456,N_8598);
nor U11718 (N_11718,N_6432,N_8829);
or U11719 (N_11719,N_7707,N_9291);
and U11720 (N_11720,N_7803,N_6949);
nand U11721 (N_11721,N_7241,N_7002);
nand U11722 (N_11722,N_6610,N_8670);
nand U11723 (N_11723,N_7491,N_7483);
nand U11724 (N_11724,N_6276,N_8963);
or U11725 (N_11725,N_7883,N_9218);
and U11726 (N_11726,N_8015,N_6644);
nand U11727 (N_11727,N_8341,N_7075);
and U11728 (N_11728,N_8924,N_9106);
nor U11729 (N_11729,N_8045,N_6995);
and U11730 (N_11730,N_6483,N_6606);
and U11731 (N_11731,N_7940,N_8141);
xor U11732 (N_11732,N_8255,N_7840);
and U11733 (N_11733,N_8631,N_7204);
xor U11734 (N_11734,N_6907,N_7016);
and U11735 (N_11735,N_7314,N_6635);
xor U11736 (N_11736,N_7586,N_7877);
nand U11737 (N_11737,N_6263,N_9216);
and U11738 (N_11738,N_8451,N_6616);
or U11739 (N_11739,N_7115,N_7722);
nor U11740 (N_11740,N_8598,N_6987);
or U11741 (N_11741,N_8789,N_7683);
and U11742 (N_11742,N_6460,N_6894);
nand U11743 (N_11743,N_7031,N_6582);
nor U11744 (N_11744,N_8145,N_6688);
and U11745 (N_11745,N_8418,N_6370);
and U11746 (N_11746,N_9005,N_6598);
and U11747 (N_11747,N_6336,N_8444);
and U11748 (N_11748,N_9124,N_6373);
nand U11749 (N_11749,N_7178,N_8962);
nor U11750 (N_11750,N_8761,N_7277);
xor U11751 (N_11751,N_7191,N_9180);
and U11752 (N_11752,N_7241,N_8470);
nand U11753 (N_11753,N_7051,N_6866);
xnor U11754 (N_11754,N_7605,N_7564);
or U11755 (N_11755,N_6790,N_6442);
and U11756 (N_11756,N_9183,N_9329);
or U11757 (N_11757,N_7686,N_8758);
nor U11758 (N_11758,N_7951,N_7479);
nand U11759 (N_11759,N_7352,N_7892);
nor U11760 (N_11760,N_7956,N_7972);
and U11761 (N_11761,N_7007,N_8089);
and U11762 (N_11762,N_7357,N_8053);
or U11763 (N_11763,N_8486,N_6471);
or U11764 (N_11764,N_7960,N_8928);
nand U11765 (N_11765,N_8273,N_8021);
and U11766 (N_11766,N_8578,N_9080);
nand U11767 (N_11767,N_7167,N_8665);
nor U11768 (N_11768,N_9134,N_8262);
or U11769 (N_11769,N_7817,N_6807);
and U11770 (N_11770,N_8349,N_6659);
xor U11771 (N_11771,N_8246,N_6385);
xor U11772 (N_11772,N_8132,N_6837);
or U11773 (N_11773,N_8924,N_9021);
and U11774 (N_11774,N_9141,N_7053);
or U11775 (N_11775,N_7377,N_9231);
and U11776 (N_11776,N_6320,N_9072);
or U11777 (N_11777,N_6712,N_7422);
xnor U11778 (N_11778,N_6256,N_9104);
nand U11779 (N_11779,N_7904,N_8868);
nand U11780 (N_11780,N_8732,N_6517);
nand U11781 (N_11781,N_8347,N_7720);
or U11782 (N_11782,N_9288,N_6629);
nand U11783 (N_11783,N_7430,N_6313);
nand U11784 (N_11784,N_9023,N_8025);
nand U11785 (N_11785,N_8970,N_9230);
and U11786 (N_11786,N_6415,N_6644);
nand U11787 (N_11787,N_9131,N_7326);
nor U11788 (N_11788,N_8688,N_6325);
xnor U11789 (N_11789,N_7314,N_9343);
and U11790 (N_11790,N_7350,N_7030);
nor U11791 (N_11791,N_8471,N_9098);
nand U11792 (N_11792,N_7192,N_9122);
nand U11793 (N_11793,N_8304,N_7300);
nor U11794 (N_11794,N_6684,N_7545);
xor U11795 (N_11795,N_7006,N_6362);
and U11796 (N_11796,N_9049,N_6398);
nand U11797 (N_11797,N_7325,N_6578);
xor U11798 (N_11798,N_8067,N_8632);
xor U11799 (N_11799,N_7250,N_6943);
or U11800 (N_11800,N_8556,N_8681);
or U11801 (N_11801,N_7518,N_8790);
or U11802 (N_11802,N_8512,N_6714);
xnor U11803 (N_11803,N_7704,N_8558);
or U11804 (N_11804,N_7978,N_7946);
and U11805 (N_11805,N_6750,N_6601);
xnor U11806 (N_11806,N_8738,N_7145);
nor U11807 (N_11807,N_9130,N_7508);
nand U11808 (N_11808,N_9244,N_9051);
and U11809 (N_11809,N_8243,N_8182);
and U11810 (N_11810,N_7160,N_6965);
or U11811 (N_11811,N_8041,N_6614);
or U11812 (N_11812,N_8752,N_9166);
and U11813 (N_11813,N_8490,N_7802);
nand U11814 (N_11814,N_8794,N_6508);
nor U11815 (N_11815,N_8865,N_7842);
nand U11816 (N_11816,N_8037,N_8627);
nor U11817 (N_11817,N_7128,N_6545);
nor U11818 (N_11818,N_6855,N_6384);
nand U11819 (N_11819,N_8408,N_7945);
nand U11820 (N_11820,N_7647,N_7116);
and U11821 (N_11821,N_7151,N_6310);
xor U11822 (N_11822,N_7906,N_8656);
nor U11823 (N_11823,N_7048,N_7151);
nor U11824 (N_11824,N_7687,N_6613);
nand U11825 (N_11825,N_8123,N_6461);
xnor U11826 (N_11826,N_6670,N_7735);
xor U11827 (N_11827,N_7359,N_7022);
nor U11828 (N_11828,N_6435,N_8098);
nor U11829 (N_11829,N_8150,N_8640);
nand U11830 (N_11830,N_8495,N_7838);
or U11831 (N_11831,N_9134,N_6477);
nand U11832 (N_11832,N_6865,N_8058);
nor U11833 (N_11833,N_8725,N_6335);
or U11834 (N_11834,N_6707,N_8821);
nand U11835 (N_11835,N_6703,N_7770);
or U11836 (N_11836,N_6893,N_7226);
and U11837 (N_11837,N_7773,N_6336);
and U11838 (N_11838,N_8417,N_7047);
nor U11839 (N_11839,N_9098,N_6669);
nor U11840 (N_11840,N_9288,N_7101);
xnor U11841 (N_11841,N_8627,N_7196);
nor U11842 (N_11842,N_8777,N_6587);
nand U11843 (N_11843,N_8439,N_8161);
xor U11844 (N_11844,N_6898,N_6506);
xor U11845 (N_11845,N_6485,N_9270);
and U11846 (N_11846,N_8431,N_8805);
nand U11847 (N_11847,N_8958,N_7500);
nor U11848 (N_11848,N_8773,N_7660);
nor U11849 (N_11849,N_8869,N_6317);
xnor U11850 (N_11850,N_6551,N_7351);
or U11851 (N_11851,N_8485,N_6699);
xnor U11852 (N_11852,N_7682,N_6520);
nor U11853 (N_11853,N_7656,N_7369);
or U11854 (N_11854,N_8467,N_8858);
xnor U11855 (N_11855,N_8390,N_6842);
and U11856 (N_11856,N_8919,N_7252);
xnor U11857 (N_11857,N_6831,N_8567);
or U11858 (N_11858,N_6486,N_9181);
or U11859 (N_11859,N_9142,N_7756);
nor U11860 (N_11860,N_9191,N_7546);
xor U11861 (N_11861,N_6487,N_8982);
and U11862 (N_11862,N_6251,N_8476);
and U11863 (N_11863,N_6401,N_9100);
xnor U11864 (N_11864,N_6903,N_9127);
nand U11865 (N_11865,N_7060,N_7730);
nand U11866 (N_11866,N_6403,N_7836);
xnor U11867 (N_11867,N_9328,N_6832);
nand U11868 (N_11868,N_7738,N_8264);
or U11869 (N_11869,N_8448,N_7608);
nand U11870 (N_11870,N_8666,N_8794);
or U11871 (N_11871,N_9335,N_8028);
xnor U11872 (N_11872,N_6672,N_8575);
nand U11873 (N_11873,N_6957,N_6267);
nor U11874 (N_11874,N_9095,N_6427);
nor U11875 (N_11875,N_9241,N_7293);
xor U11876 (N_11876,N_6681,N_7836);
nand U11877 (N_11877,N_9083,N_9332);
and U11878 (N_11878,N_8257,N_9271);
and U11879 (N_11879,N_6348,N_8007);
or U11880 (N_11880,N_6667,N_7691);
and U11881 (N_11881,N_8027,N_7296);
xnor U11882 (N_11882,N_8914,N_8003);
or U11883 (N_11883,N_9374,N_6798);
nand U11884 (N_11884,N_8643,N_7111);
nor U11885 (N_11885,N_6750,N_7486);
or U11886 (N_11886,N_7714,N_6657);
and U11887 (N_11887,N_8035,N_7912);
nand U11888 (N_11888,N_6292,N_8549);
xnor U11889 (N_11889,N_7757,N_7328);
nand U11890 (N_11890,N_6860,N_8977);
xnor U11891 (N_11891,N_8862,N_8495);
nand U11892 (N_11892,N_8627,N_7618);
nor U11893 (N_11893,N_8815,N_9110);
nand U11894 (N_11894,N_7100,N_6986);
or U11895 (N_11895,N_8353,N_6795);
nand U11896 (N_11896,N_8072,N_8561);
nand U11897 (N_11897,N_6533,N_7787);
nand U11898 (N_11898,N_8943,N_6898);
nand U11899 (N_11899,N_8729,N_9111);
xnor U11900 (N_11900,N_7270,N_6513);
nand U11901 (N_11901,N_6274,N_8078);
nor U11902 (N_11902,N_7472,N_6262);
xor U11903 (N_11903,N_9149,N_7650);
xnor U11904 (N_11904,N_6338,N_9233);
xnor U11905 (N_11905,N_8268,N_7435);
xnor U11906 (N_11906,N_6689,N_6971);
or U11907 (N_11907,N_8122,N_8759);
or U11908 (N_11908,N_8731,N_7825);
nand U11909 (N_11909,N_8165,N_7637);
xor U11910 (N_11910,N_7859,N_9285);
and U11911 (N_11911,N_8736,N_7921);
nor U11912 (N_11912,N_8393,N_7467);
nand U11913 (N_11913,N_7244,N_7683);
or U11914 (N_11914,N_7914,N_6427);
nor U11915 (N_11915,N_8237,N_9253);
or U11916 (N_11916,N_8599,N_8475);
xnor U11917 (N_11917,N_8922,N_8951);
nor U11918 (N_11918,N_9063,N_6911);
and U11919 (N_11919,N_6644,N_7355);
and U11920 (N_11920,N_9349,N_9269);
or U11921 (N_11921,N_7154,N_9332);
or U11922 (N_11922,N_8390,N_6467);
or U11923 (N_11923,N_8080,N_8878);
nor U11924 (N_11924,N_8439,N_7513);
xor U11925 (N_11925,N_7441,N_8102);
xnor U11926 (N_11926,N_7827,N_8316);
or U11927 (N_11927,N_6679,N_8941);
xnor U11928 (N_11928,N_8659,N_8367);
nor U11929 (N_11929,N_6305,N_7945);
xor U11930 (N_11930,N_6459,N_9150);
and U11931 (N_11931,N_7990,N_6793);
or U11932 (N_11932,N_8258,N_7421);
nand U11933 (N_11933,N_7015,N_8894);
nor U11934 (N_11934,N_7155,N_9321);
xor U11935 (N_11935,N_6326,N_6439);
and U11936 (N_11936,N_9025,N_6928);
nor U11937 (N_11937,N_7912,N_9327);
nand U11938 (N_11938,N_7695,N_7010);
nand U11939 (N_11939,N_6285,N_6304);
and U11940 (N_11940,N_7013,N_8001);
xor U11941 (N_11941,N_7692,N_8239);
nand U11942 (N_11942,N_7704,N_9120);
and U11943 (N_11943,N_8344,N_7250);
nor U11944 (N_11944,N_6366,N_8076);
or U11945 (N_11945,N_6724,N_6990);
and U11946 (N_11946,N_7581,N_8425);
xor U11947 (N_11947,N_8353,N_8267);
nand U11948 (N_11948,N_8333,N_6283);
nand U11949 (N_11949,N_9227,N_7372);
or U11950 (N_11950,N_8483,N_7040);
nor U11951 (N_11951,N_8087,N_6617);
nor U11952 (N_11952,N_7324,N_6845);
or U11953 (N_11953,N_8036,N_9250);
xor U11954 (N_11954,N_7568,N_8067);
nand U11955 (N_11955,N_7388,N_9370);
nand U11956 (N_11956,N_7971,N_9347);
or U11957 (N_11957,N_7062,N_6254);
nor U11958 (N_11958,N_8805,N_8456);
nand U11959 (N_11959,N_9342,N_6348);
or U11960 (N_11960,N_9042,N_8331);
and U11961 (N_11961,N_7139,N_9269);
or U11962 (N_11962,N_7207,N_8550);
xnor U11963 (N_11963,N_7337,N_6501);
nor U11964 (N_11964,N_7259,N_6350);
xnor U11965 (N_11965,N_8727,N_6589);
and U11966 (N_11966,N_7231,N_9198);
and U11967 (N_11967,N_8009,N_8877);
and U11968 (N_11968,N_7283,N_7324);
and U11969 (N_11969,N_9144,N_9272);
or U11970 (N_11970,N_7200,N_8575);
nand U11971 (N_11971,N_6733,N_6521);
nor U11972 (N_11972,N_6854,N_8105);
and U11973 (N_11973,N_8357,N_8190);
or U11974 (N_11974,N_6409,N_6437);
or U11975 (N_11975,N_6424,N_7718);
or U11976 (N_11976,N_9136,N_6292);
xor U11977 (N_11977,N_9159,N_8612);
or U11978 (N_11978,N_8720,N_8549);
nor U11979 (N_11979,N_8984,N_8606);
nand U11980 (N_11980,N_6593,N_8404);
nor U11981 (N_11981,N_7192,N_6323);
nor U11982 (N_11982,N_8736,N_7946);
or U11983 (N_11983,N_8263,N_7806);
nand U11984 (N_11984,N_8351,N_8008);
or U11985 (N_11985,N_8220,N_8549);
nand U11986 (N_11986,N_6790,N_8694);
nor U11987 (N_11987,N_6929,N_8669);
xnor U11988 (N_11988,N_9111,N_8448);
xnor U11989 (N_11989,N_8556,N_6409);
or U11990 (N_11990,N_7692,N_6626);
nor U11991 (N_11991,N_8713,N_7387);
nor U11992 (N_11992,N_8578,N_8322);
xnor U11993 (N_11993,N_6557,N_7735);
xor U11994 (N_11994,N_6774,N_6715);
and U11995 (N_11995,N_6929,N_8681);
or U11996 (N_11996,N_7881,N_7388);
nand U11997 (N_11997,N_8449,N_7814);
or U11998 (N_11998,N_8036,N_6443);
nor U11999 (N_11999,N_8256,N_8774);
nand U12000 (N_12000,N_7130,N_7505);
xor U12001 (N_12001,N_8732,N_6363);
nor U12002 (N_12002,N_9104,N_6860);
nor U12003 (N_12003,N_7712,N_8369);
nand U12004 (N_12004,N_9012,N_8572);
nor U12005 (N_12005,N_7967,N_6756);
nand U12006 (N_12006,N_6846,N_6815);
and U12007 (N_12007,N_7631,N_7862);
nor U12008 (N_12008,N_9200,N_7429);
nand U12009 (N_12009,N_8299,N_6726);
xor U12010 (N_12010,N_8623,N_6286);
nor U12011 (N_12011,N_6425,N_9309);
or U12012 (N_12012,N_7977,N_8547);
nor U12013 (N_12013,N_7337,N_6768);
nor U12014 (N_12014,N_6476,N_9057);
nand U12015 (N_12015,N_8095,N_9128);
or U12016 (N_12016,N_7971,N_9013);
xor U12017 (N_12017,N_7095,N_6707);
or U12018 (N_12018,N_6902,N_7333);
xnor U12019 (N_12019,N_9269,N_8078);
and U12020 (N_12020,N_8819,N_9352);
nor U12021 (N_12021,N_7002,N_7266);
nand U12022 (N_12022,N_7701,N_6751);
nor U12023 (N_12023,N_7197,N_6364);
nor U12024 (N_12024,N_8101,N_6884);
nor U12025 (N_12025,N_7150,N_9036);
nand U12026 (N_12026,N_9271,N_9297);
xor U12027 (N_12027,N_9083,N_6492);
or U12028 (N_12028,N_9134,N_7752);
or U12029 (N_12029,N_8344,N_7377);
xnor U12030 (N_12030,N_9257,N_8716);
and U12031 (N_12031,N_8353,N_6591);
nor U12032 (N_12032,N_8927,N_8718);
xor U12033 (N_12033,N_6835,N_6606);
xnor U12034 (N_12034,N_8249,N_6605);
or U12035 (N_12035,N_8952,N_8948);
nor U12036 (N_12036,N_8414,N_6918);
and U12037 (N_12037,N_6691,N_8143);
nor U12038 (N_12038,N_8781,N_8195);
and U12039 (N_12039,N_7927,N_9341);
nor U12040 (N_12040,N_7645,N_8771);
xnor U12041 (N_12041,N_6356,N_9125);
xnor U12042 (N_12042,N_8877,N_8625);
xnor U12043 (N_12043,N_8350,N_6381);
xnor U12044 (N_12044,N_8383,N_7374);
xnor U12045 (N_12045,N_8754,N_8263);
nand U12046 (N_12046,N_7545,N_8838);
or U12047 (N_12047,N_8245,N_9051);
xor U12048 (N_12048,N_7192,N_7160);
and U12049 (N_12049,N_9002,N_8374);
and U12050 (N_12050,N_9238,N_6777);
xor U12051 (N_12051,N_6777,N_7174);
xor U12052 (N_12052,N_6623,N_8704);
nor U12053 (N_12053,N_8833,N_8204);
xor U12054 (N_12054,N_9243,N_8083);
nor U12055 (N_12055,N_6629,N_7128);
nand U12056 (N_12056,N_7184,N_6499);
xor U12057 (N_12057,N_7839,N_6561);
and U12058 (N_12058,N_6861,N_7709);
nor U12059 (N_12059,N_6720,N_8328);
and U12060 (N_12060,N_7950,N_7919);
or U12061 (N_12061,N_6792,N_8482);
xor U12062 (N_12062,N_7481,N_7573);
nand U12063 (N_12063,N_8324,N_7227);
nand U12064 (N_12064,N_7295,N_9321);
xnor U12065 (N_12065,N_6958,N_7396);
and U12066 (N_12066,N_8210,N_7361);
and U12067 (N_12067,N_8482,N_7254);
xnor U12068 (N_12068,N_8961,N_6451);
xnor U12069 (N_12069,N_8308,N_9087);
and U12070 (N_12070,N_9254,N_7625);
nor U12071 (N_12071,N_6427,N_8371);
nand U12072 (N_12072,N_8420,N_8615);
nand U12073 (N_12073,N_9271,N_6921);
nor U12074 (N_12074,N_8696,N_8027);
nor U12075 (N_12075,N_6885,N_9135);
or U12076 (N_12076,N_7675,N_7335);
nand U12077 (N_12077,N_8965,N_9101);
nor U12078 (N_12078,N_8144,N_9101);
or U12079 (N_12079,N_8484,N_7150);
xor U12080 (N_12080,N_6330,N_8805);
xor U12081 (N_12081,N_6837,N_7537);
and U12082 (N_12082,N_8117,N_8465);
nor U12083 (N_12083,N_8619,N_7873);
nand U12084 (N_12084,N_7864,N_9229);
or U12085 (N_12085,N_8252,N_7744);
nand U12086 (N_12086,N_7427,N_9161);
nor U12087 (N_12087,N_7023,N_8611);
nand U12088 (N_12088,N_7713,N_8278);
xnor U12089 (N_12089,N_8280,N_6531);
xor U12090 (N_12090,N_9213,N_7061);
and U12091 (N_12091,N_6611,N_6333);
nand U12092 (N_12092,N_8342,N_9231);
xor U12093 (N_12093,N_7148,N_9322);
and U12094 (N_12094,N_7589,N_7749);
xor U12095 (N_12095,N_7865,N_8834);
or U12096 (N_12096,N_6913,N_8399);
nor U12097 (N_12097,N_6921,N_8750);
xor U12098 (N_12098,N_7619,N_8705);
nor U12099 (N_12099,N_9369,N_8745);
nand U12100 (N_12100,N_8730,N_9145);
nor U12101 (N_12101,N_7930,N_8802);
nor U12102 (N_12102,N_6726,N_6395);
or U12103 (N_12103,N_8753,N_7555);
nor U12104 (N_12104,N_7196,N_6751);
xnor U12105 (N_12105,N_8337,N_8070);
nor U12106 (N_12106,N_6623,N_7045);
and U12107 (N_12107,N_9014,N_7252);
xnor U12108 (N_12108,N_8983,N_7219);
and U12109 (N_12109,N_8892,N_7619);
or U12110 (N_12110,N_7708,N_6283);
xnor U12111 (N_12111,N_6726,N_6491);
xnor U12112 (N_12112,N_6577,N_6924);
or U12113 (N_12113,N_8113,N_6980);
xor U12114 (N_12114,N_9119,N_8851);
xor U12115 (N_12115,N_8310,N_8370);
nand U12116 (N_12116,N_6483,N_8528);
and U12117 (N_12117,N_7209,N_9028);
or U12118 (N_12118,N_9116,N_7351);
xnor U12119 (N_12119,N_7928,N_7005);
nand U12120 (N_12120,N_9349,N_8110);
nand U12121 (N_12121,N_6680,N_7051);
or U12122 (N_12122,N_6895,N_6449);
nand U12123 (N_12123,N_7445,N_8244);
and U12124 (N_12124,N_6350,N_9040);
and U12125 (N_12125,N_6397,N_6855);
xnor U12126 (N_12126,N_9027,N_8173);
and U12127 (N_12127,N_7824,N_6272);
nand U12128 (N_12128,N_8249,N_7663);
or U12129 (N_12129,N_9125,N_8464);
and U12130 (N_12130,N_8907,N_9353);
nor U12131 (N_12131,N_6286,N_6353);
nand U12132 (N_12132,N_7026,N_8360);
nand U12133 (N_12133,N_6345,N_7644);
or U12134 (N_12134,N_8855,N_7688);
xor U12135 (N_12135,N_6758,N_6492);
xor U12136 (N_12136,N_8029,N_8245);
xor U12137 (N_12137,N_9076,N_6258);
xnor U12138 (N_12138,N_8153,N_7286);
nand U12139 (N_12139,N_6733,N_6413);
and U12140 (N_12140,N_8421,N_9309);
nor U12141 (N_12141,N_7513,N_6987);
nor U12142 (N_12142,N_9132,N_6395);
and U12143 (N_12143,N_6825,N_6656);
and U12144 (N_12144,N_8391,N_8489);
or U12145 (N_12145,N_6977,N_7754);
or U12146 (N_12146,N_7768,N_8922);
nor U12147 (N_12147,N_7666,N_7114);
nor U12148 (N_12148,N_8001,N_6759);
or U12149 (N_12149,N_8912,N_7653);
and U12150 (N_12150,N_8897,N_8230);
nor U12151 (N_12151,N_8929,N_8095);
nor U12152 (N_12152,N_8978,N_7634);
xnor U12153 (N_12153,N_7858,N_7846);
xnor U12154 (N_12154,N_7531,N_7756);
and U12155 (N_12155,N_7347,N_7876);
nor U12156 (N_12156,N_8636,N_6887);
nand U12157 (N_12157,N_8984,N_8219);
nor U12158 (N_12158,N_8217,N_7697);
or U12159 (N_12159,N_7835,N_6616);
and U12160 (N_12160,N_9309,N_7731);
nand U12161 (N_12161,N_8347,N_9176);
xor U12162 (N_12162,N_7802,N_7295);
or U12163 (N_12163,N_8623,N_7821);
or U12164 (N_12164,N_6425,N_8814);
nand U12165 (N_12165,N_9250,N_6870);
xor U12166 (N_12166,N_6547,N_6940);
nand U12167 (N_12167,N_8190,N_6876);
nand U12168 (N_12168,N_8055,N_7577);
xnor U12169 (N_12169,N_7289,N_8908);
nor U12170 (N_12170,N_8801,N_8995);
nor U12171 (N_12171,N_7100,N_6720);
and U12172 (N_12172,N_8927,N_7894);
or U12173 (N_12173,N_9175,N_6272);
or U12174 (N_12174,N_7179,N_8889);
or U12175 (N_12175,N_6704,N_9160);
and U12176 (N_12176,N_9155,N_6838);
xor U12177 (N_12177,N_8672,N_9216);
xor U12178 (N_12178,N_7216,N_7923);
and U12179 (N_12179,N_7618,N_6539);
or U12180 (N_12180,N_7200,N_7908);
nor U12181 (N_12181,N_7044,N_7636);
or U12182 (N_12182,N_9360,N_6538);
or U12183 (N_12183,N_8750,N_8828);
nand U12184 (N_12184,N_7669,N_6909);
or U12185 (N_12185,N_8749,N_6630);
and U12186 (N_12186,N_6921,N_9361);
nand U12187 (N_12187,N_7357,N_8899);
or U12188 (N_12188,N_8858,N_6336);
and U12189 (N_12189,N_6902,N_7668);
nand U12190 (N_12190,N_7381,N_9286);
or U12191 (N_12191,N_9143,N_8734);
or U12192 (N_12192,N_6776,N_6728);
nor U12193 (N_12193,N_6828,N_7906);
nand U12194 (N_12194,N_8343,N_7252);
nor U12195 (N_12195,N_7865,N_9006);
or U12196 (N_12196,N_7225,N_6585);
or U12197 (N_12197,N_7184,N_7952);
nor U12198 (N_12198,N_7807,N_6369);
nand U12199 (N_12199,N_8380,N_6949);
or U12200 (N_12200,N_7306,N_7307);
nand U12201 (N_12201,N_9304,N_7383);
nand U12202 (N_12202,N_6935,N_7772);
and U12203 (N_12203,N_7603,N_6926);
nor U12204 (N_12204,N_7349,N_9070);
nor U12205 (N_12205,N_7755,N_8765);
and U12206 (N_12206,N_6281,N_6477);
xnor U12207 (N_12207,N_7969,N_6455);
xnor U12208 (N_12208,N_7965,N_6703);
xnor U12209 (N_12209,N_7993,N_7818);
nand U12210 (N_12210,N_8927,N_8276);
nor U12211 (N_12211,N_8355,N_8791);
nand U12212 (N_12212,N_8286,N_6957);
nand U12213 (N_12213,N_6256,N_6791);
nand U12214 (N_12214,N_6912,N_8225);
xor U12215 (N_12215,N_7972,N_6535);
xnor U12216 (N_12216,N_6869,N_7297);
nor U12217 (N_12217,N_7116,N_8405);
nor U12218 (N_12218,N_7977,N_6577);
xor U12219 (N_12219,N_6936,N_6850);
and U12220 (N_12220,N_8878,N_8447);
nor U12221 (N_12221,N_7715,N_7813);
nand U12222 (N_12222,N_7338,N_7211);
and U12223 (N_12223,N_8933,N_6390);
nor U12224 (N_12224,N_8017,N_7789);
xor U12225 (N_12225,N_8886,N_8432);
or U12226 (N_12226,N_6943,N_6648);
nand U12227 (N_12227,N_9179,N_8127);
and U12228 (N_12228,N_7286,N_7476);
nor U12229 (N_12229,N_7427,N_8833);
or U12230 (N_12230,N_6856,N_6761);
or U12231 (N_12231,N_7188,N_7112);
and U12232 (N_12232,N_8157,N_8518);
xnor U12233 (N_12233,N_8241,N_7442);
and U12234 (N_12234,N_8201,N_7186);
nand U12235 (N_12235,N_8078,N_8659);
nand U12236 (N_12236,N_8890,N_8453);
nand U12237 (N_12237,N_8652,N_7950);
or U12238 (N_12238,N_8521,N_7617);
nor U12239 (N_12239,N_7276,N_8685);
or U12240 (N_12240,N_8978,N_7151);
nor U12241 (N_12241,N_6833,N_6314);
xor U12242 (N_12242,N_8711,N_7193);
or U12243 (N_12243,N_6774,N_8744);
xnor U12244 (N_12244,N_7163,N_6612);
nor U12245 (N_12245,N_6320,N_8209);
and U12246 (N_12246,N_9282,N_6376);
and U12247 (N_12247,N_8291,N_8462);
xor U12248 (N_12248,N_8959,N_7515);
xor U12249 (N_12249,N_7004,N_9238);
and U12250 (N_12250,N_8533,N_7969);
nand U12251 (N_12251,N_7402,N_7938);
nor U12252 (N_12252,N_7253,N_9153);
xnor U12253 (N_12253,N_7061,N_8575);
or U12254 (N_12254,N_6475,N_9074);
and U12255 (N_12255,N_6479,N_7702);
or U12256 (N_12256,N_9182,N_7328);
or U12257 (N_12257,N_8119,N_6726);
xor U12258 (N_12258,N_9027,N_6968);
and U12259 (N_12259,N_7670,N_8034);
and U12260 (N_12260,N_7310,N_8662);
and U12261 (N_12261,N_7040,N_7033);
xor U12262 (N_12262,N_8218,N_8477);
or U12263 (N_12263,N_6817,N_7099);
xor U12264 (N_12264,N_7840,N_7964);
nand U12265 (N_12265,N_7331,N_8013);
nand U12266 (N_12266,N_7024,N_7010);
and U12267 (N_12267,N_7233,N_9022);
xor U12268 (N_12268,N_8550,N_8527);
and U12269 (N_12269,N_8083,N_8967);
xor U12270 (N_12270,N_8005,N_8572);
or U12271 (N_12271,N_8792,N_9008);
or U12272 (N_12272,N_7409,N_7595);
or U12273 (N_12273,N_9149,N_8954);
nand U12274 (N_12274,N_8539,N_6759);
or U12275 (N_12275,N_6836,N_6717);
and U12276 (N_12276,N_6653,N_7155);
nor U12277 (N_12277,N_7369,N_8005);
nand U12278 (N_12278,N_8773,N_9374);
nor U12279 (N_12279,N_7302,N_7973);
xnor U12280 (N_12280,N_9246,N_7321);
nor U12281 (N_12281,N_9063,N_6595);
nand U12282 (N_12282,N_6787,N_6768);
and U12283 (N_12283,N_6467,N_7752);
or U12284 (N_12284,N_7001,N_8774);
nand U12285 (N_12285,N_8455,N_7864);
nand U12286 (N_12286,N_8550,N_8909);
nor U12287 (N_12287,N_6279,N_9053);
nor U12288 (N_12288,N_6882,N_7297);
nand U12289 (N_12289,N_6746,N_9329);
or U12290 (N_12290,N_9107,N_8922);
nand U12291 (N_12291,N_7834,N_9286);
xnor U12292 (N_12292,N_7220,N_9146);
and U12293 (N_12293,N_9252,N_8862);
or U12294 (N_12294,N_6389,N_8656);
and U12295 (N_12295,N_7328,N_7726);
nand U12296 (N_12296,N_6254,N_8378);
nand U12297 (N_12297,N_7303,N_9005);
and U12298 (N_12298,N_8868,N_7404);
or U12299 (N_12299,N_8671,N_8162);
and U12300 (N_12300,N_9136,N_7152);
or U12301 (N_12301,N_7047,N_9084);
xor U12302 (N_12302,N_6565,N_7871);
and U12303 (N_12303,N_6652,N_8519);
nand U12304 (N_12304,N_8676,N_8827);
nor U12305 (N_12305,N_7926,N_7670);
xor U12306 (N_12306,N_9097,N_6337);
nor U12307 (N_12307,N_6828,N_7064);
xnor U12308 (N_12308,N_8551,N_6778);
nor U12309 (N_12309,N_7151,N_6689);
or U12310 (N_12310,N_6275,N_8484);
or U12311 (N_12311,N_9211,N_7157);
nand U12312 (N_12312,N_6807,N_6299);
nor U12313 (N_12313,N_7208,N_7223);
or U12314 (N_12314,N_6759,N_8068);
nor U12315 (N_12315,N_7498,N_7843);
xnor U12316 (N_12316,N_6481,N_7742);
nor U12317 (N_12317,N_6599,N_7120);
xor U12318 (N_12318,N_6476,N_8752);
xnor U12319 (N_12319,N_9282,N_8565);
xor U12320 (N_12320,N_7473,N_7227);
xnor U12321 (N_12321,N_8535,N_8416);
nand U12322 (N_12322,N_8198,N_7379);
xnor U12323 (N_12323,N_7343,N_9268);
nor U12324 (N_12324,N_8829,N_6597);
nand U12325 (N_12325,N_8288,N_7957);
xnor U12326 (N_12326,N_8809,N_8704);
xor U12327 (N_12327,N_9091,N_7255);
nor U12328 (N_12328,N_7253,N_6388);
and U12329 (N_12329,N_6913,N_6879);
nor U12330 (N_12330,N_6925,N_8203);
xnor U12331 (N_12331,N_7519,N_8441);
xnor U12332 (N_12332,N_6443,N_7589);
nor U12333 (N_12333,N_7798,N_7509);
nor U12334 (N_12334,N_7822,N_6757);
nand U12335 (N_12335,N_8895,N_6892);
nand U12336 (N_12336,N_8634,N_6379);
and U12337 (N_12337,N_7387,N_6781);
and U12338 (N_12338,N_6814,N_7331);
or U12339 (N_12339,N_7803,N_7184);
nand U12340 (N_12340,N_8780,N_8051);
and U12341 (N_12341,N_9033,N_7175);
nor U12342 (N_12342,N_6358,N_7366);
or U12343 (N_12343,N_8053,N_8475);
nand U12344 (N_12344,N_6287,N_6526);
nor U12345 (N_12345,N_8089,N_7124);
nand U12346 (N_12346,N_6676,N_7454);
nor U12347 (N_12347,N_9246,N_7093);
and U12348 (N_12348,N_6636,N_7193);
nor U12349 (N_12349,N_6265,N_7354);
and U12350 (N_12350,N_8401,N_6411);
nand U12351 (N_12351,N_7701,N_8205);
or U12352 (N_12352,N_8081,N_7494);
or U12353 (N_12353,N_7862,N_8776);
or U12354 (N_12354,N_7753,N_6965);
nand U12355 (N_12355,N_7902,N_6489);
xnor U12356 (N_12356,N_6930,N_8243);
and U12357 (N_12357,N_9246,N_8431);
and U12358 (N_12358,N_7786,N_9175);
and U12359 (N_12359,N_6386,N_9091);
or U12360 (N_12360,N_7467,N_6535);
xnor U12361 (N_12361,N_6275,N_7361);
nand U12362 (N_12362,N_9047,N_6990);
nand U12363 (N_12363,N_7084,N_7506);
nor U12364 (N_12364,N_7958,N_8270);
and U12365 (N_12365,N_8238,N_8673);
or U12366 (N_12366,N_7263,N_8805);
xor U12367 (N_12367,N_7476,N_7455);
xnor U12368 (N_12368,N_9034,N_6978);
xnor U12369 (N_12369,N_8196,N_7168);
or U12370 (N_12370,N_9096,N_6796);
and U12371 (N_12371,N_8859,N_7368);
xnor U12372 (N_12372,N_7079,N_6650);
nand U12373 (N_12373,N_6769,N_8859);
and U12374 (N_12374,N_7202,N_8621);
xor U12375 (N_12375,N_7194,N_6911);
and U12376 (N_12376,N_8314,N_7877);
or U12377 (N_12377,N_8017,N_7610);
and U12378 (N_12378,N_6987,N_9297);
nand U12379 (N_12379,N_7676,N_7573);
or U12380 (N_12380,N_7818,N_9074);
xor U12381 (N_12381,N_6333,N_8381);
xor U12382 (N_12382,N_7065,N_7285);
nor U12383 (N_12383,N_6671,N_7172);
xnor U12384 (N_12384,N_8122,N_6340);
nand U12385 (N_12385,N_7858,N_6676);
or U12386 (N_12386,N_6557,N_7881);
or U12387 (N_12387,N_8170,N_7568);
nor U12388 (N_12388,N_9119,N_9236);
xnor U12389 (N_12389,N_9332,N_7826);
and U12390 (N_12390,N_7406,N_8240);
and U12391 (N_12391,N_6931,N_7765);
nand U12392 (N_12392,N_6345,N_9085);
nor U12393 (N_12393,N_8243,N_7338);
nor U12394 (N_12394,N_8779,N_7958);
nor U12395 (N_12395,N_8875,N_6380);
xor U12396 (N_12396,N_7902,N_9148);
xor U12397 (N_12397,N_9076,N_8907);
xnor U12398 (N_12398,N_7908,N_8917);
nand U12399 (N_12399,N_6677,N_8411);
and U12400 (N_12400,N_6253,N_7927);
nor U12401 (N_12401,N_8999,N_6963);
xor U12402 (N_12402,N_6414,N_7799);
and U12403 (N_12403,N_6689,N_6550);
and U12404 (N_12404,N_9310,N_7463);
xor U12405 (N_12405,N_7344,N_8132);
or U12406 (N_12406,N_9019,N_9374);
xor U12407 (N_12407,N_8200,N_7464);
xor U12408 (N_12408,N_8626,N_9200);
or U12409 (N_12409,N_7602,N_6754);
nand U12410 (N_12410,N_9019,N_6452);
nor U12411 (N_12411,N_8225,N_7459);
nor U12412 (N_12412,N_7540,N_6314);
xnor U12413 (N_12413,N_6551,N_8808);
and U12414 (N_12414,N_7606,N_6252);
or U12415 (N_12415,N_7940,N_8140);
or U12416 (N_12416,N_7264,N_8882);
and U12417 (N_12417,N_8153,N_6455);
nor U12418 (N_12418,N_6748,N_7873);
nor U12419 (N_12419,N_7286,N_8779);
and U12420 (N_12420,N_8152,N_6501);
or U12421 (N_12421,N_8190,N_6459);
nand U12422 (N_12422,N_7560,N_7954);
xor U12423 (N_12423,N_7680,N_8056);
and U12424 (N_12424,N_8733,N_8901);
or U12425 (N_12425,N_7999,N_8299);
and U12426 (N_12426,N_8442,N_6513);
nand U12427 (N_12427,N_7651,N_8359);
xor U12428 (N_12428,N_7456,N_6747);
xor U12429 (N_12429,N_8052,N_7199);
nor U12430 (N_12430,N_7482,N_6561);
nand U12431 (N_12431,N_7548,N_8718);
nand U12432 (N_12432,N_9060,N_8679);
xor U12433 (N_12433,N_8479,N_7606);
xor U12434 (N_12434,N_7019,N_7375);
or U12435 (N_12435,N_9141,N_8501);
nor U12436 (N_12436,N_8077,N_9107);
and U12437 (N_12437,N_6393,N_8829);
or U12438 (N_12438,N_7798,N_6931);
nand U12439 (N_12439,N_7852,N_9115);
and U12440 (N_12440,N_7515,N_7234);
xnor U12441 (N_12441,N_7026,N_6705);
xor U12442 (N_12442,N_7710,N_9246);
nand U12443 (N_12443,N_6722,N_7039);
nor U12444 (N_12444,N_6818,N_9002);
nand U12445 (N_12445,N_7133,N_6468);
xnor U12446 (N_12446,N_9251,N_8792);
nor U12447 (N_12447,N_8629,N_6957);
nor U12448 (N_12448,N_8743,N_6310);
and U12449 (N_12449,N_8394,N_6322);
nor U12450 (N_12450,N_7243,N_7058);
and U12451 (N_12451,N_7447,N_6744);
nor U12452 (N_12452,N_8774,N_8477);
nor U12453 (N_12453,N_6415,N_8620);
or U12454 (N_12454,N_8660,N_8616);
nand U12455 (N_12455,N_9160,N_6775);
nand U12456 (N_12456,N_8215,N_7516);
and U12457 (N_12457,N_7117,N_8393);
xor U12458 (N_12458,N_9030,N_8742);
nor U12459 (N_12459,N_7675,N_8181);
or U12460 (N_12460,N_8620,N_6653);
and U12461 (N_12461,N_9269,N_7600);
and U12462 (N_12462,N_6846,N_9303);
and U12463 (N_12463,N_8129,N_7216);
xor U12464 (N_12464,N_6331,N_6315);
or U12465 (N_12465,N_7279,N_6973);
and U12466 (N_12466,N_6782,N_6592);
and U12467 (N_12467,N_7961,N_8559);
nor U12468 (N_12468,N_7498,N_7244);
and U12469 (N_12469,N_6541,N_9217);
and U12470 (N_12470,N_7077,N_8306);
and U12471 (N_12471,N_8433,N_7769);
and U12472 (N_12472,N_8241,N_7248);
nand U12473 (N_12473,N_6626,N_7529);
and U12474 (N_12474,N_9263,N_8024);
or U12475 (N_12475,N_9374,N_9184);
xor U12476 (N_12476,N_8181,N_9322);
nor U12477 (N_12477,N_7075,N_7287);
and U12478 (N_12478,N_8760,N_9321);
or U12479 (N_12479,N_8464,N_6525);
nand U12480 (N_12480,N_7036,N_7904);
nand U12481 (N_12481,N_6894,N_6795);
or U12482 (N_12482,N_8369,N_7391);
xnor U12483 (N_12483,N_8570,N_7462);
and U12484 (N_12484,N_8463,N_8857);
and U12485 (N_12485,N_7178,N_8173);
nor U12486 (N_12486,N_9209,N_8638);
xnor U12487 (N_12487,N_7700,N_6974);
nand U12488 (N_12488,N_6552,N_9278);
nor U12489 (N_12489,N_7887,N_8805);
nand U12490 (N_12490,N_9088,N_8382);
xnor U12491 (N_12491,N_8105,N_7771);
nand U12492 (N_12492,N_8488,N_9011);
or U12493 (N_12493,N_7739,N_9183);
and U12494 (N_12494,N_6593,N_6935);
or U12495 (N_12495,N_6625,N_9303);
nand U12496 (N_12496,N_7752,N_7795);
nor U12497 (N_12497,N_7348,N_8344);
xor U12498 (N_12498,N_8606,N_7085);
xor U12499 (N_12499,N_6252,N_7057);
nand U12500 (N_12500,N_11114,N_10670);
nand U12501 (N_12501,N_10004,N_11454);
or U12502 (N_12502,N_10357,N_10972);
or U12503 (N_12503,N_12201,N_12081);
or U12504 (N_12504,N_11063,N_9692);
xor U12505 (N_12505,N_12225,N_12262);
nor U12506 (N_12506,N_9887,N_11138);
or U12507 (N_12507,N_12352,N_11102);
nand U12508 (N_12508,N_10784,N_11959);
xnor U12509 (N_12509,N_12306,N_10551);
xor U12510 (N_12510,N_11061,N_9900);
nor U12511 (N_12511,N_11194,N_11319);
nor U12512 (N_12512,N_9921,N_11237);
xor U12513 (N_12513,N_12316,N_11464);
nand U12514 (N_12514,N_10309,N_9712);
nand U12515 (N_12515,N_9396,N_10960);
and U12516 (N_12516,N_11879,N_11128);
nand U12517 (N_12517,N_9731,N_10312);
or U12518 (N_12518,N_10778,N_9820);
and U12519 (N_12519,N_12180,N_10448);
xor U12520 (N_12520,N_11793,N_11487);
and U12521 (N_12521,N_9930,N_12181);
and U12522 (N_12522,N_11926,N_10292);
nor U12523 (N_12523,N_9399,N_10885);
xnor U12524 (N_12524,N_9536,N_11191);
and U12525 (N_12525,N_10411,N_10400);
or U12526 (N_12526,N_9628,N_10123);
nor U12527 (N_12527,N_9836,N_10911);
xnor U12528 (N_12528,N_9817,N_9436);
nor U12529 (N_12529,N_11505,N_10503);
or U12530 (N_12530,N_11069,N_10907);
nand U12531 (N_12531,N_11636,N_11170);
or U12532 (N_12532,N_10043,N_12458);
xor U12533 (N_12533,N_9734,N_10919);
or U12534 (N_12534,N_12084,N_12336);
nand U12535 (N_12535,N_11355,N_11028);
nor U12536 (N_12536,N_11484,N_11417);
xnor U12537 (N_12537,N_11184,N_10163);
nor U12538 (N_12538,N_9579,N_11056);
and U12539 (N_12539,N_9393,N_11157);
nand U12540 (N_12540,N_12011,N_10086);
xor U12541 (N_12541,N_12270,N_11088);
xnor U12542 (N_12542,N_12043,N_11285);
and U12543 (N_12543,N_11052,N_9658);
nor U12544 (N_12544,N_10042,N_12140);
nor U12545 (N_12545,N_9869,N_11267);
nand U12546 (N_12546,N_12328,N_10903);
xnor U12547 (N_12547,N_10208,N_10867);
nand U12548 (N_12548,N_12155,N_11305);
nand U12549 (N_12549,N_10639,N_11329);
xor U12550 (N_12550,N_11299,N_11480);
xor U12551 (N_12551,N_10101,N_9621);
and U12552 (N_12552,N_11385,N_12191);
nand U12553 (N_12553,N_10037,N_10876);
nor U12554 (N_12554,N_10809,N_10359);
nand U12555 (N_12555,N_11707,N_10017);
nor U12556 (N_12556,N_11670,N_12068);
xor U12557 (N_12557,N_10437,N_11440);
xnor U12558 (N_12558,N_11397,N_12094);
or U12559 (N_12559,N_10446,N_10317);
nor U12560 (N_12560,N_10612,N_11694);
or U12561 (N_12561,N_11593,N_11991);
or U12562 (N_12562,N_9980,N_12055);
nor U12563 (N_12563,N_10757,N_11569);
xnor U12564 (N_12564,N_12038,N_11451);
xnor U12565 (N_12565,N_10290,N_10527);
or U12566 (N_12566,N_12044,N_10112);
xor U12567 (N_12567,N_11378,N_10274);
and U12568 (N_12568,N_11485,N_9497);
and U12569 (N_12569,N_9610,N_11337);
or U12570 (N_12570,N_12331,N_9480);
or U12571 (N_12571,N_12431,N_9860);
or U12572 (N_12572,N_9433,N_10692);
nor U12573 (N_12573,N_12188,N_9764);
or U12574 (N_12574,N_10015,N_11024);
xnor U12575 (N_12575,N_12279,N_10891);
or U12576 (N_12576,N_9459,N_10439);
and U12577 (N_12577,N_10774,N_10303);
xnor U12578 (N_12578,N_10477,N_9496);
or U12579 (N_12579,N_10811,N_11546);
or U12580 (N_12580,N_11641,N_11716);
and U12581 (N_12581,N_9384,N_10839);
nand U12582 (N_12582,N_11021,N_12436);
nand U12583 (N_12583,N_11394,N_9704);
or U12584 (N_12584,N_9495,N_11403);
xnor U12585 (N_12585,N_12173,N_10873);
and U12586 (N_12586,N_11291,N_11616);
or U12587 (N_12587,N_11116,N_9729);
or U12588 (N_12588,N_9758,N_9455);
or U12589 (N_12589,N_9680,N_10151);
xor U12590 (N_12590,N_10736,N_12144);
and U12591 (N_12591,N_9924,N_10041);
xnor U12592 (N_12592,N_10080,N_9961);
or U12593 (N_12593,N_9407,N_10744);
nor U12594 (N_12594,N_12338,N_10866);
xnor U12595 (N_12595,N_11911,N_11696);
nor U12596 (N_12596,N_11055,N_9632);
nor U12597 (N_12597,N_12477,N_11025);
xnor U12598 (N_12598,N_10065,N_12227);
nand U12599 (N_12599,N_12365,N_11836);
nand U12600 (N_12600,N_10022,N_11545);
and U12601 (N_12601,N_11014,N_9504);
and U12602 (N_12602,N_11527,N_10170);
nor U12603 (N_12603,N_9406,N_9792);
or U12604 (N_12604,N_9730,N_10645);
nor U12605 (N_12605,N_11703,N_12112);
nand U12606 (N_12606,N_11441,N_9614);
and U12607 (N_12607,N_10767,N_10643);
xnor U12608 (N_12608,N_10728,N_11121);
or U12609 (N_12609,N_11995,N_9761);
or U12610 (N_12610,N_10630,N_11872);
xor U12611 (N_12611,N_10013,N_10376);
nand U12612 (N_12612,N_11691,N_9886);
xor U12613 (N_12613,N_9834,N_10030);
or U12614 (N_12614,N_9700,N_12473);
xor U12615 (N_12615,N_9772,N_10273);
nand U12616 (N_12616,N_10646,N_11969);
and U12617 (N_12617,N_10150,N_10828);
or U12618 (N_12618,N_10032,N_10063);
and U12619 (N_12619,N_11033,N_11177);
xor U12620 (N_12620,N_12080,N_11574);
nand U12621 (N_12621,N_10194,N_12162);
xnor U12622 (N_12622,N_10009,N_9796);
or U12623 (N_12623,N_10191,N_11073);
nor U12624 (N_12624,N_12207,N_10029);
xnor U12625 (N_12625,N_10501,N_12122);
nor U12626 (N_12626,N_11706,N_10351);
nor U12627 (N_12627,N_10588,N_10272);
or U12628 (N_12628,N_11017,N_10978);
or U12629 (N_12629,N_10668,N_11940);
nor U12630 (N_12630,N_11763,N_11791);
nor U12631 (N_12631,N_10936,N_11218);
or U12632 (N_12632,N_10912,N_11445);
xnor U12633 (N_12633,N_9681,N_10653);
nand U12634 (N_12634,N_11825,N_11185);
or U12635 (N_12635,N_11970,N_9460);
or U12636 (N_12636,N_10817,N_10563);
nor U12637 (N_12637,N_9677,N_9956);
or U12638 (N_12638,N_11765,N_10723);
nand U12639 (N_12639,N_11898,N_9878);
nor U12640 (N_12640,N_11475,N_9893);
nand U12641 (N_12641,N_11111,N_10768);
xnor U12642 (N_12642,N_11743,N_11284);
nor U12643 (N_12643,N_9419,N_11556);
and U12644 (N_12644,N_11080,N_11226);
nor U12645 (N_12645,N_11809,N_11346);
xor U12646 (N_12646,N_12424,N_11096);
or U12647 (N_12647,N_12102,N_10896);
xor U12648 (N_12648,N_10339,N_11684);
nor U12649 (N_12649,N_11119,N_11231);
and U12650 (N_12650,N_12493,N_9483);
or U12651 (N_12651,N_11753,N_10368);
and U12652 (N_12652,N_9951,N_10661);
nor U12653 (N_12653,N_12242,N_12288);
nor U12654 (N_12654,N_9935,N_10000);
or U12655 (N_12655,N_10350,N_12077);
or U12656 (N_12656,N_10417,N_10347);
xnor U12657 (N_12657,N_11453,N_11203);
xnor U12658 (N_12658,N_11726,N_11676);
nand U12659 (N_12659,N_10314,N_11386);
nand U12660 (N_12660,N_11018,N_10372);
nor U12661 (N_12661,N_10302,N_12375);
or U12662 (N_12662,N_10933,N_12111);
xnor U12663 (N_12663,N_9762,N_9735);
and U12664 (N_12664,N_10924,N_11223);
and U12665 (N_12665,N_10566,N_10628);
xor U12666 (N_12666,N_9911,N_11901);
or U12667 (N_12667,N_10522,N_11134);
nand U12668 (N_12668,N_10341,N_11054);
nor U12669 (N_12669,N_11927,N_10613);
xor U12670 (N_12670,N_10980,N_12048);
nor U12671 (N_12671,N_11534,N_11605);
xnor U12672 (N_12672,N_10586,N_10363);
nor U12673 (N_12673,N_12017,N_11622);
xnor U12674 (N_12674,N_11614,N_11428);
nor U12675 (N_12675,N_10199,N_9847);
or U12676 (N_12676,N_9793,N_10861);
and U12677 (N_12677,N_10326,N_10794);
xnor U12678 (N_12678,N_10733,N_9975);
and U12679 (N_12679,N_10930,N_10082);
nor U12680 (N_12680,N_12298,N_12070);
xor U12681 (N_12681,N_12009,N_9958);
and U12682 (N_12682,N_9616,N_9804);
xor U12683 (N_12683,N_10033,N_9615);
or U12684 (N_12684,N_10674,N_11795);
and U12685 (N_12685,N_9376,N_12247);
or U12686 (N_12686,N_10829,N_10633);
nor U12687 (N_12687,N_12313,N_12029);
nand U12688 (N_12688,N_10548,N_9432);
nor U12689 (N_12689,N_9840,N_10810);
and U12690 (N_12690,N_11921,N_10718);
nor U12691 (N_12691,N_9863,N_11681);
nor U12692 (N_12692,N_10739,N_9806);
or U12693 (N_12693,N_9412,N_10462);
xor U12694 (N_12694,N_10620,N_11243);
and U12695 (N_12695,N_9612,N_10178);
xnor U12696 (N_12696,N_10765,N_10556);
nor U12697 (N_12697,N_10619,N_10508);
or U12698 (N_12698,N_10815,N_12360);
or U12699 (N_12699,N_9414,N_11729);
or U12700 (N_12700,N_11235,N_11196);
nor U12701 (N_12701,N_11875,N_11234);
and U12702 (N_12702,N_11679,N_9383);
and U12703 (N_12703,N_9994,N_9623);
or U12704 (N_12704,N_12065,N_11971);
and U12705 (N_12705,N_10301,N_9583);
nor U12706 (N_12706,N_12039,N_10088);
nor U12707 (N_12707,N_10231,N_12129);
nor U12708 (N_12708,N_12350,N_11678);
or U12709 (N_12709,N_12362,N_11976);
nand U12710 (N_12710,N_12071,N_11934);
and U12711 (N_12711,N_12151,N_11294);
and U12712 (N_12712,N_9848,N_10550);
or U12713 (N_12713,N_11297,N_11816);
or U12714 (N_12714,N_10324,N_10939);
and U12715 (N_12715,N_11738,N_9776);
nor U12716 (N_12716,N_11702,N_11788);
nor U12717 (N_12717,N_9413,N_11731);
or U12718 (N_12718,N_11381,N_11987);
nor U12719 (N_12719,N_9473,N_11576);
nand U12720 (N_12720,N_11190,N_11032);
nand U12721 (N_12721,N_9919,N_9852);
nand U12722 (N_12722,N_9688,N_10313);
xor U12723 (N_12723,N_10141,N_10844);
xnor U12724 (N_12724,N_10111,N_9998);
nand U12725 (N_12725,N_10783,N_11986);
nor U12726 (N_12726,N_9589,N_10605);
and U12727 (N_12727,N_12281,N_10254);
nor U12728 (N_12728,N_10860,N_12491);
nand U12729 (N_12729,N_10971,N_11952);
or U12730 (N_12730,N_10944,N_11333);
nor U12731 (N_12731,N_12257,N_11239);
nor U12732 (N_12732,N_10246,N_10893);
xor U12733 (N_12733,N_10897,N_12303);
or U12734 (N_12734,N_11950,N_11476);
and U12735 (N_12735,N_11369,N_10460);
or U12736 (N_12736,N_11388,N_9445);
nand U12737 (N_12737,N_12294,N_12437);
or U12738 (N_12738,N_11876,N_12013);
xor U12739 (N_12739,N_9596,N_11529);
nor U12740 (N_12740,N_11800,N_10174);
nor U12741 (N_12741,N_10295,N_11640);
nand U12742 (N_12742,N_11813,N_12185);
or U12743 (N_12743,N_10571,N_11083);
nor U12744 (N_12744,N_10077,N_10489);
and U12745 (N_12745,N_12104,N_12445);
nor U12746 (N_12746,N_9894,N_10909);
nand U12747 (N_12747,N_11060,N_9442);
or U12748 (N_12748,N_12409,N_10917);
nor U12749 (N_12749,N_10179,N_11618);
or U12750 (N_12750,N_10190,N_9563);
xor U12751 (N_12751,N_10904,N_10663);
xnor U12752 (N_12752,N_11187,N_11182);
xor U12753 (N_12753,N_9953,N_10735);
or U12754 (N_12754,N_10117,N_11040);
xnor U12755 (N_12755,N_9439,N_9872);
nor U12756 (N_12756,N_10271,N_12037);
or U12757 (N_12757,N_12462,N_11361);
nor U12758 (N_12758,N_12301,N_10689);
or U12759 (N_12759,N_9524,N_11960);
and U12760 (N_12760,N_10136,N_9435);
and U12761 (N_12761,N_9744,N_11082);
xnor U12762 (N_12762,N_12145,N_11797);
xor U12763 (N_12763,N_9611,N_11515);
or U12764 (N_12764,N_10126,N_11244);
xnor U12765 (N_12765,N_11472,N_9479);
xnor U12766 (N_12766,N_11292,N_11209);
xor U12767 (N_12767,N_10127,N_10862);
nor U12768 (N_12768,N_11254,N_11581);
nor U12769 (N_12769,N_12367,N_9813);
and U12770 (N_12770,N_10717,N_10286);
nor U12771 (N_12771,N_11469,N_9945);
and U12772 (N_12772,N_10659,N_11013);
and U12773 (N_12773,N_12381,N_11078);
or U12774 (N_12774,N_12335,N_11646);
and U12775 (N_12775,N_10758,N_12098);
nand U12776 (N_12776,N_10638,N_10719);
and U12777 (N_12777,N_10852,N_11401);
nor U12778 (N_12778,N_11928,N_9661);
nor U12779 (N_12779,N_11389,N_9972);
nor U12780 (N_12780,N_10212,N_10245);
nand U12781 (N_12781,N_11195,N_10377);
nor U12782 (N_12782,N_9963,N_11003);
xnor U12783 (N_12783,N_9478,N_9683);
and U12784 (N_12784,N_11689,N_10263);
nor U12785 (N_12785,N_12230,N_10913);
or U12786 (N_12786,N_10973,N_11423);
nand U12787 (N_12787,N_10977,N_12202);
and U12788 (N_12788,N_12444,N_9475);
or U12789 (N_12789,N_12487,N_9864);
or U12790 (N_12790,N_10770,N_12382);
and U12791 (N_12791,N_10338,N_9687);
xor U12792 (N_12792,N_12333,N_12353);
nand U12793 (N_12793,N_9675,N_11568);
or U12794 (N_12794,N_9995,N_10131);
nand U12795 (N_12795,N_10511,N_11931);
or U12796 (N_12796,N_11543,N_10297);
and U12797 (N_12797,N_12378,N_9630);
and U12798 (N_12798,N_12292,N_9633);
nand U12799 (N_12799,N_11402,N_12326);
nor U12800 (N_12800,N_11784,N_9948);
or U12801 (N_12801,N_12002,N_9663);
or U12802 (N_12802,N_11540,N_11751);
nor U12803 (N_12803,N_12412,N_10435);
or U12804 (N_12804,N_12465,N_12275);
xor U12805 (N_12805,N_12170,N_9619);
nor U12806 (N_12806,N_12178,N_10564);
xor U12807 (N_12807,N_9385,N_11690);
xnor U12808 (N_12808,N_10474,N_12309);
xnor U12809 (N_12809,N_11502,N_12087);
nand U12810 (N_12810,N_11713,N_12299);
nor U12811 (N_12811,N_11156,N_9766);
nand U12812 (N_12812,N_10156,N_9666);
xnor U12813 (N_12813,N_11756,N_9588);
nor U12814 (N_12814,N_10330,N_11110);
nand U12815 (N_12815,N_11548,N_9971);
nand U12816 (N_12816,N_9853,N_10240);
nand U12817 (N_12817,N_10553,N_9855);
nor U12818 (N_12818,N_11442,N_10561);
or U12819 (N_12819,N_10076,N_9551);
and U12820 (N_12820,N_12235,N_11851);
nand U12821 (N_12821,N_10186,N_11103);
xnor U12822 (N_12822,N_12216,N_11027);
or U12823 (N_12823,N_11737,N_11698);
xor U12824 (N_12824,N_11664,N_9525);
nor U12825 (N_12825,N_12163,N_11258);
nand U12826 (N_12826,N_11984,N_10024);
nand U12827 (N_12827,N_12408,N_11070);
or U12828 (N_12828,N_11780,N_9987);
or U12829 (N_12829,N_11686,N_12269);
nor U12830 (N_12830,N_11020,N_12128);
nor U12831 (N_12831,N_10631,N_10145);
and U12832 (N_12832,N_9502,N_9990);
or U12833 (N_12833,N_11132,N_12016);
and U12834 (N_12834,N_11913,N_11871);
xor U12835 (N_12835,N_11314,N_12007);
nor U12836 (N_12836,N_10696,N_9993);
nor U12837 (N_12837,N_10075,N_10362);
nand U12838 (N_12838,N_10494,N_12236);
or U12839 (N_12839,N_11447,N_10342);
and U12840 (N_12840,N_11273,N_11095);
nor U12841 (N_12841,N_10621,N_12046);
nand U12842 (N_12842,N_11477,N_10507);
and U12843 (N_12843,N_10277,N_10622);
xnor U12844 (N_12844,N_11590,N_10836);
and U12845 (N_12845,N_11899,N_11585);
or U12846 (N_12846,N_11918,N_12416);
or U12847 (N_12847,N_11667,N_11714);
and U12848 (N_12848,N_10008,N_11942);
nor U12849 (N_12849,N_11280,N_9726);
and U12850 (N_12850,N_11635,N_10742);
nand U12851 (N_12851,N_10989,N_10028);
nand U12852 (N_12852,N_9559,N_11320);
xnor U12853 (N_12853,N_12241,N_9592);
or U12854 (N_12854,N_10050,N_11198);
nand U12855 (N_12855,N_11143,N_9597);
nand U12856 (N_12856,N_11079,N_10595);
xor U12857 (N_12857,N_12008,N_9936);
xor U12858 (N_12858,N_9561,N_10230);
and U12859 (N_12859,N_9737,N_9829);
or U12860 (N_12860,N_10214,N_10726);
nand U12861 (N_12861,N_10608,N_9646);
and U12862 (N_12862,N_12174,N_11675);
and U12863 (N_12863,N_12078,N_10666);
and U12864 (N_12864,N_9822,N_9549);
xor U12865 (N_12865,N_11236,N_10146);
nand U12866 (N_12866,N_10598,N_12000);
nand U12867 (N_12867,N_10976,N_12296);
or U12868 (N_12868,N_11777,N_11322);
nor U12869 (N_12869,N_12480,N_11775);
and U12870 (N_12870,N_10997,N_10283);
nand U12871 (N_12871,N_9421,N_9514);
or U12872 (N_12872,N_10267,N_11295);
nand U12873 (N_12873,N_10995,N_11677);
xnor U12874 (N_12874,N_12430,N_10259);
nor U12875 (N_12875,N_11507,N_12358);
or U12876 (N_12876,N_10961,N_12147);
nor U12877 (N_12877,N_11199,N_11140);
nor U12878 (N_12878,N_10442,N_12428);
xnor U12879 (N_12879,N_10014,N_10106);
nor U12880 (N_12880,N_12031,N_10821);
and U12881 (N_12881,N_9916,N_12394);
nand U12882 (N_12882,N_10496,N_10482);
and U12883 (N_12883,N_11532,N_11067);
xor U12884 (N_12884,N_9647,N_11241);
xor U12885 (N_12885,N_12448,N_10883);
or U12886 (N_12886,N_9693,N_11167);
and U12887 (N_12887,N_9574,N_10225);
or U12888 (N_12888,N_10047,N_10202);
or U12889 (N_12889,N_10902,N_10694);
xor U12890 (N_12890,N_9454,N_10011);
nor U12891 (N_12891,N_9529,N_10800);
and U12892 (N_12892,N_10470,N_10868);
xnor U12893 (N_12893,N_9839,N_9477);
and U12894 (N_12894,N_9622,N_10715);
xor U12895 (N_12895,N_9967,N_11856);
and U12896 (N_12896,N_11375,N_11782);
and U12897 (N_12897,N_9881,N_11623);
or U12898 (N_12898,N_12252,N_11988);
and U12899 (N_12899,N_9521,N_9897);
or U12900 (N_12900,N_11888,N_10617);
and U12901 (N_12901,N_10405,N_11211);
nand U12902 (N_12902,N_10266,N_11086);
and U12903 (N_12903,N_12063,N_9912);
and U12904 (N_12904,N_11606,N_10544);
xor U12905 (N_12905,N_12318,N_11098);
nand U12906 (N_12906,N_9991,N_12483);
xor U12907 (N_12907,N_9441,N_10796);
nand U12908 (N_12908,N_9444,N_10122);
and U12909 (N_12909,N_11042,N_9586);
or U12910 (N_12910,N_9748,N_11966);
or U12911 (N_12911,N_9562,N_11446);
xor U12912 (N_12912,N_11749,N_11374);
xnor U12913 (N_12913,N_12005,N_10927);
or U12914 (N_12914,N_12440,N_11123);
nor U12915 (N_12915,N_9484,N_11135);
nand U12916 (N_12916,N_10788,N_10998);
nand U12917 (N_12917,N_11761,N_12468);
nand U12918 (N_12918,N_10036,N_11947);
xnor U12919 (N_12919,N_12234,N_9835);
nor U12920 (N_12920,N_12240,N_11655);
nor U12921 (N_12921,N_10781,N_11492);
and U12922 (N_12922,N_11473,N_10224);
nor U12923 (N_12923,N_9777,N_10385);
or U12924 (N_12924,N_11838,N_9456);
nor U12925 (N_12925,N_10298,N_11961);
or U12926 (N_12926,N_9901,N_11146);
nand U12927 (N_12927,N_10092,N_11330);
or U12928 (N_12928,N_9805,N_10921);
or U12929 (N_12929,N_12066,N_9453);
and U12930 (N_12930,N_11805,N_11671);
nor U12931 (N_12931,N_10599,N_9790);
and U12932 (N_12932,N_12385,N_9398);
nor U12933 (N_12933,N_10447,N_10197);
xor U12934 (N_12934,N_10134,N_12404);
and U12935 (N_12935,N_9449,N_12276);
or U12936 (N_12936,N_10504,N_9674);
or U12937 (N_12937,N_12295,N_11719);
xnor U12938 (N_12938,N_9861,N_10062);
or U12939 (N_12939,N_11924,N_12110);
or U12940 (N_12940,N_11133,N_12157);
and U12941 (N_12941,N_11660,N_9670);
or U12942 (N_12942,N_11811,N_11818);
xor U12943 (N_12943,N_11068,N_11651);
nor U12944 (N_12944,N_9690,N_12205);
nor U12945 (N_12945,N_10284,N_9942);
nor U12946 (N_12946,N_9715,N_10819);
or U12947 (N_12947,N_12150,N_9801);
nand U12948 (N_12948,N_11362,N_9389);
or U12949 (N_12949,N_10587,N_11367);
nor U12950 (N_12950,N_11513,N_10256);
and U12951 (N_12951,N_11695,N_12167);
nand U12952 (N_12952,N_11650,N_12264);
nor U12953 (N_12953,N_10970,N_12197);
or U12954 (N_12954,N_10386,N_11154);
or U12955 (N_12955,N_10484,N_11812);
or U12956 (N_12956,N_12442,N_10443);
nor U12957 (N_12957,N_9934,N_10006);
nand U12958 (N_12958,N_11410,N_9745);
nor U12959 (N_12959,N_10841,N_12410);
xor U12960 (N_12960,N_10449,N_12001);
or U12961 (N_12961,N_9624,N_11077);
or U12962 (N_12962,N_10803,N_10493);
nand U12963 (N_12963,N_12413,N_9572);
and U12964 (N_12964,N_10974,N_10693);
nor U12965 (N_12965,N_10349,N_10346);
nand U12966 (N_12966,N_12390,N_10510);
or U12967 (N_12967,N_11748,N_10759);
nand U12968 (N_12968,N_10938,N_10276);
xor U12969 (N_12969,N_12036,N_12498);
and U12970 (N_12970,N_10328,N_10356);
xor U12971 (N_12971,N_11456,N_9962);
or U12972 (N_12972,N_9541,N_11288);
nor U12973 (N_12973,N_9605,N_12214);
xor U12974 (N_12974,N_11626,N_10205);
or U12975 (N_12975,N_11004,N_12114);
nand U12976 (N_12976,N_10196,N_10665);
xor U12977 (N_12977,N_12175,N_11864);
nand U12978 (N_12978,N_12485,N_12401);
and U12979 (N_12979,N_9686,N_9560);
and U12980 (N_12980,N_12363,N_11304);
nand U12981 (N_12981,N_12415,N_12307);
nor U12982 (N_12982,N_10573,N_11396);
xnor U12983 (N_12983,N_11256,N_11136);
xnor U12984 (N_12984,N_12120,N_9582);
xor U12985 (N_12985,N_12186,N_11552);
and U12986 (N_12986,N_11767,N_9640);
xor U12987 (N_12987,N_10589,N_11817);
nor U12988 (N_12988,N_12226,N_11064);
and U12989 (N_12989,N_9457,N_11219);
and U12990 (N_12990,N_9567,N_12291);
xnor U12991 (N_12991,N_10914,N_11604);
or U12992 (N_12992,N_10525,N_11841);
nand U12993 (N_12993,N_10591,N_10581);
and U12994 (N_12994,N_11745,N_12268);
or U12995 (N_12995,N_10116,N_11339);
or U12996 (N_12996,N_9915,N_11845);
or U12997 (N_12997,N_10857,N_12041);
nand U12998 (N_12998,N_10607,N_11326);
and U12999 (N_12999,N_11693,N_12284);
nor U13000 (N_13000,N_11559,N_10441);
nor U13001 (N_13001,N_9825,N_11332);
or U13002 (N_13002,N_9617,N_12259);
xor U13003 (N_13003,N_11302,N_11470);
and U13004 (N_13004,N_11225,N_12289);
nor U13005 (N_13005,N_11437,N_11514);
xor U13006 (N_13006,N_9889,N_11990);
nand U13007 (N_13007,N_10884,N_11257);
xor U13008 (N_13008,N_9416,N_11993);
or U13009 (N_13009,N_11450,N_9639);
xor U13010 (N_13010,N_11349,N_12190);
nand U13011 (N_13011,N_11778,N_9890);
nor U13012 (N_13012,N_10567,N_10261);
xnor U13013 (N_13013,N_10956,N_9576);
and U13014 (N_13014,N_12053,N_10155);
nand U13015 (N_13015,N_9706,N_11245);
nand U13016 (N_13016,N_11412,N_11467);
nor U13017 (N_13017,N_9824,N_10392);
nor U13018 (N_13018,N_11712,N_9699);
nand U13019 (N_13019,N_11279,N_9999);
and U13020 (N_13020,N_12361,N_9873);
and U13021 (N_13021,N_9637,N_12166);
or U13022 (N_13022,N_11922,N_10168);
nand U13023 (N_13023,N_9875,N_10020);
nand U13024 (N_13024,N_9844,N_9499);
or U13025 (N_13025,N_11594,N_11049);
nand U13026 (N_13026,N_12351,N_10031);
or U13027 (N_13027,N_12451,N_9390);
or U13028 (N_13028,N_11563,N_11935);
xor U13029 (N_13029,N_11312,N_9969);
nor U13030 (N_13030,N_11896,N_11863);
or U13031 (N_13031,N_11336,N_9550);
nand U13032 (N_13032,N_11071,N_11270);
nor U13033 (N_13033,N_10124,N_10711);
and U13034 (N_13034,N_10539,N_10918);
nor U13035 (N_13035,N_10506,N_10299);
nor U13036 (N_13036,N_9468,N_11474);
nor U13037 (N_13037,N_11956,N_10722);
nand U13038 (N_13038,N_12389,N_11353);
nor U13039 (N_13039,N_11125,N_10354);
nor U13040 (N_13040,N_9733,N_10213);
nor U13041 (N_13041,N_10204,N_9392);
and U13042 (N_13042,N_10262,N_12118);
xor U13043 (N_13043,N_10660,N_10555);
nand U13044 (N_13044,N_10644,N_10822);
xor U13045 (N_13045,N_10584,N_11461);
nand U13046 (N_13046,N_10648,N_11011);
or U13047 (N_13047,N_10130,N_10431);
or U13048 (N_13048,N_10791,N_12210);
xnor U13049 (N_13049,N_12435,N_10853);
xnor U13050 (N_13050,N_11866,N_12339);
or U13051 (N_13051,N_11321,N_10012);
xor U13052 (N_13052,N_10908,N_10325);
nor U13053 (N_13053,N_9717,N_9540);
or U13054 (N_13054,N_10228,N_10560);
or U13055 (N_13055,N_12429,N_11074);
nor U13056 (N_13056,N_10545,N_11334);
nor U13057 (N_13057,N_11720,N_9544);
nor U13058 (N_13058,N_10118,N_12274);
or U13059 (N_13059,N_11308,N_9768);
nand U13060 (N_13060,N_12198,N_11669);
nand U13061 (N_13061,N_11325,N_10672);
nor U13062 (N_13062,N_10396,N_11432);
and U13063 (N_13063,N_10152,N_11700);
and U13064 (N_13064,N_12481,N_10253);
xnor U13065 (N_13065,N_11129,N_9627);
nand U13066 (N_13066,N_11764,N_11728);
nand U13067 (N_13067,N_10922,N_10982);
nand U13068 (N_13068,N_12466,N_12425);
and U13069 (N_13069,N_9655,N_12312);
nor U13070 (N_13070,N_12074,N_10268);
and U13071 (N_13071,N_9570,N_10855);
and U13072 (N_13072,N_11708,N_10139);
nand U13073 (N_13073,N_11868,N_11518);
nor U13074 (N_13074,N_11030,N_10777);
or U13075 (N_13075,N_12158,N_10143);
and U13076 (N_13076,N_11260,N_9784);
xnor U13077 (N_13077,N_9727,N_11458);
xor U13078 (N_13078,N_10485,N_9752);
or U13079 (N_13079,N_10252,N_10623);
or U13080 (N_13080,N_11796,N_10761);
nor U13081 (N_13081,N_12194,N_11735);
or U13082 (N_13082,N_10352,N_10035);
xnor U13083 (N_13083,N_10779,N_11466);
xor U13084 (N_13084,N_10572,N_10900);
nand U13085 (N_13085,N_10872,N_10353);
xor U13086 (N_13086,N_10647,N_10335);
nand U13087 (N_13087,N_11937,N_12149);
or U13088 (N_13088,N_11705,N_11799);
or U13089 (N_13089,N_9534,N_9408);
or U13090 (N_13090,N_10958,N_9575);
nand U13091 (N_13091,N_11012,N_10307);
or U13092 (N_13092,N_12490,N_11509);
nand U13093 (N_13093,N_12438,N_11807);
xnor U13094 (N_13094,N_10071,N_11372);
and U13095 (N_13095,N_10658,N_11627);
nor U13096 (N_13096,N_9788,N_11893);
nand U13097 (N_13097,N_9914,N_11141);
nor U13098 (N_13098,N_9555,N_11085);
and U13099 (N_13099,N_12475,N_10331);
xnor U13100 (N_13100,N_9657,N_10910);
nand U13101 (N_13101,N_10153,N_12489);
nand U13102 (N_13102,N_11152,N_12423);
and U13103 (N_13103,N_11151,N_10321);
xor U13104 (N_13104,N_12137,N_10280);
nand U13105 (N_13105,N_11985,N_10601);
and U13106 (N_13106,N_11535,N_10091);
xnor U13107 (N_13107,N_11045,N_10532);
and U13108 (N_13108,N_10871,N_11373);
xnor U13109 (N_13109,N_9983,N_12320);
nand U13110 (N_13110,N_12187,N_10847);
or U13111 (N_13111,N_9974,N_11621);
nor U13112 (N_13112,N_11877,N_9469);
or U13113 (N_13113,N_9910,N_11358);
nor U13114 (N_13114,N_11122,N_9976);
nand U13115 (N_13115,N_12061,N_9425);
xnor U13116 (N_13116,N_11852,N_10189);
nand U13117 (N_13117,N_9986,N_9849);
nand U13118 (N_13118,N_10234,N_11859);
nor U13119 (N_13119,N_9489,N_9770);
or U13120 (N_13120,N_12419,N_10243);
nor U13121 (N_13121,N_10626,N_12045);
or U13122 (N_13122,N_10830,N_11592);
nand U13123 (N_13123,N_12079,N_11413);
nand U13124 (N_13124,N_9973,N_9711);
nor U13125 (N_13125,N_10678,N_12231);
and U13126 (N_13126,N_9838,N_11006);
xor U13127 (N_13127,N_9471,N_10515);
nor U13128 (N_13128,N_9517,N_11038);
nor U13129 (N_13129,N_11998,N_11923);
or U13130 (N_13130,N_11221,N_10905);
nor U13131 (N_13131,N_10060,N_11523);
nand U13132 (N_13132,N_10988,N_11521);
nand U13133 (N_13133,N_11331,N_10882);
and U13134 (N_13134,N_10099,N_10073);
or U13135 (N_13135,N_10490,N_9763);
xnor U13136 (N_13136,N_11584,N_11019);
or U13137 (N_13137,N_10557,N_11773);
nor U13138 (N_13138,N_10934,N_9789);
and U13139 (N_13139,N_9857,N_11275);
nand U13140 (N_13140,N_10825,N_9759);
nand U13141 (N_13141,N_12283,N_10824);
and U13142 (N_13142,N_9970,N_10025);
xor U13143 (N_13143,N_9831,N_9382);
and U13144 (N_13144,N_11255,N_9520);
nand U13145 (N_13145,N_9381,N_10953);
xnor U13146 (N_13146,N_11232,N_10404);
or U13147 (N_13147,N_10072,N_9654);
and U13148 (N_13148,N_10296,N_10070);
nor U13149 (N_13149,N_12086,N_9631);
and U13150 (N_13150,N_10558,N_10856);
xor U13151 (N_13151,N_11113,N_11861);
nand U13152 (N_13152,N_12103,N_10308);
nor U13153 (N_13153,N_9985,N_11164);
and U13154 (N_13154,N_12035,N_9671);
xnor U13155 (N_13155,N_11430,N_12138);
xnor U13156 (N_13156,N_11420,N_9565);
xnor U13157 (N_13157,N_11704,N_11000);
and U13158 (N_13158,N_9753,N_9742);
xor U13159 (N_13159,N_11822,N_9739);
xor U13160 (N_13160,N_9429,N_12025);
or U13161 (N_13161,N_12271,N_10258);
nor U13162 (N_13162,N_11645,N_11551);
xor U13163 (N_13163,N_9941,N_11607);
nand U13164 (N_13164,N_11043,N_10878);
or U13165 (N_13165,N_12315,N_9659);
xor U13166 (N_13166,N_10429,N_11790);
and U13167 (N_13167,N_10051,N_10656);
xor U13168 (N_13168,N_9830,N_12010);
xnor U13169 (N_13169,N_10219,N_10201);
nand U13170 (N_13170,N_11916,N_12492);
or U13171 (N_13171,N_11048,N_10344);
and U13172 (N_13172,N_9751,N_10450);
and U13173 (N_13173,N_12101,N_9388);
nand U13174 (N_13174,N_10109,N_10095);
or U13175 (N_13175,N_11031,N_11274);
xor U13176 (N_13176,N_10842,N_9649);
or U13177 (N_13177,N_12244,N_9643);
nand U13178 (N_13178,N_11005,N_10590);
nor U13179 (N_13179,N_10461,N_9573);
nor U13180 (N_13180,N_12135,N_9472);
nand U13181 (N_13181,N_10038,N_11854);
xnor U13182 (N_13182,N_10366,N_11282);
or U13183 (N_13183,N_12127,N_11920);
nand U13184 (N_13184,N_10210,N_12059);
nor U13185 (N_13185,N_12212,N_11462);
or U13186 (N_13186,N_11786,N_12267);
and U13187 (N_13187,N_9721,N_12417);
xnor U13188 (N_13188,N_12215,N_9564);
nand U13189 (N_13189,N_11820,N_9709);
or U13190 (N_13190,N_11609,N_10964);
nor U13191 (N_13191,N_11371,N_10087);
xnor U13192 (N_13192,N_9651,N_10293);
or U13193 (N_13193,N_10610,N_10200);
or U13194 (N_13194,N_12237,N_9417);
xor U13195 (N_13195,N_10901,N_12317);
nand U13196 (N_13196,N_10056,N_11526);
xnor U13197 (N_13197,N_11277,N_11999);
nand U13198 (N_13198,N_12133,N_10040);
nor U13199 (N_13199,N_12329,N_10787);
or U13200 (N_13200,N_9799,N_12290);
xnor U13201 (N_13201,N_9812,N_9827);
or U13202 (N_13202,N_11601,N_11188);
xor U13203 (N_13203,N_11853,N_9599);
nand U13204 (N_13204,N_11181,N_10949);
xor U13205 (N_13205,N_11685,N_11892);
and U13206 (N_13206,N_10054,N_11405);
or U13207 (N_13207,N_10249,N_9701);
and U13208 (N_13208,N_10509,N_9463);
nand U13209 (N_13209,N_10157,N_11204);
nor U13210 (N_13210,N_10114,N_10374);
xnor U13211 (N_13211,N_10078,N_10158);
and U13212 (N_13212,N_11290,N_12233);
or U13213 (N_13213,N_10115,N_10399);
nor U13214 (N_13214,N_11865,N_9584);
and U13215 (N_13215,N_9607,N_11015);
and U13216 (N_13216,N_12464,N_10533);
xor U13217 (N_13217,N_10414,N_11742);
or U13218 (N_13218,N_10701,N_12421);
and U13219 (N_13219,N_9394,N_10172);
nand U13220 (N_13220,N_12109,N_10520);
nor U13221 (N_13221,N_12321,N_10327);
nor U13222 (N_13222,N_10833,N_11229);
nand U13223 (N_13223,N_10473,N_10305);
nor U13224 (N_13224,N_10753,N_12471);
nor U13225 (N_13225,N_11951,N_10906);
nand U13226 (N_13226,N_10823,N_9923);
and U13227 (N_13227,N_9493,N_10103);
nand U13228 (N_13228,N_11528,N_9899);
nand U13229 (N_13229,N_12396,N_11495);
xor U13230 (N_13230,N_9403,N_11252);
or U13231 (N_13231,N_9518,N_10110);
nand U13232 (N_13232,N_10427,N_10345);
or U13233 (N_13233,N_9380,N_10052);
nor U13234 (N_13234,N_10026,N_10691);
xor U13235 (N_13235,N_11202,N_11400);
and U13236 (N_13236,N_11953,N_11633);
and U13237 (N_13237,N_10419,N_10946);
and U13238 (N_13238,N_9689,N_11972);
nor U13239 (N_13239,N_9743,N_9988);
xnor U13240 (N_13240,N_10236,N_12343);
or U13241 (N_13241,N_10864,N_10827);
nor U13242 (N_13242,N_10161,N_11666);
or U13243 (N_13243,N_12255,N_10413);
nand U13244 (N_13244,N_11519,N_11520);
nor U13245 (N_13245,N_11837,N_12020);
nor U13246 (N_13246,N_11542,N_9756);
xnor U13247 (N_13247,N_9538,N_10865);
nand U13248 (N_13248,N_10776,N_11776);
nand U13249 (N_13249,N_12325,N_10606);
nand U13250 (N_13250,N_11955,N_11907);
xnor U13251 (N_13251,N_11588,N_10066);
or U13252 (N_13252,N_11886,N_11222);
xor U13253 (N_13253,N_11798,N_12131);
or U13254 (N_13254,N_9714,N_10549);
and U13255 (N_13255,N_12232,N_11586);
nor U13256 (N_13256,N_12113,N_10732);
xor U13257 (N_13257,N_12450,N_11001);
and U13258 (N_13258,N_10994,N_12200);
or U13259 (N_13259,N_11338,N_10843);
and U13260 (N_13260,N_11307,N_9785);
nor U13261 (N_13261,N_11393,N_10979);
and U13262 (N_13262,N_10614,N_9375);
or U13263 (N_13263,N_10164,N_10720);
nor U13264 (N_13264,N_10001,N_11978);
xnor U13265 (N_13265,N_11183,N_11459);
nand U13266 (N_13266,N_9966,N_10090);
xnor U13267 (N_13267,N_10579,N_10445);
nand U13268 (N_13268,N_11429,N_11380);
xnor U13269 (N_13269,N_12033,N_11227);
nor U13270 (N_13270,N_11653,N_10764);
nor U13271 (N_13271,N_9841,N_11827);
or U13272 (N_13272,N_9823,N_12452);
xor U13273 (N_13273,N_11624,N_11180);
or U13274 (N_13274,N_11957,N_12051);
or U13275 (N_13275,N_11878,N_12314);
and U13276 (N_13276,N_12199,N_9673);
nor U13277 (N_13277,N_11050,N_11200);
or U13278 (N_13278,N_10806,N_11766);
and U13279 (N_13279,N_9797,N_10048);
and U13280 (N_13280,N_10569,N_11755);
and U13281 (N_13281,N_12324,N_10752);
xor U13282 (N_13282,N_12141,N_10053);
nor U13283 (N_13283,N_12311,N_11870);
xor U13284 (N_13284,N_12261,N_11557);
nand U13285 (N_13285,N_12023,N_10257);
and U13286 (N_13286,N_10870,N_12391);
xnor U13287 (N_13287,N_10387,N_9826);
nand U13288 (N_13288,N_10812,N_11908);
xor U13289 (N_13289,N_9862,N_10481);
nor U13290 (N_13290,N_12297,N_12482);
nand U13291 (N_13291,N_11281,N_11328);
xor U13292 (N_13292,N_11630,N_10578);
xor U13293 (N_13293,N_10169,N_9809);
and U13294 (N_13294,N_11982,N_10772);
nand U13295 (N_13295,N_11486,N_11710);
xor U13296 (N_13296,N_11214,N_12347);
nor U13297 (N_13297,N_11503,N_9918);
xnor U13298 (N_13298,N_11855,N_9926);
and U13299 (N_13299,N_11846,N_9641);
nor U13300 (N_13300,N_9780,N_11938);
or U13301 (N_13301,N_11169,N_11632);
or U13302 (N_13302,N_12092,N_10393);
nand U13303 (N_13303,N_11327,N_11538);
nor U13304 (N_13304,N_12287,N_10055);
nor U13305 (N_13305,N_9907,N_11084);
nand U13306 (N_13306,N_9888,N_10173);
nor U13307 (N_13307,N_10671,N_11810);
nand U13308 (N_13308,N_9626,N_11099);
nor U13309 (N_13309,N_9867,N_11106);
nor U13310 (N_13310,N_11341,N_10932);
xnor U13311 (N_13311,N_12014,N_11016);
or U13312 (N_13312,N_12486,N_11407);
nand U13313 (N_13313,N_10554,N_11271);
and U13314 (N_13314,N_10512,N_9905);
or U13315 (N_13315,N_12062,N_12310);
or U13316 (N_13316,N_10336,N_9779);
nor U13317 (N_13317,N_12243,N_11301);
and U13318 (N_13318,N_11148,N_12497);
and U13319 (N_13319,N_11230,N_11849);
and U13320 (N_13320,N_9532,N_10627);
nand U13321 (N_13321,N_11491,N_11137);
or U13322 (N_13322,N_11560,N_10415);
and U13323 (N_13323,N_12460,N_12411);
or U13324 (N_13324,N_12433,N_9604);
xor U13325 (N_13325,N_9997,N_9378);
nor U13326 (N_13326,N_9754,N_11697);
xnor U13327 (N_13327,N_10840,N_12047);
or U13328 (N_13328,N_11364,N_11828);
xnor U13329 (N_13329,N_10754,N_10687);
nor U13330 (N_13330,N_11975,N_10651);
nand U13331 (N_13331,N_11561,N_11286);
and U13332 (N_13332,N_11212,N_10642);
and U13333 (N_13333,N_11309,N_11479);
and U13334 (N_13334,N_9856,N_10250);
or U13335 (N_13335,N_12136,N_11263);
nand U13336 (N_13336,N_9509,N_12072);
or U13337 (N_13337,N_11674,N_9707);
nand U13338 (N_13338,N_9482,N_10316);
xnor U13339 (N_13339,N_11269,N_11112);
xor U13340 (N_13340,N_9685,N_10834);
xnor U13341 (N_13341,N_10067,N_9928);
nand U13342 (N_13342,N_12239,N_9832);
xnor U13343 (N_13343,N_12015,N_10990);
and U13344 (N_13344,N_11435,N_9736);
and U13345 (N_13345,N_11382,N_10104);
xor U13346 (N_13346,N_12091,N_11652);
xor U13347 (N_13347,N_9740,N_11730);
nor U13348 (N_13348,N_9874,N_10962);
nand U13349 (N_13349,N_11408,N_9723);
nor U13350 (N_13350,N_10129,N_11489);
nand U13351 (N_13351,N_11162,N_10275);
and U13352 (N_13352,N_10688,N_10680);
xor U13353 (N_13353,N_11419,N_10538);
or U13354 (N_13354,N_12388,N_10928);
and U13355 (N_13355,N_12213,N_10987);
and U13356 (N_13356,N_9548,N_9587);
nor U13357 (N_13357,N_10709,N_9868);
nor U13358 (N_13358,N_9846,N_10102);
or U13359 (N_13359,N_9466,N_9906);
nor U13360 (N_13360,N_10813,N_10416);
and U13361 (N_13361,N_12184,N_9946);
and U13362 (N_13362,N_10412,N_11583);
xor U13363 (N_13363,N_11351,N_10209);
and U13364 (N_13364,N_9430,N_11501);
nor U13365 (N_13365,N_11354,N_10467);
and U13366 (N_13366,N_11945,N_11059);
nand U13367 (N_13367,N_11324,N_11468);
nand U13368 (N_13368,N_11567,N_11457);
and U13369 (N_13369,N_12300,N_12455);
nand U13370 (N_13370,N_11220,N_10681);
nor U13371 (N_13371,N_11634,N_10452);
nor U13372 (N_13372,N_10543,N_11598);
nand U13373 (N_13373,N_9557,N_10269);
xor U13374 (N_13374,N_10233,N_10981);
nand U13375 (N_13375,N_12403,N_11832);
nor U13376 (N_13376,N_11008,N_9512);
and U13377 (N_13377,N_10966,N_9578);
xor U13378 (N_13378,N_11278,N_11035);
nand U13379 (N_13379,N_10021,N_10242);
xnor U13380 (N_13380,N_12470,N_9870);
and U13381 (N_13381,N_9667,N_10725);
and U13382 (N_13382,N_11081,N_12345);
and U13383 (N_13383,N_10138,N_9925);
nand U13384 (N_13384,N_10641,N_10238);
xnor U13385 (N_13385,N_10513,N_12168);
and U13386 (N_13386,N_10534,N_12399);
or U13387 (N_13387,N_10655,N_12469);
nor U13388 (N_13388,N_9884,N_12349);
and U13389 (N_13389,N_12018,N_9814);
and U13390 (N_13390,N_11847,N_9917);
or U13391 (N_13391,N_10807,N_9505);
nor U13392 (N_13392,N_12152,N_12334);
nor U13393 (N_13393,N_10007,N_10814);
nor U13394 (N_13394,N_10529,N_10583);
and U13395 (N_13395,N_12246,N_11962);
or U13396 (N_13396,N_10967,N_11497);
xor U13397 (N_13397,N_10596,N_10888);
xor U13398 (N_13398,N_12090,N_10265);
or U13399 (N_13399,N_11860,N_12323);
xor U13400 (N_13400,N_11912,N_11897);
xnor U13401 (N_13401,N_11874,N_12383);
xor U13402 (N_13402,N_9871,N_9877);
nor U13403 (N_13403,N_11261,N_10378);
and U13404 (N_13404,N_10089,N_9526);
or U13405 (N_13405,N_12453,N_9650);
nor U13406 (N_13406,N_10585,N_10367);
nand U13407 (N_13407,N_12052,N_12083);
nand U13408 (N_13408,N_11692,N_10334);
or U13409 (N_13409,N_11089,N_10820);
and U13410 (N_13410,N_11149,N_10355);
nor U13411 (N_13411,N_12277,N_11512);
xnor U13412 (N_13412,N_11770,N_10023);
or U13413 (N_13413,N_11216,N_10611);
nor U13414 (N_13414,N_10371,N_11481);
nand U13415 (N_13415,N_10664,N_11037);
and U13416 (N_13416,N_10218,N_11318);
nor U13417 (N_13417,N_11582,N_10108);
or U13418 (N_13418,N_12049,N_11340);
xnor U13419 (N_13419,N_11734,N_10027);
and U13420 (N_13420,N_11053,N_12305);
xor U13421 (N_13421,N_12097,N_10952);
nand U13422 (N_13422,N_12148,N_10604);
and U13423 (N_13423,N_10923,N_10388);
and U13424 (N_13424,N_10837,N_10472);
and U13425 (N_13425,N_12165,N_11421);
nand U13426 (N_13426,N_10851,N_11347);
and U13427 (N_13427,N_11287,N_10887);
xnor U13428 (N_13428,N_9668,N_12405);
and U13429 (N_13429,N_9503,N_11163);
nand U13430 (N_13430,N_12164,N_11758);
or U13431 (N_13431,N_10756,N_10079);
and U13432 (N_13432,N_10180,N_10890);
xnor U13433 (N_13433,N_10808,N_11504);
or U13434 (N_13434,N_11390,N_11733);
and U13435 (N_13435,N_12374,N_11883);
nand U13436 (N_13436,N_9882,N_11439);
nand U13437 (N_13437,N_10592,N_9510);
nor U13438 (N_13438,N_10061,N_12293);
and U13439 (N_13439,N_12060,N_12108);
nand U13440 (N_13440,N_12393,N_9426);
nand U13441 (N_13441,N_12407,N_11010);
nand U13442 (N_13442,N_10113,N_10749);
nor U13443 (N_13443,N_10499,N_10925);
and U13444 (N_13444,N_11939,N_9718);
nor U13445 (N_13445,N_11482,N_11873);
or U13446 (N_13446,N_10712,N_12330);
and U13447 (N_13447,N_9880,N_10975);
nor U13448 (N_13448,N_10546,N_12126);
xor U13449 (N_13449,N_11803,N_9932);
nand U13450 (N_13450,N_11723,N_10502);
or U13451 (N_13451,N_11980,N_12116);
or U13452 (N_13452,N_11431,N_11783);
and U13453 (N_13453,N_11904,N_9490);
or U13454 (N_13454,N_10329,N_12426);
nor U13455 (N_13455,N_11903,N_9697);
nand U13456 (N_13456,N_11639,N_11572);
nor U13457 (N_13457,N_11794,N_10348);
or U13458 (N_13458,N_11591,N_12208);
nor U13459 (N_13459,N_9858,N_12395);
xor U13460 (N_13460,N_10310,N_9719);
and U13461 (N_13461,N_9608,N_9750);
nand U13462 (N_13462,N_9415,N_10562);
or U13463 (N_13463,N_12156,N_10528);
or U13464 (N_13464,N_9648,N_9978);
and U13465 (N_13465,N_10285,N_12245);
and U13466 (N_13466,N_9546,N_11426);
nor U13467 (N_13467,N_11142,N_9815);
and U13468 (N_13468,N_11422,N_12107);
or U13469 (N_13469,N_10241,N_11197);
nor U13470 (N_13470,N_12377,N_10747);
xnor U13471 (N_13471,N_11100,N_10710);
xnor U13472 (N_13472,N_11739,N_9695);
and U13473 (N_13473,N_12238,N_12461);
nand U13474 (N_13474,N_10315,N_10288);
xor U13475 (N_13475,N_11418,N_11611);
nor U13476 (N_13476,N_12386,N_11600);
or U13477 (N_13477,N_12253,N_9462);
nand U13478 (N_13478,N_10323,N_10690);
nand U13479 (N_13479,N_12332,N_11240);
or U13480 (N_13480,N_11580,N_10343);
nor U13481 (N_13481,N_11174,N_11296);
nand U13482 (N_13482,N_11046,N_11233);
nand U13483 (N_13483,N_9828,N_10369);
nor U13484 (N_13484,N_11259,N_12341);
xor U13485 (N_13485,N_9807,N_10478);
xnor U13486 (N_13486,N_12285,N_10526);
nor U13487 (N_13487,N_11944,N_9908);
nand U13488 (N_13488,N_11996,N_10034);
or U13489 (N_13489,N_12004,N_11208);
xor U13490 (N_13490,N_12319,N_12478);
nand U13491 (N_13491,N_9965,N_10700);
xor U13492 (N_13492,N_10521,N_9428);
or U13493 (N_13493,N_9865,N_10045);
xnor U13494 (N_13494,N_11835,N_10935);
or U13495 (N_13495,N_10603,N_11994);
xnor U13496 (N_13496,N_10797,N_10705);
nand U13497 (N_13497,N_9554,N_11092);
nand U13498 (N_13498,N_10193,N_12146);
and U13499 (N_13499,N_9811,N_10471);
xnor U13500 (N_13500,N_12398,N_10340);
xor U13501 (N_13501,N_10624,N_11815);
and U13502 (N_13502,N_10750,N_9944);
nor U13503 (N_13503,N_10565,N_10418);
nor U13504 (N_13504,N_9710,N_10858);
xnor U13505 (N_13505,N_11310,N_10333);
or U13506 (N_13506,N_11090,N_12256);
nand U13507 (N_13507,N_12474,N_10279);
and U13508 (N_13508,N_11620,N_10383);
nand U13509 (N_13509,N_11508,N_11130);
or U13510 (N_13510,N_12447,N_9423);
or U13511 (N_13511,N_10898,N_11109);
nand U13512 (N_13512,N_10636,N_11902);
nor U13513 (N_13513,N_9566,N_12364);
or U13514 (N_13514,N_9474,N_11663);
nand U13515 (N_13515,N_10432,N_10547);
and U13516 (N_13516,N_10916,N_11746);
xor U13517 (N_13517,N_10398,N_11406);
and U13518 (N_13518,N_11701,N_11145);
and U13519 (N_13519,N_12499,N_11885);
xor U13520 (N_13520,N_10826,N_9996);
nor U13521 (N_13521,N_10018,N_11754);
or U13522 (N_13522,N_9461,N_12075);
xor U13523 (N_13523,N_10875,N_11126);
or U13524 (N_13524,N_10945,N_10360);
xor U13525 (N_13525,N_10364,N_10406);
xnor U13526 (N_13526,N_9879,N_11768);
xor U13527 (N_13527,N_9539,N_10818);
or U13528 (N_13528,N_10832,N_12115);
nor U13529 (N_13529,N_11890,N_11589);
nor U13530 (N_13530,N_11740,N_9747);
nor U13531 (N_13531,N_11566,N_11168);
and U13532 (N_13532,N_11313,N_10379);
nand U13533 (N_13533,N_11603,N_9920);
xor U13534 (N_13534,N_12251,N_12057);
nor U13535 (N_13535,N_11242,N_9843);
nand U13536 (N_13536,N_11343,N_9749);
nand U13537 (N_13537,N_11483,N_11680);
and U13538 (N_13538,N_11759,N_11752);
xnor U13539 (N_13539,N_10167,N_11531);
nor U13540 (N_13540,N_10282,N_12132);
nand U13541 (N_13541,N_12344,N_11009);
nor U13542 (N_13542,N_10792,N_11022);
xor U13543 (N_13543,N_11072,N_11303);
nand U13544 (N_13544,N_10859,N_10391);
or U13545 (N_13545,N_10593,N_10574);
nand U13546 (N_13546,N_11023,N_9959);
nand U13547 (N_13547,N_11834,N_11887);
nor U13548 (N_13548,N_12153,N_10454);
or U13549 (N_13549,N_9850,N_11051);
nand U13550 (N_13550,N_9638,N_9732);
or U13551 (N_13551,N_10985,N_10049);
xnor U13552 (N_13552,N_11175,N_10542);
and U13553 (N_13553,N_12124,N_10003);
nand U13554 (N_13554,N_12130,N_12085);
nor U13555 (N_13555,N_11895,N_9724);
nand U13556 (N_13556,N_9728,N_12384);
and U13557 (N_13557,N_10708,N_11357);
or U13558 (N_13558,N_10456,N_10483);
or U13559 (N_13559,N_10105,N_11724);
nand U13560 (N_13560,N_9678,N_11317);
or U13561 (N_13561,N_11804,N_10786);
or U13562 (N_13562,N_9448,N_12355);
nand U13563 (N_13563,N_10084,N_11127);
nor U13564 (N_13564,N_11041,N_11725);
xor U13565 (N_13565,N_10746,N_12139);
xnor U13566 (N_13566,N_10673,N_11414);
and U13567 (N_13567,N_10183,N_9402);
or U13568 (N_13568,N_10451,N_11525);
nand U13569 (N_13569,N_11760,N_9577);
xor U13570 (N_13570,N_10675,N_9778);
or U13571 (N_13571,N_9927,N_11833);
nor U13572 (N_13572,N_12456,N_10886);
xnor U13573 (N_13573,N_10395,N_12076);
and U13574 (N_13574,N_10798,N_12142);
nand U13575 (N_13575,N_12272,N_10165);
nand U13576 (N_13576,N_10453,N_11744);
nand U13577 (N_13577,N_9705,N_10093);
and U13578 (N_13578,N_11750,N_12286);
and U13579 (N_13579,N_9613,N_10789);
or U13580 (N_13580,N_10760,N_9903);
xnor U13581 (N_13581,N_10954,N_11044);
and U13582 (N_13582,N_11101,N_12406);
nor U13583 (N_13583,N_10695,N_11602);
xor U13584 (N_13584,N_11398,N_10602);
xor U13585 (N_13585,N_9845,N_10941);
nor U13586 (N_13586,N_11436,N_12273);
nor U13587 (N_13587,N_9606,N_10175);
nand U13588 (N_13588,N_11463,N_12034);
nand U13589 (N_13589,N_9431,N_10306);
nor U13590 (N_13590,N_11662,N_10010);
and U13591 (N_13591,N_9603,N_10148);
and U13592 (N_13592,N_10185,N_10730);
nor U13593 (N_13593,N_10947,N_10120);
nor U13594 (N_13594,N_10931,N_9795);
xor U13595 (N_13595,N_12176,N_11736);
xor U13596 (N_13596,N_10519,N_12125);
nand U13597 (N_13597,N_9760,N_9896);
xnor U13598 (N_13598,N_10652,N_9537);
or U13599 (N_13599,N_9487,N_10703);
or U13600 (N_13600,N_11392,N_11595);
and U13601 (N_13601,N_11617,N_10068);
nor U13602 (N_13602,N_11153,N_10319);
nand U13603 (N_13603,N_11356,N_11656);
nand U13604 (N_13604,N_11105,N_11547);
nor U13605 (N_13605,N_10094,N_10479);
or U13606 (N_13606,N_10570,N_11108);
nor U13607 (N_13607,N_10577,N_10877);
xnor U13608 (N_13608,N_9452,N_11631);
xor U13609 (N_13609,N_11718,N_10215);
nand U13610 (N_13610,N_10444,N_10128);
or U13611 (N_13611,N_11826,N_10140);
nand U13612 (N_13612,N_10217,N_9774);
nand U13613 (N_13613,N_12459,N_11228);
and U13614 (N_13614,N_12117,N_10016);
xor U13615 (N_13615,N_11683,N_10920);
or U13616 (N_13616,N_11465,N_10248);
nor U13617 (N_13617,N_10420,N_11311);
nor U13618 (N_13618,N_11802,N_12446);
or U13619 (N_13619,N_9876,N_11409);
nor U13620 (N_13620,N_12099,N_12169);
and U13621 (N_13621,N_12302,N_11383);
and U13622 (N_13622,N_9556,N_12418);
nand U13623 (N_13623,N_11158,N_10436);
nor U13624 (N_13624,N_9500,N_10176);
nand U13625 (N_13625,N_9418,N_11654);
nor U13626 (N_13626,N_12143,N_11499);
or U13627 (N_13627,N_10790,N_10763);
nor U13628 (N_13628,N_11658,N_10848);
xor U13629 (N_13629,N_11500,N_11554);
nor U13630 (N_13630,N_11806,N_11210);
xnor U13631 (N_13631,N_9738,N_11065);
nor U13632 (N_13632,N_12054,N_10940);
xnor U13633 (N_13633,N_11544,N_11249);
nand U13634 (N_13634,N_11115,N_11964);
or U13635 (N_13635,N_10679,N_10375);
and U13636 (N_13636,N_12195,N_9767);
and U13637 (N_13637,N_11510,N_11889);
xnor U13638 (N_13638,N_10332,N_12434);
xor U13639 (N_13639,N_12019,N_10475);
and U13640 (N_13640,N_11411,N_12106);
nor U13641 (N_13641,N_10637,N_10300);
or U13642 (N_13642,N_9800,N_10854);
and U13643 (N_13643,N_11687,N_9922);
nor U13644 (N_13644,N_10039,N_9818);
nor U13645 (N_13645,N_11506,N_9786);
nand U13646 (N_13646,N_9465,N_11266);
and U13647 (N_13647,N_9773,N_9989);
nor U13648 (N_13648,N_10046,N_11173);
xnor U13649 (N_13649,N_12182,N_11831);
nand U13650 (N_13650,N_10096,N_10320);
or U13651 (N_13651,N_11391,N_11608);
and U13652 (N_13652,N_9645,N_11298);
xnor U13653 (N_13653,N_10264,N_11306);
and U13654 (N_13654,N_10222,N_11262);
xor U13655 (N_13655,N_10575,N_9672);
xor U13656 (N_13656,N_10963,N_11002);
nand U13657 (N_13657,N_11120,N_11124);
or U13658 (N_13658,N_12449,N_9581);
nand U13659 (N_13659,N_10950,N_9506);
nand U13660 (N_13660,N_10992,N_11404);
nor U13661 (N_13661,N_9594,N_11399);
and U13662 (N_13662,N_11929,N_10465);
xnor U13663 (N_13663,N_10540,N_11438);
nand U13664 (N_13664,N_12204,N_9782);
xor U13665 (N_13665,N_10795,N_9422);
nor U13666 (N_13666,N_12161,N_10771);
xor U13667 (N_13667,N_11118,N_10486);
or U13668 (N_13668,N_11342,N_9434);
and U13669 (N_13669,N_9451,N_10959);
xor U13670 (N_13670,N_10991,N_10382);
nor U13671 (N_13671,N_12370,N_10831);
and U13672 (N_13672,N_10121,N_11619);
and U13673 (N_13673,N_10488,N_12266);
and U13674 (N_13674,N_9440,N_11844);
nor U13675 (N_13675,N_9955,N_11370);
xor U13676 (N_13676,N_11424,N_10899);
nor U13677 (N_13677,N_10229,N_9542);
and U13678 (N_13678,N_9783,N_11747);
and U13679 (N_13679,N_9653,N_11840);
xnor U13680 (N_13680,N_9595,N_11062);
xnor U13681 (N_13681,N_11363,N_11034);
or U13682 (N_13682,N_10469,N_10667);
or U13683 (N_13683,N_10239,N_10677);
and U13684 (N_13684,N_12380,N_10983);
nor U13685 (N_13685,N_9943,N_11824);
xnor U13686 (N_13686,N_9580,N_11647);
nor U13687 (N_13687,N_9939,N_11007);
or U13688 (N_13688,N_12359,N_10287);
or U13689 (N_13689,N_10100,N_9866);
xor U13690 (N_13690,N_9464,N_10171);
and U13691 (N_13691,N_11178,N_9982);
nand U13692 (N_13692,N_11925,N_10107);
xnor U13693 (N_13693,N_11785,N_10497);
nand U13694 (N_13694,N_11891,N_10894);
xnor U13695 (N_13695,N_11524,N_12003);
nor U13696 (N_13696,N_10500,N_11771);
nand U13697 (N_13697,N_12093,N_10278);
and U13698 (N_13698,N_9937,N_9819);
and U13699 (N_13699,N_10805,N_11425);
or U13700 (N_13700,N_11821,N_11289);
and U13701 (N_13701,N_11036,N_9981);
nand U13702 (N_13702,N_12088,N_11536);
nand U13703 (N_13703,N_10188,N_11932);
nor U13704 (N_13704,N_11914,N_9902);
xor U13705 (N_13705,N_9447,N_9386);
and U13706 (N_13706,N_11348,N_11579);
nor U13707 (N_13707,N_11207,N_11573);
xnor U13708 (N_13708,N_9507,N_11179);
xnor U13709 (N_13709,N_11427,N_9703);
and U13710 (N_13710,N_10773,N_12392);
nand U13711 (N_13711,N_10083,N_12265);
nor U13712 (N_13712,N_10487,N_12248);
or U13713 (N_13713,N_11711,N_12476);
and U13714 (N_13714,N_10698,N_10394);
nand U13715 (N_13715,N_12228,N_9765);
xor U13716 (N_13716,N_11910,N_12121);
xnor U13717 (N_13717,N_11206,N_9522);
nand U13718 (N_13718,N_11026,N_9508);
nor U13719 (N_13719,N_9810,N_12494);
or U13720 (N_13720,N_11272,N_9694);
xnor U13721 (N_13721,N_10438,N_12134);
nand U13722 (N_13722,N_12218,N_11498);
nand U13723 (N_13723,N_10782,N_10181);
or U13724 (N_13724,N_12027,N_9620);
xnor U13725 (N_13725,N_11201,N_9895);
nor U13726 (N_13726,N_9391,N_11565);
or U13727 (N_13727,N_10476,N_12095);
or U13728 (N_13728,N_9602,N_9984);
xor U13729 (N_13729,N_11858,N_11974);
or U13730 (N_13730,N_11682,N_12422);
nand U13731 (N_13731,N_11555,N_12217);
xor U13732 (N_13732,N_11558,N_12040);
nand U13733 (N_13733,N_11848,N_11571);
or U13734 (N_13734,N_11478,N_9533);
xor U13735 (N_13735,N_11384,N_11839);
or U13736 (N_13736,N_10915,N_10430);
or U13737 (N_13737,N_9949,N_9535);
nor U13738 (N_13738,N_10421,N_9954);
nand U13739 (N_13739,N_9977,N_11379);
nand U13740 (N_13740,N_10850,N_9437);
nor U13741 (N_13741,N_12089,N_11300);
or U13742 (N_13742,N_9669,N_11665);
xor U13743 (N_13743,N_12193,N_11850);
and U13744 (N_13744,N_11192,N_10597);
or U13745 (N_13745,N_10192,N_11917);
and U13746 (N_13746,N_10211,N_11715);
and U13747 (N_13747,N_11823,N_10650);
and U13748 (N_13748,N_10743,N_10780);
xor U13749 (N_13749,N_10270,N_9395);
nor U13750 (N_13750,N_11881,N_10044);
nand U13751 (N_13751,N_10942,N_9545);
nor U13752 (N_13752,N_11448,N_9775);
nand U13753 (N_13753,N_9821,N_11147);
xnor U13754 (N_13754,N_9833,N_11789);
nand U13755 (N_13755,N_11104,N_9601);
nor U13756 (N_13756,N_11150,N_9960);
or U13757 (N_13757,N_11808,N_9629);
nor U13758 (N_13758,N_9400,N_11977);
or U13759 (N_13759,N_12488,N_9957);
and U13760 (N_13760,N_12250,N_9511);
xor U13761 (N_13761,N_10220,N_10874);
and U13762 (N_13762,N_11039,N_12258);
nand U13763 (N_13763,N_9771,N_10969);
xnor U13764 (N_13764,N_11661,N_12067);
and U13765 (N_13765,N_11612,N_10707);
xor U13766 (N_13766,N_10731,N_12206);
xnor U13767 (N_13767,N_11915,N_10002);
nand U13768 (N_13768,N_10654,N_10737);
nor U13769 (N_13769,N_12379,N_9938);
and U13770 (N_13770,N_10247,N_11792);
nor U13771 (N_13771,N_10738,N_12119);
nor U13772 (N_13772,N_9591,N_10294);
nand U13773 (N_13773,N_11250,N_12454);
nand U13774 (N_13774,N_11587,N_10580);
xnor U13775 (N_13775,N_10289,N_9929);
nor U13776 (N_13776,N_10069,N_9450);
and U13777 (N_13777,N_10762,N_10880);
and U13778 (N_13778,N_10433,N_10434);
nand U13779 (N_13779,N_10410,N_12050);
nand U13780 (N_13780,N_9691,N_11075);
nand U13781 (N_13781,N_9485,N_10615);
or U13782 (N_13782,N_10702,N_12472);
nor U13783 (N_13783,N_10568,N_9722);
or U13784 (N_13784,N_12342,N_11983);
nor U13785 (N_13785,N_10766,N_10322);
or U13786 (N_13786,N_10074,N_12260);
and U13787 (N_13787,N_11909,N_10618);
nand U13788 (N_13788,N_12123,N_11869);
nand U13789 (N_13789,N_10203,N_11189);
or U13790 (N_13790,N_11638,N_11649);
and U13791 (N_13791,N_11857,N_12006);
nand U13792 (N_13792,N_11455,N_12400);
nand U13793 (N_13793,N_10166,N_11246);
xor U13794 (N_13794,N_10802,N_12024);
nor U13795 (N_13795,N_12484,N_10699);
nor U13796 (N_13796,N_9427,N_12322);
xor U13797 (N_13797,N_10704,N_10801);
nand U13798 (N_13798,N_11539,N_12223);
xor U13799 (N_13799,N_9702,N_11787);
nand U13800 (N_13800,N_12211,N_12096);
nor U13801 (N_13801,N_12012,N_11172);
nor U13802 (N_13802,N_9527,N_10409);
and U13803 (N_13803,N_10463,N_10740);
nor U13804 (N_13804,N_10640,N_11315);
or U13805 (N_13805,N_11131,N_11516);
xor U13806 (N_13806,N_11268,N_10119);
and U13807 (N_13807,N_10401,N_11238);
and U13808 (N_13808,N_10536,N_10984);
nand U13809 (N_13809,N_11517,N_9494);
nor U13810 (N_13810,N_9696,N_11335);
and U13811 (N_13811,N_12100,N_11625);
and U13812 (N_13812,N_11176,N_9851);
xor U13813 (N_13813,N_9679,N_11668);
and U13814 (N_13814,N_9746,N_9660);
nand U13815 (N_13815,N_11160,N_10713);
xnor U13816 (N_13816,N_9904,N_9665);
xnor U13817 (N_13817,N_9404,N_11537);
nand U13818 (N_13818,N_10996,N_12278);
or U13819 (N_13819,N_12354,N_11657);
or U13820 (N_13820,N_9755,N_9625);
nand U13821 (N_13821,N_9569,N_11829);
or U13822 (N_13822,N_10676,N_9682);
xor U13823 (N_13823,N_11066,N_9553);
nand U13824 (N_13824,N_10838,N_12177);
and U13825 (N_13825,N_11511,N_11989);
and U13826 (N_13826,N_11265,N_11943);
or U13827 (N_13827,N_10849,N_11144);
nand U13828 (N_13828,N_12439,N_10634);
xor U13829 (N_13829,N_11741,N_10498);
and U13830 (N_13830,N_11900,N_12373);
or U13831 (N_13831,N_12183,N_12154);
nor U13832 (N_13832,N_10135,N_9476);
or U13833 (N_13833,N_11097,N_10142);
nor U13834 (N_13834,N_11460,N_11936);
and U13835 (N_13835,N_9644,N_10576);
nor U13836 (N_13836,N_12304,N_11159);
or U13837 (N_13837,N_10863,N_11530);
nand U13838 (N_13838,N_9854,N_10361);
and U13839 (N_13839,N_12189,N_10706);
nand U13840 (N_13840,N_11376,N_12229);
xnor U13841 (N_13841,N_9713,N_10440);
xor U13842 (N_13842,N_10255,N_11365);
and U13843 (N_13843,N_10381,N_11283);
or U13844 (N_13844,N_11444,N_10869);
or U13845 (N_13845,N_9698,N_11345);
and U13846 (N_13846,N_9931,N_12282);
or U13847 (N_13847,N_10745,N_9913);
nand U13848 (N_13848,N_11673,N_9593);
nor U13849 (N_13849,N_10495,N_10304);
nor U13850 (N_13850,N_10207,N_10993);
and U13851 (N_13851,N_12366,N_11366);
nand U13852 (N_13852,N_10727,N_11884);
xnor U13853 (N_13853,N_12376,N_12348);
nor U13854 (N_13854,N_11377,N_10177);
or U13855 (N_13855,N_9794,N_10530);
nand U13856 (N_13856,N_11597,N_11253);
nand U13857 (N_13857,N_11087,N_11643);
nand U13858 (N_13858,N_9501,N_11488);
nor U13859 (N_13859,N_10716,N_11613);
xnor U13860 (N_13860,N_9618,N_9492);
nor U13861 (N_13861,N_12356,N_11644);
xor U13862 (N_13862,N_10098,N_11293);
or U13863 (N_13863,N_9787,N_12467);
xor U13864 (N_13864,N_11166,N_10492);
nand U13865 (N_13865,N_11057,N_12219);
nand U13866 (N_13866,N_10965,N_10895);
xor U13867 (N_13867,N_12159,N_10423);
xor U13868 (N_13868,N_9642,N_9808);
xor U13869 (N_13869,N_10748,N_10198);
nor U13870 (N_13870,N_9410,N_9950);
nand U13871 (N_13871,N_9467,N_11948);
nor U13872 (N_13872,N_11648,N_9662);
or U13873 (N_13873,N_11452,N_11213);
and U13874 (N_13874,N_10216,N_11659);
xor U13875 (N_13875,N_10133,N_11205);
xnor U13876 (N_13876,N_10892,N_10516);
and U13877 (N_13877,N_10162,N_11867);
xor U13878 (N_13878,N_10144,N_12022);
xor U13879 (N_13879,N_11880,N_10955);
nor U13880 (N_13880,N_10244,N_11091);
xnor U13881 (N_13881,N_11248,N_9405);
nand U13882 (N_13882,N_10755,N_11801);
xnor U13883 (N_13883,N_10951,N_9379);
nand U13884 (N_13884,N_9842,N_9634);
nand U13885 (N_13885,N_9443,N_10468);
xnor U13886 (N_13886,N_11076,N_11954);
and U13887 (N_13887,N_11058,N_10403);
xnor U13888 (N_13888,N_10147,N_10889);
nand U13889 (N_13889,N_11709,N_12171);
nor U13890 (N_13890,N_11171,N_11779);
or U13891 (N_13891,N_10531,N_11493);
xor U13892 (N_13892,N_12058,N_11979);
and U13893 (N_13893,N_12443,N_10537);
nand U13894 (N_13894,N_10132,N_11415);
nand U13895 (N_13895,N_11772,N_9883);
nor U13896 (N_13896,N_11958,N_9716);
and U13897 (N_13897,N_11862,N_9708);
nand U13898 (N_13898,N_9892,N_10466);
nand U13899 (N_13899,N_10251,N_10397);
or U13900 (N_13900,N_10721,N_10184);
nor U13901 (N_13901,N_10669,N_12369);
and U13902 (N_13902,N_10064,N_10227);
nand U13903 (N_13903,N_9781,N_9600);
nor U13904 (N_13904,N_11967,N_12209);
nor U13905 (N_13905,N_9741,N_10682);
nand U13906 (N_13906,N_11047,N_12254);
nand U13907 (N_13907,N_10260,N_10235);
nor U13908 (N_13908,N_10793,N_11494);
nor U13909 (N_13909,N_11316,N_12327);
nor U13910 (N_13910,N_11963,N_11433);
nand U13911 (N_13911,N_10480,N_11352);
xnor U13912 (N_13912,N_12224,N_12441);
or U13913 (N_13913,N_12337,N_11395);
nand U13914 (N_13914,N_10734,N_11905);
and U13915 (N_13915,N_10881,N_10629);
xnor U13916 (N_13916,N_9636,N_10684);
xor U13917 (N_13917,N_9947,N_11155);
xor U13918 (N_13918,N_10232,N_10390);
nor U13919 (N_13919,N_9791,N_9519);
nor U13920 (N_13920,N_10559,N_11919);
or U13921 (N_13921,N_12069,N_11247);
and U13922 (N_13922,N_11161,N_12371);
and U13923 (N_13923,N_11757,N_10389);
xnor U13924 (N_13924,N_10986,N_11717);
xor U13925 (N_13925,N_10505,N_12203);
xnor U13926 (N_13926,N_11387,N_10311);
and U13927 (N_13927,N_10804,N_10365);
nor U13928 (N_13928,N_10775,N_11610);
xor U13929 (N_13929,N_9798,N_12220);
nor U13930 (N_13930,N_10632,N_10206);
and U13931 (N_13931,N_10195,N_11949);
xor U13932 (N_13932,N_11672,N_9531);
or U13933 (N_13933,N_11688,N_12280);
or U13934 (N_13934,N_11449,N_11930);
or U13935 (N_13935,N_10491,N_9571);
xnor U13936 (N_13936,N_12372,N_11637);
nand U13937 (N_13937,N_12221,N_10769);
or U13938 (N_13938,N_11819,N_12432);
nor U13939 (N_13939,N_9720,N_9909);
nand U13940 (N_13940,N_10455,N_11215);
nand U13941 (N_13941,N_9816,N_12032);
xnor U13942 (N_13942,N_9933,N_10518);
nor U13943 (N_13943,N_12263,N_10373);
and U13944 (N_13944,N_9470,N_10221);
nor U13945 (N_13945,N_12427,N_11416);
nand U13946 (N_13946,N_9488,N_9515);
and U13947 (N_13947,N_10957,N_11570);
or U13948 (N_13948,N_10384,N_12105);
or U13949 (N_13949,N_11323,N_10154);
and U13950 (N_13950,N_11642,N_9656);
and U13951 (N_13951,N_11094,N_10281);
or U13952 (N_13952,N_12308,N_9968);
and U13953 (N_13953,N_11541,N_9424);
or U13954 (N_13954,N_11578,N_11941);
and U13955 (N_13955,N_9438,N_11906);
nor U13956 (N_13956,N_11965,N_9558);
nor U13957 (N_13957,N_11165,N_11564);
nor U13958 (N_13958,N_9420,N_12222);
xnor U13959 (N_13959,N_11029,N_10685);
xnor U13960 (N_13960,N_11553,N_10724);
nor U13961 (N_13961,N_9528,N_10929);
nand U13962 (N_13962,N_9486,N_9898);
and U13963 (N_13963,N_10159,N_10662);
nand U13964 (N_13964,N_11882,N_10459);
or U13965 (N_13965,N_9498,N_11842);
and U13966 (N_13966,N_12357,N_11562);
and U13967 (N_13967,N_11615,N_12026);
xor U13968 (N_13968,N_10714,N_9757);
nor U13969 (N_13969,N_12196,N_12073);
nand U13970 (N_13970,N_10657,N_10058);
xnor U13971 (N_13971,N_11360,N_10425);
or U13972 (N_13972,N_9652,N_10187);
nand U13973 (N_13973,N_10948,N_12056);
xnor U13974 (N_13974,N_11093,N_10879);
and U13975 (N_13975,N_10514,N_11721);
nand U13976 (N_13976,N_10799,N_11997);
xor U13977 (N_13977,N_11471,N_10524);
and U13978 (N_13978,N_12192,N_9979);
and U13979 (N_13979,N_9635,N_9891);
xnor U13980 (N_13980,N_10846,N_9769);
nor U13981 (N_13981,N_11107,N_11774);
nor U13982 (N_13982,N_11933,N_9513);
xor U13983 (N_13983,N_11722,N_10686);
and U13984 (N_13984,N_10816,N_10402);
and U13985 (N_13985,N_10999,N_12346);
nand U13986 (N_13986,N_10426,N_10337);
xnor U13987 (N_13987,N_10408,N_10937);
and U13988 (N_13988,N_9397,N_9568);
and U13989 (N_13989,N_10380,N_10845);
and U13990 (N_13990,N_11946,N_9409);
nor U13991 (N_13991,N_10182,N_10458);
and U13992 (N_13992,N_9590,N_12402);
nand U13993 (N_13993,N_12028,N_11769);
nor U13994 (N_13994,N_9543,N_11973);
or U13995 (N_13995,N_11629,N_10600);
nor U13996 (N_13996,N_9401,N_10523);
nand U13997 (N_13997,N_9885,N_9585);
nor U13998 (N_13998,N_10149,N_9952);
or U13999 (N_13999,N_10097,N_12172);
xnor U14000 (N_14000,N_10751,N_10552);
xor U14001 (N_14001,N_12479,N_11117);
nand U14002 (N_14002,N_10160,N_9676);
and U14003 (N_14003,N_12463,N_10635);
or U14004 (N_14004,N_11217,N_9491);
xor U14005 (N_14005,N_10535,N_12042);
nand U14006 (N_14006,N_11139,N_11550);
or U14007 (N_14007,N_9803,N_9664);
or U14008 (N_14008,N_10226,N_10457);
xnor U14009 (N_14009,N_9609,N_10318);
and U14010 (N_14010,N_10237,N_12030);
and U14011 (N_14011,N_10517,N_11549);
nand U14012 (N_14012,N_9992,N_10729);
nand U14013 (N_14013,N_10582,N_10081);
and U14014 (N_14014,N_11762,N_11781);
nor U14015 (N_14015,N_9859,N_11732);
xnor U14016 (N_14016,N_11443,N_10019);
or U14017 (N_14017,N_11224,N_11490);
and U14018 (N_14018,N_11368,N_11596);
xnor U14019 (N_14019,N_10370,N_10291);
nor U14020 (N_14020,N_12179,N_9964);
or U14021 (N_14021,N_10428,N_12495);
xnor U14022 (N_14022,N_11350,N_11522);
nor U14023 (N_14023,N_10541,N_11699);
nor U14024 (N_14024,N_10616,N_10625);
xor U14025 (N_14025,N_10649,N_9684);
nand U14026 (N_14026,N_11186,N_9516);
xor U14027 (N_14027,N_10223,N_9481);
nand U14028 (N_14028,N_11628,N_11533);
nor U14029 (N_14029,N_11830,N_11968);
nor U14030 (N_14030,N_12160,N_9458);
xor U14031 (N_14031,N_10785,N_11981);
or U14032 (N_14032,N_12021,N_12397);
xor U14033 (N_14033,N_12340,N_9940);
nor U14034 (N_14034,N_9530,N_11843);
nand U14035 (N_14035,N_10609,N_9377);
nand U14036 (N_14036,N_9598,N_12414);
xor U14037 (N_14037,N_12387,N_9725);
nand U14038 (N_14038,N_10683,N_12064);
nor U14039 (N_14039,N_10125,N_9547);
and U14040 (N_14040,N_9802,N_9411);
nand U14041 (N_14041,N_10137,N_11814);
nor U14042 (N_14042,N_11575,N_11894);
and U14043 (N_14043,N_11276,N_10594);
xor U14044 (N_14044,N_10085,N_11599);
nor U14045 (N_14045,N_12457,N_9837);
nand U14046 (N_14046,N_11251,N_10358);
xnor U14047 (N_14047,N_11344,N_10005);
nand U14048 (N_14048,N_10835,N_12368);
nand U14049 (N_14049,N_12082,N_10697);
nand U14050 (N_14050,N_9446,N_10057);
xor U14051 (N_14051,N_11727,N_11992);
nor U14052 (N_14052,N_10464,N_12249);
nor U14053 (N_14053,N_11577,N_11496);
and U14054 (N_14054,N_11193,N_10968);
xnor U14055 (N_14055,N_10943,N_11434);
nand U14056 (N_14056,N_12496,N_11359);
nor U14057 (N_14057,N_9552,N_9387);
xnor U14058 (N_14058,N_10741,N_11264);
xor U14059 (N_14059,N_10926,N_12420);
nor U14060 (N_14060,N_10422,N_9523);
and U14061 (N_14061,N_10059,N_10407);
nand U14062 (N_14062,N_10424,N_10950);
or U14063 (N_14063,N_11973,N_10012);
xor U14064 (N_14064,N_10227,N_9562);
nand U14065 (N_14065,N_11319,N_12328);
nand U14066 (N_14066,N_9681,N_9563);
nand U14067 (N_14067,N_10175,N_11738);
xnor U14068 (N_14068,N_12215,N_12190);
or U14069 (N_14069,N_9627,N_10600);
or U14070 (N_14070,N_10098,N_11908);
xor U14071 (N_14071,N_10126,N_11327);
or U14072 (N_14072,N_11784,N_10356);
nor U14073 (N_14073,N_12408,N_9917);
or U14074 (N_14074,N_11323,N_12266);
nor U14075 (N_14075,N_10246,N_10401);
nand U14076 (N_14076,N_10199,N_9884);
xor U14077 (N_14077,N_9800,N_12394);
nor U14078 (N_14078,N_11748,N_11138);
and U14079 (N_14079,N_12361,N_10818);
and U14080 (N_14080,N_9702,N_10196);
nand U14081 (N_14081,N_11003,N_9492);
and U14082 (N_14082,N_10368,N_10462);
xnor U14083 (N_14083,N_11026,N_12468);
nor U14084 (N_14084,N_9519,N_11283);
and U14085 (N_14085,N_11448,N_10679);
nor U14086 (N_14086,N_11636,N_11639);
xor U14087 (N_14087,N_11959,N_9896);
or U14088 (N_14088,N_9385,N_11078);
nor U14089 (N_14089,N_10480,N_11777);
nand U14090 (N_14090,N_11074,N_10628);
nand U14091 (N_14091,N_9592,N_12413);
or U14092 (N_14092,N_11295,N_11580);
and U14093 (N_14093,N_11125,N_11070);
nor U14094 (N_14094,N_11358,N_10442);
and U14095 (N_14095,N_11912,N_10046);
or U14096 (N_14096,N_9747,N_9421);
nand U14097 (N_14097,N_9466,N_9639);
or U14098 (N_14098,N_12303,N_12341);
nor U14099 (N_14099,N_9505,N_10183);
nor U14100 (N_14100,N_9634,N_11220);
nand U14101 (N_14101,N_9567,N_12122);
or U14102 (N_14102,N_11619,N_9470);
nand U14103 (N_14103,N_10552,N_9411);
nand U14104 (N_14104,N_9843,N_10059);
nor U14105 (N_14105,N_12078,N_9759);
nand U14106 (N_14106,N_11838,N_9631);
xor U14107 (N_14107,N_12037,N_12030);
or U14108 (N_14108,N_12256,N_10110);
and U14109 (N_14109,N_11378,N_10527);
nor U14110 (N_14110,N_11291,N_11067);
nand U14111 (N_14111,N_9627,N_10928);
and U14112 (N_14112,N_9895,N_11308);
nand U14113 (N_14113,N_10690,N_11274);
nand U14114 (N_14114,N_10953,N_11566);
xnor U14115 (N_14115,N_11683,N_11739);
xor U14116 (N_14116,N_11723,N_9986);
or U14117 (N_14117,N_10214,N_11476);
xnor U14118 (N_14118,N_10664,N_11199);
nor U14119 (N_14119,N_10149,N_10023);
nand U14120 (N_14120,N_11158,N_12115);
and U14121 (N_14121,N_9909,N_12087);
or U14122 (N_14122,N_11712,N_11388);
nor U14123 (N_14123,N_10868,N_11351);
or U14124 (N_14124,N_9814,N_12249);
or U14125 (N_14125,N_12276,N_10450);
nand U14126 (N_14126,N_11362,N_10709);
nand U14127 (N_14127,N_10893,N_11479);
or U14128 (N_14128,N_11581,N_11532);
and U14129 (N_14129,N_11730,N_9512);
nor U14130 (N_14130,N_10089,N_11983);
xnor U14131 (N_14131,N_12338,N_9560);
nand U14132 (N_14132,N_9737,N_9393);
xnor U14133 (N_14133,N_11141,N_10891);
xor U14134 (N_14134,N_10744,N_11152);
or U14135 (N_14135,N_10420,N_11152);
and U14136 (N_14136,N_10857,N_9711);
or U14137 (N_14137,N_9723,N_11965);
nor U14138 (N_14138,N_9441,N_10779);
nand U14139 (N_14139,N_11131,N_10450);
xnor U14140 (N_14140,N_11867,N_10796);
and U14141 (N_14141,N_11775,N_12442);
and U14142 (N_14142,N_12215,N_10005);
xor U14143 (N_14143,N_11908,N_9675);
xnor U14144 (N_14144,N_9611,N_12406);
or U14145 (N_14145,N_9398,N_11368);
or U14146 (N_14146,N_11859,N_11394);
nor U14147 (N_14147,N_11786,N_11753);
and U14148 (N_14148,N_9705,N_12173);
or U14149 (N_14149,N_12447,N_11472);
nand U14150 (N_14150,N_9940,N_11186);
or U14151 (N_14151,N_11101,N_12159);
nor U14152 (N_14152,N_10565,N_11223);
or U14153 (N_14153,N_9410,N_11245);
or U14154 (N_14154,N_10731,N_10055);
nand U14155 (N_14155,N_11719,N_10820);
or U14156 (N_14156,N_11635,N_11000);
and U14157 (N_14157,N_10404,N_10691);
nor U14158 (N_14158,N_12262,N_9459);
or U14159 (N_14159,N_12251,N_10133);
or U14160 (N_14160,N_12114,N_12361);
nor U14161 (N_14161,N_11120,N_11030);
nand U14162 (N_14162,N_9874,N_11505);
nand U14163 (N_14163,N_11818,N_11503);
nor U14164 (N_14164,N_9786,N_9915);
nor U14165 (N_14165,N_10069,N_10411);
xor U14166 (N_14166,N_12228,N_12359);
or U14167 (N_14167,N_9756,N_10491);
nand U14168 (N_14168,N_11415,N_12318);
nand U14169 (N_14169,N_9411,N_12232);
nor U14170 (N_14170,N_9745,N_11884);
or U14171 (N_14171,N_10385,N_12496);
and U14172 (N_14172,N_12138,N_10678);
and U14173 (N_14173,N_10325,N_10216);
and U14174 (N_14174,N_12158,N_10560);
and U14175 (N_14175,N_10190,N_12286);
xor U14176 (N_14176,N_9820,N_12240);
or U14177 (N_14177,N_10273,N_9992);
and U14178 (N_14178,N_11975,N_11968);
or U14179 (N_14179,N_11074,N_10278);
xor U14180 (N_14180,N_10184,N_9666);
nor U14181 (N_14181,N_11023,N_10666);
nand U14182 (N_14182,N_10039,N_10901);
nor U14183 (N_14183,N_10911,N_12237);
xnor U14184 (N_14184,N_12314,N_10155);
nand U14185 (N_14185,N_11103,N_9384);
nand U14186 (N_14186,N_11589,N_12032);
nor U14187 (N_14187,N_11479,N_11599);
nor U14188 (N_14188,N_10246,N_11714);
and U14189 (N_14189,N_12095,N_12486);
or U14190 (N_14190,N_10182,N_11845);
and U14191 (N_14191,N_9692,N_11661);
xnor U14192 (N_14192,N_11851,N_9743);
xnor U14193 (N_14193,N_9455,N_11931);
nor U14194 (N_14194,N_11534,N_11182);
or U14195 (N_14195,N_11286,N_11548);
or U14196 (N_14196,N_11047,N_10301);
xnor U14197 (N_14197,N_11505,N_11191);
or U14198 (N_14198,N_9951,N_10551);
nand U14199 (N_14199,N_12146,N_12064);
or U14200 (N_14200,N_12079,N_11046);
or U14201 (N_14201,N_12463,N_11693);
or U14202 (N_14202,N_11573,N_10549);
and U14203 (N_14203,N_10769,N_11545);
xor U14204 (N_14204,N_10954,N_9831);
xnor U14205 (N_14205,N_9740,N_9742);
or U14206 (N_14206,N_9745,N_12041);
xor U14207 (N_14207,N_11101,N_11642);
or U14208 (N_14208,N_11488,N_12064);
and U14209 (N_14209,N_11647,N_11349);
or U14210 (N_14210,N_9519,N_11994);
nand U14211 (N_14211,N_10356,N_10930);
and U14212 (N_14212,N_9972,N_12065);
xnor U14213 (N_14213,N_10824,N_11950);
nor U14214 (N_14214,N_11954,N_10937);
nor U14215 (N_14215,N_10418,N_12310);
nand U14216 (N_14216,N_11355,N_11922);
or U14217 (N_14217,N_11011,N_10042);
xor U14218 (N_14218,N_11054,N_12017);
nand U14219 (N_14219,N_11385,N_12227);
nor U14220 (N_14220,N_11757,N_11095);
nand U14221 (N_14221,N_11160,N_9804);
or U14222 (N_14222,N_11355,N_11925);
or U14223 (N_14223,N_11163,N_11613);
or U14224 (N_14224,N_11935,N_10125);
nand U14225 (N_14225,N_11270,N_9812);
nand U14226 (N_14226,N_10105,N_11043);
or U14227 (N_14227,N_12263,N_10936);
nor U14228 (N_14228,N_9756,N_12254);
nor U14229 (N_14229,N_10743,N_12079);
xnor U14230 (N_14230,N_11510,N_10683);
or U14231 (N_14231,N_12103,N_12395);
nand U14232 (N_14232,N_10788,N_9731);
and U14233 (N_14233,N_12164,N_11223);
and U14234 (N_14234,N_9730,N_10497);
nand U14235 (N_14235,N_12375,N_9507);
nor U14236 (N_14236,N_10603,N_9405);
or U14237 (N_14237,N_10613,N_12432);
nor U14238 (N_14238,N_10291,N_11950);
nor U14239 (N_14239,N_10889,N_12244);
and U14240 (N_14240,N_9589,N_10835);
and U14241 (N_14241,N_10364,N_12478);
nand U14242 (N_14242,N_9818,N_10529);
or U14243 (N_14243,N_12187,N_10249);
or U14244 (N_14244,N_9811,N_12259);
or U14245 (N_14245,N_12360,N_9609);
xor U14246 (N_14246,N_11753,N_11814);
nor U14247 (N_14247,N_10770,N_12445);
nand U14248 (N_14248,N_10821,N_9929);
and U14249 (N_14249,N_10957,N_9396);
nor U14250 (N_14250,N_12042,N_11016);
xnor U14251 (N_14251,N_11513,N_11433);
xor U14252 (N_14252,N_10346,N_10915);
nor U14253 (N_14253,N_9483,N_9857);
xnor U14254 (N_14254,N_10251,N_10041);
xnor U14255 (N_14255,N_11968,N_10871);
nor U14256 (N_14256,N_11851,N_10084);
nand U14257 (N_14257,N_12415,N_10460);
and U14258 (N_14258,N_9468,N_10490);
xor U14259 (N_14259,N_9717,N_10834);
xor U14260 (N_14260,N_12343,N_9630);
and U14261 (N_14261,N_11944,N_12459);
and U14262 (N_14262,N_12075,N_10170);
nor U14263 (N_14263,N_11955,N_10883);
nor U14264 (N_14264,N_11303,N_9923);
or U14265 (N_14265,N_10765,N_10292);
and U14266 (N_14266,N_9902,N_10141);
and U14267 (N_14267,N_11856,N_11437);
nor U14268 (N_14268,N_9582,N_10611);
or U14269 (N_14269,N_11360,N_10624);
nand U14270 (N_14270,N_10949,N_10516);
nand U14271 (N_14271,N_11014,N_10152);
or U14272 (N_14272,N_11588,N_9940);
nor U14273 (N_14273,N_10427,N_10159);
nand U14274 (N_14274,N_11327,N_10847);
or U14275 (N_14275,N_10729,N_11258);
or U14276 (N_14276,N_12127,N_11260);
or U14277 (N_14277,N_10915,N_11777);
nor U14278 (N_14278,N_12439,N_11909);
xnor U14279 (N_14279,N_10231,N_10247);
xnor U14280 (N_14280,N_10367,N_10952);
and U14281 (N_14281,N_11778,N_11032);
or U14282 (N_14282,N_10045,N_9559);
nor U14283 (N_14283,N_10209,N_10093);
nor U14284 (N_14284,N_9590,N_11830);
nand U14285 (N_14285,N_10531,N_11393);
nor U14286 (N_14286,N_11793,N_9464);
and U14287 (N_14287,N_9890,N_12181);
nand U14288 (N_14288,N_10128,N_11168);
xnor U14289 (N_14289,N_10232,N_12044);
xor U14290 (N_14290,N_11061,N_12365);
and U14291 (N_14291,N_12472,N_9711);
or U14292 (N_14292,N_10974,N_12486);
nand U14293 (N_14293,N_9784,N_9383);
or U14294 (N_14294,N_11923,N_11361);
nand U14295 (N_14295,N_11348,N_10068);
or U14296 (N_14296,N_9464,N_10508);
nor U14297 (N_14297,N_11799,N_9553);
and U14298 (N_14298,N_11704,N_11278);
or U14299 (N_14299,N_11955,N_9940);
or U14300 (N_14300,N_10719,N_12393);
nand U14301 (N_14301,N_10797,N_12105);
xnor U14302 (N_14302,N_11222,N_10745);
or U14303 (N_14303,N_12275,N_10975);
nor U14304 (N_14304,N_9780,N_10840);
xnor U14305 (N_14305,N_10488,N_11418);
xnor U14306 (N_14306,N_11113,N_10118);
and U14307 (N_14307,N_9951,N_11900);
xnor U14308 (N_14308,N_11644,N_10361);
xor U14309 (N_14309,N_9887,N_10230);
and U14310 (N_14310,N_10631,N_10580);
nor U14311 (N_14311,N_10452,N_12219);
xor U14312 (N_14312,N_9995,N_11849);
or U14313 (N_14313,N_12434,N_10795);
and U14314 (N_14314,N_10188,N_9712);
nor U14315 (N_14315,N_12292,N_11321);
xor U14316 (N_14316,N_11377,N_11003);
nor U14317 (N_14317,N_11712,N_9749);
xor U14318 (N_14318,N_11879,N_12458);
nand U14319 (N_14319,N_12027,N_11537);
and U14320 (N_14320,N_10506,N_11717);
xor U14321 (N_14321,N_12355,N_12399);
and U14322 (N_14322,N_11216,N_9576);
and U14323 (N_14323,N_10172,N_11933);
nor U14324 (N_14324,N_9860,N_11274);
xnor U14325 (N_14325,N_10055,N_9870);
and U14326 (N_14326,N_12040,N_9983);
nand U14327 (N_14327,N_12378,N_10704);
or U14328 (N_14328,N_10625,N_12046);
nor U14329 (N_14329,N_9425,N_10467);
or U14330 (N_14330,N_10345,N_12462);
xnor U14331 (N_14331,N_9491,N_10177);
or U14332 (N_14332,N_10695,N_10537);
or U14333 (N_14333,N_11819,N_9988);
or U14334 (N_14334,N_11195,N_11872);
nor U14335 (N_14335,N_11549,N_11675);
xnor U14336 (N_14336,N_10750,N_10817);
xor U14337 (N_14337,N_9561,N_11623);
or U14338 (N_14338,N_12107,N_11809);
xor U14339 (N_14339,N_10712,N_11337);
or U14340 (N_14340,N_10411,N_11624);
and U14341 (N_14341,N_10427,N_10167);
nand U14342 (N_14342,N_9412,N_10073);
and U14343 (N_14343,N_11974,N_11842);
xnor U14344 (N_14344,N_12243,N_11424);
and U14345 (N_14345,N_11595,N_10567);
nand U14346 (N_14346,N_9559,N_12084);
and U14347 (N_14347,N_10000,N_11996);
or U14348 (N_14348,N_9536,N_11792);
or U14349 (N_14349,N_9398,N_11456);
or U14350 (N_14350,N_10638,N_11612);
nand U14351 (N_14351,N_9533,N_10048);
nand U14352 (N_14352,N_10782,N_10105);
nand U14353 (N_14353,N_12378,N_12278);
nand U14354 (N_14354,N_9934,N_11200);
or U14355 (N_14355,N_12253,N_9772);
nand U14356 (N_14356,N_10751,N_9714);
xor U14357 (N_14357,N_12309,N_12147);
nand U14358 (N_14358,N_10332,N_12115);
nor U14359 (N_14359,N_9396,N_9750);
or U14360 (N_14360,N_11118,N_10085);
nor U14361 (N_14361,N_9415,N_10020);
nor U14362 (N_14362,N_10758,N_10235);
nor U14363 (N_14363,N_11877,N_11702);
nor U14364 (N_14364,N_10813,N_9458);
nor U14365 (N_14365,N_11675,N_12258);
nand U14366 (N_14366,N_9709,N_11471);
and U14367 (N_14367,N_10749,N_12025);
xor U14368 (N_14368,N_12024,N_10644);
and U14369 (N_14369,N_10157,N_10463);
xnor U14370 (N_14370,N_10145,N_10206);
and U14371 (N_14371,N_10779,N_11349);
nand U14372 (N_14372,N_10081,N_9760);
or U14373 (N_14373,N_9699,N_9960);
nand U14374 (N_14374,N_11412,N_10873);
xor U14375 (N_14375,N_12405,N_10926);
and U14376 (N_14376,N_11617,N_9456);
or U14377 (N_14377,N_9858,N_10336);
nand U14378 (N_14378,N_11782,N_9745);
xor U14379 (N_14379,N_12379,N_10277);
nand U14380 (N_14380,N_10049,N_12397);
nand U14381 (N_14381,N_11028,N_9787);
nand U14382 (N_14382,N_9536,N_10801);
nor U14383 (N_14383,N_11036,N_10926);
or U14384 (N_14384,N_9865,N_10181);
xnor U14385 (N_14385,N_10577,N_10327);
or U14386 (N_14386,N_9395,N_10096);
or U14387 (N_14387,N_11115,N_10788);
or U14388 (N_14388,N_9375,N_11248);
nor U14389 (N_14389,N_9701,N_9375);
or U14390 (N_14390,N_10112,N_11486);
and U14391 (N_14391,N_11831,N_12480);
and U14392 (N_14392,N_9557,N_11990);
or U14393 (N_14393,N_11254,N_9653);
and U14394 (N_14394,N_11046,N_10547);
and U14395 (N_14395,N_11223,N_10069);
and U14396 (N_14396,N_12467,N_10769);
and U14397 (N_14397,N_10543,N_10947);
nor U14398 (N_14398,N_9416,N_12290);
nand U14399 (N_14399,N_12193,N_9677);
and U14400 (N_14400,N_12327,N_9970);
xor U14401 (N_14401,N_10107,N_10974);
and U14402 (N_14402,N_10517,N_11110);
nor U14403 (N_14403,N_11983,N_10256);
xnor U14404 (N_14404,N_11024,N_10225);
nor U14405 (N_14405,N_9600,N_12126);
or U14406 (N_14406,N_10991,N_9507);
and U14407 (N_14407,N_10909,N_10726);
xor U14408 (N_14408,N_10589,N_9944);
nand U14409 (N_14409,N_10688,N_9961);
nor U14410 (N_14410,N_10684,N_11184);
nor U14411 (N_14411,N_10066,N_11688);
nor U14412 (N_14412,N_10720,N_10776);
nand U14413 (N_14413,N_10546,N_12483);
or U14414 (N_14414,N_10669,N_10636);
xnor U14415 (N_14415,N_12113,N_12320);
xor U14416 (N_14416,N_10075,N_9448);
xnor U14417 (N_14417,N_12291,N_10395);
xnor U14418 (N_14418,N_10861,N_11001);
xnor U14419 (N_14419,N_12180,N_12007);
or U14420 (N_14420,N_9647,N_12432);
nor U14421 (N_14421,N_12258,N_12035);
or U14422 (N_14422,N_10692,N_11359);
xor U14423 (N_14423,N_9557,N_12177);
xnor U14424 (N_14424,N_9437,N_11518);
nand U14425 (N_14425,N_10528,N_10752);
and U14426 (N_14426,N_11164,N_10017);
and U14427 (N_14427,N_10060,N_11146);
or U14428 (N_14428,N_11805,N_12041);
xor U14429 (N_14429,N_12269,N_10030);
and U14430 (N_14430,N_12150,N_12422);
and U14431 (N_14431,N_10677,N_12199);
or U14432 (N_14432,N_10402,N_10931);
and U14433 (N_14433,N_10914,N_10575);
xor U14434 (N_14434,N_9962,N_9902);
and U14435 (N_14435,N_10038,N_11778);
or U14436 (N_14436,N_12098,N_12180);
nor U14437 (N_14437,N_10730,N_12213);
nor U14438 (N_14438,N_10269,N_12023);
nor U14439 (N_14439,N_11411,N_12443);
xor U14440 (N_14440,N_9512,N_10078);
xnor U14441 (N_14441,N_10393,N_10038);
and U14442 (N_14442,N_12342,N_11287);
and U14443 (N_14443,N_10352,N_10385);
nand U14444 (N_14444,N_10710,N_10388);
and U14445 (N_14445,N_11521,N_9691);
xnor U14446 (N_14446,N_11547,N_10454);
and U14447 (N_14447,N_11570,N_9684);
nor U14448 (N_14448,N_9719,N_12092);
nor U14449 (N_14449,N_10127,N_10080);
or U14450 (N_14450,N_11269,N_11771);
and U14451 (N_14451,N_12410,N_11801);
nor U14452 (N_14452,N_10155,N_9930);
nand U14453 (N_14453,N_10355,N_10725);
nor U14454 (N_14454,N_11772,N_11439);
or U14455 (N_14455,N_11160,N_10642);
nor U14456 (N_14456,N_10281,N_10412);
nand U14457 (N_14457,N_11956,N_11536);
nor U14458 (N_14458,N_9973,N_11483);
or U14459 (N_14459,N_12089,N_9462);
nand U14460 (N_14460,N_10719,N_11863);
xor U14461 (N_14461,N_11086,N_9697);
or U14462 (N_14462,N_12149,N_10194);
nand U14463 (N_14463,N_11590,N_10515);
nor U14464 (N_14464,N_10801,N_12261);
nor U14465 (N_14465,N_9444,N_10307);
nand U14466 (N_14466,N_10226,N_10353);
and U14467 (N_14467,N_10737,N_10608);
nand U14468 (N_14468,N_11200,N_11965);
nand U14469 (N_14469,N_11656,N_12418);
or U14470 (N_14470,N_10322,N_11052);
or U14471 (N_14471,N_10552,N_11399);
nor U14472 (N_14472,N_9871,N_10553);
nor U14473 (N_14473,N_12160,N_10333);
nand U14474 (N_14474,N_10097,N_11103);
nand U14475 (N_14475,N_9872,N_11613);
and U14476 (N_14476,N_11647,N_10897);
nand U14477 (N_14477,N_11273,N_12410);
or U14478 (N_14478,N_10305,N_11574);
and U14479 (N_14479,N_9587,N_11869);
or U14480 (N_14480,N_10061,N_9455);
xnor U14481 (N_14481,N_11543,N_11980);
or U14482 (N_14482,N_11401,N_9705);
nor U14483 (N_14483,N_11629,N_10885);
nor U14484 (N_14484,N_10420,N_11501);
xor U14485 (N_14485,N_11361,N_11700);
xnor U14486 (N_14486,N_10770,N_10358);
and U14487 (N_14487,N_11660,N_10914);
nor U14488 (N_14488,N_11560,N_10142);
nor U14489 (N_14489,N_9602,N_9645);
or U14490 (N_14490,N_9784,N_12202);
nor U14491 (N_14491,N_10335,N_9747);
and U14492 (N_14492,N_10500,N_10675);
xnor U14493 (N_14493,N_11590,N_10463);
nand U14494 (N_14494,N_9584,N_11481);
xor U14495 (N_14495,N_11163,N_10138);
xnor U14496 (N_14496,N_10544,N_11313);
or U14497 (N_14497,N_11271,N_11275);
nor U14498 (N_14498,N_10144,N_10168);
or U14499 (N_14499,N_9495,N_12483);
nand U14500 (N_14500,N_11232,N_9773);
and U14501 (N_14501,N_10505,N_10732);
nor U14502 (N_14502,N_10760,N_9930);
and U14503 (N_14503,N_10891,N_11996);
xnor U14504 (N_14504,N_10326,N_11065);
nand U14505 (N_14505,N_10937,N_11868);
or U14506 (N_14506,N_11676,N_9975);
nor U14507 (N_14507,N_12153,N_10238);
nor U14508 (N_14508,N_11819,N_11666);
and U14509 (N_14509,N_10925,N_9588);
xnor U14510 (N_14510,N_10941,N_10156);
nor U14511 (N_14511,N_10364,N_11311);
xor U14512 (N_14512,N_10079,N_11626);
and U14513 (N_14513,N_10107,N_12093);
nand U14514 (N_14514,N_11453,N_9735);
xor U14515 (N_14515,N_11239,N_10129);
and U14516 (N_14516,N_11746,N_12215);
nor U14517 (N_14517,N_11737,N_11887);
nand U14518 (N_14518,N_11716,N_9989);
nor U14519 (N_14519,N_11065,N_9439);
nor U14520 (N_14520,N_10460,N_11595);
xor U14521 (N_14521,N_11616,N_10629);
or U14522 (N_14522,N_9490,N_9824);
nand U14523 (N_14523,N_11559,N_12292);
or U14524 (N_14524,N_11440,N_10731);
and U14525 (N_14525,N_10841,N_11386);
xor U14526 (N_14526,N_11876,N_11587);
nand U14527 (N_14527,N_11208,N_9389);
xor U14528 (N_14528,N_10114,N_10878);
or U14529 (N_14529,N_12381,N_11453);
nand U14530 (N_14530,N_10109,N_12319);
nor U14531 (N_14531,N_9619,N_10181);
xnor U14532 (N_14532,N_10387,N_11879);
or U14533 (N_14533,N_10924,N_9411);
or U14534 (N_14534,N_10529,N_9378);
nor U14535 (N_14535,N_9764,N_10849);
xnor U14536 (N_14536,N_11939,N_10313);
nor U14537 (N_14537,N_9783,N_10869);
or U14538 (N_14538,N_11108,N_11495);
or U14539 (N_14539,N_11024,N_12135);
nor U14540 (N_14540,N_11251,N_10400);
nor U14541 (N_14541,N_9389,N_11065);
nor U14542 (N_14542,N_10502,N_12277);
or U14543 (N_14543,N_11343,N_12284);
and U14544 (N_14544,N_10506,N_11818);
or U14545 (N_14545,N_11283,N_11253);
nor U14546 (N_14546,N_12010,N_11982);
xnor U14547 (N_14547,N_10760,N_9645);
xnor U14548 (N_14548,N_10013,N_9436);
nor U14549 (N_14549,N_9580,N_11867);
and U14550 (N_14550,N_11553,N_11030);
or U14551 (N_14551,N_12246,N_11821);
nand U14552 (N_14552,N_12428,N_12018);
nor U14553 (N_14553,N_10634,N_10674);
nor U14554 (N_14554,N_9637,N_9969);
xor U14555 (N_14555,N_11322,N_11005);
nor U14556 (N_14556,N_11650,N_10357);
nor U14557 (N_14557,N_11811,N_9617);
and U14558 (N_14558,N_11814,N_11170);
or U14559 (N_14559,N_11126,N_11506);
or U14560 (N_14560,N_11931,N_11522);
nand U14561 (N_14561,N_10863,N_10073);
xor U14562 (N_14562,N_12187,N_11993);
nand U14563 (N_14563,N_12332,N_9564);
nor U14564 (N_14564,N_10750,N_11976);
nor U14565 (N_14565,N_11239,N_12484);
nand U14566 (N_14566,N_11785,N_11927);
and U14567 (N_14567,N_11369,N_11445);
or U14568 (N_14568,N_10377,N_10451);
nand U14569 (N_14569,N_11806,N_11058);
or U14570 (N_14570,N_10077,N_9713);
nand U14571 (N_14571,N_12397,N_9557);
nor U14572 (N_14572,N_11410,N_12387);
nor U14573 (N_14573,N_11841,N_12450);
xnor U14574 (N_14574,N_9945,N_12181);
xnor U14575 (N_14575,N_10476,N_11222);
nand U14576 (N_14576,N_11333,N_11932);
or U14577 (N_14577,N_12361,N_9837);
nand U14578 (N_14578,N_11125,N_11735);
xnor U14579 (N_14579,N_10747,N_11968);
xor U14580 (N_14580,N_10871,N_10729);
nor U14581 (N_14581,N_10626,N_9679);
nand U14582 (N_14582,N_12124,N_10441);
nor U14583 (N_14583,N_12366,N_11602);
nand U14584 (N_14584,N_12473,N_11855);
nor U14585 (N_14585,N_9948,N_12473);
nor U14586 (N_14586,N_12278,N_10505);
xor U14587 (N_14587,N_9535,N_11358);
and U14588 (N_14588,N_12246,N_10906);
xor U14589 (N_14589,N_9787,N_10450);
or U14590 (N_14590,N_10152,N_11708);
nor U14591 (N_14591,N_11529,N_10243);
and U14592 (N_14592,N_10972,N_12425);
and U14593 (N_14593,N_10871,N_9571);
and U14594 (N_14594,N_12276,N_11209);
xnor U14595 (N_14595,N_11872,N_10123);
nand U14596 (N_14596,N_11977,N_9724);
nor U14597 (N_14597,N_10419,N_11442);
and U14598 (N_14598,N_9768,N_9778);
nand U14599 (N_14599,N_11652,N_11393);
xor U14600 (N_14600,N_10804,N_10418);
and U14601 (N_14601,N_12186,N_12321);
nand U14602 (N_14602,N_11360,N_10085);
nand U14603 (N_14603,N_11226,N_9810);
or U14604 (N_14604,N_9641,N_10690);
and U14605 (N_14605,N_10137,N_9871);
or U14606 (N_14606,N_10299,N_11487);
nand U14607 (N_14607,N_10968,N_10604);
xnor U14608 (N_14608,N_11124,N_9554);
or U14609 (N_14609,N_12342,N_10255);
nor U14610 (N_14610,N_11751,N_10657);
xor U14611 (N_14611,N_10464,N_11883);
nor U14612 (N_14612,N_12314,N_10878);
nor U14613 (N_14613,N_10449,N_9610);
or U14614 (N_14614,N_10002,N_9684);
and U14615 (N_14615,N_10941,N_10714);
and U14616 (N_14616,N_11814,N_11487);
xor U14617 (N_14617,N_11293,N_10911);
xor U14618 (N_14618,N_9610,N_10410);
nand U14619 (N_14619,N_9991,N_11402);
xnor U14620 (N_14620,N_12334,N_10386);
nor U14621 (N_14621,N_11501,N_10460);
nor U14622 (N_14622,N_11500,N_10893);
nand U14623 (N_14623,N_11495,N_9424);
nand U14624 (N_14624,N_9599,N_11264);
nor U14625 (N_14625,N_9874,N_11118);
nor U14626 (N_14626,N_12081,N_11856);
nand U14627 (N_14627,N_11308,N_11323);
nand U14628 (N_14628,N_10599,N_11068);
nand U14629 (N_14629,N_9444,N_11388);
nand U14630 (N_14630,N_10075,N_9928);
xor U14631 (N_14631,N_12247,N_11938);
and U14632 (N_14632,N_9775,N_11044);
nor U14633 (N_14633,N_12179,N_10378);
nor U14634 (N_14634,N_11678,N_10892);
or U14635 (N_14635,N_11423,N_11923);
nor U14636 (N_14636,N_11606,N_11402);
and U14637 (N_14637,N_11099,N_11749);
nor U14638 (N_14638,N_10357,N_11459);
xor U14639 (N_14639,N_11680,N_9564);
or U14640 (N_14640,N_10753,N_11885);
nor U14641 (N_14641,N_10817,N_9711);
and U14642 (N_14642,N_10114,N_9958);
nand U14643 (N_14643,N_11804,N_11273);
nor U14644 (N_14644,N_10593,N_9733);
and U14645 (N_14645,N_12013,N_12390);
xnor U14646 (N_14646,N_9690,N_11525);
and U14647 (N_14647,N_11959,N_11427);
nor U14648 (N_14648,N_10237,N_11156);
or U14649 (N_14649,N_11117,N_10182);
xor U14650 (N_14650,N_12146,N_11153);
xnor U14651 (N_14651,N_11844,N_11549);
xor U14652 (N_14652,N_11713,N_11481);
nor U14653 (N_14653,N_11184,N_11100);
nor U14654 (N_14654,N_9633,N_9809);
or U14655 (N_14655,N_10116,N_11874);
and U14656 (N_14656,N_9526,N_12126);
and U14657 (N_14657,N_9939,N_10139);
xor U14658 (N_14658,N_9850,N_9939);
xnor U14659 (N_14659,N_11038,N_10537);
nor U14660 (N_14660,N_10764,N_12048);
and U14661 (N_14661,N_9920,N_10410);
xor U14662 (N_14662,N_10155,N_9686);
and U14663 (N_14663,N_9632,N_11927);
and U14664 (N_14664,N_9931,N_10838);
and U14665 (N_14665,N_12374,N_11223);
nand U14666 (N_14666,N_11293,N_11881);
nand U14667 (N_14667,N_9671,N_11575);
nand U14668 (N_14668,N_11792,N_9754);
xnor U14669 (N_14669,N_11472,N_9717);
and U14670 (N_14670,N_10719,N_9941);
and U14671 (N_14671,N_9398,N_11551);
or U14672 (N_14672,N_11891,N_10008);
nor U14673 (N_14673,N_12436,N_9475);
or U14674 (N_14674,N_10958,N_10657);
nor U14675 (N_14675,N_9495,N_10602);
and U14676 (N_14676,N_11112,N_11515);
nor U14677 (N_14677,N_10946,N_12279);
nand U14678 (N_14678,N_9879,N_9833);
xor U14679 (N_14679,N_11998,N_12229);
nor U14680 (N_14680,N_11206,N_11205);
or U14681 (N_14681,N_11121,N_9747);
or U14682 (N_14682,N_12349,N_11068);
nor U14683 (N_14683,N_10408,N_9417);
nand U14684 (N_14684,N_11464,N_10214);
nand U14685 (N_14685,N_10732,N_11460);
nor U14686 (N_14686,N_9996,N_11988);
nor U14687 (N_14687,N_10759,N_11957);
nand U14688 (N_14688,N_9961,N_12143);
or U14689 (N_14689,N_9854,N_10877);
nor U14690 (N_14690,N_12115,N_10082);
or U14691 (N_14691,N_11991,N_10120);
xor U14692 (N_14692,N_12229,N_9502);
nand U14693 (N_14693,N_11641,N_10190);
nand U14694 (N_14694,N_11236,N_9934);
and U14695 (N_14695,N_9769,N_10440);
or U14696 (N_14696,N_10184,N_10081);
nor U14697 (N_14697,N_11976,N_12024);
and U14698 (N_14698,N_11371,N_11356);
nor U14699 (N_14699,N_11344,N_11980);
and U14700 (N_14700,N_9380,N_12152);
or U14701 (N_14701,N_9696,N_9468);
xnor U14702 (N_14702,N_11264,N_11990);
nand U14703 (N_14703,N_11595,N_10394);
xnor U14704 (N_14704,N_10460,N_10277);
and U14705 (N_14705,N_9565,N_9654);
nor U14706 (N_14706,N_11810,N_9990);
xor U14707 (N_14707,N_11753,N_12408);
nor U14708 (N_14708,N_10900,N_12014);
xor U14709 (N_14709,N_10259,N_11356);
nor U14710 (N_14710,N_11428,N_9749);
nand U14711 (N_14711,N_12369,N_9714);
or U14712 (N_14712,N_10902,N_9719);
nor U14713 (N_14713,N_11429,N_9904);
xor U14714 (N_14714,N_11725,N_11902);
nand U14715 (N_14715,N_10286,N_11852);
or U14716 (N_14716,N_10587,N_10988);
xor U14717 (N_14717,N_9559,N_10837);
nand U14718 (N_14718,N_9726,N_12302);
and U14719 (N_14719,N_10103,N_10255);
xnor U14720 (N_14720,N_9414,N_10864);
xor U14721 (N_14721,N_9939,N_12331);
nand U14722 (N_14722,N_11108,N_10119);
nand U14723 (N_14723,N_11738,N_10257);
nor U14724 (N_14724,N_11674,N_9684);
nand U14725 (N_14725,N_10052,N_10756);
nand U14726 (N_14726,N_10826,N_9962);
xnor U14727 (N_14727,N_11780,N_11468);
xnor U14728 (N_14728,N_12419,N_9833);
nor U14729 (N_14729,N_10111,N_10854);
or U14730 (N_14730,N_10554,N_9992);
and U14731 (N_14731,N_11607,N_11614);
and U14732 (N_14732,N_10053,N_12203);
or U14733 (N_14733,N_11231,N_11024);
and U14734 (N_14734,N_11915,N_9717);
nand U14735 (N_14735,N_9575,N_10968);
or U14736 (N_14736,N_12121,N_10737);
and U14737 (N_14737,N_11144,N_11071);
nand U14738 (N_14738,N_11673,N_9835);
or U14739 (N_14739,N_12006,N_10451);
xnor U14740 (N_14740,N_10721,N_10265);
or U14741 (N_14741,N_11513,N_12323);
or U14742 (N_14742,N_9906,N_12202);
xor U14743 (N_14743,N_10236,N_11534);
nand U14744 (N_14744,N_10375,N_11410);
and U14745 (N_14745,N_12435,N_10347);
nor U14746 (N_14746,N_9784,N_10969);
or U14747 (N_14747,N_10059,N_12073);
and U14748 (N_14748,N_9870,N_10737);
xor U14749 (N_14749,N_11672,N_11762);
nor U14750 (N_14750,N_11966,N_9648);
or U14751 (N_14751,N_11493,N_12054);
and U14752 (N_14752,N_10470,N_10184);
xnor U14753 (N_14753,N_11388,N_11065);
and U14754 (N_14754,N_10678,N_10802);
and U14755 (N_14755,N_9872,N_12336);
nor U14756 (N_14756,N_10667,N_11099);
xnor U14757 (N_14757,N_11222,N_9576);
xor U14758 (N_14758,N_11865,N_11720);
nor U14759 (N_14759,N_10419,N_12271);
and U14760 (N_14760,N_11809,N_9580);
and U14761 (N_14761,N_9502,N_11801);
xnor U14762 (N_14762,N_10818,N_11269);
nor U14763 (N_14763,N_10359,N_9555);
xor U14764 (N_14764,N_11497,N_11119);
nand U14765 (N_14765,N_10014,N_10547);
nor U14766 (N_14766,N_11914,N_11962);
nand U14767 (N_14767,N_11474,N_11180);
nand U14768 (N_14768,N_12256,N_10381);
nand U14769 (N_14769,N_10167,N_11434);
and U14770 (N_14770,N_10019,N_10414);
nand U14771 (N_14771,N_12053,N_10301);
nor U14772 (N_14772,N_11819,N_10579);
xnor U14773 (N_14773,N_12404,N_9543);
or U14774 (N_14774,N_11196,N_11209);
nand U14775 (N_14775,N_11601,N_9708);
nand U14776 (N_14776,N_9971,N_10563);
nand U14777 (N_14777,N_10704,N_11896);
nand U14778 (N_14778,N_11149,N_9944);
nand U14779 (N_14779,N_11459,N_12246);
xnor U14780 (N_14780,N_9663,N_12122);
nand U14781 (N_14781,N_9385,N_12291);
and U14782 (N_14782,N_9510,N_12132);
and U14783 (N_14783,N_11124,N_9973);
and U14784 (N_14784,N_11566,N_12101);
xor U14785 (N_14785,N_12148,N_9985);
and U14786 (N_14786,N_11974,N_10710);
and U14787 (N_14787,N_10719,N_10552);
nand U14788 (N_14788,N_12430,N_9683);
nand U14789 (N_14789,N_11096,N_12374);
nand U14790 (N_14790,N_10256,N_11046);
and U14791 (N_14791,N_12426,N_11138);
or U14792 (N_14792,N_12323,N_12013);
nor U14793 (N_14793,N_11972,N_10039);
nand U14794 (N_14794,N_10690,N_12261);
nand U14795 (N_14795,N_9924,N_11536);
nand U14796 (N_14796,N_12329,N_11775);
nor U14797 (N_14797,N_11064,N_11990);
or U14798 (N_14798,N_11656,N_11641);
xor U14799 (N_14799,N_10639,N_10382);
or U14800 (N_14800,N_11046,N_10108);
or U14801 (N_14801,N_9971,N_10588);
nor U14802 (N_14802,N_12485,N_12223);
nor U14803 (N_14803,N_11450,N_10693);
nor U14804 (N_14804,N_9581,N_10635);
nor U14805 (N_14805,N_11433,N_11256);
xor U14806 (N_14806,N_9807,N_12248);
nor U14807 (N_14807,N_11947,N_10095);
xnor U14808 (N_14808,N_12376,N_11068);
nor U14809 (N_14809,N_9604,N_9470);
and U14810 (N_14810,N_11510,N_9874);
nor U14811 (N_14811,N_11606,N_9456);
or U14812 (N_14812,N_11224,N_12313);
and U14813 (N_14813,N_10442,N_12164);
nor U14814 (N_14814,N_11393,N_10863);
nor U14815 (N_14815,N_9643,N_11476);
nor U14816 (N_14816,N_9645,N_12052);
nand U14817 (N_14817,N_11921,N_9627);
xor U14818 (N_14818,N_11615,N_11493);
xor U14819 (N_14819,N_10772,N_12013);
or U14820 (N_14820,N_9619,N_12339);
or U14821 (N_14821,N_11534,N_10320);
nand U14822 (N_14822,N_12169,N_10819);
nand U14823 (N_14823,N_10511,N_11749);
nand U14824 (N_14824,N_9460,N_11160);
nor U14825 (N_14825,N_11693,N_9773);
xnor U14826 (N_14826,N_11004,N_10098);
nand U14827 (N_14827,N_10411,N_12327);
and U14828 (N_14828,N_10589,N_11944);
and U14829 (N_14829,N_12077,N_11249);
and U14830 (N_14830,N_9836,N_10332);
xor U14831 (N_14831,N_11466,N_9813);
or U14832 (N_14832,N_11934,N_11518);
xor U14833 (N_14833,N_12404,N_11359);
nor U14834 (N_14834,N_11415,N_11354);
xnor U14835 (N_14835,N_10444,N_11329);
nor U14836 (N_14836,N_11198,N_11336);
and U14837 (N_14837,N_11555,N_10646);
xnor U14838 (N_14838,N_11071,N_9892);
xor U14839 (N_14839,N_10432,N_10729);
and U14840 (N_14840,N_10069,N_10463);
xnor U14841 (N_14841,N_9928,N_11574);
nand U14842 (N_14842,N_11634,N_9859);
and U14843 (N_14843,N_10411,N_10727);
or U14844 (N_14844,N_9662,N_12358);
or U14845 (N_14845,N_10889,N_10417);
xor U14846 (N_14846,N_11823,N_11416);
and U14847 (N_14847,N_9602,N_10807);
nor U14848 (N_14848,N_11405,N_10750);
nor U14849 (N_14849,N_10620,N_10604);
or U14850 (N_14850,N_12122,N_12316);
nand U14851 (N_14851,N_10148,N_12351);
xnor U14852 (N_14852,N_11313,N_9908);
or U14853 (N_14853,N_10111,N_12104);
or U14854 (N_14854,N_10601,N_11241);
or U14855 (N_14855,N_12455,N_9454);
or U14856 (N_14856,N_10688,N_12268);
and U14857 (N_14857,N_10544,N_12486);
nor U14858 (N_14858,N_11617,N_9641);
nand U14859 (N_14859,N_10747,N_10314);
and U14860 (N_14860,N_10042,N_11054);
or U14861 (N_14861,N_9433,N_10943);
or U14862 (N_14862,N_10276,N_11717);
nor U14863 (N_14863,N_11507,N_9648);
or U14864 (N_14864,N_10565,N_10687);
nor U14865 (N_14865,N_11185,N_9597);
nor U14866 (N_14866,N_10398,N_9890);
nand U14867 (N_14867,N_11155,N_12461);
nand U14868 (N_14868,N_10342,N_11616);
nand U14869 (N_14869,N_9756,N_11299);
nand U14870 (N_14870,N_10629,N_10327);
xor U14871 (N_14871,N_9996,N_12082);
or U14872 (N_14872,N_10904,N_9804);
and U14873 (N_14873,N_10566,N_9578);
nand U14874 (N_14874,N_10638,N_9630);
and U14875 (N_14875,N_9823,N_12324);
or U14876 (N_14876,N_11068,N_11210);
or U14877 (N_14877,N_9388,N_12301);
nand U14878 (N_14878,N_12120,N_9980);
or U14879 (N_14879,N_11230,N_11783);
xnor U14880 (N_14880,N_12050,N_11216);
nor U14881 (N_14881,N_11292,N_11074);
and U14882 (N_14882,N_10828,N_10420);
and U14883 (N_14883,N_10713,N_10753);
and U14884 (N_14884,N_10392,N_9671);
or U14885 (N_14885,N_11129,N_10899);
xnor U14886 (N_14886,N_10262,N_10923);
or U14887 (N_14887,N_10550,N_10470);
xor U14888 (N_14888,N_11373,N_10231);
nor U14889 (N_14889,N_10254,N_9753);
xnor U14890 (N_14890,N_11224,N_9967);
nor U14891 (N_14891,N_9849,N_12063);
and U14892 (N_14892,N_9901,N_10839);
or U14893 (N_14893,N_10774,N_9401);
and U14894 (N_14894,N_10670,N_11823);
xnor U14895 (N_14895,N_10062,N_10897);
nor U14896 (N_14896,N_11125,N_10772);
or U14897 (N_14897,N_11056,N_10839);
nand U14898 (N_14898,N_12432,N_10331);
or U14899 (N_14899,N_12365,N_9490);
xnor U14900 (N_14900,N_11082,N_11231);
xor U14901 (N_14901,N_12275,N_9508);
nor U14902 (N_14902,N_11401,N_9673);
or U14903 (N_14903,N_11426,N_11514);
and U14904 (N_14904,N_10209,N_10890);
and U14905 (N_14905,N_11765,N_10509);
or U14906 (N_14906,N_10673,N_12476);
or U14907 (N_14907,N_9429,N_10593);
nand U14908 (N_14908,N_12308,N_11371);
and U14909 (N_14909,N_9753,N_9979);
or U14910 (N_14910,N_10359,N_10045);
and U14911 (N_14911,N_11802,N_10648);
and U14912 (N_14912,N_11851,N_10936);
or U14913 (N_14913,N_9889,N_12057);
xnor U14914 (N_14914,N_10190,N_9430);
and U14915 (N_14915,N_11521,N_10704);
nor U14916 (N_14916,N_11583,N_12329);
and U14917 (N_14917,N_9481,N_11107);
xor U14918 (N_14918,N_10762,N_11028);
nand U14919 (N_14919,N_11341,N_10793);
xor U14920 (N_14920,N_10050,N_9555);
and U14921 (N_14921,N_9577,N_11659);
nand U14922 (N_14922,N_10998,N_12302);
nand U14923 (N_14923,N_10886,N_10203);
nand U14924 (N_14924,N_11540,N_10884);
nor U14925 (N_14925,N_10124,N_9908);
or U14926 (N_14926,N_12416,N_9725);
nor U14927 (N_14927,N_11498,N_12021);
or U14928 (N_14928,N_11912,N_11071);
nor U14929 (N_14929,N_10824,N_9510);
or U14930 (N_14930,N_11134,N_10610);
xnor U14931 (N_14931,N_12180,N_11525);
nor U14932 (N_14932,N_10557,N_10378);
or U14933 (N_14933,N_10651,N_10453);
or U14934 (N_14934,N_12234,N_10913);
and U14935 (N_14935,N_11974,N_10678);
and U14936 (N_14936,N_9942,N_12412);
nand U14937 (N_14937,N_10586,N_11487);
nand U14938 (N_14938,N_9974,N_10308);
and U14939 (N_14939,N_10514,N_11083);
or U14940 (N_14940,N_12473,N_12187);
nor U14941 (N_14941,N_11740,N_10240);
and U14942 (N_14942,N_11562,N_11195);
or U14943 (N_14943,N_10987,N_11201);
and U14944 (N_14944,N_9399,N_9987);
nand U14945 (N_14945,N_10194,N_12234);
and U14946 (N_14946,N_10344,N_11486);
nand U14947 (N_14947,N_11795,N_10218);
nand U14948 (N_14948,N_10785,N_11078);
nand U14949 (N_14949,N_10541,N_12237);
nor U14950 (N_14950,N_11074,N_11711);
or U14951 (N_14951,N_9504,N_9499);
and U14952 (N_14952,N_10298,N_11233);
xnor U14953 (N_14953,N_10344,N_10555);
and U14954 (N_14954,N_11677,N_11262);
nor U14955 (N_14955,N_10121,N_11423);
xor U14956 (N_14956,N_9638,N_11060);
or U14957 (N_14957,N_11419,N_10138);
and U14958 (N_14958,N_11891,N_9824);
nor U14959 (N_14959,N_10668,N_11546);
nand U14960 (N_14960,N_11384,N_9955);
or U14961 (N_14961,N_12416,N_11433);
and U14962 (N_14962,N_10437,N_9980);
nand U14963 (N_14963,N_9568,N_11256);
nand U14964 (N_14964,N_10008,N_10338);
or U14965 (N_14965,N_11420,N_12401);
nand U14966 (N_14966,N_9592,N_12192);
nor U14967 (N_14967,N_10970,N_10607);
or U14968 (N_14968,N_10902,N_11581);
nand U14969 (N_14969,N_11987,N_10124);
nor U14970 (N_14970,N_10942,N_10543);
nand U14971 (N_14971,N_10155,N_10579);
nand U14972 (N_14972,N_11207,N_10015);
or U14973 (N_14973,N_11283,N_9721);
and U14974 (N_14974,N_9899,N_11896);
or U14975 (N_14975,N_10358,N_10719);
and U14976 (N_14976,N_10105,N_11624);
nor U14977 (N_14977,N_10599,N_10388);
nor U14978 (N_14978,N_10575,N_10337);
or U14979 (N_14979,N_12080,N_11830);
and U14980 (N_14980,N_9720,N_11622);
nand U14981 (N_14981,N_9509,N_10829);
or U14982 (N_14982,N_9893,N_10255);
nand U14983 (N_14983,N_12001,N_9991);
nand U14984 (N_14984,N_9660,N_10904);
nor U14985 (N_14985,N_12359,N_10276);
or U14986 (N_14986,N_9922,N_12282);
or U14987 (N_14987,N_11488,N_11370);
and U14988 (N_14988,N_11737,N_10184);
or U14989 (N_14989,N_12339,N_10801);
or U14990 (N_14990,N_10777,N_10640);
or U14991 (N_14991,N_10021,N_9447);
xnor U14992 (N_14992,N_11678,N_10415);
and U14993 (N_14993,N_11168,N_9459);
and U14994 (N_14994,N_11135,N_9979);
or U14995 (N_14995,N_10313,N_9819);
nor U14996 (N_14996,N_9926,N_10745);
and U14997 (N_14997,N_12229,N_11821);
and U14998 (N_14998,N_10003,N_9980);
nor U14999 (N_14999,N_12298,N_11617);
nor U15000 (N_15000,N_10875,N_11090);
xnor U15001 (N_15001,N_10475,N_9917);
nor U15002 (N_15002,N_11116,N_11693);
nand U15003 (N_15003,N_9965,N_10744);
nor U15004 (N_15004,N_12460,N_10655);
and U15005 (N_15005,N_11281,N_11373);
and U15006 (N_15006,N_11460,N_9408);
and U15007 (N_15007,N_11557,N_10255);
and U15008 (N_15008,N_10185,N_11044);
or U15009 (N_15009,N_10900,N_9722);
nor U15010 (N_15010,N_10055,N_11429);
nand U15011 (N_15011,N_11392,N_9986);
nand U15012 (N_15012,N_11295,N_10472);
nor U15013 (N_15013,N_9700,N_11883);
nor U15014 (N_15014,N_12396,N_10334);
or U15015 (N_15015,N_11193,N_11630);
xnor U15016 (N_15016,N_12299,N_11539);
or U15017 (N_15017,N_9832,N_9943);
nor U15018 (N_15018,N_9521,N_10178);
xnor U15019 (N_15019,N_10763,N_10292);
nor U15020 (N_15020,N_9685,N_11613);
xnor U15021 (N_15021,N_11790,N_9544);
nand U15022 (N_15022,N_12473,N_10124);
nor U15023 (N_15023,N_11416,N_12346);
nand U15024 (N_15024,N_10964,N_10123);
nand U15025 (N_15025,N_12175,N_9640);
nor U15026 (N_15026,N_11232,N_9835);
nand U15027 (N_15027,N_10360,N_10163);
or U15028 (N_15028,N_10880,N_9840);
nand U15029 (N_15029,N_12064,N_12398);
nand U15030 (N_15030,N_12084,N_10983);
xor U15031 (N_15031,N_11197,N_9718);
xor U15032 (N_15032,N_11633,N_12346);
or U15033 (N_15033,N_10154,N_10459);
xnor U15034 (N_15034,N_9422,N_11535);
nor U15035 (N_15035,N_9982,N_9655);
or U15036 (N_15036,N_10165,N_11714);
xor U15037 (N_15037,N_11059,N_11285);
nand U15038 (N_15038,N_11471,N_11391);
nor U15039 (N_15039,N_12382,N_10761);
xor U15040 (N_15040,N_10778,N_9649);
nand U15041 (N_15041,N_10406,N_12032);
nor U15042 (N_15042,N_11581,N_11092);
and U15043 (N_15043,N_11258,N_9893);
or U15044 (N_15044,N_10080,N_10880);
or U15045 (N_15045,N_9495,N_10253);
nor U15046 (N_15046,N_9691,N_11791);
nand U15047 (N_15047,N_11895,N_11545);
or U15048 (N_15048,N_11672,N_11710);
nand U15049 (N_15049,N_11781,N_11856);
and U15050 (N_15050,N_10221,N_10862);
or U15051 (N_15051,N_10983,N_10112);
or U15052 (N_15052,N_10889,N_11419);
or U15053 (N_15053,N_10509,N_10130);
nand U15054 (N_15054,N_12098,N_10596);
nand U15055 (N_15055,N_11580,N_12306);
and U15056 (N_15056,N_11265,N_11985);
nor U15057 (N_15057,N_10447,N_12457);
or U15058 (N_15058,N_10469,N_10126);
and U15059 (N_15059,N_10591,N_10095);
xnor U15060 (N_15060,N_12073,N_11176);
xnor U15061 (N_15061,N_9800,N_11065);
and U15062 (N_15062,N_11665,N_12166);
nand U15063 (N_15063,N_9913,N_9888);
xnor U15064 (N_15064,N_10730,N_11165);
nand U15065 (N_15065,N_9819,N_9489);
nor U15066 (N_15066,N_10031,N_9583);
and U15067 (N_15067,N_11857,N_11783);
xor U15068 (N_15068,N_11828,N_11165);
or U15069 (N_15069,N_12496,N_11156);
and U15070 (N_15070,N_12455,N_12000);
nand U15071 (N_15071,N_9898,N_10647);
or U15072 (N_15072,N_9913,N_10373);
and U15073 (N_15073,N_11482,N_9891);
and U15074 (N_15074,N_10752,N_10778);
xnor U15075 (N_15075,N_10638,N_12450);
xor U15076 (N_15076,N_9923,N_10361);
nor U15077 (N_15077,N_11708,N_9779);
or U15078 (N_15078,N_11663,N_10880);
nor U15079 (N_15079,N_12099,N_12006);
or U15080 (N_15080,N_10557,N_10912);
nand U15081 (N_15081,N_11364,N_9934);
and U15082 (N_15082,N_9472,N_9544);
nor U15083 (N_15083,N_11181,N_9655);
nand U15084 (N_15084,N_9447,N_11242);
or U15085 (N_15085,N_10225,N_10141);
nand U15086 (N_15086,N_11342,N_11491);
xor U15087 (N_15087,N_11906,N_9567);
nor U15088 (N_15088,N_11641,N_10252);
and U15089 (N_15089,N_11006,N_10535);
and U15090 (N_15090,N_11756,N_9759);
nand U15091 (N_15091,N_9834,N_12176);
xnor U15092 (N_15092,N_9899,N_10912);
and U15093 (N_15093,N_12216,N_12310);
nor U15094 (N_15094,N_11832,N_11005);
xor U15095 (N_15095,N_9613,N_11874);
xnor U15096 (N_15096,N_9394,N_11049);
xor U15097 (N_15097,N_10077,N_10679);
or U15098 (N_15098,N_11596,N_11468);
nand U15099 (N_15099,N_10371,N_11279);
and U15100 (N_15100,N_10134,N_9469);
or U15101 (N_15101,N_10053,N_9484);
nor U15102 (N_15102,N_12416,N_10905);
xor U15103 (N_15103,N_11488,N_11213);
xor U15104 (N_15104,N_10884,N_12169);
and U15105 (N_15105,N_9859,N_10910);
and U15106 (N_15106,N_12100,N_9790);
nor U15107 (N_15107,N_10835,N_10656);
xor U15108 (N_15108,N_11100,N_12305);
or U15109 (N_15109,N_9428,N_11978);
nand U15110 (N_15110,N_9434,N_10007);
nor U15111 (N_15111,N_9381,N_11116);
xnor U15112 (N_15112,N_9630,N_10688);
nor U15113 (N_15113,N_12146,N_10954);
and U15114 (N_15114,N_10572,N_9668);
or U15115 (N_15115,N_10864,N_12068);
or U15116 (N_15116,N_11206,N_10695);
nand U15117 (N_15117,N_12177,N_11475);
nand U15118 (N_15118,N_11452,N_10272);
or U15119 (N_15119,N_11686,N_11352);
nor U15120 (N_15120,N_12474,N_11125);
and U15121 (N_15121,N_9592,N_11396);
xor U15122 (N_15122,N_10916,N_10776);
xnor U15123 (N_15123,N_9425,N_10003);
nor U15124 (N_15124,N_11436,N_11309);
nor U15125 (N_15125,N_9962,N_10548);
xnor U15126 (N_15126,N_11571,N_11913);
or U15127 (N_15127,N_9878,N_12464);
nand U15128 (N_15128,N_12279,N_10874);
or U15129 (N_15129,N_11595,N_10259);
nand U15130 (N_15130,N_9650,N_9726);
or U15131 (N_15131,N_9830,N_10245);
and U15132 (N_15132,N_11181,N_12268);
nor U15133 (N_15133,N_11463,N_11445);
or U15134 (N_15134,N_10683,N_11077);
xor U15135 (N_15135,N_12026,N_12087);
or U15136 (N_15136,N_9490,N_10874);
nand U15137 (N_15137,N_10709,N_11642);
xnor U15138 (N_15138,N_10056,N_10601);
or U15139 (N_15139,N_12494,N_11555);
or U15140 (N_15140,N_9953,N_11535);
or U15141 (N_15141,N_9429,N_11185);
and U15142 (N_15142,N_11754,N_11455);
xor U15143 (N_15143,N_12426,N_11765);
or U15144 (N_15144,N_10095,N_9431);
nand U15145 (N_15145,N_10335,N_9894);
nand U15146 (N_15146,N_11770,N_9475);
nand U15147 (N_15147,N_10906,N_10558);
nand U15148 (N_15148,N_9641,N_12358);
and U15149 (N_15149,N_10420,N_10925);
nand U15150 (N_15150,N_9562,N_10060);
nor U15151 (N_15151,N_11802,N_12107);
nor U15152 (N_15152,N_9422,N_11391);
nand U15153 (N_15153,N_10606,N_11625);
nor U15154 (N_15154,N_12112,N_11321);
and U15155 (N_15155,N_11110,N_11441);
nor U15156 (N_15156,N_10576,N_11974);
or U15157 (N_15157,N_10130,N_12225);
or U15158 (N_15158,N_12290,N_11791);
nand U15159 (N_15159,N_9673,N_10981);
nor U15160 (N_15160,N_12355,N_12160);
nand U15161 (N_15161,N_9647,N_10460);
nand U15162 (N_15162,N_10590,N_11659);
and U15163 (N_15163,N_10727,N_12390);
nor U15164 (N_15164,N_9499,N_11294);
xor U15165 (N_15165,N_9839,N_11568);
and U15166 (N_15166,N_11056,N_12132);
or U15167 (N_15167,N_12111,N_10709);
nand U15168 (N_15168,N_9843,N_11734);
xor U15169 (N_15169,N_12293,N_10165);
nand U15170 (N_15170,N_11697,N_9388);
or U15171 (N_15171,N_12333,N_10936);
xnor U15172 (N_15172,N_9648,N_10786);
nor U15173 (N_15173,N_11129,N_11681);
nand U15174 (N_15174,N_10569,N_10214);
nand U15175 (N_15175,N_10347,N_11465);
nand U15176 (N_15176,N_12312,N_10799);
nand U15177 (N_15177,N_11999,N_9785);
xnor U15178 (N_15178,N_9980,N_9931);
xnor U15179 (N_15179,N_12100,N_11535);
or U15180 (N_15180,N_10978,N_10499);
nor U15181 (N_15181,N_11585,N_11832);
xor U15182 (N_15182,N_10811,N_10133);
and U15183 (N_15183,N_11724,N_11600);
xnor U15184 (N_15184,N_9936,N_10144);
nand U15185 (N_15185,N_10593,N_9998);
nand U15186 (N_15186,N_11606,N_9927);
nor U15187 (N_15187,N_12449,N_10426);
or U15188 (N_15188,N_9996,N_10079);
or U15189 (N_15189,N_11837,N_10981);
nand U15190 (N_15190,N_9676,N_9422);
and U15191 (N_15191,N_12109,N_9799);
or U15192 (N_15192,N_9810,N_12087);
and U15193 (N_15193,N_10916,N_9980);
xnor U15194 (N_15194,N_10865,N_10750);
and U15195 (N_15195,N_12334,N_10275);
xor U15196 (N_15196,N_10281,N_11368);
or U15197 (N_15197,N_9931,N_9922);
nor U15198 (N_15198,N_9889,N_12379);
and U15199 (N_15199,N_9803,N_11686);
nor U15200 (N_15200,N_11437,N_12194);
nor U15201 (N_15201,N_11126,N_9987);
or U15202 (N_15202,N_11661,N_11748);
nor U15203 (N_15203,N_11663,N_11406);
nand U15204 (N_15204,N_11585,N_9451);
and U15205 (N_15205,N_10799,N_12107);
nand U15206 (N_15206,N_11332,N_9457);
or U15207 (N_15207,N_11883,N_10825);
and U15208 (N_15208,N_10509,N_11965);
nand U15209 (N_15209,N_10409,N_9633);
xor U15210 (N_15210,N_10126,N_11496);
nor U15211 (N_15211,N_10635,N_11242);
xor U15212 (N_15212,N_10748,N_11626);
xnor U15213 (N_15213,N_9874,N_11259);
nor U15214 (N_15214,N_11234,N_9476);
xnor U15215 (N_15215,N_9915,N_9535);
nand U15216 (N_15216,N_11544,N_12239);
nor U15217 (N_15217,N_12334,N_11499);
nor U15218 (N_15218,N_12321,N_11290);
nor U15219 (N_15219,N_10604,N_12113);
and U15220 (N_15220,N_10675,N_10367);
or U15221 (N_15221,N_11133,N_9750);
xor U15222 (N_15222,N_11416,N_11628);
or U15223 (N_15223,N_11460,N_11199);
nand U15224 (N_15224,N_9859,N_10422);
nor U15225 (N_15225,N_11732,N_10971);
or U15226 (N_15226,N_10017,N_11162);
nor U15227 (N_15227,N_10946,N_12415);
nor U15228 (N_15228,N_10657,N_11256);
nor U15229 (N_15229,N_9715,N_10702);
xor U15230 (N_15230,N_11039,N_11955);
and U15231 (N_15231,N_10702,N_11797);
nor U15232 (N_15232,N_11860,N_10406);
nor U15233 (N_15233,N_10056,N_11185);
xnor U15234 (N_15234,N_11485,N_9953);
or U15235 (N_15235,N_11126,N_9686);
nand U15236 (N_15236,N_10499,N_11777);
nor U15237 (N_15237,N_10884,N_11036);
nor U15238 (N_15238,N_11377,N_10612);
nand U15239 (N_15239,N_11622,N_10415);
and U15240 (N_15240,N_11307,N_11862);
and U15241 (N_15241,N_12332,N_12330);
nand U15242 (N_15242,N_10000,N_11587);
nor U15243 (N_15243,N_11870,N_11260);
xnor U15244 (N_15244,N_12358,N_10354);
nand U15245 (N_15245,N_9559,N_9379);
and U15246 (N_15246,N_10586,N_11141);
and U15247 (N_15247,N_11835,N_11205);
nor U15248 (N_15248,N_10394,N_12209);
and U15249 (N_15249,N_11038,N_11363);
nand U15250 (N_15250,N_11972,N_11246);
xnor U15251 (N_15251,N_11326,N_11004);
nor U15252 (N_15252,N_10740,N_9428);
nor U15253 (N_15253,N_11394,N_10078);
or U15254 (N_15254,N_11813,N_12059);
xnor U15255 (N_15255,N_11619,N_11473);
nor U15256 (N_15256,N_11292,N_11313);
and U15257 (N_15257,N_10957,N_12488);
or U15258 (N_15258,N_10410,N_11280);
nand U15259 (N_15259,N_10423,N_11721);
xor U15260 (N_15260,N_11685,N_11536);
and U15261 (N_15261,N_11877,N_10676);
nand U15262 (N_15262,N_10193,N_10168);
xnor U15263 (N_15263,N_10819,N_11349);
and U15264 (N_15264,N_12215,N_11669);
xor U15265 (N_15265,N_11125,N_9878);
xnor U15266 (N_15266,N_10195,N_12210);
nor U15267 (N_15267,N_12134,N_10555);
and U15268 (N_15268,N_11402,N_9506);
xnor U15269 (N_15269,N_11307,N_12149);
nor U15270 (N_15270,N_9647,N_10934);
or U15271 (N_15271,N_9825,N_10124);
xnor U15272 (N_15272,N_10978,N_9716);
or U15273 (N_15273,N_11883,N_12187);
xnor U15274 (N_15274,N_11542,N_9511);
and U15275 (N_15275,N_11467,N_12023);
or U15276 (N_15276,N_11568,N_12035);
and U15277 (N_15277,N_10252,N_9381);
nor U15278 (N_15278,N_12037,N_12467);
xnor U15279 (N_15279,N_10492,N_12119);
and U15280 (N_15280,N_9703,N_10788);
or U15281 (N_15281,N_10401,N_10137);
or U15282 (N_15282,N_10386,N_10132);
xor U15283 (N_15283,N_10281,N_10584);
nor U15284 (N_15284,N_9978,N_9433);
and U15285 (N_15285,N_10945,N_11866);
and U15286 (N_15286,N_10534,N_12095);
nor U15287 (N_15287,N_10637,N_10106);
nand U15288 (N_15288,N_10240,N_9700);
nand U15289 (N_15289,N_10697,N_9462);
or U15290 (N_15290,N_10158,N_11897);
and U15291 (N_15291,N_10005,N_12412);
or U15292 (N_15292,N_12077,N_12013);
or U15293 (N_15293,N_10833,N_9761);
nor U15294 (N_15294,N_10870,N_9768);
nand U15295 (N_15295,N_10204,N_9872);
nor U15296 (N_15296,N_12065,N_10014);
or U15297 (N_15297,N_12135,N_9793);
or U15298 (N_15298,N_11572,N_12495);
nor U15299 (N_15299,N_9575,N_10259);
and U15300 (N_15300,N_10064,N_10099);
or U15301 (N_15301,N_9477,N_11401);
nand U15302 (N_15302,N_12053,N_12221);
nor U15303 (N_15303,N_10361,N_9379);
and U15304 (N_15304,N_9798,N_10851);
or U15305 (N_15305,N_11489,N_10662);
and U15306 (N_15306,N_10258,N_12324);
xor U15307 (N_15307,N_12249,N_10911);
xor U15308 (N_15308,N_11735,N_12433);
nor U15309 (N_15309,N_9587,N_9595);
xor U15310 (N_15310,N_11761,N_10206);
xnor U15311 (N_15311,N_12021,N_11242);
and U15312 (N_15312,N_9413,N_11179);
or U15313 (N_15313,N_11443,N_11996);
xnor U15314 (N_15314,N_10358,N_9390);
or U15315 (N_15315,N_11227,N_11560);
nor U15316 (N_15316,N_10082,N_11057);
or U15317 (N_15317,N_9875,N_9620);
xor U15318 (N_15318,N_12485,N_12059);
nand U15319 (N_15319,N_12291,N_11465);
xnor U15320 (N_15320,N_12477,N_10630);
nor U15321 (N_15321,N_12128,N_10773);
nand U15322 (N_15322,N_10618,N_9397);
xor U15323 (N_15323,N_10285,N_9817);
xnor U15324 (N_15324,N_9396,N_11690);
and U15325 (N_15325,N_11474,N_9674);
nor U15326 (N_15326,N_11943,N_10993);
or U15327 (N_15327,N_9690,N_11764);
and U15328 (N_15328,N_12062,N_10744);
nand U15329 (N_15329,N_11379,N_11884);
nand U15330 (N_15330,N_10344,N_11018);
and U15331 (N_15331,N_11097,N_12299);
and U15332 (N_15332,N_10037,N_11130);
nor U15333 (N_15333,N_11349,N_12462);
or U15334 (N_15334,N_12077,N_11444);
or U15335 (N_15335,N_10455,N_9935);
nand U15336 (N_15336,N_9532,N_10905);
or U15337 (N_15337,N_9883,N_11235);
or U15338 (N_15338,N_11653,N_12280);
nor U15339 (N_15339,N_12207,N_9680);
or U15340 (N_15340,N_12099,N_11682);
nor U15341 (N_15341,N_11233,N_12313);
and U15342 (N_15342,N_9846,N_10490);
nand U15343 (N_15343,N_10304,N_12151);
xnor U15344 (N_15344,N_10709,N_12271);
xnor U15345 (N_15345,N_10156,N_9559);
or U15346 (N_15346,N_11612,N_9946);
or U15347 (N_15347,N_12055,N_10289);
or U15348 (N_15348,N_10129,N_11222);
nand U15349 (N_15349,N_10698,N_9398);
nand U15350 (N_15350,N_11575,N_10365);
or U15351 (N_15351,N_10039,N_10967);
nand U15352 (N_15352,N_10801,N_10459);
nor U15353 (N_15353,N_10917,N_12428);
nand U15354 (N_15354,N_11004,N_12390);
nand U15355 (N_15355,N_11432,N_10226);
or U15356 (N_15356,N_9634,N_11528);
xor U15357 (N_15357,N_10615,N_10084);
nor U15358 (N_15358,N_11170,N_11867);
and U15359 (N_15359,N_9378,N_11467);
nand U15360 (N_15360,N_10145,N_11035);
nor U15361 (N_15361,N_10501,N_12106);
or U15362 (N_15362,N_11226,N_10805);
and U15363 (N_15363,N_10545,N_9688);
and U15364 (N_15364,N_9718,N_11199);
or U15365 (N_15365,N_11663,N_11567);
or U15366 (N_15366,N_11030,N_10369);
nor U15367 (N_15367,N_11957,N_9773);
nor U15368 (N_15368,N_9691,N_10099);
nor U15369 (N_15369,N_10608,N_10877);
xor U15370 (N_15370,N_10750,N_10006);
xor U15371 (N_15371,N_12223,N_11733);
or U15372 (N_15372,N_10966,N_12408);
nand U15373 (N_15373,N_10562,N_9992);
or U15374 (N_15374,N_10701,N_11179);
nor U15375 (N_15375,N_10588,N_10300);
and U15376 (N_15376,N_10468,N_11282);
nand U15377 (N_15377,N_11008,N_10075);
xnor U15378 (N_15378,N_10820,N_11074);
or U15379 (N_15379,N_10297,N_11156);
nand U15380 (N_15380,N_9537,N_11599);
and U15381 (N_15381,N_10639,N_9377);
xnor U15382 (N_15382,N_10097,N_11180);
or U15383 (N_15383,N_10639,N_10685);
xor U15384 (N_15384,N_9814,N_9376);
nand U15385 (N_15385,N_10996,N_9705);
nand U15386 (N_15386,N_11339,N_11390);
nor U15387 (N_15387,N_11169,N_12160);
nor U15388 (N_15388,N_11656,N_12306);
or U15389 (N_15389,N_12407,N_9429);
xnor U15390 (N_15390,N_12417,N_11061);
nor U15391 (N_15391,N_10629,N_10988);
xor U15392 (N_15392,N_9969,N_9631);
nand U15393 (N_15393,N_11087,N_11724);
or U15394 (N_15394,N_11685,N_11496);
nand U15395 (N_15395,N_10410,N_10232);
and U15396 (N_15396,N_10853,N_11897);
nor U15397 (N_15397,N_10926,N_10748);
xnor U15398 (N_15398,N_10265,N_11381);
or U15399 (N_15399,N_12117,N_12355);
or U15400 (N_15400,N_12097,N_11729);
or U15401 (N_15401,N_11858,N_10262);
and U15402 (N_15402,N_10439,N_9392);
and U15403 (N_15403,N_12080,N_11831);
and U15404 (N_15404,N_10776,N_10636);
and U15405 (N_15405,N_11223,N_10830);
xor U15406 (N_15406,N_10151,N_9451);
or U15407 (N_15407,N_11567,N_9518);
xnor U15408 (N_15408,N_10987,N_12197);
and U15409 (N_15409,N_9511,N_10075);
xor U15410 (N_15410,N_10233,N_10683);
nor U15411 (N_15411,N_9669,N_9624);
nor U15412 (N_15412,N_9911,N_10661);
xor U15413 (N_15413,N_11062,N_10336);
nand U15414 (N_15414,N_12009,N_11194);
or U15415 (N_15415,N_11061,N_11564);
or U15416 (N_15416,N_11309,N_11085);
nor U15417 (N_15417,N_10524,N_11357);
xor U15418 (N_15418,N_12205,N_11832);
nor U15419 (N_15419,N_11859,N_10124);
or U15420 (N_15420,N_10674,N_10174);
xnor U15421 (N_15421,N_11585,N_9704);
and U15422 (N_15422,N_12438,N_10874);
or U15423 (N_15423,N_11271,N_10146);
xor U15424 (N_15424,N_11873,N_11079);
xor U15425 (N_15425,N_10398,N_11470);
nor U15426 (N_15426,N_10110,N_11809);
nand U15427 (N_15427,N_10572,N_11234);
xnor U15428 (N_15428,N_11321,N_12272);
nand U15429 (N_15429,N_10149,N_12349);
or U15430 (N_15430,N_9543,N_12170);
or U15431 (N_15431,N_10898,N_11604);
nand U15432 (N_15432,N_11868,N_12085);
or U15433 (N_15433,N_9561,N_10576);
nor U15434 (N_15434,N_10065,N_11914);
nand U15435 (N_15435,N_10488,N_11244);
or U15436 (N_15436,N_11904,N_12300);
xor U15437 (N_15437,N_10224,N_11870);
or U15438 (N_15438,N_10986,N_10722);
nand U15439 (N_15439,N_10881,N_10753);
xnor U15440 (N_15440,N_12006,N_10575);
or U15441 (N_15441,N_10066,N_11523);
xor U15442 (N_15442,N_10071,N_12320);
nor U15443 (N_15443,N_11454,N_10467);
nor U15444 (N_15444,N_11626,N_12082);
xor U15445 (N_15445,N_11828,N_10532);
nand U15446 (N_15446,N_11302,N_12224);
xor U15447 (N_15447,N_11910,N_10269);
or U15448 (N_15448,N_11695,N_11158);
and U15449 (N_15449,N_11263,N_11497);
and U15450 (N_15450,N_12391,N_11606);
and U15451 (N_15451,N_10547,N_10149);
and U15452 (N_15452,N_10171,N_11049);
nand U15453 (N_15453,N_12430,N_9577);
or U15454 (N_15454,N_12028,N_10259);
and U15455 (N_15455,N_12131,N_11710);
xnor U15456 (N_15456,N_10679,N_10869);
and U15457 (N_15457,N_10646,N_10319);
and U15458 (N_15458,N_9569,N_11237);
nor U15459 (N_15459,N_11613,N_11731);
and U15460 (N_15460,N_11362,N_11729);
or U15461 (N_15461,N_10588,N_11298);
nand U15462 (N_15462,N_9764,N_10049);
nor U15463 (N_15463,N_11287,N_11009);
and U15464 (N_15464,N_10649,N_11097);
and U15465 (N_15465,N_10526,N_12341);
xnor U15466 (N_15466,N_11647,N_11381);
xor U15467 (N_15467,N_10575,N_11199);
nor U15468 (N_15468,N_11498,N_10000);
or U15469 (N_15469,N_9956,N_9720);
and U15470 (N_15470,N_9529,N_10134);
or U15471 (N_15471,N_10857,N_11465);
nor U15472 (N_15472,N_9678,N_12026);
or U15473 (N_15473,N_11411,N_12058);
xor U15474 (N_15474,N_11088,N_11439);
and U15475 (N_15475,N_10662,N_11221);
nand U15476 (N_15476,N_9810,N_11969);
nand U15477 (N_15477,N_10119,N_11550);
or U15478 (N_15478,N_10424,N_12386);
xnor U15479 (N_15479,N_9936,N_11665);
nor U15480 (N_15480,N_9720,N_9706);
nand U15481 (N_15481,N_9921,N_10178);
nor U15482 (N_15482,N_10339,N_11053);
nand U15483 (N_15483,N_10113,N_9441);
nor U15484 (N_15484,N_12158,N_12300);
nand U15485 (N_15485,N_9746,N_11438);
or U15486 (N_15486,N_10073,N_9690);
or U15487 (N_15487,N_11181,N_12403);
and U15488 (N_15488,N_11421,N_9648);
xnor U15489 (N_15489,N_10076,N_10522);
xnor U15490 (N_15490,N_12005,N_9652);
nor U15491 (N_15491,N_9964,N_10621);
and U15492 (N_15492,N_11304,N_9840);
nor U15493 (N_15493,N_11222,N_12381);
or U15494 (N_15494,N_10302,N_9502);
or U15495 (N_15495,N_11059,N_11428);
nand U15496 (N_15496,N_9592,N_11407);
or U15497 (N_15497,N_11778,N_9650);
and U15498 (N_15498,N_10128,N_11124);
nor U15499 (N_15499,N_10961,N_11487);
nand U15500 (N_15500,N_11408,N_12068);
xor U15501 (N_15501,N_11840,N_10016);
nand U15502 (N_15502,N_10243,N_12235);
or U15503 (N_15503,N_12422,N_11477);
nor U15504 (N_15504,N_9627,N_12397);
and U15505 (N_15505,N_9542,N_10747);
and U15506 (N_15506,N_10051,N_11000);
nand U15507 (N_15507,N_10408,N_10163);
and U15508 (N_15508,N_9633,N_12374);
or U15509 (N_15509,N_9504,N_11037);
nor U15510 (N_15510,N_11325,N_11329);
nor U15511 (N_15511,N_12208,N_10561);
and U15512 (N_15512,N_12492,N_9956);
nor U15513 (N_15513,N_11154,N_11782);
and U15514 (N_15514,N_9626,N_12371);
or U15515 (N_15515,N_11594,N_12111);
nand U15516 (N_15516,N_10641,N_10681);
or U15517 (N_15517,N_9387,N_10920);
and U15518 (N_15518,N_9717,N_10091);
and U15519 (N_15519,N_9572,N_9717);
nand U15520 (N_15520,N_11568,N_11701);
xnor U15521 (N_15521,N_9826,N_11422);
xnor U15522 (N_15522,N_10764,N_10479);
or U15523 (N_15523,N_10990,N_12436);
xnor U15524 (N_15524,N_11803,N_11218);
xor U15525 (N_15525,N_9463,N_11065);
or U15526 (N_15526,N_11558,N_9445);
or U15527 (N_15527,N_12439,N_10759);
and U15528 (N_15528,N_10725,N_9455);
and U15529 (N_15529,N_12238,N_11422);
nor U15530 (N_15530,N_11317,N_11794);
nor U15531 (N_15531,N_11164,N_10269);
and U15532 (N_15532,N_11957,N_10362);
or U15533 (N_15533,N_11983,N_10455);
nand U15534 (N_15534,N_11759,N_11312);
nor U15535 (N_15535,N_11273,N_11481);
or U15536 (N_15536,N_11760,N_10470);
and U15537 (N_15537,N_10951,N_10330);
or U15538 (N_15538,N_11500,N_9673);
xnor U15539 (N_15539,N_10023,N_11011);
xnor U15540 (N_15540,N_12150,N_11349);
nand U15541 (N_15541,N_9448,N_9952);
xor U15542 (N_15542,N_10155,N_12492);
or U15543 (N_15543,N_9992,N_11851);
and U15544 (N_15544,N_11143,N_11111);
xnor U15545 (N_15545,N_10314,N_11853);
nor U15546 (N_15546,N_9887,N_10496);
and U15547 (N_15547,N_10814,N_10682);
nor U15548 (N_15548,N_11499,N_11855);
and U15549 (N_15549,N_12088,N_10005);
nand U15550 (N_15550,N_10160,N_11115);
and U15551 (N_15551,N_11449,N_10822);
xor U15552 (N_15552,N_9885,N_10252);
and U15553 (N_15553,N_11653,N_10655);
xor U15554 (N_15554,N_9827,N_11885);
nand U15555 (N_15555,N_10892,N_9748);
nand U15556 (N_15556,N_12386,N_9991);
and U15557 (N_15557,N_11619,N_10284);
or U15558 (N_15558,N_9979,N_10775);
or U15559 (N_15559,N_9783,N_11206);
nor U15560 (N_15560,N_9783,N_11537);
or U15561 (N_15561,N_10343,N_10053);
or U15562 (N_15562,N_9433,N_10407);
nand U15563 (N_15563,N_10501,N_9710);
nor U15564 (N_15564,N_11470,N_10580);
xnor U15565 (N_15565,N_11024,N_12213);
or U15566 (N_15566,N_10184,N_10583);
nand U15567 (N_15567,N_10342,N_11761);
nor U15568 (N_15568,N_12497,N_10937);
xor U15569 (N_15569,N_9418,N_9595);
xnor U15570 (N_15570,N_11006,N_11036);
nand U15571 (N_15571,N_11948,N_12457);
nor U15572 (N_15572,N_9815,N_10604);
and U15573 (N_15573,N_10483,N_9898);
nand U15574 (N_15574,N_10575,N_12208);
xnor U15575 (N_15575,N_10182,N_10534);
or U15576 (N_15576,N_11472,N_10087);
xor U15577 (N_15577,N_11413,N_10949);
nor U15578 (N_15578,N_9450,N_9933);
xor U15579 (N_15579,N_10037,N_9630);
nor U15580 (N_15580,N_12263,N_10567);
nand U15581 (N_15581,N_11013,N_11821);
or U15582 (N_15582,N_12360,N_12258);
xnor U15583 (N_15583,N_9625,N_9773);
nand U15584 (N_15584,N_12053,N_9880);
nor U15585 (N_15585,N_11185,N_10471);
xor U15586 (N_15586,N_12413,N_12205);
xnor U15587 (N_15587,N_9730,N_9492);
nor U15588 (N_15588,N_9967,N_9618);
xnor U15589 (N_15589,N_9726,N_9767);
nand U15590 (N_15590,N_10962,N_11465);
nand U15591 (N_15591,N_9797,N_12264);
xor U15592 (N_15592,N_9721,N_11799);
or U15593 (N_15593,N_9909,N_9649);
and U15594 (N_15594,N_12204,N_10857);
xnor U15595 (N_15595,N_11865,N_12283);
xnor U15596 (N_15596,N_12130,N_11089);
xor U15597 (N_15597,N_10248,N_10306);
nand U15598 (N_15598,N_11810,N_10137);
xnor U15599 (N_15599,N_10945,N_11599);
and U15600 (N_15600,N_9411,N_12077);
or U15601 (N_15601,N_11118,N_11359);
nor U15602 (N_15602,N_11286,N_10681);
nor U15603 (N_15603,N_11166,N_11636);
xor U15604 (N_15604,N_12459,N_10161);
nor U15605 (N_15605,N_11916,N_9470);
xor U15606 (N_15606,N_11829,N_12197);
xor U15607 (N_15607,N_9996,N_9420);
xor U15608 (N_15608,N_11284,N_10703);
and U15609 (N_15609,N_11633,N_9440);
nand U15610 (N_15610,N_12486,N_9467);
nand U15611 (N_15611,N_11448,N_10890);
xor U15612 (N_15612,N_11926,N_11804);
nor U15613 (N_15613,N_11153,N_12022);
and U15614 (N_15614,N_9636,N_11806);
xnor U15615 (N_15615,N_9446,N_9614);
and U15616 (N_15616,N_11524,N_10823);
nor U15617 (N_15617,N_9925,N_11643);
or U15618 (N_15618,N_11785,N_11147);
and U15619 (N_15619,N_11213,N_10077);
nand U15620 (N_15620,N_11311,N_10102);
nor U15621 (N_15621,N_9733,N_11757);
or U15622 (N_15622,N_10363,N_10537);
nand U15623 (N_15623,N_10827,N_11289);
xnor U15624 (N_15624,N_10602,N_10316);
or U15625 (N_15625,N_12630,N_12897);
nor U15626 (N_15626,N_13278,N_13127);
nor U15627 (N_15627,N_13651,N_12570);
nand U15628 (N_15628,N_13062,N_13186);
and U15629 (N_15629,N_15238,N_13953);
or U15630 (N_15630,N_13320,N_14361);
nand U15631 (N_15631,N_13302,N_15057);
nor U15632 (N_15632,N_15018,N_13284);
xnor U15633 (N_15633,N_14209,N_13585);
or U15634 (N_15634,N_13670,N_14268);
xor U15635 (N_15635,N_15390,N_15250);
nor U15636 (N_15636,N_12958,N_12770);
and U15637 (N_15637,N_14971,N_13477);
nor U15638 (N_15638,N_15232,N_14937);
or U15639 (N_15639,N_14002,N_14043);
xor U15640 (N_15640,N_14530,N_13531);
nand U15641 (N_15641,N_15564,N_13885);
and U15642 (N_15642,N_14348,N_13222);
or U15643 (N_15643,N_12542,N_14048);
nor U15644 (N_15644,N_14683,N_13747);
or U15645 (N_15645,N_13895,N_13425);
nand U15646 (N_15646,N_15046,N_12774);
nand U15647 (N_15647,N_13577,N_12724);
nor U15648 (N_15648,N_14944,N_14239);
xnor U15649 (N_15649,N_15227,N_14916);
xor U15650 (N_15650,N_12930,N_14691);
and U15651 (N_15651,N_14791,N_15084);
nor U15652 (N_15652,N_14198,N_15460);
or U15653 (N_15653,N_14872,N_14474);
or U15654 (N_15654,N_14514,N_13767);
nor U15655 (N_15655,N_15059,N_14203);
xnor U15656 (N_15656,N_14140,N_13815);
or U15657 (N_15657,N_13117,N_13824);
or U15658 (N_15658,N_13015,N_15619);
nand U15659 (N_15659,N_13305,N_15357);
and U15660 (N_15660,N_15408,N_12628);
xor U15661 (N_15661,N_14248,N_15544);
nand U15662 (N_15662,N_14958,N_14966);
and U15663 (N_15663,N_13264,N_13259);
or U15664 (N_15664,N_14995,N_14339);
nand U15665 (N_15665,N_14484,N_13109);
xnor U15666 (N_15666,N_15079,N_14125);
or U15667 (N_15667,N_14420,N_15085);
nand U15668 (N_15668,N_14614,N_15493);
or U15669 (N_15669,N_15511,N_14572);
nor U15670 (N_15670,N_13751,N_13151);
or U15671 (N_15671,N_12689,N_12504);
and U15672 (N_15672,N_15299,N_13846);
nor U15673 (N_15673,N_14708,N_14697);
or U15674 (N_15674,N_14347,N_14032);
nand U15675 (N_15675,N_14326,N_14765);
xor U15676 (N_15676,N_13635,N_13737);
nand U15677 (N_15677,N_14724,N_14055);
or U15678 (N_15678,N_14928,N_14289);
and U15679 (N_15679,N_13503,N_14781);
xor U15680 (N_15680,N_13311,N_13066);
nand U15681 (N_15681,N_15533,N_14386);
nand U15682 (N_15682,N_12988,N_15108);
nor U15683 (N_15683,N_14495,N_15172);
nand U15684 (N_15684,N_13816,N_14573);
and U15685 (N_15685,N_12808,N_14416);
and U15686 (N_15686,N_15450,N_14899);
nand U15687 (N_15687,N_14360,N_13628);
nor U15688 (N_15688,N_12629,N_14739);
nor U15689 (N_15689,N_14030,N_12766);
or U15690 (N_15690,N_13756,N_15235);
nor U15691 (N_15691,N_13123,N_15008);
nand U15692 (N_15692,N_12878,N_14210);
xnor U15693 (N_15693,N_14445,N_13579);
nor U15694 (N_15694,N_14143,N_12627);
nand U15695 (N_15695,N_14710,N_12926);
nor U15696 (N_15696,N_14828,N_13605);
nand U15697 (N_15697,N_14450,N_14687);
xnor U15698 (N_15698,N_14852,N_13021);
nand U15699 (N_15699,N_15548,N_15590);
or U15700 (N_15700,N_12508,N_14806);
nor U15701 (N_15701,N_14517,N_14776);
xor U15702 (N_15702,N_12718,N_15483);
nor U15703 (N_15703,N_13408,N_13580);
or U15704 (N_15704,N_13656,N_13863);
or U15705 (N_15705,N_15394,N_12530);
or U15706 (N_15706,N_12967,N_15426);
and U15707 (N_15707,N_12756,N_14940);
or U15708 (N_15708,N_14583,N_14258);
nor U15709 (N_15709,N_15141,N_13060);
or U15710 (N_15710,N_15127,N_13958);
xor U15711 (N_15711,N_15262,N_15410);
nor U15712 (N_15712,N_14058,N_15479);
nand U15713 (N_15713,N_13493,N_13598);
nor U15714 (N_15714,N_13698,N_13052);
or U15715 (N_15715,N_15582,N_13257);
xnor U15716 (N_15716,N_12875,N_13215);
xnor U15717 (N_15717,N_15516,N_13592);
nor U15718 (N_15718,N_13188,N_13119);
or U15719 (N_15719,N_14300,N_14723);
or U15720 (N_15720,N_13560,N_14242);
xor U15721 (N_15721,N_12747,N_15505);
nand U15722 (N_15722,N_13378,N_14110);
nand U15723 (N_15723,N_14667,N_14840);
nor U15724 (N_15724,N_14423,N_14369);
nand U15725 (N_15725,N_14991,N_14458);
nor U15726 (N_15726,N_15346,N_14276);
and U15727 (N_15727,N_14205,N_14860);
nand U15728 (N_15728,N_15024,N_14431);
and U15729 (N_15729,N_15324,N_14149);
nor U15730 (N_15730,N_13349,N_15029);
or U15731 (N_15731,N_12996,N_14465);
nor U15732 (N_15732,N_14603,N_15060);
xnor U15733 (N_15733,N_14640,N_14615);
nor U15734 (N_15734,N_15378,N_12802);
nor U15735 (N_15735,N_14936,N_13999);
nor U15736 (N_15736,N_13202,N_12914);
xor U15737 (N_15737,N_15451,N_13943);
xnor U15738 (N_15738,N_14832,N_13083);
or U15739 (N_15739,N_12782,N_14858);
nand U15740 (N_15740,N_14690,N_14113);
nand U15741 (N_15741,N_13982,N_15209);
nor U15742 (N_15742,N_13399,N_13865);
and U15743 (N_15743,N_15092,N_14882);
xnor U15744 (N_15744,N_14174,N_13969);
and U15745 (N_15745,N_13325,N_14673);
and U15746 (N_15746,N_14121,N_14146);
xor U15747 (N_15747,N_13498,N_13077);
or U15748 (N_15748,N_15102,N_13534);
and U15749 (N_15749,N_13744,N_13867);
nor U15750 (N_15750,N_15143,N_15443);
nor U15751 (N_15751,N_14275,N_15555);
nor U15752 (N_15752,N_12859,N_14972);
and U15753 (N_15753,N_14273,N_14492);
nand U15754 (N_15754,N_13415,N_14421);
or U15755 (N_15755,N_15195,N_12863);
and U15756 (N_15756,N_12688,N_15042);
xnor U15757 (N_15757,N_14631,N_14750);
xor U15758 (N_15758,N_13100,N_14184);
nand U15759 (N_15759,N_12745,N_13307);
and U15760 (N_15760,N_14227,N_14861);
and U15761 (N_15761,N_14133,N_12963);
or U15762 (N_15762,N_13096,N_14062);
nor U15763 (N_15763,N_15362,N_13804);
xor U15764 (N_15764,N_13900,N_15184);
nor U15765 (N_15765,N_14969,N_14853);
nand U15766 (N_15766,N_13960,N_13382);
and U15767 (N_15767,N_13819,N_13987);
nand U15768 (N_15768,N_13207,N_14986);
xor U15769 (N_15769,N_12757,N_13921);
and U15770 (N_15770,N_14012,N_15325);
and U15771 (N_15771,N_12526,N_14760);
nand U15772 (N_15772,N_15167,N_14523);
and U15773 (N_15773,N_15306,N_15570);
nor U15774 (N_15774,N_15313,N_13221);
or U15775 (N_15775,N_14443,N_14512);
xor U15776 (N_15776,N_14357,N_13682);
or U15777 (N_15777,N_12719,N_13770);
nor U15778 (N_15778,N_14060,N_12590);
or U15779 (N_15779,N_15597,N_15407);
nand U15780 (N_15780,N_14897,N_15073);
nor U15781 (N_15781,N_13028,N_14112);
xor U15782 (N_15782,N_14315,N_14929);
nand U15783 (N_15783,N_15069,N_14437);
or U15784 (N_15784,N_14827,N_13704);
and U15785 (N_15785,N_14201,N_14306);
nor U15786 (N_15786,N_14282,N_14575);
nor U15787 (N_15787,N_12890,N_13891);
nor U15788 (N_15788,N_13140,N_13687);
and U15789 (N_15789,N_15448,N_13099);
nor U15790 (N_15790,N_14130,N_13888);
nor U15791 (N_15791,N_15000,N_15043);
nand U15792 (N_15792,N_13013,N_15269);
nand U15793 (N_15793,N_13396,N_13169);
and U15794 (N_15794,N_14411,N_14727);
and U15795 (N_15795,N_15484,N_14496);
or U15796 (N_15796,N_14483,N_14934);
nor U15797 (N_15797,N_13679,N_12806);
or U15798 (N_15798,N_15157,N_12877);
nor U15799 (N_15799,N_12812,N_13993);
or U15800 (N_15800,N_14438,N_14824);
and U15801 (N_15801,N_13936,N_13516);
or U15802 (N_15802,N_15005,N_14223);
or U15803 (N_15803,N_14435,N_13225);
nand U15804 (N_15804,N_12917,N_14666);
xnor U15805 (N_15805,N_12998,N_13512);
or U15806 (N_15806,N_13492,N_15497);
and U15807 (N_15807,N_14122,N_13803);
nor U15808 (N_15808,N_13525,N_13977);
xor U15809 (N_15809,N_14606,N_13287);
and U15810 (N_15810,N_13097,N_13184);
nor U15811 (N_15811,N_12631,N_14733);
and U15812 (N_15812,N_12973,N_13283);
and U15813 (N_15813,N_14429,N_14188);
nand U15814 (N_15814,N_15583,N_13041);
or U15815 (N_15815,N_12676,N_15298);
or U15816 (N_15816,N_12610,N_15180);
or U15817 (N_15817,N_13262,N_13250);
and U15818 (N_15818,N_15183,N_15251);
nand U15819 (N_15819,N_15429,N_13175);
xor U15820 (N_15820,N_15521,N_13589);
nor U15821 (N_15821,N_13912,N_14358);
nor U15822 (N_15822,N_15297,N_15502);
xor U15823 (N_15823,N_14237,N_14625);
or U15824 (N_15824,N_13347,N_13734);
nand U15825 (N_15825,N_12667,N_15240);
and U15826 (N_15826,N_13044,N_12891);
and U15827 (N_15827,N_14243,N_12726);
nand U15828 (N_15828,N_15602,N_13495);
nor U15829 (N_15829,N_13718,N_13812);
and U15830 (N_15830,N_13848,N_14975);
or U15831 (N_15831,N_15565,N_15427);
nand U15832 (N_15832,N_13572,N_15228);
nor U15833 (N_15833,N_15500,N_13575);
and U15834 (N_15834,N_13335,N_14678);
and U15835 (N_15835,N_15016,N_14427);
and U15836 (N_15836,N_15503,N_14904);
nand U15837 (N_15837,N_15418,N_14368);
nand U15838 (N_15838,N_15271,N_13456);
or U15839 (N_15839,N_15011,N_13561);
xnor U15840 (N_15840,N_13065,N_15424);
nand U15841 (N_15841,N_14096,N_12920);
nor U15842 (N_15842,N_15488,N_13590);
xnor U15843 (N_15843,N_14881,N_14428);
nor U15844 (N_15844,N_15101,N_12528);
nand U15845 (N_15845,N_13925,N_15136);
xor U15846 (N_15846,N_15222,N_14865);
and U15847 (N_15847,N_12866,N_13798);
xnor U15848 (N_15848,N_14085,N_13586);
nand U15849 (N_15849,N_14323,N_12636);
nor U15850 (N_15850,N_14912,N_14365);
or U15851 (N_15851,N_14703,N_15139);
or U15852 (N_15852,N_12635,N_15224);
nor U15853 (N_15853,N_12584,N_12686);
nand U15854 (N_15854,N_14291,N_14328);
and U15855 (N_15855,N_15428,N_13149);
or U15856 (N_15856,N_15571,N_13604);
or U15857 (N_15857,N_13595,N_12641);
or U15858 (N_15858,N_13289,N_14221);
nand U15859 (N_15859,N_14079,N_14228);
xnor U15860 (N_15860,N_13741,N_14153);
xnor U15861 (N_15861,N_13719,N_14324);
or U15862 (N_15862,N_15463,N_12503);
nand U15863 (N_15863,N_12941,N_15036);
and U15864 (N_15864,N_14651,N_14592);
or U15865 (N_15865,N_13797,N_15098);
nor U15866 (N_15866,N_14815,N_15051);
and U15867 (N_15867,N_14453,N_14773);
nor U15868 (N_15868,N_13872,N_12614);
xnor U15869 (N_15869,N_14871,N_14548);
nor U15870 (N_15870,N_13363,N_13124);
or U15871 (N_15871,N_14455,N_14259);
xor U15872 (N_15872,N_14745,N_14023);
xor U15873 (N_15873,N_14747,N_15517);
xnor U15874 (N_15874,N_14756,N_13050);
or U15875 (N_15875,N_13392,N_15121);
and U15876 (N_15876,N_15064,N_13762);
or U15877 (N_15877,N_14290,N_12512);
xor U15878 (N_15878,N_12715,N_13893);
or U15879 (N_15879,N_13954,N_15458);
and U15880 (N_15880,N_13959,N_14219);
xor U15881 (N_15881,N_14325,N_13114);
and U15882 (N_15882,N_12516,N_15310);
and U15883 (N_15883,N_13432,N_13963);
nor U15884 (N_15884,N_13781,N_15540);
or U15885 (N_15885,N_14805,N_13419);
and U15886 (N_15886,N_13272,N_14684);
or U15887 (N_15887,N_14531,N_13198);
xnor U15888 (N_15888,N_14758,N_13765);
and U15889 (N_15889,N_13986,N_14304);
xor U15890 (N_15890,N_15004,N_14843);
nand U15891 (N_15891,N_14907,N_14749);
xor U15892 (N_15892,N_13655,N_13989);
nor U15893 (N_15893,N_14610,N_13535);
nand U15894 (N_15894,N_14895,N_14519);
nand U15895 (N_15895,N_14217,N_13648);
nand U15896 (N_15896,N_15027,N_15604);
nand U15897 (N_15897,N_14891,N_13312);
or U15898 (N_15898,N_13915,N_14561);
and U15899 (N_15899,N_12502,N_15320);
xnor U15900 (N_15900,N_12569,N_14620);
nand U15901 (N_15901,N_13908,N_12984);
xor U15902 (N_15902,N_13717,N_14281);
xnor U15903 (N_15903,N_13134,N_14554);
nor U15904 (N_15904,N_12674,N_13552);
or U15905 (N_15905,N_14500,N_13506);
or U15906 (N_15906,N_13111,N_13540);
nor U15907 (N_15907,N_13564,N_12799);
nand U15908 (N_15908,N_13983,N_15417);
nand U15909 (N_15909,N_15332,N_15515);
nor U15910 (N_15910,N_14501,N_14105);
nand U15911 (N_15911,N_12952,N_14446);
and U15912 (N_15912,N_13243,N_13829);
nor U15913 (N_15913,N_14337,N_14231);
and U15914 (N_15914,N_13563,N_14064);
nor U15915 (N_15915,N_13514,N_15389);
or U15916 (N_15916,N_15203,N_12831);
and U15917 (N_15917,N_13092,N_14200);
and U15918 (N_15918,N_15076,N_13513);
or U15919 (N_15919,N_12558,N_15137);
nor U15920 (N_15920,N_14587,N_15591);
xor U15921 (N_15921,N_12607,N_13693);
and U15922 (N_15922,N_15193,N_12826);
nor U15923 (N_15923,N_14535,N_13645);
nor U15924 (N_15924,N_14588,N_15566);
nor U15925 (N_15925,N_13821,N_14378);
nor U15926 (N_15926,N_14999,N_13505);
or U15927 (N_15927,N_15214,N_13774);
and U15928 (N_15928,N_13219,N_13583);
nor U15929 (N_15929,N_15363,N_14809);
xnor U15930 (N_15930,N_14212,N_13245);
or U15931 (N_15931,N_13542,N_15411);
xnor U15932 (N_15932,N_14783,N_13735);
or U15933 (N_15933,N_15386,N_14537);
and U15934 (N_15934,N_12677,N_15416);
nand U15935 (N_15935,N_15531,N_13389);
and U15936 (N_15936,N_12637,N_14641);
and U15937 (N_15937,N_13814,N_14810);
or U15938 (N_15938,N_14700,N_12560);
nand U15939 (N_15939,N_14726,N_15163);
and U15940 (N_15940,N_13026,N_12972);
and U15941 (N_15941,N_13402,N_13509);
nand U15942 (N_15942,N_14468,N_12580);
nor U15943 (N_15943,N_13897,N_13275);
nand U15944 (N_15944,N_14179,N_13546);
or U15945 (N_15945,N_14399,N_14367);
nor U15946 (N_15946,N_12749,N_14308);
xor U15947 (N_15947,N_13253,N_12652);
nor U15948 (N_15948,N_14329,N_14345);
or U15949 (N_15949,N_14844,N_12978);
nand U15950 (N_15950,N_12969,N_12994);
and U15951 (N_15951,N_14473,N_13608);
and U15952 (N_15952,N_13852,N_15278);
or U15953 (N_15953,N_14441,N_14772);
xor U15954 (N_15954,N_12804,N_13520);
and U15955 (N_15955,N_14014,N_14471);
nor U15956 (N_15956,N_13268,N_14195);
xnor U15957 (N_15957,N_14662,N_13014);
nor U15958 (N_15958,N_12778,N_14470);
and U15959 (N_15959,N_12595,N_15159);
or U15960 (N_15960,N_13632,N_13429);
or U15961 (N_15961,N_14129,N_15091);
and U15962 (N_15962,N_14340,N_12723);
xor U15963 (N_15963,N_13183,N_15430);
or U15964 (N_15964,N_14370,N_12999);
nor U15965 (N_15965,N_13733,N_13457);
nand U15966 (N_15966,N_13355,N_14284);
and U15967 (N_15967,N_15245,N_14759);
nor U15968 (N_15968,N_12795,N_13005);
xor U15969 (N_15969,N_12644,N_13136);
xor U15970 (N_15970,N_14364,N_14654);
xnor U15971 (N_15971,N_12820,N_15265);
nor U15972 (N_15972,N_12990,N_14754);
and U15973 (N_15973,N_13214,N_13381);
nor U15974 (N_15974,N_14511,N_12781);
nor U15975 (N_15975,N_13935,N_14351);
nand U15976 (N_15976,N_12609,N_14033);
nand U15977 (N_15977,N_15551,N_13971);
or U15978 (N_15978,N_12698,N_12603);
and U15979 (N_15979,N_12514,N_14283);
or U15980 (N_15980,N_13417,N_13692);
nand U15981 (N_15981,N_12733,N_13864);
or U15982 (N_15982,N_14480,N_15044);
nand U15983 (N_15983,N_14863,N_14037);
or U15984 (N_15984,N_14746,N_14056);
xor U15985 (N_15985,N_13967,N_13837);
nand U15986 (N_15986,N_13955,N_14743);
nand U15987 (N_15987,N_14106,N_14959);
nand U15988 (N_15988,N_12505,N_15223);
nor U15989 (N_15989,N_15274,N_14158);
nor U15990 (N_15990,N_12983,N_13163);
nand U15991 (N_15991,N_13773,N_14265);
or U15992 (N_15992,N_15315,N_14857);
or U15993 (N_15993,N_15616,N_13614);
or U15994 (N_15994,N_13370,N_12763);
nand U15995 (N_15995,N_14230,N_13602);
xnor U15996 (N_15996,N_14960,N_15623);
xor U15997 (N_15997,N_13448,N_15525);
nand U15998 (N_15998,N_13988,N_12912);
xnor U15999 (N_15999,N_15498,N_12814);
or U16000 (N_16000,N_13333,N_15490);
nor U16001 (N_16001,N_15581,N_13058);
nor U16002 (N_16002,N_13462,N_13676);
or U16003 (N_16003,N_14344,N_14080);
or U16004 (N_16004,N_14714,N_14178);
nand U16005 (N_16005,N_13106,N_15436);
nor U16006 (N_16006,N_14917,N_12670);
nor U16007 (N_16007,N_12851,N_13004);
and U16008 (N_16008,N_12791,N_14981);
nand U16009 (N_16009,N_15066,N_13771);
xnor U16010 (N_16010,N_14199,N_12964);
or U16011 (N_16011,N_13182,N_15049);
xor U16012 (N_16012,N_13532,N_15096);
or U16013 (N_16013,N_14003,N_13965);
and U16014 (N_16014,N_15208,N_13095);
xnor U16015 (N_16015,N_15617,N_13410);
nor U16016 (N_16016,N_15321,N_14327);
xor U16017 (N_16017,N_14638,N_15070);
and U16018 (N_16018,N_15021,N_12617);
xnor U16019 (N_16019,N_14257,N_12679);
xor U16020 (N_16020,N_13481,N_13633);
nor U16021 (N_16021,N_12571,N_12828);
nor U16022 (N_16022,N_13623,N_14868);
or U16023 (N_16023,N_13420,N_13414);
xnor U16024 (N_16024,N_13899,N_14396);
or U16025 (N_16025,N_15094,N_13145);
nand U16026 (N_16026,N_15100,N_13887);
nor U16027 (N_16027,N_12907,N_15355);
nor U16028 (N_16028,N_12700,N_12697);
xor U16029 (N_16029,N_15175,N_14333);
or U16030 (N_16030,N_14494,N_13424);
nand U16031 (N_16031,N_12622,N_14187);
nor U16032 (N_16032,N_13466,N_14142);
nor U16033 (N_16033,N_12929,N_15155);
or U16034 (N_16034,N_13430,N_14639);
and U16035 (N_16035,N_14689,N_15348);
and U16036 (N_16036,N_13139,N_13686);
xnor U16037 (N_16037,N_15494,N_13851);
or U16038 (N_16038,N_15618,N_14036);
nor U16039 (N_16039,N_12764,N_13385);
nor U16040 (N_16040,N_13806,N_14287);
and U16041 (N_16041,N_15400,N_13056);
or U16042 (N_16042,N_12611,N_14309);
and U16043 (N_16043,N_15557,N_12665);
or U16044 (N_16044,N_15572,N_13240);
and U16045 (N_16045,N_14655,N_12663);
xnor U16046 (N_16046,N_15152,N_12661);
or U16047 (N_16047,N_12892,N_15541);
nand U16048 (N_16048,N_12816,N_14504);
xnor U16049 (N_16049,N_12721,N_12903);
nor U16050 (N_16050,N_13581,N_13295);
or U16051 (N_16051,N_14649,N_13500);
nor U16052 (N_16052,N_13384,N_13856);
xnor U16053 (N_16053,N_12675,N_14108);
nor U16054 (N_16054,N_13968,N_14078);
nand U16055 (N_16055,N_15063,N_13779);
nor U16056 (N_16056,N_14070,N_14288);
or U16057 (N_16057,N_12710,N_14883);
or U16058 (N_16058,N_13539,N_13059);
nor U16059 (N_16059,N_12754,N_12691);
and U16060 (N_16060,N_14921,N_12813);
xor U16061 (N_16061,N_12669,N_15439);
nand U16062 (N_16062,N_14634,N_15034);
nand U16063 (N_16063,N_13388,N_13413);
nor U16064 (N_16064,N_14586,N_14788);
and U16065 (N_16065,N_13880,N_13528);
or U16066 (N_16066,N_15048,N_14628);
or U16067 (N_16067,N_12807,N_13533);
nor U16068 (N_16068,N_14608,N_12784);
or U16069 (N_16069,N_13665,N_14041);
xnor U16070 (N_16070,N_14925,N_15485);
or U16071 (N_16071,N_14543,N_15077);
and U16072 (N_16072,N_15267,N_14100);
or U16073 (N_16073,N_14251,N_15384);
nor U16074 (N_16074,N_14763,N_12953);
nand U16075 (N_16075,N_15622,N_13593);
or U16076 (N_16076,N_13016,N_14366);
or U16077 (N_16077,N_15349,N_13494);
nand U16078 (N_16078,N_14677,N_14799);
nand U16079 (N_16079,N_15206,N_14401);
nor U16080 (N_16080,N_14464,N_13033);
or U16081 (N_16081,N_13716,N_13434);
nor U16082 (N_16082,N_13913,N_13437);
xor U16083 (N_16083,N_15329,N_13511);
and U16084 (N_16084,N_12780,N_13637);
nor U16085 (N_16085,N_12906,N_14409);
and U16086 (N_16086,N_12575,N_13951);
and U16087 (N_16087,N_14529,N_15431);
nor U16088 (N_16088,N_14850,N_14139);
xnor U16089 (N_16089,N_13952,N_13387);
and U16090 (N_16090,N_13337,N_13715);
or U16091 (N_16091,N_13342,N_14695);
or U16092 (N_16092,N_12752,N_14600);
and U16093 (N_16093,N_14965,N_13085);
nor U16094 (N_16094,N_13091,N_13950);
or U16095 (N_16095,N_12989,N_14215);
or U16096 (N_16096,N_14155,N_13193);
nor U16097 (N_16097,N_14701,N_14109);
nand U16098 (N_16098,N_14757,N_13909);
and U16099 (N_16099,N_13650,N_15162);
nor U16100 (N_16100,N_15556,N_15268);
or U16101 (N_16101,N_12800,N_13990);
and U16102 (N_16102,N_13757,N_14922);
nand U16103 (N_16103,N_12787,N_14102);
xor U16104 (N_16104,N_13423,N_13019);
nor U16105 (N_16105,N_14157,N_14152);
or U16106 (N_16106,N_14945,N_12948);
nor U16107 (N_16107,N_14225,N_13201);
xor U16108 (N_16108,N_13543,N_13195);
and U16109 (N_16109,N_13159,N_14256);
xor U16110 (N_16110,N_13927,N_14415);
or U16111 (N_16111,N_14138,N_13017);
xnor U16112 (N_16112,N_13991,N_12913);
or U16113 (N_16113,N_12779,N_13914);
and U16114 (N_16114,N_14766,N_14088);
and U16115 (N_16115,N_14982,N_13619);
or U16116 (N_16116,N_14162,N_13673);
xor U16117 (N_16117,N_13850,N_14376);
xnor U16118 (N_16118,N_14597,N_15402);
or U16119 (N_16119,N_12654,N_15512);
or U16120 (N_16120,N_12775,N_15560);
or U16121 (N_16121,N_13522,N_14132);
xor U16122 (N_16122,N_13164,N_14838);
nor U16123 (N_16123,N_14616,N_12860);
nand U16124 (N_16124,N_13435,N_13728);
and U16125 (N_16125,N_14576,N_14424);
nor U16126 (N_16126,N_13588,N_13246);
and U16127 (N_16127,N_12918,N_15302);
or U16128 (N_16128,N_15218,N_12740);
or U16129 (N_16129,N_14035,N_12773);
or U16130 (N_16130,N_12511,N_12600);
nor U16131 (N_16131,N_12884,N_15606);
xor U16132 (N_16132,N_14910,N_14855);
nand U16133 (N_16133,N_13365,N_15535);
nand U16134 (N_16134,N_13334,N_14027);
nor U16135 (N_16135,N_12815,N_13055);
nor U16136 (N_16136,N_13035,N_12729);
nand U16137 (N_16137,N_15520,N_13671);
xor U16138 (N_16138,N_13087,N_15605);
nor U16139 (N_16139,N_15519,N_14569);
or U16140 (N_16140,N_15381,N_13051);
xor U16141 (N_16141,N_12872,N_13775);
nand U16142 (N_16142,N_14104,N_13764);
xor U16143 (N_16143,N_15133,N_15241);
and U16144 (N_16144,N_14440,N_15481);
nand U16145 (N_16145,N_13553,N_15586);
nor U16146 (N_16146,N_12620,N_15499);
xor U16147 (N_16147,N_13267,N_13981);
or U16148 (N_16148,N_13700,N_13544);
or U16149 (N_16149,N_13249,N_15339);
nand U16150 (N_16150,N_14211,N_12666);
or U16151 (N_16151,N_15052,N_13922);
or U16152 (N_16152,N_15154,N_13636);
and U16153 (N_16153,N_14833,N_14042);
or U16154 (N_16154,N_12685,N_14970);
xor U16155 (N_16155,N_14029,N_12761);
and U16156 (N_16156,N_13801,N_12772);
or U16157 (N_16157,N_14900,N_12541);
nor U16158 (N_16158,N_12762,N_14202);
nand U16159 (N_16159,N_14964,N_14000);
and U16160 (N_16160,N_14154,N_15219);
or U16161 (N_16161,N_15595,N_13296);
nor U16162 (N_16162,N_12982,N_14709);
xor U16163 (N_16163,N_12657,N_12659);
nand U16164 (N_16164,N_14528,N_14571);
nor U16165 (N_16165,N_15473,N_13074);
nand U16166 (N_16166,N_15112,N_13233);
nand U16167 (N_16167,N_14527,N_13631);
and U16168 (N_16168,N_14878,N_13144);
nor U16169 (N_16169,N_14564,N_15388);
or U16170 (N_16170,N_14508,N_12845);
xor U16171 (N_16171,N_13230,N_13873);
and U16172 (N_16172,N_15412,N_12529);
nand U16173 (N_16173,N_15372,N_13234);
and U16174 (N_16174,N_15151,N_12934);
nor U16175 (N_16175,N_12653,N_14604);
and U16176 (N_16176,N_12844,N_12577);
nor U16177 (N_16177,N_13618,N_13446);
xnor U16178 (N_16178,N_14842,N_14009);
nand U16179 (N_16179,N_14880,N_13323);
or U16180 (N_16180,N_14623,N_15285);
and U16181 (N_16181,N_15086,N_15446);
and U16182 (N_16182,N_14831,N_13465);
and U16183 (N_16183,N_12701,N_12753);
nand U16184 (N_16184,N_13732,N_14968);
nor U16185 (N_16185,N_13088,N_14692);
nor U16186 (N_16186,N_13607,N_13625);
and U16187 (N_16187,N_15263,N_15472);
or U16188 (N_16188,N_15194,N_12728);
nand U16189 (N_16189,N_14661,N_15374);
xnor U16190 (N_16190,N_13792,N_14755);
or U16191 (N_16191,N_14807,N_14417);
xnor U16192 (N_16192,N_13763,N_15338);
and U16193 (N_16193,N_15530,N_13600);
xor U16194 (N_16194,N_13366,N_12940);
nor U16195 (N_16195,N_14867,N_15317);
and U16196 (N_16196,N_14332,N_14206);
nand U16197 (N_16197,N_13354,N_13131);
xnor U16198 (N_16198,N_13181,N_14598);
nor U16199 (N_16199,N_14343,N_14076);
nor U16200 (N_16200,N_12991,N_13079);
nor U16201 (N_16201,N_13871,N_15253);
nor U16202 (N_16202,N_13556,N_12894);
xor U16203 (N_16203,N_14083,N_13978);
or U16204 (N_16204,N_12895,N_12959);
xnor U16205 (N_16205,N_13937,N_14238);
nand U16206 (N_16206,N_14456,N_12896);
nor U16207 (N_16207,N_12974,N_15449);
and U16208 (N_16208,N_13726,N_14717);
nor U16209 (N_16209,N_13362,N_12722);
and U16210 (N_16210,N_15182,N_12809);
nand U16211 (N_16211,N_14404,N_13428);
nand U16212 (N_16212,N_14374,N_13105);
or U16213 (N_16213,N_13573,N_14901);
nand U16214 (N_16214,N_13597,N_15248);
nand U16215 (N_16215,N_14434,N_15435);
or U16216 (N_16216,N_14224,N_15397);
or U16217 (N_16217,N_13176,N_12975);
and U16218 (N_16218,N_14522,N_14905);
nor U16219 (N_16219,N_13835,N_12794);
nor U16220 (N_16220,N_14736,N_13723);
and U16221 (N_16221,N_13216,N_14516);
xnor U16222 (N_16222,N_12846,N_13314);
xnor U16223 (N_16223,N_13304,N_14353);
nand U16224 (N_16224,N_14558,N_14071);
and U16225 (N_16225,N_13301,N_15165);
nor U16226 (N_16226,N_15153,N_14408);
xnor U16227 (N_16227,N_12801,N_14478);
nand U16228 (N_16228,N_14118,N_15191);
xor U16229 (N_16229,N_14172,N_14059);
nor U16230 (N_16230,N_15161,N_12738);
nor U16231 (N_16231,N_13439,N_13209);
and U16232 (N_16232,N_15326,N_14702);
nor U16233 (N_16233,N_15495,N_13223);
nand U16234 (N_16234,N_13906,N_13197);
nor U16235 (N_16235,N_12915,N_13158);
or U16236 (N_16236,N_15456,N_13433);
nor U16237 (N_16237,N_13461,N_14356);
and U16238 (N_16238,N_13269,N_13211);
or U16239 (N_16239,N_14075,N_15038);
xnor U16240 (N_16240,N_14476,N_12619);
xor U16241 (N_16241,N_12898,N_14646);
xor U16242 (N_16242,N_15466,N_14979);
and U16243 (N_16243,N_12605,N_13566);
xor U16244 (N_16244,N_15244,N_15065);
nand U16245 (N_16245,N_14270,N_14957);
nand U16246 (N_16246,N_12857,N_13321);
nor U16247 (N_16247,N_14941,N_15442);
nor U16248 (N_16248,N_13190,N_15489);
or U16249 (N_16249,N_14253,N_14862);
and U16250 (N_16250,N_14706,N_15453);
xnor U16251 (N_16251,N_13591,N_13155);
or U16252 (N_16252,N_14864,N_14650);
nor U16253 (N_16253,N_12797,N_13098);
or U16254 (N_16254,N_14542,N_12925);
and U16255 (N_16255,N_15095,N_12707);
or U16256 (N_16256,N_13213,N_15188);
and U16257 (N_16257,N_13752,N_14311);
and U16258 (N_16258,N_14039,N_13386);
or U16259 (N_16259,N_14119,N_13046);
nand U16260 (N_16260,N_12885,N_13394);
nand U16261 (N_16261,N_15190,N_12827);
xnor U16262 (N_16262,N_15536,N_14980);
and U16263 (N_16263,N_15620,N_14412);
or U16264 (N_16264,N_12551,N_13086);
nand U16265 (N_16265,N_15196,N_13029);
nand U16266 (N_16266,N_14741,N_12868);
nand U16267 (N_16267,N_14389,N_15025);
and U16268 (N_16268,N_15461,N_14159);
and U16269 (N_16269,N_12519,N_13319);
or U16270 (N_16270,N_14025,N_13358);
nand U16271 (N_16271,N_12832,N_14241);
xor U16272 (N_16272,N_13787,N_14385);
nor U16273 (N_16273,N_13710,N_15259);
xnor U16274 (N_16274,N_14590,N_13263);
nand U16275 (N_16275,N_12594,N_13836);
nand U16276 (N_16276,N_15061,N_14919);
and U16277 (N_16277,N_14835,N_13875);
nand U16278 (N_16278,N_14019,N_15546);
xnor U16279 (N_16279,N_15385,N_15547);
and U16280 (N_16280,N_14787,N_14540);
xor U16281 (N_16281,N_13724,N_13657);
or U16282 (N_16282,N_13789,N_13992);
or U16283 (N_16283,N_14681,N_13081);
nand U16284 (N_16284,N_12696,N_14939);
and U16285 (N_16285,N_12817,N_14988);
and U16286 (N_16286,N_13043,N_15083);
nor U16287 (N_16287,N_15072,N_14992);
nand U16288 (N_16288,N_13638,N_13818);
nand U16289 (N_16289,N_13426,N_14653);
nand U16290 (N_16290,N_14107,N_14873);
nor U16291 (N_16291,N_13568,N_15323);
or U16292 (N_16292,N_13045,N_12935);
nand U16293 (N_16293,N_13020,N_15007);
and U16294 (N_16294,N_14151,N_14682);
nor U16295 (N_16295,N_12871,N_14216);
or U16296 (N_16296,N_14254,N_14047);
xor U16297 (N_16297,N_15090,N_15258);
and U16298 (N_16298,N_14320,N_12852);
nor U16299 (N_16299,N_15020,N_15358);
or U16300 (N_16300,N_15147,N_13518);
xnor U16301 (N_16301,N_13248,N_14720);
xnor U16302 (N_16302,N_14156,N_13459);
nand U16303 (N_16303,N_14447,N_14321);
nand U16304 (N_16304,N_14262,N_13761);
and U16305 (N_16305,N_15452,N_14595);
nand U16306 (N_16306,N_15211,N_15352);
nor U16307 (N_16307,N_13449,N_13832);
and U16308 (N_16308,N_15176,N_15131);
or U16309 (N_16309,N_15236,N_15598);
nand U16310 (N_16310,N_14596,N_14169);
and U16311 (N_16311,N_14593,N_15111);
and U16312 (N_16312,N_14095,N_13907);
xnor U16313 (N_16313,N_12955,N_14084);
nor U16314 (N_16314,N_14567,N_15469);
xor U16315 (N_16315,N_15266,N_13788);
nand U16316 (N_16316,N_15334,N_15361);
nor U16317 (N_16317,N_13048,N_13599);
and U16318 (N_16318,N_12638,N_13063);
and U16319 (N_16319,N_15158,N_13854);
xor U16320 (N_16320,N_14026,N_15088);
nand U16321 (N_16321,N_14189,N_12650);
nand U16322 (N_16322,N_13611,N_14004);
xor U16323 (N_16323,N_13006,N_12730);
nand U16324 (N_16324,N_13427,N_14444);
xnor U16325 (N_16325,N_13270,N_13748);
nor U16326 (N_16326,N_12919,N_13403);
nor U16327 (N_16327,N_12905,N_14196);
nand U16328 (N_16328,N_15082,N_13758);
xor U16329 (N_16329,N_14630,N_13808);
nor U16330 (N_16330,N_12938,N_14821);
and U16331 (N_16331,N_14830,N_15233);
and U16332 (N_16332,N_14814,N_13212);
nand U16333 (N_16333,N_12690,N_15146);
nor U16334 (N_16334,N_14279,N_13003);
xnor U16335 (N_16335,N_15523,N_15199);
and U16336 (N_16336,N_13293,N_14920);
nand U16337 (N_16337,N_15392,N_15440);
and U16338 (N_16338,N_15406,N_12767);
xnor U16339 (N_16339,N_13994,N_12694);
xnor U16340 (N_16340,N_14930,N_12567);
nand U16341 (N_16341,N_14260,N_15433);
and U16342 (N_16342,N_15078,N_14208);
and U16343 (N_16343,N_12849,N_12513);
nor U16344 (N_16344,N_13147,N_14552);
or U16345 (N_16345,N_14619,N_15031);
xor U16346 (N_16346,N_13876,N_15242);
or U16347 (N_16347,N_12587,N_14297);
and U16348 (N_16348,N_14674,N_13578);
xor U16349 (N_16349,N_14675,N_14485);
and U16350 (N_16350,N_13467,N_13903);
and U16351 (N_16351,N_14301,N_12618);
nand U16352 (N_16352,N_15423,N_12976);
xnor U16353 (N_16353,N_14069,N_14851);
and U16354 (N_16354,N_13738,N_12612);
or U16355 (N_16355,N_14698,N_13675);
nor U16356 (N_16356,N_14730,N_14591);
or U16357 (N_16357,N_15584,N_13142);
nand U16358 (N_16358,N_15296,N_13450);
nand U16359 (N_16359,N_13622,N_13527);
and U16360 (N_16360,N_14601,N_14915);
and U16361 (N_16361,N_13554,N_15023);
nor U16362 (N_16362,N_13911,N_13931);
nor U16363 (N_16363,N_12838,N_14081);
nand U16364 (N_16364,N_14668,N_12899);
and U16365 (N_16365,N_14927,N_14050);
or U16366 (N_16366,N_13881,N_13179);
xnor U16367 (N_16367,N_13928,N_12586);
nor U16368 (N_16368,N_12702,N_15396);
or U16369 (N_16369,N_15122,N_12573);
nand U16370 (N_16370,N_15080,N_14777);
nor U16371 (N_16371,N_13691,N_15264);
or U16372 (N_16372,N_15003,N_12744);
or U16373 (N_16373,N_13218,N_15395);
and U16374 (N_16374,N_15212,N_13236);
xor U16375 (N_16375,N_14679,N_15026);
nor U16376 (N_16376,N_13652,N_14082);
or U16377 (N_16377,N_15316,N_14911);
or U16378 (N_16378,N_12572,N_13431);
nand U16379 (N_16379,N_14711,N_13330);
xnor U16380 (N_16380,N_15149,N_13156);
xor U16381 (N_16381,N_14562,N_15134);
or U16382 (N_16382,N_13485,N_14780);
or U16383 (N_16383,N_13972,N_14602);
and U16384 (N_16384,N_14336,N_13833);
and U16385 (N_16385,N_13277,N_13480);
and U16386 (N_16386,N_13956,N_14264);
nor U16387 (N_16387,N_13910,N_12509);
xnor U16388 (N_16388,N_14252,N_13783);
xor U16389 (N_16389,N_13879,N_15478);
nand U16390 (N_16390,N_13714,N_14317);
nor U16391 (N_16391,N_13501,N_14135);
nor U16392 (N_16392,N_13104,N_14489);
or U16393 (N_16393,N_14987,N_13576);
nand U16394 (N_16394,N_13537,N_14218);
or U16395 (N_16395,N_13438,N_15301);
nor U16396 (N_16396,N_12709,N_15017);
nand U16397 (N_16397,N_14165,N_12943);
or U16398 (N_16398,N_15342,N_15056);
or U16399 (N_16399,N_12870,N_13242);
or U16400 (N_16400,N_12841,N_13476);
nor U16401 (N_16401,N_12500,N_13550);
nor U16402 (N_16402,N_13229,N_13807);
and U16403 (N_16403,N_15425,N_15075);
and U16404 (N_16404,N_15518,N_15012);
or U16405 (N_16405,N_14737,N_12944);
nor U16406 (N_16406,N_14466,N_13310);
and U16407 (N_16407,N_12986,N_13942);
xnor U16408 (N_16408,N_13499,N_13300);
or U16409 (N_16409,N_15128,N_14973);
or U16410 (N_16410,N_14207,N_14463);
nand U16411 (N_16411,N_14952,N_13776);
nor U16412 (N_16412,N_12501,N_14044);
nor U16413 (N_16413,N_15553,N_13360);
and U16414 (N_16414,N_13778,N_14949);
and U16415 (N_16415,N_13750,N_14914);
xor U16416 (N_16416,N_14645,N_13082);
nor U16417 (N_16417,N_15047,N_14715);
or U16418 (N_16418,N_14823,N_13228);
nor U16419 (N_16419,N_14477,N_15014);
and U16420 (N_16420,N_14665,N_12591);
and U16421 (N_16421,N_13348,N_13660);
nand U16422 (N_16422,N_15609,N_13397);
or U16423 (N_16423,N_14185,N_12874);
nor U16424 (N_16424,N_14359,N_14166);
nand U16425 (N_16425,N_14018,N_15567);
and U16426 (N_16426,N_14642,N_14797);
xor U16427 (N_16427,N_13421,N_15380);
xnor U16428 (N_16428,N_14770,N_15001);
nand U16429 (N_16429,N_13708,N_13641);
or U16430 (N_16430,N_14874,N_15015);
or U16431 (N_16431,N_13721,N_14233);
and U16432 (N_16432,N_12554,N_15539);
xor U16433 (N_16433,N_12995,N_12506);
nor U16434 (N_16434,N_15327,N_12693);
nor U16435 (N_16435,N_15561,N_14719);
and U16436 (N_16436,N_13084,N_12981);
xnor U16437 (N_16437,N_12527,N_14379);
or U16438 (N_16438,N_12865,N_13727);
or U16439 (N_16439,N_15607,N_15257);
xnor U16440 (N_16440,N_13547,N_14846);
xor U16441 (N_16441,N_15107,N_12678);
xor U16442 (N_16442,N_14618,N_13146);
and U16443 (N_16443,N_14051,N_14285);
and U16444 (N_16444,N_12985,N_13565);
and U16445 (N_16445,N_12880,N_13024);
nor U16446 (N_16446,N_13407,N_15364);
nor U16447 (N_16447,N_14295,N_13811);
nand U16448 (N_16448,N_13007,N_15198);
and U16449 (N_16449,N_15596,N_14924);
or U16450 (N_16450,N_13038,N_14394);
and U16451 (N_16451,N_13094,N_13064);
nor U16452 (N_16452,N_14768,N_13487);
nor U16453 (N_16453,N_15370,N_13472);
or U16454 (N_16454,N_14875,N_14704);
nand U16455 (N_16455,N_14688,N_12786);
and U16456 (N_16456,N_15538,N_13115);
or U16457 (N_16457,N_14335,N_14375);
and U16458 (N_16458,N_14676,N_13866);
xor U16459 (N_16459,N_14538,N_15506);
nand U16460 (N_16460,N_14559,N_14120);
xor U16461 (N_16461,N_15563,N_12727);
nand U16462 (N_16462,N_12823,N_12660);
xor U16463 (N_16463,N_14136,N_14547);
nor U16464 (N_16464,N_12649,N_12792);
xor U16465 (N_16465,N_14950,N_14580);
nor U16466 (N_16466,N_12658,N_14232);
or U16467 (N_16467,N_15371,N_15345);
xor U16468 (N_16468,N_13180,N_14976);
nand U16469 (N_16469,N_15621,N_13702);
or U16470 (N_16470,N_14574,N_12965);
and U16471 (N_16471,N_15552,N_14330);
and U16472 (N_16472,N_15110,N_15405);
nor U16473 (N_16473,N_13343,N_12672);
xor U16474 (N_16474,N_13868,N_15197);
nand U16475 (N_16475,N_12927,N_13009);
and U16476 (N_16476,N_13995,N_13352);
xor U16477 (N_16477,N_12555,N_13884);
nand U16478 (N_16478,N_13877,N_12540);
nand U16479 (N_16479,N_14903,N_13271);
and U16480 (N_16480,N_15230,N_14406);
nand U16481 (N_16481,N_14557,N_13336);
or U16482 (N_16482,N_15099,N_12951);
or U16483 (N_16483,N_14486,N_14013);
xnor U16484 (N_16484,N_15513,N_12993);
or U16485 (N_16485,N_13672,N_12647);
or U16486 (N_16486,N_13227,N_12583);
or U16487 (N_16487,N_14390,N_14685);
and U16488 (N_16488,N_14097,N_15543);
xor U16489 (N_16489,N_14391,N_14247);
or U16490 (N_16490,N_13120,N_13025);
or U16491 (N_16491,N_15252,N_14826);
nor U16492 (N_16492,N_13627,N_13345);
xnor U16493 (N_16493,N_13130,N_15295);
nor U16494 (N_16494,N_15496,N_13766);
xnor U16495 (N_16495,N_14789,N_14007);
nor U16496 (N_16496,N_13265,N_15035);
and U16497 (N_16497,N_15294,N_13647);
or U16498 (N_16498,N_14460,N_13722);
or U16499 (N_16499,N_12921,N_13559);
nor U16500 (N_16500,N_12746,N_15116);
or U16501 (N_16501,N_15282,N_12805);
and U16502 (N_16502,N_14782,N_14061);
and U16503 (N_16503,N_15229,N_13782);
and U16504 (N_16504,N_15367,N_14128);
xor U16505 (N_16505,N_12888,N_14658);
nor U16506 (N_16506,N_14250,N_12793);
or U16507 (N_16507,N_14906,N_15032);
nor U16508 (N_16508,N_13453,N_14294);
and U16509 (N_16509,N_14180,N_15050);
and U16510 (N_16510,N_12643,N_13557);
nor U16511 (N_16511,N_14718,N_14277);
or U16512 (N_16512,N_13274,N_13479);
or U16513 (N_16513,N_15120,N_14546);
xor U16514 (N_16514,N_14859,N_13371);
nor U16515 (N_16515,N_14452,N_15105);
nor U16516 (N_16516,N_13961,N_13309);
xnor U16517 (N_16517,N_14488,N_15166);
or U16518 (N_16518,N_14407,N_14672);
nand U16519 (N_16519,N_14457,N_14487);
nor U16520 (N_16520,N_12613,N_13842);
and U16521 (N_16521,N_13210,N_15213);
xnor U16522 (N_16522,N_14150,N_13957);
nor U16523 (N_16523,N_13235,N_14779);
or U16524 (N_16524,N_14963,N_13316);
or U16525 (N_16525,N_12510,N_13662);
nor U16526 (N_16526,N_13444,N_13667);
xnor U16527 (N_16527,N_15087,N_15246);
and U16528 (N_16528,N_15273,N_15055);
nand U16529 (N_16529,N_14933,N_12854);
xnor U16530 (N_16530,N_13101,N_13497);
xnor U16531 (N_16531,N_13121,N_15603);
and U16532 (N_16532,N_12515,N_12632);
nand U16533 (N_16533,N_13206,N_15359);
or U16534 (N_16534,N_15375,N_13356);
nand U16535 (N_16535,N_14555,N_13890);
and U16536 (N_16536,N_12789,N_13830);
xor U16537 (N_16537,N_15376,N_15576);
nand U16538 (N_16538,N_14341,N_12833);
nand U16539 (N_16539,N_14380,N_13241);
nor U16540 (N_16540,N_13285,N_14998);
nand U16541 (N_16541,N_14889,N_14475);
nand U16542 (N_16542,N_12957,N_13634);
and U16543 (N_16543,N_12521,N_12768);
xor U16544 (N_16544,N_14005,N_14024);
or U16545 (N_16545,N_13047,N_14578);
nor U16546 (N_16546,N_15054,N_12830);
or U16547 (N_16547,N_15447,N_15300);
or U16548 (N_16548,N_12538,N_12742);
nor U16549 (N_16549,N_13189,N_15256);
nor U16550 (N_16550,N_15413,N_12552);
nor U16551 (N_16551,N_13464,N_14214);
or U16552 (N_16552,N_13713,N_15577);
and U16553 (N_16553,N_14643,N_13137);
xor U16554 (N_16554,N_14545,N_14182);
nand U16555 (N_16555,N_14467,N_14731);
nor U16556 (N_16556,N_13649,N_12671);
nor U16557 (N_16557,N_15178,N_13282);
nand U16558 (N_16558,N_12576,N_12687);
xnor U16559 (N_16559,N_14656,N_15575);
xor U16560 (N_16560,N_14808,N_13469);
or U16561 (N_16561,N_13739,N_13549);
nor U16562 (N_16562,N_12853,N_12534);
and U16563 (N_16563,N_14953,N_14034);
or U16564 (N_16564,N_12977,N_14204);
nand U16565 (N_16565,N_15568,N_12543);
nor U16566 (N_16566,N_15314,N_13162);
or U16567 (N_16567,N_15398,N_13658);
and U16568 (N_16568,N_14053,N_12705);
nor U16569 (N_16569,N_13601,N_13582);
xnor U16570 (N_16570,N_14414,N_13508);
or U16571 (N_16571,N_13697,N_12673);
xor U16572 (N_16572,N_14313,N_12550);
nand U16573 (N_16573,N_14570,N_13523);
or U16574 (N_16574,N_14869,N_14803);
and U16575 (N_16575,N_13820,N_12589);
or U16576 (N_16576,N_13690,N_14893);
nor U16577 (N_16577,N_15368,N_14994);
nand U16578 (N_16578,N_15476,N_15524);
nand U16579 (N_16579,N_15528,N_12623);
xnor U16580 (N_16580,N_12731,N_14381);
nor U16581 (N_16581,N_14292,N_13373);
and U16582 (N_16582,N_15504,N_12939);
and U16583 (N_16583,N_13754,N_13377);
nand U16584 (N_16584,N_15097,N_12602);
nand U16585 (N_16585,N_14892,N_13422);
nor U16586 (N_16586,N_14094,N_14269);
nor U16587 (N_16587,N_15304,N_14722);
nand U16588 (N_16588,N_12585,N_15592);
nor U16589 (N_16589,N_13976,N_14073);
or U16590 (N_16590,N_13496,N_14621);
nor U16591 (N_16591,N_14192,N_13933);
nor U16592 (N_16592,N_14350,N_14439);
and U16593 (N_16593,N_13680,N_14131);
or U16594 (N_16594,N_14644,N_14314);
nand U16595 (N_16595,N_15201,N_13939);
xnor U16596 (N_16596,N_13839,N_13869);
xnor U16597 (N_16597,N_12545,N_15331);
nor U16598 (N_16598,N_15286,N_15231);
nor U16599 (N_16599,N_12810,N_15341);
xor U16600 (N_16600,N_14183,N_14967);
or U16601 (N_16601,N_13571,N_15600);
nor U16602 (N_16602,N_13141,N_12992);
xnor U16603 (N_16603,N_13793,N_13862);
nand U16604 (N_16604,N_12524,N_14031);
nor U16605 (N_16605,N_13669,N_14001);
nor U16606 (N_16606,N_14349,N_14767);
nor U16607 (N_16607,N_13203,N_13329);
nand U16608 (N_16608,N_13185,N_14175);
or U16609 (N_16609,N_15216,N_13068);
nand U16610 (N_16610,N_15373,N_12549);
nand U16611 (N_16611,N_15309,N_15117);
or U16612 (N_16612,N_14261,N_13570);
xnor U16613 (N_16613,N_14479,N_14093);
and U16614 (N_16614,N_13478,N_14267);
and U16615 (N_16615,N_15171,N_15580);
nand U16616 (N_16616,N_15404,N_14331);
nor U16617 (N_16617,N_15192,N_15220);
nor U16618 (N_16618,N_15579,N_14886);
nand U16619 (N_16619,N_15534,N_14249);
nor U16620 (N_16620,N_14854,N_13122);
and U16621 (N_16621,N_13266,N_13883);
xor U16622 (N_16622,N_12601,N_13736);
or U16623 (N_16623,N_14802,N_13237);
or U16624 (N_16624,N_12883,N_13859);
and U16625 (N_16625,N_14091,N_13102);
xnor U16626 (N_16626,N_15243,N_13313);
and U16627 (N_16627,N_13173,N_15573);
nor U16628 (N_16628,N_13753,N_14134);
nor U16629 (N_16629,N_14299,N_13383);
nor U16630 (N_16630,N_14738,N_15283);
xnor U16631 (N_16631,N_12822,N_15421);
xor U16632 (N_16632,N_15391,N_12625);
or U16633 (N_16633,N_14334,N_14908);
and U16634 (N_16634,N_15140,N_15454);
xor U16635 (N_16635,N_15138,N_13664);
and U16636 (N_16636,N_13929,N_13521);
nand U16637 (N_16637,N_14255,N_14896);
or U16638 (N_16638,N_12856,N_15477);
or U16639 (N_16639,N_14469,N_13125);
nand U16640 (N_16640,N_12759,N_15135);
nand U16641 (N_16641,N_14876,N_12933);
or U16642 (N_16642,N_15255,N_13072);
or U16643 (N_16643,N_13966,N_15434);
and U16644 (N_16644,N_13441,N_14790);
nand U16645 (N_16645,N_14637,N_13400);
nor U16646 (N_16646,N_13252,N_14197);
xnor U16647 (N_16647,N_14271,N_15118);
nor U16648 (N_16648,N_15403,N_13232);
and U16649 (N_16649,N_12855,N_14115);
or U16650 (N_16650,N_13076,N_13548);
nor U16651 (N_16651,N_12869,N_13870);
and U16652 (N_16652,N_15593,N_14664);
or U16653 (N_16653,N_12758,N_13442);
nand U16654 (N_16654,N_13409,N_12563);
nor U16655 (N_16655,N_15150,N_14371);
nand U16656 (N_16656,N_14812,N_14753);
nor U16657 (N_16657,N_13281,N_15106);
and U16658 (N_16658,N_13152,N_14114);
and U16659 (N_16659,N_12597,N_12824);
xnor U16660 (N_16660,N_13484,N_14978);
nor U16661 (N_16661,N_15550,N_13502);
nor U16662 (N_16662,N_14887,N_14984);
and U16663 (N_16663,N_12777,N_13322);
and U16664 (N_16664,N_14461,N_14099);
xor U16665 (N_16665,N_14699,N_14948);
or U16666 (N_16666,N_14734,N_13475);
nor U16667 (N_16667,N_15132,N_13894);
and U16668 (N_16668,N_12769,N_13328);
xor U16669 (N_16669,N_12867,N_12564);
and U16670 (N_16670,N_13941,N_13196);
nand U16671 (N_16671,N_14190,N_15009);
nand U16672 (N_16672,N_12692,N_14186);
xor U16673 (N_16673,N_12980,N_12624);
nand U16674 (N_16674,N_12517,N_14160);
xor U16675 (N_16675,N_13367,N_13113);
or U16676 (N_16676,N_13678,N_14707);
nor U16677 (N_16677,N_14680,N_13945);
and U16678 (N_16678,N_14740,N_13012);
and U16679 (N_16679,N_12664,N_12956);
nand U16680 (N_16680,N_13170,N_13157);
nor U16681 (N_16681,N_13725,N_13054);
and U16682 (N_16682,N_14792,N_13317);
nor U16683 (N_16683,N_14613,N_13078);
nand U16684 (N_16684,N_14054,N_15202);
xnor U16685 (N_16685,N_13488,N_14422);
xor U16686 (N_16686,N_14898,N_15465);
or U16687 (N_16687,N_14063,N_13351);
and U16688 (N_16688,N_15475,N_14090);
xor U16689 (N_16689,N_14520,N_13780);
or U16690 (N_16690,N_14235,N_13332);
nand U16691 (N_16691,N_13194,N_12683);
nor U16692 (N_16692,N_14599,N_13364);
nand U16693 (N_16693,N_14167,N_13023);
xor U16694 (N_16694,N_15610,N_13541);
xor U16695 (N_16695,N_15045,N_15491);
or U16696 (N_16696,N_14498,N_12608);
or U16697 (N_16697,N_15333,N_13412);
xnor U16698 (N_16698,N_13840,N_14550);
nand U16699 (N_16699,N_13646,N_15330);
nor U16700 (N_16700,N_15204,N_15281);
and U16701 (N_16701,N_13745,N_14010);
and U16702 (N_16702,N_14518,N_14974);
nand U16703 (N_16703,N_12960,N_14541);
or U16704 (N_16704,N_13297,N_13261);
xor U16705 (N_16705,N_14515,N_13529);
or U16706 (N_16706,N_15170,N_13276);
nor U16707 (N_16707,N_13545,N_15114);
nand U16708 (N_16708,N_15487,N_14813);
nand U16709 (N_16709,N_13849,N_12699);
or U16710 (N_16710,N_13684,N_14493);
xnor U16711 (N_16711,N_14398,N_13640);
nand U16712 (N_16712,N_14605,N_13855);
and U16713 (N_16713,N_14449,N_13749);
and U16714 (N_16714,N_13831,N_15322);
nand U16715 (N_16715,N_14046,N_14497);
xnor U16716 (N_16716,N_14923,N_12971);
or U16717 (N_16717,N_13844,N_15053);
and U16718 (N_16718,N_12924,N_12547);
and U16719 (N_16719,N_13612,N_12736);
and U16720 (N_16720,N_13126,N_13777);
nor U16721 (N_16721,N_14017,N_15369);
nand U16722 (N_16722,N_15613,N_13061);
and U16723 (N_16723,N_12708,N_14532);
xnor U16724 (N_16724,N_12864,N_14732);
nor U16725 (N_16725,N_14045,N_15508);
nor U16726 (N_16726,N_12522,N_14553);
nor U16727 (N_16727,N_12886,N_13073);
xnor U16728 (N_16728,N_14384,N_14240);
and U16729 (N_16729,N_13447,N_13154);
nor U16730 (N_16730,N_13401,N_15119);
nand U16731 (N_16731,N_15340,N_13683);
or U16732 (N_16732,N_15247,N_12765);
nand U16733 (N_16733,N_12537,N_14395);
xnor U16734 (N_16734,N_15537,N_14392);
nand U16735 (N_16735,N_15002,N_13372);
nand U16736 (N_16736,N_13668,N_12748);
nor U16737 (N_16737,N_12796,N_14565);
nand U16738 (N_16738,N_14997,N_15468);
or U16739 (N_16739,N_15438,N_14622);
nor U16740 (N_16740,N_14116,N_13504);
and U16741 (N_16741,N_15187,N_12928);
nand U16742 (N_16742,N_12599,N_13624);
or U16743 (N_16743,N_13490,N_15415);
nor U16744 (N_16744,N_14961,N_12548);
nor U16745 (N_16745,N_14459,N_15614);
nor U16746 (N_16746,N_14845,N_12566);
and U16747 (N_16747,N_15145,N_14686);
xnor U16748 (N_16748,N_14246,N_13949);
nor U16749 (N_16749,N_13174,N_13440);
nand U16750 (N_16750,N_14089,N_14161);
nor U16751 (N_16751,N_13135,N_14436);
or U16752 (N_16752,N_13292,N_13290);
xor U16753 (N_16753,N_13191,N_13350);
xor U16754 (N_16754,N_13344,N_14837);
nand U16755 (N_16755,N_15156,N_13526);
and U16756 (N_16756,N_12862,N_13620);
and U16757 (N_16757,N_14648,N_13615);
nand U16758 (N_16758,N_13160,N_15569);
and U16759 (N_16759,N_15328,N_14405);
nor U16760 (N_16760,N_14123,N_15312);
xor U16761 (N_16761,N_14632,N_13208);
nor U16762 (N_16762,N_12717,N_13743);
or U16763 (N_16763,N_13166,N_15275);
or U16764 (N_16764,N_13709,N_12840);
nand U16765 (N_16765,N_13251,N_15422);
nand U16766 (N_16766,N_15444,N_12893);
nand U16767 (N_16767,N_13799,N_13010);
nand U16768 (N_16768,N_14926,N_14652);
xor U16769 (N_16769,N_13555,N_14086);
or U16770 (N_16770,N_15611,N_13609);
nand U16771 (N_16771,N_14549,N_13630);
nor U16772 (N_16772,N_15270,N_14551);
and U16773 (N_16773,N_14293,N_12842);
or U16774 (N_16774,N_14181,N_14748);
nor U16775 (N_16775,N_15360,N_15464);
and U16776 (N_16776,N_15366,N_14996);
and U16777 (N_16777,N_12588,N_13760);
nand U16778 (N_16778,N_12716,N_13165);
and U16779 (N_16779,N_15284,N_13486);
or U16780 (N_16780,N_13416,N_12950);
and U16781 (N_16781,N_13594,N_13376);
or U16782 (N_16782,N_15225,N_14418);
nor U16783 (N_16783,N_15081,N_14935);
xor U16784 (N_16784,N_12850,N_14266);
or U16785 (N_16785,N_15526,N_15033);
nand U16786 (N_16786,N_14177,N_15303);
xnor U16787 (N_16787,N_15089,N_13551);
or U16788 (N_16788,N_12942,N_15432);
xor U16789 (N_16789,N_14303,N_14098);
xnor U16790 (N_16790,N_14363,N_12725);
or U16791 (N_16791,N_14020,N_15068);
nor U16792 (N_16792,N_13769,N_14006);
xnor U16793 (N_16793,N_14946,N_13374);
and U16794 (N_16794,N_15343,N_13606);
nor U16795 (N_16795,N_13805,N_14499);
nand U16796 (N_16796,N_12936,N_14534);
nor U16797 (N_16797,N_12539,N_14509);
nor U16798 (N_16798,N_14705,N_14067);
nor U16799 (N_16799,N_12785,N_14877);
xor U16800 (N_16800,N_13069,N_14663);
or U16801 (N_16801,N_15559,N_14794);
and U16802 (N_16802,N_13711,N_13902);
xnor U16803 (N_16803,N_13280,N_15307);
xnor U16804 (N_16804,N_13616,N_13795);
nand U16805 (N_16805,N_12561,N_14913);
xnor U16806 (N_16806,N_13980,N_15509);
nor U16807 (N_16807,N_13458,N_14627);
and U16808 (N_16808,N_14539,N_13053);
and U16809 (N_16809,N_15382,N_15601);
or U16810 (N_16810,N_15419,N_14170);
and U16811 (N_16811,N_14111,N_12633);
or U16812 (N_16812,N_13730,N_12811);
and U16813 (N_16813,N_15179,N_12642);
nand U16814 (N_16814,N_14068,N_13817);
nor U16815 (N_16815,N_12593,N_14425);
nand U16816 (N_16816,N_15109,N_13940);
and U16817 (N_16817,N_14764,N_15353);
nor U16818 (N_16818,N_14065,N_13857);
nand U16819 (N_16819,N_13898,N_12911);
and U16820 (N_16820,N_12592,N_15189);
xnor U16821 (N_16821,N_13153,N_12879);
nor U16822 (N_16822,N_13040,N_13103);
or U16823 (N_16823,N_13226,N_14274);
or U16824 (N_16824,N_12604,N_14077);
or U16825 (N_16825,N_15510,N_14786);
nor U16826 (N_16826,N_12518,N_14947);
and U16827 (N_16827,N_13845,N_13742);
nor U16828 (N_16828,N_13454,N_14028);
xor U16829 (N_16829,N_13712,N_14955);
nor U16830 (N_16830,N_13731,N_15612);
or U16831 (N_16831,N_13932,N_13663);
or U16832 (N_16832,N_15006,N_15594);
or U16833 (N_16833,N_15126,N_13794);
xnor U16834 (N_16834,N_12847,N_14725);
and U16835 (N_16835,N_15337,N_12634);
or U16836 (N_16836,N_15558,N_13603);
nand U16837 (N_16837,N_14506,N_13491);
nor U16838 (N_16838,N_13997,N_14954);
or U16839 (N_16839,N_14938,N_14693);
xor U16840 (N_16840,N_14513,N_14581);
xnor U16841 (N_16841,N_12682,N_12562);
or U16842 (N_16842,N_15200,N_15549);
nand U16843 (N_16843,N_12532,N_15527);
xnor U16844 (N_16844,N_15288,N_14383);
and U16845 (N_16845,N_13031,N_14943);
nand U16846 (N_16846,N_13626,N_14176);
nor U16847 (N_16847,N_14346,N_15168);
nor U16848 (N_16848,N_14373,N_12606);
xnor U16849 (N_16849,N_13379,N_14890);
and U16850 (N_16850,N_12755,N_12581);
nor U16851 (N_16851,N_12732,N_14563);
xnor U16852 (N_16852,N_14879,N_13089);
and U16853 (N_16853,N_15462,N_13008);
nor U16854 (N_16854,N_15186,N_14074);
or U16855 (N_16855,N_12902,N_13375);
nor U16856 (N_16856,N_14505,N_13294);
and U16857 (N_16857,N_14507,N_13244);
and U16858 (N_16858,N_15169,N_14962);
and U16859 (N_16859,N_13562,N_15028);
nand U16860 (N_16860,N_14052,N_12574);
xnor U16861 (N_16861,N_13455,N_12646);
nor U16862 (N_16862,N_12655,N_14318);
nand U16863 (N_16863,N_12680,N_12656);
nor U16864 (N_16864,N_13944,N_14402);
and U16865 (N_16865,N_13057,N_14918);
or U16866 (N_16866,N_15437,N_13861);
or U16867 (N_16867,N_12743,N_12932);
and U16868 (N_16868,N_15585,N_15074);
or U16869 (N_16869,N_13621,N_14319);
or U16870 (N_16870,N_14191,N_15185);
or U16871 (N_16871,N_15260,N_13445);
nor U16872 (N_16872,N_13298,N_15480);
and U16873 (N_16873,N_14671,N_13858);
xor U16874 (N_16874,N_14117,N_12720);
nor U16875 (N_16875,N_12835,N_13204);
and U16876 (N_16876,N_13706,N_14298);
xnor U16877 (N_16877,N_14316,N_12848);
nor U16878 (N_16878,N_13398,N_13042);
nand U16879 (N_16879,N_15261,N_14413);
and U16880 (N_16880,N_13695,N_14145);
nand U16881 (N_16881,N_14585,N_14577);
xnor U16882 (N_16882,N_14822,N_13341);
nor U16883 (N_16883,N_14942,N_12711);
and U16884 (N_16884,N_15142,N_14784);
xnor U16885 (N_16885,N_13224,N_13610);
nor U16886 (N_16886,N_15471,N_14312);
xnor U16887 (N_16887,N_13030,N_15393);
nand U16888 (N_16888,N_14236,N_13694);
xnor U16889 (N_16889,N_13705,N_13644);
or U16890 (N_16890,N_14066,N_13524);
nor U16891 (N_16891,N_14171,N_14659);
xnor U16892 (N_16892,N_13629,N_13411);
nor U16893 (N_16893,N_13359,N_14629);
nor U16894 (N_16894,N_15319,N_13483);
xor U16895 (N_16895,N_13759,N_12887);
nand U16896 (N_16896,N_14433,N_13286);
and U16897 (N_16897,N_13901,N_12734);
nor U16898 (N_16898,N_14482,N_13468);
nor U16899 (N_16899,N_12966,N_14397);
or U16900 (N_16900,N_15356,N_13200);
and U16901 (N_16901,N_15311,N_13974);
and U16902 (N_16902,N_15277,N_12970);
and U16903 (N_16903,N_14194,N_14016);
nor U16904 (N_16904,N_15414,N_12565);
nand U16905 (N_16905,N_12544,N_13979);
or U16906 (N_16906,N_15067,N_13810);
and U16907 (N_16907,N_13133,N_15467);
xnor U16908 (N_16908,N_13569,N_13674);
xor U16909 (N_16909,N_13791,N_13889);
nand U16910 (N_16910,N_15215,N_15234);
nand U16911 (N_16911,N_14836,N_13258);
nor U16912 (N_16912,N_13489,N_15482);
or U16913 (N_16913,N_12662,N_14426);
xnor U16914 (N_16914,N_13326,N_14989);
and U16915 (N_16915,N_14778,N_13654);
nand U16916 (N_16916,N_14751,N_13327);
xor U16917 (N_16917,N_15492,N_13538);
xor U16918 (N_16918,N_13247,N_13032);
and U16919 (N_16919,N_13574,N_12961);
nand U16920 (N_16920,N_14841,N_15292);
nand U16921 (N_16921,N_15071,N_13217);
xor U16922 (N_16922,N_13405,N_14793);
or U16923 (N_16923,N_14568,N_14594);
and U16924 (N_16924,N_12776,N_13639);
nor U16925 (N_16925,N_13071,N_13701);
nand U16926 (N_16926,N_12945,N_14524);
and U16927 (N_16927,N_13515,N_13391);
nand U16928 (N_16928,N_15093,N_15280);
or U16929 (N_16929,N_15445,N_12507);
xor U16930 (N_16930,N_14902,N_15529);
or U16931 (N_16931,N_12836,N_15123);
and U16932 (N_16932,N_13587,N_12579);
xor U16933 (N_16933,N_15210,N_14168);
and U16934 (N_16934,N_13150,N_14579);
nor U16935 (N_16935,N_14774,N_14263);
nor U16936 (N_16936,N_14769,N_13380);
or U16937 (N_16937,N_14403,N_13129);
nand U16938 (N_16938,N_13002,N_13393);
or U16939 (N_16939,N_13946,N_14372);
xor U16940 (N_16940,N_15470,N_12858);
xnor U16941 (N_16941,N_13346,N_15104);
xnor U16942 (N_16942,N_15545,N_12553);
nor U16943 (N_16943,N_15226,N_15587);
nor U16944 (N_16944,N_12536,N_15562);
xor U16945 (N_16945,N_13740,N_12582);
and U16946 (N_16946,N_13918,N_13255);
nand U16947 (N_16947,N_15144,N_12703);
xor U16948 (N_16948,N_14669,N_14362);
and U16949 (N_16949,N_15058,N_14696);
or U16950 (N_16950,N_12790,N_13860);
and U16951 (N_16951,N_14848,N_14735);
nand U16952 (N_16952,N_12596,N_12834);
xnor U16953 (N_16953,N_13110,N_13303);
or U16954 (N_16954,N_14022,N_14087);
xnor U16955 (N_16955,N_13331,N_14015);
and U16956 (N_16956,N_14817,N_14296);
and U16957 (N_16957,N_15522,N_14278);
xnor U16958 (N_16958,N_14536,N_12559);
and U16959 (N_16959,N_13108,N_12987);
nor U16960 (N_16960,N_14816,N_14193);
or U16961 (N_16961,N_13279,N_12616);
nand U16962 (N_16962,N_13596,N_14607);
or U16963 (N_16963,N_14101,N_12997);
or U16964 (N_16964,N_13075,N_13177);
or U16965 (N_16965,N_14382,N_13707);
nor U16966 (N_16966,N_14354,N_12916);
or U16967 (N_16967,N_13677,N_12962);
xor U16968 (N_16968,N_13934,N_13199);
nand U16969 (N_16969,N_14387,N_14410);
or U16970 (N_16970,N_13847,N_14400);
nand U16971 (N_16971,N_12937,N_13938);
or U16972 (N_16972,N_12979,N_14626);
nor U16973 (N_16973,N_15164,N_13451);
and U16974 (N_16974,N_13171,N_13168);
xor U16975 (N_16975,N_14011,N_13904);
xnor U16976 (N_16976,N_14660,N_12639);
nor U16977 (N_16977,N_14544,N_15239);
and U16978 (N_16978,N_15335,N_14647);
nor U16979 (N_16979,N_14801,N_13948);
and U16980 (N_16980,N_13369,N_13653);
xnor U16981 (N_16981,N_13143,N_13696);
nor U16982 (N_16982,N_12668,N_15130);
nor U16983 (N_16983,N_15608,N_15177);
or U16984 (N_16984,N_13703,N_12640);
nand U16985 (N_16985,N_15457,N_14072);
xor U16986 (N_16986,N_15459,N_14322);
nand U16987 (N_16987,N_15237,N_14286);
xor U16988 (N_16988,N_15486,N_13470);
xnor U16989 (N_16989,N_15401,N_14040);
and U16990 (N_16990,N_14609,N_12648);
or U16991 (N_16991,N_14584,N_13536);
or U16992 (N_16992,N_13874,N_13790);
xnor U16993 (N_16993,N_13039,N_13132);
and U16994 (N_16994,N_13473,N_14589);
and U16995 (N_16995,N_12760,N_13809);
xnor U16996 (N_16996,N_12803,N_15615);
and U16997 (N_16997,N_15041,N_14977);
and U16998 (N_16998,N_13128,N_15318);
or U16999 (N_16999,N_14856,N_13919);
xor U17000 (N_17000,N_12949,N_14222);
xnor U17001 (N_17001,N_13138,N_12741);
and U17002 (N_17002,N_13785,N_13172);
nor U17003 (N_17003,N_13260,N_12783);
and U17004 (N_17004,N_13452,N_14993);
or U17005 (N_17005,N_13567,N_14103);
nand U17006 (N_17006,N_14728,N_13930);
xnor U17007 (N_17007,N_12908,N_15554);
and U17008 (N_17008,N_13517,N_13220);
and U17009 (N_17009,N_13338,N_14800);
nand U17010 (N_17010,N_13843,N_15308);
xor U17011 (N_17011,N_13318,N_12578);
or U17012 (N_17012,N_13167,N_15129);
nor U17013 (N_17013,N_15574,N_15113);
and U17014 (N_17014,N_15305,N_14849);
and U17015 (N_17015,N_14525,N_12876);
or U17016 (N_17016,N_15181,N_13882);
nand U17017 (N_17017,N_14985,N_13720);
nor U17018 (N_17018,N_13037,N_13746);
or U17019 (N_17019,N_15022,N_12771);
xor U17020 (N_17020,N_13000,N_15115);
nand U17021 (N_17021,N_13729,N_14377);
nor U17022 (N_17022,N_13905,N_13418);
xnor U17023 (N_17023,N_13507,N_14213);
or U17024 (N_17024,N_14310,N_14820);
and U17025 (N_17025,N_14526,N_14742);
nor U17026 (N_17026,N_13916,N_14847);
nor U17027 (N_17027,N_13436,N_13187);
and U17028 (N_17028,N_12882,N_14503);
nand U17029 (N_17029,N_13661,N_13357);
and U17030 (N_17030,N_13975,N_14951);
nand U17031 (N_17031,N_13962,N_15377);
or U17032 (N_17032,N_13642,N_15290);
xnor U17033 (N_17033,N_15420,N_12839);
and U17034 (N_17034,N_13826,N_15399);
nand U17035 (N_17035,N_13834,N_13254);
nor U17036 (N_17036,N_12704,N_14811);
and U17037 (N_17037,N_15160,N_14352);
and U17038 (N_17038,N_14280,N_13299);
or U17039 (N_17039,N_12598,N_15588);
nand U17040 (N_17040,N_13238,N_14894);
nor U17041 (N_17041,N_15578,N_13340);
xnor U17042 (N_17042,N_15354,N_12651);
nor U17043 (N_17043,N_12873,N_13291);
xor U17044 (N_17044,N_15347,N_14008);
or U17045 (N_17045,N_13584,N_15383);
nand U17046 (N_17046,N_13460,N_14566);
nand U17047 (N_17047,N_13339,N_12798);
or U17048 (N_17048,N_14490,N_14729);
nand U17049 (N_17049,N_12531,N_13666);
nand U17050 (N_17050,N_14533,N_14870);
nor U17051 (N_17051,N_14582,N_13796);
or U17052 (N_17052,N_13828,N_13892);
and U17053 (N_17053,N_12819,N_13368);
and U17054 (N_17054,N_15542,N_13011);
or U17055 (N_17055,N_15289,N_12923);
xnor U17056 (N_17056,N_15387,N_12712);
nand U17057 (N_17057,N_13823,N_14244);
or U17058 (N_17058,N_14819,N_14633);
and U17059 (N_17059,N_15039,N_14338);
or U17060 (N_17060,N_12829,N_12922);
or U17061 (N_17061,N_13558,N_15365);
xnor U17062 (N_17062,N_15148,N_12615);
xnor U17063 (N_17063,N_13482,N_13924);
nand U17064 (N_17064,N_14694,N_12954);
xnor U17065 (N_17065,N_13800,N_14229);
nor U17066 (N_17066,N_13353,N_15217);
and U17067 (N_17067,N_13613,N_14983);
xnor U17068 (N_17068,N_15409,N_14021);
or U17069 (N_17069,N_12946,N_15279);
and U17070 (N_17070,N_12825,N_13288);
nor U17071 (N_17071,N_14305,N_13395);
or U17072 (N_17072,N_13688,N_13886);
or U17073 (N_17073,N_13256,N_15589);
and U17074 (N_17074,N_13920,N_12910);
nand U17075 (N_17075,N_15205,N_13917);
nand U17076 (N_17076,N_12626,N_12901);
and U17077 (N_17077,N_14670,N_12568);
and U17078 (N_17078,N_13530,N_15037);
or U17079 (N_17079,N_15455,N_14234);
or U17080 (N_17080,N_15350,N_14798);
nand U17081 (N_17081,N_13802,N_14137);
nand U17082 (N_17082,N_14038,N_13827);
or U17083 (N_17083,N_14220,N_14775);
nor U17084 (N_17084,N_14839,N_12881);
and U17085 (N_17085,N_13231,N_12931);
or U17086 (N_17086,N_14657,N_12818);
or U17087 (N_17087,N_15379,N_12684);
and U17088 (N_17088,N_13878,N_13324);
and U17089 (N_17089,N_14884,N_14556);
xnor U17090 (N_17090,N_13841,N_13107);
nor U17091 (N_17091,N_15514,N_13001);
or U17092 (N_17092,N_13070,N_14785);
or U17093 (N_17093,N_15624,N_14990);
and U17094 (N_17094,N_13838,N_13406);
nand U17095 (N_17095,N_12737,N_14393);
or U17096 (N_17096,N_12556,N_14560);
nor U17097 (N_17097,N_14472,N_12645);
xor U17098 (N_17098,N_15174,N_12681);
nor U17099 (N_17099,N_13964,N_12535);
nand U17100 (N_17100,N_13027,N_14419);
nand U17101 (N_17101,N_14825,N_14771);
and U17102 (N_17102,N_14829,N_14635);
nand U17103 (N_17103,N_15287,N_13643);
nand U17104 (N_17104,N_14956,N_13699);
nor U17105 (N_17105,N_14866,N_13361);
and U17106 (N_17106,N_12751,N_14909);
nor U17107 (N_17107,N_12904,N_13685);
xor U17108 (N_17108,N_13996,N_14762);
nor U17109 (N_17109,N_15507,N_14611);
or U17110 (N_17110,N_13067,N_13970);
and U17111 (N_17111,N_15207,N_13947);
nand U17112 (N_17112,N_14818,N_13659);
and U17113 (N_17113,N_14617,N_15336);
nand U17114 (N_17114,N_13926,N_13036);
and U17115 (N_17115,N_13985,N_14716);
and U17116 (N_17116,N_13973,N_14430);
nor U17117 (N_17117,N_14795,N_14888);
xor U17118 (N_17118,N_12523,N_14127);
or U17119 (N_17119,N_12947,N_14147);
or U17120 (N_17120,N_14144,N_13768);
nand U17121 (N_17121,N_14163,N_14226);
or U17122 (N_17122,N_14712,N_13093);
xnor U17123 (N_17123,N_15276,N_12837);
nand U17124 (N_17124,N_13772,N_13148);
and U17125 (N_17125,N_12843,N_14502);
nand U17126 (N_17126,N_12520,N_14448);
or U17127 (N_17127,N_14355,N_14245);
nand U17128 (N_17128,N_12750,N_13273);
nor U17129 (N_17129,N_13034,N_15221);
nor U17130 (N_17130,N_14752,N_14462);
nand U17131 (N_17131,N_15124,N_12900);
or U17132 (N_17132,N_14442,N_13923);
or U17133 (N_17133,N_14636,N_13998);
or U17134 (N_17134,N_12788,N_14834);
xnor U17135 (N_17135,N_15344,N_13112);
or U17136 (N_17136,N_14931,N_14388);
xor U17137 (N_17137,N_12739,N_14932);
or U17138 (N_17138,N_15254,N_14624);
nor U17139 (N_17139,N_13896,N_13755);
xnor U17140 (N_17140,N_13471,N_14307);
and U17141 (N_17141,N_15599,N_12735);
and U17142 (N_17142,N_13080,N_13822);
nor U17143 (N_17143,N_13853,N_13825);
xor U17144 (N_17144,N_15351,N_13306);
and U17145 (N_17145,N_13510,N_12706);
or U17146 (N_17146,N_12889,N_12909);
or U17147 (N_17147,N_15441,N_14124);
nand U17148 (N_17148,N_15532,N_14521);
nor U17149 (N_17149,N_14173,N_13049);
and U17150 (N_17150,N_14885,N_14761);
nand U17151 (N_17151,N_13474,N_14481);
or U17152 (N_17152,N_14148,N_13308);
xnor U17153 (N_17153,N_15040,N_12713);
xor U17154 (N_17154,N_13784,N_13390);
and U17155 (N_17155,N_13178,N_13022);
and U17156 (N_17156,N_13205,N_13681);
and U17157 (N_17157,N_13813,N_15019);
or U17158 (N_17158,N_14049,N_12714);
or U17159 (N_17159,N_14804,N_15125);
nand U17160 (N_17160,N_13617,N_15013);
and U17161 (N_17161,N_14302,N_13463);
and U17162 (N_17162,N_12968,N_14744);
or U17163 (N_17163,N_15272,N_15010);
nor U17164 (N_17164,N_13315,N_13239);
and U17165 (N_17165,N_13018,N_12557);
nand U17166 (N_17166,N_14454,N_12546);
nand U17167 (N_17167,N_12861,N_13984);
and U17168 (N_17168,N_13786,N_13689);
and U17169 (N_17169,N_14721,N_15501);
xor U17170 (N_17170,N_14432,N_14164);
nor U17171 (N_17171,N_15293,N_15062);
nor U17172 (N_17172,N_12525,N_13519);
nor U17173 (N_17173,N_13090,N_15173);
nand U17174 (N_17174,N_15249,N_15103);
or U17175 (N_17175,N_14612,N_14796);
or U17176 (N_17176,N_14092,N_13116);
nor U17177 (N_17177,N_12695,N_15030);
or U17178 (N_17178,N_12533,N_14272);
xor U17179 (N_17179,N_14713,N_13161);
and U17180 (N_17180,N_14491,N_14510);
and U17181 (N_17181,N_12821,N_14342);
or U17182 (N_17182,N_14451,N_13404);
or U17183 (N_17183,N_13192,N_14126);
and U17184 (N_17184,N_12621,N_13443);
nor U17185 (N_17185,N_15474,N_15291);
nor U17186 (N_17186,N_13118,N_14141);
nor U17187 (N_17187,N_14057,N_13211);
or U17188 (N_17188,N_13433,N_13844);
xnor U17189 (N_17189,N_14192,N_15549);
and U17190 (N_17190,N_12875,N_14902);
and U17191 (N_17191,N_13483,N_13667);
or U17192 (N_17192,N_14188,N_13983);
or U17193 (N_17193,N_13444,N_15498);
nand U17194 (N_17194,N_15294,N_14314);
nand U17195 (N_17195,N_12988,N_13434);
nand U17196 (N_17196,N_13968,N_14937);
nor U17197 (N_17197,N_15271,N_13050);
xnor U17198 (N_17198,N_13574,N_15095);
nand U17199 (N_17199,N_15081,N_14584);
or U17200 (N_17200,N_12727,N_12568);
xor U17201 (N_17201,N_13254,N_15337);
nand U17202 (N_17202,N_15490,N_15512);
and U17203 (N_17203,N_14691,N_15216);
or U17204 (N_17204,N_12846,N_15004);
and U17205 (N_17205,N_13734,N_13489);
and U17206 (N_17206,N_15171,N_14504);
nand U17207 (N_17207,N_14420,N_13604);
and U17208 (N_17208,N_13677,N_14184);
nand U17209 (N_17209,N_13214,N_15503);
xor U17210 (N_17210,N_12577,N_15107);
or U17211 (N_17211,N_14323,N_14411);
and U17212 (N_17212,N_13605,N_12523);
and U17213 (N_17213,N_12507,N_14020);
nor U17214 (N_17214,N_13711,N_12913);
and U17215 (N_17215,N_14010,N_13677);
nand U17216 (N_17216,N_13979,N_15423);
nor U17217 (N_17217,N_14870,N_15126);
and U17218 (N_17218,N_15467,N_15590);
nor U17219 (N_17219,N_14916,N_14828);
xor U17220 (N_17220,N_15310,N_15159);
nor U17221 (N_17221,N_12525,N_12721);
and U17222 (N_17222,N_12960,N_15170);
xor U17223 (N_17223,N_15435,N_13502);
nor U17224 (N_17224,N_14895,N_14169);
xnor U17225 (N_17225,N_13390,N_13096);
and U17226 (N_17226,N_12589,N_13376);
xnor U17227 (N_17227,N_14351,N_15113);
nor U17228 (N_17228,N_14318,N_12708);
or U17229 (N_17229,N_12578,N_15331);
or U17230 (N_17230,N_15236,N_14371);
and U17231 (N_17231,N_14765,N_12590);
or U17232 (N_17232,N_13916,N_13696);
or U17233 (N_17233,N_12664,N_12820);
nand U17234 (N_17234,N_12916,N_15609);
and U17235 (N_17235,N_14197,N_13958);
xor U17236 (N_17236,N_14033,N_15271);
xnor U17237 (N_17237,N_14776,N_14990);
nor U17238 (N_17238,N_14584,N_13449);
and U17239 (N_17239,N_13403,N_14506);
and U17240 (N_17240,N_14775,N_13275);
and U17241 (N_17241,N_13893,N_15189);
nor U17242 (N_17242,N_15002,N_14112);
nor U17243 (N_17243,N_14281,N_14706);
or U17244 (N_17244,N_12954,N_14882);
nor U17245 (N_17245,N_13792,N_13723);
nand U17246 (N_17246,N_15283,N_15007);
nor U17247 (N_17247,N_13205,N_15255);
nor U17248 (N_17248,N_13239,N_12981);
and U17249 (N_17249,N_15030,N_15421);
nand U17250 (N_17250,N_15372,N_13782);
nand U17251 (N_17251,N_13607,N_15584);
or U17252 (N_17252,N_15359,N_14627);
and U17253 (N_17253,N_12653,N_14259);
nand U17254 (N_17254,N_14177,N_13845);
nor U17255 (N_17255,N_13853,N_14897);
and U17256 (N_17256,N_14368,N_15412);
or U17257 (N_17257,N_12630,N_12963);
nand U17258 (N_17258,N_15308,N_14516);
nand U17259 (N_17259,N_14445,N_12764);
nor U17260 (N_17260,N_13674,N_14385);
or U17261 (N_17261,N_14625,N_15517);
xor U17262 (N_17262,N_13127,N_14813);
nor U17263 (N_17263,N_13789,N_13886);
xor U17264 (N_17264,N_14471,N_15064);
nor U17265 (N_17265,N_12504,N_13963);
xor U17266 (N_17266,N_12923,N_12953);
nand U17267 (N_17267,N_12699,N_13283);
xor U17268 (N_17268,N_13994,N_13169);
and U17269 (N_17269,N_13841,N_13649);
and U17270 (N_17270,N_12897,N_14870);
nor U17271 (N_17271,N_13229,N_14272);
or U17272 (N_17272,N_13612,N_12699);
nand U17273 (N_17273,N_14380,N_13489);
and U17274 (N_17274,N_13543,N_13740);
or U17275 (N_17275,N_13507,N_14424);
xnor U17276 (N_17276,N_15137,N_15554);
xnor U17277 (N_17277,N_13713,N_13920);
xor U17278 (N_17278,N_14842,N_13684);
nand U17279 (N_17279,N_15304,N_12628);
nand U17280 (N_17280,N_12565,N_14179);
xnor U17281 (N_17281,N_13017,N_13075);
nor U17282 (N_17282,N_15072,N_15584);
and U17283 (N_17283,N_12683,N_14843);
or U17284 (N_17284,N_15464,N_15090);
and U17285 (N_17285,N_13232,N_15245);
nor U17286 (N_17286,N_15081,N_13898);
or U17287 (N_17287,N_13470,N_13953);
or U17288 (N_17288,N_14629,N_13163);
or U17289 (N_17289,N_15379,N_15333);
nand U17290 (N_17290,N_12892,N_13308);
nand U17291 (N_17291,N_13342,N_14320);
nor U17292 (N_17292,N_12872,N_13756);
and U17293 (N_17293,N_13664,N_12520);
or U17294 (N_17294,N_14509,N_12983);
and U17295 (N_17295,N_15182,N_13830);
nor U17296 (N_17296,N_15119,N_13041);
xnor U17297 (N_17297,N_14815,N_13953);
and U17298 (N_17298,N_13955,N_12630);
and U17299 (N_17299,N_13902,N_13027);
nand U17300 (N_17300,N_13735,N_13172);
and U17301 (N_17301,N_13514,N_14035);
nor U17302 (N_17302,N_13610,N_14213);
xor U17303 (N_17303,N_13861,N_14327);
nor U17304 (N_17304,N_12782,N_14038);
nor U17305 (N_17305,N_14534,N_14828);
nand U17306 (N_17306,N_13770,N_12591);
or U17307 (N_17307,N_14235,N_13776);
and U17308 (N_17308,N_14211,N_14183);
or U17309 (N_17309,N_14737,N_12947);
nor U17310 (N_17310,N_12754,N_12683);
and U17311 (N_17311,N_13716,N_13598);
nor U17312 (N_17312,N_13655,N_13243);
and U17313 (N_17313,N_15260,N_14581);
xnor U17314 (N_17314,N_14983,N_13401);
nor U17315 (N_17315,N_13190,N_13479);
nor U17316 (N_17316,N_12572,N_13268);
or U17317 (N_17317,N_14995,N_13018);
nor U17318 (N_17318,N_14576,N_13476);
nand U17319 (N_17319,N_13159,N_13390);
nor U17320 (N_17320,N_15456,N_13930);
or U17321 (N_17321,N_13289,N_13195);
or U17322 (N_17322,N_14559,N_14430);
or U17323 (N_17323,N_12513,N_15249);
or U17324 (N_17324,N_13719,N_13495);
xor U17325 (N_17325,N_15411,N_15428);
and U17326 (N_17326,N_13825,N_14707);
nand U17327 (N_17327,N_14786,N_15048);
xnor U17328 (N_17328,N_14097,N_14863);
or U17329 (N_17329,N_13753,N_15606);
and U17330 (N_17330,N_13385,N_14005);
or U17331 (N_17331,N_14461,N_12851);
xnor U17332 (N_17332,N_15355,N_12668);
xor U17333 (N_17333,N_15457,N_14596);
nand U17334 (N_17334,N_14637,N_15473);
nor U17335 (N_17335,N_13606,N_14695);
nor U17336 (N_17336,N_12734,N_14002);
nand U17337 (N_17337,N_12848,N_13457);
nand U17338 (N_17338,N_15614,N_14868);
or U17339 (N_17339,N_13646,N_13225);
nor U17340 (N_17340,N_12994,N_12892);
nand U17341 (N_17341,N_15571,N_15557);
nor U17342 (N_17342,N_14254,N_13585);
or U17343 (N_17343,N_15059,N_15295);
nor U17344 (N_17344,N_13367,N_13518);
nor U17345 (N_17345,N_13243,N_15096);
nor U17346 (N_17346,N_15198,N_14962);
nand U17347 (N_17347,N_13672,N_14012);
and U17348 (N_17348,N_14515,N_14878);
nor U17349 (N_17349,N_14159,N_13033);
nand U17350 (N_17350,N_13509,N_13122);
nand U17351 (N_17351,N_14890,N_13894);
and U17352 (N_17352,N_13923,N_13443);
or U17353 (N_17353,N_15222,N_12566);
nor U17354 (N_17354,N_12914,N_14010);
or U17355 (N_17355,N_13078,N_13045);
and U17356 (N_17356,N_14670,N_13966);
and U17357 (N_17357,N_15055,N_15027);
or U17358 (N_17358,N_14399,N_14703);
or U17359 (N_17359,N_15302,N_12667);
xor U17360 (N_17360,N_14333,N_12954);
nand U17361 (N_17361,N_12600,N_12893);
xor U17362 (N_17362,N_14618,N_15390);
nand U17363 (N_17363,N_15319,N_14929);
xor U17364 (N_17364,N_13802,N_14698);
nand U17365 (N_17365,N_15596,N_13428);
nand U17366 (N_17366,N_14184,N_13994);
nor U17367 (N_17367,N_13259,N_12988);
and U17368 (N_17368,N_14655,N_14354);
nor U17369 (N_17369,N_14272,N_14723);
nor U17370 (N_17370,N_13753,N_14042);
nor U17371 (N_17371,N_14841,N_13317);
nand U17372 (N_17372,N_13260,N_14580);
xnor U17373 (N_17373,N_15520,N_12845);
or U17374 (N_17374,N_13614,N_14690);
or U17375 (N_17375,N_12804,N_13146);
nand U17376 (N_17376,N_14859,N_13369);
nor U17377 (N_17377,N_14005,N_13413);
xor U17378 (N_17378,N_13256,N_12881);
nor U17379 (N_17379,N_15085,N_12517);
and U17380 (N_17380,N_14588,N_14030);
or U17381 (N_17381,N_13233,N_12860);
or U17382 (N_17382,N_13018,N_12504);
or U17383 (N_17383,N_12541,N_14772);
nor U17384 (N_17384,N_14691,N_14492);
and U17385 (N_17385,N_13878,N_15025);
nand U17386 (N_17386,N_12718,N_14732);
or U17387 (N_17387,N_13251,N_14900);
nor U17388 (N_17388,N_14775,N_13133);
and U17389 (N_17389,N_15062,N_15250);
nand U17390 (N_17390,N_14966,N_13871);
or U17391 (N_17391,N_14506,N_14886);
xnor U17392 (N_17392,N_15606,N_15435);
and U17393 (N_17393,N_12772,N_15522);
nor U17394 (N_17394,N_12514,N_14808);
xor U17395 (N_17395,N_12618,N_13202);
xor U17396 (N_17396,N_13752,N_13038);
or U17397 (N_17397,N_13754,N_13149);
xor U17398 (N_17398,N_12899,N_15022);
and U17399 (N_17399,N_14362,N_14205);
or U17400 (N_17400,N_13814,N_13519);
or U17401 (N_17401,N_15328,N_15135);
and U17402 (N_17402,N_14018,N_13288);
or U17403 (N_17403,N_14486,N_15460);
xor U17404 (N_17404,N_15085,N_13061);
nor U17405 (N_17405,N_14679,N_14983);
xor U17406 (N_17406,N_13565,N_14674);
nand U17407 (N_17407,N_14832,N_14369);
nor U17408 (N_17408,N_13323,N_15317);
or U17409 (N_17409,N_13869,N_13301);
nor U17410 (N_17410,N_14938,N_12858);
nand U17411 (N_17411,N_14731,N_14739);
nand U17412 (N_17412,N_14748,N_14914);
or U17413 (N_17413,N_15034,N_15032);
xor U17414 (N_17414,N_14837,N_13094);
or U17415 (N_17415,N_14474,N_14472);
or U17416 (N_17416,N_15171,N_14566);
and U17417 (N_17417,N_12942,N_12806);
and U17418 (N_17418,N_13959,N_13838);
xor U17419 (N_17419,N_15182,N_15178);
or U17420 (N_17420,N_12991,N_12670);
nor U17421 (N_17421,N_13926,N_15335);
and U17422 (N_17422,N_12749,N_12674);
xor U17423 (N_17423,N_13659,N_12825);
nand U17424 (N_17424,N_15495,N_12954);
xor U17425 (N_17425,N_15216,N_14502);
and U17426 (N_17426,N_15352,N_14552);
nor U17427 (N_17427,N_14409,N_12584);
xnor U17428 (N_17428,N_13874,N_13311);
nand U17429 (N_17429,N_13252,N_15538);
nor U17430 (N_17430,N_12670,N_15600);
nor U17431 (N_17431,N_13055,N_14494);
nor U17432 (N_17432,N_14492,N_14426);
nand U17433 (N_17433,N_12840,N_14945);
xnor U17434 (N_17434,N_12615,N_12672);
nor U17435 (N_17435,N_14017,N_14398);
and U17436 (N_17436,N_12840,N_14267);
nor U17437 (N_17437,N_14119,N_13772);
nor U17438 (N_17438,N_14928,N_15068);
and U17439 (N_17439,N_15015,N_13738);
and U17440 (N_17440,N_14154,N_13439);
nor U17441 (N_17441,N_13984,N_13531);
or U17442 (N_17442,N_13622,N_12523);
or U17443 (N_17443,N_14363,N_13766);
xor U17444 (N_17444,N_13838,N_14760);
xnor U17445 (N_17445,N_14811,N_13493);
xor U17446 (N_17446,N_14669,N_13399);
nand U17447 (N_17447,N_13574,N_13388);
or U17448 (N_17448,N_12763,N_14025);
nor U17449 (N_17449,N_15276,N_14753);
or U17450 (N_17450,N_14647,N_15250);
and U17451 (N_17451,N_13709,N_14437);
xor U17452 (N_17452,N_15229,N_13896);
nand U17453 (N_17453,N_12946,N_12868);
nor U17454 (N_17454,N_15345,N_13370);
nor U17455 (N_17455,N_13033,N_13612);
or U17456 (N_17456,N_12647,N_12878);
xor U17457 (N_17457,N_14360,N_15176);
nand U17458 (N_17458,N_12509,N_12526);
or U17459 (N_17459,N_15069,N_13044);
nand U17460 (N_17460,N_15143,N_13431);
xnor U17461 (N_17461,N_14896,N_15030);
or U17462 (N_17462,N_15305,N_14428);
and U17463 (N_17463,N_14920,N_13913);
xnor U17464 (N_17464,N_13030,N_15286);
nand U17465 (N_17465,N_15605,N_15512);
and U17466 (N_17466,N_15536,N_15559);
nor U17467 (N_17467,N_15084,N_12516);
nand U17468 (N_17468,N_14903,N_13625);
and U17469 (N_17469,N_13058,N_15598);
or U17470 (N_17470,N_15405,N_14886);
nor U17471 (N_17471,N_14236,N_15443);
nor U17472 (N_17472,N_12596,N_14514);
or U17473 (N_17473,N_13200,N_14587);
xor U17474 (N_17474,N_12674,N_13576);
xnor U17475 (N_17475,N_13428,N_12677);
and U17476 (N_17476,N_14945,N_14735);
xor U17477 (N_17477,N_15396,N_12738);
nor U17478 (N_17478,N_13783,N_15098);
nor U17479 (N_17479,N_14171,N_13436);
or U17480 (N_17480,N_13486,N_14707);
xor U17481 (N_17481,N_14817,N_13490);
nor U17482 (N_17482,N_15354,N_13134);
or U17483 (N_17483,N_13314,N_13536);
nand U17484 (N_17484,N_14331,N_13956);
xor U17485 (N_17485,N_15093,N_14707);
xnor U17486 (N_17486,N_13099,N_14378);
nand U17487 (N_17487,N_14286,N_15589);
nand U17488 (N_17488,N_14721,N_15119);
xnor U17489 (N_17489,N_13269,N_12970);
nor U17490 (N_17490,N_14628,N_15597);
nor U17491 (N_17491,N_14800,N_13244);
and U17492 (N_17492,N_13665,N_14448);
or U17493 (N_17493,N_13335,N_15084);
nor U17494 (N_17494,N_15077,N_15024);
and U17495 (N_17495,N_14607,N_13211);
and U17496 (N_17496,N_14674,N_14768);
xnor U17497 (N_17497,N_14261,N_13039);
xnor U17498 (N_17498,N_14880,N_13928);
xor U17499 (N_17499,N_13210,N_12817);
and U17500 (N_17500,N_14949,N_13802);
nor U17501 (N_17501,N_13435,N_14875);
nand U17502 (N_17502,N_12729,N_15220);
and U17503 (N_17503,N_15574,N_14210);
xor U17504 (N_17504,N_15254,N_15366);
xnor U17505 (N_17505,N_12584,N_14778);
nand U17506 (N_17506,N_15171,N_14808);
nor U17507 (N_17507,N_15141,N_14044);
or U17508 (N_17508,N_15030,N_13562);
xor U17509 (N_17509,N_12557,N_13308);
and U17510 (N_17510,N_14882,N_13610);
nand U17511 (N_17511,N_15326,N_15424);
nand U17512 (N_17512,N_14499,N_15140);
nor U17513 (N_17513,N_13154,N_14816);
xnor U17514 (N_17514,N_12984,N_14030);
nand U17515 (N_17515,N_14028,N_13748);
or U17516 (N_17516,N_14342,N_14145);
and U17517 (N_17517,N_13050,N_13766);
xor U17518 (N_17518,N_14165,N_14001);
xnor U17519 (N_17519,N_13119,N_15034);
or U17520 (N_17520,N_14655,N_14134);
xnor U17521 (N_17521,N_15557,N_13774);
or U17522 (N_17522,N_13899,N_12940);
or U17523 (N_17523,N_13568,N_12991);
nor U17524 (N_17524,N_13034,N_14925);
nand U17525 (N_17525,N_13841,N_13898);
nor U17526 (N_17526,N_12833,N_14926);
or U17527 (N_17527,N_14325,N_13306);
and U17528 (N_17528,N_13249,N_14938);
nand U17529 (N_17529,N_14828,N_13049);
nand U17530 (N_17530,N_12658,N_13273);
or U17531 (N_17531,N_13395,N_13195);
and U17532 (N_17532,N_12661,N_13029);
or U17533 (N_17533,N_15617,N_13117);
and U17534 (N_17534,N_15012,N_13801);
nor U17535 (N_17535,N_12727,N_14724);
xnor U17536 (N_17536,N_13002,N_13536);
nor U17537 (N_17537,N_13860,N_13578);
and U17538 (N_17538,N_13842,N_13563);
nand U17539 (N_17539,N_14849,N_13031);
xnor U17540 (N_17540,N_14622,N_15236);
xnor U17541 (N_17541,N_12781,N_14062);
nor U17542 (N_17542,N_12881,N_14158);
or U17543 (N_17543,N_13273,N_15290);
nor U17544 (N_17544,N_14824,N_12982);
nor U17545 (N_17545,N_12664,N_14225);
nand U17546 (N_17546,N_12685,N_13757);
and U17547 (N_17547,N_14699,N_14998);
xor U17548 (N_17548,N_14567,N_15130);
nor U17549 (N_17549,N_13145,N_13406);
xnor U17550 (N_17550,N_13979,N_13512);
xor U17551 (N_17551,N_14709,N_14007);
xnor U17552 (N_17552,N_14238,N_14068);
nand U17553 (N_17553,N_13497,N_14248);
or U17554 (N_17554,N_14239,N_13643);
or U17555 (N_17555,N_14446,N_13693);
nand U17556 (N_17556,N_12589,N_14023);
nand U17557 (N_17557,N_15066,N_15057);
and U17558 (N_17558,N_14677,N_13419);
or U17559 (N_17559,N_15558,N_15588);
nand U17560 (N_17560,N_13473,N_15104);
nand U17561 (N_17561,N_14974,N_12683);
nor U17562 (N_17562,N_14807,N_15393);
nand U17563 (N_17563,N_14938,N_13843);
nor U17564 (N_17564,N_12883,N_15079);
nor U17565 (N_17565,N_12750,N_12968);
nor U17566 (N_17566,N_14945,N_14614);
xor U17567 (N_17567,N_14090,N_15416);
nor U17568 (N_17568,N_12948,N_12888);
and U17569 (N_17569,N_14826,N_15374);
xnor U17570 (N_17570,N_13102,N_14113);
and U17571 (N_17571,N_13076,N_14279);
nor U17572 (N_17572,N_15368,N_12982);
and U17573 (N_17573,N_14378,N_12700);
nor U17574 (N_17574,N_13477,N_13345);
nor U17575 (N_17575,N_12541,N_12678);
or U17576 (N_17576,N_14452,N_14861);
xor U17577 (N_17577,N_13604,N_12719);
and U17578 (N_17578,N_14023,N_15033);
or U17579 (N_17579,N_15230,N_12637);
and U17580 (N_17580,N_15276,N_14877);
nand U17581 (N_17581,N_12522,N_14756);
nand U17582 (N_17582,N_15366,N_12874);
or U17583 (N_17583,N_12811,N_12568);
nand U17584 (N_17584,N_13152,N_15059);
xor U17585 (N_17585,N_13748,N_13389);
nand U17586 (N_17586,N_13648,N_13271);
nand U17587 (N_17587,N_15525,N_13359);
and U17588 (N_17588,N_14860,N_14525);
and U17589 (N_17589,N_14667,N_12834);
xor U17590 (N_17590,N_12547,N_14667);
nor U17591 (N_17591,N_13430,N_15208);
and U17592 (N_17592,N_12785,N_14992);
and U17593 (N_17593,N_12845,N_12704);
nand U17594 (N_17594,N_13808,N_13343);
and U17595 (N_17595,N_14230,N_12833);
nand U17596 (N_17596,N_12595,N_12707);
nor U17597 (N_17597,N_12794,N_13659);
xnor U17598 (N_17598,N_14940,N_14427);
xnor U17599 (N_17599,N_14161,N_15219);
nand U17600 (N_17600,N_14956,N_14712);
and U17601 (N_17601,N_13307,N_14903);
nand U17602 (N_17602,N_13895,N_14120);
and U17603 (N_17603,N_13769,N_13445);
nor U17604 (N_17604,N_14351,N_13879);
or U17605 (N_17605,N_12508,N_13541);
nand U17606 (N_17606,N_14496,N_13103);
and U17607 (N_17607,N_14302,N_12834);
and U17608 (N_17608,N_14342,N_14975);
and U17609 (N_17609,N_13910,N_15364);
nor U17610 (N_17610,N_14715,N_13473);
and U17611 (N_17611,N_13330,N_15464);
xor U17612 (N_17612,N_14207,N_13290);
and U17613 (N_17613,N_12945,N_15193);
xor U17614 (N_17614,N_15058,N_15097);
nor U17615 (N_17615,N_13179,N_13036);
and U17616 (N_17616,N_12602,N_13749);
nor U17617 (N_17617,N_14368,N_13115);
nor U17618 (N_17618,N_14941,N_14949);
and U17619 (N_17619,N_14250,N_13746);
or U17620 (N_17620,N_13997,N_12584);
and U17621 (N_17621,N_12990,N_13790);
nand U17622 (N_17622,N_14241,N_15090);
or U17623 (N_17623,N_14533,N_13222);
and U17624 (N_17624,N_15253,N_13711);
xnor U17625 (N_17625,N_14866,N_13733);
nand U17626 (N_17626,N_14011,N_14032);
nor U17627 (N_17627,N_13689,N_13825);
or U17628 (N_17628,N_13903,N_14151);
nor U17629 (N_17629,N_15565,N_14740);
or U17630 (N_17630,N_14463,N_14671);
nor U17631 (N_17631,N_15391,N_15238);
nand U17632 (N_17632,N_15172,N_14881);
and U17633 (N_17633,N_12914,N_15573);
nand U17634 (N_17634,N_14972,N_13411);
nor U17635 (N_17635,N_14808,N_14023);
nand U17636 (N_17636,N_12918,N_13285);
nand U17637 (N_17637,N_13631,N_13067);
or U17638 (N_17638,N_13258,N_15341);
xnor U17639 (N_17639,N_12919,N_14177);
or U17640 (N_17640,N_14052,N_14494);
xor U17641 (N_17641,N_14796,N_13320);
or U17642 (N_17642,N_14629,N_13820);
and U17643 (N_17643,N_13985,N_15611);
nand U17644 (N_17644,N_13385,N_13066);
xnor U17645 (N_17645,N_15093,N_13503);
xnor U17646 (N_17646,N_15150,N_12519);
or U17647 (N_17647,N_13729,N_12661);
nor U17648 (N_17648,N_13078,N_15182);
or U17649 (N_17649,N_15230,N_13173);
or U17650 (N_17650,N_14538,N_14266);
nor U17651 (N_17651,N_14101,N_13339);
nor U17652 (N_17652,N_14445,N_15420);
nand U17653 (N_17653,N_13998,N_15547);
nor U17654 (N_17654,N_14424,N_12899);
and U17655 (N_17655,N_14175,N_13914);
xor U17656 (N_17656,N_15492,N_13656);
or U17657 (N_17657,N_14341,N_15327);
xnor U17658 (N_17658,N_14239,N_12720);
xor U17659 (N_17659,N_14430,N_13956);
nor U17660 (N_17660,N_14835,N_13190);
nand U17661 (N_17661,N_15560,N_15375);
or U17662 (N_17662,N_13232,N_14564);
and U17663 (N_17663,N_12765,N_13453);
or U17664 (N_17664,N_15149,N_13891);
and U17665 (N_17665,N_15524,N_12519);
or U17666 (N_17666,N_13806,N_12843);
nand U17667 (N_17667,N_12731,N_12892);
xnor U17668 (N_17668,N_15394,N_12836);
nand U17669 (N_17669,N_15150,N_13652);
xor U17670 (N_17670,N_12965,N_15504);
nor U17671 (N_17671,N_14241,N_13337);
or U17672 (N_17672,N_14997,N_15085);
and U17673 (N_17673,N_15356,N_12974);
nand U17674 (N_17674,N_14026,N_13506);
and U17675 (N_17675,N_13993,N_15021);
or U17676 (N_17676,N_14051,N_12556);
nand U17677 (N_17677,N_13459,N_14380);
nand U17678 (N_17678,N_15369,N_15509);
and U17679 (N_17679,N_13482,N_14437);
or U17680 (N_17680,N_13125,N_13070);
and U17681 (N_17681,N_15218,N_12765);
and U17682 (N_17682,N_14295,N_14445);
nor U17683 (N_17683,N_13662,N_15189);
or U17684 (N_17684,N_12976,N_14619);
or U17685 (N_17685,N_14613,N_14927);
nor U17686 (N_17686,N_12921,N_15205);
or U17687 (N_17687,N_15300,N_13347);
or U17688 (N_17688,N_13230,N_14278);
nor U17689 (N_17689,N_14975,N_13666);
and U17690 (N_17690,N_13540,N_12954);
and U17691 (N_17691,N_14127,N_13396);
nor U17692 (N_17692,N_13905,N_13696);
nand U17693 (N_17693,N_14881,N_14513);
nor U17694 (N_17694,N_13869,N_14105);
nor U17695 (N_17695,N_14829,N_12908);
and U17696 (N_17696,N_12840,N_15305);
nor U17697 (N_17697,N_15363,N_13667);
or U17698 (N_17698,N_13971,N_13328);
or U17699 (N_17699,N_15314,N_15515);
or U17700 (N_17700,N_13971,N_13853);
nor U17701 (N_17701,N_13439,N_13605);
nor U17702 (N_17702,N_14001,N_15431);
and U17703 (N_17703,N_12538,N_12572);
xor U17704 (N_17704,N_13948,N_14954);
xor U17705 (N_17705,N_13438,N_14523);
and U17706 (N_17706,N_13496,N_13304);
and U17707 (N_17707,N_15465,N_14726);
xor U17708 (N_17708,N_13883,N_15573);
nand U17709 (N_17709,N_13545,N_12575);
xnor U17710 (N_17710,N_13756,N_14789);
and U17711 (N_17711,N_14382,N_13890);
and U17712 (N_17712,N_15570,N_14298);
and U17713 (N_17713,N_13012,N_12663);
or U17714 (N_17714,N_15481,N_13178);
xnor U17715 (N_17715,N_15350,N_14481);
or U17716 (N_17716,N_14405,N_15245);
xor U17717 (N_17717,N_15182,N_13505);
or U17718 (N_17718,N_14153,N_12718);
xnor U17719 (N_17719,N_14862,N_14931);
and U17720 (N_17720,N_14256,N_14854);
and U17721 (N_17721,N_13719,N_13168);
xnor U17722 (N_17722,N_13756,N_13757);
xnor U17723 (N_17723,N_12823,N_14289);
nand U17724 (N_17724,N_13650,N_15528);
or U17725 (N_17725,N_14542,N_12532);
nand U17726 (N_17726,N_12602,N_13282);
nor U17727 (N_17727,N_14303,N_14002);
and U17728 (N_17728,N_14882,N_12540);
and U17729 (N_17729,N_15482,N_14937);
nand U17730 (N_17730,N_13515,N_14830);
nor U17731 (N_17731,N_15203,N_14562);
or U17732 (N_17732,N_15042,N_14999);
and U17733 (N_17733,N_12608,N_12986);
or U17734 (N_17734,N_14712,N_14468);
xor U17735 (N_17735,N_14587,N_15302);
or U17736 (N_17736,N_13484,N_15512);
and U17737 (N_17737,N_12870,N_15613);
or U17738 (N_17738,N_12983,N_14103);
xnor U17739 (N_17739,N_15232,N_14123);
nor U17740 (N_17740,N_14925,N_13388);
nand U17741 (N_17741,N_12815,N_13014);
nand U17742 (N_17742,N_14514,N_14175);
nand U17743 (N_17743,N_13659,N_13168);
xor U17744 (N_17744,N_13671,N_13750);
xnor U17745 (N_17745,N_13752,N_13648);
nor U17746 (N_17746,N_14557,N_12675);
nand U17747 (N_17747,N_15374,N_13308);
nor U17748 (N_17748,N_14376,N_14741);
nor U17749 (N_17749,N_13115,N_14284);
and U17750 (N_17750,N_14955,N_12626);
nor U17751 (N_17751,N_15156,N_13524);
nor U17752 (N_17752,N_14927,N_12712);
or U17753 (N_17753,N_12503,N_12655);
xor U17754 (N_17754,N_14823,N_13900);
and U17755 (N_17755,N_13381,N_14487);
and U17756 (N_17756,N_15428,N_14789);
and U17757 (N_17757,N_12858,N_14374);
nor U17758 (N_17758,N_13624,N_15556);
nand U17759 (N_17759,N_13839,N_13028);
xnor U17760 (N_17760,N_14262,N_13079);
nand U17761 (N_17761,N_13445,N_15005);
nand U17762 (N_17762,N_14901,N_14736);
nor U17763 (N_17763,N_15187,N_15412);
nand U17764 (N_17764,N_15610,N_13978);
xor U17765 (N_17765,N_15282,N_14066);
nand U17766 (N_17766,N_13265,N_13721);
or U17767 (N_17767,N_15435,N_14907);
nor U17768 (N_17768,N_12556,N_12641);
nand U17769 (N_17769,N_14760,N_15386);
and U17770 (N_17770,N_12971,N_14089);
and U17771 (N_17771,N_15559,N_13795);
or U17772 (N_17772,N_12572,N_12580);
nand U17773 (N_17773,N_12999,N_14983);
or U17774 (N_17774,N_13580,N_15188);
xnor U17775 (N_17775,N_12574,N_13076);
nand U17776 (N_17776,N_14604,N_15559);
xnor U17777 (N_17777,N_13742,N_13724);
nor U17778 (N_17778,N_12879,N_14197);
or U17779 (N_17779,N_13346,N_15124);
and U17780 (N_17780,N_15517,N_13250);
xnor U17781 (N_17781,N_14896,N_14433);
xor U17782 (N_17782,N_15059,N_14659);
xor U17783 (N_17783,N_13276,N_14534);
nand U17784 (N_17784,N_12799,N_15060);
and U17785 (N_17785,N_14270,N_14039);
and U17786 (N_17786,N_15525,N_13936);
nand U17787 (N_17787,N_13947,N_12671);
xor U17788 (N_17788,N_13021,N_15133);
or U17789 (N_17789,N_14457,N_15556);
nor U17790 (N_17790,N_12768,N_12842);
or U17791 (N_17791,N_15004,N_13814);
nor U17792 (N_17792,N_14633,N_12926);
xnor U17793 (N_17793,N_14434,N_13797);
or U17794 (N_17794,N_15359,N_14625);
nand U17795 (N_17795,N_13569,N_13558);
and U17796 (N_17796,N_13843,N_13221);
nand U17797 (N_17797,N_15353,N_15573);
nor U17798 (N_17798,N_13013,N_12592);
and U17799 (N_17799,N_15586,N_13704);
or U17800 (N_17800,N_15557,N_14444);
xor U17801 (N_17801,N_14879,N_13266);
or U17802 (N_17802,N_15465,N_13262);
xor U17803 (N_17803,N_14553,N_12851);
nand U17804 (N_17804,N_14627,N_13118);
nand U17805 (N_17805,N_15457,N_12635);
nor U17806 (N_17806,N_13502,N_13524);
nor U17807 (N_17807,N_13755,N_14156);
and U17808 (N_17808,N_12943,N_14346);
and U17809 (N_17809,N_14687,N_12641);
and U17810 (N_17810,N_15607,N_15577);
and U17811 (N_17811,N_14396,N_14341);
xnor U17812 (N_17812,N_15026,N_15472);
xnor U17813 (N_17813,N_15074,N_13346);
nor U17814 (N_17814,N_14770,N_13329);
nand U17815 (N_17815,N_14310,N_13349);
nor U17816 (N_17816,N_14362,N_15135);
nor U17817 (N_17817,N_14089,N_13447);
and U17818 (N_17818,N_13265,N_13112);
nand U17819 (N_17819,N_15424,N_13420);
xor U17820 (N_17820,N_14190,N_12829);
nor U17821 (N_17821,N_14253,N_13454);
and U17822 (N_17822,N_14754,N_14820);
or U17823 (N_17823,N_15525,N_12919);
nand U17824 (N_17824,N_14513,N_13687);
nand U17825 (N_17825,N_13883,N_13868);
or U17826 (N_17826,N_13807,N_15100);
nand U17827 (N_17827,N_13553,N_14743);
nand U17828 (N_17828,N_14207,N_14929);
or U17829 (N_17829,N_15176,N_12698);
xnor U17830 (N_17830,N_14274,N_14521);
or U17831 (N_17831,N_13281,N_13634);
nor U17832 (N_17832,N_13580,N_14341);
or U17833 (N_17833,N_14507,N_12904);
nand U17834 (N_17834,N_12543,N_12785);
xor U17835 (N_17835,N_13939,N_15288);
xor U17836 (N_17836,N_14832,N_15168);
or U17837 (N_17837,N_13626,N_13656);
and U17838 (N_17838,N_13540,N_15485);
and U17839 (N_17839,N_13034,N_15458);
xor U17840 (N_17840,N_14357,N_14998);
nand U17841 (N_17841,N_12703,N_12974);
nor U17842 (N_17842,N_14800,N_13441);
nor U17843 (N_17843,N_12900,N_14124);
nand U17844 (N_17844,N_13401,N_13632);
nand U17845 (N_17845,N_14519,N_12710);
nor U17846 (N_17846,N_14682,N_13098);
nand U17847 (N_17847,N_12759,N_15046);
xor U17848 (N_17848,N_12606,N_15404);
xnor U17849 (N_17849,N_14656,N_14391);
nand U17850 (N_17850,N_14031,N_14264);
and U17851 (N_17851,N_14906,N_15374);
nand U17852 (N_17852,N_15057,N_15218);
and U17853 (N_17853,N_13295,N_14382);
nand U17854 (N_17854,N_13626,N_15481);
nor U17855 (N_17855,N_13401,N_14333);
nor U17856 (N_17856,N_14275,N_13452);
or U17857 (N_17857,N_15017,N_13174);
or U17858 (N_17858,N_13214,N_15256);
xor U17859 (N_17859,N_14572,N_14760);
nand U17860 (N_17860,N_15368,N_14361);
and U17861 (N_17861,N_13797,N_14450);
nor U17862 (N_17862,N_13329,N_14630);
xor U17863 (N_17863,N_15474,N_12621);
nand U17864 (N_17864,N_13724,N_14990);
or U17865 (N_17865,N_14452,N_12601);
or U17866 (N_17866,N_14099,N_13299);
or U17867 (N_17867,N_14992,N_13942);
and U17868 (N_17868,N_15386,N_13237);
nor U17869 (N_17869,N_13010,N_14768);
nor U17870 (N_17870,N_15502,N_13904);
and U17871 (N_17871,N_13776,N_13780);
or U17872 (N_17872,N_12653,N_14047);
or U17873 (N_17873,N_13684,N_13061);
xnor U17874 (N_17874,N_13781,N_13146);
and U17875 (N_17875,N_13502,N_15105);
or U17876 (N_17876,N_15435,N_13037);
nand U17877 (N_17877,N_14942,N_14190);
and U17878 (N_17878,N_14383,N_15492);
and U17879 (N_17879,N_12954,N_14599);
xnor U17880 (N_17880,N_15315,N_13536);
xor U17881 (N_17881,N_14037,N_13265);
or U17882 (N_17882,N_14270,N_13516);
or U17883 (N_17883,N_13736,N_12918);
nand U17884 (N_17884,N_12780,N_13694);
nand U17885 (N_17885,N_12721,N_15476);
nand U17886 (N_17886,N_14481,N_15235);
xnor U17887 (N_17887,N_12746,N_13491);
or U17888 (N_17888,N_12632,N_14668);
nand U17889 (N_17889,N_13384,N_12832);
nand U17890 (N_17890,N_14881,N_14901);
or U17891 (N_17891,N_14613,N_14427);
or U17892 (N_17892,N_15238,N_15594);
or U17893 (N_17893,N_13097,N_14752);
xor U17894 (N_17894,N_14177,N_12918);
xor U17895 (N_17895,N_12901,N_13737);
or U17896 (N_17896,N_14781,N_13964);
nor U17897 (N_17897,N_15624,N_14924);
nand U17898 (N_17898,N_12902,N_13402);
nand U17899 (N_17899,N_12837,N_13899);
xor U17900 (N_17900,N_14095,N_14631);
nor U17901 (N_17901,N_13082,N_15124);
nor U17902 (N_17902,N_15453,N_13653);
xnor U17903 (N_17903,N_15421,N_14745);
or U17904 (N_17904,N_15257,N_13433);
xor U17905 (N_17905,N_12625,N_13136);
nor U17906 (N_17906,N_13963,N_15283);
or U17907 (N_17907,N_14350,N_14169);
xor U17908 (N_17908,N_12603,N_14699);
nand U17909 (N_17909,N_12709,N_13036);
or U17910 (N_17910,N_15344,N_14016);
or U17911 (N_17911,N_13181,N_13895);
and U17912 (N_17912,N_15277,N_13530);
and U17913 (N_17913,N_13363,N_13100);
nand U17914 (N_17914,N_14798,N_14498);
xnor U17915 (N_17915,N_14424,N_15169);
or U17916 (N_17916,N_14433,N_15501);
or U17917 (N_17917,N_15274,N_15567);
xor U17918 (N_17918,N_14813,N_14115);
nor U17919 (N_17919,N_14285,N_14810);
or U17920 (N_17920,N_14779,N_13818);
and U17921 (N_17921,N_14129,N_14402);
or U17922 (N_17922,N_13276,N_13840);
xnor U17923 (N_17923,N_12596,N_14277);
or U17924 (N_17924,N_14230,N_15251);
or U17925 (N_17925,N_13680,N_14842);
or U17926 (N_17926,N_14256,N_12858);
and U17927 (N_17927,N_14214,N_15208);
or U17928 (N_17928,N_15370,N_12876);
nand U17929 (N_17929,N_13044,N_15501);
nor U17930 (N_17930,N_14228,N_13183);
or U17931 (N_17931,N_14542,N_13704);
and U17932 (N_17932,N_13855,N_15166);
xor U17933 (N_17933,N_13447,N_13045);
xnor U17934 (N_17934,N_12507,N_15381);
and U17935 (N_17935,N_15090,N_15048);
nand U17936 (N_17936,N_13941,N_14932);
xnor U17937 (N_17937,N_15565,N_15215);
or U17938 (N_17938,N_14010,N_12697);
xnor U17939 (N_17939,N_15270,N_13609);
nor U17940 (N_17940,N_15351,N_13694);
xor U17941 (N_17941,N_14606,N_14352);
nor U17942 (N_17942,N_14185,N_14928);
nor U17943 (N_17943,N_12894,N_13762);
or U17944 (N_17944,N_12827,N_14810);
and U17945 (N_17945,N_14922,N_14160);
xor U17946 (N_17946,N_12697,N_14423);
or U17947 (N_17947,N_14033,N_13393);
nor U17948 (N_17948,N_14499,N_13459);
xnor U17949 (N_17949,N_14029,N_13763);
or U17950 (N_17950,N_14473,N_15295);
nand U17951 (N_17951,N_14423,N_15198);
and U17952 (N_17952,N_14180,N_12525);
nand U17953 (N_17953,N_14313,N_14405);
xnor U17954 (N_17954,N_15027,N_14465);
and U17955 (N_17955,N_15435,N_12590);
and U17956 (N_17956,N_13133,N_14548);
xnor U17957 (N_17957,N_12797,N_14651);
or U17958 (N_17958,N_13687,N_14869);
xor U17959 (N_17959,N_14302,N_12854);
and U17960 (N_17960,N_15019,N_13269);
nor U17961 (N_17961,N_13105,N_13835);
nand U17962 (N_17962,N_12699,N_15049);
or U17963 (N_17963,N_14072,N_14583);
and U17964 (N_17964,N_12999,N_14073);
nand U17965 (N_17965,N_14879,N_14525);
xor U17966 (N_17966,N_13055,N_14794);
and U17967 (N_17967,N_14309,N_13080);
xor U17968 (N_17968,N_15105,N_15350);
and U17969 (N_17969,N_14750,N_14087);
nor U17970 (N_17970,N_13791,N_13803);
xnor U17971 (N_17971,N_13005,N_12669);
xor U17972 (N_17972,N_15365,N_13400);
nor U17973 (N_17973,N_14595,N_13280);
nand U17974 (N_17974,N_14275,N_15620);
xnor U17975 (N_17975,N_13808,N_13453);
xnor U17976 (N_17976,N_15202,N_15300);
nor U17977 (N_17977,N_14662,N_13266);
xor U17978 (N_17978,N_14122,N_14115);
nor U17979 (N_17979,N_12572,N_12520);
and U17980 (N_17980,N_13836,N_12940);
nand U17981 (N_17981,N_14859,N_15211);
and U17982 (N_17982,N_15518,N_14997);
or U17983 (N_17983,N_12870,N_14490);
and U17984 (N_17984,N_13233,N_14980);
nor U17985 (N_17985,N_12980,N_14426);
nor U17986 (N_17986,N_14936,N_13737);
nand U17987 (N_17987,N_15134,N_14189);
nor U17988 (N_17988,N_15616,N_14159);
nand U17989 (N_17989,N_14238,N_12563);
and U17990 (N_17990,N_13404,N_13205);
and U17991 (N_17991,N_14987,N_12568);
xnor U17992 (N_17992,N_15273,N_14011);
and U17993 (N_17993,N_14691,N_12511);
or U17994 (N_17994,N_14218,N_12963);
xnor U17995 (N_17995,N_15399,N_12940);
nand U17996 (N_17996,N_15016,N_14776);
or U17997 (N_17997,N_14376,N_13683);
nand U17998 (N_17998,N_12516,N_13689);
xor U17999 (N_17999,N_12844,N_15076);
or U18000 (N_18000,N_14159,N_13896);
and U18001 (N_18001,N_15396,N_13807);
and U18002 (N_18002,N_13312,N_13463);
nand U18003 (N_18003,N_12727,N_13633);
or U18004 (N_18004,N_14045,N_13624);
xor U18005 (N_18005,N_13556,N_13211);
or U18006 (N_18006,N_13864,N_13884);
nor U18007 (N_18007,N_14592,N_13335);
nor U18008 (N_18008,N_14127,N_15465);
nor U18009 (N_18009,N_14136,N_14237);
xnor U18010 (N_18010,N_14608,N_12738);
xor U18011 (N_18011,N_15340,N_13057);
nand U18012 (N_18012,N_14753,N_15274);
xnor U18013 (N_18013,N_15330,N_15621);
nand U18014 (N_18014,N_14606,N_12874);
and U18015 (N_18015,N_13132,N_13218);
or U18016 (N_18016,N_14426,N_15294);
and U18017 (N_18017,N_15376,N_14115);
and U18018 (N_18018,N_13977,N_12827);
and U18019 (N_18019,N_15602,N_12972);
or U18020 (N_18020,N_14423,N_13640);
nand U18021 (N_18021,N_15137,N_13798);
xnor U18022 (N_18022,N_14690,N_12771);
xnor U18023 (N_18023,N_14496,N_14843);
and U18024 (N_18024,N_12701,N_15074);
and U18025 (N_18025,N_15249,N_14551);
nor U18026 (N_18026,N_12905,N_12783);
or U18027 (N_18027,N_13156,N_12592);
or U18028 (N_18028,N_14987,N_15321);
nand U18029 (N_18029,N_12599,N_13391);
nand U18030 (N_18030,N_15045,N_14550);
nor U18031 (N_18031,N_13484,N_14750);
or U18032 (N_18032,N_14047,N_14247);
or U18033 (N_18033,N_15418,N_14656);
nand U18034 (N_18034,N_14184,N_15513);
nor U18035 (N_18035,N_15047,N_15390);
or U18036 (N_18036,N_14408,N_15382);
nor U18037 (N_18037,N_14378,N_13432);
nand U18038 (N_18038,N_14103,N_14330);
and U18039 (N_18039,N_12977,N_13944);
nand U18040 (N_18040,N_15067,N_12823);
xor U18041 (N_18041,N_13618,N_13803);
and U18042 (N_18042,N_12878,N_14023);
nand U18043 (N_18043,N_14979,N_15493);
or U18044 (N_18044,N_13499,N_12813);
xor U18045 (N_18045,N_15399,N_13283);
nand U18046 (N_18046,N_12554,N_15407);
nand U18047 (N_18047,N_12847,N_13849);
or U18048 (N_18048,N_12876,N_13965);
nand U18049 (N_18049,N_13619,N_14988);
or U18050 (N_18050,N_13609,N_15547);
nor U18051 (N_18051,N_12782,N_12594);
xor U18052 (N_18052,N_13292,N_15405);
or U18053 (N_18053,N_12896,N_15476);
nor U18054 (N_18054,N_12826,N_14800);
nand U18055 (N_18055,N_15315,N_14271);
nor U18056 (N_18056,N_13180,N_12951);
or U18057 (N_18057,N_14835,N_13920);
xnor U18058 (N_18058,N_15059,N_13189);
nor U18059 (N_18059,N_13981,N_14926);
xnor U18060 (N_18060,N_12852,N_14427);
xnor U18061 (N_18061,N_14073,N_15617);
xor U18062 (N_18062,N_15025,N_15429);
nand U18063 (N_18063,N_13025,N_15446);
nor U18064 (N_18064,N_15305,N_13564);
or U18065 (N_18065,N_14594,N_12632);
xor U18066 (N_18066,N_13044,N_14545);
nand U18067 (N_18067,N_14420,N_14288);
or U18068 (N_18068,N_13027,N_12578);
or U18069 (N_18069,N_13435,N_14996);
nand U18070 (N_18070,N_14165,N_13778);
nand U18071 (N_18071,N_12620,N_14849);
nand U18072 (N_18072,N_12742,N_14981);
or U18073 (N_18073,N_12966,N_13394);
nor U18074 (N_18074,N_14116,N_13301);
or U18075 (N_18075,N_13331,N_13176);
or U18076 (N_18076,N_14355,N_15100);
and U18077 (N_18077,N_15556,N_15495);
or U18078 (N_18078,N_15351,N_15543);
and U18079 (N_18079,N_15513,N_12639);
and U18080 (N_18080,N_13109,N_12785);
or U18081 (N_18081,N_13710,N_13690);
and U18082 (N_18082,N_13980,N_15555);
nand U18083 (N_18083,N_14259,N_12901);
nor U18084 (N_18084,N_13677,N_13175);
nor U18085 (N_18085,N_14272,N_13592);
and U18086 (N_18086,N_14797,N_14009);
or U18087 (N_18087,N_12787,N_12790);
or U18088 (N_18088,N_12506,N_14389);
nor U18089 (N_18089,N_13866,N_13254);
or U18090 (N_18090,N_13931,N_14800);
nor U18091 (N_18091,N_14100,N_15195);
nor U18092 (N_18092,N_15172,N_14085);
nor U18093 (N_18093,N_12634,N_14900);
or U18094 (N_18094,N_14640,N_12954);
nand U18095 (N_18095,N_13385,N_13458);
xor U18096 (N_18096,N_15142,N_12904);
nor U18097 (N_18097,N_15016,N_13417);
or U18098 (N_18098,N_13678,N_13725);
or U18099 (N_18099,N_14618,N_14239);
nor U18100 (N_18100,N_15537,N_14098);
xnor U18101 (N_18101,N_13180,N_12626);
xor U18102 (N_18102,N_13137,N_13253);
nor U18103 (N_18103,N_13732,N_13280);
nand U18104 (N_18104,N_15170,N_14435);
and U18105 (N_18105,N_13565,N_14568);
and U18106 (N_18106,N_14756,N_12565);
and U18107 (N_18107,N_13646,N_15561);
nor U18108 (N_18108,N_15071,N_14543);
nand U18109 (N_18109,N_15413,N_14300);
or U18110 (N_18110,N_13176,N_13059);
nand U18111 (N_18111,N_13968,N_13037);
xnor U18112 (N_18112,N_12866,N_12904);
nand U18113 (N_18113,N_14808,N_14371);
nand U18114 (N_18114,N_13878,N_13872);
or U18115 (N_18115,N_12997,N_12859);
or U18116 (N_18116,N_12605,N_13504);
xor U18117 (N_18117,N_13828,N_14245);
nor U18118 (N_18118,N_15323,N_12989);
nand U18119 (N_18119,N_15228,N_14872);
nor U18120 (N_18120,N_12626,N_12585);
xor U18121 (N_18121,N_14134,N_15282);
nand U18122 (N_18122,N_14286,N_13906);
xnor U18123 (N_18123,N_14451,N_15276);
or U18124 (N_18124,N_14471,N_14800);
or U18125 (N_18125,N_12644,N_13434);
nor U18126 (N_18126,N_13717,N_15591);
nor U18127 (N_18127,N_12781,N_14265);
xnor U18128 (N_18128,N_13205,N_13249);
or U18129 (N_18129,N_15177,N_13185);
and U18130 (N_18130,N_13039,N_15292);
nand U18131 (N_18131,N_14819,N_13473);
nand U18132 (N_18132,N_13223,N_13662);
nand U18133 (N_18133,N_14446,N_13607);
nor U18134 (N_18134,N_14805,N_14546);
and U18135 (N_18135,N_14486,N_12733);
and U18136 (N_18136,N_15557,N_13114);
and U18137 (N_18137,N_15191,N_13038);
and U18138 (N_18138,N_15104,N_13606);
or U18139 (N_18139,N_15453,N_14948);
xor U18140 (N_18140,N_13349,N_13020);
nor U18141 (N_18141,N_14210,N_15342);
nor U18142 (N_18142,N_14499,N_13709);
xnor U18143 (N_18143,N_12925,N_12726);
nand U18144 (N_18144,N_15475,N_14336);
or U18145 (N_18145,N_13762,N_12538);
xnor U18146 (N_18146,N_13660,N_12808);
nor U18147 (N_18147,N_13274,N_14897);
nor U18148 (N_18148,N_14385,N_14047);
xor U18149 (N_18149,N_13358,N_12692);
nor U18150 (N_18150,N_14758,N_12885);
nor U18151 (N_18151,N_13631,N_13436);
nor U18152 (N_18152,N_14101,N_13521);
and U18153 (N_18153,N_13373,N_14615);
or U18154 (N_18154,N_15233,N_13859);
or U18155 (N_18155,N_15117,N_12718);
nand U18156 (N_18156,N_13014,N_14693);
nand U18157 (N_18157,N_15506,N_14389);
nand U18158 (N_18158,N_13251,N_13973);
xnor U18159 (N_18159,N_14756,N_12876);
or U18160 (N_18160,N_13291,N_15270);
or U18161 (N_18161,N_14716,N_15140);
or U18162 (N_18162,N_15579,N_14901);
and U18163 (N_18163,N_14500,N_12505);
nor U18164 (N_18164,N_15618,N_13782);
and U18165 (N_18165,N_13972,N_13879);
and U18166 (N_18166,N_14369,N_14694);
nand U18167 (N_18167,N_13210,N_13461);
and U18168 (N_18168,N_12751,N_13291);
xnor U18169 (N_18169,N_13755,N_13701);
and U18170 (N_18170,N_14948,N_12766);
or U18171 (N_18171,N_14334,N_14004);
nor U18172 (N_18172,N_12907,N_14909);
xnor U18173 (N_18173,N_15393,N_15128);
xnor U18174 (N_18174,N_15338,N_13279);
and U18175 (N_18175,N_13944,N_12605);
nand U18176 (N_18176,N_13210,N_15260);
or U18177 (N_18177,N_13223,N_14982);
or U18178 (N_18178,N_15406,N_15384);
or U18179 (N_18179,N_14624,N_15236);
and U18180 (N_18180,N_14084,N_14740);
or U18181 (N_18181,N_14184,N_13257);
xnor U18182 (N_18182,N_15031,N_15020);
nand U18183 (N_18183,N_15382,N_13471);
nor U18184 (N_18184,N_12714,N_12984);
nand U18185 (N_18185,N_12664,N_14834);
xor U18186 (N_18186,N_13289,N_14568);
and U18187 (N_18187,N_15260,N_14926);
or U18188 (N_18188,N_14486,N_15599);
nor U18189 (N_18189,N_13558,N_14837);
xor U18190 (N_18190,N_14592,N_15134);
and U18191 (N_18191,N_14798,N_12619);
nand U18192 (N_18192,N_14163,N_13756);
xor U18193 (N_18193,N_12849,N_15254);
nand U18194 (N_18194,N_15009,N_14647);
xor U18195 (N_18195,N_13713,N_15061);
nand U18196 (N_18196,N_14990,N_14861);
nand U18197 (N_18197,N_13924,N_15181);
and U18198 (N_18198,N_14063,N_14058);
and U18199 (N_18199,N_12685,N_12940);
xnor U18200 (N_18200,N_14855,N_15573);
nor U18201 (N_18201,N_13715,N_12861);
xor U18202 (N_18202,N_12704,N_14556);
and U18203 (N_18203,N_13525,N_14357);
nand U18204 (N_18204,N_13175,N_15117);
nand U18205 (N_18205,N_13408,N_12732);
nor U18206 (N_18206,N_15578,N_14203);
and U18207 (N_18207,N_14650,N_14637);
xor U18208 (N_18208,N_13045,N_12872);
nor U18209 (N_18209,N_12914,N_15460);
and U18210 (N_18210,N_15606,N_13570);
nand U18211 (N_18211,N_13401,N_12568);
nor U18212 (N_18212,N_14762,N_13456);
and U18213 (N_18213,N_12940,N_12528);
or U18214 (N_18214,N_14868,N_13359);
and U18215 (N_18215,N_14351,N_14804);
xnor U18216 (N_18216,N_15189,N_13654);
and U18217 (N_18217,N_14531,N_12825);
xor U18218 (N_18218,N_14423,N_13134);
nand U18219 (N_18219,N_12539,N_14243);
nand U18220 (N_18220,N_14631,N_15568);
nand U18221 (N_18221,N_14319,N_13620);
xnor U18222 (N_18222,N_13190,N_13421);
nand U18223 (N_18223,N_13973,N_15307);
and U18224 (N_18224,N_15447,N_15002);
nor U18225 (N_18225,N_14432,N_12521);
nor U18226 (N_18226,N_15551,N_14127);
nor U18227 (N_18227,N_14286,N_13731);
xnor U18228 (N_18228,N_15137,N_14416);
and U18229 (N_18229,N_13850,N_13368);
nor U18230 (N_18230,N_13351,N_12699);
nor U18231 (N_18231,N_13020,N_14690);
or U18232 (N_18232,N_12980,N_14408);
xor U18233 (N_18233,N_14090,N_12564);
nand U18234 (N_18234,N_15024,N_12614);
and U18235 (N_18235,N_13673,N_12633);
nor U18236 (N_18236,N_15271,N_12606);
or U18237 (N_18237,N_13580,N_13174);
and U18238 (N_18238,N_15323,N_14087);
nand U18239 (N_18239,N_15154,N_13871);
nand U18240 (N_18240,N_13429,N_15065);
nand U18241 (N_18241,N_12856,N_14114);
xor U18242 (N_18242,N_13791,N_15019);
nor U18243 (N_18243,N_13697,N_14732);
or U18244 (N_18244,N_13715,N_14672);
and U18245 (N_18245,N_13344,N_14808);
and U18246 (N_18246,N_13904,N_15227);
nand U18247 (N_18247,N_14571,N_12585);
nand U18248 (N_18248,N_12781,N_13238);
xnor U18249 (N_18249,N_13077,N_14806);
nor U18250 (N_18250,N_14306,N_13277);
and U18251 (N_18251,N_13116,N_12933);
xor U18252 (N_18252,N_15238,N_13267);
xnor U18253 (N_18253,N_13929,N_15056);
or U18254 (N_18254,N_12695,N_13646);
or U18255 (N_18255,N_15161,N_14398);
nor U18256 (N_18256,N_14806,N_14105);
nor U18257 (N_18257,N_13703,N_15253);
xor U18258 (N_18258,N_14034,N_15553);
and U18259 (N_18259,N_13889,N_13011);
or U18260 (N_18260,N_12936,N_13018);
nor U18261 (N_18261,N_13761,N_14759);
or U18262 (N_18262,N_13466,N_13706);
nand U18263 (N_18263,N_14555,N_14325);
nor U18264 (N_18264,N_14419,N_15522);
nor U18265 (N_18265,N_14251,N_12546);
or U18266 (N_18266,N_15532,N_14957);
or U18267 (N_18267,N_14500,N_15594);
nor U18268 (N_18268,N_13775,N_12528);
and U18269 (N_18269,N_13527,N_13550);
and U18270 (N_18270,N_13655,N_14891);
or U18271 (N_18271,N_14411,N_15376);
or U18272 (N_18272,N_15251,N_13895);
and U18273 (N_18273,N_12806,N_13990);
nor U18274 (N_18274,N_14204,N_14686);
and U18275 (N_18275,N_14781,N_12904);
xor U18276 (N_18276,N_15573,N_15508);
and U18277 (N_18277,N_12792,N_13425);
nand U18278 (N_18278,N_12933,N_14712);
nor U18279 (N_18279,N_12842,N_14189);
nand U18280 (N_18280,N_13097,N_13014);
or U18281 (N_18281,N_13653,N_13548);
nor U18282 (N_18282,N_15280,N_15583);
nand U18283 (N_18283,N_15102,N_13412);
nor U18284 (N_18284,N_13761,N_12671);
nor U18285 (N_18285,N_14734,N_12908);
and U18286 (N_18286,N_15432,N_13000);
xnor U18287 (N_18287,N_13741,N_14433);
nor U18288 (N_18288,N_14928,N_14929);
and U18289 (N_18289,N_13933,N_14373);
and U18290 (N_18290,N_15357,N_14120);
xor U18291 (N_18291,N_13351,N_14230);
xor U18292 (N_18292,N_14383,N_14966);
xor U18293 (N_18293,N_14368,N_13827);
or U18294 (N_18294,N_14420,N_15212);
nand U18295 (N_18295,N_13043,N_14358);
or U18296 (N_18296,N_14366,N_14779);
xor U18297 (N_18297,N_13353,N_15484);
nor U18298 (N_18298,N_13515,N_12867);
and U18299 (N_18299,N_13019,N_13830);
and U18300 (N_18300,N_13259,N_15455);
nor U18301 (N_18301,N_14738,N_12560);
nand U18302 (N_18302,N_13946,N_15577);
or U18303 (N_18303,N_13128,N_14371);
xnor U18304 (N_18304,N_14163,N_14154);
or U18305 (N_18305,N_13237,N_14168);
xnor U18306 (N_18306,N_13638,N_13109);
xor U18307 (N_18307,N_14223,N_12728);
xnor U18308 (N_18308,N_12767,N_14073);
and U18309 (N_18309,N_13746,N_12522);
and U18310 (N_18310,N_15050,N_13335);
nor U18311 (N_18311,N_13372,N_13564);
or U18312 (N_18312,N_14471,N_15114);
and U18313 (N_18313,N_13836,N_15392);
xnor U18314 (N_18314,N_15312,N_12695);
nand U18315 (N_18315,N_13505,N_13144);
and U18316 (N_18316,N_12784,N_14581);
and U18317 (N_18317,N_12953,N_15320);
nor U18318 (N_18318,N_13676,N_15584);
and U18319 (N_18319,N_14994,N_14724);
and U18320 (N_18320,N_12977,N_15006);
and U18321 (N_18321,N_13587,N_15303);
xnor U18322 (N_18322,N_14431,N_13596);
or U18323 (N_18323,N_13682,N_15331);
or U18324 (N_18324,N_14437,N_14920);
xor U18325 (N_18325,N_12906,N_14552);
xor U18326 (N_18326,N_15584,N_13812);
and U18327 (N_18327,N_13771,N_12962);
and U18328 (N_18328,N_13894,N_12517);
nand U18329 (N_18329,N_12576,N_12722);
and U18330 (N_18330,N_13985,N_14683);
or U18331 (N_18331,N_13437,N_12550);
and U18332 (N_18332,N_15372,N_13366);
or U18333 (N_18333,N_13414,N_13933);
xor U18334 (N_18334,N_14750,N_15262);
nor U18335 (N_18335,N_14985,N_13097);
or U18336 (N_18336,N_14108,N_14692);
or U18337 (N_18337,N_14452,N_14977);
xnor U18338 (N_18338,N_14460,N_13732);
nand U18339 (N_18339,N_15446,N_15440);
xnor U18340 (N_18340,N_15527,N_13191);
and U18341 (N_18341,N_14353,N_14346);
nand U18342 (N_18342,N_13253,N_15258);
nor U18343 (N_18343,N_12800,N_15548);
or U18344 (N_18344,N_14844,N_15613);
or U18345 (N_18345,N_13732,N_13605);
nor U18346 (N_18346,N_14580,N_15171);
nor U18347 (N_18347,N_14886,N_12729);
nand U18348 (N_18348,N_13994,N_15139);
and U18349 (N_18349,N_14505,N_14443);
or U18350 (N_18350,N_15198,N_13257);
xor U18351 (N_18351,N_13923,N_13658);
xnor U18352 (N_18352,N_13235,N_13877);
or U18353 (N_18353,N_14604,N_15438);
or U18354 (N_18354,N_13358,N_15030);
xor U18355 (N_18355,N_14753,N_13875);
or U18356 (N_18356,N_13776,N_13304);
and U18357 (N_18357,N_13554,N_14875);
and U18358 (N_18358,N_12808,N_12502);
nand U18359 (N_18359,N_14411,N_13227);
nor U18360 (N_18360,N_13810,N_14634);
xnor U18361 (N_18361,N_13759,N_14523);
nor U18362 (N_18362,N_12812,N_15168);
nand U18363 (N_18363,N_14555,N_15447);
nand U18364 (N_18364,N_15091,N_14105);
nor U18365 (N_18365,N_15580,N_14149);
or U18366 (N_18366,N_13468,N_14688);
nand U18367 (N_18367,N_13061,N_14692);
nor U18368 (N_18368,N_14873,N_12515);
xnor U18369 (N_18369,N_12876,N_14336);
and U18370 (N_18370,N_13489,N_14043);
or U18371 (N_18371,N_15550,N_13962);
or U18372 (N_18372,N_15096,N_14135);
nand U18373 (N_18373,N_12878,N_14650);
or U18374 (N_18374,N_14664,N_13220);
xor U18375 (N_18375,N_12896,N_13218);
and U18376 (N_18376,N_14203,N_13932);
xnor U18377 (N_18377,N_14356,N_14275);
or U18378 (N_18378,N_12712,N_13613);
xnor U18379 (N_18379,N_13152,N_13550);
or U18380 (N_18380,N_15194,N_13080);
or U18381 (N_18381,N_15430,N_12940);
nor U18382 (N_18382,N_15514,N_14769);
and U18383 (N_18383,N_15424,N_15388);
or U18384 (N_18384,N_13524,N_13395);
nand U18385 (N_18385,N_15428,N_14313);
xnor U18386 (N_18386,N_13994,N_13445);
nor U18387 (N_18387,N_14304,N_13689);
nand U18388 (N_18388,N_15308,N_15048);
nand U18389 (N_18389,N_13797,N_13166);
nor U18390 (N_18390,N_12883,N_13018);
xor U18391 (N_18391,N_14761,N_13221);
nor U18392 (N_18392,N_13886,N_14989);
and U18393 (N_18393,N_13925,N_13532);
nor U18394 (N_18394,N_13058,N_15304);
xnor U18395 (N_18395,N_15109,N_12745);
or U18396 (N_18396,N_14684,N_14137);
and U18397 (N_18397,N_13927,N_12931);
nor U18398 (N_18398,N_14312,N_14214);
nand U18399 (N_18399,N_12549,N_13694);
nor U18400 (N_18400,N_13499,N_15379);
nor U18401 (N_18401,N_15506,N_15162);
nand U18402 (N_18402,N_12710,N_12796);
nand U18403 (N_18403,N_12656,N_12803);
nor U18404 (N_18404,N_15482,N_13875);
xnor U18405 (N_18405,N_15314,N_15085);
or U18406 (N_18406,N_13973,N_12772);
xor U18407 (N_18407,N_14990,N_13129);
and U18408 (N_18408,N_14384,N_15294);
and U18409 (N_18409,N_15621,N_14690);
nor U18410 (N_18410,N_14617,N_13180);
xor U18411 (N_18411,N_14281,N_14971);
xnor U18412 (N_18412,N_14301,N_15554);
or U18413 (N_18413,N_14959,N_12586);
or U18414 (N_18414,N_13667,N_15402);
nor U18415 (N_18415,N_15058,N_14776);
or U18416 (N_18416,N_14651,N_13680);
xnor U18417 (N_18417,N_13615,N_14676);
nor U18418 (N_18418,N_14668,N_12505);
or U18419 (N_18419,N_14493,N_13583);
nand U18420 (N_18420,N_13632,N_15212);
xnor U18421 (N_18421,N_14849,N_12812);
xnor U18422 (N_18422,N_13714,N_13067);
xnor U18423 (N_18423,N_14594,N_15444);
xor U18424 (N_18424,N_14654,N_15074);
or U18425 (N_18425,N_13029,N_12998);
nor U18426 (N_18426,N_12996,N_14563);
and U18427 (N_18427,N_14246,N_12685);
xnor U18428 (N_18428,N_13519,N_14188);
or U18429 (N_18429,N_13245,N_14385);
or U18430 (N_18430,N_13506,N_13867);
nand U18431 (N_18431,N_15159,N_15160);
and U18432 (N_18432,N_12534,N_15014);
xor U18433 (N_18433,N_14656,N_14196);
and U18434 (N_18434,N_15506,N_15408);
xnor U18435 (N_18435,N_15080,N_15361);
nor U18436 (N_18436,N_13362,N_13314);
and U18437 (N_18437,N_14266,N_13877);
nand U18438 (N_18438,N_14706,N_12921);
xor U18439 (N_18439,N_14875,N_13280);
nand U18440 (N_18440,N_13121,N_13655);
nor U18441 (N_18441,N_15247,N_12662);
nand U18442 (N_18442,N_15326,N_13742);
or U18443 (N_18443,N_15578,N_13841);
nor U18444 (N_18444,N_13970,N_12618);
or U18445 (N_18445,N_13037,N_14732);
or U18446 (N_18446,N_14329,N_13448);
nand U18447 (N_18447,N_15311,N_14368);
or U18448 (N_18448,N_14102,N_14285);
nor U18449 (N_18449,N_14343,N_14216);
nand U18450 (N_18450,N_15430,N_13070);
or U18451 (N_18451,N_14028,N_15037);
and U18452 (N_18452,N_13547,N_15127);
nand U18453 (N_18453,N_15474,N_15554);
nand U18454 (N_18454,N_13916,N_13848);
nor U18455 (N_18455,N_14379,N_13750);
or U18456 (N_18456,N_12864,N_15519);
and U18457 (N_18457,N_14534,N_15364);
nand U18458 (N_18458,N_13293,N_14122);
nand U18459 (N_18459,N_12565,N_13924);
and U18460 (N_18460,N_13372,N_14055);
and U18461 (N_18461,N_15502,N_15574);
nand U18462 (N_18462,N_13221,N_15171);
nor U18463 (N_18463,N_12858,N_12608);
nor U18464 (N_18464,N_14452,N_14120);
and U18465 (N_18465,N_15489,N_13471);
and U18466 (N_18466,N_13057,N_13981);
and U18467 (N_18467,N_14105,N_12853);
xnor U18468 (N_18468,N_14362,N_14817);
xnor U18469 (N_18469,N_14113,N_13030);
nor U18470 (N_18470,N_15523,N_14184);
nor U18471 (N_18471,N_14952,N_15324);
nand U18472 (N_18472,N_13696,N_13911);
nand U18473 (N_18473,N_14937,N_14412);
xor U18474 (N_18474,N_13158,N_14652);
nor U18475 (N_18475,N_14723,N_14875);
nand U18476 (N_18476,N_14316,N_14257);
or U18477 (N_18477,N_12650,N_14854);
or U18478 (N_18478,N_15157,N_13764);
and U18479 (N_18479,N_13160,N_15062);
xnor U18480 (N_18480,N_12890,N_13725);
or U18481 (N_18481,N_14942,N_12721);
and U18482 (N_18482,N_14803,N_14327);
xor U18483 (N_18483,N_14722,N_14667);
nor U18484 (N_18484,N_14901,N_14686);
nor U18485 (N_18485,N_14932,N_14128);
or U18486 (N_18486,N_13887,N_14709);
nor U18487 (N_18487,N_15439,N_14347);
or U18488 (N_18488,N_12597,N_13260);
and U18489 (N_18489,N_15566,N_14220);
and U18490 (N_18490,N_12863,N_15110);
and U18491 (N_18491,N_14606,N_15572);
or U18492 (N_18492,N_13393,N_13686);
nand U18493 (N_18493,N_14273,N_14091);
and U18494 (N_18494,N_15466,N_13876);
nand U18495 (N_18495,N_12759,N_15160);
or U18496 (N_18496,N_13829,N_14137);
nand U18497 (N_18497,N_14272,N_14648);
nor U18498 (N_18498,N_14569,N_12600);
nand U18499 (N_18499,N_14442,N_14616);
and U18500 (N_18500,N_13422,N_13633);
or U18501 (N_18501,N_13433,N_14161);
or U18502 (N_18502,N_13578,N_14655);
and U18503 (N_18503,N_14227,N_12911);
nor U18504 (N_18504,N_15172,N_14953);
or U18505 (N_18505,N_14127,N_15262);
nand U18506 (N_18506,N_13880,N_15340);
xor U18507 (N_18507,N_13093,N_13289);
nand U18508 (N_18508,N_15204,N_14167);
nor U18509 (N_18509,N_14557,N_13678);
and U18510 (N_18510,N_15523,N_13444);
or U18511 (N_18511,N_13671,N_15060);
nor U18512 (N_18512,N_14544,N_15084);
xnor U18513 (N_18513,N_14522,N_14850);
and U18514 (N_18514,N_13478,N_13970);
nor U18515 (N_18515,N_13598,N_14215);
and U18516 (N_18516,N_15085,N_13073);
or U18517 (N_18517,N_13274,N_13382);
nand U18518 (N_18518,N_15002,N_14933);
nand U18519 (N_18519,N_14854,N_12504);
nor U18520 (N_18520,N_14970,N_14118);
xnor U18521 (N_18521,N_15147,N_14733);
xnor U18522 (N_18522,N_14208,N_15200);
xor U18523 (N_18523,N_14831,N_15150);
xor U18524 (N_18524,N_14633,N_12903);
or U18525 (N_18525,N_12788,N_13897);
or U18526 (N_18526,N_13549,N_12833);
or U18527 (N_18527,N_12695,N_13600);
nor U18528 (N_18528,N_12565,N_14971);
nand U18529 (N_18529,N_13387,N_15058);
nand U18530 (N_18530,N_14393,N_14232);
xnor U18531 (N_18531,N_13092,N_13689);
nor U18532 (N_18532,N_13767,N_14116);
nor U18533 (N_18533,N_13729,N_12551);
or U18534 (N_18534,N_15011,N_13165);
or U18535 (N_18535,N_13246,N_13801);
or U18536 (N_18536,N_12524,N_15315);
nand U18537 (N_18537,N_14020,N_13145);
nor U18538 (N_18538,N_13845,N_15605);
nand U18539 (N_18539,N_15282,N_13189);
xnor U18540 (N_18540,N_13868,N_15382);
nor U18541 (N_18541,N_13515,N_15492);
nand U18542 (N_18542,N_15100,N_13507);
xor U18543 (N_18543,N_13605,N_12576);
and U18544 (N_18544,N_12939,N_13575);
xnor U18545 (N_18545,N_14721,N_14949);
xnor U18546 (N_18546,N_14702,N_12971);
nor U18547 (N_18547,N_13234,N_14354);
and U18548 (N_18548,N_15206,N_15229);
nor U18549 (N_18549,N_13869,N_15144);
and U18550 (N_18550,N_13370,N_13242);
and U18551 (N_18551,N_14686,N_13073);
or U18552 (N_18552,N_15355,N_13539);
nor U18553 (N_18553,N_12904,N_14022);
nor U18554 (N_18554,N_13118,N_13572);
xor U18555 (N_18555,N_12974,N_12817);
and U18556 (N_18556,N_12934,N_14027);
and U18557 (N_18557,N_15048,N_13976);
and U18558 (N_18558,N_14002,N_12811);
nand U18559 (N_18559,N_14996,N_15054);
and U18560 (N_18560,N_13552,N_13446);
or U18561 (N_18561,N_13106,N_14114);
or U18562 (N_18562,N_15297,N_12539);
nor U18563 (N_18563,N_13563,N_15485);
or U18564 (N_18564,N_14923,N_14755);
xor U18565 (N_18565,N_15483,N_14392);
and U18566 (N_18566,N_13761,N_12640);
nand U18567 (N_18567,N_13967,N_13171);
and U18568 (N_18568,N_14370,N_13734);
nor U18569 (N_18569,N_12602,N_13524);
or U18570 (N_18570,N_12973,N_12525);
or U18571 (N_18571,N_13386,N_13896);
or U18572 (N_18572,N_12616,N_14351);
nor U18573 (N_18573,N_13795,N_12642);
or U18574 (N_18574,N_12857,N_13328);
nand U18575 (N_18575,N_13144,N_14238);
and U18576 (N_18576,N_13421,N_14456);
or U18577 (N_18577,N_13022,N_13570);
nand U18578 (N_18578,N_13623,N_13664);
nand U18579 (N_18579,N_12857,N_12807);
xor U18580 (N_18580,N_15415,N_14612);
xor U18581 (N_18581,N_12890,N_15589);
nor U18582 (N_18582,N_14196,N_14587);
xor U18583 (N_18583,N_14100,N_13736);
nand U18584 (N_18584,N_14579,N_15513);
xnor U18585 (N_18585,N_13666,N_15034);
and U18586 (N_18586,N_14525,N_13599);
nor U18587 (N_18587,N_13923,N_13038);
xnor U18588 (N_18588,N_14693,N_14337);
nand U18589 (N_18589,N_13258,N_14034);
or U18590 (N_18590,N_14621,N_13899);
and U18591 (N_18591,N_14928,N_12529);
and U18592 (N_18592,N_12621,N_13411);
and U18593 (N_18593,N_13698,N_15348);
and U18594 (N_18594,N_15213,N_13368);
or U18595 (N_18595,N_13037,N_13740);
and U18596 (N_18596,N_13666,N_15442);
and U18597 (N_18597,N_13560,N_12874);
nand U18598 (N_18598,N_14554,N_13169);
and U18599 (N_18599,N_14438,N_14464);
nand U18600 (N_18600,N_15499,N_14427);
xor U18601 (N_18601,N_14120,N_13439);
nor U18602 (N_18602,N_13289,N_13142);
xnor U18603 (N_18603,N_14890,N_13270);
nor U18604 (N_18604,N_13149,N_15390);
xnor U18605 (N_18605,N_14684,N_13209);
or U18606 (N_18606,N_15204,N_14266);
or U18607 (N_18607,N_15621,N_13354);
nand U18608 (N_18608,N_12631,N_14934);
or U18609 (N_18609,N_15507,N_13641);
xnor U18610 (N_18610,N_14276,N_12548);
nand U18611 (N_18611,N_14655,N_13532);
or U18612 (N_18612,N_13362,N_12960);
nor U18613 (N_18613,N_13033,N_15151);
or U18614 (N_18614,N_14892,N_13140);
nand U18615 (N_18615,N_15557,N_13653);
nand U18616 (N_18616,N_13371,N_14702);
and U18617 (N_18617,N_14330,N_12610);
nand U18618 (N_18618,N_14120,N_13051);
xnor U18619 (N_18619,N_13794,N_13526);
and U18620 (N_18620,N_13235,N_15198);
or U18621 (N_18621,N_13978,N_14836);
and U18622 (N_18622,N_13924,N_14039);
nor U18623 (N_18623,N_14990,N_12559);
nand U18624 (N_18624,N_13608,N_13688);
xnor U18625 (N_18625,N_12731,N_13051);
nand U18626 (N_18626,N_14549,N_14816);
xor U18627 (N_18627,N_14223,N_15523);
or U18628 (N_18628,N_14155,N_12740);
nor U18629 (N_18629,N_14830,N_15290);
xor U18630 (N_18630,N_14775,N_14585);
or U18631 (N_18631,N_15529,N_14149);
xnor U18632 (N_18632,N_13672,N_13737);
nand U18633 (N_18633,N_14175,N_15003);
and U18634 (N_18634,N_14287,N_14929);
nor U18635 (N_18635,N_12578,N_12720);
xnor U18636 (N_18636,N_15234,N_14281);
and U18637 (N_18637,N_14537,N_15251);
xor U18638 (N_18638,N_13993,N_15223);
and U18639 (N_18639,N_15450,N_13838);
nand U18640 (N_18640,N_12694,N_15559);
nand U18641 (N_18641,N_13933,N_14660);
nand U18642 (N_18642,N_13241,N_12947);
and U18643 (N_18643,N_13970,N_15575);
nor U18644 (N_18644,N_13117,N_14474);
or U18645 (N_18645,N_13520,N_14388);
or U18646 (N_18646,N_13127,N_15022);
and U18647 (N_18647,N_15053,N_13381);
and U18648 (N_18648,N_13532,N_13216);
nor U18649 (N_18649,N_14179,N_15323);
nand U18650 (N_18650,N_12971,N_12779);
nor U18651 (N_18651,N_14064,N_12887);
and U18652 (N_18652,N_13114,N_14458);
or U18653 (N_18653,N_13616,N_12946);
xnor U18654 (N_18654,N_13575,N_13045);
nor U18655 (N_18655,N_12605,N_13047);
or U18656 (N_18656,N_13437,N_12851);
nand U18657 (N_18657,N_13235,N_13217);
nor U18658 (N_18658,N_14770,N_13103);
nand U18659 (N_18659,N_14223,N_12969);
nand U18660 (N_18660,N_12946,N_13574);
nor U18661 (N_18661,N_14129,N_13505);
nand U18662 (N_18662,N_13546,N_14622);
nor U18663 (N_18663,N_14950,N_15437);
nand U18664 (N_18664,N_13106,N_12954);
nor U18665 (N_18665,N_13993,N_12729);
nand U18666 (N_18666,N_12759,N_14621);
or U18667 (N_18667,N_12897,N_12772);
nand U18668 (N_18668,N_13476,N_12572);
xnor U18669 (N_18669,N_12552,N_13505);
xor U18670 (N_18670,N_13489,N_15270);
nor U18671 (N_18671,N_14185,N_14247);
and U18672 (N_18672,N_15372,N_15566);
or U18673 (N_18673,N_15441,N_13780);
nand U18674 (N_18674,N_14313,N_14471);
xnor U18675 (N_18675,N_12835,N_12710);
or U18676 (N_18676,N_12522,N_13566);
or U18677 (N_18677,N_12706,N_15338);
nor U18678 (N_18678,N_13457,N_14123);
and U18679 (N_18679,N_13658,N_12835);
nor U18680 (N_18680,N_15604,N_13495);
nand U18681 (N_18681,N_14689,N_14596);
xnor U18682 (N_18682,N_13781,N_14433);
nand U18683 (N_18683,N_14414,N_15275);
xor U18684 (N_18684,N_14410,N_15495);
or U18685 (N_18685,N_13977,N_13231);
nand U18686 (N_18686,N_14456,N_14842);
nor U18687 (N_18687,N_13907,N_15624);
and U18688 (N_18688,N_13292,N_13778);
or U18689 (N_18689,N_15309,N_15622);
xnor U18690 (N_18690,N_14482,N_13855);
xnor U18691 (N_18691,N_12732,N_14243);
nor U18692 (N_18692,N_13556,N_13879);
nor U18693 (N_18693,N_13438,N_13119);
xor U18694 (N_18694,N_12672,N_12863);
or U18695 (N_18695,N_13388,N_14254);
xor U18696 (N_18696,N_12955,N_13213);
nor U18697 (N_18697,N_12897,N_14287);
nor U18698 (N_18698,N_13272,N_12788);
or U18699 (N_18699,N_13221,N_13667);
nor U18700 (N_18700,N_14312,N_12592);
or U18701 (N_18701,N_15254,N_13743);
xor U18702 (N_18702,N_13519,N_13867);
xnor U18703 (N_18703,N_13662,N_13041);
and U18704 (N_18704,N_13044,N_14787);
nand U18705 (N_18705,N_13089,N_12550);
nor U18706 (N_18706,N_14702,N_13229);
or U18707 (N_18707,N_14695,N_13775);
or U18708 (N_18708,N_15511,N_14750);
nor U18709 (N_18709,N_13171,N_14730);
nor U18710 (N_18710,N_15024,N_14294);
and U18711 (N_18711,N_15568,N_14895);
or U18712 (N_18712,N_14422,N_13496);
nor U18713 (N_18713,N_15015,N_15514);
nand U18714 (N_18714,N_13296,N_14594);
and U18715 (N_18715,N_13202,N_15497);
and U18716 (N_18716,N_14916,N_13564);
or U18717 (N_18717,N_14822,N_13939);
nand U18718 (N_18718,N_15107,N_13776);
or U18719 (N_18719,N_14790,N_14037);
and U18720 (N_18720,N_13375,N_13156);
and U18721 (N_18721,N_13400,N_13390);
nor U18722 (N_18722,N_15057,N_15299);
nor U18723 (N_18723,N_14987,N_15159);
nand U18724 (N_18724,N_13738,N_12740);
and U18725 (N_18725,N_14636,N_13437);
and U18726 (N_18726,N_13353,N_13225);
or U18727 (N_18727,N_14303,N_12538);
xnor U18728 (N_18728,N_14782,N_15557);
nor U18729 (N_18729,N_13014,N_15250);
nor U18730 (N_18730,N_12812,N_14843);
nor U18731 (N_18731,N_12829,N_14453);
nor U18732 (N_18732,N_14709,N_12511);
xnor U18733 (N_18733,N_14852,N_13035);
nor U18734 (N_18734,N_13446,N_13784);
xnor U18735 (N_18735,N_12520,N_13692);
and U18736 (N_18736,N_12855,N_15484);
and U18737 (N_18737,N_13037,N_15541);
and U18738 (N_18738,N_12684,N_13080);
nand U18739 (N_18739,N_15468,N_14438);
nor U18740 (N_18740,N_12877,N_15045);
nand U18741 (N_18741,N_13784,N_14357);
nand U18742 (N_18742,N_13365,N_13611);
xor U18743 (N_18743,N_15296,N_13570);
or U18744 (N_18744,N_12837,N_14904);
or U18745 (N_18745,N_12682,N_14312);
nor U18746 (N_18746,N_13935,N_15277);
xor U18747 (N_18747,N_14629,N_13618);
or U18748 (N_18748,N_14105,N_13619);
nand U18749 (N_18749,N_12992,N_13595);
nor U18750 (N_18750,N_15813,N_16400);
and U18751 (N_18751,N_17165,N_18437);
nand U18752 (N_18752,N_17293,N_15738);
nand U18753 (N_18753,N_15675,N_17312);
nor U18754 (N_18754,N_16410,N_18659);
xor U18755 (N_18755,N_17722,N_17936);
xor U18756 (N_18756,N_15944,N_17693);
xor U18757 (N_18757,N_18190,N_15788);
xnor U18758 (N_18758,N_17100,N_17814);
or U18759 (N_18759,N_16172,N_18554);
or U18760 (N_18760,N_18738,N_16541);
nand U18761 (N_18761,N_15817,N_16710);
or U18762 (N_18762,N_17506,N_17347);
xnor U18763 (N_18763,N_16074,N_16553);
nor U18764 (N_18764,N_15643,N_18090);
nand U18765 (N_18765,N_15692,N_18185);
nor U18766 (N_18766,N_17295,N_16649);
xnor U18767 (N_18767,N_17116,N_15902);
and U18768 (N_18768,N_18639,N_18407);
nand U18769 (N_18769,N_16918,N_18003);
nand U18770 (N_18770,N_15665,N_15967);
nor U18771 (N_18771,N_16264,N_16489);
xor U18772 (N_18772,N_17589,N_18710);
and U18773 (N_18773,N_17039,N_18178);
and U18774 (N_18774,N_16542,N_18174);
nand U18775 (N_18775,N_16164,N_16549);
or U18776 (N_18776,N_18233,N_18573);
or U18777 (N_18777,N_18094,N_16513);
nor U18778 (N_18778,N_17508,N_16680);
or U18779 (N_18779,N_16149,N_17567);
nand U18780 (N_18780,N_18244,N_18087);
nor U18781 (N_18781,N_15983,N_17530);
nor U18782 (N_18782,N_18705,N_18541);
nand U18783 (N_18783,N_16405,N_17690);
nand U18784 (N_18784,N_17282,N_16810);
or U18785 (N_18785,N_18609,N_18347);
nand U18786 (N_18786,N_17573,N_15686);
xnor U18787 (N_18787,N_18108,N_17301);
nand U18788 (N_18788,N_18026,N_16162);
nand U18789 (N_18789,N_16547,N_17665);
and U18790 (N_18790,N_17096,N_16881);
nand U18791 (N_18791,N_16749,N_18579);
nand U18792 (N_18792,N_17972,N_16579);
nor U18793 (N_18793,N_16317,N_17405);
nand U18794 (N_18794,N_17812,N_16033);
nor U18795 (N_18795,N_18259,N_17911);
nand U18796 (N_18796,N_18651,N_18505);
or U18797 (N_18797,N_18392,N_18458);
nand U18798 (N_18798,N_18455,N_16141);
nand U18799 (N_18799,N_18621,N_16893);
or U18800 (N_18800,N_16548,N_15880);
nand U18801 (N_18801,N_17237,N_18613);
xor U18802 (N_18802,N_18631,N_18715);
and U18803 (N_18803,N_17559,N_18535);
xor U18804 (N_18804,N_17526,N_17873);
and U18805 (N_18805,N_16577,N_17473);
nand U18806 (N_18806,N_16560,N_15696);
nor U18807 (N_18807,N_15844,N_16084);
and U18808 (N_18808,N_16118,N_16169);
nand U18809 (N_18809,N_17804,N_17168);
nand U18810 (N_18810,N_17860,N_18476);
and U18811 (N_18811,N_17923,N_15825);
and U18812 (N_18812,N_17871,N_18559);
nor U18813 (N_18813,N_18694,N_16017);
nor U18814 (N_18814,N_15921,N_17501);
nor U18815 (N_18815,N_17497,N_18276);
or U18816 (N_18816,N_18404,N_16021);
and U18817 (N_18817,N_15945,N_15805);
nor U18818 (N_18818,N_16100,N_17599);
and U18819 (N_18819,N_16699,N_17525);
or U18820 (N_18820,N_18585,N_16319);
nor U18821 (N_18821,N_17944,N_15943);
or U18822 (N_18822,N_16497,N_17635);
and U18823 (N_18823,N_17761,N_16004);
nand U18824 (N_18824,N_16965,N_16873);
nor U18825 (N_18825,N_18263,N_16380);
or U18826 (N_18826,N_17798,N_18568);
or U18827 (N_18827,N_18401,N_18221);
and U18828 (N_18828,N_17462,N_17064);
and U18829 (N_18829,N_16154,N_16146);
and U18830 (N_18830,N_16874,N_17715);
or U18831 (N_18831,N_16471,N_17042);
or U18832 (N_18832,N_18046,N_18132);
xor U18833 (N_18833,N_17957,N_17374);
and U18834 (N_18834,N_16960,N_18195);
xor U18835 (N_18835,N_16241,N_17359);
or U18836 (N_18836,N_16569,N_18733);
xor U18837 (N_18837,N_18663,N_17638);
xnor U18838 (N_18838,N_17218,N_15942);
and U18839 (N_18839,N_17037,N_18092);
and U18840 (N_18840,N_15707,N_17515);
and U18841 (N_18841,N_15915,N_16727);
or U18842 (N_18842,N_17421,N_16768);
or U18843 (N_18843,N_16199,N_17117);
or U18844 (N_18844,N_17284,N_16833);
and U18845 (N_18845,N_18084,N_15963);
or U18846 (N_18846,N_15977,N_16103);
nand U18847 (N_18847,N_18691,N_17631);
or U18848 (N_18848,N_17794,N_17514);
xnor U18849 (N_18849,N_17843,N_17894);
xnor U18850 (N_18850,N_17256,N_16813);
and U18851 (N_18851,N_17740,N_15918);
or U18852 (N_18852,N_17674,N_17054);
xnor U18853 (N_18853,N_18469,N_18723);
nor U18854 (N_18854,N_18575,N_17652);
nor U18855 (N_18855,N_16260,N_18745);
and U18856 (N_18856,N_16466,N_18329);
and U18857 (N_18857,N_17443,N_16282);
or U18858 (N_18858,N_18236,N_17148);
xnor U18859 (N_18859,N_17060,N_15973);
xor U18860 (N_18860,N_17420,N_16249);
nor U18861 (N_18861,N_18219,N_16205);
or U18862 (N_18862,N_17705,N_16627);
xor U18863 (N_18863,N_18297,N_16136);
or U18864 (N_18864,N_17830,N_17142);
nand U18865 (N_18865,N_16292,N_17906);
nor U18866 (N_18866,N_17430,N_18557);
nand U18867 (N_18867,N_18207,N_15782);
xnor U18868 (N_18868,N_18686,N_17095);
or U18869 (N_18869,N_18346,N_16895);
nor U18870 (N_18870,N_16878,N_17952);
and U18871 (N_18871,N_16481,N_16412);
or U18872 (N_18872,N_18293,N_16616);
xor U18873 (N_18873,N_18016,N_16907);
nand U18874 (N_18874,N_17363,N_18354);
and U18875 (N_18875,N_15925,N_18169);
or U18876 (N_18876,N_16515,N_17387);
xor U18877 (N_18877,N_18369,N_15689);
nand U18878 (N_18878,N_16558,N_16590);
or U18879 (N_18879,N_18604,N_17130);
or U18880 (N_18880,N_18319,N_17826);
nor U18881 (N_18881,N_17551,N_16611);
nor U18882 (N_18882,N_16739,N_16863);
and U18883 (N_18883,N_16805,N_16433);
nand U18884 (N_18884,N_15989,N_18035);
or U18885 (N_18885,N_15786,N_17545);
nand U18886 (N_18886,N_17220,N_17101);
or U18887 (N_18887,N_16885,N_17482);
nand U18888 (N_18888,N_17580,N_16736);
or U18889 (N_18889,N_17030,N_16682);
nor U18890 (N_18890,N_18038,N_18363);
and U18891 (N_18891,N_15980,N_17783);
or U18892 (N_18892,N_18413,N_16786);
xnor U18893 (N_18893,N_17157,N_17186);
nand U18894 (N_18894,N_17935,N_17194);
nor U18895 (N_18895,N_17166,N_18361);
nor U18896 (N_18896,N_16914,N_18634);
nor U18897 (N_18897,N_17498,N_17544);
xnor U18898 (N_18898,N_15857,N_17388);
nor U18899 (N_18899,N_16479,N_17953);
nand U18900 (N_18900,N_18685,N_16673);
nand U18901 (N_18901,N_18111,N_17024);
xor U18902 (N_18902,N_18146,N_16493);
nor U18903 (N_18903,N_15706,N_18483);
xor U18904 (N_18904,N_16189,N_16543);
nor U18905 (N_18905,N_16254,N_17524);
or U18906 (N_18906,N_16564,N_16028);
xor U18907 (N_18907,N_16753,N_15975);
or U18908 (N_18908,N_16638,N_16315);
nand U18909 (N_18909,N_16185,N_16061);
and U18910 (N_18910,N_15929,N_17605);
and U18911 (N_18911,N_18472,N_18421);
nor U18912 (N_18912,N_15759,N_16959);
nand U18913 (N_18913,N_16617,N_16465);
nor U18914 (N_18914,N_18479,N_18488);
or U18915 (N_18915,N_15896,N_15781);
nand U18916 (N_18916,N_16670,N_18167);
or U18917 (N_18917,N_17931,N_16689);
and U18918 (N_18918,N_15678,N_15911);
nor U18919 (N_18919,N_18569,N_16953);
or U18920 (N_18920,N_18417,N_16843);
xnor U18921 (N_18921,N_17590,N_16218);
or U18922 (N_18922,N_18310,N_16495);
nor U18923 (N_18923,N_15655,N_17307);
nand U18924 (N_18924,N_17193,N_16795);
and U18925 (N_18925,N_16429,N_15843);
or U18926 (N_18926,N_15995,N_17925);
or U18927 (N_18927,N_18571,N_17057);
and U18928 (N_18928,N_16018,N_17639);
nand U18929 (N_18929,N_16411,N_18306);
nor U18930 (N_18930,N_17283,N_16243);
or U18931 (N_18931,N_17769,N_17625);
xnor U18932 (N_18932,N_16123,N_17485);
xnor U18933 (N_18933,N_15819,N_18556);
xnor U18934 (N_18934,N_17822,N_17774);
or U18935 (N_18935,N_15672,N_17341);
xnor U18936 (N_18936,N_18398,N_15820);
and U18937 (N_18937,N_17091,N_15868);
and U18938 (N_18938,N_17464,N_16394);
nor U18939 (N_18939,N_18484,N_16178);
xnor U18940 (N_18940,N_17300,N_16781);
or U18941 (N_18941,N_17771,N_16356);
or U18942 (N_18942,N_18021,N_18203);
and U18943 (N_18943,N_17044,N_17147);
nor U18944 (N_18944,N_17720,N_16402);
and U18945 (N_18945,N_17512,N_15654);
and U18946 (N_18946,N_16663,N_16568);
or U18947 (N_18947,N_17909,N_16993);
and U18948 (N_18948,N_17302,N_17770);
nor U18949 (N_18949,N_16016,N_18352);
or U18950 (N_18950,N_15766,N_18578);
nand U18951 (N_18951,N_16206,N_17303);
xor U18952 (N_18952,N_17452,N_17160);
nor U18953 (N_18953,N_15684,N_16053);
and U18954 (N_18954,N_16083,N_15681);
xnor U18955 (N_18955,N_15808,N_17324);
and U18956 (N_18956,N_17948,N_17615);
and U18957 (N_18957,N_17831,N_17681);
nand U18958 (N_18958,N_17731,N_16963);
nand U18959 (N_18959,N_15970,N_16803);
xnor U18960 (N_18960,N_16764,N_16269);
nand U18961 (N_18961,N_16335,N_17048);
xor U18962 (N_18962,N_18296,N_17242);
nor U18963 (N_18963,N_16476,N_16656);
nand U18964 (N_18964,N_18591,N_18457);
or U18965 (N_18965,N_17466,N_16195);
or U18966 (N_18966,N_16737,N_16514);
xor U18967 (N_18967,N_16439,N_15688);
nand U18968 (N_18968,N_18532,N_18561);
and U18969 (N_18969,N_17745,N_18282);
and U18970 (N_18970,N_15834,N_16355);
or U18971 (N_18971,N_16448,N_18172);
or U18972 (N_18972,N_17431,N_16460);
nand U18973 (N_18973,N_16387,N_18365);
xor U18974 (N_18974,N_15869,N_16068);
or U18975 (N_18975,N_17358,N_17565);
nor U18976 (N_18976,N_18223,N_17691);
or U18977 (N_18977,N_16790,N_15953);
nor U18978 (N_18978,N_17434,N_16823);
or U18979 (N_18979,N_17719,N_18622);
and U18980 (N_18980,N_15905,N_17829);
xor U18981 (N_18981,N_16116,N_16272);
nor U18982 (N_18982,N_16897,N_18136);
and U18983 (N_18983,N_16425,N_15683);
nor U18984 (N_18984,N_16721,N_17992);
nor U18985 (N_18985,N_16209,N_17739);
nand U18986 (N_18986,N_16486,N_16720);
and U18987 (N_18987,N_18510,N_18058);
nor U18988 (N_18988,N_17110,N_18030);
or U18989 (N_18989,N_18529,N_17672);
and U18990 (N_18990,N_18272,N_18381);
nand U18991 (N_18991,N_18372,N_17252);
nand U18992 (N_18992,N_16950,N_16855);
xnor U18993 (N_18993,N_17627,N_15711);
or U18994 (N_18994,N_17213,N_18180);
or U18995 (N_18995,N_18465,N_15709);
and U18996 (N_18996,N_15893,N_15949);
and U18997 (N_18997,N_16392,N_16921);
and U18998 (N_18998,N_17913,N_18312);
and U18999 (N_18999,N_16593,N_15815);
and U19000 (N_19000,N_16107,N_16762);
or U19001 (N_19001,N_16703,N_17248);
nor U19002 (N_19002,N_18615,N_17854);
or U19003 (N_19003,N_16211,N_17081);
nand U19004 (N_19004,N_17476,N_16019);
and U19005 (N_19005,N_18545,N_16139);
or U19006 (N_19006,N_16728,N_16231);
nand U19007 (N_19007,N_18656,N_15889);
xnor U19008 (N_19008,N_15888,N_18491);
or U19009 (N_19009,N_18338,N_16712);
nand U19010 (N_19010,N_17576,N_16113);
or U19011 (N_19011,N_18340,N_16485);
xnor U19012 (N_19012,N_17225,N_15745);
xor U19013 (N_19013,N_16414,N_16785);
nor U19014 (N_19014,N_18506,N_16353);
or U19015 (N_19015,N_17195,N_17063);
or U19016 (N_19016,N_17239,N_17093);
xor U19017 (N_19017,N_17103,N_16247);
nand U19018 (N_19018,N_17296,N_16299);
or U19019 (N_19019,N_18268,N_18082);
or U19020 (N_19020,N_18358,N_17172);
nor U19021 (N_19021,N_16257,N_17177);
nor U19022 (N_19022,N_17072,N_16540);
and U19023 (N_19023,N_15724,N_17883);
or U19024 (N_19024,N_18537,N_16181);
or U19025 (N_19025,N_17052,N_17088);
and U19026 (N_19026,N_18144,N_18524);
and U19027 (N_19027,N_18238,N_15669);
and U19028 (N_19028,N_15884,N_18333);
and U19029 (N_19029,N_16995,N_17268);
nor U19030 (N_19030,N_17958,N_17173);
xor U19031 (N_19031,N_15685,N_18355);
xor U19032 (N_19032,N_16370,N_17566);
nand U19033 (N_19033,N_18580,N_16002);
and U19034 (N_19034,N_18431,N_16659);
or U19035 (N_19035,N_15785,N_15793);
nand U19036 (N_19036,N_16979,N_18447);
and U19037 (N_19037,N_17999,N_18749);
and U19038 (N_19038,N_18139,N_18106);
and U19039 (N_19039,N_16253,N_16098);
nor U19040 (N_19040,N_16738,N_16233);
and U19041 (N_19041,N_16182,N_18245);
nor U19042 (N_19042,N_17281,N_15703);
nand U19043 (N_19043,N_17269,N_18641);
nand U19044 (N_19044,N_17721,N_16403);
nor U19045 (N_19045,N_16436,N_18370);
nand U19046 (N_19046,N_16800,N_17694);
xnor U19047 (N_19047,N_18034,N_15900);
nor U19048 (N_19048,N_17034,N_18643);
xnor U19049 (N_19049,N_17276,N_15926);
or U19050 (N_19050,N_17089,N_18513);
nor U19051 (N_19051,N_17345,N_17973);
or U19052 (N_19052,N_16364,N_17577);
nand U19053 (N_19053,N_18145,N_18316);
or U19054 (N_19054,N_17151,N_16046);
xnor U19055 (N_19055,N_17868,N_17141);
or U19056 (N_19056,N_18104,N_17942);
nand U19057 (N_19057,N_16801,N_16916);
nand U19058 (N_19058,N_18116,N_15798);
xor U19059 (N_19059,N_18043,N_18662);
nand U19060 (N_19060,N_17976,N_17112);
xor U19061 (N_19061,N_16188,N_16134);
or U19062 (N_19062,N_18270,N_17823);
or U19063 (N_19063,N_16071,N_18160);
or U19064 (N_19064,N_17688,N_17092);
or U19065 (N_19065,N_16262,N_17384);
and U19066 (N_19066,N_15679,N_16610);
and U19067 (N_19067,N_15891,N_16420);
nor U19068 (N_19068,N_16445,N_16902);
nand U19069 (N_19069,N_18019,N_16310);
or U19070 (N_19070,N_17575,N_16912);
nand U19071 (N_19071,N_18448,N_16361);
nor U19072 (N_19072,N_17333,N_16418);
and U19073 (N_19073,N_17067,N_17987);
nor U19074 (N_19074,N_16362,N_16242);
nor U19075 (N_19075,N_17964,N_18273);
or U19076 (N_19076,N_15879,N_17755);
xor U19077 (N_19077,N_16975,N_17483);
xnor U19078 (N_19078,N_18383,N_16605);
and U19079 (N_19079,N_18708,N_17344);
nor U19080 (N_19080,N_18191,N_16120);
and U19081 (N_19081,N_15837,N_17912);
nand U19082 (N_19082,N_17777,N_18013);
nor U19083 (N_19083,N_18577,N_18228);
and U19084 (N_19084,N_15705,N_18657);
xor U19085 (N_19085,N_17241,N_16693);
or U19086 (N_19086,N_15850,N_16731);
xor U19087 (N_19087,N_18216,N_15840);
nor U19088 (N_19088,N_17107,N_16093);
nor U19089 (N_19089,N_17586,N_16075);
nand U19090 (N_19090,N_18017,N_16308);
nor U19091 (N_19091,N_15846,N_17529);
nor U19092 (N_19092,N_17983,N_17569);
nor U19093 (N_19093,N_18549,N_18331);
nor U19094 (N_19094,N_16760,N_18307);
xor U19095 (N_19095,N_16911,N_16634);
or U19096 (N_19096,N_15872,N_17538);
nand U19097 (N_19097,N_18667,N_16284);
xnor U19098 (N_19098,N_17175,N_16557);
xor U19099 (N_19099,N_16115,N_16860);
nor U19100 (N_19100,N_16326,N_15882);
nand U19101 (N_19101,N_16092,N_15658);
nand U19102 (N_19102,N_16849,N_17204);
and U19103 (N_19103,N_17841,N_18714);
xor U19104 (N_19104,N_15634,N_18423);
xor U19105 (N_19105,N_16121,N_17588);
nand U19106 (N_19106,N_16857,N_18600);
xor U19107 (N_19107,N_17730,N_17409);
nand U19108 (N_19108,N_17278,N_17206);
or U19109 (N_19109,N_15969,N_16322);
or U19110 (N_19110,N_15919,N_16684);
and U19111 (N_19111,N_18120,N_15797);
and U19112 (N_19112,N_17535,N_16475);
nor U19113 (N_19113,N_15659,N_17929);
nand U19114 (N_19114,N_17402,N_16102);
nand U19115 (N_19115,N_15957,N_17233);
xor U19116 (N_19116,N_18385,N_18635);
and U19117 (N_19117,N_18161,N_17671);
or U19118 (N_19118,N_16551,N_16578);
nor U19119 (N_19119,N_16038,N_18220);
xnor U19120 (N_19120,N_16328,N_17087);
and U19121 (N_19121,N_17439,N_17159);
xnor U19122 (N_19122,N_17955,N_17616);
and U19123 (N_19123,N_16161,N_16831);
nor U19124 (N_19124,N_16759,N_18623);
and U19125 (N_19125,N_17758,N_16904);
nor U19126 (N_19126,N_18747,N_17310);
and U19127 (N_19127,N_16286,N_18496);
nor U19128 (N_19128,N_16691,N_16001);
and U19129 (N_19129,N_15742,N_17306);
nand U19130 (N_19130,N_16382,N_18237);
and U19131 (N_19131,N_15976,N_17271);
nor U19132 (N_19132,N_15767,N_17121);
or U19133 (N_19133,N_17540,N_18428);
nor U19134 (N_19134,N_18462,N_15756);
xnor U19135 (N_19135,N_16629,N_16419);
xor U19136 (N_19136,N_15674,N_17946);
nor U19137 (N_19137,N_16406,N_16915);
and U19138 (N_19138,N_16201,N_18408);
nor U19139 (N_19139,N_15694,N_18485);
nor U19140 (N_19140,N_18375,N_17267);
or U19141 (N_19141,N_17910,N_18239);
nand U19142 (N_19142,N_17863,N_18041);
nand U19143 (N_19143,N_16342,N_16457);
xor U19144 (N_19144,N_15736,N_16794);
nor U19145 (N_19145,N_18425,N_17880);
nand U19146 (N_19146,N_16806,N_17188);
xor U19147 (N_19147,N_17712,N_17375);
xnor U19148 (N_19148,N_16646,N_17872);
or U19149 (N_19149,N_18677,N_18504);
and U19150 (N_19150,N_17005,N_16138);
nor U19151 (N_19151,N_18005,N_17620);
and U19152 (N_19152,N_16072,N_18069);
or U19153 (N_19153,N_18079,N_16056);
nand U19154 (N_19154,N_16451,N_18054);
xor U19155 (N_19155,N_18155,N_17596);
or U19156 (N_19156,N_16086,N_16500);
nand U19157 (N_19157,N_18251,N_16051);
nand U19158 (N_19158,N_16179,N_15752);
or U19159 (N_19159,N_17025,N_18587);
nand U19160 (N_19160,N_15719,N_15871);
or U19161 (N_19161,N_15633,N_17549);
xnor U19162 (N_19162,N_16746,N_16430);
or U19163 (N_19163,N_16844,N_18743);
or U19164 (N_19164,N_18616,N_16517);
and U19165 (N_19165,N_17069,N_16996);
or U19166 (N_19166,N_17299,N_17680);
nor U19167 (N_19167,N_16776,N_17998);
nor U19168 (N_19168,N_16129,N_16652);
nand U19169 (N_19169,N_16359,N_18397);
and U19170 (N_19170,N_16478,N_18748);
xnor U19171 (N_19171,N_16148,N_18117);
nand U19172 (N_19172,N_18304,N_16705);
or U19173 (N_19173,N_15885,N_17416);
and U19174 (N_19174,N_17417,N_18502);
or U19175 (N_19175,N_16741,N_18480);
or U19176 (N_19176,N_18521,N_17008);
or U19177 (N_19177,N_16811,N_15717);
nor U19178 (N_19178,N_18739,N_17624);
and U19179 (N_19179,N_16596,N_18027);
or U19180 (N_19180,N_17918,N_18525);
nor U19181 (N_19181,N_16064,N_18687);
nand U19182 (N_19182,N_18552,N_18164);
xor U19183 (N_19183,N_17372,N_16039);
nand U19184 (N_19184,N_18309,N_18343);
and U19185 (N_19185,N_18512,N_17046);
xnor U19186 (N_19186,N_17898,N_17710);
and U19187 (N_19187,N_16440,N_16345);
or U19188 (N_19188,N_18429,N_18519);
nor U19189 (N_19189,N_16059,N_18689);
xnor U19190 (N_19190,N_18159,N_16240);
xnor U19191 (N_19191,N_18435,N_17723);
nor U19192 (N_19192,N_18308,N_16274);
nand U19193 (N_19193,N_16399,N_18068);
nand U19194 (N_19194,N_18494,N_16055);
nand U19195 (N_19195,N_16839,N_18114);
or U19196 (N_19196,N_18224,N_17356);
and U19197 (N_19197,N_18498,N_18241);
nand U19198 (N_19198,N_15795,N_16556);
nor U19199 (N_19199,N_18332,N_16648);
nand U19200 (N_19200,N_17090,N_17040);
or U19201 (N_19201,N_16255,N_17634);
nand U19202 (N_19202,N_16922,N_17629);
nor U19203 (N_19203,N_16528,N_18563);
nand U19204 (N_19204,N_18590,N_18603);
and U19205 (N_19205,N_17463,N_18493);
xnor U19206 (N_19206,N_18258,N_16330);
and U19207 (N_19207,N_17288,N_18152);
or U19208 (N_19208,N_15930,N_17633);
and U19209 (N_19209,N_18105,N_18154);
or U19210 (N_19210,N_17029,N_17821);
or U19211 (N_19211,N_17904,N_18594);
nor U19212 (N_19212,N_18170,N_16105);
nor U19213 (N_19213,N_18345,N_16283);
xor U19214 (N_19214,N_17180,N_17606);
nand U19215 (N_19215,N_16381,N_16957);
xnor U19216 (N_19216,N_18255,N_16078);
xnor U19217 (N_19217,N_16932,N_17594);
and U19218 (N_19218,N_17015,N_18101);
nand U19219 (N_19219,N_16170,N_16091);
nand U19220 (N_19220,N_16334,N_16119);
and U19221 (N_19221,N_18071,N_17051);
nand U19222 (N_19222,N_16751,N_15833);
nand U19223 (N_19223,N_17686,N_17169);
or U19224 (N_19224,N_17297,N_16314);
nand U19225 (N_19225,N_17663,N_18254);
nor U19226 (N_19226,N_15762,N_18344);
nor U19227 (N_19227,N_17158,N_18729);
xor U19228 (N_19228,N_18211,N_18311);
nand U19229 (N_19229,N_17820,N_17746);
nand U19230 (N_19230,N_16939,N_16802);
and U19231 (N_19231,N_17571,N_18489);
or U19232 (N_19232,N_16943,N_16640);
and U19233 (N_19233,N_15961,N_18162);
and U19234 (N_19234,N_17539,N_18374);
or U19235 (N_19235,N_15959,N_17718);
nor U19236 (N_19236,N_17533,N_17438);
nand U19237 (N_19237,N_17348,N_17410);
nor U19238 (N_19238,N_16415,N_15830);
nand U19239 (N_19239,N_17810,N_16725);
xnor U19240 (N_19240,N_18547,N_17143);
nand U19241 (N_19241,N_17198,N_16155);
xnor U19242 (N_19242,N_18324,N_18225);
and U19243 (N_19243,N_18638,N_18567);
nor U19244 (N_19244,N_15647,N_15722);
nor U19245 (N_19245,N_16413,N_17009);
nand U19246 (N_19246,N_16770,N_17311);
nor U19247 (N_19247,N_17289,N_17689);
or U19248 (N_19248,N_16045,N_16608);
nor U19249 (N_19249,N_16934,N_17668);
nand U19250 (N_19250,N_17486,N_16888);
nor U19251 (N_19251,N_17662,N_16667);
and U19252 (N_19252,N_17853,N_18107);
nand U19253 (N_19253,N_15865,N_17313);
xnor U19254 (N_19254,N_16349,N_16836);
xor U19255 (N_19255,N_16900,N_18460);
nor U19256 (N_19256,N_18436,N_17655);
or U19257 (N_19257,N_18628,N_18039);
nor U19258 (N_19258,N_18446,N_16966);
or U19259 (N_19259,N_15641,N_15861);
or U19260 (N_19260,N_16396,N_16585);
or U19261 (N_19261,N_18672,N_17768);
nand U19262 (N_19262,N_17677,N_17189);
and U19263 (N_19263,N_16550,N_18110);
nand U19264 (N_19264,N_18468,N_16982);
or U19265 (N_19265,N_15881,N_17098);
nor U19266 (N_19266,N_16398,N_18097);
nor U19267 (N_19267,N_16031,N_16085);
nand U19268 (N_19268,N_18349,N_18133);
xor U19269 (N_19269,N_17626,N_18452);
and U19270 (N_19270,N_16069,N_17450);
nand U19271 (N_19271,N_17390,N_16826);
or U19272 (N_19272,N_16899,N_15894);
nor U19273 (N_19273,N_16278,N_17162);
or U19274 (N_19274,N_18416,N_17527);
xor U19275 (N_19275,N_16070,N_16559);
nor U19276 (N_19276,N_17725,N_17587);
or U19277 (N_19277,N_16490,N_18647);
or U19278 (N_19278,N_17484,N_16407);
xor U19279 (N_19279,N_18031,N_16789);
xnor U19280 (N_19280,N_18607,N_15790);
and U19281 (N_19281,N_16344,N_17200);
and U19282 (N_19282,N_17021,N_17389);
nor U19283 (N_19283,N_18696,N_16645);
and U19284 (N_19284,N_17458,N_18362);
and U19285 (N_19285,N_17342,N_17800);
and U19286 (N_19286,N_17340,N_16232);
and U19287 (N_19287,N_18551,N_18222);
nand U19288 (N_19288,N_18119,N_16301);
or U19289 (N_19289,N_16861,N_17703);
or U19290 (N_19290,N_17002,N_17471);
xnor U19291 (N_19291,N_15870,N_18495);
and U19292 (N_19292,N_15860,N_17236);
xnor U19293 (N_19293,N_16223,N_17553);
and U19294 (N_19294,N_16563,N_16225);
xnor U19295 (N_19295,N_15666,N_17479);
nor U19296 (N_19296,N_18684,N_18206);
and U19297 (N_19297,N_18722,N_16467);
xor U19298 (N_19298,N_15739,N_17809);
nor U19299 (N_19299,N_18321,N_18095);
and U19300 (N_19300,N_17139,N_16862);
or U19301 (N_19301,N_17790,N_18189);
and U19302 (N_19302,N_16298,N_17637);
xnor U19303 (N_19303,N_16941,N_15859);
and U19304 (N_19304,N_16988,N_17349);
xnor U19305 (N_19305,N_16048,N_18010);
nor U19306 (N_19306,N_16850,N_17630);
or U19307 (N_19307,N_18023,N_18018);
or U19308 (N_19308,N_17031,N_16245);
xnor U19309 (N_19309,N_17145,N_18266);
nand U19310 (N_19310,N_17032,N_17604);
xnor U19311 (N_19311,N_17924,N_17305);
xnor U19312 (N_19312,N_16300,N_15673);
xnor U19313 (N_19313,N_15948,N_16722);
and U19314 (N_19314,N_17897,N_17207);
nand U19315 (N_19315,N_16780,N_15854);
nor U19316 (N_19316,N_16820,N_15780);
or U19317 (N_19317,N_16393,N_18250);
and U19318 (N_19318,N_18192,N_18313);
and U19319 (N_19319,N_16819,N_17163);
and U19320 (N_19320,N_17510,N_16229);
nor U19321 (N_19321,N_16088,N_16073);
and U19322 (N_19322,N_15715,N_18433);
nand U19323 (N_19323,N_17201,N_17982);
and U19324 (N_19324,N_18492,N_16830);
xor U19325 (N_19325,N_17673,N_16054);
and U19326 (N_19326,N_16026,N_17612);
nand U19327 (N_19327,N_16951,N_18430);
nor U19328 (N_19328,N_15940,N_16384);
nand U19329 (N_19329,N_18654,N_16470);
nor U19330 (N_19330,N_16847,N_16688);
or U19331 (N_19331,N_18536,N_18396);
xnor U19332 (N_19332,N_16156,N_17669);
nand U19333 (N_19333,N_17859,N_18049);
nor U19334 (N_19334,N_16367,N_16665);
nor U19335 (N_19335,N_16213,N_18232);
and U19336 (N_19336,N_16639,N_17554);
nor U19337 (N_19337,N_18546,N_15814);
nand U19338 (N_19338,N_18405,N_16664);
or U19339 (N_19339,N_18720,N_18171);
nor U19340 (N_19340,N_17377,N_16432);
nor U19341 (N_19341,N_18072,N_16327);
xnor U19342 (N_19342,N_18231,N_18281);
nand U19343 (N_19343,N_17058,N_15855);
or U19344 (N_19344,N_17321,N_16887);
nor U19345 (N_19345,N_16586,N_16125);
nand U19346 (N_19346,N_15858,N_15751);
and U19347 (N_19347,N_17751,N_18009);
nor U19348 (N_19348,N_15687,N_18692);
or U19349 (N_19349,N_16952,N_17732);
xor U19350 (N_19350,N_18342,N_17645);
nand U19351 (N_19351,N_16158,N_17971);
or U19352 (N_19352,N_16783,N_15804);
nor U19353 (N_19353,N_16961,N_15892);
or U19354 (N_19354,N_18326,N_17546);
or U19355 (N_19355,N_16463,N_18475);
and U19356 (N_19356,N_17273,N_16130);
nand U19357 (N_19357,N_18045,N_16618);
xnor U19358 (N_19358,N_18412,N_16456);
and U19359 (N_19359,N_16877,N_16769);
or U19360 (N_19360,N_17876,N_18012);
nand U19361 (N_19361,N_17916,N_15628);
and U19362 (N_19362,N_17235,N_18713);
nand U19363 (N_19363,N_15791,N_18390);
and U19364 (N_19364,N_17418,N_17555);
and U19365 (N_19365,N_17350,N_16812);
and U19366 (N_19366,N_16743,N_16408);
nand U19367 (N_19367,N_18707,N_16816);
nand U19368 (N_19368,N_18001,N_15629);
and U19369 (N_19369,N_16369,N_16654);
xor U19370 (N_19370,N_17436,N_15981);
or U19371 (N_19371,N_16437,N_16390);
xnor U19372 (N_19372,N_17702,N_16894);
nand U19373 (N_19373,N_15667,N_18295);
and U19374 (N_19374,N_17865,N_17257);
nor U19375 (N_19375,N_16097,N_17981);
or U19376 (N_19376,N_15996,N_17613);
nor U19377 (N_19377,N_15699,N_16313);
nand U19378 (N_19378,N_17807,N_18098);
nand U19379 (N_19379,N_18063,N_17222);
nor U19380 (N_19380,N_17759,N_15775);
xnor U19381 (N_19381,N_16677,N_18008);
nand U19382 (N_19382,N_16679,N_16305);
nand U19383 (N_19383,N_18439,N_17579);
and U19384 (N_19384,N_17294,N_16938);
or U19385 (N_19385,N_16416,N_15809);
nor U19386 (N_19386,N_16891,N_18240);
nor U19387 (N_19387,N_17563,N_18608);
nor U19388 (N_19388,N_18499,N_15730);
xnor U19389 (N_19389,N_16261,N_18006);
or U19390 (N_19390,N_17989,N_17813);
nor U19391 (N_19391,N_15800,N_17423);
nor U19392 (N_19392,N_15773,N_15744);
xnor U19393 (N_19393,N_16009,N_18061);
or U19394 (N_19394,N_18015,N_16307);
and U19395 (N_19395,N_15652,N_16234);
or U19396 (N_19396,N_18066,N_16793);
nor U19397 (N_19397,N_16999,N_15839);
nand U19398 (N_19398,N_17152,N_16389);
nand U19399 (N_19399,N_16374,N_17914);
nand U19400 (N_19400,N_16835,N_18235);
nand U19401 (N_19401,N_17435,N_16666);
and U19402 (N_19402,N_15890,N_18193);
and U19403 (N_19403,N_17414,N_16527);
xnor U19404 (N_19404,N_17764,N_16455);
and U19405 (N_19405,N_17076,N_17399);
nand U19406 (N_19406,N_17601,N_17011);
and U19407 (N_19407,N_18626,N_16846);
and U19408 (N_19408,N_17393,N_15690);
xnor U19409 (N_19409,N_16000,N_15994);
or U19410 (N_19410,N_16626,N_15928);
nor U19411 (N_19411,N_16754,N_18718);
nor U19412 (N_19412,N_16864,N_17683);
nand U19413 (N_19413,N_17792,N_16525);
xor U19414 (N_19414,N_15645,N_17136);
or U19415 (N_19415,N_16409,N_17199);
or U19416 (N_19416,N_16338,N_18242);
nor U19417 (N_19417,N_15877,N_16520);
and U19418 (N_19418,N_18700,N_18540);
or U19419 (N_19419,N_17017,N_16131);
xor U19420 (N_19420,N_17517,N_18330);
nor U19421 (N_19421,N_18466,N_16395);
nand U19422 (N_19422,N_17857,N_16530);
nand U19423 (N_19423,N_17453,N_16944);
and U19424 (N_19424,N_15939,N_15913);
xnor U19425 (N_19425,N_15741,N_17653);
or U19426 (N_19426,N_17270,N_15851);
xnor U19427 (N_19427,N_18366,N_17891);
nand U19428 (N_19428,N_17650,N_15960);
nand U19429 (N_19429,N_17308,N_16876);
nand U19430 (N_19430,N_16773,N_17899);
xnor U19431 (N_19431,N_15769,N_16291);
or U19432 (N_19432,N_18102,N_17932);
and U19433 (N_19433,N_16295,N_17724);
xor U19434 (N_19434,N_15657,N_17757);
and U19435 (N_19435,N_17700,N_18454);
or U19436 (N_19436,N_17851,N_17124);
and U19437 (N_19437,N_17697,N_15763);
nor U19438 (N_19438,N_18115,N_16336);
xor U19439 (N_19439,N_16312,N_17685);
or U19440 (N_19440,N_15632,N_18688);
or U19441 (N_19441,N_17259,N_15799);
xnor U19442 (N_19442,N_17503,N_18302);
and U19443 (N_19443,N_16477,N_17552);
xor U19444 (N_19444,N_17582,N_18611);
nor U19445 (N_19445,N_17219,N_16469);
nor U19446 (N_19446,N_16329,N_16837);
or U19447 (N_19447,N_17304,N_17361);
and U19448 (N_19448,N_18373,N_18292);
and U19449 (N_19449,N_17767,N_18384);
or U19450 (N_19450,N_17119,N_18198);
or U19451 (N_19451,N_16620,N_18438);
xnor U19452 (N_19452,N_16007,N_16065);
nand U19453 (N_19453,N_16732,N_15796);
nand U19454 (N_19454,N_18217,N_16333);
nand U19455 (N_19455,N_18166,N_16650);
xor U19456 (N_19456,N_18056,N_16983);
xor U19457 (N_19457,N_15824,N_16175);
xnor U19458 (N_19458,N_17028,N_17229);
nor U19459 (N_19459,N_18278,N_16742);
and U19460 (N_19460,N_15876,N_17640);
nor U19461 (N_19461,N_17461,N_17354);
or U19462 (N_19462,N_17698,N_17424);
and U19463 (N_19463,N_18177,N_15901);
and U19464 (N_19464,N_17903,N_16521);
xor U19465 (N_19465,N_17502,N_16267);
and U19466 (N_19466,N_18618,N_15991);
xor U19467 (N_19467,N_15802,N_17205);
and U19468 (N_19468,N_15777,N_17997);
and U19469 (N_19469,N_17542,N_15886);
nand U19470 (N_19470,N_18393,N_18737);
or U19471 (N_19471,N_15863,N_18062);
or U19472 (N_19472,N_17656,N_18218);
nand U19473 (N_19473,N_18674,N_16422);
and U19474 (N_19474,N_17977,N_18267);
or U19475 (N_19475,N_16832,N_17223);
nand U19476 (N_19476,N_16576,N_16948);
xnor U19477 (N_19477,N_17286,N_16987);
and U19478 (N_19478,N_16150,N_17993);
xnor U19479 (N_19479,N_15958,N_16095);
nand U19480 (N_19480,N_16371,N_16582);
and U19481 (N_19481,N_16279,N_17889);
nor U19482 (N_19482,N_18305,N_18645);
xnor U19483 (N_19483,N_17202,N_15662);
xor U19484 (N_19484,N_17970,N_17791);
nand U19485 (N_19485,N_18695,N_16079);
and U19486 (N_19486,N_16972,N_17844);
xnor U19487 (N_19487,N_18036,N_15646);
nand U19488 (N_19488,N_16076,N_17848);
xor U19489 (N_19489,N_18325,N_15932);
and U19490 (N_19490,N_16708,N_18142);
xor U19491 (N_19491,N_16535,N_17934);
nand U19492 (N_19492,N_16706,N_16510);
or U19493 (N_19493,N_15899,N_18130);
nor U19494 (N_19494,N_17109,N_17138);
nor U19495 (N_19495,N_18188,N_15768);
nor U19496 (N_19496,N_18424,N_15821);
and U19497 (N_19497,N_17741,N_16502);
and U19498 (N_19498,N_15664,N_16447);
and U19499 (N_19499,N_17317,N_15704);
and U19500 (N_19500,N_16554,N_18746);
nand U19501 (N_19501,N_17351,N_18353);
xor U19502 (N_19502,N_17684,N_16464);
nor U19503 (N_19503,N_17398,N_16931);
or U19504 (N_19504,N_18050,N_15826);
and U19505 (N_19505,N_17658,N_16967);
or U19506 (N_19506,N_16435,N_17480);
and U19507 (N_19507,N_17750,N_16929);
nand U19508 (N_19508,N_18121,N_16946);
nor U19509 (N_19509,N_18507,N_18173);
nand U19510 (N_19510,N_15754,N_17245);
nor U19511 (N_19511,N_17756,N_18359);
or U19512 (N_19512,N_16251,N_18261);
xnor U19513 (N_19513,N_18735,N_18123);
and U19514 (N_19514,N_15812,N_17752);
nand U19515 (N_19515,N_17263,N_16144);
or U19516 (N_19516,N_18025,N_15728);
or U19517 (N_19517,N_16718,N_18299);
and U19518 (N_19518,N_15986,N_16174);
or U19519 (N_19519,N_18456,N_18697);
or U19520 (N_19520,N_15716,N_16397);
xor U19521 (N_19521,N_16145,N_17460);
nand U19522 (N_19522,N_16632,N_16133);
and U19523 (N_19523,N_17679,N_18088);
nand U19524 (N_19524,N_17135,N_18197);
nand U19525 (N_19525,N_18514,N_17187);
and U19526 (N_19526,N_17734,N_17364);
or U19527 (N_19527,N_17670,N_17266);
xor U19528 (N_19528,N_18350,N_17727);
or U19529 (N_19529,N_17651,N_16207);
nor U19530 (N_19530,N_17699,N_17919);
xor U19531 (N_19531,N_16454,N_16200);
and U19532 (N_19532,N_16219,N_15908);
nor U19533 (N_19533,N_16020,N_17447);
nor U19534 (N_19534,N_18427,N_16602);
and U19535 (N_19535,N_17659,N_17446);
nand U19536 (N_19536,N_17144,N_18655);
nor U19537 (N_19537,N_16373,N_17832);
and U19538 (N_19538,N_18553,N_16662);
or U19539 (N_19539,N_16964,N_15907);
xor U19540 (N_19540,N_16230,N_15648);
xnor U19541 (N_19541,N_16488,N_18356);
xor U19542 (N_19542,N_15822,N_16003);
nor U19543 (N_19543,N_18002,N_16239);
nor U19544 (N_19544,N_18007,N_18287);
or U19545 (N_19545,N_16224,N_18523);
nor U19546 (N_19546,N_16194,N_17940);
nor U19547 (N_19547,N_17966,N_18403);
or U19548 (N_19548,N_16082,N_17558);
or U19549 (N_19549,N_17819,N_18165);
xor U19550 (N_19550,N_17570,N_17041);
xor U19551 (N_19551,N_17901,N_17711);
and U19552 (N_19552,N_16782,N_18052);
nor U19553 (N_19553,N_16426,N_16719);
or U19554 (N_19554,N_15779,N_16594);
nor U19555 (N_19555,N_18637,N_16378);
nand U19556 (N_19556,N_17984,N_16655);
and U19557 (N_19557,N_18555,N_17607);
or U19558 (N_19558,N_18434,N_17956);
and U19559 (N_19559,N_16949,N_17619);
or U19560 (N_19560,N_18464,N_17019);
xor U19561 (N_19561,N_18522,N_17915);
xor U19562 (N_19562,N_16544,N_16702);
xor U19563 (N_19563,N_15727,N_16077);
or U19564 (N_19564,N_18364,N_17026);
and U19565 (N_19565,N_17118,N_16289);
nand U19566 (N_19566,N_15829,N_17850);
xor U19567 (N_19567,N_17413,N_16717);
xor U19568 (N_19568,N_16767,N_15626);
nand U19569 (N_19569,N_17185,N_18627);
and U19570 (N_19570,N_18400,N_16112);
or U19571 (N_19571,N_16624,N_16675);
nor U19572 (N_19572,N_17675,N_16986);
or U19573 (N_19573,N_17793,N_17660);
and U19574 (N_19574,N_17006,N_17621);
nor U19575 (N_19575,N_18204,N_18158);
xor U19576 (N_19576,N_16962,N_18683);
and U19577 (N_19577,N_18560,N_18679);
or U19578 (N_19578,N_18652,N_16755);
or U19579 (N_19579,N_16235,N_17747);
xnor U19580 (N_19580,N_18426,N_16365);
and U19581 (N_19581,N_18336,N_17521);
and U19582 (N_19582,N_18011,N_17326);
nand U19583 (N_19583,N_16094,N_16332);
xor U19584 (N_19584,N_15650,N_16192);
xor U19585 (N_19585,N_17818,N_16700);
nor U19586 (N_19586,N_18044,N_18128);
nor U19587 (N_19587,N_17403,N_17392);
or U19588 (N_19588,N_18264,N_16715);
xor U19589 (N_19589,N_17368,N_17706);
and U19590 (N_19590,N_18124,N_17714);
or U19591 (N_19591,N_17370,N_17816);
and U19592 (N_19592,N_17386,N_18382);
nand U19593 (N_19593,N_17789,N_17995);
xor U19594 (N_19594,N_17362,N_17961);
xor U19595 (N_19595,N_17828,N_16750);
nand U19596 (N_19596,N_16592,N_18704);
nand U19597 (N_19597,N_17742,N_15842);
xnor U19598 (N_19598,N_17507,N_16265);
nor U19599 (N_19599,N_18624,N_16580);
xor U19600 (N_19600,N_15627,N_16815);
nand U19601 (N_19601,N_17128,N_16117);
nand U19602 (N_19602,N_18371,N_16049);
or U19603 (N_19603,N_17261,N_16884);
or U19604 (N_19604,N_15636,N_18143);
or U19605 (N_19605,N_16066,N_17766);
and U19606 (N_19606,N_16190,N_17164);
or U19607 (N_19607,N_15644,N_16023);
xnor U19608 (N_19608,N_17753,N_15923);
xor U19609 (N_19609,N_17622,N_16660);
and U19610 (N_19610,N_16210,N_18736);
or U19611 (N_19611,N_18409,N_16184);
or U19612 (N_19612,N_18134,N_18368);
and U19613 (N_19613,N_18574,N_17773);
nand U19614 (N_19614,N_17077,N_17885);
nand U19615 (N_19615,N_17441,N_16062);
nor U19616 (N_19616,N_15818,N_18029);
nand U19617 (N_19617,N_16137,N_18077);
nand U19618 (N_19618,N_16871,N_17817);
nor U19619 (N_19619,N_17845,N_17490);
nor U19620 (N_19620,N_18257,N_18558);
nor U19621 (N_19621,N_18320,N_16503);
xnor U19622 (N_19622,N_17465,N_17240);
xnor U19623 (N_19623,N_15649,N_15954);
nor U19624 (N_19624,N_17837,N_16865);
or U19625 (N_19625,N_17114,N_17082);
nand U19626 (N_19626,N_17133,N_15897);
xor U19627 (N_19627,N_15631,N_16607);
xor U19628 (N_19628,N_15990,N_16124);
or U19629 (N_19629,N_17943,N_16954);
nor U19630 (N_19630,N_17230,N_16880);
nand U19631 (N_19631,N_16797,N_18149);
nand U19632 (N_19632,N_17523,N_18387);
and U19633 (N_19633,N_15867,N_16507);
and U19634 (N_19634,N_18246,N_17557);
nand U19635 (N_19635,N_18660,N_15952);
or U19636 (N_19636,N_16920,N_18402);
nand U19637 (N_19637,N_18042,N_17890);
or U19638 (N_19638,N_16404,N_18070);
xnor U19639 (N_19639,N_16343,N_18277);
nor U19640 (N_19640,N_16766,N_16603);
and U19641 (N_19641,N_17428,N_15758);
and U19642 (N_19642,N_16573,N_17537);
or U19643 (N_19643,N_16216,N_17228);
xnor U19644 (N_19644,N_17332,N_17796);
xor U19645 (N_19645,N_16446,N_16609);
nand U19646 (N_19646,N_17949,N_17801);
nand U19647 (N_19647,N_17716,N_18583);
and U19648 (N_19648,N_16694,N_18544);
nor U19649 (N_19649,N_16879,N_16994);
nand U19650 (N_19650,N_16350,N_16372);
xor U19651 (N_19651,N_18665,N_18612);
nand U19652 (N_19652,N_17227,N_16883);
nor U19653 (N_19653,N_17055,N_17426);
nor U19654 (N_19654,N_17648,N_17073);
nand U19655 (N_19655,N_17422,N_15845);
and U19656 (N_19656,N_16591,N_16143);
or U19657 (N_19657,N_17105,N_17255);
xor U19658 (N_19658,N_16034,N_17968);
xor U19659 (N_19659,N_17996,N_18265);
xnor U19660 (N_19660,N_15732,N_16752);
nor U19661 (N_19661,N_18528,N_16196);
or U19662 (N_19662,N_18678,N_18210);
and U19663 (N_19663,N_18140,N_17954);
and U19664 (N_19664,N_15637,N_17728);
and U19665 (N_19665,N_18706,N_16010);
or U19666 (N_19666,N_16152,N_18247);
and U19667 (N_19667,N_17004,N_15691);
xor U19668 (N_19668,N_16930,N_16533);
and U19669 (N_19669,N_16221,N_16352);
nand U19670 (N_19670,N_17331,N_18085);
xor U19671 (N_19671,N_17469,N_16587);
nor U19672 (N_19672,N_17713,N_18125);
or U19673 (N_19673,N_16159,N_18477);
nor U19674 (N_19674,N_16992,N_16980);
nand U19675 (N_19675,N_18716,N_16052);
xnor U19676 (N_19676,N_18461,N_18734);
nand U19677 (N_19677,N_15660,N_17595);
nand U19678 (N_19678,N_17395,N_18644);
and U19679 (N_19679,N_16379,N_16537);
or U19680 (N_19680,N_17491,N_16208);
nor U19681 (N_19681,N_18213,N_17419);
or U19682 (N_19682,N_18151,N_17824);
or U19683 (N_19683,N_17085,N_15852);
nor U19684 (N_19684,N_17882,N_18445);
or U19685 (N_19685,N_17990,N_16180);
nand U19686 (N_19686,N_15898,N_17707);
nor U19687 (N_19687,N_15962,N_16157);
xor U19688 (N_19688,N_16368,N_16275);
or U19689 (N_19689,N_18596,N_16698);
nor U19690 (N_19690,N_17786,N_17183);
and U19691 (N_19691,N_17318,N_16671);
and U19692 (N_19692,N_15874,N_18059);
or U19693 (N_19693,N_16252,N_16505);
nor U19694 (N_19694,N_16892,N_18262);
xor U19695 (N_19695,N_17215,N_18253);
or U19696 (N_19696,N_17646,N_18543);
nor U19697 (N_19697,N_18208,N_15979);
and U19698 (N_19698,N_17592,N_17456);
and U19699 (N_19699,N_17687,N_18184);
xor U19700 (N_19700,N_15816,N_16281);
nor U19701 (N_19701,N_18542,N_17444);
or U19702 (N_19702,N_18020,N_15941);
and U19703 (N_19703,N_16104,N_17528);
xor U19704 (N_19704,N_17743,N_15671);
nor U19705 (N_19705,N_17760,N_17591);
nor U19706 (N_19706,N_15701,N_15640);
and U19707 (N_19707,N_16701,N_16761);
xor U19708 (N_19708,N_16108,N_18175);
xor U19709 (N_19709,N_16526,N_18335);
and U19710 (N_19710,N_17695,N_16106);
and U19711 (N_19711,N_17736,N_16516);
and U19712 (N_19712,N_18509,N_16268);
or U19713 (N_19713,N_16127,N_17161);
nand U19714 (N_19714,N_17534,N_18187);
or U19715 (N_19715,N_17666,N_17560);
xor U19716 (N_19716,N_18318,N_16323);
nand U19717 (N_19717,N_16942,N_17099);
nor U19718 (N_19718,N_15801,N_18399);
xnor U19719 (N_19719,N_18701,N_15936);
and U19720 (N_19720,N_17881,N_18562);
or U19721 (N_19721,N_16937,N_16653);
and U19722 (N_19722,N_16177,N_15789);
nor U19723 (N_19723,N_16401,N_16779);
and U19724 (N_19724,N_17251,N_17967);
nand U19725 (N_19725,N_18004,N_15924);
xor U19726 (N_19726,N_16276,N_17181);
xnor U19727 (N_19727,N_18157,N_15726);
and U19728 (N_19728,N_16856,N_16827);
or U19729 (N_19729,N_16866,N_17945);
xnor U19730 (N_19730,N_15783,N_17578);
nor U19731 (N_19731,N_16523,N_16758);
xor U19732 (N_19732,N_18410,N_18520);
or U19733 (N_19733,N_18096,N_17867);
nor U19734 (N_19734,N_17781,N_17170);
nand U19735 (N_19735,N_18163,N_15933);
or U19736 (N_19736,N_17649,N_15625);
or U19737 (N_19737,N_16747,N_18482);
xnor U19738 (N_19738,N_17196,N_16765);
xnor U19739 (N_19739,N_16822,N_16037);
nand U19740 (N_19740,N_17709,N_16204);
xnor U19741 (N_19741,N_16644,N_15832);
and U19742 (N_19742,N_18640,N_15748);
or U19743 (N_19743,N_17314,N_18279);
nor U19744 (N_19744,N_17678,N_17806);
or U19745 (N_19745,N_16035,N_17023);
nand U19746 (N_19746,N_15713,N_16792);
xnor U19747 (N_19747,N_16459,N_18109);
and U19748 (N_19748,N_18086,N_17126);
xnor U19749 (N_19749,N_16567,N_18065);
nor U19750 (N_19750,N_18515,N_18595);
xnor U19751 (N_19751,N_15753,N_18081);
nor U19752 (N_19752,N_16923,N_15746);
nand U19753 (N_19753,N_18315,N_17799);
xor U19754 (N_19754,N_17962,N_15931);
or U19755 (N_19755,N_17352,N_16834);
nor U19756 (N_19756,N_17585,N_18284);
or U19757 (N_19757,N_16615,N_18614);
and U19758 (N_19758,N_16976,N_17505);
nor U19759 (N_19759,N_18470,N_16637);
nor U19760 (N_19760,N_16989,N_17287);
nand U19761 (N_19761,N_17855,N_16633);
or U19762 (N_19762,N_17084,N_17738);
nor U19763 (N_19763,N_18099,N_17325);
xor U19764 (N_19764,N_17437,N_15841);
nand U19765 (N_19765,N_17224,N_15964);
nor U19766 (N_19766,N_15828,N_17536);
and U19767 (N_19767,N_17154,N_17140);
nand U19768 (N_19768,N_15831,N_18712);
nand U19769 (N_19769,N_15974,N_17038);
or U19770 (N_19770,N_15639,N_17000);
and U19771 (N_19771,N_18256,N_16925);
xor U19772 (N_19772,N_17737,N_17415);
and U19773 (N_19773,N_18548,N_18053);
or U19774 (N_19774,N_17744,N_17775);
xor U19775 (N_19775,N_15787,N_17938);
or U19776 (N_19776,N_18646,N_18550);
or U19777 (N_19777,N_16340,N_18620);
and U19778 (N_19778,N_18032,N_16140);
nand U19779 (N_19779,N_17550,N_16220);
and U19780 (N_19780,N_18078,N_18539);
and U19781 (N_19781,N_16566,N_15848);
and U19782 (N_19782,N_16025,N_18724);
nor U19783 (N_19783,N_18339,N_16524);
xor U19784 (N_19784,N_16777,N_15873);
nor U19785 (N_19785,N_15772,N_18422);
nor U19786 (N_19786,N_16013,N_16461);
or U19787 (N_19787,N_16599,N_18449);
and U19788 (N_19788,N_18290,N_17211);
xnor U19789 (N_19789,N_16625,N_16101);
nor U19790 (N_19790,N_16022,N_17879);
nand U19791 (N_19791,N_17643,N_18083);
nor U19792 (N_19792,N_17869,N_18658);
nand U19793 (N_19793,N_17068,N_18376);
nor U19794 (N_19794,N_15700,N_16748);
xnor U19795 (N_19795,N_16858,N_15866);
and U19796 (N_19796,N_18378,N_18075);
and U19797 (N_19797,N_17329,N_15776);
nor U19798 (N_19798,N_16614,N_17323);
nand U19799 (N_19799,N_16581,N_15914);
nor U19800 (N_19800,N_16772,N_18274);
or U19801 (N_19801,N_17214,N_18565);
nand U19802 (N_19802,N_18661,N_17380);
nor U19803 (N_19803,N_17780,N_18726);
and U19804 (N_19804,N_17827,N_18147);
or U19805 (N_19805,N_18711,N_16814);
and U19806 (N_19806,N_18599,N_16595);
xor U19807 (N_19807,N_15653,N_18322);
nor U19808 (N_19808,N_17190,N_15984);
nand U19809 (N_19809,N_17315,N_16099);
xnor U19810 (N_19810,N_17132,N_17197);
xnor U19811 (N_19811,N_15982,N_18415);
nor U19812 (N_19812,N_17547,N_17600);
and U19813 (N_19813,N_16331,N_16977);
xor U19814 (N_19814,N_16388,N_18234);
nor U19815 (N_19815,N_18642,N_16882);
and U19816 (N_19816,N_15955,N_18597);
or U19817 (N_19817,N_17895,N_17597);
xnor U19818 (N_19818,N_15680,N_17926);
or U19819 (N_19819,N_16956,N_17264);
xor U19820 (N_19820,N_17383,N_17013);
or U19821 (N_19821,N_16044,N_18406);
or U19822 (N_19822,N_16259,N_16324);
and U19823 (N_19823,N_18538,N_17115);
nor U19824 (N_19824,N_16187,N_18709);
nand U19825 (N_19825,N_16658,N_17246);
and U19826 (N_19826,N_15635,N_18269);
or U19827 (N_19827,N_18379,N_17488);
nor U19828 (N_19828,N_15856,N_17762);
xor U19829 (N_19829,N_17888,N_15985);
nand U19830 (N_19830,N_18601,N_17614);
or U19831 (N_19831,N_18632,N_18629);
nor U19832 (N_19832,N_16357,N_17155);
or U19833 (N_19833,N_16641,N_16443);
xnor U19834 (N_19834,N_17980,N_15682);
or U19835 (N_19835,N_17249,N_18420);
or U19836 (N_19836,N_16484,N_17852);
xor U19837 (N_19837,N_15778,N_18289);
or U19838 (N_19838,N_16726,N_17896);
and U19839 (N_19839,N_16248,N_16325);
and U19840 (N_19840,N_15972,N_18000);
or U19841 (N_19841,N_17581,N_18300);
and U19842 (N_19842,N_15937,N_16940);
or U19843 (N_19843,N_18014,N_16015);
or U19844 (N_19844,N_17511,N_17951);
xor U19845 (N_19845,N_17861,N_18650);
or U19846 (N_19846,N_18047,N_18617);
nand U19847 (N_19847,N_17062,N_15630);
and U19848 (N_19848,N_17192,N_17338);
xor U19849 (N_19849,N_17027,N_16474);
or U19850 (N_19850,N_17644,N_16280);
nor U19851 (N_19851,N_17884,N_17811);
and U19852 (N_19852,N_18681,N_17319);
xnor U19853 (N_19853,N_15642,N_15917);
nor U19854 (N_19854,N_18486,N_17900);
xor U19855 (N_19855,N_18653,N_17455);
nand U19856 (N_19856,N_18741,N_18463);
xor U19857 (N_19857,N_16775,N_15909);
nor U19858 (N_19858,N_16619,N_16287);
and U19859 (N_19859,N_15875,N_17279);
and U19860 (N_19860,N_15735,N_16511);
and U19861 (N_19861,N_17564,N_18028);
or U19862 (N_19862,N_15749,N_16147);
and U19863 (N_19863,N_18201,N_15950);
or U19864 (N_19864,N_16160,N_18699);
xor U19865 (N_19865,N_16845,N_17014);
nand U19866 (N_19866,N_16868,N_17097);
nand U19867 (N_19867,N_16636,N_16774);
nand U19868 (N_19868,N_17583,N_18394);
nand U19869 (N_19869,N_16428,N_16729);
or U19870 (N_19870,N_18260,N_16024);
nand U19871 (N_19871,N_17922,N_17070);
xor U19872 (N_19872,N_15740,N_16583);
and U19873 (N_19873,N_18500,N_18728);
nand U19874 (N_19874,N_18357,N_16730);
xnor U19875 (N_19875,N_18360,N_18196);
and U19876 (N_19876,N_17369,N_16621);
and U19877 (N_19877,N_16375,N_15920);
xor U19878 (N_19878,N_17184,N_16552);
and U19879 (N_19879,N_18666,N_16690);
and U19880 (N_19880,N_16997,N_18633);
xor U19881 (N_19881,N_16128,N_16238);
nor U19882 (N_19882,N_17043,N_18033);
xnor U19883 (N_19883,N_16354,N_17445);
or U19884 (N_19884,N_16990,N_16909);
xor U19885 (N_19885,N_17086,N_15747);
xnor U19886 (N_19886,N_18527,N_16494);
nor U19887 (N_19887,N_16444,N_15757);
xor U19888 (N_19888,N_15951,N_17226);
and U19889 (N_19889,N_17153,N_17156);
or U19890 (N_19890,N_18100,N_16453);
xor U19891 (N_19891,N_18721,N_16132);
and U19892 (N_19892,N_17532,N_16538);
nor U19893 (N_19893,N_15734,N_16854);
nor U19894 (N_19894,N_16491,N_16531);
nor U19895 (N_19895,N_16063,N_16043);
and U19896 (N_19896,N_17210,N_18473);
nand U19897 (N_19897,N_17078,N_16935);
xnor U19898 (N_19898,N_18586,N_17772);
and U19899 (N_19899,N_17928,N_17500);
nand U19900 (N_19900,N_17149,N_18619);
and U19901 (N_19901,N_15938,N_16841);
and U19902 (N_19902,N_16896,N_18610);
or U19903 (N_19903,N_17137,N_16842);
and U19904 (N_19904,N_18285,N_16236);
nor U19905 (N_19905,N_16417,N_17950);
and U19906 (N_19906,N_18459,N_17941);
nand U19907 (N_19907,N_17216,N_17986);
xnor U19908 (N_19908,N_17921,N_16933);
and U19909 (N_19909,N_18212,N_17834);
or U19910 (N_19910,N_16163,N_17481);
and U19911 (N_19911,N_16166,N_17642);
xor U19912 (N_19912,N_18067,N_18113);
xor U19913 (N_19913,N_15693,N_18605);
xnor U19914 (N_19914,N_18693,N_17309);
nand U19915 (N_19915,N_16651,N_16391);
or U19916 (N_19916,N_16442,N_18337);
xor U19917 (N_19917,N_18126,N_15656);
and U19918 (N_19918,N_15965,N_16936);
or U19919 (N_19919,N_18419,N_16744);
xnor U19920 (N_19920,N_16183,N_17933);
nand U19921 (N_19921,N_18732,N_16109);
or U19922 (N_19922,N_18444,N_18411);
nand U19923 (N_19923,N_15910,N_18103);
or U19924 (N_19924,N_18593,N_17509);
or U19925 (N_19925,N_18440,N_16227);
nand U19926 (N_19926,N_16434,N_16297);
nand U19927 (N_19927,N_17134,N_18636);
and U19928 (N_19928,N_17797,N_16643);
nand U19929 (N_19929,N_18389,N_16246);
xor U19930 (N_19930,N_16588,N_17878);
xnor U19931 (N_19931,N_17825,N_17182);
or U19932 (N_19932,N_16657,N_18451);
xor U19933 (N_19933,N_17033,N_16692);
or U19934 (N_19934,N_17568,N_18283);
or U19935 (N_19935,N_17232,N_16903);
nor U19936 (N_19936,N_17203,N_15714);
and U19937 (N_19937,N_18508,N_18249);
and U19938 (N_19938,N_16851,N_18719);
nand U19939 (N_19939,N_17234,N_16828);
and U19940 (N_19940,N_17065,N_17893);
xnor U19941 (N_19941,N_16575,N_15720);
nand U19942 (N_19942,N_17696,N_17874);
or U19943 (N_19943,N_18731,N_17036);
xnor U19944 (N_19944,N_15761,N_18668);
and U19945 (N_19945,N_18481,N_16804);
or U19946 (N_19946,N_17866,N_17661);
or U19947 (N_19947,N_16635,N_17320);
and U19948 (N_19948,N_17487,N_16606);
or U19949 (N_19949,N_17012,N_17127);
nor U19950 (N_19950,N_18602,N_17150);
or U19951 (N_19951,N_18503,N_16890);
nor U19952 (N_19952,N_17858,N_15864);
nand U19953 (N_19953,N_16347,N_17113);
xor U19954 (N_19954,N_16173,N_16029);
xor U19955 (N_19955,N_16288,N_16506);
or U19956 (N_19956,N_16006,N_16687);
xor U19957 (N_19957,N_16709,N_17875);
nand U19958 (N_19958,N_18037,N_18377);
xnor U19959 (N_19959,N_17905,N_15847);
and U19960 (N_19960,N_17692,N_18414);
or U19961 (N_19961,N_18202,N_18280);
nor U19962 (N_19962,N_16126,N_16886);
nand U19963 (N_19963,N_18294,N_16421);
or U19964 (N_19964,N_16202,N_16462);
and U19965 (N_19965,N_18205,N_16818);
nor U19966 (N_19966,N_17862,N_15934);
nand U19967 (N_19967,N_15718,N_18670);
nor U19968 (N_19968,N_16974,N_16217);
or U19969 (N_19969,N_18564,N_16309);
or U19970 (N_19970,N_17056,N_17122);
nand U19971 (N_19971,N_15883,N_18742);
and U19972 (N_19972,N_17254,N_17451);
and U19973 (N_19973,N_16927,N_16176);
or U19974 (N_19974,N_17381,N_18589);
nand U19975 (N_19975,N_16711,N_18497);
xnor U19976 (N_19976,N_15638,N_16955);
nand U19977 (N_19977,N_18129,N_17969);
xnor U19978 (N_19978,N_15904,N_17053);
and U19979 (N_19979,N_15670,N_16919);
xor U19980 (N_19980,N_17754,N_16825);
or U19981 (N_19981,N_17835,N_16589);
nor U19982 (N_19982,N_17603,N_16853);
nand U19983 (N_19983,N_16926,N_16696);
or U19984 (N_19984,N_18487,N_17965);
xnor U19985 (N_19985,N_16947,N_17209);
nor U19986 (N_19986,N_17131,N_18200);
xnor U19987 (N_19987,N_18248,N_17171);
or U19988 (N_19988,N_15971,N_17519);
xnor U19989 (N_19989,N_18275,N_16674);
and U19990 (N_19990,N_17125,N_16271);
xor U19991 (N_19991,N_17355,N_17429);
nor U19992 (N_19992,N_18584,N_18471);
nor U19993 (N_19993,N_18051,N_17250);
xnor U19994 (N_19994,N_15661,N_16142);
and U19995 (N_19995,N_15733,N_16906);
or U19996 (N_19996,N_17050,N_16168);
xnor U19997 (N_19997,N_17495,N_18675);
nand U19998 (N_19998,N_18630,N_16165);
nand U19999 (N_19999,N_18194,N_16198);
xnor U20000 (N_20000,N_16784,N_18717);
or U20001 (N_20001,N_16791,N_17035);
nor U20002 (N_20002,N_16763,N_17274);
nor U20003 (N_20003,N_17459,N_17336);
nor U20004 (N_20004,N_17959,N_16186);
nand U20005 (N_20005,N_15887,N_17886);
or U20006 (N_20006,N_16501,N_16058);
xnor U20007 (N_20007,N_17449,N_15729);
nand U20008 (N_20008,N_17217,N_17244);
and U20009 (N_20009,N_16539,N_15770);
or U20010 (N_20010,N_17994,N_16011);
or U20011 (N_20011,N_17877,N_17975);
xor U20012 (N_20012,N_15668,N_17493);
nor U20013 (N_20013,N_16041,N_18022);
or U20014 (N_20014,N_17397,N_16306);
nor U20015 (N_20015,N_17432,N_16509);
nand U20016 (N_20016,N_15708,N_16151);
nand U20017 (N_20017,N_16756,N_15992);
or U20018 (N_20018,N_18080,N_18730);
xnor U20019 (N_20019,N_17978,N_17337);
nor U20020 (N_20020,N_15968,N_18351);
nand U20021 (N_20021,N_18531,N_16348);
xnor U20022 (N_20022,N_17632,N_18229);
xor U20023 (N_20023,N_18150,N_18148);
and U20024 (N_20024,N_18671,N_16508);
and U20025 (N_20025,N_18303,N_17623);
or U20026 (N_20026,N_17408,N_16320);
and U20027 (N_20027,N_18501,N_16047);
nor U20028 (N_20028,N_17016,N_17346);
nand U20029 (N_20029,N_18288,N_16898);
nand U20030 (N_20030,N_16807,N_16984);
nand U20031 (N_20031,N_15810,N_15803);
nor U20032 (N_20032,N_16212,N_16087);
xor U20033 (N_20033,N_18432,N_18089);
or U20034 (N_20034,N_18450,N_16067);
xor U20035 (N_20035,N_17376,N_17636);
xor U20036 (N_20036,N_16498,N_16707);
and U20037 (N_20037,N_17864,N_18533);
xnor U20038 (N_20038,N_16135,N_16740);
and U20039 (N_20039,N_17840,N_15806);
or U20040 (N_20040,N_15956,N_15823);
xor U20041 (N_20041,N_17272,N_16250);
or U20042 (N_20042,N_17457,N_17628);
nor U20043 (N_20043,N_16256,N_17729);
and U20044 (N_20044,N_16452,N_17401);
xnor U20045 (N_20045,N_16438,N_17763);
xor U20046 (N_20046,N_18074,N_18673);
nor U20047 (N_20047,N_16601,N_17275);
or U20048 (N_20048,N_18298,N_17733);
xnor U20049 (N_20049,N_16005,N_16294);
nand U20050 (N_20050,N_15946,N_17108);
nor U20051 (N_20051,N_16910,N_17787);
nor U20052 (N_20052,N_16244,N_16669);
nor U20053 (N_20053,N_16423,N_16612);
nor U20054 (N_20054,N_15743,N_16985);
or U20055 (N_20055,N_16193,N_17778);
nor U20056 (N_20056,N_15750,N_16050);
nor U20057 (N_20057,N_16277,N_16318);
nor U20058 (N_20058,N_17360,N_16012);
or U20059 (N_20059,N_16532,N_15702);
or U20060 (N_20060,N_16973,N_18664);
nor U20061 (N_20061,N_18676,N_17020);
nor U20062 (N_20062,N_16153,N_17394);
nand U20063 (N_20063,N_16546,N_15774);
or U20064 (N_20064,N_17765,N_15760);
nor U20065 (N_20065,N_17676,N_18199);
nor U20066 (N_20066,N_16504,N_16499);
and U20067 (N_20067,N_16668,N_18060);
or U20068 (N_20068,N_16704,N_18179);
nor U20069 (N_20069,N_17123,N_17427);
or U20070 (N_20070,N_17022,N_16971);
nand U20071 (N_20071,N_17475,N_18442);
and U20072 (N_20072,N_17253,N_17593);
nand U20073 (N_20073,N_16386,N_18690);
or U20074 (N_20074,N_17477,N_17513);
nor U20075 (N_20075,N_17470,N_17335);
nor U20076 (N_20076,N_16998,N_16676);
or U20077 (N_20077,N_16171,N_16917);
or U20078 (N_20078,N_17327,N_15999);
or U20079 (N_20079,N_16441,N_17191);
and U20080 (N_20080,N_17472,N_18112);
nand U20081 (N_20081,N_16901,N_16562);
nor U20082 (N_20082,N_16483,N_16341);
nor U20083 (N_20083,N_18588,N_17667);
nor U20084 (N_20084,N_18418,N_17803);
nand U20085 (N_20085,N_16745,N_17396);
nor U20086 (N_20086,N_18702,N_16778);
xnor U20087 (N_20087,N_17003,N_17075);
and U20088 (N_20088,N_17238,N_17548);
nor U20089 (N_20089,N_16681,N_17618);
or U20090 (N_20090,N_17815,N_17425);
nand U20091 (N_20091,N_17007,N_15922);
and U20092 (N_20092,N_17277,N_17010);
or U20093 (N_20093,N_15721,N_16848);
xor U20094 (N_20094,N_16869,N_16981);
xnor U20095 (N_20095,N_17339,N_16480);
nor U20096 (N_20096,N_15878,N_17385);
nand U20097 (N_20097,N_17584,N_18137);
nor U20098 (N_20098,N_16114,N_18317);
or U20099 (N_20099,N_16215,N_16799);
and U20100 (N_20100,N_17371,N_16574);
or U20101 (N_20101,N_18680,N_18328);
or U20102 (N_20102,N_18516,N_17947);
xor U20103 (N_20103,N_15676,N_17907);
or U20104 (N_20104,N_17522,N_15988);
or U20105 (N_20105,N_18566,N_16266);
xnor U20106 (N_20106,N_17179,N_15755);
xor U20107 (N_20107,N_17574,N_17059);
nor U20108 (N_20108,N_17839,N_17788);
xnor U20109 (N_20109,N_16628,N_16529);
or U20110 (N_20110,N_17178,N_18024);
or U20111 (N_20111,N_17930,N_18271);
nand U20112 (N_20112,N_16817,N_18186);
nor U20113 (N_20113,N_18127,N_17001);
xor U20114 (N_20114,N_15835,N_18648);
nand U20115 (N_20115,N_16889,N_16647);
nand U20116 (N_20116,N_15811,N_16111);
or U20117 (N_20117,N_16351,N_17920);
nand U20118 (N_20118,N_15903,N_16366);
and U20119 (N_20119,N_18334,N_16714);
xor U20120 (N_20120,N_18048,N_15906);
or U20121 (N_20121,N_17353,N_16080);
and U20122 (N_20122,N_16824,N_16346);
nor U20123 (N_20123,N_15723,N_18091);
nor U20124 (N_20124,N_16518,N_18441);
and U20125 (N_20125,N_16968,N_17489);
nand U20126 (N_20126,N_15764,N_15912);
xnor U20127 (N_20127,N_16302,N_16360);
nor U20128 (N_20128,N_15697,N_15895);
nor U20129 (N_20129,N_17988,N_16970);
nor U20130 (N_20130,N_15725,N_17937);
and U20131 (N_20131,N_17782,N_18243);
nand U20132 (N_20132,N_16623,N_16377);
xnor U20133 (N_20133,N_18176,N_17102);
or U20134 (N_20134,N_18725,N_16697);
and U20135 (N_20135,N_16431,N_17367);
or U20136 (N_20136,N_17991,N_17330);
and U20137 (N_20137,N_17902,N_17440);
nor U20138 (N_20138,N_16376,N_17208);
or U20139 (N_20139,N_17520,N_17617);
or U20140 (N_20140,N_15698,N_16661);
and U20141 (N_20141,N_17979,N_16081);
nor U20142 (N_20142,N_18209,N_18252);
and U20143 (N_20143,N_16032,N_18474);
and U20144 (N_20144,N_16316,N_16492);
xor U20145 (N_20145,N_17749,N_17836);
xor U20146 (N_20146,N_17018,N_17784);
and U20147 (N_20147,N_15997,N_17247);
nor U20148 (N_20148,N_16472,N_17221);
xnor U20149 (N_20149,N_17856,N_16631);
and U20150 (N_20150,N_18064,N_16008);
or U20151 (N_20151,N_18592,N_16572);
nor U20152 (N_20152,N_16337,N_16339);
or U20153 (N_20153,N_17641,N_15695);
xor U20154 (N_20154,N_18323,N_18314);
or U20155 (N_20155,N_17927,N_16859);
nand U20156 (N_20156,N_17735,N_16808);
nand U20157 (N_20157,N_17322,N_15935);
nor U20158 (N_20158,N_16473,N_16798);
and U20159 (N_20159,N_16096,N_18181);
and U20160 (N_20160,N_16630,N_17849);
or U20161 (N_20161,N_17496,N_17870);
or U20162 (N_20162,N_16030,N_17960);
nor U20163 (N_20163,N_16723,N_17079);
or U20164 (N_20164,N_18341,N_15807);
and U20165 (N_20165,N_16584,N_16672);
and U20166 (N_20166,N_17985,N_17406);
nor U20167 (N_20167,N_18598,N_15987);
xnor U20168 (N_20168,N_18625,N_17111);
xnor U20169 (N_20169,N_16036,N_16027);
or U20170 (N_20170,N_16290,N_15731);
nand U20171 (N_20171,N_16040,N_18168);
or U20172 (N_20172,N_16928,N_18367);
and U20173 (N_20173,N_16809,N_16512);
or U20174 (N_20174,N_17805,N_18669);
nor U20175 (N_20175,N_18467,N_16296);
nand U20176 (N_20176,N_16226,N_15710);
and U20177 (N_20177,N_18327,N_17701);
and U20178 (N_20178,N_17467,N_16913);
nand U20179 (N_20179,N_16424,N_16304);
and U20180 (N_20180,N_16622,N_17917);
xnor U20181 (N_20181,N_17343,N_17608);
xor U20182 (N_20182,N_18698,N_16821);
and U20183 (N_20183,N_18286,N_16565);
nor U20184 (N_20184,N_15651,N_17129);
or U20185 (N_20185,N_18740,N_18391);
or U20186 (N_20186,N_15836,N_15794);
xor U20187 (N_20187,N_16458,N_15737);
nor U20188 (N_20188,N_18153,N_16273);
xnor U20189 (N_20189,N_17474,N_16222);
or U20190 (N_20190,N_16057,N_16285);
nor U20191 (N_20191,N_17492,N_17407);
and U20192 (N_20192,N_16683,N_16838);
or U20193 (N_20193,N_16311,N_18226);
nand U20194 (N_20194,N_17454,N_17080);
xor U20195 (N_20195,N_15947,N_17717);
nand U20196 (N_20196,N_18380,N_18122);
nor U20197 (N_20197,N_17748,N_17262);
and U20198 (N_20198,N_17657,N_16089);
nor U20199 (N_20199,N_17292,N_17061);
or U20200 (N_20200,N_16969,N_16468);
or U20201 (N_20201,N_16924,N_16678);
or U20202 (N_20202,N_18490,N_17365);
nand U20203 (N_20203,N_17174,N_16427);
and U20204 (N_20204,N_18388,N_17433);
and U20205 (N_20205,N_15998,N_17231);
nand U20206 (N_20206,N_16735,N_16787);
or U20207 (N_20207,N_17066,N_17779);
nor U20208 (N_20208,N_17556,N_16450);
or U20209 (N_20209,N_17808,N_16796);
nand U20210 (N_20210,N_18156,N_17776);
or U20211 (N_20211,N_16534,N_17892);
nor U20212 (N_20212,N_17939,N_16536);
xnor U20213 (N_20213,N_16958,N_18301);
and U20214 (N_20214,N_16496,N_17094);
xnor U20215 (N_20215,N_18530,N_17543);
and U20216 (N_20216,N_16522,N_17704);
and U20217 (N_20217,N_16561,N_17611);
and U20218 (N_20218,N_16724,N_18478);
or U20219 (N_20219,N_17572,N_16945);
or U20220 (N_20220,N_16991,N_17243);
and U20221 (N_20221,N_16167,N_15784);
or U20222 (N_20222,N_17562,N_17785);
or U20223 (N_20223,N_16042,N_16060);
xor U20224 (N_20224,N_15771,N_17074);
nand U20225 (N_20225,N_17378,N_17802);
and U20226 (N_20226,N_18606,N_18703);
nor U20227 (N_20227,N_16604,N_16571);
or U20228 (N_20228,N_18118,N_17838);
nand U20229 (N_20229,N_17400,N_18453);
nand U20230 (N_20230,N_17541,N_15853);
xor U20231 (N_20231,N_17561,N_18744);
nand U20232 (N_20232,N_16872,N_18131);
nand U20233 (N_20233,N_16870,N_16716);
and U20234 (N_20234,N_17382,N_17531);
nor U20235 (N_20235,N_18443,N_17404);
nand U20236 (N_20236,N_17120,N_18214);
nand U20237 (N_20237,N_17212,N_17602);
nand U20238 (N_20238,N_17045,N_18215);
and U20239 (N_20239,N_17328,N_16642);
nand U20240 (N_20240,N_16303,N_17411);
and U20241 (N_20241,N_16122,N_17442);
nand U20242 (N_20242,N_17795,N_17499);
nor U20243 (N_20243,N_16228,N_17285);
xnor U20244 (N_20244,N_16685,N_17518);
nor U20245 (N_20245,N_17071,N_16197);
nand U20246 (N_20246,N_17104,N_16840);
xnor U20247 (N_20247,N_18076,N_16487);
xor U20248 (N_20248,N_18649,N_16449);
xor U20249 (N_20249,N_17412,N_18183);
nand U20250 (N_20250,N_16733,N_16771);
xnor U20251 (N_20251,N_16270,N_17846);
nor U20252 (N_20252,N_17504,N_18135);
nor U20253 (N_20253,N_16570,N_16191);
and U20254 (N_20254,N_16321,N_17598);
or U20255 (N_20255,N_17468,N_16757);
and U20256 (N_20256,N_17290,N_17478);
nor U20257 (N_20257,N_16978,N_17280);
nand U20258 (N_20258,N_15993,N_18570);
nand U20259 (N_20259,N_16597,N_15849);
and U20260 (N_20260,N_17357,N_17334);
nand U20261 (N_20261,N_17265,N_17610);
and U20262 (N_20262,N_17047,N_17647);
or U20263 (N_20263,N_15927,N_16263);
or U20264 (N_20264,N_17516,N_16014);
and U20265 (N_20265,N_17842,N_17654);
nor U20266 (N_20266,N_15862,N_18581);
xnor U20267 (N_20267,N_16867,N_18518);
or U20268 (N_20268,N_16555,N_16293);
and U20269 (N_20269,N_17291,N_17258);
nand U20270 (N_20270,N_16110,N_18682);
nand U20271 (N_20271,N_16383,N_16788);
or U20272 (N_20272,N_17391,N_17963);
xor U20273 (N_20273,N_18348,N_15765);
or U20274 (N_20274,N_17833,N_18534);
xor U20275 (N_20275,N_18141,N_18572);
xor U20276 (N_20276,N_15712,N_15677);
nor U20277 (N_20277,N_18517,N_15916);
and U20278 (N_20278,N_17609,N_16613);
nor U20279 (N_20279,N_17146,N_15792);
and U20280 (N_20280,N_17908,N_17682);
xor U20281 (N_20281,N_18057,N_16363);
and U20282 (N_20282,N_16237,N_16519);
xnor U20283 (N_20283,N_18526,N_17049);
and U20284 (N_20284,N_18073,N_17494);
nand U20285 (N_20285,N_17366,N_16686);
nor U20286 (N_20286,N_18040,N_18291);
or U20287 (N_20287,N_15838,N_16829);
or U20288 (N_20288,N_17708,N_17448);
nand U20289 (N_20289,N_16090,N_18582);
or U20290 (N_20290,N_16214,N_15663);
nand U20291 (N_20291,N_16908,N_18138);
or U20292 (N_20292,N_17379,N_15827);
or U20293 (N_20293,N_16600,N_16203);
and U20294 (N_20294,N_17106,N_15978);
nand U20295 (N_20295,N_17887,N_16385);
nand U20296 (N_20296,N_18395,N_18511);
nor U20297 (N_20297,N_17847,N_17726);
nand U20298 (N_20298,N_17664,N_18227);
nor U20299 (N_20299,N_18230,N_18576);
nand U20300 (N_20300,N_18055,N_16713);
xnor U20301 (N_20301,N_18727,N_17316);
xnor U20302 (N_20302,N_16482,N_16545);
nand U20303 (N_20303,N_16905,N_17260);
xnor U20304 (N_20304,N_17167,N_16358);
and U20305 (N_20305,N_16258,N_16852);
and U20306 (N_20306,N_18182,N_16695);
or U20307 (N_20307,N_17298,N_17083);
nor U20308 (N_20308,N_16598,N_17373);
nor U20309 (N_20309,N_17974,N_18386);
nand U20310 (N_20310,N_17176,N_18093);
nor U20311 (N_20311,N_16734,N_16875);
nand U20312 (N_20312,N_15966,N_18369);
nor U20313 (N_20313,N_17752,N_18390);
or U20314 (N_20314,N_16237,N_17472);
xor U20315 (N_20315,N_15865,N_16033);
xnor U20316 (N_20316,N_16650,N_16451);
nand U20317 (N_20317,N_18407,N_17462);
nand U20318 (N_20318,N_18409,N_16412);
xnor U20319 (N_20319,N_17239,N_15633);
xor U20320 (N_20320,N_16902,N_18159);
xnor U20321 (N_20321,N_18648,N_15945);
or U20322 (N_20322,N_17486,N_17758);
xor U20323 (N_20323,N_16723,N_15851);
or U20324 (N_20324,N_16024,N_17211);
or U20325 (N_20325,N_17050,N_18492);
nand U20326 (N_20326,N_16590,N_16755);
or U20327 (N_20327,N_16908,N_18451);
nand U20328 (N_20328,N_18208,N_16509);
or U20329 (N_20329,N_16224,N_18649);
or U20330 (N_20330,N_18170,N_16073);
nor U20331 (N_20331,N_17083,N_17533);
xor U20332 (N_20332,N_15758,N_17840);
and U20333 (N_20333,N_17355,N_17090);
nor U20334 (N_20334,N_17480,N_16561);
and U20335 (N_20335,N_17405,N_16971);
nor U20336 (N_20336,N_16812,N_18065);
xnor U20337 (N_20337,N_18335,N_18473);
xor U20338 (N_20338,N_17256,N_16792);
nor U20339 (N_20339,N_18068,N_17735);
or U20340 (N_20340,N_16737,N_16825);
nand U20341 (N_20341,N_17474,N_17909);
xnor U20342 (N_20342,N_15872,N_15768);
or U20343 (N_20343,N_17370,N_15905);
nand U20344 (N_20344,N_17201,N_16781);
nand U20345 (N_20345,N_18190,N_17394);
and U20346 (N_20346,N_15675,N_15968);
nor U20347 (N_20347,N_18586,N_16773);
nand U20348 (N_20348,N_17387,N_16284);
nor U20349 (N_20349,N_17963,N_15775);
nor U20350 (N_20350,N_18125,N_16283);
nor U20351 (N_20351,N_15831,N_17165);
xnor U20352 (N_20352,N_17062,N_16443);
nor U20353 (N_20353,N_16437,N_17295);
nor U20354 (N_20354,N_16634,N_18046);
nor U20355 (N_20355,N_18116,N_16756);
nor U20356 (N_20356,N_17594,N_16930);
xor U20357 (N_20357,N_16576,N_15653);
or U20358 (N_20358,N_18488,N_15696);
nor U20359 (N_20359,N_17783,N_18707);
nor U20360 (N_20360,N_15703,N_16129);
nor U20361 (N_20361,N_16041,N_18718);
nand U20362 (N_20362,N_17975,N_17525);
or U20363 (N_20363,N_16019,N_16186);
or U20364 (N_20364,N_16646,N_15844);
nand U20365 (N_20365,N_16248,N_15629);
xor U20366 (N_20366,N_18620,N_18476);
and U20367 (N_20367,N_17982,N_16265);
and U20368 (N_20368,N_16627,N_17292);
xor U20369 (N_20369,N_18407,N_17330);
xnor U20370 (N_20370,N_16770,N_16950);
nor U20371 (N_20371,N_17122,N_16606);
nand U20372 (N_20372,N_18672,N_18193);
xnor U20373 (N_20373,N_15921,N_18149);
and U20374 (N_20374,N_17710,N_17891);
or U20375 (N_20375,N_17765,N_18435);
and U20376 (N_20376,N_15989,N_16323);
nor U20377 (N_20377,N_17854,N_16190);
and U20378 (N_20378,N_15834,N_16773);
nand U20379 (N_20379,N_15739,N_17386);
or U20380 (N_20380,N_18093,N_18233);
nand U20381 (N_20381,N_17162,N_17516);
xor U20382 (N_20382,N_16738,N_17956);
and U20383 (N_20383,N_16512,N_15813);
xor U20384 (N_20384,N_16900,N_15913);
xnor U20385 (N_20385,N_17661,N_15847);
or U20386 (N_20386,N_17871,N_15881);
and U20387 (N_20387,N_17658,N_18194);
and U20388 (N_20388,N_15861,N_18709);
xor U20389 (N_20389,N_17507,N_16812);
and U20390 (N_20390,N_17877,N_18328);
or U20391 (N_20391,N_18203,N_18746);
xnor U20392 (N_20392,N_15990,N_18735);
or U20393 (N_20393,N_15653,N_18020);
and U20394 (N_20394,N_16985,N_16901);
nand U20395 (N_20395,N_16165,N_17228);
or U20396 (N_20396,N_17726,N_16309);
and U20397 (N_20397,N_16230,N_16822);
or U20398 (N_20398,N_18643,N_16573);
nor U20399 (N_20399,N_15834,N_18004);
nor U20400 (N_20400,N_17477,N_15784);
nor U20401 (N_20401,N_15901,N_18722);
xor U20402 (N_20402,N_16450,N_17684);
nor U20403 (N_20403,N_18203,N_16831);
nor U20404 (N_20404,N_16829,N_18118);
nor U20405 (N_20405,N_15667,N_18178);
or U20406 (N_20406,N_17526,N_16438);
and U20407 (N_20407,N_18693,N_16665);
nor U20408 (N_20408,N_15966,N_15923);
nand U20409 (N_20409,N_17193,N_17853);
nand U20410 (N_20410,N_17287,N_16296);
or U20411 (N_20411,N_17949,N_17448);
or U20412 (N_20412,N_16918,N_17004);
nor U20413 (N_20413,N_18280,N_18433);
nand U20414 (N_20414,N_18595,N_18374);
or U20415 (N_20415,N_18184,N_16130);
nor U20416 (N_20416,N_17314,N_16537);
nor U20417 (N_20417,N_16750,N_17944);
or U20418 (N_20418,N_17732,N_18623);
xor U20419 (N_20419,N_18668,N_16544);
nand U20420 (N_20420,N_16915,N_17822);
nor U20421 (N_20421,N_17244,N_17226);
and U20422 (N_20422,N_17921,N_15998);
nor U20423 (N_20423,N_18283,N_17015);
xor U20424 (N_20424,N_17155,N_18501);
or U20425 (N_20425,N_17631,N_17525);
xor U20426 (N_20426,N_15789,N_16575);
and U20427 (N_20427,N_16983,N_17597);
or U20428 (N_20428,N_18526,N_16501);
xor U20429 (N_20429,N_16938,N_17810);
nand U20430 (N_20430,N_17285,N_16404);
nand U20431 (N_20431,N_16196,N_17068);
nand U20432 (N_20432,N_16492,N_16800);
nor U20433 (N_20433,N_17370,N_16341);
xor U20434 (N_20434,N_18561,N_16672);
xor U20435 (N_20435,N_15745,N_17377);
or U20436 (N_20436,N_17680,N_16508);
xor U20437 (N_20437,N_17696,N_17320);
nor U20438 (N_20438,N_16427,N_18442);
or U20439 (N_20439,N_17989,N_18074);
and U20440 (N_20440,N_16979,N_17440);
xor U20441 (N_20441,N_18703,N_18191);
nor U20442 (N_20442,N_16558,N_17029);
nor U20443 (N_20443,N_18413,N_18218);
nand U20444 (N_20444,N_16458,N_18103);
xor U20445 (N_20445,N_18515,N_17589);
nand U20446 (N_20446,N_16942,N_16882);
or U20447 (N_20447,N_16495,N_17789);
and U20448 (N_20448,N_16101,N_17526);
nor U20449 (N_20449,N_16548,N_16180);
and U20450 (N_20450,N_16481,N_18060);
xor U20451 (N_20451,N_17977,N_16450);
nand U20452 (N_20452,N_18724,N_17885);
and U20453 (N_20453,N_16256,N_17688);
xnor U20454 (N_20454,N_16232,N_17051);
xnor U20455 (N_20455,N_16537,N_16914);
and U20456 (N_20456,N_17461,N_16994);
or U20457 (N_20457,N_17654,N_17963);
nor U20458 (N_20458,N_18323,N_17154);
or U20459 (N_20459,N_16011,N_16724);
xor U20460 (N_20460,N_18202,N_15788);
and U20461 (N_20461,N_17084,N_15741);
nor U20462 (N_20462,N_15821,N_16213);
and U20463 (N_20463,N_16587,N_16247);
xor U20464 (N_20464,N_16498,N_17649);
or U20465 (N_20465,N_17200,N_17527);
and U20466 (N_20466,N_17917,N_15631);
and U20467 (N_20467,N_17714,N_17830);
nor U20468 (N_20468,N_18665,N_18186);
or U20469 (N_20469,N_16910,N_16361);
xor U20470 (N_20470,N_16491,N_17896);
nor U20471 (N_20471,N_17128,N_18125);
and U20472 (N_20472,N_17084,N_17202);
and U20473 (N_20473,N_18172,N_15824);
and U20474 (N_20474,N_18497,N_18292);
nand U20475 (N_20475,N_17396,N_16276);
nand U20476 (N_20476,N_18243,N_15718);
or U20477 (N_20477,N_18138,N_17779);
nor U20478 (N_20478,N_17352,N_17541);
nor U20479 (N_20479,N_16257,N_16298);
nand U20480 (N_20480,N_15825,N_16290);
or U20481 (N_20481,N_18002,N_18182);
xor U20482 (N_20482,N_15713,N_16402);
xnor U20483 (N_20483,N_18251,N_17025);
xor U20484 (N_20484,N_17526,N_17710);
or U20485 (N_20485,N_16033,N_15829);
and U20486 (N_20486,N_17297,N_18004);
xor U20487 (N_20487,N_16783,N_16376);
nor U20488 (N_20488,N_15854,N_17323);
or U20489 (N_20489,N_18099,N_17467);
or U20490 (N_20490,N_16363,N_17406);
nor U20491 (N_20491,N_15662,N_16923);
or U20492 (N_20492,N_17925,N_16269);
and U20493 (N_20493,N_17703,N_16137);
and U20494 (N_20494,N_17212,N_17512);
and U20495 (N_20495,N_18367,N_18629);
and U20496 (N_20496,N_16364,N_17784);
xor U20497 (N_20497,N_16584,N_17542);
nor U20498 (N_20498,N_16131,N_16343);
xnor U20499 (N_20499,N_17195,N_16757);
nor U20500 (N_20500,N_17734,N_18095);
nand U20501 (N_20501,N_16925,N_16420);
and U20502 (N_20502,N_16905,N_17184);
and U20503 (N_20503,N_17683,N_16054);
nor U20504 (N_20504,N_16528,N_15880);
nor U20505 (N_20505,N_17891,N_17893);
xor U20506 (N_20506,N_17950,N_16375);
nor U20507 (N_20507,N_15855,N_16872);
nand U20508 (N_20508,N_17281,N_16226);
nand U20509 (N_20509,N_17178,N_16023);
nor U20510 (N_20510,N_17617,N_16653);
nand U20511 (N_20511,N_17395,N_17343);
or U20512 (N_20512,N_17589,N_16998);
xnor U20513 (N_20513,N_18199,N_16552);
and U20514 (N_20514,N_15641,N_17267);
nor U20515 (N_20515,N_16959,N_17178);
or U20516 (N_20516,N_16201,N_18477);
nand U20517 (N_20517,N_16063,N_17147);
nand U20518 (N_20518,N_15870,N_16292);
nand U20519 (N_20519,N_16955,N_18521);
or U20520 (N_20520,N_18397,N_15980);
or U20521 (N_20521,N_18165,N_18714);
xnor U20522 (N_20522,N_17425,N_17060);
or U20523 (N_20523,N_17192,N_16120);
nand U20524 (N_20524,N_16696,N_16672);
xor U20525 (N_20525,N_15992,N_17239);
xor U20526 (N_20526,N_18332,N_17759);
or U20527 (N_20527,N_18533,N_16697);
and U20528 (N_20528,N_15758,N_15683);
xnor U20529 (N_20529,N_18206,N_17850);
or U20530 (N_20530,N_16578,N_18244);
and U20531 (N_20531,N_17499,N_16287);
nand U20532 (N_20532,N_17246,N_16303);
and U20533 (N_20533,N_16390,N_18338);
nor U20534 (N_20534,N_18132,N_18450);
xor U20535 (N_20535,N_15732,N_18405);
nand U20536 (N_20536,N_18625,N_17275);
nor U20537 (N_20537,N_17333,N_17479);
and U20538 (N_20538,N_18324,N_16707);
and U20539 (N_20539,N_16863,N_16464);
xor U20540 (N_20540,N_15819,N_18624);
nor U20541 (N_20541,N_16015,N_16024);
nor U20542 (N_20542,N_16244,N_18172);
or U20543 (N_20543,N_17751,N_15674);
and U20544 (N_20544,N_15913,N_16788);
nand U20545 (N_20545,N_17748,N_17166);
xor U20546 (N_20546,N_18050,N_16356);
and U20547 (N_20547,N_16803,N_16952);
nand U20548 (N_20548,N_16679,N_16933);
nand U20549 (N_20549,N_16605,N_18003);
nor U20550 (N_20550,N_16351,N_18658);
xor U20551 (N_20551,N_16749,N_16486);
xnor U20552 (N_20552,N_15746,N_16401);
nor U20553 (N_20553,N_16264,N_18554);
or U20554 (N_20554,N_16481,N_18312);
xor U20555 (N_20555,N_15763,N_17679);
and U20556 (N_20556,N_18038,N_17482);
nand U20557 (N_20557,N_17778,N_16363);
and U20558 (N_20558,N_17500,N_17542);
nand U20559 (N_20559,N_16719,N_18682);
and U20560 (N_20560,N_17486,N_17273);
and U20561 (N_20561,N_17026,N_16983);
xor U20562 (N_20562,N_15770,N_17333);
xor U20563 (N_20563,N_15837,N_16687);
xnor U20564 (N_20564,N_18323,N_18341);
xor U20565 (N_20565,N_18394,N_16877);
xnor U20566 (N_20566,N_18155,N_15696);
and U20567 (N_20567,N_15867,N_17095);
nor U20568 (N_20568,N_18366,N_18677);
or U20569 (N_20569,N_15655,N_17390);
and U20570 (N_20570,N_17246,N_17623);
xor U20571 (N_20571,N_16268,N_18587);
xor U20572 (N_20572,N_16363,N_16466);
xnor U20573 (N_20573,N_17751,N_16778);
and U20574 (N_20574,N_16990,N_18593);
nor U20575 (N_20575,N_16190,N_16305);
xnor U20576 (N_20576,N_16297,N_16514);
or U20577 (N_20577,N_16136,N_16462);
nor U20578 (N_20578,N_17920,N_18363);
or U20579 (N_20579,N_17056,N_16456);
and U20580 (N_20580,N_15950,N_17009);
nor U20581 (N_20581,N_15699,N_18008);
nand U20582 (N_20582,N_18128,N_16918);
nor U20583 (N_20583,N_17995,N_16112);
or U20584 (N_20584,N_18156,N_17353);
and U20585 (N_20585,N_17391,N_18147);
xnor U20586 (N_20586,N_16556,N_18507);
nand U20587 (N_20587,N_18233,N_18196);
nand U20588 (N_20588,N_17899,N_17321);
and U20589 (N_20589,N_16331,N_17828);
xor U20590 (N_20590,N_16062,N_16543);
and U20591 (N_20591,N_15786,N_16196);
or U20592 (N_20592,N_16765,N_16563);
or U20593 (N_20593,N_17495,N_17912);
xnor U20594 (N_20594,N_18621,N_17326);
nand U20595 (N_20595,N_15753,N_16865);
nor U20596 (N_20596,N_18706,N_16856);
xnor U20597 (N_20597,N_18093,N_18306);
or U20598 (N_20598,N_17076,N_16844);
and U20599 (N_20599,N_18576,N_17346);
or U20600 (N_20600,N_15797,N_16564);
xnor U20601 (N_20601,N_17543,N_17749);
nor U20602 (N_20602,N_17003,N_17872);
xor U20603 (N_20603,N_16785,N_18735);
and U20604 (N_20604,N_16920,N_16965);
nand U20605 (N_20605,N_16744,N_16480);
nor U20606 (N_20606,N_17442,N_18540);
xnor U20607 (N_20607,N_17463,N_16803);
nand U20608 (N_20608,N_17294,N_17730);
and U20609 (N_20609,N_18252,N_16600);
xor U20610 (N_20610,N_18305,N_16679);
nand U20611 (N_20611,N_16935,N_18484);
nor U20612 (N_20612,N_18626,N_15749);
and U20613 (N_20613,N_16756,N_17115);
xor U20614 (N_20614,N_18677,N_16320);
nor U20615 (N_20615,N_15836,N_18313);
and U20616 (N_20616,N_16229,N_15704);
nor U20617 (N_20617,N_18300,N_16133);
nand U20618 (N_20618,N_16353,N_17683);
xnor U20619 (N_20619,N_17129,N_18461);
xor U20620 (N_20620,N_18593,N_17702);
nand U20621 (N_20621,N_17722,N_18601);
nand U20622 (N_20622,N_18388,N_16539);
nor U20623 (N_20623,N_16427,N_18174);
xor U20624 (N_20624,N_15904,N_15657);
nor U20625 (N_20625,N_18706,N_16690);
or U20626 (N_20626,N_18111,N_17175);
xnor U20627 (N_20627,N_16494,N_16095);
nand U20628 (N_20628,N_16612,N_17134);
nor U20629 (N_20629,N_17117,N_17688);
nand U20630 (N_20630,N_17502,N_17085);
or U20631 (N_20631,N_18478,N_17351);
and U20632 (N_20632,N_17427,N_16834);
xor U20633 (N_20633,N_17676,N_18334);
or U20634 (N_20634,N_16314,N_16467);
nor U20635 (N_20635,N_15632,N_18512);
nand U20636 (N_20636,N_18278,N_16511);
xor U20637 (N_20637,N_16982,N_16057);
xnor U20638 (N_20638,N_16817,N_16916);
and U20639 (N_20639,N_18415,N_17073);
nor U20640 (N_20640,N_17037,N_16118);
xor U20641 (N_20641,N_16988,N_17348);
nand U20642 (N_20642,N_17685,N_15693);
xor U20643 (N_20643,N_17270,N_17620);
nand U20644 (N_20644,N_17246,N_16831);
or U20645 (N_20645,N_15682,N_16659);
xor U20646 (N_20646,N_16100,N_16393);
nor U20647 (N_20647,N_15648,N_18045);
and U20648 (N_20648,N_15892,N_16556);
and U20649 (N_20649,N_16778,N_17268);
xnor U20650 (N_20650,N_18429,N_16724);
nor U20651 (N_20651,N_17010,N_16921);
nor U20652 (N_20652,N_16481,N_16083);
and U20653 (N_20653,N_17759,N_17512);
or U20654 (N_20654,N_17862,N_16515);
xnor U20655 (N_20655,N_17265,N_16993);
nor U20656 (N_20656,N_17858,N_16884);
or U20657 (N_20657,N_16966,N_16853);
and U20658 (N_20658,N_16111,N_16044);
nand U20659 (N_20659,N_15891,N_17502);
xnor U20660 (N_20660,N_18118,N_17564);
nand U20661 (N_20661,N_18269,N_17426);
nand U20662 (N_20662,N_17253,N_18082);
nor U20663 (N_20663,N_18154,N_15698);
and U20664 (N_20664,N_18089,N_15689);
xor U20665 (N_20665,N_16287,N_15816);
or U20666 (N_20666,N_17159,N_15906);
or U20667 (N_20667,N_17925,N_16487);
nand U20668 (N_20668,N_17256,N_15938);
or U20669 (N_20669,N_16663,N_16194);
or U20670 (N_20670,N_17809,N_16845);
nand U20671 (N_20671,N_17511,N_18194);
nand U20672 (N_20672,N_17190,N_17475);
nor U20673 (N_20673,N_18445,N_17482);
xor U20674 (N_20674,N_17537,N_15799);
or U20675 (N_20675,N_18630,N_16972);
nand U20676 (N_20676,N_18740,N_17676);
xor U20677 (N_20677,N_17211,N_16520);
nand U20678 (N_20678,N_17593,N_15908);
xor U20679 (N_20679,N_16951,N_17163);
nor U20680 (N_20680,N_18351,N_18325);
nand U20681 (N_20681,N_17107,N_17337);
nor U20682 (N_20682,N_18728,N_17462);
nor U20683 (N_20683,N_18199,N_16072);
nor U20684 (N_20684,N_15807,N_16633);
xnor U20685 (N_20685,N_18102,N_15656);
nor U20686 (N_20686,N_17841,N_15731);
or U20687 (N_20687,N_17637,N_17082);
nand U20688 (N_20688,N_17711,N_17437);
and U20689 (N_20689,N_16561,N_18086);
nor U20690 (N_20690,N_18430,N_17677);
and U20691 (N_20691,N_17889,N_17509);
and U20692 (N_20692,N_15927,N_16383);
nor U20693 (N_20693,N_18381,N_17956);
nand U20694 (N_20694,N_16357,N_18290);
xor U20695 (N_20695,N_16694,N_15836);
and U20696 (N_20696,N_17473,N_16721);
and U20697 (N_20697,N_16475,N_17753);
nand U20698 (N_20698,N_15668,N_16726);
and U20699 (N_20699,N_15992,N_16831);
xor U20700 (N_20700,N_15993,N_17817);
nor U20701 (N_20701,N_17623,N_18178);
and U20702 (N_20702,N_17548,N_16802);
and U20703 (N_20703,N_18668,N_17651);
or U20704 (N_20704,N_18236,N_16683);
or U20705 (N_20705,N_18538,N_17545);
xnor U20706 (N_20706,N_17828,N_16598);
or U20707 (N_20707,N_16225,N_18611);
nor U20708 (N_20708,N_17927,N_17392);
and U20709 (N_20709,N_15769,N_17967);
xor U20710 (N_20710,N_15962,N_18370);
nor U20711 (N_20711,N_17909,N_16451);
xor U20712 (N_20712,N_15996,N_16696);
or U20713 (N_20713,N_17483,N_18258);
nand U20714 (N_20714,N_17590,N_16103);
nor U20715 (N_20715,N_18087,N_16122);
nand U20716 (N_20716,N_16601,N_15937);
nor U20717 (N_20717,N_16758,N_16292);
nor U20718 (N_20718,N_17399,N_16385);
nor U20719 (N_20719,N_18038,N_17816);
and U20720 (N_20720,N_17659,N_16011);
nand U20721 (N_20721,N_17380,N_16154);
nand U20722 (N_20722,N_18526,N_17350);
or U20723 (N_20723,N_16613,N_17126);
nor U20724 (N_20724,N_16398,N_16452);
nor U20725 (N_20725,N_15807,N_17607);
xor U20726 (N_20726,N_16781,N_17610);
nand U20727 (N_20727,N_17901,N_16677);
or U20728 (N_20728,N_16070,N_16278);
nor U20729 (N_20729,N_18003,N_18010);
nand U20730 (N_20730,N_16590,N_16078);
xnor U20731 (N_20731,N_18590,N_18723);
nor U20732 (N_20732,N_16044,N_15834);
nand U20733 (N_20733,N_15932,N_18689);
xnor U20734 (N_20734,N_16240,N_16241);
nand U20735 (N_20735,N_15810,N_15703);
or U20736 (N_20736,N_16679,N_18474);
nand U20737 (N_20737,N_18504,N_18351);
xor U20738 (N_20738,N_16812,N_18061);
or U20739 (N_20739,N_17937,N_16340);
and U20740 (N_20740,N_15651,N_15881);
nor U20741 (N_20741,N_15981,N_17599);
and U20742 (N_20742,N_17362,N_18184);
nor U20743 (N_20743,N_16864,N_16163);
xnor U20744 (N_20744,N_16310,N_16429);
nand U20745 (N_20745,N_15785,N_16940);
nor U20746 (N_20746,N_18588,N_17153);
or U20747 (N_20747,N_17319,N_17796);
and U20748 (N_20748,N_17240,N_16429);
nand U20749 (N_20749,N_18154,N_17247);
nor U20750 (N_20750,N_17633,N_16440);
nor U20751 (N_20751,N_16061,N_18547);
nand U20752 (N_20752,N_17840,N_16789);
or U20753 (N_20753,N_17687,N_18507);
and U20754 (N_20754,N_17437,N_17260);
or U20755 (N_20755,N_17623,N_18211);
xnor U20756 (N_20756,N_18385,N_15680);
nand U20757 (N_20757,N_15769,N_17043);
nand U20758 (N_20758,N_17652,N_18150);
nor U20759 (N_20759,N_17501,N_16771);
or U20760 (N_20760,N_17644,N_16307);
or U20761 (N_20761,N_16831,N_17672);
nand U20762 (N_20762,N_16020,N_16278);
nand U20763 (N_20763,N_18264,N_17321);
nand U20764 (N_20764,N_15928,N_17609);
and U20765 (N_20765,N_18001,N_17852);
nand U20766 (N_20766,N_16486,N_17566);
nor U20767 (N_20767,N_17392,N_16016);
and U20768 (N_20768,N_16142,N_17133);
or U20769 (N_20769,N_18537,N_16682);
nand U20770 (N_20770,N_15718,N_17949);
xnor U20771 (N_20771,N_18267,N_17599);
nand U20772 (N_20772,N_17531,N_18680);
nand U20773 (N_20773,N_16256,N_16572);
or U20774 (N_20774,N_16398,N_16016);
nand U20775 (N_20775,N_16374,N_16198);
nor U20776 (N_20776,N_17869,N_17730);
nor U20777 (N_20777,N_16327,N_18689);
xor U20778 (N_20778,N_16326,N_15803);
nor U20779 (N_20779,N_18681,N_17462);
and U20780 (N_20780,N_17314,N_16109);
or U20781 (N_20781,N_16855,N_16287);
or U20782 (N_20782,N_16667,N_18013);
xnor U20783 (N_20783,N_18376,N_17462);
nor U20784 (N_20784,N_15802,N_16447);
nor U20785 (N_20785,N_16078,N_15732);
or U20786 (N_20786,N_16182,N_18504);
and U20787 (N_20787,N_16465,N_17809);
and U20788 (N_20788,N_16203,N_17230);
or U20789 (N_20789,N_18587,N_18134);
nand U20790 (N_20790,N_17433,N_16989);
xnor U20791 (N_20791,N_18041,N_17210);
and U20792 (N_20792,N_17633,N_15665);
xor U20793 (N_20793,N_17195,N_15727);
and U20794 (N_20794,N_17973,N_17317);
xor U20795 (N_20795,N_17999,N_15908);
and U20796 (N_20796,N_15958,N_15805);
xnor U20797 (N_20797,N_16726,N_16809);
nand U20798 (N_20798,N_17766,N_18343);
or U20799 (N_20799,N_17270,N_18092);
and U20800 (N_20800,N_16393,N_17096);
and U20801 (N_20801,N_18525,N_17299);
and U20802 (N_20802,N_18578,N_16795);
xnor U20803 (N_20803,N_17109,N_17409);
and U20804 (N_20804,N_17891,N_16058);
or U20805 (N_20805,N_18289,N_18236);
nor U20806 (N_20806,N_16277,N_16932);
or U20807 (N_20807,N_18561,N_16835);
and U20808 (N_20808,N_18691,N_15665);
nand U20809 (N_20809,N_17963,N_15732);
nor U20810 (N_20810,N_17125,N_18275);
nand U20811 (N_20811,N_16471,N_16362);
or U20812 (N_20812,N_17565,N_17146);
and U20813 (N_20813,N_17366,N_17966);
and U20814 (N_20814,N_17851,N_18720);
nor U20815 (N_20815,N_18204,N_16404);
and U20816 (N_20816,N_15767,N_18068);
or U20817 (N_20817,N_16812,N_17612);
or U20818 (N_20818,N_18221,N_16865);
xnor U20819 (N_20819,N_16071,N_16266);
or U20820 (N_20820,N_15904,N_16684);
xnor U20821 (N_20821,N_17984,N_17383);
or U20822 (N_20822,N_16672,N_16357);
and U20823 (N_20823,N_15665,N_16523);
nand U20824 (N_20824,N_17063,N_16664);
or U20825 (N_20825,N_15651,N_16568);
or U20826 (N_20826,N_17446,N_18711);
nand U20827 (N_20827,N_16093,N_17299);
xnor U20828 (N_20828,N_18602,N_16689);
xor U20829 (N_20829,N_17700,N_16077);
and U20830 (N_20830,N_17161,N_18560);
nor U20831 (N_20831,N_17845,N_17857);
xor U20832 (N_20832,N_18217,N_18546);
nand U20833 (N_20833,N_18085,N_17174);
nand U20834 (N_20834,N_16406,N_17727);
nor U20835 (N_20835,N_17738,N_16209);
xor U20836 (N_20836,N_18157,N_16342);
and U20837 (N_20837,N_18175,N_16712);
nand U20838 (N_20838,N_17163,N_17385);
nor U20839 (N_20839,N_17891,N_17699);
xnor U20840 (N_20840,N_16864,N_16481);
nand U20841 (N_20841,N_16470,N_17224);
nand U20842 (N_20842,N_18065,N_16383);
nor U20843 (N_20843,N_16644,N_16443);
xor U20844 (N_20844,N_17069,N_17701);
nor U20845 (N_20845,N_17908,N_18510);
nand U20846 (N_20846,N_17981,N_17472);
xnor U20847 (N_20847,N_17541,N_18085);
nand U20848 (N_20848,N_17107,N_18262);
or U20849 (N_20849,N_15989,N_17781);
and U20850 (N_20850,N_15954,N_16606);
nor U20851 (N_20851,N_17352,N_17965);
nor U20852 (N_20852,N_16135,N_17064);
xnor U20853 (N_20853,N_17758,N_18442);
xnor U20854 (N_20854,N_18037,N_16872);
nand U20855 (N_20855,N_17679,N_16877);
xor U20856 (N_20856,N_17679,N_16077);
xor U20857 (N_20857,N_17822,N_16843);
xor U20858 (N_20858,N_17603,N_16355);
xor U20859 (N_20859,N_17747,N_16621);
and U20860 (N_20860,N_16985,N_17379);
and U20861 (N_20861,N_17358,N_17627);
or U20862 (N_20862,N_16938,N_18732);
nand U20863 (N_20863,N_17832,N_17041);
or U20864 (N_20864,N_17249,N_16466);
nand U20865 (N_20865,N_17009,N_15653);
and U20866 (N_20866,N_15678,N_16321);
and U20867 (N_20867,N_16795,N_17620);
nand U20868 (N_20868,N_17270,N_18167);
and U20869 (N_20869,N_16428,N_16418);
and U20870 (N_20870,N_16785,N_16693);
or U20871 (N_20871,N_18608,N_17503);
nor U20872 (N_20872,N_18560,N_18075);
nor U20873 (N_20873,N_15644,N_16200);
or U20874 (N_20874,N_17998,N_17540);
and U20875 (N_20875,N_17658,N_18413);
xor U20876 (N_20876,N_16692,N_15711);
nand U20877 (N_20877,N_18363,N_16299);
and U20878 (N_20878,N_18554,N_17583);
or U20879 (N_20879,N_18481,N_15629);
or U20880 (N_20880,N_15817,N_16771);
or U20881 (N_20881,N_17726,N_16884);
or U20882 (N_20882,N_17035,N_16624);
or U20883 (N_20883,N_18387,N_18285);
xnor U20884 (N_20884,N_16626,N_16542);
nor U20885 (N_20885,N_16050,N_17438);
or U20886 (N_20886,N_18055,N_17721);
nand U20887 (N_20887,N_15907,N_16872);
and U20888 (N_20888,N_16889,N_18067);
and U20889 (N_20889,N_16906,N_18588);
or U20890 (N_20890,N_18330,N_16321);
xnor U20891 (N_20891,N_18386,N_16819);
and U20892 (N_20892,N_15959,N_16327);
or U20893 (N_20893,N_17106,N_16123);
xnor U20894 (N_20894,N_15932,N_17601);
or U20895 (N_20895,N_16024,N_16358);
and U20896 (N_20896,N_18602,N_18084);
xor U20897 (N_20897,N_16178,N_17979);
xnor U20898 (N_20898,N_16761,N_16240);
nand U20899 (N_20899,N_18633,N_18133);
and U20900 (N_20900,N_18239,N_16217);
xor U20901 (N_20901,N_15983,N_18404);
xor U20902 (N_20902,N_15644,N_17477);
or U20903 (N_20903,N_18112,N_18295);
or U20904 (N_20904,N_16214,N_18069);
xor U20905 (N_20905,N_17207,N_16646);
and U20906 (N_20906,N_17287,N_15717);
and U20907 (N_20907,N_15955,N_15778);
xnor U20908 (N_20908,N_15807,N_17087);
nand U20909 (N_20909,N_15961,N_15683);
nand U20910 (N_20910,N_16956,N_17337);
nand U20911 (N_20911,N_17456,N_18730);
and U20912 (N_20912,N_17019,N_16265);
xor U20913 (N_20913,N_18139,N_17464);
nor U20914 (N_20914,N_17104,N_18615);
and U20915 (N_20915,N_17895,N_17957);
or U20916 (N_20916,N_17755,N_15820);
nand U20917 (N_20917,N_17002,N_15843);
or U20918 (N_20918,N_17140,N_17089);
nand U20919 (N_20919,N_18326,N_18371);
or U20920 (N_20920,N_16878,N_16599);
nor U20921 (N_20921,N_16702,N_17702);
and U20922 (N_20922,N_17405,N_18434);
or U20923 (N_20923,N_15837,N_16273);
and U20924 (N_20924,N_15851,N_16945);
nor U20925 (N_20925,N_17516,N_15958);
xnor U20926 (N_20926,N_17019,N_17136);
and U20927 (N_20927,N_16900,N_16111);
or U20928 (N_20928,N_16561,N_16098);
nand U20929 (N_20929,N_17479,N_17886);
or U20930 (N_20930,N_17879,N_17721);
nor U20931 (N_20931,N_17099,N_18117);
nor U20932 (N_20932,N_17636,N_17001);
or U20933 (N_20933,N_16182,N_17466);
xnor U20934 (N_20934,N_15821,N_17204);
nand U20935 (N_20935,N_16853,N_16247);
xnor U20936 (N_20936,N_16344,N_18583);
xnor U20937 (N_20937,N_18144,N_18293);
nor U20938 (N_20938,N_15767,N_18210);
nand U20939 (N_20939,N_18733,N_16368);
and U20940 (N_20940,N_17850,N_18269);
xor U20941 (N_20941,N_16680,N_18605);
nand U20942 (N_20942,N_16499,N_17274);
and U20943 (N_20943,N_16078,N_15980);
xnor U20944 (N_20944,N_18342,N_16983);
or U20945 (N_20945,N_18163,N_16774);
or U20946 (N_20946,N_17337,N_16039);
nor U20947 (N_20947,N_16745,N_17729);
and U20948 (N_20948,N_17392,N_17258);
or U20949 (N_20949,N_16187,N_18171);
or U20950 (N_20950,N_17398,N_15743);
nor U20951 (N_20951,N_15995,N_17833);
or U20952 (N_20952,N_18381,N_16440);
nor U20953 (N_20953,N_18482,N_16450);
nor U20954 (N_20954,N_15680,N_18113);
and U20955 (N_20955,N_17542,N_18708);
nand U20956 (N_20956,N_16167,N_17877);
nand U20957 (N_20957,N_18367,N_17529);
or U20958 (N_20958,N_16702,N_16865);
and U20959 (N_20959,N_16327,N_17394);
xnor U20960 (N_20960,N_17986,N_17155);
nor U20961 (N_20961,N_17240,N_17994);
xor U20962 (N_20962,N_16610,N_15665);
or U20963 (N_20963,N_15765,N_15722);
and U20964 (N_20964,N_15765,N_16246);
nor U20965 (N_20965,N_15859,N_17212);
nand U20966 (N_20966,N_15671,N_15646);
nor U20967 (N_20967,N_17203,N_17720);
nor U20968 (N_20968,N_15874,N_16827);
nor U20969 (N_20969,N_16526,N_16345);
xnor U20970 (N_20970,N_17808,N_17976);
and U20971 (N_20971,N_16219,N_17792);
and U20972 (N_20972,N_17959,N_16366);
or U20973 (N_20973,N_18124,N_17425);
or U20974 (N_20974,N_16478,N_16237);
nand U20975 (N_20975,N_17265,N_18005);
nor U20976 (N_20976,N_17321,N_18488);
nor U20977 (N_20977,N_18597,N_17396);
or U20978 (N_20978,N_17162,N_15880);
nand U20979 (N_20979,N_15803,N_16530);
or U20980 (N_20980,N_17803,N_17532);
or U20981 (N_20981,N_16169,N_17737);
nand U20982 (N_20982,N_18011,N_17595);
and U20983 (N_20983,N_15843,N_16022);
or U20984 (N_20984,N_15683,N_16174);
nand U20985 (N_20985,N_16584,N_17249);
nor U20986 (N_20986,N_18238,N_17657);
nand U20987 (N_20987,N_16639,N_17012);
nor U20988 (N_20988,N_17580,N_16977);
xor U20989 (N_20989,N_15770,N_16845);
nor U20990 (N_20990,N_17287,N_16641);
nor U20991 (N_20991,N_16811,N_15724);
nand U20992 (N_20992,N_18098,N_18198);
nor U20993 (N_20993,N_18594,N_17997);
xnor U20994 (N_20994,N_16540,N_16458);
nor U20995 (N_20995,N_18384,N_16383);
nor U20996 (N_20996,N_17132,N_16541);
nand U20997 (N_20997,N_18079,N_18242);
or U20998 (N_20998,N_17525,N_17215);
and U20999 (N_20999,N_17289,N_18579);
and U21000 (N_21000,N_16023,N_15778);
or U21001 (N_21001,N_18004,N_16574);
and U21002 (N_21002,N_15664,N_16305);
xor U21003 (N_21003,N_18467,N_17131);
or U21004 (N_21004,N_18390,N_15846);
xor U21005 (N_21005,N_17876,N_15870);
nor U21006 (N_21006,N_18577,N_16299);
or U21007 (N_21007,N_17145,N_15943);
or U21008 (N_21008,N_18026,N_16391);
or U21009 (N_21009,N_18511,N_17289);
and U21010 (N_21010,N_17728,N_17067);
xnor U21011 (N_21011,N_18625,N_17831);
nor U21012 (N_21012,N_17582,N_15656);
and U21013 (N_21013,N_15923,N_17317);
nor U21014 (N_21014,N_18441,N_18742);
nand U21015 (N_21015,N_16739,N_17249);
and U21016 (N_21016,N_16757,N_16142);
nand U21017 (N_21017,N_18069,N_15946);
xor U21018 (N_21018,N_16720,N_16948);
or U21019 (N_21019,N_16123,N_16514);
nor U21020 (N_21020,N_17463,N_18197);
nor U21021 (N_21021,N_16722,N_16554);
nand U21022 (N_21022,N_17583,N_18623);
nand U21023 (N_21023,N_16487,N_18205);
and U21024 (N_21024,N_17034,N_17186);
nand U21025 (N_21025,N_17641,N_18566);
or U21026 (N_21026,N_15756,N_16790);
nand U21027 (N_21027,N_17456,N_16803);
and U21028 (N_21028,N_16667,N_18477);
and U21029 (N_21029,N_17196,N_16200);
nand U21030 (N_21030,N_16154,N_16964);
nand U21031 (N_21031,N_16536,N_18491);
nand U21032 (N_21032,N_15784,N_17162);
xor U21033 (N_21033,N_16492,N_15656);
nor U21034 (N_21034,N_17548,N_16002);
nor U21035 (N_21035,N_17514,N_15910);
xnor U21036 (N_21036,N_18147,N_17358);
and U21037 (N_21037,N_17385,N_16355);
nor U21038 (N_21038,N_16036,N_16265);
and U21039 (N_21039,N_16002,N_17224);
nor U21040 (N_21040,N_17256,N_17088);
nor U21041 (N_21041,N_18083,N_18237);
and U21042 (N_21042,N_18722,N_17002);
or U21043 (N_21043,N_17461,N_16132);
nand U21044 (N_21044,N_16443,N_15647);
and U21045 (N_21045,N_17750,N_18068);
nand U21046 (N_21046,N_16904,N_17844);
nor U21047 (N_21047,N_18165,N_15991);
xnor U21048 (N_21048,N_15805,N_16246);
nor U21049 (N_21049,N_18445,N_17467);
xor U21050 (N_21050,N_17864,N_15844);
xnor U21051 (N_21051,N_16131,N_18671);
xnor U21052 (N_21052,N_18602,N_17224);
or U21053 (N_21053,N_18227,N_17321);
nand U21054 (N_21054,N_17585,N_18376);
nor U21055 (N_21055,N_17652,N_16000);
nand U21056 (N_21056,N_18071,N_18418);
and U21057 (N_21057,N_17828,N_17988);
nand U21058 (N_21058,N_16210,N_17850);
nor U21059 (N_21059,N_15761,N_17094);
xnor U21060 (N_21060,N_16544,N_18406);
xor U21061 (N_21061,N_17258,N_18616);
xor U21062 (N_21062,N_18561,N_17430);
or U21063 (N_21063,N_18301,N_15764);
nor U21064 (N_21064,N_17115,N_17067);
xor U21065 (N_21065,N_18173,N_17630);
or U21066 (N_21066,N_17646,N_17682);
nand U21067 (N_21067,N_15911,N_17469);
and U21068 (N_21068,N_16860,N_16483);
and U21069 (N_21069,N_16995,N_17552);
nand U21070 (N_21070,N_17472,N_18502);
and U21071 (N_21071,N_17437,N_15875);
and U21072 (N_21072,N_17887,N_17352);
nand U21073 (N_21073,N_18604,N_16863);
or U21074 (N_21074,N_16882,N_17993);
and U21075 (N_21075,N_18339,N_15764);
and U21076 (N_21076,N_16576,N_15682);
or U21077 (N_21077,N_18677,N_16585);
nand U21078 (N_21078,N_18148,N_17012);
nor U21079 (N_21079,N_16189,N_16837);
nor U21080 (N_21080,N_16389,N_16477);
nand U21081 (N_21081,N_17324,N_17207);
xnor U21082 (N_21082,N_16079,N_17860);
nand U21083 (N_21083,N_17501,N_18329);
xnor U21084 (N_21084,N_17980,N_16861);
or U21085 (N_21085,N_17355,N_17072);
xor U21086 (N_21086,N_16966,N_17968);
nand U21087 (N_21087,N_17346,N_18291);
and U21088 (N_21088,N_16057,N_17157);
or U21089 (N_21089,N_18192,N_18597);
nor U21090 (N_21090,N_18140,N_18594);
nand U21091 (N_21091,N_18477,N_18181);
xor U21092 (N_21092,N_18642,N_17546);
nor U21093 (N_21093,N_17195,N_17855);
nor U21094 (N_21094,N_17358,N_17851);
nor U21095 (N_21095,N_15857,N_18238);
and U21096 (N_21096,N_16712,N_17158);
nor U21097 (N_21097,N_16942,N_18135);
and U21098 (N_21098,N_17615,N_17594);
nand U21099 (N_21099,N_15984,N_17613);
or U21100 (N_21100,N_17953,N_16060);
xor U21101 (N_21101,N_17443,N_15938);
nand U21102 (N_21102,N_17612,N_17005);
xnor U21103 (N_21103,N_15661,N_17896);
or U21104 (N_21104,N_17412,N_18074);
or U21105 (N_21105,N_17996,N_17590);
and U21106 (N_21106,N_16299,N_16011);
nor U21107 (N_21107,N_17734,N_17758);
xor U21108 (N_21108,N_17609,N_16064);
or U21109 (N_21109,N_17705,N_17200);
and U21110 (N_21110,N_17441,N_16853);
xnor U21111 (N_21111,N_18492,N_16681);
xnor U21112 (N_21112,N_16861,N_17859);
nor U21113 (N_21113,N_18313,N_18103);
or U21114 (N_21114,N_17948,N_16160);
or U21115 (N_21115,N_17495,N_17371);
nor U21116 (N_21116,N_15695,N_15999);
or U21117 (N_21117,N_17180,N_17072);
xnor U21118 (N_21118,N_17300,N_16703);
nand U21119 (N_21119,N_17701,N_18616);
nand U21120 (N_21120,N_17700,N_17299);
nand U21121 (N_21121,N_16457,N_18642);
and U21122 (N_21122,N_15776,N_18044);
xor U21123 (N_21123,N_16768,N_18576);
nor U21124 (N_21124,N_17455,N_16882);
or U21125 (N_21125,N_15675,N_17457);
or U21126 (N_21126,N_17676,N_17708);
nor U21127 (N_21127,N_16375,N_15755);
or U21128 (N_21128,N_15832,N_17134);
nor U21129 (N_21129,N_15880,N_18330);
or U21130 (N_21130,N_17794,N_16493);
nor U21131 (N_21131,N_16410,N_15992);
nor U21132 (N_21132,N_17389,N_16654);
nand U21133 (N_21133,N_16418,N_16971);
xnor U21134 (N_21134,N_16690,N_16643);
nor U21135 (N_21135,N_16962,N_16504);
nand U21136 (N_21136,N_17799,N_17296);
and U21137 (N_21137,N_15640,N_15876);
or U21138 (N_21138,N_18124,N_15828);
nand U21139 (N_21139,N_15758,N_15835);
or U21140 (N_21140,N_18056,N_15650);
and U21141 (N_21141,N_18355,N_17315);
or U21142 (N_21142,N_17288,N_16711);
nor U21143 (N_21143,N_18107,N_17115);
nand U21144 (N_21144,N_15956,N_16193);
and U21145 (N_21145,N_17476,N_15877);
nor U21146 (N_21146,N_16980,N_16266);
nor U21147 (N_21147,N_16886,N_16092);
nand U21148 (N_21148,N_16438,N_17901);
xnor U21149 (N_21149,N_18034,N_17466);
nor U21150 (N_21150,N_18168,N_17787);
xor U21151 (N_21151,N_15856,N_17637);
and U21152 (N_21152,N_17826,N_16695);
nor U21153 (N_21153,N_16632,N_16043);
nor U21154 (N_21154,N_18742,N_15889);
nor U21155 (N_21155,N_16417,N_16255);
or U21156 (N_21156,N_16266,N_17716);
nand U21157 (N_21157,N_15852,N_17206);
nor U21158 (N_21158,N_15793,N_17740);
or U21159 (N_21159,N_16397,N_16052);
nor U21160 (N_21160,N_18026,N_17840);
or U21161 (N_21161,N_17337,N_16470);
and U21162 (N_21162,N_17172,N_16166);
and U21163 (N_21163,N_17141,N_16431);
nor U21164 (N_21164,N_15729,N_16410);
nand U21165 (N_21165,N_17297,N_16332);
nor U21166 (N_21166,N_17335,N_18142);
or U21167 (N_21167,N_18335,N_16522);
nor U21168 (N_21168,N_16606,N_18138);
or U21169 (N_21169,N_18348,N_15916);
nor U21170 (N_21170,N_17855,N_15906);
and U21171 (N_21171,N_17871,N_18165);
or U21172 (N_21172,N_16246,N_18393);
and U21173 (N_21173,N_16297,N_16184);
and U21174 (N_21174,N_17653,N_18572);
or U21175 (N_21175,N_16004,N_16352);
nand U21176 (N_21176,N_18513,N_17679);
nor U21177 (N_21177,N_18116,N_16838);
or U21178 (N_21178,N_17687,N_17208);
nor U21179 (N_21179,N_15729,N_18204);
nand U21180 (N_21180,N_17008,N_17019);
nor U21181 (N_21181,N_17411,N_15707);
nand U21182 (N_21182,N_15948,N_17434);
nor U21183 (N_21183,N_15700,N_17603);
nor U21184 (N_21184,N_17763,N_17856);
or U21185 (N_21185,N_15658,N_18630);
nand U21186 (N_21186,N_16759,N_16887);
xor U21187 (N_21187,N_17605,N_18427);
or U21188 (N_21188,N_16539,N_16338);
nor U21189 (N_21189,N_18353,N_18741);
nand U21190 (N_21190,N_17313,N_18306);
nor U21191 (N_21191,N_17855,N_15689);
xnor U21192 (N_21192,N_17577,N_18144);
xor U21193 (N_21193,N_18631,N_17485);
xnor U21194 (N_21194,N_17842,N_18007);
nand U21195 (N_21195,N_18567,N_18219);
nor U21196 (N_21196,N_18222,N_16418);
nor U21197 (N_21197,N_16192,N_18572);
nor U21198 (N_21198,N_16112,N_15647);
nand U21199 (N_21199,N_17928,N_16120);
and U21200 (N_21200,N_17781,N_16847);
nor U21201 (N_21201,N_17431,N_17180);
nand U21202 (N_21202,N_16505,N_18706);
or U21203 (N_21203,N_17954,N_16066);
nand U21204 (N_21204,N_15901,N_16703);
nor U21205 (N_21205,N_17094,N_16199);
and U21206 (N_21206,N_17747,N_17275);
and U21207 (N_21207,N_15748,N_17364);
or U21208 (N_21208,N_16452,N_18538);
and U21209 (N_21209,N_16807,N_18220);
xnor U21210 (N_21210,N_16060,N_16153);
and U21211 (N_21211,N_18608,N_18552);
and U21212 (N_21212,N_18514,N_17599);
nor U21213 (N_21213,N_15941,N_18174);
nor U21214 (N_21214,N_15673,N_17378);
xnor U21215 (N_21215,N_15746,N_16125);
nor U21216 (N_21216,N_16137,N_18312);
and U21217 (N_21217,N_15952,N_17415);
nor U21218 (N_21218,N_18508,N_18634);
nor U21219 (N_21219,N_18467,N_17431);
xor U21220 (N_21220,N_15803,N_18347);
or U21221 (N_21221,N_16327,N_16835);
or U21222 (N_21222,N_15959,N_18625);
or U21223 (N_21223,N_18616,N_16460);
nand U21224 (N_21224,N_15872,N_17372);
or U21225 (N_21225,N_18377,N_18542);
xor U21226 (N_21226,N_17569,N_18295);
or U21227 (N_21227,N_16126,N_16665);
xor U21228 (N_21228,N_18379,N_15741);
xor U21229 (N_21229,N_16868,N_16271);
and U21230 (N_21230,N_16749,N_17001);
and U21231 (N_21231,N_18514,N_16400);
or U21232 (N_21232,N_17264,N_16512);
nand U21233 (N_21233,N_17777,N_18730);
xor U21234 (N_21234,N_18546,N_16740);
nand U21235 (N_21235,N_16366,N_15921);
nand U21236 (N_21236,N_16782,N_18389);
nor U21237 (N_21237,N_17030,N_16297);
nand U21238 (N_21238,N_16919,N_16008);
and U21239 (N_21239,N_15723,N_17387);
nand U21240 (N_21240,N_18121,N_15723);
and U21241 (N_21241,N_17141,N_18235);
or U21242 (N_21242,N_17158,N_16175);
nor U21243 (N_21243,N_16024,N_16738);
xor U21244 (N_21244,N_16248,N_16384);
xnor U21245 (N_21245,N_16394,N_17894);
and U21246 (N_21246,N_16420,N_18294);
xnor U21247 (N_21247,N_15989,N_17824);
xor U21248 (N_21248,N_16481,N_16048);
or U21249 (N_21249,N_16962,N_17266);
nor U21250 (N_21250,N_15692,N_16598);
nor U21251 (N_21251,N_17167,N_17692);
or U21252 (N_21252,N_18398,N_18126);
nand U21253 (N_21253,N_15967,N_16221);
nor U21254 (N_21254,N_16597,N_17442);
or U21255 (N_21255,N_18370,N_15661);
nand U21256 (N_21256,N_15661,N_17061);
xor U21257 (N_21257,N_16100,N_15647);
and U21258 (N_21258,N_16679,N_17313);
nor U21259 (N_21259,N_16157,N_18711);
xor U21260 (N_21260,N_16688,N_16921);
xnor U21261 (N_21261,N_16411,N_16449);
or U21262 (N_21262,N_18538,N_18130);
and U21263 (N_21263,N_17506,N_18178);
or U21264 (N_21264,N_18178,N_17484);
xor U21265 (N_21265,N_16017,N_16322);
and U21266 (N_21266,N_16628,N_17244);
or U21267 (N_21267,N_18202,N_17436);
xnor U21268 (N_21268,N_16546,N_17723);
nand U21269 (N_21269,N_18582,N_18309);
nand U21270 (N_21270,N_16951,N_17571);
xor U21271 (N_21271,N_16009,N_17629);
or U21272 (N_21272,N_16921,N_18397);
nand U21273 (N_21273,N_16776,N_16116);
nand U21274 (N_21274,N_18481,N_17171);
or U21275 (N_21275,N_17423,N_17797);
and U21276 (N_21276,N_17979,N_15745);
xnor U21277 (N_21277,N_18698,N_17592);
and U21278 (N_21278,N_17521,N_18050);
and U21279 (N_21279,N_16178,N_15723);
nand U21280 (N_21280,N_18741,N_16524);
or U21281 (N_21281,N_17382,N_18173);
nand U21282 (N_21282,N_16012,N_16502);
xor U21283 (N_21283,N_18047,N_16226);
xnor U21284 (N_21284,N_17287,N_16413);
nand U21285 (N_21285,N_17511,N_15975);
or U21286 (N_21286,N_17384,N_16363);
or U21287 (N_21287,N_15878,N_16626);
and U21288 (N_21288,N_16965,N_18011);
nand U21289 (N_21289,N_18172,N_17843);
nand U21290 (N_21290,N_17437,N_18076);
nor U21291 (N_21291,N_16426,N_17154);
and U21292 (N_21292,N_17986,N_16792);
xor U21293 (N_21293,N_17348,N_18650);
and U21294 (N_21294,N_17212,N_18402);
nand U21295 (N_21295,N_18491,N_16103);
nand U21296 (N_21296,N_17147,N_17764);
nor U21297 (N_21297,N_18240,N_16584);
xor U21298 (N_21298,N_16903,N_15768);
xor U21299 (N_21299,N_18395,N_16044);
xnor U21300 (N_21300,N_17665,N_17572);
nor U21301 (N_21301,N_16965,N_17597);
or U21302 (N_21302,N_18019,N_18128);
and U21303 (N_21303,N_15702,N_18333);
xor U21304 (N_21304,N_17723,N_16806);
nor U21305 (N_21305,N_16012,N_17115);
or U21306 (N_21306,N_17770,N_16633);
xor U21307 (N_21307,N_16798,N_18673);
xor U21308 (N_21308,N_18260,N_16169);
and U21309 (N_21309,N_18654,N_17322);
and U21310 (N_21310,N_17531,N_15860);
nand U21311 (N_21311,N_17681,N_16015);
or U21312 (N_21312,N_18098,N_17621);
or U21313 (N_21313,N_15877,N_15963);
or U21314 (N_21314,N_18704,N_17284);
and U21315 (N_21315,N_16840,N_16666);
and U21316 (N_21316,N_16210,N_16153);
and U21317 (N_21317,N_15761,N_15829);
nor U21318 (N_21318,N_17841,N_16258);
nand U21319 (N_21319,N_16372,N_17038);
or U21320 (N_21320,N_18121,N_16206);
and U21321 (N_21321,N_18716,N_17138);
nand U21322 (N_21322,N_18144,N_17017);
and U21323 (N_21323,N_16308,N_18555);
nand U21324 (N_21324,N_16201,N_17374);
and U21325 (N_21325,N_15742,N_18583);
nor U21326 (N_21326,N_16460,N_16351);
xnor U21327 (N_21327,N_15642,N_17083);
nand U21328 (N_21328,N_18579,N_15975);
nor U21329 (N_21329,N_17612,N_18519);
and U21330 (N_21330,N_18728,N_18092);
xor U21331 (N_21331,N_17910,N_15922);
xnor U21332 (N_21332,N_15754,N_17718);
and U21333 (N_21333,N_16953,N_17367);
and U21334 (N_21334,N_16120,N_17596);
xnor U21335 (N_21335,N_15721,N_16594);
nor U21336 (N_21336,N_18526,N_18496);
or U21337 (N_21337,N_18331,N_17870);
or U21338 (N_21338,N_17955,N_18063);
or U21339 (N_21339,N_17180,N_17374);
or U21340 (N_21340,N_16250,N_16855);
or U21341 (N_21341,N_15989,N_18748);
or U21342 (N_21342,N_16500,N_17222);
or U21343 (N_21343,N_17384,N_16168);
and U21344 (N_21344,N_17406,N_17588);
xor U21345 (N_21345,N_16893,N_17012);
xor U21346 (N_21346,N_16170,N_18404);
nand U21347 (N_21347,N_16391,N_18540);
and U21348 (N_21348,N_16664,N_17905);
nand U21349 (N_21349,N_17273,N_18477);
and U21350 (N_21350,N_17845,N_18667);
and U21351 (N_21351,N_18502,N_16084);
nor U21352 (N_21352,N_17248,N_17673);
and U21353 (N_21353,N_18503,N_17865);
and U21354 (N_21354,N_18310,N_17745);
or U21355 (N_21355,N_18133,N_17724);
nand U21356 (N_21356,N_18235,N_18187);
xor U21357 (N_21357,N_15937,N_18224);
and U21358 (N_21358,N_16135,N_16294);
nor U21359 (N_21359,N_17428,N_18639);
and U21360 (N_21360,N_16641,N_17355);
or U21361 (N_21361,N_18232,N_16303);
xor U21362 (N_21362,N_18007,N_16324);
nand U21363 (N_21363,N_18370,N_17008);
nor U21364 (N_21364,N_16719,N_18322);
or U21365 (N_21365,N_17680,N_18400);
and U21366 (N_21366,N_17751,N_18625);
nor U21367 (N_21367,N_17889,N_15680);
and U21368 (N_21368,N_16137,N_18522);
or U21369 (N_21369,N_18018,N_17545);
or U21370 (N_21370,N_16768,N_17801);
and U21371 (N_21371,N_15949,N_17313);
nand U21372 (N_21372,N_17998,N_15681);
and U21373 (N_21373,N_16454,N_16140);
xnor U21374 (N_21374,N_16125,N_18325);
and U21375 (N_21375,N_16074,N_17477);
nand U21376 (N_21376,N_18509,N_16677);
xnor U21377 (N_21377,N_16977,N_17452);
nand U21378 (N_21378,N_18444,N_18602);
nor U21379 (N_21379,N_18103,N_17954);
nor U21380 (N_21380,N_18459,N_17789);
xor U21381 (N_21381,N_16239,N_18042);
and U21382 (N_21382,N_16812,N_15842);
nor U21383 (N_21383,N_17520,N_16907);
xor U21384 (N_21384,N_17978,N_18443);
xnor U21385 (N_21385,N_18722,N_16393);
nand U21386 (N_21386,N_15980,N_17413);
xnor U21387 (N_21387,N_16695,N_17769);
nor U21388 (N_21388,N_17893,N_18720);
and U21389 (N_21389,N_17514,N_17596);
xor U21390 (N_21390,N_16863,N_18045);
xor U21391 (N_21391,N_18613,N_17460);
or U21392 (N_21392,N_16915,N_17490);
nand U21393 (N_21393,N_16196,N_16638);
nor U21394 (N_21394,N_18071,N_17359);
xor U21395 (N_21395,N_15893,N_17221);
nand U21396 (N_21396,N_16732,N_18353);
nor U21397 (N_21397,N_16628,N_18052);
nor U21398 (N_21398,N_15940,N_16704);
nand U21399 (N_21399,N_16135,N_18705);
nor U21400 (N_21400,N_16183,N_16858);
and U21401 (N_21401,N_17744,N_16441);
xor U21402 (N_21402,N_17587,N_17417);
nor U21403 (N_21403,N_15868,N_16752);
nand U21404 (N_21404,N_17867,N_18097);
and U21405 (N_21405,N_18588,N_15836);
or U21406 (N_21406,N_16646,N_16020);
and U21407 (N_21407,N_16558,N_15684);
nor U21408 (N_21408,N_18119,N_17301);
or U21409 (N_21409,N_16868,N_16491);
xnor U21410 (N_21410,N_17586,N_17605);
xnor U21411 (N_21411,N_16290,N_16085);
xnor U21412 (N_21412,N_16043,N_16291);
and U21413 (N_21413,N_18361,N_18628);
or U21414 (N_21414,N_17671,N_16304);
and U21415 (N_21415,N_15626,N_16562);
and U21416 (N_21416,N_16303,N_16848);
xor U21417 (N_21417,N_17473,N_16414);
nor U21418 (N_21418,N_17079,N_17735);
xor U21419 (N_21419,N_17962,N_15984);
and U21420 (N_21420,N_16992,N_16725);
xnor U21421 (N_21421,N_17968,N_16301);
nor U21422 (N_21422,N_16054,N_17899);
and U21423 (N_21423,N_18356,N_16148);
or U21424 (N_21424,N_18247,N_15636);
nand U21425 (N_21425,N_15923,N_16939);
nand U21426 (N_21426,N_17057,N_17076);
xnor U21427 (N_21427,N_17860,N_18557);
and U21428 (N_21428,N_16018,N_17188);
nor U21429 (N_21429,N_17996,N_17501);
xnor U21430 (N_21430,N_16593,N_18150);
or U21431 (N_21431,N_15692,N_16056);
nand U21432 (N_21432,N_18334,N_16918);
xor U21433 (N_21433,N_18125,N_18316);
nor U21434 (N_21434,N_15671,N_18110);
nor U21435 (N_21435,N_18587,N_16301);
nor U21436 (N_21436,N_18356,N_18157);
nand U21437 (N_21437,N_17923,N_18206);
and U21438 (N_21438,N_15652,N_18292);
nor U21439 (N_21439,N_15964,N_18201);
and U21440 (N_21440,N_17262,N_17901);
or U21441 (N_21441,N_16486,N_17191);
nand U21442 (N_21442,N_15812,N_18237);
and U21443 (N_21443,N_18723,N_15671);
nand U21444 (N_21444,N_17846,N_18557);
and U21445 (N_21445,N_18164,N_18576);
nand U21446 (N_21446,N_17662,N_17053);
and U21447 (N_21447,N_18368,N_17196);
xnor U21448 (N_21448,N_16012,N_15707);
xor U21449 (N_21449,N_16937,N_16395);
nor U21450 (N_21450,N_15931,N_18251);
xnor U21451 (N_21451,N_18727,N_17463);
nor U21452 (N_21452,N_16137,N_17967);
nor U21453 (N_21453,N_17682,N_18289);
nand U21454 (N_21454,N_15763,N_18568);
nor U21455 (N_21455,N_15775,N_15640);
or U21456 (N_21456,N_18471,N_16264);
and U21457 (N_21457,N_18192,N_18075);
or U21458 (N_21458,N_17007,N_18509);
nand U21459 (N_21459,N_17480,N_16005);
nand U21460 (N_21460,N_15700,N_18700);
and U21461 (N_21461,N_16361,N_18603);
and U21462 (N_21462,N_18081,N_17242);
nor U21463 (N_21463,N_18645,N_15933);
and U21464 (N_21464,N_16984,N_18181);
nor U21465 (N_21465,N_18402,N_18654);
nor U21466 (N_21466,N_15691,N_18473);
and U21467 (N_21467,N_18657,N_17630);
or U21468 (N_21468,N_17634,N_16072);
or U21469 (N_21469,N_18101,N_16278);
or U21470 (N_21470,N_17089,N_16683);
xor U21471 (N_21471,N_18413,N_16127);
or U21472 (N_21472,N_16436,N_17043);
or U21473 (N_21473,N_16647,N_16353);
xnor U21474 (N_21474,N_17254,N_17373);
nand U21475 (N_21475,N_18174,N_18090);
or U21476 (N_21476,N_17459,N_15663);
or U21477 (N_21477,N_15809,N_18586);
and U21478 (N_21478,N_18014,N_17987);
xnor U21479 (N_21479,N_16624,N_15910);
nand U21480 (N_21480,N_16299,N_17106);
or U21481 (N_21481,N_16337,N_17176);
nand U21482 (N_21482,N_17762,N_16892);
xnor U21483 (N_21483,N_17966,N_17731);
nand U21484 (N_21484,N_16334,N_17986);
or U21485 (N_21485,N_16901,N_16088);
nand U21486 (N_21486,N_17512,N_17809);
and U21487 (N_21487,N_15756,N_17332);
xor U21488 (N_21488,N_17529,N_17720);
nor U21489 (N_21489,N_16080,N_17390);
and U21490 (N_21490,N_17507,N_16540);
xor U21491 (N_21491,N_17580,N_17307);
nor U21492 (N_21492,N_17244,N_16560);
and U21493 (N_21493,N_17130,N_17095);
xor U21494 (N_21494,N_17413,N_18513);
xnor U21495 (N_21495,N_16388,N_17699);
nand U21496 (N_21496,N_16286,N_16434);
xnor U21497 (N_21497,N_18625,N_17260);
nand U21498 (N_21498,N_17318,N_16294);
xnor U21499 (N_21499,N_15766,N_17189);
nand U21500 (N_21500,N_17671,N_18638);
xnor U21501 (N_21501,N_17731,N_17893);
or U21502 (N_21502,N_16070,N_18146);
and U21503 (N_21503,N_17788,N_16828);
nor U21504 (N_21504,N_16029,N_15740);
nor U21505 (N_21505,N_16281,N_17755);
or U21506 (N_21506,N_17438,N_17611);
nor U21507 (N_21507,N_18663,N_16543);
or U21508 (N_21508,N_18580,N_17037);
nor U21509 (N_21509,N_17105,N_18585);
xnor U21510 (N_21510,N_16668,N_17088);
xnor U21511 (N_21511,N_17365,N_17283);
xor U21512 (N_21512,N_18190,N_16449);
xnor U21513 (N_21513,N_16456,N_18622);
and U21514 (N_21514,N_18165,N_16954);
nor U21515 (N_21515,N_17081,N_18296);
nand U21516 (N_21516,N_16713,N_17136);
nor U21517 (N_21517,N_17579,N_16004);
xnor U21518 (N_21518,N_16995,N_18311);
and U21519 (N_21519,N_17086,N_16382);
nor U21520 (N_21520,N_18538,N_16898);
and U21521 (N_21521,N_16646,N_16286);
nand U21522 (N_21522,N_17460,N_16673);
nand U21523 (N_21523,N_16875,N_16026);
xnor U21524 (N_21524,N_16698,N_15736);
or U21525 (N_21525,N_18419,N_16997);
nand U21526 (N_21526,N_15959,N_17604);
xnor U21527 (N_21527,N_18575,N_17729);
xnor U21528 (N_21528,N_16053,N_17431);
nor U21529 (N_21529,N_18594,N_18018);
nor U21530 (N_21530,N_18480,N_17927);
nand U21531 (N_21531,N_18676,N_17638);
nor U21532 (N_21532,N_16554,N_17171);
nand U21533 (N_21533,N_16656,N_18732);
and U21534 (N_21534,N_18730,N_18275);
nor U21535 (N_21535,N_16695,N_17511);
and U21536 (N_21536,N_17855,N_17627);
xnor U21537 (N_21537,N_18114,N_17744);
and U21538 (N_21538,N_17337,N_18306);
and U21539 (N_21539,N_18617,N_17433);
xor U21540 (N_21540,N_15714,N_16076);
nand U21541 (N_21541,N_15916,N_16220);
or U21542 (N_21542,N_17137,N_17422);
nor U21543 (N_21543,N_18385,N_15947);
nand U21544 (N_21544,N_16916,N_16739);
nand U21545 (N_21545,N_18738,N_17606);
or U21546 (N_21546,N_16617,N_17169);
xor U21547 (N_21547,N_17444,N_17534);
or U21548 (N_21548,N_16743,N_16076);
nor U21549 (N_21549,N_18035,N_16784);
and U21550 (N_21550,N_16622,N_16953);
nor U21551 (N_21551,N_15703,N_18545);
and U21552 (N_21552,N_18206,N_17211);
xnor U21553 (N_21553,N_18633,N_16644);
and U21554 (N_21554,N_16593,N_16058);
nor U21555 (N_21555,N_16739,N_16345);
nor U21556 (N_21556,N_15651,N_18658);
xnor U21557 (N_21557,N_16597,N_18657);
nor U21558 (N_21558,N_18331,N_16104);
nand U21559 (N_21559,N_15761,N_18402);
xor U21560 (N_21560,N_16517,N_17745);
and U21561 (N_21561,N_16529,N_18690);
nand U21562 (N_21562,N_18691,N_18308);
xnor U21563 (N_21563,N_17321,N_15632);
nand U21564 (N_21564,N_16446,N_17295);
xor U21565 (N_21565,N_15741,N_17662);
or U21566 (N_21566,N_16264,N_16838);
nor U21567 (N_21567,N_17745,N_18117);
or U21568 (N_21568,N_17083,N_16268);
nor U21569 (N_21569,N_15963,N_17537);
or U21570 (N_21570,N_18255,N_17592);
xnor U21571 (N_21571,N_15906,N_17938);
and U21572 (N_21572,N_16129,N_18114);
and U21573 (N_21573,N_16960,N_15911);
nand U21574 (N_21574,N_17921,N_16851);
xor U21575 (N_21575,N_17910,N_18272);
or U21576 (N_21576,N_16144,N_16554);
nor U21577 (N_21577,N_18432,N_17910);
nand U21578 (N_21578,N_16203,N_17702);
nor U21579 (N_21579,N_18019,N_16414);
or U21580 (N_21580,N_16228,N_15977);
nand U21581 (N_21581,N_17625,N_16019);
and U21582 (N_21582,N_16617,N_18178);
or U21583 (N_21583,N_18738,N_15928);
or U21584 (N_21584,N_17671,N_16823);
nand U21585 (N_21585,N_17648,N_18492);
xnor U21586 (N_21586,N_17439,N_17671);
nand U21587 (N_21587,N_17141,N_17732);
and U21588 (N_21588,N_16448,N_17307);
and U21589 (N_21589,N_18680,N_17643);
and U21590 (N_21590,N_17067,N_16932);
or U21591 (N_21591,N_17756,N_17741);
nor U21592 (N_21592,N_16967,N_18246);
nor U21593 (N_21593,N_16632,N_18205);
or U21594 (N_21594,N_16398,N_15994);
nand U21595 (N_21595,N_18180,N_15653);
nor U21596 (N_21596,N_17185,N_18327);
nor U21597 (N_21597,N_16237,N_18388);
nor U21598 (N_21598,N_15716,N_16889);
nor U21599 (N_21599,N_17933,N_17964);
nand U21600 (N_21600,N_16861,N_17061);
or U21601 (N_21601,N_15631,N_16636);
nand U21602 (N_21602,N_15988,N_16383);
and U21603 (N_21603,N_17877,N_18376);
nor U21604 (N_21604,N_17048,N_17154);
xor U21605 (N_21605,N_18139,N_16591);
and U21606 (N_21606,N_16835,N_16335);
and U21607 (N_21607,N_16116,N_18021);
or U21608 (N_21608,N_16397,N_16846);
xor U21609 (N_21609,N_15961,N_15633);
nand U21610 (N_21610,N_17715,N_17859);
or U21611 (N_21611,N_18427,N_17514);
and U21612 (N_21612,N_17770,N_18365);
nor U21613 (N_21613,N_17382,N_18418);
nand U21614 (N_21614,N_16763,N_17995);
or U21615 (N_21615,N_18164,N_18744);
nand U21616 (N_21616,N_16003,N_16904);
xnor U21617 (N_21617,N_16865,N_15800);
nand U21618 (N_21618,N_17728,N_17028);
nor U21619 (N_21619,N_17435,N_16591);
nand U21620 (N_21620,N_17023,N_16025);
xor U21621 (N_21621,N_15767,N_16036);
and U21622 (N_21622,N_16327,N_15713);
nand U21623 (N_21623,N_15973,N_18015);
xor U21624 (N_21624,N_18017,N_15751);
nand U21625 (N_21625,N_17575,N_17205);
nand U21626 (N_21626,N_17576,N_17811);
xor U21627 (N_21627,N_18583,N_18063);
and U21628 (N_21628,N_17467,N_17119);
nor U21629 (N_21629,N_15651,N_16516);
nor U21630 (N_21630,N_17943,N_18151);
nor U21631 (N_21631,N_15921,N_18638);
or U21632 (N_21632,N_17350,N_18591);
and U21633 (N_21633,N_17216,N_18737);
nand U21634 (N_21634,N_16875,N_18581);
and U21635 (N_21635,N_17984,N_17507);
and U21636 (N_21636,N_18231,N_17544);
nand U21637 (N_21637,N_16544,N_17810);
xnor U21638 (N_21638,N_15907,N_17837);
nor U21639 (N_21639,N_18361,N_18196);
xor U21640 (N_21640,N_17647,N_16020);
and U21641 (N_21641,N_16992,N_16731);
and U21642 (N_21642,N_17228,N_15765);
and U21643 (N_21643,N_18167,N_18200);
nor U21644 (N_21644,N_18138,N_16209);
and U21645 (N_21645,N_17888,N_18317);
and U21646 (N_21646,N_15684,N_18572);
nand U21647 (N_21647,N_18373,N_17241);
nand U21648 (N_21648,N_18089,N_18272);
or U21649 (N_21649,N_16828,N_18493);
xor U21650 (N_21650,N_16801,N_18648);
nor U21651 (N_21651,N_16131,N_16421);
xor U21652 (N_21652,N_15710,N_16496);
nand U21653 (N_21653,N_17640,N_18047);
xnor U21654 (N_21654,N_16039,N_16158);
nand U21655 (N_21655,N_15689,N_16366);
nand U21656 (N_21656,N_18653,N_17318);
and U21657 (N_21657,N_16412,N_17851);
and U21658 (N_21658,N_17016,N_17487);
nand U21659 (N_21659,N_16430,N_16464);
xor U21660 (N_21660,N_18445,N_15695);
nand U21661 (N_21661,N_16524,N_15831);
nor U21662 (N_21662,N_17086,N_17347);
xor U21663 (N_21663,N_17013,N_17248);
or U21664 (N_21664,N_18596,N_16189);
xnor U21665 (N_21665,N_16731,N_16016);
nor U21666 (N_21666,N_16558,N_18172);
nor U21667 (N_21667,N_17810,N_18208);
or U21668 (N_21668,N_16414,N_16828);
or U21669 (N_21669,N_17952,N_18092);
nor U21670 (N_21670,N_18025,N_17939);
nor U21671 (N_21671,N_18494,N_16443);
nor U21672 (N_21672,N_16353,N_17444);
xnor U21673 (N_21673,N_17428,N_17945);
nor U21674 (N_21674,N_17373,N_16690);
xor U21675 (N_21675,N_16657,N_17675);
xnor U21676 (N_21676,N_16636,N_18330);
nand U21677 (N_21677,N_17307,N_16458);
xnor U21678 (N_21678,N_16070,N_15806);
and U21679 (N_21679,N_18658,N_16609);
xor U21680 (N_21680,N_16233,N_18262);
xnor U21681 (N_21681,N_16217,N_16904);
nor U21682 (N_21682,N_17337,N_16603);
xnor U21683 (N_21683,N_17210,N_17175);
nand U21684 (N_21684,N_16227,N_16781);
xor U21685 (N_21685,N_15685,N_17679);
xor U21686 (N_21686,N_16433,N_15851);
and U21687 (N_21687,N_16299,N_16106);
xnor U21688 (N_21688,N_15946,N_15690);
nor U21689 (N_21689,N_17000,N_17559);
and U21690 (N_21690,N_16371,N_17457);
xnor U21691 (N_21691,N_18302,N_17823);
and U21692 (N_21692,N_16167,N_16034);
or U21693 (N_21693,N_17501,N_18432);
or U21694 (N_21694,N_16400,N_17655);
nor U21695 (N_21695,N_16441,N_18422);
xnor U21696 (N_21696,N_17390,N_17428);
and U21697 (N_21697,N_18211,N_15985);
nor U21698 (N_21698,N_16639,N_17343);
nand U21699 (N_21699,N_18097,N_16210);
and U21700 (N_21700,N_18265,N_18689);
or U21701 (N_21701,N_18314,N_18303);
xor U21702 (N_21702,N_18613,N_16391);
and U21703 (N_21703,N_15711,N_16550);
nor U21704 (N_21704,N_16374,N_17996);
nor U21705 (N_21705,N_17283,N_18145);
and U21706 (N_21706,N_17699,N_17301);
xor U21707 (N_21707,N_18510,N_17726);
nor U21708 (N_21708,N_15745,N_17873);
nor U21709 (N_21709,N_18550,N_18270);
and U21710 (N_21710,N_18130,N_17483);
nand U21711 (N_21711,N_16529,N_16364);
or U21712 (N_21712,N_18574,N_16735);
xor U21713 (N_21713,N_16400,N_17003);
nand U21714 (N_21714,N_16606,N_16918);
xnor U21715 (N_21715,N_17400,N_16434);
and U21716 (N_21716,N_16495,N_16204);
nor U21717 (N_21717,N_18156,N_17062);
nand U21718 (N_21718,N_17302,N_18397);
nor U21719 (N_21719,N_18023,N_15968);
and U21720 (N_21720,N_16248,N_16060);
nand U21721 (N_21721,N_16531,N_17026);
nor U21722 (N_21722,N_16639,N_17017);
nor U21723 (N_21723,N_18241,N_18429);
and U21724 (N_21724,N_18370,N_16823);
nand U21725 (N_21725,N_16690,N_18311);
nand U21726 (N_21726,N_17463,N_17976);
or U21727 (N_21727,N_15999,N_16207);
and U21728 (N_21728,N_15944,N_16816);
and U21729 (N_21729,N_18415,N_16795);
or U21730 (N_21730,N_18638,N_17697);
nand U21731 (N_21731,N_18610,N_17301);
nand U21732 (N_21732,N_16562,N_18739);
nand U21733 (N_21733,N_18097,N_17485);
and U21734 (N_21734,N_15840,N_17139);
or U21735 (N_21735,N_16329,N_17115);
nand U21736 (N_21736,N_17147,N_15707);
nand U21737 (N_21737,N_17877,N_15810);
nand U21738 (N_21738,N_16352,N_16185);
or U21739 (N_21739,N_17716,N_18359);
xor U21740 (N_21740,N_17916,N_18256);
and U21741 (N_21741,N_17612,N_17227);
nand U21742 (N_21742,N_17038,N_16954);
and U21743 (N_21743,N_17078,N_18248);
xnor U21744 (N_21744,N_18617,N_16702);
xor U21745 (N_21745,N_16358,N_16071);
nand U21746 (N_21746,N_17997,N_17612);
and U21747 (N_21747,N_18081,N_16263);
and U21748 (N_21748,N_16000,N_17813);
xor U21749 (N_21749,N_15708,N_16924);
xnor U21750 (N_21750,N_17135,N_17643);
nor U21751 (N_21751,N_17258,N_17594);
nor U21752 (N_21752,N_17101,N_17731);
xor U21753 (N_21753,N_17304,N_18369);
or U21754 (N_21754,N_17949,N_15638);
and U21755 (N_21755,N_17442,N_17028);
and U21756 (N_21756,N_18353,N_17521);
nand U21757 (N_21757,N_17793,N_16042);
xor U21758 (N_21758,N_18357,N_18039);
nand U21759 (N_21759,N_15626,N_16554);
and U21760 (N_21760,N_16549,N_16222);
and U21761 (N_21761,N_18291,N_17463);
nor U21762 (N_21762,N_17416,N_18285);
xnor U21763 (N_21763,N_17918,N_16709);
nor U21764 (N_21764,N_15673,N_17855);
nand U21765 (N_21765,N_17711,N_17340);
nor U21766 (N_21766,N_17112,N_15632);
and U21767 (N_21767,N_17135,N_15732);
nor U21768 (N_21768,N_18501,N_17578);
nor U21769 (N_21769,N_16804,N_18041);
or U21770 (N_21770,N_16366,N_18534);
nand U21771 (N_21771,N_16678,N_15740);
xnor U21772 (N_21772,N_15913,N_18610);
nand U21773 (N_21773,N_18083,N_16685);
xnor U21774 (N_21774,N_17993,N_17868);
or U21775 (N_21775,N_15785,N_16910);
nand U21776 (N_21776,N_17545,N_17450);
nor U21777 (N_21777,N_18376,N_17141);
nand U21778 (N_21778,N_16322,N_15980);
xor U21779 (N_21779,N_17676,N_17053);
xnor U21780 (N_21780,N_15888,N_16530);
and U21781 (N_21781,N_16122,N_16929);
xor U21782 (N_21782,N_17687,N_18128);
and U21783 (N_21783,N_17972,N_16107);
xnor U21784 (N_21784,N_16944,N_18027);
or U21785 (N_21785,N_16041,N_17086);
or U21786 (N_21786,N_16156,N_15762);
xnor U21787 (N_21787,N_17519,N_17793);
or U21788 (N_21788,N_16046,N_18122);
nand U21789 (N_21789,N_16033,N_18400);
xor U21790 (N_21790,N_15905,N_16603);
and U21791 (N_21791,N_17527,N_18715);
xor U21792 (N_21792,N_16843,N_18335);
nand U21793 (N_21793,N_16566,N_15693);
xor U21794 (N_21794,N_17380,N_16774);
nor U21795 (N_21795,N_16903,N_17561);
or U21796 (N_21796,N_16574,N_18205);
and U21797 (N_21797,N_17920,N_17136);
xor U21798 (N_21798,N_17764,N_18096);
nand U21799 (N_21799,N_18344,N_16695);
and U21800 (N_21800,N_17995,N_18124);
nor U21801 (N_21801,N_16046,N_17200);
and U21802 (N_21802,N_16179,N_15754);
nand U21803 (N_21803,N_17244,N_17581);
or U21804 (N_21804,N_17754,N_18321);
or U21805 (N_21805,N_18230,N_18613);
and U21806 (N_21806,N_18544,N_17684);
and U21807 (N_21807,N_16162,N_18671);
xnor U21808 (N_21808,N_17078,N_16300);
xor U21809 (N_21809,N_16510,N_16121);
and U21810 (N_21810,N_16208,N_16712);
or U21811 (N_21811,N_18249,N_17538);
xor U21812 (N_21812,N_17483,N_18137);
and U21813 (N_21813,N_17624,N_18454);
nand U21814 (N_21814,N_16222,N_17814);
and U21815 (N_21815,N_17977,N_17897);
xnor U21816 (N_21816,N_16782,N_16242);
nand U21817 (N_21817,N_18600,N_18319);
xor U21818 (N_21818,N_17241,N_17187);
nor U21819 (N_21819,N_18586,N_17490);
xnor U21820 (N_21820,N_17057,N_16025);
nand U21821 (N_21821,N_17336,N_16110);
or U21822 (N_21822,N_17233,N_16849);
or U21823 (N_21823,N_16628,N_17194);
nand U21824 (N_21824,N_17836,N_18124);
xor U21825 (N_21825,N_16391,N_17722);
and U21826 (N_21826,N_17161,N_17908);
or U21827 (N_21827,N_16067,N_18216);
or U21828 (N_21828,N_18737,N_17382);
xnor U21829 (N_21829,N_18580,N_15654);
nor U21830 (N_21830,N_15704,N_17453);
xor U21831 (N_21831,N_15655,N_15770);
and U21832 (N_21832,N_15682,N_15989);
nand U21833 (N_21833,N_17691,N_16890);
nand U21834 (N_21834,N_16915,N_17772);
and U21835 (N_21835,N_15828,N_18583);
and U21836 (N_21836,N_17281,N_16510);
or U21837 (N_21837,N_16480,N_16851);
or U21838 (N_21838,N_17274,N_17500);
and U21839 (N_21839,N_17249,N_16718);
nor U21840 (N_21840,N_16497,N_18257);
nand U21841 (N_21841,N_17096,N_16867);
xor U21842 (N_21842,N_16740,N_17643);
nand U21843 (N_21843,N_18098,N_16241);
nor U21844 (N_21844,N_16098,N_15989);
xnor U21845 (N_21845,N_17731,N_18618);
and U21846 (N_21846,N_15725,N_16364);
xnor U21847 (N_21847,N_17773,N_17416);
or U21848 (N_21848,N_15679,N_18038);
nor U21849 (N_21849,N_16417,N_17443);
nand U21850 (N_21850,N_15899,N_17483);
and U21851 (N_21851,N_16520,N_16516);
nand U21852 (N_21852,N_16265,N_15674);
and U21853 (N_21853,N_18007,N_18690);
and U21854 (N_21854,N_17802,N_18368);
nor U21855 (N_21855,N_17754,N_16831);
nor U21856 (N_21856,N_18576,N_17034);
and U21857 (N_21857,N_15675,N_15924);
and U21858 (N_21858,N_17697,N_17686);
and U21859 (N_21859,N_18422,N_17505);
and U21860 (N_21860,N_17657,N_18310);
xor U21861 (N_21861,N_18341,N_18675);
nor U21862 (N_21862,N_17817,N_18397);
nand U21863 (N_21863,N_17981,N_17667);
and U21864 (N_21864,N_18483,N_15708);
xnor U21865 (N_21865,N_17757,N_16028);
xor U21866 (N_21866,N_18386,N_16763);
nand U21867 (N_21867,N_17635,N_18320);
nand U21868 (N_21868,N_15644,N_18089);
and U21869 (N_21869,N_17163,N_18681);
nor U21870 (N_21870,N_17536,N_16706);
nand U21871 (N_21871,N_15884,N_16509);
nand U21872 (N_21872,N_16121,N_18566);
xor U21873 (N_21873,N_16609,N_16720);
nand U21874 (N_21874,N_18463,N_17883);
or U21875 (N_21875,N_19044,N_20421);
and U21876 (N_21876,N_20559,N_21836);
nand U21877 (N_21877,N_20253,N_20019);
xor U21878 (N_21878,N_20143,N_21196);
nor U21879 (N_21879,N_20504,N_21038);
nand U21880 (N_21880,N_21316,N_18764);
xor U21881 (N_21881,N_20121,N_20003);
nand U21882 (N_21882,N_19047,N_21711);
nor U21883 (N_21883,N_21515,N_21347);
nand U21884 (N_21884,N_21425,N_19775);
and U21885 (N_21885,N_19178,N_21848);
and U21886 (N_21886,N_21719,N_20079);
xnor U21887 (N_21887,N_21050,N_19256);
and U21888 (N_21888,N_20746,N_20583);
nor U21889 (N_21889,N_20795,N_20387);
nor U21890 (N_21890,N_20759,N_20651);
and U21891 (N_21891,N_19018,N_20441);
nand U21892 (N_21892,N_19680,N_19569);
nand U21893 (N_21893,N_20500,N_21390);
or U21894 (N_21894,N_19165,N_21784);
nand U21895 (N_21895,N_19006,N_21767);
nand U21896 (N_21896,N_20896,N_19110);
nor U21897 (N_21897,N_20198,N_21583);
or U21898 (N_21898,N_21227,N_19790);
nand U21899 (N_21899,N_20577,N_19619);
and U21900 (N_21900,N_20955,N_19304);
nor U21901 (N_21901,N_20111,N_18924);
nand U21902 (N_21902,N_21676,N_20957);
xnor U21903 (N_21903,N_21803,N_19345);
and U21904 (N_21904,N_19016,N_19895);
and U21905 (N_21905,N_20765,N_20215);
or U21906 (N_21906,N_20308,N_20952);
nor U21907 (N_21907,N_20332,N_19405);
nor U21908 (N_21908,N_21539,N_20794);
xnor U21909 (N_21909,N_21060,N_19161);
and U21910 (N_21910,N_20021,N_20417);
nor U21911 (N_21911,N_19782,N_21604);
or U21912 (N_21912,N_18968,N_20047);
and U21913 (N_21913,N_20467,N_21426);
or U21914 (N_21914,N_18915,N_19787);
nand U21915 (N_21915,N_19396,N_21269);
nand U21916 (N_21916,N_19003,N_19336);
nand U21917 (N_21917,N_21482,N_19556);
nand U21918 (N_21918,N_21234,N_20035);
xor U21919 (N_21919,N_20127,N_20989);
nand U21920 (N_21920,N_20146,N_19261);
nand U21921 (N_21921,N_19363,N_19102);
xor U21922 (N_21922,N_21845,N_21627);
nor U21923 (N_21923,N_19733,N_19633);
or U21924 (N_21924,N_18964,N_20644);
xnor U21925 (N_21925,N_20083,N_20687);
or U21926 (N_21926,N_19966,N_19111);
or U21927 (N_21927,N_19947,N_21802);
nor U21928 (N_21928,N_19411,N_20766);
nand U21929 (N_21929,N_18965,N_20106);
or U21930 (N_21930,N_21785,N_20109);
or U21931 (N_21931,N_21669,N_20945);
or U21932 (N_21932,N_20597,N_19313);
nor U21933 (N_21933,N_21260,N_19464);
nand U21934 (N_21934,N_21643,N_21157);
or U21935 (N_21935,N_20565,N_20623);
nor U21936 (N_21936,N_21186,N_18894);
nor U21937 (N_21937,N_19788,N_20114);
xor U21938 (N_21938,N_19539,N_20407);
or U21939 (N_21939,N_19082,N_20562);
and U21940 (N_21940,N_20844,N_20991);
or U21941 (N_21941,N_19154,N_20921);
nand U21942 (N_21942,N_19192,N_19855);
nor U21943 (N_21943,N_20434,N_20399);
xnor U21944 (N_21944,N_19439,N_20339);
nand U21945 (N_21945,N_18853,N_21179);
nand U21946 (N_21946,N_18805,N_21221);
nand U21947 (N_21947,N_19284,N_19393);
xor U21948 (N_21948,N_19766,N_21026);
or U21949 (N_21949,N_21014,N_20133);
nor U21950 (N_21950,N_20272,N_19061);
nand U21951 (N_21951,N_19862,N_19104);
and U21952 (N_21952,N_21144,N_20684);
nor U21953 (N_21953,N_19942,N_20920);
nor U21954 (N_21954,N_20700,N_18937);
nor U21955 (N_21955,N_19728,N_18942);
or U21956 (N_21956,N_20251,N_20400);
xor U21957 (N_21957,N_20942,N_20428);
or U21958 (N_21958,N_20784,N_21125);
and U21959 (N_21959,N_21183,N_20906);
nor U21960 (N_21960,N_21556,N_21531);
nor U21961 (N_21961,N_19786,N_20908);
xnor U21962 (N_21962,N_20476,N_19287);
nor U21963 (N_21963,N_20134,N_21790);
or U21964 (N_21964,N_20309,N_19605);
and U21965 (N_21965,N_18847,N_21695);
xor U21966 (N_21966,N_19751,N_21787);
nor U21967 (N_21967,N_19199,N_19837);
nand U21968 (N_21968,N_21015,N_20981);
nand U21969 (N_21969,N_21549,N_19524);
nand U21970 (N_21970,N_21085,N_20255);
nor U21971 (N_21971,N_19635,N_19993);
or U21972 (N_21972,N_19435,N_20674);
nand U21973 (N_21973,N_21619,N_19239);
nor U21974 (N_21974,N_19298,N_21121);
or U21975 (N_21975,N_19921,N_20474);
nand U21976 (N_21976,N_21297,N_18836);
xor U21977 (N_21977,N_21609,N_21670);
nor U21978 (N_21978,N_20691,N_18833);
or U21979 (N_21979,N_20136,N_21587);
and U21980 (N_21980,N_19692,N_20366);
nor U21981 (N_21981,N_19586,N_20120);
nand U21982 (N_21982,N_21516,N_19241);
nor U21983 (N_21983,N_20196,N_20786);
xor U21984 (N_21984,N_19606,N_20837);
or U21985 (N_21985,N_20201,N_20773);
or U21986 (N_21986,N_18825,N_19931);
and U21987 (N_21987,N_21341,N_21285);
nand U21988 (N_21988,N_21830,N_19528);
and U21989 (N_21989,N_20665,N_21766);
xnor U21990 (N_21990,N_19328,N_20987);
xor U21991 (N_21991,N_21352,N_19088);
nand U21992 (N_21992,N_19231,N_20066);
xnor U21993 (N_21993,N_18835,N_19317);
and U21994 (N_21994,N_18898,N_20688);
nand U21995 (N_21995,N_19505,N_20246);
nand U21996 (N_21996,N_21206,N_19449);
nor U21997 (N_21997,N_19355,N_20963);
or U21998 (N_21998,N_20697,N_21419);
or U21999 (N_21999,N_19567,N_19615);
and U22000 (N_22000,N_19932,N_19901);
nand U22001 (N_22001,N_19098,N_20333);
nand U22002 (N_22002,N_19688,N_21646);
nand U22003 (N_22003,N_19040,N_20866);
and U22004 (N_22004,N_20703,N_20226);
and U22005 (N_22005,N_21118,N_19598);
or U22006 (N_22006,N_19209,N_21422);
nand U22007 (N_22007,N_21020,N_18930);
xnor U22008 (N_22008,N_21872,N_20254);
nor U22009 (N_22009,N_21454,N_18954);
and U22010 (N_22010,N_19202,N_20154);
and U22011 (N_22011,N_19525,N_20704);
xnor U22012 (N_22012,N_21493,N_21280);
xor U22013 (N_22013,N_18990,N_19011);
or U22014 (N_22014,N_19080,N_20639);
and U22015 (N_22015,N_18786,N_19059);
and U22016 (N_22016,N_19371,N_19024);
and U22017 (N_22017,N_19297,N_20429);
xor U22018 (N_22018,N_19455,N_20926);
xor U22019 (N_22019,N_21483,N_19235);
and U22020 (N_22020,N_21415,N_18939);
and U22021 (N_22021,N_19395,N_20596);
nor U22022 (N_22022,N_19268,N_20600);
and U22023 (N_22023,N_21374,N_18840);
xnor U22024 (N_22024,N_20884,N_21017);
nor U22025 (N_22025,N_20064,N_19175);
and U22026 (N_22026,N_20128,N_21601);
xnor U22027 (N_22027,N_21624,N_19714);
or U22028 (N_22028,N_19697,N_21197);
nor U22029 (N_22029,N_20473,N_21431);
xnor U22030 (N_22030,N_19206,N_21355);
nand U22031 (N_22031,N_20498,N_21674);
or U22032 (N_22032,N_20548,N_20809);
xor U22033 (N_22033,N_21198,N_19112);
xor U22034 (N_22034,N_20078,N_20401);
or U22035 (N_22035,N_21473,N_21294);
nand U22036 (N_22036,N_20449,N_20211);
and U22037 (N_22037,N_19547,N_19283);
or U22038 (N_22038,N_19715,N_20444);
and U22039 (N_22039,N_20274,N_21725);
nand U22040 (N_22040,N_19427,N_18986);
or U22041 (N_22041,N_19866,N_20937);
xnor U22042 (N_22042,N_19276,N_20068);
nor U22043 (N_22043,N_21520,N_21292);
or U22044 (N_22044,N_19307,N_20291);
xnor U22045 (N_22045,N_18839,N_20698);
and U22046 (N_22046,N_20129,N_21598);
or U22047 (N_22047,N_19578,N_19172);
and U22048 (N_22048,N_20002,N_19867);
nand U22049 (N_22049,N_21545,N_19211);
or U22050 (N_22050,N_20769,N_20184);
xor U22051 (N_22051,N_19538,N_20280);
nand U22052 (N_22052,N_20220,N_19094);
and U22053 (N_22053,N_21450,N_20005);
and U22054 (N_22054,N_19327,N_20203);
or U22055 (N_22055,N_21019,N_20119);
xor U22056 (N_22056,N_20414,N_18961);
nand U22057 (N_22057,N_19764,N_21841);
nor U22058 (N_22058,N_18953,N_19353);
or U22059 (N_22059,N_21332,N_19067);
nor U22060 (N_22060,N_19968,N_19823);
nor U22061 (N_22061,N_20459,N_21022);
or U22062 (N_22062,N_20008,N_21456);
or U22063 (N_22063,N_19919,N_19724);
xor U22064 (N_22064,N_20774,N_20526);
nand U22065 (N_22065,N_19796,N_20994);
xor U22066 (N_22066,N_18903,N_21046);
nor U22067 (N_22067,N_20566,N_19999);
and U22068 (N_22068,N_19233,N_19720);
nor U22069 (N_22069,N_20607,N_21595);
nand U22070 (N_22070,N_20797,N_20673);
xnor U22071 (N_22071,N_19099,N_19700);
or U22072 (N_22072,N_19851,N_21180);
nor U22073 (N_22073,N_21187,N_21247);
xor U22074 (N_22074,N_20663,N_19017);
nor U22075 (N_22075,N_19789,N_20675);
xnor U22076 (N_22076,N_19669,N_21164);
and U22077 (N_22077,N_20683,N_21055);
nand U22078 (N_22078,N_21647,N_20237);
or U22079 (N_22079,N_19526,N_21690);
or U22080 (N_22080,N_21145,N_21857);
xnor U22081 (N_22081,N_19458,N_20368);
or U22082 (N_22082,N_20167,N_19169);
nor U22083 (N_22083,N_20988,N_20581);
nor U22084 (N_22084,N_19792,N_21555);
nand U22085 (N_22085,N_19873,N_18802);
or U22086 (N_22086,N_20158,N_21402);
xor U22087 (N_22087,N_19509,N_21066);
nor U22088 (N_22088,N_19021,N_19708);
nand U22089 (N_22089,N_18871,N_20568);
nor U22090 (N_22090,N_19058,N_19618);
or U22091 (N_22091,N_21165,N_19709);
and U22092 (N_22092,N_19254,N_21650);
nor U22093 (N_22093,N_19324,N_21827);
xnor U22094 (N_22094,N_20325,N_20445);
nand U22095 (N_22095,N_21585,N_21272);
nand U22096 (N_22096,N_20218,N_19632);
nand U22097 (N_22097,N_19779,N_21692);
or U22098 (N_22098,N_21448,N_20686);
or U22099 (N_22099,N_20446,N_21253);
nand U22100 (N_22100,N_20488,N_19773);
nand U22101 (N_22101,N_21252,N_21840);
or U22102 (N_22102,N_19426,N_21447);
xnor U22103 (N_22103,N_19945,N_21632);
xor U22104 (N_22104,N_20013,N_21308);
xor U22105 (N_22105,N_20372,N_20398);
nand U22106 (N_22106,N_18778,N_20865);
or U22107 (N_22107,N_21811,N_19188);
and U22108 (N_22108,N_19460,N_21392);
xor U22109 (N_22109,N_20749,N_20670);
and U22110 (N_22110,N_19753,N_21514);
nor U22111 (N_22111,N_20599,N_20553);
or U22112 (N_22112,N_20560,N_20163);
or U22113 (N_22113,N_21789,N_20277);
and U22114 (N_22114,N_21133,N_21207);
and U22115 (N_22115,N_19335,N_19760);
nand U22116 (N_22116,N_21867,N_20102);
nand U22117 (N_22117,N_20880,N_20397);
nand U22118 (N_22118,N_20307,N_21574);
nor U22119 (N_22119,N_21863,N_19711);
nand U22120 (N_22120,N_20931,N_21455);
or U22121 (N_22121,N_20721,N_18974);
nor U22122 (N_22122,N_18977,N_19886);
nor U22123 (N_22123,N_19988,N_20854);
xnor U22124 (N_22124,N_19656,N_20071);
nor U22125 (N_22125,N_19983,N_18820);
xnor U22126 (N_22126,N_19349,N_21758);
and U22127 (N_22127,N_19332,N_20739);
or U22128 (N_22128,N_20725,N_21522);
nand U22129 (N_22129,N_21652,N_21502);
nand U22130 (N_22130,N_20629,N_20057);
and U22131 (N_22131,N_19022,N_21255);
nor U22132 (N_22132,N_19486,N_19212);
or U22133 (N_22133,N_20342,N_20415);
or U22134 (N_22134,N_20477,N_20744);
nand U22135 (N_22135,N_20084,N_19592);
and U22136 (N_22136,N_21034,N_19330);
xor U22137 (N_22137,N_20023,N_21077);
and U22138 (N_22138,N_19684,N_19155);
nand U22139 (N_22139,N_20267,N_21788);
and U22140 (N_22140,N_20585,N_21365);
or U22141 (N_22141,N_21833,N_19950);
or U22142 (N_22142,N_19035,N_19874);
nand U22143 (N_22143,N_21203,N_20048);
xnor U22144 (N_22144,N_19593,N_19951);
nor U22145 (N_22145,N_19809,N_20879);
and U22146 (N_22146,N_21656,N_19713);
nand U22147 (N_22147,N_19638,N_21813);
and U22148 (N_22148,N_19127,N_20259);
and U22149 (N_22149,N_20666,N_21527);
and U22150 (N_22150,N_21101,N_18900);
and U22151 (N_22151,N_21375,N_21156);
nand U22152 (N_22152,N_19833,N_21357);
nor U22153 (N_22153,N_20935,N_20932);
xor U22154 (N_22154,N_21391,N_21128);
nand U22155 (N_22155,N_20614,N_21293);
nor U22156 (N_22156,N_20507,N_20485);
or U22157 (N_22157,N_20223,N_19323);
and U22158 (N_22158,N_20505,N_19816);
or U22159 (N_22159,N_18982,N_19939);
nand U22160 (N_22160,N_21302,N_19604);
nor U22161 (N_22161,N_19534,N_19431);
nand U22162 (N_22162,N_20524,N_21074);
nor U22163 (N_22163,N_21139,N_19845);
nand U22164 (N_22164,N_20609,N_21136);
or U22165 (N_22165,N_19038,N_19875);
nand U22166 (N_22166,N_21846,N_19574);
and U22167 (N_22167,N_21562,N_19506);
nand U22168 (N_22168,N_19594,N_21258);
xnor U22169 (N_22169,N_20189,N_20409);
nor U22170 (N_22170,N_20723,N_21437);
xnor U22171 (N_22171,N_20925,N_21579);
nand U22172 (N_22172,N_19027,N_18843);
and U22173 (N_22173,N_21218,N_20338);
nor U22174 (N_22174,N_20099,N_20902);
and U22175 (N_22175,N_18766,N_19634);
nor U22176 (N_22176,N_19914,N_20802);
or U22177 (N_22177,N_21608,N_20382);
or U22178 (N_22178,N_21873,N_20443);
xnor U22179 (N_22179,N_19726,N_20039);
nor U22180 (N_22180,N_21773,N_19275);
and U22181 (N_22181,N_21501,N_21205);
and U22182 (N_22182,N_19761,N_21148);
nand U22183 (N_22183,N_18812,N_19041);
nor U22184 (N_22184,N_21305,N_19143);
or U22185 (N_22185,N_19191,N_20849);
nand U22186 (N_22186,N_18969,N_19938);
nand U22187 (N_22187,N_20710,N_21404);
or U22188 (N_22188,N_20360,N_20394);
nor U22189 (N_22189,N_19544,N_21052);
nand U22190 (N_22190,N_20539,N_21720);
nor U22191 (N_22191,N_20895,N_18884);
xor U22192 (N_22192,N_20395,N_19471);
xnor U22193 (N_22193,N_21783,N_21622);
and U22194 (N_22194,N_20017,N_20391);
and U22195 (N_22195,N_19401,N_19470);
and U22196 (N_22196,N_21409,N_19358);
nand U22197 (N_22197,N_18854,N_21572);
or U22198 (N_22198,N_19805,N_21508);
nand U22199 (N_22199,N_19677,N_21786);
and U22200 (N_22200,N_20363,N_19810);
nor U22201 (N_22201,N_19870,N_20516);
nor U22202 (N_22202,N_20883,N_19923);
nand U22203 (N_22203,N_21770,N_20601);
xor U22204 (N_22204,N_20617,N_21487);
and U22205 (N_22205,N_21781,N_20751);
nand U22206 (N_22206,N_19438,N_18760);
nand U22207 (N_22207,N_20501,N_21538);
nand U22208 (N_22208,N_20521,N_21368);
or U22209 (N_22209,N_21801,N_21058);
and U22210 (N_22210,N_19571,N_18856);
nand U22211 (N_22211,N_19124,N_20091);
or U22212 (N_22212,N_19179,N_20475);
nor U22213 (N_22213,N_19889,N_21199);
nor U22214 (N_22214,N_20640,N_19797);
or U22215 (N_22215,N_19767,N_21263);
and U22216 (N_22216,N_19693,N_21828);
nand U22217 (N_22217,N_19280,N_19882);
xor U22218 (N_22218,N_19636,N_19665);
nand U22219 (N_22219,N_18978,N_19650);
nor U22220 (N_22220,N_21230,N_21703);
xnor U22221 (N_22221,N_21212,N_21648);
and U22222 (N_22222,N_19387,N_21742);
or U22223 (N_22223,N_21819,N_20904);
xnor U22224 (N_22224,N_20555,N_19356);
nand U22225 (N_22225,N_21868,N_19857);
xnor U22226 (N_22226,N_18851,N_18813);
and U22227 (N_22227,N_21581,N_19519);
nand U22228 (N_22228,N_18777,N_21712);
and U22229 (N_22229,N_19483,N_20734);
nand U22230 (N_22230,N_19613,N_20396);
xnor U22231 (N_22231,N_20460,N_20612);
nor U22232 (N_22232,N_20826,N_21701);
or U22233 (N_22233,N_21638,N_19595);
and U22234 (N_22234,N_20388,N_20692);
or U22235 (N_22235,N_19050,N_18941);
or U22236 (N_22236,N_19031,N_19842);
and U22237 (N_22237,N_20043,N_20205);
nand U22238 (N_22238,N_21382,N_20406);
xor U22239 (N_22239,N_18866,N_19236);
nand U22240 (N_22240,N_21797,N_21244);
xnor U22241 (N_22241,N_20798,N_21492);
nor U22242 (N_22242,N_20719,N_20430);
nand U22243 (N_22243,N_21159,N_19351);
xor U22244 (N_22244,N_19272,N_18781);
nor U22245 (N_22245,N_20789,N_21043);
or U22246 (N_22246,N_19529,N_19090);
nor U22247 (N_22247,N_20094,N_20537);
nor U22248 (N_22248,N_21189,N_19601);
and U22249 (N_22249,N_19116,N_21548);
and U22250 (N_22250,N_20520,N_19830);
or U22251 (N_22251,N_21319,N_21132);
xor U22252 (N_22252,N_21488,N_21268);
xor U22253 (N_22253,N_21698,N_20860);
nand U22254 (N_22254,N_20953,N_19091);
xor U22255 (N_22255,N_21223,N_19461);
nand U22256 (N_22256,N_20660,N_21000);
xnor U22257 (N_22257,N_21045,N_19156);
xor U22258 (N_22258,N_20727,N_20918);
nor U22259 (N_22259,N_19844,N_19648);
xor U22260 (N_22260,N_20210,N_21644);
nor U22261 (N_22261,N_21405,N_20310);
and U22262 (N_22262,N_19400,N_20871);
nand U22263 (N_22263,N_19074,N_21340);
and U22264 (N_22264,N_21109,N_20040);
or U22265 (N_22265,N_19681,N_21284);
nor U22266 (N_22266,N_19294,N_21602);
or U22267 (N_22267,N_20060,N_21612);
and U22268 (N_22268,N_21339,N_20208);
or U22269 (N_22269,N_21182,N_20052);
xnor U22270 (N_22270,N_21024,N_19360);
xor U22271 (N_22271,N_21710,N_21202);
nor U22272 (N_22272,N_18882,N_21591);
and U22273 (N_22273,N_20911,N_21168);
xnor U22274 (N_22274,N_19368,N_20236);
nor U22275 (N_22275,N_20682,N_20243);
or U22276 (N_22276,N_21705,N_20404);
nor U22277 (N_22277,N_19570,N_18928);
and U22278 (N_22278,N_18842,N_19247);
nor U22279 (N_22279,N_20074,N_19030);
and U22280 (N_22280,N_19777,N_21664);
and U22281 (N_22281,N_19558,N_20392);
nand U22282 (N_22282,N_19279,N_20062);
xnor U22283 (N_22283,N_19694,N_21370);
nor U22284 (N_22284,N_20100,N_19992);
or U22285 (N_22285,N_20293,N_21858);
xor U22286 (N_22286,N_19144,N_19496);
or U22287 (N_22287,N_20875,N_20093);
nor U22288 (N_22288,N_21775,N_20820);
nand U22289 (N_22289,N_20534,N_20419);
and U22290 (N_22290,N_18792,N_19442);
xor U22291 (N_22291,N_20736,N_19630);
and U22292 (N_22292,N_20606,N_21233);
nand U22293 (N_22293,N_20993,N_20341);
nor U22294 (N_22294,N_20910,N_20265);
nor U22295 (N_22295,N_19004,N_19293);
or U22296 (N_22296,N_20178,N_19002);
nor U22297 (N_22297,N_20768,N_21700);
and U22298 (N_22298,N_19884,N_20235);
or U22299 (N_22299,N_18877,N_18796);
nor U22300 (N_22300,N_21717,N_18826);
nand U22301 (N_22301,N_20353,N_19549);
xor U22302 (N_22302,N_19955,N_18962);
nand U22303 (N_22303,N_19057,N_19226);
nor U22304 (N_22304,N_21411,N_21076);
or U22305 (N_22305,N_21418,N_19434);
nand U22306 (N_22306,N_20536,N_19652);
xor U22307 (N_22307,N_19214,N_19820);
and U22308 (N_22308,N_19671,N_19954);
nand U22309 (N_22309,N_20648,N_19913);
nand U22310 (N_22310,N_19063,N_20668);
nand U22311 (N_22311,N_21095,N_19367);
or U22312 (N_22312,N_19893,N_21800);
xor U22313 (N_22313,N_21304,N_19085);
nand U22314 (N_22314,N_19150,N_21185);
and U22315 (N_22315,N_18875,N_18799);
and U22316 (N_22316,N_21265,N_21861);
nor U22317 (N_22317,N_21016,N_21238);
nand U22318 (N_22318,N_20222,N_18996);
or U22319 (N_22319,N_20365,N_19487);
or U22320 (N_22320,N_19748,N_20279);
nor U22321 (N_22321,N_21373,N_21603);
xor U22322 (N_22322,N_19871,N_18992);
nand U22323 (N_22323,N_21350,N_19778);
or U22324 (N_22324,N_19900,N_19987);
nand U22325 (N_22325,N_19846,N_21540);
nand U22326 (N_22326,N_19252,N_21542);
nand U22327 (N_22327,N_21772,N_19507);
nand U22328 (N_22328,N_19457,N_21140);
nor U22329 (N_22329,N_20224,N_21636);
xnor U22330 (N_22330,N_18972,N_21249);
and U22331 (N_22331,N_20888,N_20130);
nand U22332 (N_22332,N_18838,N_19488);
xor U22333 (N_22333,N_19702,N_19691);
nor U22334 (N_22334,N_20929,N_19357);
nand U22335 (N_22335,N_18780,N_20087);
xnor U22336 (N_22336,N_19131,N_20499);
and U22337 (N_22337,N_21310,N_20138);
nor U22338 (N_22338,N_18989,N_21831);
or U22339 (N_22339,N_19645,N_21315);
and U22340 (N_22340,N_19614,N_19537);
nor U22341 (N_22341,N_19465,N_20627);
xnor U22342 (N_22342,N_20861,N_21311);
and U22343 (N_22343,N_20755,N_19213);
nand U22344 (N_22344,N_18862,N_19958);
xnor U22345 (N_22345,N_19642,N_20761);
or U22346 (N_22346,N_21554,N_19278);
and U22347 (N_22347,N_20076,N_21414);
nor U22348 (N_22348,N_19736,N_21250);
and U22349 (N_22349,N_21408,N_21459);
and U22350 (N_22350,N_19459,N_21222);
or U22351 (N_22351,N_20800,N_21287);
and U22352 (N_22352,N_19666,N_19164);
xor U22353 (N_22353,N_19072,N_19557);
nor U22354 (N_22354,N_18929,N_21283);
xnor U22355 (N_22355,N_20180,N_19291);
xnor U22356 (N_22356,N_21081,N_21178);
or U22357 (N_22357,N_20016,N_21626);
or U22358 (N_22358,N_19667,N_20266);
and U22359 (N_22359,N_19429,N_20225);
nor U22360 (N_22360,N_19474,N_19783);
nand U22361 (N_22361,N_20233,N_19548);
xnor U22362 (N_22362,N_18897,N_20461);
and U22363 (N_22363,N_20190,N_19589);
nor U22364 (N_22364,N_19916,N_20113);
or U22365 (N_22365,N_20754,N_20436);
xnor U22366 (N_22366,N_18943,N_21855);
nand U22367 (N_22367,N_20695,N_20056);
xor U22368 (N_22368,N_21033,N_20662);
nand U22369 (N_22369,N_20028,N_18869);
nor U22370 (N_22370,N_20029,N_20359);
nand U22371 (N_22371,N_21281,N_20781);
nor U22372 (N_22372,N_20077,N_19503);
nor U22373 (N_22373,N_21557,N_20856);
or U22374 (N_22374,N_19378,N_19477);
nor U22375 (N_22375,N_19971,N_19300);
or U22376 (N_22376,N_21429,N_21433);
nor U22377 (N_22377,N_18754,N_21398);
nand U22378 (N_22378,N_19189,N_20250);
nor U22379 (N_22379,N_19695,N_19927);
and U22380 (N_22380,N_21093,N_20709);
or U22381 (N_22381,N_19575,N_21778);
nor U22382 (N_22382,N_21423,N_20960);
or U22383 (N_22383,N_20822,N_19026);
nor U22384 (N_22384,N_21291,N_20081);
and U22385 (N_22385,N_21078,N_20045);
and U22386 (N_22386,N_21737,N_19303);
or U22387 (N_22387,N_19746,N_20635);
or U22388 (N_22388,N_20491,N_21177);
and U22389 (N_22389,N_19984,N_19649);
xor U22390 (N_22390,N_21843,N_20095);
nor U22391 (N_22391,N_21678,N_20801);
nand U22392 (N_22392,N_21615,N_21477);
or U22393 (N_22393,N_21239,N_21677);
nor U22394 (N_22394,N_19129,N_20864);
nand U22395 (N_22395,N_19204,N_19655);
and U22396 (N_22396,N_21449,N_21734);
nand U22397 (N_22397,N_20364,N_21842);
nor U22398 (N_22398,N_21560,N_21796);
nand U22399 (N_22399,N_19196,N_20869);
and U22400 (N_22400,N_21641,N_19877);
xor U22401 (N_22401,N_21282,N_20729);
and U22402 (N_22402,N_21289,N_19141);
or U22403 (N_22403,N_21353,N_21062);
or U22404 (N_22404,N_18770,N_19086);
or U22405 (N_22405,N_20484,N_20448);
or U22406 (N_22406,N_20027,N_21823);
xnor U22407 (N_22407,N_21577,N_20540);
or U22408 (N_22408,N_20641,N_20142);
nor U22409 (N_22409,N_21485,N_21427);
nand U22410 (N_22410,N_19218,N_19568);
nand U22411 (N_22411,N_20815,N_21529);
or U22412 (N_22412,N_20447,N_21495);
nor U22413 (N_22413,N_20916,N_20104);
and U22414 (N_22414,N_20433,N_19977);
nor U22415 (N_22415,N_18795,N_19705);
or U22416 (N_22416,N_19499,N_21306);
xor U22417 (N_22417,N_19182,N_18815);
xnor U22418 (N_22418,N_19282,N_21759);
nand U22419 (N_22419,N_18931,N_19314);
xor U22420 (N_22420,N_19450,N_19223);
or U22421 (N_22421,N_20361,N_19066);
nand U22422 (N_22422,N_21479,N_19696);
nor U22423 (N_22423,N_21388,N_19333);
and U22424 (N_22424,N_19013,N_21816);
nor U22425 (N_22425,N_19140,N_20979);
and U22426 (N_22426,N_19784,N_21290);
or U22427 (N_22427,N_19361,N_19180);
or U22428 (N_22428,N_19685,N_21143);
and U22429 (N_22429,N_20328,N_19743);
and U22430 (N_22430,N_21063,N_19139);
nand U22431 (N_22431,N_18787,N_20069);
nor U22432 (N_22432,N_21752,N_19508);
nand U22433 (N_22433,N_19924,N_19577);
and U22434 (N_22434,N_21175,N_20531);
nand U22435 (N_22435,N_21003,N_18950);
nand U22436 (N_22436,N_20490,N_19626);
nand U22437 (N_22437,N_19344,N_19420);
nand U22438 (N_22438,N_19195,N_19663);
or U22439 (N_22439,N_20978,N_21172);
nor U22440 (N_22440,N_19602,N_20118);
nor U22441 (N_22441,N_20227,N_20735);
or U22442 (N_22442,N_20164,N_19679);
nor U22443 (N_22443,N_19852,N_20285);
nand U22444 (N_22444,N_20466,N_19305);
nand U22445 (N_22445,N_20296,N_19564);
nor U22446 (N_22446,N_21457,N_19222);
xnor U22447 (N_22447,N_18864,N_21381);
and U22448 (N_22448,N_18967,N_19801);
nor U22449 (N_22449,N_21444,N_20219);
xor U22450 (N_22450,N_20938,N_21662);
and U22451 (N_22451,N_18790,N_20271);
xor U22452 (N_22452,N_21617,N_20669);
xnor U22453 (N_22453,N_19944,N_19237);
and U22454 (N_22454,N_19868,N_19600);
xnor U22455 (N_22455,N_21163,N_19288);
nand U22456 (N_22456,N_19840,N_19745);
nor U22457 (N_22457,N_20785,N_19064);
nand U22458 (N_22458,N_20252,N_18819);
nor U22459 (N_22459,N_20713,N_19676);
and U22460 (N_22460,N_19473,N_20453);
nor U22461 (N_22461,N_21166,N_20405);
nand U22462 (N_22462,N_19398,N_20913);
nand U22463 (N_22463,N_19814,N_19969);
and U22464 (N_22464,N_20284,N_19070);
nand U22465 (N_22465,N_21537,N_21860);
or U22466 (N_22466,N_19770,N_20427);
xor U22467 (N_22467,N_19976,N_20728);
xor U22468 (N_22468,N_19385,N_20179);
or U22469 (N_22469,N_21035,N_19512);
nor U22470 (N_22470,N_21401,N_21707);
or U22471 (N_22471,N_18858,N_21683);
or U22472 (N_22472,N_19390,N_20563);
xnor U22473 (N_22473,N_19535,N_18973);
or U22474 (N_22474,N_19416,N_19045);
nand U22475 (N_22475,N_19117,N_21771);
xnor U22476 (N_22476,N_19012,N_19566);
or U22477 (N_22477,N_21413,N_19979);
or U22478 (N_22478,N_20796,N_21174);
or U22479 (N_22479,N_20711,N_20137);
xor U22480 (N_22480,N_19707,N_19682);
xor U22481 (N_22481,N_21826,N_20901);
and U22482 (N_22482,N_19301,N_19170);
nand U22483 (N_22483,N_18895,N_18959);
and U22484 (N_22484,N_19103,N_21318);
or U22485 (N_22485,N_20980,N_19253);
xnor U22486 (N_22486,N_20589,N_21573);
xor U22487 (N_22487,N_19885,N_20232);
and U22488 (N_22488,N_21259,N_20780);
or U22489 (N_22489,N_20408,N_19492);
and U22490 (N_22490,N_19186,N_20385);
xnor U22491 (N_22491,N_21322,N_20197);
and U22492 (N_22492,N_19953,N_19948);
xor U22493 (N_22493,N_19752,N_20637);
nor U22494 (N_22494,N_20229,N_20495);
or U22495 (N_22495,N_21605,N_21478);
nand U22496 (N_22496,N_21517,N_20943);
or U22497 (N_22497,N_21243,N_18920);
nor U22498 (N_22498,N_20506,N_20671);
xor U22499 (N_22499,N_19409,N_19960);
nand U22500 (N_22500,N_21649,N_21503);
or U22501 (N_22501,N_19037,N_20956);
and U22502 (N_22502,N_21051,N_21181);
and U22503 (N_22503,N_21443,N_19262);
nand U22504 (N_22504,N_19629,N_21614);
xnor U22505 (N_22505,N_19310,N_19019);
xnor U22506 (N_22506,N_21822,N_21718);
and U22507 (N_22507,N_20107,N_19453);
xnor U22508 (N_22508,N_20206,N_20298);
nand U22509 (N_22509,N_18910,N_20489);
and U22510 (N_22510,N_21465,N_20304);
and U22511 (N_22511,N_21735,N_18841);
or U22512 (N_22512,N_19126,N_19599);
nor U22513 (N_22513,N_20630,N_18951);
and U22514 (N_22514,N_20792,N_19590);
xor U22515 (N_22515,N_21592,N_21681);
or U22516 (N_22516,N_21580,N_20973);
nand U22517 (N_22517,N_21792,N_21151);
and U22518 (N_22518,N_19065,N_21805);
xor U22519 (N_22519,N_20986,N_20098);
and U22520 (N_22520,N_21853,N_18948);
nand U22521 (N_22521,N_21336,N_21847);
or U22522 (N_22522,N_21300,N_19440);
nor U22523 (N_22523,N_19163,N_21486);
or U22524 (N_22524,N_21748,N_21214);
or U22525 (N_22525,N_20603,N_20275);
or U22526 (N_22526,N_21131,N_21254);
nor U22527 (N_22527,N_21729,N_19125);
nor U22528 (N_22528,N_19407,N_21558);
nor U22529 (N_22529,N_18911,N_19631);
xnor U22530 (N_22530,N_19798,N_18985);
or U22531 (N_22531,N_19430,N_18873);
nand U22532 (N_22532,N_18837,N_21006);
or U22533 (N_22533,N_19005,N_20649);
and U22534 (N_22534,N_19068,N_18800);
xnor U22535 (N_22535,N_19121,N_19772);
or U22536 (N_22536,N_20699,N_19145);
or U22537 (N_22537,N_21025,N_19551);
nor U22538 (N_22538,N_18785,N_21687);
or U22539 (N_22539,N_20533,N_19408);
or U22540 (N_22540,N_20667,N_20481);
or U22541 (N_22541,N_20633,N_20140);
nand U22542 (N_22542,N_21526,N_19325);
and U22543 (N_22543,N_20645,N_19580);
or U22544 (N_22544,N_20878,N_19270);
or U22545 (N_22545,N_19978,N_20714);
nor U22546 (N_22546,N_19831,N_20230);
nand U22547 (N_22547,N_21642,N_21476);
xnor U22548 (N_22548,N_21730,N_19498);
xor U22549 (N_22549,N_21470,N_18776);
xnor U22550 (N_22550,N_19114,N_19083);
and U22551 (N_22551,N_21468,N_19274);
or U22552 (N_22552,N_20439,N_21523);
nand U22553 (N_22553,N_20462,N_18773);
and U22554 (N_22554,N_19716,N_19095);
and U22555 (N_22555,N_21056,N_21395);
nand U22556 (N_22556,N_21835,N_20335);
nor U22557 (N_22557,N_19641,N_19029);
nand U22558 (N_22558,N_18827,N_19319);
and U22559 (N_22559,N_20092,N_19957);
nor U22560 (N_22560,N_19122,N_21680);
nand U22561 (N_22561,N_20750,N_21507);
nand U22562 (N_22562,N_21256,N_19725);
and U22563 (N_22563,N_19972,N_19827);
xnor U22564 (N_22564,N_20131,N_21071);
nand U22565 (N_22565,N_21428,N_20833);
and U22566 (N_22566,N_21596,N_20483);
nand U22567 (N_22567,N_20200,N_19166);
xnor U22568 (N_22568,N_21432,N_21551);
xor U22569 (N_22569,N_20044,N_19732);
and U22570 (N_22570,N_20550,N_21458);
or U22571 (N_22571,N_19173,N_19384);
nand U22572 (N_22572,N_20492,N_19468);
or U22573 (N_22573,N_19952,N_19136);
or U22574 (N_22574,N_19119,N_20316);
nand U22575 (N_22575,N_20182,N_21521);
xor U22576 (N_22576,N_21870,N_21070);
and U22577 (N_22577,N_21371,N_20974);
nor U22578 (N_22578,N_20166,N_19936);
nor U22579 (N_22579,N_19187,N_20080);
nor U22580 (N_22580,N_19706,N_18861);
nor U22581 (N_22581,N_20753,N_18863);
nand U22582 (N_22582,N_21195,N_19853);
and U22583 (N_22583,N_19109,N_18907);
nor U22584 (N_22584,N_18947,N_19824);
or U22585 (N_22585,N_20384,N_20996);
and U22586 (N_22586,N_18824,N_19234);
nor U22587 (N_22587,N_20141,N_19185);
nor U22588 (N_22588,N_20281,N_21864);
nor U22589 (N_22589,N_20337,N_20717);
xor U22590 (N_22590,N_19795,N_21645);
or U22591 (N_22591,N_20187,N_20881);
and U22592 (N_22592,N_19160,N_21471);
nor U22593 (N_22593,N_20241,N_21584);
nor U22594 (N_22594,N_20613,N_21777);
nor U22595 (N_22595,N_20162,N_20248);
nand U22596 (N_22596,N_20465,N_20193);
or U22597 (N_22597,N_20816,N_21682);
xor U22598 (N_22598,N_19502,N_20297);
or U22599 (N_22599,N_20763,N_20959);
nor U22600 (N_22600,N_20435,N_19322);
and U22601 (N_22601,N_21820,N_20456);
and U22602 (N_22602,N_18899,N_21838);
and U22603 (N_22603,N_20544,N_20242);
and U22604 (N_22604,N_20848,N_19536);
or U22605 (N_22605,N_20156,N_20969);
nand U22606 (N_22606,N_21654,N_20160);
xnor U22607 (N_22607,N_20478,N_19079);
and U22608 (N_22608,N_19864,N_20580);
nor U22609 (N_22609,N_21779,N_19309);
nor U22610 (N_22610,N_19230,N_21170);
xor U22611 (N_22611,N_20031,N_20381);
xor U22612 (N_22612,N_21029,N_21383);
and U22613 (N_22613,N_19905,N_20517);
xor U22614 (N_22614,N_21671,N_20086);
xor U22615 (N_22615,N_21342,N_20195);
and U22616 (N_22616,N_20186,N_19299);
xor U22617 (N_22617,N_21774,N_21012);
or U22618 (N_22618,N_20503,N_19466);
xnor U22619 (N_22619,N_19856,N_21693);
xor U22620 (N_22620,N_21768,N_19073);
nand U22621 (N_22621,N_20657,N_20174);
and U22622 (N_22622,N_19818,N_20602);
nand U22623 (N_22623,N_18994,N_19008);
nor U22624 (N_22624,N_19264,N_19739);
xor U22625 (N_22625,N_20842,N_21201);
nor U22626 (N_22626,N_19201,N_18921);
and U22627 (N_22627,N_20862,N_20070);
xor U22628 (N_22628,N_19834,N_19422);
nand U22629 (N_22629,N_19482,N_20522);
nor U22630 (N_22630,N_20982,N_20269);
nand U22631 (N_22631,N_18828,N_18814);
nand U22632 (N_22632,N_20829,N_19554);
xor U22633 (N_22633,N_20819,N_20006);
or U22634 (N_22634,N_19591,N_19563);
xor U22635 (N_22635,N_18914,N_18845);
xnor U22636 (N_22636,N_20634,N_21505);
or U22637 (N_22637,N_20523,N_19249);
xnor U22638 (N_22638,N_20760,N_20420);
xnor U22639 (N_22639,N_19561,N_21358);
nor U22640 (N_22640,N_21008,N_20859);
nor U22641 (N_22641,N_19998,N_20181);
xnor U22642 (N_22642,N_18922,N_21702);
and U22643 (N_22643,N_19134,N_18917);
nor U22644 (N_22644,N_19970,N_20374);
nand U22645 (N_22645,N_21491,N_21832);
nor U22646 (N_22646,N_20096,N_21713);
or U22647 (N_22647,N_21146,N_20513);
nand U22648 (N_22648,N_18831,N_20055);
nor U22649 (N_22649,N_19245,N_19883);
nand U22650 (N_22650,N_18999,N_21704);
nor U22651 (N_22651,N_20689,N_21082);
nand U22652 (N_22652,N_21817,N_19478);
or U22653 (N_22653,N_20053,N_21399);
nand U22654 (N_22654,N_20432,N_21048);
xor U22655 (N_22655,N_21571,N_20850);
or U22656 (N_22656,N_21073,N_19722);
and U22657 (N_22657,N_21634,N_21149);
or U22658 (N_22658,N_21111,N_21467);
or U22659 (N_22659,N_19263,N_21866);
xor U22660 (N_22660,N_21324,N_21756);
or U22661 (N_22661,N_21075,N_21335);
and U22662 (N_22662,N_20970,N_21031);
xor U22663 (N_22663,N_18925,N_19042);
xnor U22664 (N_22664,N_21072,N_21049);
or U22665 (N_22665,N_21791,N_20282);
and U22666 (N_22666,N_21103,N_19391);
and U22667 (N_22667,N_19579,N_19928);
nand U22668 (N_22668,N_19758,N_21041);
nand U22669 (N_22669,N_21794,N_19887);
and U22670 (N_22670,N_21098,N_19985);
nand U22671 (N_22671,N_19847,N_21750);
or U22672 (N_22672,N_20571,N_20349);
nor U22673 (N_22673,N_18918,N_21732);
nor U22674 (N_22674,N_20681,N_20371);
nor U22675 (N_22675,N_20741,N_19908);
and U22676 (N_22676,N_21262,N_21525);
or U22677 (N_22677,N_19243,N_19352);
nor U22678 (N_22678,N_18855,N_19159);
and U22679 (N_22679,N_19898,N_20032);
and U22680 (N_22680,N_21229,N_20838);
xnor U22681 (N_22681,N_19774,N_20303);
nor U22682 (N_22682,N_19892,N_21059);
and U22683 (N_22683,N_20870,N_19785);
and U22684 (N_22684,N_20075,N_21240);
xnor U22685 (N_22685,N_20595,N_20632);
nand U22686 (N_22686,N_21593,N_19559);
and U22687 (N_22687,N_18874,N_20840);
nor U22688 (N_22688,N_18885,N_19190);
or U22689 (N_22689,N_19089,N_21688);
or U22690 (N_22690,N_20590,N_19093);
nand U22691 (N_22691,N_19904,N_19296);
nand U22692 (N_22692,N_19819,N_20839);
nand U22693 (N_22693,N_20678,N_20356);
nand U22694 (N_22694,N_19690,N_20574);
nand U22695 (N_22695,N_19811,N_20510);
nor U22696 (N_22696,N_20194,N_19286);
xor U22697 (N_22697,N_21141,N_19501);
or U22698 (N_22698,N_21528,N_20748);
xor U22699 (N_22699,N_20917,N_20355);
nor U22700 (N_22700,N_20647,N_20437);
nand U22701 (N_22701,N_20294,N_21804);
xnor U22702 (N_22702,N_19238,N_20376);
xor U22703 (N_22703,N_20587,N_19318);
nor U22704 (N_22704,N_18782,N_19532);
or U22705 (N_22705,N_19740,N_19392);
or U22706 (N_22706,N_21709,N_19436);
xor U22707 (N_22707,N_19704,N_19376);
and U22708 (N_22708,N_20535,N_19545);
or U22709 (N_22709,N_20680,N_20287);
nor U22710 (N_22710,N_20262,N_19653);
xnor U22711 (N_22711,N_18984,N_20611);
and U22712 (N_22712,N_20496,N_19107);
xor U22713 (N_22713,N_21829,N_19826);
nor U22714 (N_22714,N_18817,N_19120);
and U22715 (N_22715,N_21466,N_20899);
and U22716 (N_22716,N_20313,N_19316);
and U22717 (N_22717,N_19043,N_21658);
nor U22718 (N_22718,N_20038,N_21824);
nand U22719 (N_22719,N_21333,N_18902);
nor U22720 (N_22720,N_21245,N_19020);
or U22721 (N_22721,N_20030,N_19861);
nand U22722 (N_22722,N_18980,N_20557);
and U22723 (N_22723,N_20997,N_19915);
nand U22724 (N_22724,N_20827,N_19719);
or U22725 (N_22725,N_20732,N_21463);
xor U22726 (N_22726,N_21869,N_19415);
nand U22727 (N_22727,N_20605,N_20874);
xnor U22728 (N_22728,N_19513,N_20416);
nor U22729 (N_22729,N_20694,N_20089);
or U22730 (N_22730,N_21102,N_21535);
or U22731 (N_22731,N_19359,N_21251);
xnor U22732 (N_22732,N_21117,N_20199);
xor U22733 (N_22733,N_21566,N_19611);
nand U22734 (N_22734,N_19374,N_18752);
nor U22735 (N_22735,N_19321,N_20050);
and U22736 (N_22736,N_21389,N_21190);
nor U22737 (N_22737,N_21270,N_20217);
and U22738 (N_22738,N_20812,N_19754);
and U22739 (N_22739,N_21323,N_20915);
or U22740 (N_22740,N_20063,N_20998);
nand U22741 (N_22741,N_20463,N_19075);
xnor U22742 (N_22742,N_20743,N_21754);
nand U22743 (N_22743,N_19907,N_21325);
xor U22744 (N_22744,N_21552,N_20933);
xor U22745 (N_22745,N_20440,N_21576);
xnor U22746 (N_22746,N_21810,N_19829);
xnor U22747 (N_22747,N_19147,N_21162);
and U22748 (N_22748,N_21400,N_21607);
or U22749 (N_22749,N_19698,N_21173);
and U22750 (N_22750,N_21628,N_19612);
nand U22751 (N_22751,N_19639,N_20012);
nand U22752 (N_22752,N_19183,N_20851);
xor U22753 (N_22753,N_20946,N_20515);
nand U22754 (N_22754,N_21047,N_20924);
or U22755 (N_22755,N_19654,N_19331);
nand U22756 (N_22756,N_20835,N_20610);
or U22757 (N_22757,N_20821,N_20188);
or U22758 (N_22758,N_21689,N_19273);
nor U22759 (N_22759,N_20320,N_20811);
and U22760 (N_22760,N_20212,N_19366);
nor U22761 (N_22761,N_19338,N_19025);
xor U22762 (N_22762,N_19097,N_21147);
and U22763 (N_22763,N_21104,N_21372);
nand U22764 (N_22764,N_21723,N_21613);
nor U22765 (N_22765,N_20808,N_20659);
or U22766 (N_22766,N_19060,N_21406);
nor U22767 (N_22767,N_20054,N_18913);
nor U22768 (N_22768,N_19151,N_20014);
nor U22769 (N_22769,N_18893,N_19176);
or U22770 (N_22770,N_21279,N_21348);
nor U22771 (N_22771,N_19660,N_20810);
and U22772 (N_22772,N_20509,N_20756);
nor U22773 (N_22773,N_19221,N_18906);
and U22774 (N_22774,N_20772,N_19980);
and U22775 (N_22775,N_20655,N_19646);
and U22776 (N_22776,N_20302,N_20967);
or U22777 (N_22777,N_20947,N_18767);
nand U22778 (N_22778,N_19001,N_19472);
or U22779 (N_22779,N_20706,N_20247);
or U22780 (N_22780,N_21795,N_20001);
nand U22781 (N_22781,N_19917,N_21589);
nand U22782 (N_22782,N_19622,N_20369);
or U22783 (N_22783,N_19135,N_21242);
xor U22784 (N_22784,N_19271,N_20238);
and U22785 (N_22785,N_19703,N_20628);
xnor U22786 (N_22786,N_19912,N_20558);
and U22787 (N_22787,N_20985,N_19876);
xor U22788 (N_22788,N_19490,N_19963);
and U22789 (N_22789,N_19937,N_19872);
nand U22790 (N_22790,N_21851,N_19863);
nand U22791 (N_22791,N_21610,N_19721);
and U22792 (N_22792,N_21764,N_20793);
and U22793 (N_22793,N_19014,N_20567);
xnor U22794 (N_22794,N_18867,N_19817);
and U22795 (N_22795,N_19804,N_20745);
or U22796 (N_22796,N_19807,N_18821);
and U22797 (N_22797,N_20438,N_19315);
xnor U22798 (N_22798,N_19881,N_20144);
nor U22799 (N_22799,N_19219,N_18971);
nand U22800 (N_22800,N_18944,N_21161);
nor U22801 (N_22801,N_20132,N_20928);
nand U22802 (N_22802,N_18849,N_18935);
or U22803 (N_22803,N_21360,N_19494);
nor U22804 (N_22804,N_21621,N_21200);
xor U22805 (N_22805,N_21679,N_19664);
or U22806 (N_22806,N_18859,N_19888);
and U22807 (N_22807,N_21561,N_19768);
or U22808 (N_22808,N_20314,N_18807);
nor U22809 (N_22809,N_20170,N_19056);
nor U22810 (N_22810,N_21445,N_19445);
xnor U22811 (N_22811,N_21191,N_20552);
xor U22812 (N_22812,N_19347,N_21158);
or U22813 (N_22813,N_21359,N_21821);
and U22814 (N_22814,N_19454,N_21039);
nor U22815 (N_22815,N_18865,N_20579);
nand U22816 (N_22816,N_20886,N_20426);
and U22817 (N_22817,N_21594,N_19967);
xor U22818 (N_22818,N_21807,N_20770);
or U22819 (N_22819,N_18834,N_19053);
nand U22820 (N_22820,N_20941,N_18793);
and U22821 (N_22821,N_20940,N_21312);
or U22822 (N_22822,N_19389,N_19897);
nand U22823 (N_22823,N_20788,N_19010);
nor U22824 (N_22824,N_19277,N_19152);
nand U22825 (N_22825,N_18759,N_19674);
or U22826 (N_22826,N_20469,N_19576);
nor U22827 (N_22827,N_18788,N_21751);
xor U22828 (N_22828,N_20868,N_20726);
or U22829 (N_22829,N_21728,N_20646);
nor U22830 (N_22830,N_20930,N_21116);
or U22831 (N_22831,N_18801,N_19608);
and U22832 (N_22832,N_20737,N_19158);
and U22833 (N_22833,N_19910,N_19295);
xor U22834 (N_22834,N_20290,N_19850);
or U22835 (N_22835,N_21506,N_21660);
and U22836 (N_22836,N_18909,N_21686);
or U22837 (N_22837,N_19203,N_20067);
nand U22838 (N_22838,N_19130,N_19062);
nor U22839 (N_22839,N_18765,N_18860);
nor U22840 (N_22840,N_18905,N_18857);
nand U22841 (N_22841,N_21657,N_20482);
nor U22842 (N_22842,N_18783,N_19138);
and U22843 (N_22843,N_19585,N_20730);
or U22844 (N_22844,N_21150,N_20551);
nor U22845 (N_22845,N_19935,N_20890);
xnor U22846 (N_22846,N_19346,N_20393);
and U22847 (N_22847,N_20234,N_21209);
nand U22848 (N_22848,N_20346,N_19675);
xnor U22849 (N_22849,N_21536,N_21839);
xor U22850 (N_22850,N_21124,N_21738);
or U22851 (N_22851,N_19941,N_21193);
nand U22852 (N_22852,N_19934,N_21871);
xnor U22853 (N_22853,N_20367,N_19806);
xor U22854 (N_22854,N_21666,N_21442);
nor U22855 (N_22855,N_20958,N_19447);
nand U22856 (N_22856,N_19087,N_21724);
and U22857 (N_22857,N_21530,N_20493);
and U22858 (N_22858,N_20889,N_21441);
xor U22859 (N_22859,N_19485,N_21298);
and U22860 (N_22860,N_21213,N_20323);
nor U22861 (N_22861,N_21780,N_19329);
and U22862 (N_22862,N_18908,N_21494);
or U22863 (N_22863,N_21407,N_19738);
nand U22864 (N_22864,N_20636,N_18804);
or U22865 (N_22865,N_18878,N_19444);
nand U22866 (N_22866,N_19032,N_21460);
xnor U22867 (N_22867,N_19880,N_18850);
nand U22868 (N_22868,N_19517,N_20126);
and U22869 (N_22869,N_19377,N_20033);
or U22870 (N_22870,N_20638,N_19133);
or U22871 (N_22871,N_20834,N_20321);
or U22872 (N_22872,N_18888,N_19765);
or U22873 (N_22873,N_20273,N_21084);
nor U22874 (N_22874,N_18889,N_20872);
xor U22875 (N_22875,N_21261,N_19402);
nor U22876 (N_22876,N_20715,N_20042);
and U22877 (N_22877,N_21731,N_21160);
and U22878 (N_22878,N_21859,N_19340);
or U22879 (N_22879,N_20412,N_20283);
nand U22880 (N_22880,N_21274,N_19100);
nor U22881 (N_22881,N_21036,N_20900);
or U22882 (N_22882,N_19637,N_19878);
xor U22883 (N_22883,N_21714,N_21564);
nor U22884 (N_22884,N_19251,N_20288);
nor U22885 (N_22885,N_19583,N_20454);
xor U22886 (N_22886,N_19365,N_21299);
and U22887 (N_22887,N_19054,N_21030);
and U22888 (N_22888,N_19596,N_20707);
nand U22889 (N_22889,N_20778,N_19546);
nor U22890 (N_22890,N_18868,N_20541);
and U22891 (N_22891,N_20919,N_19975);
and U22892 (N_22892,N_19879,N_19205);
xor U22893 (N_22893,N_20344,N_21874);
nand U22894 (N_22894,N_18823,N_20679);
nand U22895 (N_22895,N_19723,N_21435);
nor U22896 (N_22896,N_21578,N_19153);
nand U22897 (N_22897,N_20317,N_19762);
or U22898 (N_22898,N_20846,N_21480);
or U22899 (N_22899,N_19573,N_18979);
and U22900 (N_22900,N_18983,N_19712);
nand U22901 (N_22901,N_19670,N_21518);
or U22902 (N_22902,N_18958,N_20572);
and U22903 (N_22903,N_21675,N_20370);
and U22904 (N_22904,N_18934,N_21497);
and U22905 (N_22905,N_19480,N_20480);
or U22906 (N_22906,N_21553,N_20939);
and U22907 (N_22907,N_21798,N_21114);
nand U22908 (N_22908,N_21565,N_20036);
nand U22909 (N_22909,N_21760,N_19092);
nand U22910 (N_22910,N_20122,N_20318);
or U22911 (N_22911,N_18832,N_20348);
xnor U22912 (N_22912,N_20575,N_20159);
xnor U22913 (N_22913,N_19039,N_20716);
or U22914 (N_22914,N_19543,N_19891);
and U22915 (N_22915,N_19265,N_21410);
or U22916 (N_22916,N_21533,N_18960);
nor U22917 (N_22917,N_19899,N_21386);
and U22918 (N_22918,N_20270,N_18876);
xor U22919 (N_22919,N_18927,N_19990);
nand U22920 (N_22920,N_20431,N_21273);
and U22921 (N_22921,N_19157,N_21167);
or U22922 (N_22922,N_21512,N_19168);
or U22923 (N_22923,N_21765,N_19423);
nor U22924 (N_22924,N_19896,N_19710);
nand U22925 (N_22925,N_20378,N_21380);
nand U22926 (N_22926,N_19046,N_20245);
nand U22927 (N_22927,N_21667,N_19200);
nor U22928 (N_22928,N_20085,N_19193);
xnor U22929 (N_22929,N_19800,N_21067);
and U22930 (N_22930,N_21384,N_18919);
or U22931 (N_22931,N_19742,N_20814);
and U22932 (N_22932,N_19207,N_19484);
nor U22933 (N_22933,N_20147,N_19381);
nor U22934 (N_22934,N_21080,N_20799);
and U22935 (N_22935,N_21309,N_19248);
or U22936 (N_22936,N_19781,N_21665);
nor U22937 (N_22937,N_21744,N_19489);
and U22938 (N_22938,N_21018,N_21474);
xor U22939 (N_22939,N_20450,N_21762);
nand U22940 (N_22940,N_20858,N_19078);
nor U22941 (N_22941,N_20326,N_21007);
nand U22942 (N_22942,N_19052,N_21749);
and U22943 (N_22943,N_21328,N_18846);
nor U22944 (N_22944,N_20813,N_18879);
nand U22945 (N_22945,N_21013,N_21286);
nor U22946 (N_22946,N_19607,N_21575);
nand U22947 (N_22947,N_19306,N_19364);
xnor U22948 (N_22948,N_20764,N_21532);
nand U22949 (N_22949,N_18904,N_21745);
and U22950 (N_22950,N_19531,N_20887);
or U22951 (N_22951,N_21231,N_19552);
xor U22952 (N_22952,N_19388,N_21317);
nor U22953 (N_22953,N_20776,N_21096);
or U22954 (N_22954,N_20936,N_20139);
nand U22955 (N_22955,N_20258,N_21219);
or U22956 (N_22956,N_20312,N_19982);
xnor U22957 (N_22957,N_21089,N_19755);
nand U22958 (N_22958,N_19727,N_19399);
nand U22959 (N_22959,N_21743,N_19658);
or U22960 (N_22960,N_21761,N_21394);
or U22961 (N_22961,N_21267,N_21028);
nor U22962 (N_22962,N_20892,N_20653);
and U22963 (N_22963,N_19668,N_20806);
nand U22964 (N_22964,N_20025,N_20390);
nor U22965 (N_22965,N_21747,N_18830);
and U22966 (N_22966,N_20157,N_19744);
nand U22967 (N_22967,N_20584,N_19515);
and U22968 (N_22968,N_21228,N_20951);
nor U22969 (N_22969,N_21094,N_20037);
nor U22970 (N_22970,N_20891,N_20525);
nand U22971 (N_22971,N_21307,N_20542);
xnor U22972 (N_22972,N_19731,N_21630);
or U22973 (N_22973,N_19930,N_21590);
and U22974 (N_22974,N_20051,N_19839);
and U22975 (N_22975,N_20169,N_20757);
nor U22976 (N_22976,N_19902,N_19510);
or U22977 (N_22977,N_21119,N_20165);
nand U22978 (N_22978,N_21484,N_21338);
xnor U22979 (N_22979,N_21220,N_20554);
xor U22980 (N_22980,N_18753,N_19757);
or U22981 (N_22981,N_21027,N_21733);
nor U22982 (N_22982,N_20747,N_20962);
xor U22983 (N_22983,N_20024,N_21844);
and U22984 (N_22984,N_20582,N_21354);
xnor U22985 (N_22985,N_19475,N_20824);
nand U22986 (N_22986,N_18896,N_19813);
nor U22987 (N_22987,N_18998,N_20591);
and U22988 (N_22988,N_18970,N_18768);
xor U22989 (N_22989,N_20950,N_19216);
nand U22990 (N_22990,N_20289,N_20616);
or U22991 (N_22991,N_19240,N_21367);
xnor U22992 (N_22992,N_18955,N_19617);
and U22993 (N_22993,N_20841,N_20362);
xor U22994 (N_22994,N_21716,N_20545);
nor U22995 (N_22995,N_21715,N_19869);
nand U22996 (N_22996,N_18803,N_19113);
xor U22997 (N_22997,N_20173,N_20976);
and U22998 (N_22998,N_21640,N_20594);
or U22999 (N_22999,N_20733,N_19949);
nand U23000 (N_23000,N_20549,N_19267);
nor U23001 (N_23001,N_21337,N_21069);
nor U23002 (N_23002,N_21635,N_21344);
or U23003 (N_23003,N_19933,N_18791);
or U23004 (N_23004,N_18771,N_20153);
or U23005 (N_23005,N_20508,N_20046);
xnor U23006 (N_23006,N_20598,N_18750);
and U23007 (N_23007,N_20340,N_21815);
nand U23008 (N_23008,N_19028,N_21755);
nand U23009 (N_23009,N_19749,N_19302);
or U23010 (N_23010,N_20152,N_18755);
or U23011 (N_23011,N_18762,N_19382);
nand U23012 (N_23012,N_20803,N_19521);
nor U23013 (N_23013,N_21706,N_20992);
or U23014 (N_23014,N_21155,N_20472);
xnor U23015 (N_23015,N_19049,N_19616);
xnor U23016 (N_23016,N_21023,N_19918);
nor U23017 (N_23017,N_19572,N_19981);
xor U23018 (N_23018,N_21440,N_20642);
nand U23019 (N_23019,N_21127,N_18848);
xnor U23020 (N_23020,N_21672,N_20116);
nand U23021 (N_23021,N_21475,N_20845);
nand U23022 (N_23022,N_21490,N_20984);
nor U23023 (N_23023,N_19403,N_19962);
nand U23024 (N_23024,N_20175,N_21115);
or U23025 (N_23025,N_21570,N_18883);
and U23026 (N_23026,N_19776,N_19959);
xor U23027 (N_23027,N_21452,N_19808);
xnor U23028 (N_23028,N_20204,N_20777);
or U23029 (N_23029,N_18891,N_20720);
and U23030 (N_23030,N_19146,N_21153);
and U23031 (N_23031,N_19311,N_19339);
and U23032 (N_23032,N_19463,N_21769);
or U23033 (N_23033,N_19822,N_21808);
nor U23034 (N_23034,N_21044,N_19348);
nand U23035 (N_23035,N_21546,N_19281);
and U23036 (N_23036,N_20783,N_21278);
nand U23037 (N_23037,N_18769,N_21266);
and U23038 (N_23038,N_20701,N_20305);
nand U23039 (N_23039,N_20231,N_21126);
or U23040 (N_23040,N_20015,N_19825);
and U23041 (N_23041,N_20442,N_20990);
nor U23042 (N_23042,N_20072,N_20652);
xor U23043 (N_23043,N_20625,N_19246);
and U23044 (N_23044,N_20103,N_21850);
or U23045 (N_23045,N_21763,N_20299);
nor U23046 (N_23046,N_20315,N_21296);
or U23047 (N_23047,N_18940,N_20972);
nor U23048 (N_23048,N_19848,N_21361);
or U23049 (N_23049,N_20257,N_19162);
nand U23050 (N_23050,N_19511,N_20295);
nor U23051 (N_23051,N_19076,N_20561);
nand U23052 (N_23052,N_19007,N_19718);
nor U23053 (N_23053,N_21496,N_21684);
xnor U23054 (N_23054,N_21623,N_20519);
and U23055 (N_23055,N_20148,N_19343);
and U23056 (N_23056,N_20620,N_20377);
and U23057 (N_23057,N_19523,N_20823);
xnor U23058 (N_23058,N_19550,N_21142);
nand U23059 (N_23059,N_21834,N_19451);
nor U23060 (N_23060,N_19197,N_18872);
and U23061 (N_23061,N_19149,N_19000);
nor U23062 (N_23062,N_21547,N_21631);
and U23063 (N_23063,N_20324,N_19609);
nand U23064 (N_23064,N_20588,N_20358);
xnor U23065 (N_23065,N_21009,N_19362);
and U23066 (N_23066,N_19441,N_20497);
or U23067 (N_23067,N_21288,N_21852);
and U23068 (N_23068,N_19257,N_19424);
nand U23069 (N_23069,N_18806,N_21037);
nor U23070 (N_23070,N_20817,N_20041);
nand U23071 (N_23071,N_21451,N_20345);
nor U23072 (N_23072,N_20479,N_18952);
nand U23073 (N_23073,N_19350,N_20065);
xnor U23074 (N_23074,N_21424,N_19181);
xor U23075 (N_23075,N_19925,N_21511);
or U23076 (N_23076,N_20873,N_21088);
xor U23077 (N_23077,N_20615,N_19414);
nand U23078 (N_23078,N_19228,N_20624);
nand U23079 (N_23079,N_19890,N_19269);
xor U23080 (N_23080,N_19894,N_19354);
or U23081 (N_23081,N_20977,N_19922);
xnor U23082 (N_23082,N_21563,N_21064);
nor U23083 (N_23083,N_20767,N_19326);
and U23084 (N_23084,N_19224,N_20319);
xnor U23085 (N_23085,N_21618,N_21192);
or U23086 (N_23086,N_19581,N_21184);
and U23087 (N_23087,N_20422,N_21417);
nand U23088 (N_23088,N_20268,N_20161);
xnor U23089 (N_23089,N_20592,N_19217);
and U23090 (N_23090,N_20619,N_18932);
nand U23091 (N_23091,N_18844,N_21611);
or U23092 (N_23092,N_20151,N_20804);
xnor U23093 (N_23093,N_19763,N_19860);
nor U23094 (N_23094,N_21135,N_18763);
xnor U23095 (N_23095,N_21462,N_21079);
xor U23096 (N_23096,N_19137,N_21314);
nand U23097 (N_23097,N_19432,N_20357);
xor U23098 (N_23098,N_20088,N_18774);
or U23099 (N_23099,N_19965,N_19920);
and U23100 (N_23100,N_18887,N_20125);
nor U23101 (N_23101,N_19735,N_21122);
nor U23102 (N_23102,N_21513,N_19997);
nand U23103 (N_23103,N_20049,N_21865);
nor U23104 (N_23104,N_20604,N_20244);
xor U23105 (N_23105,N_19479,N_19413);
xor U23106 (N_23106,N_20425,N_21385);
nand U23107 (N_23107,N_20424,N_19015);
or U23108 (N_23108,N_18751,N_21498);
nand U23109 (N_23109,N_19106,N_19342);
or U23110 (N_23110,N_19597,N_20423);
and U23111 (N_23111,N_21257,N_19194);
xor U23112 (N_23112,N_20073,N_19312);
xnor U23113 (N_23113,N_20762,N_19603);
and U23114 (N_23114,N_21110,N_19560);
and U23115 (N_23115,N_20547,N_19956);
nand U23116 (N_23116,N_20221,N_21331);
or U23117 (N_23117,N_19255,N_21210);
or U23118 (N_23118,N_21625,N_20090);
nand U23119 (N_23119,N_19964,N_21313);
or U23120 (N_23120,N_21364,N_21472);
and U23121 (N_23121,N_19659,N_19009);
and U23122 (N_23122,N_21837,N_21377);
or U23123 (N_23123,N_21362,N_21236);
nand U23124 (N_23124,N_19812,N_21694);
xor U23125 (N_23125,N_19514,N_18956);
nand U23126 (N_23126,N_20885,N_21137);
and U23127 (N_23127,N_19421,N_19433);
or U23128 (N_23128,N_21519,N_21097);
or U23129 (N_23129,N_21002,N_19428);
and U23130 (N_23130,N_20836,N_19394);
nand U23131 (N_23131,N_18988,N_21500);
nor U23132 (N_23132,N_21434,N_20329);
nand U23133 (N_23133,N_21606,N_20909);
and U23134 (N_23134,N_21224,N_19909);
or U23135 (N_23135,N_19540,N_20213);
nor U23136 (N_23136,N_19341,N_21087);
xnor U23137 (N_23137,N_20690,N_19627);
and U23138 (N_23138,N_21464,N_20693);
xnor U23139 (N_23139,N_21378,N_20468);
xnor U23140 (N_23140,N_21345,N_19123);
xnor U23141 (N_23141,N_20458,N_19926);
nor U23142 (N_23142,N_18997,N_21356);
or U23143 (N_23143,N_21320,N_20877);
or U23144 (N_23144,N_20018,N_19260);
and U23145 (N_23145,N_21271,N_21397);
nand U23146 (N_23146,N_20286,N_20528);
nor U23147 (N_23147,N_21091,N_19493);
nand U23148 (N_23148,N_20101,N_20192);
xnor U23149 (N_23149,N_20261,N_20322);
and U23150 (N_23150,N_21741,N_19412);
nor U23151 (N_23151,N_21346,N_21349);
and U23152 (N_23152,N_21849,N_20383);
nand U23153 (N_23153,N_18852,N_20964);
xor U23154 (N_23154,N_19071,N_21567);
xnor U23155 (N_23155,N_20135,N_19662);
and U23156 (N_23156,N_20712,N_19794);
and U23157 (N_23157,N_21134,N_20292);
and U23158 (N_23158,N_21276,N_20828);
or U23159 (N_23159,N_20779,N_19683);
nor U23160 (N_23160,N_20907,N_20026);
nor U23161 (N_23161,N_20656,N_18976);
or U23162 (N_23162,N_20975,N_20782);
and U23163 (N_23163,N_20514,N_21569);
xnor U23164 (N_23164,N_21721,N_18926);
or U23165 (N_23165,N_21083,N_19369);
xor U23166 (N_23166,N_20758,N_18901);
or U23167 (N_23167,N_20593,N_20389);
nor U23168 (N_23168,N_19943,N_21691);
nand U23169 (N_23169,N_18797,N_21001);
or U23170 (N_23170,N_19244,N_21854);
or U23171 (N_23171,N_19425,N_21685);
nor U23172 (N_23172,N_21739,N_20790);
or U23173 (N_23173,N_21776,N_20334);
or U23174 (N_23174,N_20511,N_20622);
nand U23175 (N_23175,N_20944,N_19419);
xor U23176 (N_23176,N_21108,N_20207);
or U23177 (N_23177,N_19208,N_21225);
nand U23178 (N_23178,N_19285,N_19734);
xnor U23179 (N_23179,N_20740,N_19437);
or U23180 (N_23180,N_21054,N_19258);
xnor U23181 (N_23181,N_21204,N_19991);
or U23182 (N_23182,N_21040,N_19791);
xor U23183 (N_23183,N_19836,N_19108);
nand U23184 (N_23184,N_19961,N_21061);
nand U23185 (N_23185,N_19854,N_20350);
and U23186 (N_23186,N_19373,N_19588);
nor U23187 (N_23187,N_19686,N_20905);
nor U23188 (N_23188,N_18975,N_19034);
and U23189 (N_23189,N_21226,N_18809);
nand U23190 (N_23190,N_20149,N_19220);
and U23191 (N_23191,N_19225,N_20995);
xor U23192 (N_23192,N_19620,N_21862);
xnor U23193 (N_23193,N_20965,N_21330);
xnor U23194 (N_23194,N_18808,N_18798);
nand U23195 (N_23195,N_19308,N_20576);
and U23196 (N_23196,N_19320,N_20949);
and U23197 (N_23197,N_18794,N_21651);
xnor U23198 (N_23198,N_20347,N_20124);
or U23199 (N_23199,N_21782,N_19105);
xor U23200 (N_23200,N_20863,N_20009);
and U23201 (N_23201,N_21264,N_18880);
nor U23202 (N_23202,N_20787,N_21100);
nand U23203 (N_23203,N_21005,N_18993);
or U23204 (N_23204,N_21588,N_19555);
nor U23205 (N_23205,N_20403,N_19802);
nor U23206 (N_23206,N_20775,N_20664);
xnor U23207 (N_23207,N_20239,N_20455);
nand U23208 (N_23208,N_18757,N_21504);
and U23209 (N_23209,N_20059,N_21129);
or U23210 (N_23210,N_20708,N_21099);
and U23211 (N_23211,N_21232,N_20457);
or U23212 (N_23212,N_19741,N_20183);
nand U23213 (N_23213,N_20061,N_21154);
and U23214 (N_23214,N_19379,N_19469);
nand U23215 (N_23215,N_19417,N_21032);
nand U23216 (N_23216,N_21436,N_19096);
nor U23217 (N_23217,N_19337,N_20082);
xor U23218 (N_23218,N_20914,N_20852);
nor U23219 (N_23219,N_21469,N_21582);
or U23220 (N_23220,N_21130,N_20155);
nor U23221 (N_23221,N_19292,N_21248);
xnor U23222 (N_23222,N_19497,N_19815);
xnor U23223 (N_23223,N_19448,N_19989);
nor U23224 (N_23224,N_20264,N_20112);
xor U23225 (N_23225,N_19184,N_20311);
nor U23226 (N_23226,N_20202,N_18949);
xnor U23227 (N_23227,N_20894,N_20752);
or U23228 (N_23228,N_20529,N_21327);
nand U23229 (N_23229,N_19452,N_19259);
nor U23230 (N_23230,N_20882,N_21321);
nor U23231 (N_23231,N_18957,N_20643);
nor U23232 (N_23232,N_19250,N_20578);
nand U23233 (N_23233,N_20527,N_20240);
nand U23234 (N_23234,N_21633,N_21176);
nor U23235 (N_23235,N_19266,N_19289);
and U23236 (N_23236,N_19730,N_20586);
and U23237 (N_23237,N_20818,N_19858);
nand U23238 (N_23238,N_20379,N_21550);
or U23239 (N_23239,N_21722,N_20300);
nand U23240 (N_23240,N_19986,N_20354);
xor U23241 (N_23241,N_21004,N_21481);
or U23242 (N_23242,N_21659,N_19865);
xnor U23243 (N_23243,N_20150,N_19048);
nand U23244 (N_23244,N_21620,N_21453);
nor U23245 (N_23245,N_18916,N_18829);
nand U23246 (N_23246,N_20847,N_20968);
xnor U23247 (N_23247,N_19750,N_21068);
and U23248 (N_23248,N_21799,N_21246);
nor U23249 (N_23249,N_21329,N_19229);
nor U23250 (N_23250,N_18890,N_21740);
nand U23251 (N_23251,N_20705,N_19242);
or U23252 (N_23252,N_19210,N_21461);
nand U23253 (N_23253,N_20256,N_21326);
or U23254 (N_23254,N_18779,N_21138);
and U23255 (N_23255,N_20331,N_19996);
or U23256 (N_23256,N_19410,N_19443);
and U23257 (N_23257,N_19565,N_18775);
nor U23258 (N_23258,N_19077,N_19689);
or U23259 (N_23259,N_20411,N_20000);
nor U23260 (N_23260,N_21541,N_20857);
xnor U23261 (N_23261,N_20123,N_19036);
nor U23262 (N_23262,N_18816,N_20658);
and U23263 (N_23263,N_20145,N_20452);
nor U23264 (N_23264,N_20934,N_21053);
nand U23265 (N_23265,N_19527,N_20564);
nor U23266 (N_23266,N_20954,N_19495);
xor U23267 (N_23267,N_19476,N_20464);
nand U23268 (N_23268,N_20570,N_19838);
nor U23269 (N_23269,N_18981,N_20410);
or U23270 (N_23270,N_19587,N_19661);
nor U23271 (N_23271,N_20807,N_18963);
nand U23272 (N_23272,N_19406,N_19177);
nor U23273 (N_23273,N_21696,N_21438);
nand U23274 (N_23274,N_21655,N_21303);
or U23275 (N_23275,N_20380,N_21708);
nor U23276 (N_23276,N_19462,N_21673);
or U23277 (N_23277,N_19584,N_19647);
or U23278 (N_23278,N_21559,N_19033);
nand U23279 (N_23279,N_20058,N_19542);
xor U23280 (N_23280,N_19828,N_18886);
or U23281 (N_23281,N_20115,N_20855);
xnor U23282 (N_23282,N_21393,N_19625);
and U23283 (N_23283,N_20418,N_20263);
xor U23284 (N_23284,N_20948,N_21235);
nand U23285 (N_23285,N_21653,N_21543);
and U23286 (N_23286,N_21107,N_20343);
nand U23287 (N_23287,N_19640,N_20171);
nand U23288 (N_23288,N_21237,N_20923);
or U23289 (N_23289,N_20853,N_18881);
xnor U23290 (N_23290,N_20512,N_18945);
and U23291 (N_23291,N_19148,N_20494);
and U23292 (N_23292,N_19404,N_19383);
nor U23293 (N_23293,N_19372,N_19446);
xnor U23294 (N_23294,N_20676,N_20742);
xnor U23295 (N_23295,N_19759,N_19530);
xnor U23296 (N_23296,N_20927,N_21812);
and U23297 (N_23297,N_19651,N_19946);
xor U23298 (N_23298,N_20971,N_20922);
nand U23299 (N_23299,N_20004,N_19610);
nand U23300 (N_23300,N_21334,N_20898);
nand U23301 (N_23301,N_20260,N_21217);
xnor U23302 (N_23302,N_19672,N_21403);
or U23303 (N_23303,N_19769,N_19849);
or U23304 (N_23304,N_19624,N_19481);
or U23305 (N_23305,N_20168,N_21215);
nand U23306 (N_23306,N_20228,N_21668);
xor U23307 (N_23307,N_21629,N_19518);
and U23308 (N_23308,N_21152,N_20413);
nand U23309 (N_23309,N_19227,N_20375);
and U23310 (N_23310,N_21793,N_20654);
nor U23311 (N_23311,N_21600,N_20843);
and U23312 (N_23312,N_20825,N_20718);
and U23313 (N_23313,N_19995,N_21188);
and U23314 (N_23314,N_21746,N_19644);
and U23315 (N_23315,N_21489,N_19101);
xor U23316 (N_23316,N_20722,N_20471);
or U23317 (N_23317,N_20386,N_21809);
xnor U23318 (N_23318,N_21421,N_18938);
nor U23319 (N_23319,N_21753,N_19370);
nand U23320 (N_23320,N_20556,N_20532);
nor U23321 (N_23321,N_21637,N_19491);
or U23322 (N_23322,N_19835,N_20216);
and U23323 (N_23323,N_20724,N_20301);
and U23324 (N_23324,N_20117,N_21534);
or U23325 (N_23325,N_20702,N_20278);
xnor U23326 (N_23326,N_18987,N_20893);
or U23327 (N_23327,N_19737,N_19167);
or U23328 (N_23328,N_21568,N_19973);
or U23329 (N_23329,N_20373,N_20831);
nand U23330 (N_23330,N_20306,N_20983);
nand U23331 (N_23331,N_21439,N_19903);
or U23332 (N_23332,N_20830,N_19128);
nand U23333 (N_23333,N_20672,N_19699);
xor U23334 (N_23334,N_21818,N_20731);
xor U23335 (N_23335,N_20626,N_19171);
nor U23336 (N_23336,N_19841,N_19803);
nor U23337 (N_23337,N_21275,N_20185);
nand U23338 (N_23338,N_20276,N_21510);
nand U23339 (N_23339,N_18912,N_20330);
nand U23340 (N_23340,N_21105,N_20867);
and U23341 (N_23341,N_21599,N_21169);
and U23342 (N_23342,N_21277,N_19380);
and U23343 (N_23343,N_20543,N_19132);
nor U23344 (N_23344,N_21010,N_19747);
nand U23345 (N_23345,N_20999,N_19793);
or U23346 (N_23346,N_19500,N_18772);
xor U23347 (N_23347,N_21856,N_19522);
xnor U23348 (N_23348,N_20685,N_20573);
xor U23349 (N_23349,N_21301,N_20805);
nand U23350 (N_23350,N_21387,N_19232);
xor U23351 (N_23351,N_20108,N_20177);
nand U23352 (N_23352,N_18892,N_21211);
or U23353 (N_23353,N_21171,N_19467);
nor U23354 (N_23354,N_19541,N_21369);
or U23355 (N_23355,N_19198,N_19657);
nor U23356 (N_23356,N_21806,N_21208);
nand U23357 (N_23357,N_19055,N_20034);
nor U23358 (N_23358,N_19687,N_19174);
or U23359 (N_23359,N_20738,N_20961);
nand U23360 (N_23360,N_20010,N_21065);
xor U23361 (N_23361,N_20661,N_20022);
xnor U23362 (N_23362,N_20903,N_21351);
nor U23363 (N_23363,N_21106,N_21586);
nor U23364 (N_23364,N_21499,N_19729);
or U23365 (N_23365,N_20402,N_20538);
nor U23366 (N_23366,N_19562,N_21086);
nand U23367 (N_23367,N_20502,N_18923);
nor U23368 (N_23368,N_20696,N_19397);
nand U23369 (N_23369,N_20110,N_21699);
or U23370 (N_23370,N_21376,N_19504);
and U23371 (N_23371,N_19843,N_19520);
and U23372 (N_23372,N_21396,N_18810);
xnor U23373 (N_23373,N_20336,N_20451);
and U23374 (N_23374,N_20007,N_21112);
xor U23375 (N_23375,N_18818,N_21295);
or U23376 (N_23376,N_21524,N_20966);
xor U23377 (N_23377,N_19215,N_18756);
xor U23378 (N_23378,N_21825,N_19643);
and U23379 (N_23379,N_18789,N_19628);
xnor U23380 (N_23380,N_21343,N_19799);
or U23381 (N_23381,N_21021,N_20912);
nor U23382 (N_23382,N_18811,N_19533);
and U23383 (N_23383,N_18991,N_18936);
or U23384 (N_23384,N_19859,N_19023);
or U23385 (N_23385,N_20011,N_19081);
and U23386 (N_23386,N_20832,N_21736);
nor U23387 (N_23387,N_20191,N_19621);
nor U23388 (N_23388,N_20608,N_21416);
nor U23389 (N_23389,N_20352,N_20897);
xor U23390 (N_23390,N_19974,N_21011);
and U23391 (N_23391,N_21090,N_19084);
nor U23392 (N_23392,N_18966,N_18761);
and U23393 (N_23393,N_20020,N_21697);
xor U23394 (N_23394,N_21814,N_20518);
nor U23395 (N_23395,N_21757,N_19051);
nor U23396 (N_23396,N_20546,N_19386);
or U23397 (N_23397,N_20487,N_21663);
xnor U23398 (N_23398,N_19911,N_20249);
or U23399 (N_23399,N_19418,N_20209);
nor U23400 (N_23400,N_20105,N_21120);
xor U23401 (N_23401,N_21420,N_18784);
nand U23402 (N_23402,N_21597,N_19456);
and U23403 (N_23403,N_20631,N_21092);
xnor U23404 (N_23404,N_21726,N_20618);
and U23405 (N_23405,N_20791,N_18933);
xor U23406 (N_23406,N_21509,N_19290);
xor U23407 (N_23407,N_20172,N_21363);
nand U23408 (N_23408,N_19994,N_21216);
nand U23409 (N_23409,N_21113,N_19069);
and U23410 (N_23410,N_21366,N_21379);
nor U23411 (N_23411,N_21544,N_20470);
nand U23412 (N_23412,N_20327,N_21616);
nor U23413 (N_23413,N_19832,N_19929);
and U23414 (N_23414,N_19623,N_19142);
nor U23415 (N_23415,N_19821,N_20650);
or U23416 (N_23416,N_19582,N_21123);
or U23417 (N_23417,N_20097,N_19118);
or U23418 (N_23418,N_20351,N_21042);
nor U23419 (N_23419,N_21661,N_20771);
and U23420 (N_23420,N_19940,N_18995);
and U23421 (N_23421,N_20530,N_19756);
and U23422 (N_23422,N_19771,N_19375);
nand U23423 (N_23423,N_20569,N_21241);
and U23424 (N_23424,N_19678,N_20876);
and U23425 (N_23425,N_19701,N_21194);
and U23426 (N_23426,N_20176,N_21639);
and U23427 (N_23427,N_20214,N_19115);
and U23428 (N_23428,N_19780,N_18822);
nand U23429 (N_23429,N_20621,N_20486);
xor U23430 (N_23430,N_18758,N_21057);
or U23431 (N_23431,N_18946,N_19334);
and U23432 (N_23432,N_19516,N_21412);
nor U23433 (N_23433,N_20677,N_19906);
or U23434 (N_23434,N_21446,N_19553);
nor U23435 (N_23435,N_21430,N_18870);
nand U23436 (N_23436,N_21727,N_19673);
or U23437 (N_23437,N_19717,N_20719);
nand U23438 (N_23438,N_21442,N_20197);
xor U23439 (N_23439,N_20239,N_19906);
and U23440 (N_23440,N_19925,N_19539);
or U23441 (N_23441,N_21474,N_19366);
and U23442 (N_23442,N_19264,N_20420);
and U23443 (N_23443,N_19123,N_19319);
or U23444 (N_23444,N_19660,N_18766);
nand U23445 (N_23445,N_21554,N_20728);
nand U23446 (N_23446,N_21689,N_19931);
and U23447 (N_23447,N_21223,N_19781);
xnor U23448 (N_23448,N_20338,N_21518);
xnor U23449 (N_23449,N_19592,N_20433);
xor U23450 (N_23450,N_19215,N_19080);
nor U23451 (N_23451,N_21764,N_21103);
and U23452 (N_23452,N_21208,N_20911);
xor U23453 (N_23453,N_21527,N_21041);
or U23454 (N_23454,N_21526,N_19938);
nand U23455 (N_23455,N_21729,N_20763);
nor U23456 (N_23456,N_19181,N_19653);
xor U23457 (N_23457,N_20499,N_20255);
or U23458 (N_23458,N_19924,N_19646);
and U23459 (N_23459,N_21513,N_19983);
and U23460 (N_23460,N_20316,N_20394);
nor U23461 (N_23461,N_20640,N_20006);
nand U23462 (N_23462,N_18790,N_20260);
xor U23463 (N_23463,N_21139,N_19257);
nand U23464 (N_23464,N_18752,N_19627);
and U23465 (N_23465,N_19298,N_19780);
nand U23466 (N_23466,N_21671,N_20769);
nor U23467 (N_23467,N_21163,N_20713);
or U23468 (N_23468,N_19982,N_19181);
or U23469 (N_23469,N_19715,N_21333);
xor U23470 (N_23470,N_21283,N_20328);
xor U23471 (N_23471,N_21047,N_20496);
xor U23472 (N_23472,N_21512,N_19338);
xor U23473 (N_23473,N_18929,N_19791);
and U23474 (N_23474,N_20498,N_19793);
and U23475 (N_23475,N_18796,N_19062);
nand U23476 (N_23476,N_19206,N_19846);
and U23477 (N_23477,N_21322,N_20395);
nand U23478 (N_23478,N_21311,N_20454);
nor U23479 (N_23479,N_19117,N_19475);
nor U23480 (N_23480,N_20362,N_21194);
xor U23481 (N_23481,N_20691,N_21343);
nand U23482 (N_23482,N_19886,N_20512);
and U23483 (N_23483,N_19628,N_19590);
and U23484 (N_23484,N_19441,N_19098);
nor U23485 (N_23485,N_20885,N_19247);
xnor U23486 (N_23486,N_21033,N_20420);
nand U23487 (N_23487,N_20420,N_21017);
and U23488 (N_23488,N_20933,N_20692);
or U23489 (N_23489,N_21754,N_21116);
nand U23490 (N_23490,N_19738,N_20470);
or U23491 (N_23491,N_20958,N_18858);
and U23492 (N_23492,N_20345,N_19537);
nor U23493 (N_23493,N_19137,N_20116);
or U23494 (N_23494,N_21020,N_21084);
nand U23495 (N_23495,N_21037,N_20340);
xnor U23496 (N_23496,N_21736,N_20526);
nor U23497 (N_23497,N_21204,N_20485);
and U23498 (N_23498,N_20914,N_21201);
nor U23499 (N_23499,N_18772,N_21128);
or U23500 (N_23500,N_19879,N_19661);
nand U23501 (N_23501,N_20578,N_19381);
nor U23502 (N_23502,N_20137,N_19638);
or U23503 (N_23503,N_20104,N_21264);
and U23504 (N_23504,N_21206,N_19567);
nor U23505 (N_23505,N_19440,N_21531);
nand U23506 (N_23506,N_20841,N_20074);
nand U23507 (N_23507,N_19906,N_19596);
nor U23508 (N_23508,N_19451,N_21775);
and U23509 (N_23509,N_20213,N_20466);
nand U23510 (N_23510,N_19221,N_20519);
nand U23511 (N_23511,N_19576,N_18763);
nand U23512 (N_23512,N_21012,N_20145);
nor U23513 (N_23513,N_19697,N_20424);
and U23514 (N_23514,N_21554,N_21537);
or U23515 (N_23515,N_21202,N_21051);
xnor U23516 (N_23516,N_20586,N_19232);
xnor U23517 (N_23517,N_19947,N_20878);
nand U23518 (N_23518,N_21854,N_19903);
and U23519 (N_23519,N_19387,N_18907);
and U23520 (N_23520,N_19719,N_18946);
and U23521 (N_23521,N_19563,N_19749);
nor U23522 (N_23522,N_21106,N_19262);
xnor U23523 (N_23523,N_18942,N_19043);
and U23524 (N_23524,N_19859,N_20055);
nand U23525 (N_23525,N_21509,N_19746);
and U23526 (N_23526,N_20524,N_19995);
nor U23527 (N_23527,N_20688,N_19402);
or U23528 (N_23528,N_18920,N_20647);
xor U23529 (N_23529,N_20143,N_19364);
nor U23530 (N_23530,N_19351,N_20904);
and U23531 (N_23531,N_20894,N_18805);
or U23532 (N_23532,N_19753,N_20939);
nand U23533 (N_23533,N_19055,N_19291);
and U23534 (N_23534,N_19201,N_20924);
nand U23535 (N_23535,N_21470,N_19309);
and U23536 (N_23536,N_21556,N_19656);
or U23537 (N_23537,N_20190,N_19111);
nor U23538 (N_23538,N_20109,N_20315);
nor U23539 (N_23539,N_19061,N_19216);
xor U23540 (N_23540,N_20227,N_21454);
and U23541 (N_23541,N_20714,N_20909);
nor U23542 (N_23542,N_21382,N_20502);
or U23543 (N_23543,N_21758,N_20655);
nand U23544 (N_23544,N_19737,N_19038);
xor U23545 (N_23545,N_20026,N_21529);
or U23546 (N_23546,N_19123,N_19820);
nor U23547 (N_23547,N_20974,N_20289);
nand U23548 (N_23548,N_18914,N_19042);
xor U23549 (N_23549,N_21113,N_19285);
and U23550 (N_23550,N_20834,N_20193);
nand U23551 (N_23551,N_21154,N_21134);
nor U23552 (N_23552,N_18977,N_21310);
xor U23553 (N_23553,N_21585,N_21854);
and U23554 (N_23554,N_19120,N_20401);
nor U23555 (N_23555,N_19196,N_19264);
nand U23556 (N_23556,N_21305,N_20576);
xnor U23557 (N_23557,N_21085,N_21740);
or U23558 (N_23558,N_19352,N_19864);
and U23559 (N_23559,N_20417,N_19646);
nor U23560 (N_23560,N_21738,N_19790);
xor U23561 (N_23561,N_19228,N_20362);
nand U23562 (N_23562,N_20991,N_21449);
and U23563 (N_23563,N_20782,N_21497);
and U23564 (N_23564,N_19989,N_18863);
xnor U23565 (N_23565,N_19492,N_18850);
or U23566 (N_23566,N_18940,N_19409);
nand U23567 (N_23567,N_19741,N_19948);
and U23568 (N_23568,N_19909,N_20402);
nand U23569 (N_23569,N_20392,N_19810);
or U23570 (N_23570,N_20504,N_19311);
or U23571 (N_23571,N_19304,N_19170);
nand U23572 (N_23572,N_20827,N_20366);
xnor U23573 (N_23573,N_21763,N_21515);
nor U23574 (N_23574,N_21540,N_21643);
nor U23575 (N_23575,N_20149,N_20649);
xnor U23576 (N_23576,N_21681,N_21750);
nor U23577 (N_23577,N_20015,N_21747);
or U23578 (N_23578,N_18798,N_19145);
nand U23579 (N_23579,N_21815,N_20281);
nand U23580 (N_23580,N_20963,N_21237);
and U23581 (N_23581,N_21605,N_19300);
xor U23582 (N_23582,N_19910,N_21130);
and U23583 (N_23583,N_20749,N_21758);
and U23584 (N_23584,N_21520,N_18956);
or U23585 (N_23585,N_20590,N_21160);
and U23586 (N_23586,N_21489,N_21628);
or U23587 (N_23587,N_21831,N_21539);
and U23588 (N_23588,N_21100,N_19466);
and U23589 (N_23589,N_21285,N_19926);
nand U23590 (N_23590,N_19606,N_20505);
nand U23591 (N_23591,N_19056,N_19321);
xnor U23592 (N_23592,N_18863,N_20193);
nand U23593 (N_23593,N_18787,N_21634);
nor U23594 (N_23594,N_21489,N_19515);
nand U23595 (N_23595,N_21141,N_19402);
nor U23596 (N_23596,N_20509,N_21246);
and U23597 (N_23597,N_20139,N_20967);
xnor U23598 (N_23598,N_19677,N_21141);
nand U23599 (N_23599,N_21396,N_21690);
xor U23600 (N_23600,N_19724,N_21081);
and U23601 (N_23601,N_21315,N_20890);
nor U23602 (N_23602,N_19605,N_19356);
xor U23603 (N_23603,N_20474,N_19587);
nand U23604 (N_23604,N_19197,N_19258);
xor U23605 (N_23605,N_21555,N_19798);
or U23606 (N_23606,N_18993,N_19148);
and U23607 (N_23607,N_19456,N_19198);
xnor U23608 (N_23608,N_19624,N_21161);
xnor U23609 (N_23609,N_18795,N_20675);
xnor U23610 (N_23610,N_21136,N_21710);
xor U23611 (N_23611,N_19111,N_18750);
nand U23612 (N_23612,N_19624,N_20892);
or U23613 (N_23613,N_21706,N_20801);
nor U23614 (N_23614,N_19735,N_18890);
or U23615 (N_23615,N_19427,N_20198);
or U23616 (N_23616,N_19059,N_18787);
xor U23617 (N_23617,N_20185,N_21261);
and U23618 (N_23618,N_21376,N_21811);
nand U23619 (N_23619,N_21398,N_18993);
nor U23620 (N_23620,N_21202,N_19871);
and U23621 (N_23621,N_19497,N_20682);
xnor U23622 (N_23622,N_20630,N_20423);
or U23623 (N_23623,N_19534,N_19263);
and U23624 (N_23624,N_21351,N_19184);
xnor U23625 (N_23625,N_21286,N_20941);
nor U23626 (N_23626,N_21368,N_19615);
nor U23627 (N_23627,N_21190,N_19677);
xnor U23628 (N_23628,N_21828,N_20244);
or U23629 (N_23629,N_19970,N_20695);
nand U23630 (N_23630,N_21231,N_21211);
or U23631 (N_23631,N_21482,N_19722);
nor U23632 (N_23632,N_19708,N_20290);
nand U23633 (N_23633,N_19323,N_21425);
or U23634 (N_23634,N_19685,N_21277);
nand U23635 (N_23635,N_19318,N_19261);
nand U23636 (N_23636,N_20258,N_20687);
xor U23637 (N_23637,N_19493,N_20244);
nor U23638 (N_23638,N_20779,N_19009);
nand U23639 (N_23639,N_18851,N_20036);
nor U23640 (N_23640,N_19028,N_20277);
and U23641 (N_23641,N_20321,N_18798);
nor U23642 (N_23642,N_20241,N_19410);
nor U23643 (N_23643,N_21180,N_19405);
nor U23644 (N_23644,N_20938,N_19274);
xnor U23645 (N_23645,N_21064,N_19852);
nand U23646 (N_23646,N_19605,N_19215);
xnor U23647 (N_23647,N_21431,N_21535);
nand U23648 (N_23648,N_21749,N_19807);
or U23649 (N_23649,N_19466,N_18902);
xnor U23650 (N_23650,N_18906,N_20363);
nor U23651 (N_23651,N_18975,N_21137);
nand U23652 (N_23652,N_20969,N_19380);
or U23653 (N_23653,N_20978,N_18853);
nand U23654 (N_23654,N_19381,N_21693);
nand U23655 (N_23655,N_21647,N_19071);
xnor U23656 (N_23656,N_20616,N_20005);
or U23657 (N_23657,N_21641,N_21553);
nor U23658 (N_23658,N_20318,N_18851);
nand U23659 (N_23659,N_20226,N_18904);
nand U23660 (N_23660,N_19393,N_19238);
xor U23661 (N_23661,N_21427,N_21158);
nand U23662 (N_23662,N_21758,N_19233);
nor U23663 (N_23663,N_21359,N_20132);
xnor U23664 (N_23664,N_21186,N_19852);
nor U23665 (N_23665,N_20120,N_19868);
xor U23666 (N_23666,N_21280,N_21835);
nor U23667 (N_23667,N_20118,N_20166);
nand U23668 (N_23668,N_21122,N_19045);
nand U23669 (N_23669,N_19503,N_19890);
xnor U23670 (N_23670,N_19770,N_19216);
xor U23671 (N_23671,N_21356,N_20557);
and U23672 (N_23672,N_21639,N_18790);
xnor U23673 (N_23673,N_20857,N_20338);
nand U23674 (N_23674,N_20290,N_18942);
nand U23675 (N_23675,N_19956,N_21304);
xnor U23676 (N_23676,N_18901,N_19444);
xor U23677 (N_23677,N_19383,N_19059);
or U23678 (N_23678,N_20663,N_20506);
xnor U23679 (N_23679,N_21765,N_19896);
and U23680 (N_23680,N_19669,N_19022);
or U23681 (N_23681,N_18780,N_19697);
nand U23682 (N_23682,N_20989,N_19703);
and U23683 (N_23683,N_19954,N_19738);
nor U23684 (N_23684,N_21589,N_19865);
nor U23685 (N_23685,N_21459,N_19981);
and U23686 (N_23686,N_20711,N_21234);
and U23687 (N_23687,N_18859,N_18756);
and U23688 (N_23688,N_20051,N_21028);
or U23689 (N_23689,N_21024,N_20167);
or U23690 (N_23690,N_21078,N_19347);
nand U23691 (N_23691,N_21846,N_20284);
xor U23692 (N_23692,N_21657,N_21764);
and U23693 (N_23693,N_20208,N_21701);
nand U23694 (N_23694,N_20416,N_21181);
and U23695 (N_23695,N_21240,N_18920);
nand U23696 (N_23696,N_21418,N_21073);
xnor U23697 (N_23697,N_21668,N_20049);
or U23698 (N_23698,N_21195,N_21263);
nor U23699 (N_23699,N_21683,N_19357);
nand U23700 (N_23700,N_19172,N_19823);
nand U23701 (N_23701,N_19222,N_19060);
nand U23702 (N_23702,N_19924,N_20993);
xnor U23703 (N_23703,N_19854,N_20241);
nor U23704 (N_23704,N_21603,N_21581);
xnor U23705 (N_23705,N_19948,N_20064);
xor U23706 (N_23706,N_19584,N_19879);
nor U23707 (N_23707,N_20634,N_20443);
nand U23708 (N_23708,N_20785,N_18912);
and U23709 (N_23709,N_18802,N_21112);
nor U23710 (N_23710,N_21052,N_20009);
nand U23711 (N_23711,N_20091,N_21115);
or U23712 (N_23712,N_19671,N_20375);
nor U23713 (N_23713,N_21172,N_19292);
or U23714 (N_23714,N_21160,N_20863);
xor U23715 (N_23715,N_20248,N_19671);
xor U23716 (N_23716,N_19918,N_19420);
nand U23717 (N_23717,N_20948,N_19189);
nor U23718 (N_23718,N_18932,N_21743);
or U23719 (N_23719,N_18969,N_21464);
nor U23720 (N_23720,N_20035,N_20739);
and U23721 (N_23721,N_21265,N_19882);
and U23722 (N_23722,N_21182,N_19574);
xor U23723 (N_23723,N_20630,N_19585);
xnor U23724 (N_23724,N_20721,N_19013);
or U23725 (N_23725,N_20259,N_19612);
or U23726 (N_23726,N_19807,N_20221);
or U23727 (N_23727,N_20751,N_20596);
and U23728 (N_23728,N_20307,N_18876);
xor U23729 (N_23729,N_21666,N_21384);
nand U23730 (N_23730,N_20350,N_19725);
or U23731 (N_23731,N_21454,N_19955);
xor U23732 (N_23732,N_19300,N_20110);
nor U23733 (N_23733,N_21444,N_21731);
or U23734 (N_23734,N_19785,N_19078);
and U23735 (N_23735,N_20419,N_20244);
nor U23736 (N_23736,N_21782,N_19284);
or U23737 (N_23737,N_20672,N_21500);
nor U23738 (N_23738,N_21194,N_20293);
or U23739 (N_23739,N_21413,N_21280);
nand U23740 (N_23740,N_20354,N_20241);
and U23741 (N_23741,N_21370,N_20370);
or U23742 (N_23742,N_20208,N_21167);
nand U23743 (N_23743,N_19395,N_21818);
or U23744 (N_23744,N_20483,N_19283);
or U23745 (N_23745,N_19143,N_21221);
and U23746 (N_23746,N_20207,N_21607);
or U23747 (N_23747,N_20620,N_21197);
nand U23748 (N_23748,N_19696,N_20635);
nand U23749 (N_23749,N_21299,N_21414);
and U23750 (N_23750,N_21521,N_19222);
or U23751 (N_23751,N_20361,N_19528);
or U23752 (N_23752,N_21172,N_18805);
nor U23753 (N_23753,N_18769,N_18968);
nand U23754 (N_23754,N_18805,N_18882);
or U23755 (N_23755,N_20620,N_19394);
nand U23756 (N_23756,N_18790,N_19432);
or U23757 (N_23757,N_21111,N_19101);
and U23758 (N_23758,N_19470,N_21155);
nand U23759 (N_23759,N_19566,N_19569);
or U23760 (N_23760,N_21185,N_19033);
xor U23761 (N_23761,N_20208,N_20661);
xor U23762 (N_23762,N_21753,N_20885);
nor U23763 (N_23763,N_20480,N_18792);
nand U23764 (N_23764,N_19785,N_20068);
or U23765 (N_23765,N_18877,N_21031);
and U23766 (N_23766,N_20820,N_21605);
or U23767 (N_23767,N_20331,N_19592);
nand U23768 (N_23768,N_19846,N_19707);
or U23769 (N_23769,N_21863,N_19003);
or U23770 (N_23770,N_21655,N_21059);
nor U23771 (N_23771,N_19691,N_20357);
xor U23772 (N_23772,N_21792,N_21300);
nor U23773 (N_23773,N_19574,N_19218);
nand U23774 (N_23774,N_19847,N_19231);
or U23775 (N_23775,N_20605,N_21777);
xor U23776 (N_23776,N_20793,N_19257);
nor U23777 (N_23777,N_20544,N_19403);
or U23778 (N_23778,N_20808,N_19916);
nand U23779 (N_23779,N_20798,N_20310);
nor U23780 (N_23780,N_20157,N_20196);
nand U23781 (N_23781,N_20015,N_19187);
and U23782 (N_23782,N_21729,N_18820);
xor U23783 (N_23783,N_19324,N_19135);
nand U23784 (N_23784,N_20439,N_19389);
nor U23785 (N_23785,N_20561,N_20537);
and U23786 (N_23786,N_19385,N_18876);
nor U23787 (N_23787,N_19102,N_21833);
or U23788 (N_23788,N_20961,N_21841);
xnor U23789 (N_23789,N_21518,N_20153);
and U23790 (N_23790,N_20846,N_21341);
or U23791 (N_23791,N_21708,N_19395);
nand U23792 (N_23792,N_21562,N_19316);
or U23793 (N_23793,N_20440,N_20678);
or U23794 (N_23794,N_19170,N_19956);
nand U23795 (N_23795,N_20649,N_21126);
xnor U23796 (N_23796,N_19316,N_20889);
and U23797 (N_23797,N_18851,N_20888);
nor U23798 (N_23798,N_20810,N_19029);
nand U23799 (N_23799,N_20846,N_21694);
xnor U23800 (N_23800,N_21373,N_21153);
xor U23801 (N_23801,N_20147,N_20403);
and U23802 (N_23802,N_21414,N_21560);
and U23803 (N_23803,N_21215,N_19937);
and U23804 (N_23804,N_20693,N_19955);
xor U23805 (N_23805,N_19629,N_20672);
nand U23806 (N_23806,N_19961,N_21193);
nor U23807 (N_23807,N_19708,N_20154);
or U23808 (N_23808,N_19554,N_20577);
nand U23809 (N_23809,N_21180,N_20362);
nand U23810 (N_23810,N_19481,N_20087);
and U23811 (N_23811,N_21664,N_18750);
nor U23812 (N_23812,N_21387,N_20602);
xnor U23813 (N_23813,N_20655,N_20799);
nor U23814 (N_23814,N_20116,N_19263);
and U23815 (N_23815,N_20482,N_20056);
or U23816 (N_23816,N_20012,N_20815);
nor U23817 (N_23817,N_21402,N_20135);
xnor U23818 (N_23818,N_19061,N_21474);
nand U23819 (N_23819,N_19956,N_21477);
xor U23820 (N_23820,N_20337,N_21174);
xor U23821 (N_23821,N_20545,N_21438);
nor U23822 (N_23822,N_21149,N_20072);
nand U23823 (N_23823,N_20810,N_21868);
xor U23824 (N_23824,N_20856,N_19152);
or U23825 (N_23825,N_20926,N_19750);
nand U23826 (N_23826,N_19320,N_18901);
xor U23827 (N_23827,N_19756,N_21790);
nand U23828 (N_23828,N_19899,N_19986);
nor U23829 (N_23829,N_19309,N_19723);
nor U23830 (N_23830,N_19311,N_19768);
or U23831 (N_23831,N_19685,N_19776);
and U23832 (N_23832,N_19819,N_18937);
nand U23833 (N_23833,N_21482,N_20583);
xnor U23834 (N_23834,N_19521,N_21601);
xor U23835 (N_23835,N_20782,N_20327);
xnor U23836 (N_23836,N_20959,N_21561);
nand U23837 (N_23837,N_18852,N_18863);
and U23838 (N_23838,N_19798,N_21663);
nor U23839 (N_23839,N_21849,N_20087);
nand U23840 (N_23840,N_18778,N_20078);
nor U23841 (N_23841,N_21153,N_21056);
nor U23842 (N_23842,N_21530,N_19851);
nand U23843 (N_23843,N_20207,N_19975);
nor U23844 (N_23844,N_20652,N_21541);
or U23845 (N_23845,N_18971,N_19971);
nor U23846 (N_23846,N_21160,N_20618);
nand U23847 (N_23847,N_19865,N_19153);
nand U23848 (N_23848,N_20803,N_20678);
xor U23849 (N_23849,N_20953,N_20725);
nand U23850 (N_23850,N_19164,N_20846);
or U23851 (N_23851,N_18947,N_20987);
xor U23852 (N_23852,N_21401,N_18786);
or U23853 (N_23853,N_20053,N_19451);
or U23854 (N_23854,N_19641,N_20596);
or U23855 (N_23855,N_18845,N_20435);
nand U23856 (N_23856,N_19323,N_20029);
nand U23857 (N_23857,N_20945,N_21694);
xor U23858 (N_23858,N_20838,N_19447);
nor U23859 (N_23859,N_19195,N_19244);
nor U23860 (N_23860,N_19484,N_20166);
nor U23861 (N_23861,N_19657,N_21494);
nor U23862 (N_23862,N_19592,N_21398);
nor U23863 (N_23863,N_19410,N_19369);
or U23864 (N_23864,N_20548,N_19538);
nand U23865 (N_23865,N_19627,N_21183);
or U23866 (N_23866,N_20418,N_21698);
nand U23867 (N_23867,N_19069,N_18954);
and U23868 (N_23868,N_19775,N_21511);
xnor U23869 (N_23869,N_19062,N_20240);
or U23870 (N_23870,N_20664,N_20685);
nand U23871 (N_23871,N_21029,N_21799);
nor U23872 (N_23872,N_20223,N_20986);
xor U23873 (N_23873,N_19810,N_20409);
or U23874 (N_23874,N_21714,N_19348);
nand U23875 (N_23875,N_21680,N_21137);
nor U23876 (N_23876,N_21564,N_20256);
and U23877 (N_23877,N_19420,N_21344);
nand U23878 (N_23878,N_19763,N_18767);
and U23879 (N_23879,N_20119,N_20103);
or U23880 (N_23880,N_19078,N_19782);
or U23881 (N_23881,N_19710,N_21700);
xor U23882 (N_23882,N_21849,N_21519);
and U23883 (N_23883,N_19435,N_21546);
nand U23884 (N_23884,N_20511,N_20840);
and U23885 (N_23885,N_20005,N_19654);
and U23886 (N_23886,N_19064,N_19055);
xnor U23887 (N_23887,N_20003,N_21650);
and U23888 (N_23888,N_20948,N_21489);
nor U23889 (N_23889,N_19421,N_19827);
nand U23890 (N_23890,N_21735,N_21575);
or U23891 (N_23891,N_19787,N_20415);
and U23892 (N_23892,N_19726,N_19792);
and U23893 (N_23893,N_20162,N_21187);
and U23894 (N_23894,N_18808,N_21676);
or U23895 (N_23895,N_20130,N_19034);
nand U23896 (N_23896,N_20621,N_20693);
xnor U23897 (N_23897,N_20404,N_19136);
or U23898 (N_23898,N_20345,N_19304);
and U23899 (N_23899,N_20282,N_19542);
or U23900 (N_23900,N_21728,N_18935);
nand U23901 (N_23901,N_20710,N_19998);
nand U23902 (N_23902,N_18861,N_19523);
nor U23903 (N_23903,N_20536,N_21863);
xnor U23904 (N_23904,N_21162,N_19357);
or U23905 (N_23905,N_19943,N_19315);
and U23906 (N_23906,N_21707,N_21359);
and U23907 (N_23907,N_19704,N_19587);
and U23908 (N_23908,N_20054,N_20353);
nand U23909 (N_23909,N_21038,N_21701);
or U23910 (N_23910,N_20093,N_20334);
and U23911 (N_23911,N_19664,N_19457);
or U23912 (N_23912,N_19128,N_21799);
nor U23913 (N_23913,N_19601,N_20416);
and U23914 (N_23914,N_20473,N_21063);
and U23915 (N_23915,N_19535,N_21538);
nand U23916 (N_23916,N_19121,N_19759);
nor U23917 (N_23917,N_20764,N_21448);
nor U23918 (N_23918,N_20623,N_20087);
or U23919 (N_23919,N_18816,N_19305);
nand U23920 (N_23920,N_20661,N_19307);
and U23921 (N_23921,N_21356,N_21095);
nand U23922 (N_23922,N_20684,N_18982);
or U23923 (N_23923,N_18940,N_20611);
and U23924 (N_23924,N_19973,N_20149);
nor U23925 (N_23925,N_19654,N_19460);
nand U23926 (N_23926,N_21567,N_19253);
and U23927 (N_23927,N_20703,N_21482);
xor U23928 (N_23928,N_19766,N_21577);
or U23929 (N_23929,N_21190,N_19390);
nand U23930 (N_23930,N_21686,N_20724);
xor U23931 (N_23931,N_19312,N_21530);
nand U23932 (N_23932,N_18942,N_20752);
and U23933 (N_23933,N_21641,N_21146);
or U23934 (N_23934,N_21859,N_21380);
and U23935 (N_23935,N_20360,N_20536);
and U23936 (N_23936,N_20964,N_21458);
xor U23937 (N_23937,N_20074,N_19865);
or U23938 (N_23938,N_20503,N_21775);
xnor U23939 (N_23939,N_20482,N_18981);
xnor U23940 (N_23940,N_20912,N_20903);
nor U23941 (N_23941,N_19343,N_20877);
nand U23942 (N_23942,N_20347,N_19338);
and U23943 (N_23943,N_19140,N_21586);
nand U23944 (N_23944,N_20877,N_21068);
xnor U23945 (N_23945,N_19503,N_20638);
or U23946 (N_23946,N_20736,N_20720);
nand U23947 (N_23947,N_20481,N_21842);
nor U23948 (N_23948,N_20987,N_20953);
nand U23949 (N_23949,N_20761,N_19085);
or U23950 (N_23950,N_20924,N_20933);
nand U23951 (N_23951,N_20787,N_19856);
nand U23952 (N_23952,N_21036,N_20091);
and U23953 (N_23953,N_20309,N_18839);
and U23954 (N_23954,N_21628,N_19489);
and U23955 (N_23955,N_21779,N_21752);
nor U23956 (N_23956,N_20984,N_19376);
xnor U23957 (N_23957,N_21739,N_18765);
xnor U23958 (N_23958,N_19510,N_19595);
and U23959 (N_23959,N_21801,N_19237);
nor U23960 (N_23960,N_20870,N_19455);
and U23961 (N_23961,N_19545,N_19540);
nor U23962 (N_23962,N_20757,N_20911);
or U23963 (N_23963,N_19144,N_21767);
and U23964 (N_23964,N_20800,N_19891);
nor U23965 (N_23965,N_21332,N_21129);
xnor U23966 (N_23966,N_20332,N_20331);
and U23967 (N_23967,N_21463,N_21803);
or U23968 (N_23968,N_21449,N_21011);
and U23969 (N_23969,N_20998,N_20799);
nor U23970 (N_23970,N_21741,N_18803);
nand U23971 (N_23971,N_21009,N_21526);
or U23972 (N_23972,N_19147,N_21635);
nor U23973 (N_23973,N_18945,N_21851);
or U23974 (N_23974,N_20662,N_20634);
and U23975 (N_23975,N_19424,N_21032);
nand U23976 (N_23976,N_20440,N_19184);
nand U23977 (N_23977,N_21023,N_19112);
nor U23978 (N_23978,N_21181,N_19856);
xnor U23979 (N_23979,N_21502,N_18899);
xor U23980 (N_23980,N_18950,N_20180);
xnor U23981 (N_23981,N_21657,N_21517);
or U23982 (N_23982,N_19648,N_19215);
and U23983 (N_23983,N_19875,N_19490);
nor U23984 (N_23984,N_21471,N_21059);
nor U23985 (N_23985,N_21323,N_19658);
nor U23986 (N_23986,N_19314,N_19965);
nand U23987 (N_23987,N_20273,N_19359);
or U23988 (N_23988,N_20959,N_21768);
xnor U23989 (N_23989,N_19131,N_18994);
nand U23990 (N_23990,N_20665,N_20795);
nor U23991 (N_23991,N_19905,N_19377);
or U23992 (N_23992,N_20784,N_19813);
and U23993 (N_23993,N_21051,N_19817);
and U23994 (N_23994,N_20238,N_19983);
and U23995 (N_23995,N_19032,N_19221);
and U23996 (N_23996,N_19471,N_20516);
nand U23997 (N_23997,N_18810,N_21302);
and U23998 (N_23998,N_20202,N_19070);
or U23999 (N_23999,N_21632,N_20317);
nand U24000 (N_24000,N_20835,N_19884);
nor U24001 (N_24001,N_18769,N_20310);
nor U24002 (N_24002,N_21752,N_21488);
nor U24003 (N_24003,N_19837,N_21462);
xnor U24004 (N_24004,N_21871,N_20896);
xnor U24005 (N_24005,N_20514,N_19940);
xor U24006 (N_24006,N_19243,N_21394);
nand U24007 (N_24007,N_20415,N_21190);
nand U24008 (N_24008,N_20546,N_19749);
nor U24009 (N_24009,N_21395,N_19267);
or U24010 (N_24010,N_20521,N_20168);
nor U24011 (N_24011,N_19445,N_21867);
and U24012 (N_24012,N_21424,N_21527);
or U24013 (N_24013,N_20777,N_20600);
nand U24014 (N_24014,N_20589,N_20497);
nor U24015 (N_24015,N_19214,N_20108);
nand U24016 (N_24016,N_20047,N_19365);
and U24017 (N_24017,N_20923,N_20883);
xnor U24018 (N_24018,N_21645,N_21192);
nand U24019 (N_24019,N_20375,N_21263);
or U24020 (N_24020,N_21751,N_21383);
nor U24021 (N_24021,N_19358,N_18841);
xnor U24022 (N_24022,N_19097,N_20084);
nor U24023 (N_24023,N_21617,N_21525);
nor U24024 (N_24024,N_19630,N_20273);
or U24025 (N_24025,N_20003,N_19343);
nand U24026 (N_24026,N_21221,N_20438);
nand U24027 (N_24027,N_19725,N_19501);
nor U24028 (N_24028,N_21851,N_20469);
or U24029 (N_24029,N_18833,N_20381);
nor U24030 (N_24030,N_21039,N_20890);
nand U24031 (N_24031,N_19060,N_19298);
nor U24032 (N_24032,N_20210,N_21728);
nand U24033 (N_24033,N_18763,N_21044);
and U24034 (N_24034,N_21351,N_20991);
xnor U24035 (N_24035,N_21750,N_20395);
nand U24036 (N_24036,N_19921,N_21069);
nor U24037 (N_24037,N_21536,N_20650);
or U24038 (N_24038,N_21237,N_21120);
nand U24039 (N_24039,N_19727,N_19636);
or U24040 (N_24040,N_20618,N_18990);
and U24041 (N_24041,N_21798,N_19575);
or U24042 (N_24042,N_21783,N_21343);
nand U24043 (N_24043,N_21291,N_20974);
nand U24044 (N_24044,N_20929,N_19061);
nor U24045 (N_24045,N_19366,N_20545);
nand U24046 (N_24046,N_21446,N_20294);
nand U24047 (N_24047,N_19636,N_20674);
and U24048 (N_24048,N_19652,N_20702);
nand U24049 (N_24049,N_19157,N_20312);
nand U24050 (N_24050,N_19365,N_20840);
and U24051 (N_24051,N_19482,N_19264);
nand U24052 (N_24052,N_18782,N_21750);
nand U24053 (N_24053,N_20496,N_19802);
or U24054 (N_24054,N_19983,N_21358);
nor U24055 (N_24055,N_19745,N_19803);
nand U24056 (N_24056,N_21112,N_20551);
xnor U24057 (N_24057,N_21772,N_21830);
nor U24058 (N_24058,N_19384,N_19846);
and U24059 (N_24059,N_20163,N_19656);
nor U24060 (N_24060,N_19054,N_20126);
nand U24061 (N_24061,N_19622,N_20298);
nor U24062 (N_24062,N_20650,N_19977);
xor U24063 (N_24063,N_19978,N_21848);
xnor U24064 (N_24064,N_19516,N_21364);
nand U24065 (N_24065,N_20878,N_19203);
nand U24066 (N_24066,N_20806,N_21616);
nor U24067 (N_24067,N_19212,N_21216);
or U24068 (N_24068,N_19489,N_20133);
xnor U24069 (N_24069,N_21151,N_19160);
or U24070 (N_24070,N_18790,N_21062);
nor U24071 (N_24071,N_20229,N_21090);
and U24072 (N_24072,N_19986,N_19480);
nor U24073 (N_24073,N_21658,N_20783);
or U24074 (N_24074,N_21428,N_21026);
xnor U24075 (N_24075,N_20657,N_21392);
nand U24076 (N_24076,N_19377,N_20015);
or U24077 (N_24077,N_20434,N_20882);
and U24078 (N_24078,N_19032,N_19526);
or U24079 (N_24079,N_19958,N_19927);
nand U24080 (N_24080,N_19980,N_19127);
xnor U24081 (N_24081,N_18830,N_20437);
xnor U24082 (N_24082,N_20092,N_21735);
xnor U24083 (N_24083,N_20295,N_21322);
xor U24084 (N_24084,N_21545,N_21803);
and U24085 (N_24085,N_19388,N_20798);
or U24086 (N_24086,N_21030,N_18765);
nand U24087 (N_24087,N_20710,N_19839);
or U24088 (N_24088,N_20196,N_21153);
xor U24089 (N_24089,N_21503,N_20845);
xnor U24090 (N_24090,N_20699,N_19388);
xnor U24091 (N_24091,N_21345,N_20897);
and U24092 (N_24092,N_20295,N_19993);
nor U24093 (N_24093,N_21545,N_21826);
and U24094 (N_24094,N_19811,N_20065);
nand U24095 (N_24095,N_21324,N_20892);
nand U24096 (N_24096,N_20816,N_19804);
nand U24097 (N_24097,N_19062,N_18904);
or U24098 (N_24098,N_21522,N_20344);
nand U24099 (N_24099,N_19537,N_21230);
or U24100 (N_24100,N_20799,N_21732);
nand U24101 (N_24101,N_20964,N_21151);
xor U24102 (N_24102,N_19683,N_21398);
or U24103 (N_24103,N_21317,N_18865);
xor U24104 (N_24104,N_19164,N_19896);
or U24105 (N_24105,N_20305,N_20802);
and U24106 (N_24106,N_20306,N_19490);
nor U24107 (N_24107,N_20309,N_18868);
xnor U24108 (N_24108,N_20573,N_19301);
nor U24109 (N_24109,N_19604,N_20321);
and U24110 (N_24110,N_19777,N_21484);
or U24111 (N_24111,N_20130,N_20738);
nand U24112 (N_24112,N_19330,N_21345);
or U24113 (N_24113,N_20050,N_21347);
and U24114 (N_24114,N_19958,N_21654);
and U24115 (N_24115,N_19797,N_18897);
xnor U24116 (N_24116,N_21032,N_18777);
or U24117 (N_24117,N_19796,N_19915);
nand U24118 (N_24118,N_21693,N_20618);
nor U24119 (N_24119,N_19279,N_21345);
xnor U24120 (N_24120,N_20700,N_20438);
nor U24121 (N_24121,N_18950,N_21037);
nor U24122 (N_24122,N_18762,N_20375);
nor U24123 (N_24123,N_19075,N_20987);
and U24124 (N_24124,N_19596,N_20785);
or U24125 (N_24125,N_20575,N_20942);
and U24126 (N_24126,N_19262,N_19816);
xnor U24127 (N_24127,N_18899,N_19715);
nand U24128 (N_24128,N_21250,N_19290);
and U24129 (N_24129,N_20669,N_21419);
nand U24130 (N_24130,N_19262,N_20370);
nor U24131 (N_24131,N_21239,N_20752);
nand U24132 (N_24132,N_20186,N_20332);
nand U24133 (N_24133,N_20751,N_20092);
nand U24134 (N_24134,N_21679,N_20388);
nor U24135 (N_24135,N_20978,N_20466);
nor U24136 (N_24136,N_21314,N_20577);
nor U24137 (N_24137,N_20617,N_21668);
nand U24138 (N_24138,N_20959,N_19779);
and U24139 (N_24139,N_18837,N_20284);
and U24140 (N_24140,N_21247,N_20149);
or U24141 (N_24141,N_20290,N_21541);
nand U24142 (N_24142,N_20304,N_19191);
xor U24143 (N_24143,N_21854,N_18850);
nor U24144 (N_24144,N_20280,N_21197);
nand U24145 (N_24145,N_19264,N_20284);
and U24146 (N_24146,N_19974,N_18808);
and U24147 (N_24147,N_20538,N_21474);
nor U24148 (N_24148,N_20583,N_19804);
nand U24149 (N_24149,N_19805,N_21377);
and U24150 (N_24150,N_21112,N_21460);
nor U24151 (N_24151,N_20189,N_19099);
and U24152 (N_24152,N_20763,N_20496);
or U24153 (N_24153,N_20703,N_21194);
nand U24154 (N_24154,N_19853,N_20041);
or U24155 (N_24155,N_19466,N_21431);
xor U24156 (N_24156,N_21127,N_18880);
and U24157 (N_24157,N_19304,N_19072);
xor U24158 (N_24158,N_19705,N_21867);
nand U24159 (N_24159,N_20041,N_20928);
nor U24160 (N_24160,N_20713,N_20270);
and U24161 (N_24161,N_21149,N_19754);
or U24162 (N_24162,N_21812,N_19019);
xor U24163 (N_24163,N_21603,N_20438);
and U24164 (N_24164,N_19497,N_19032);
and U24165 (N_24165,N_21495,N_21864);
nand U24166 (N_24166,N_21588,N_19148);
nor U24167 (N_24167,N_19619,N_19004);
or U24168 (N_24168,N_20376,N_18781);
or U24169 (N_24169,N_21426,N_20704);
or U24170 (N_24170,N_20761,N_19517);
nor U24171 (N_24171,N_20241,N_19565);
xnor U24172 (N_24172,N_21245,N_20817);
and U24173 (N_24173,N_21770,N_18837);
xnor U24174 (N_24174,N_20724,N_18759);
or U24175 (N_24175,N_20119,N_20625);
or U24176 (N_24176,N_19456,N_19629);
nand U24177 (N_24177,N_20917,N_19440);
and U24178 (N_24178,N_20730,N_20264);
and U24179 (N_24179,N_21338,N_19137);
or U24180 (N_24180,N_19816,N_20445);
and U24181 (N_24181,N_19060,N_20366);
xor U24182 (N_24182,N_18957,N_21039);
or U24183 (N_24183,N_21268,N_19311);
nand U24184 (N_24184,N_21650,N_20868);
or U24185 (N_24185,N_19335,N_21297);
and U24186 (N_24186,N_21372,N_21221);
xnor U24187 (N_24187,N_20851,N_20799);
nand U24188 (N_24188,N_21080,N_19477);
or U24189 (N_24189,N_19389,N_21058);
nand U24190 (N_24190,N_20047,N_20926);
nand U24191 (N_24191,N_19979,N_21268);
and U24192 (N_24192,N_21372,N_19793);
nand U24193 (N_24193,N_21699,N_19071);
or U24194 (N_24194,N_20856,N_20841);
nor U24195 (N_24195,N_20044,N_20907);
nand U24196 (N_24196,N_20077,N_20250);
nand U24197 (N_24197,N_20694,N_20405);
xor U24198 (N_24198,N_19392,N_19281);
xor U24199 (N_24199,N_19279,N_20972);
nand U24200 (N_24200,N_21690,N_20355);
xor U24201 (N_24201,N_19652,N_21677);
nor U24202 (N_24202,N_19032,N_20369);
nand U24203 (N_24203,N_20553,N_19008);
nand U24204 (N_24204,N_19534,N_19774);
and U24205 (N_24205,N_21316,N_20781);
nand U24206 (N_24206,N_19803,N_19169);
nand U24207 (N_24207,N_19601,N_19618);
nand U24208 (N_24208,N_21181,N_20304);
xor U24209 (N_24209,N_21873,N_19568);
nor U24210 (N_24210,N_19172,N_20111);
and U24211 (N_24211,N_21003,N_19750);
or U24212 (N_24212,N_21145,N_20409);
xnor U24213 (N_24213,N_19988,N_20272);
xor U24214 (N_24214,N_19528,N_19708);
nor U24215 (N_24215,N_18908,N_19772);
nand U24216 (N_24216,N_20260,N_21550);
nor U24217 (N_24217,N_21443,N_21181);
nand U24218 (N_24218,N_18783,N_19243);
or U24219 (N_24219,N_19588,N_19897);
and U24220 (N_24220,N_20750,N_20321);
and U24221 (N_24221,N_20043,N_19907);
nor U24222 (N_24222,N_21080,N_20605);
nor U24223 (N_24223,N_20340,N_20559);
nor U24224 (N_24224,N_19787,N_20827);
nor U24225 (N_24225,N_21265,N_20755);
nor U24226 (N_24226,N_19252,N_19869);
or U24227 (N_24227,N_21780,N_19928);
nor U24228 (N_24228,N_19312,N_19731);
or U24229 (N_24229,N_21792,N_19059);
xnor U24230 (N_24230,N_20460,N_18811);
or U24231 (N_24231,N_20602,N_19504);
and U24232 (N_24232,N_19098,N_20483);
and U24233 (N_24233,N_19335,N_21182);
and U24234 (N_24234,N_21718,N_21079);
or U24235 (N_24235,N_21377,N_19328);
and U24236 (N_24236,N_18929,N_21266);
nor U24237 (N_24237,N_18803,N_19482);
xor U24238 (N_24238,N_21869,N_19758);
nand U24239 (N_24239,N_18910,N_20418);
nor U24240 (N_24240,N_21390,N_21810);
nand U24241 (N_24241,N_20816,N_20114);
or U24242 (N_24242,N_18974,N_20446);
or U24243 (N_24243,N_21192,N_21165);
nor U24244 (N_24244,N_20499,N_21810);
nor U24245 (N_24245,N_21160,N_20801);
and U24246 (N_24246,N_19260,N_18771);
nand U24247 (N_24247,N_20527,N_19178);
nor U24248 (N_24248,N_20663,N_20766);
nand U24249 (N_24249,N_19213,N_21752);
and U24250 (N_24250,N_21195,N_19343);
or U24251 (N_24251,N_19178,N_20018);
and U24252 (N_24252,N_19149,N_19228);
and U24253 (N_24253,N_21846,N_19476);
xnor U24254 (N_24254,N_18777,N_19323);
nand U24255 (N_24255,N_20254,N_20513);
and U24256 (N_24256,N_18929,N_20668);
or U24257 (N_24257,N_19934,N_20450);
nand U24258 (N_24258,N_20745,N_19267);
or U24259 (N_24259,N_19920,N_20576);
or U24260 (N_24260,N_20742,N_20864);
and U24261 (N_24261,N_20806,N_21435);
nor U24262 (N_24262,N_19336,N_21135);
xnor U24263 (N_24263,N_20884,N_19670);
xor U24264 (N_24264,N_21231,N_20994);
and U24265 (N_24265,N_19198,N_19283);
nor U24266 (N_24266,N_20028,N_21518);
or U24267 (N_24267,N_19270,N_20831);
xor U24268 (N_24268,N_21115,N_21645);
or U24269 (N_24269,N_19693,N_21666);
and U24270 (N_24270,N_18880,N_21018);
or U24271 (N_24271,N_21015,N_21394);
nor U24272 (N_24272,N_18761,N_19956);
xnor U24273 (N_24273,N_21019,N_20954);
and U24274 (N_24274,N_20238,N_19356);
nor U24275 (N_24275,N_19925,N_21207);
and U24276 (N_24276,N_21084,N_21502);
xnor U24277 (N_24277,N_18803,N_18930);
nand U24278 (N_24278,N_20542,N_19332);
nor U24279 (N_24279,N_21540,N_19215);
nand U24280 (N_24280,N_19023,N_20655);
xnor U24281 (N_24281,N_21539,N_20013);
and U24282 (N_24282,N_20631,N_20395);
or U24283 (N_24283,N_19694,N_20147);
xor U24284 (N_24284,N_21311,N_18854);
nand U24285 (N_24285,N_19637,N_20534);
and U24286 (N_24286,N_20622,N_21051);
and U24287 (N_24287,N_19302,N_21057);
xor U24288 (N_24288,N_19003,N_19174);
nor U24289 (N_24289,N_18877,N_20788);
nand U24290 (N_24290,N_21423,N_20011);
xor U24291 (N_24291,N_20583,N_19744);
and U24292 (N_24292,N_18786,N_20068);
or U24293 (N_24293,N_19183,N_21491);
or U24294 (N_24294,N_20824,N_21673);
and U24295 (N_24295,N_18848,N_19441);
nand U24296 (N_24296,N_20948,N_20141);
or U24297 (N_24297,N_19589,N_19398);
nand U24298 (N_24298,N_18952,N_19879);
and U24299 (N_24299,N_21504,N_19648);
xnor U24300 (N_24300,N_18943,N_21532);
xor U24301 (N_24301,N_19177,N_21342);
nand U24302 (N_24302,N_21581,N_20504);
or U24303 (N_24303,N_19767,N_19142);
or U24304 (N_24304,N_19277,N_21287);
and U24305 (N_24305,N_21219,N_18824);
or U24306 (N_24306,N_19454,N_21453);
and U24307 (N_24307,N_19855,N_19097);
nand U24308 (N_24308,N_21328,N_20413);
nand U24309 (N_24309,N_21059,N_20396);
nor U24310 (N_24310,N_19776,N_21093);
xor U24311 (N_24311,N_19150,N_21594);
and U24312 (N_24312,N_20330,N_19718);
and U24313 (N_24313,N_19356,N_20104);
xor U24314 (N_24314,N_19619,N_21400);
or U24315 (N_24315,N_19490,N_20268);
nor U24316 (N_24316,N_19782,N_21145);
or U24317 (N_24317,N_21477,N_19686);
or U24318 (N_24318,N_20395,N_19657);
or U24319 (N_24319,N_20984,N_21100);
nand U24320 (N_24320,N_20623,N_20427);
nor U24321 (N_24321,N_20022,N_20833);
nand U24322 (N_24322,N_20648,N_21599);
or U24323 (N_24323,N_21183,N_21811);
xnor U24324 (N_24324,N_20078,N_20118);
nand U24325 (N_24325,N_20801,N_20494);
nor U24326 (N_24326,N_21855,N_20203);
nor U24327 (N_24327,N_20500,N_20968);
nand U24328 (N_24328,N_21217,N_19725);
xnor U24329 (N_24329,N_20237,N_20351);
xor U24330 (N_24330,N_21503,N_19696);
or U24331 (N_24331,N_19449,N_20389);
xnor U24332 (N_24332,N_20715,N_20653);
xor U24333 (N_24333,N_20996,N_18975);
or U24334 (N_24334,N_20151,N_20200);
xnor U24335 (N_24335,N_19848,N_19729);
and U24336 (N_24336,N_19816,N_21715);
and U24337 (N_24337,N_19286,N_20685);
nand U24338 (N_24338,N_19313,N_21851);
and U24339 (N_24339,N_21147,N_19805);
and U24340 (N_24340,N_19777,N_19455);
xnor U24341 (N_24341,N_21309,N_19154);
or U24342 (N_24342,N_19543,N_19288);
or U24343 (N_24343,N_19031,N_18881);
or U24344 (N_24344,N_19381,N_20161);
or U24345 (N_24345,N_19185,N_21030);
nor U24346 (N_24346,N_21573,N_21040);
xor U24347 (N_24347,N_19513,N_19276);
nor U24348 (N_24348,N_18916,N_20576);
or U24349 (N_24349,N_19774,N_21748);
and U24350 (N_24350,N_19264,N_21022);
xnor U24351 (N_24351,N_20117,N_19273);
or U24352 (N_24352,N_21744,N_19643);
nand U24353 (N_24353,N_19319,N_19330);
xor U24354 (N_24354,N_20042,N_19019);
nand U24355 (N_24355,N_21241,N_20330);
or U24356 (N_24356,N_20620,N_19567);
nand U24357 (N_24357,N_20371,N_20901);
and U24358 (N_24358,N_21354,N_19622);
nand U24359 (N_24359,N_19984,N_21242);
nor U24360 (N_24360,N_21424,N_20041);
and U24361 (N_24361,N_18884,N_20423);
or U24362 (N_24362,N_21380,N_21050);
or U24363 (N_24363,N_19442,N_18779);
nor U24364 (N_24364,N_20882,N_20940);
or U24365 (N_24365,N_19861,N_19903);
nand U24366 (N_24366,N_20585,N_21352);
xnor U24367 (N_24367,N_20327,N_19920);
xor U24368 (N_24368,N_20724,N_21022);
nor U24369 (N_24369,N_20314,N_21488);
nor U24370 (N_24370,N_20913,N_21360);
nand U24371 (N_24371,N_19493,N_19425);
xor U24372 (N_24372,N_19126,N_20309);
nand U24373 (N_24373,N_18951,N_20245);
nor U24374 (N_24374,N_18879,N_19232);
and U24375 (N_24375,N_21031,N_19726);
xnor U24376 (N_24376,N_21447,N_19339);
nand U24377 (N_24377,N_21686,N_20459);
nor U24378 (N_24378,N_20718,N_20153);
nand U24379 (N_24379,N_19532,N_19733);
and U24380 (N_24380,N_21473,N_20446);
nor U24381 (N_24381,N_18883,N_19588);
nand U24382 (N_24382,N_19449,N_18994);
or U24383 (N_24383,N_20290,N_19063);
or U24384 (N_24384,N_21392,N_20094);
nor U24385 (N_24385,N_19449,N_19359);
nand U24386 (N_24386,N_21557,N_20214);
nor U24387 (N_24387,N_21327,N_21117);
or U24388 (N_24388,N_18934,N_20723);
or U24389 (N_24389,N_18984,N_20166);
nand U24390 (N_24390,N_19327,N_21481);
nor U24391 (N_24391,N_18943,N_19627);
nor U24392 (N_24392,N_19180,N_18827);
and U24393 (N_24393,N_19555,N_18939);
xor U24394 (N_24394,N_21144,N_20270);
xnor U24395 (N_24395,N_20581,N_20515);
nand U24396 (N_24396,N_20354,N_21541);
xnor U24397 (N_24397,N_18888,N_21153);
nor U24398 (N_24398,N_20150,N_20731);
and U24399 (N_24399,N_20669,N_19253);
and U24400 (N_24400,N_19614,N_21548);
nor U24401 (N_24401,N_19750,N_19933);
or U24402 (N_24402,N_21739,N_18963);
xor U24403 (N_24403,N_21539,N_21421);
and U24404 (N_24404,N_20263,N_21332);
or U24405 (N_24405,N_20593,N_21611);
xnor U24406 (N_24406,N_20231,N_18879);
nand U24407 (N_24407,N_20527,N_21869);
nand U24408 (N_24408,N_20703,N_21484);
nor U24409 (N_24409,N_21096,N_19840);
and U24410 (N_24410,N_21389,N_21810);
xor U24411 (N_24411,N_20690,N_20861);
or U24412 (N_24412,N_19020,N_19967);
nor U24413 (N_24413,N_21008,N_21110);
and U24414 (N_24414,N_19144,N_19695);
xnor U24415 (N_24415,N_21674,N_21311);
xnor U24416 (N_24416,N_19275,N_20670);
xnor U24417 (N_24417,N_21614,N_20176);
xor U24418 (N_24418,N_19052,N_20601);
xor U24419 (N_24419,N_20608,N_21282);
nor U24420 (N_24420,N_19221,N_20593);
or U24421 (N_24421,N_21150,N_19779);
and U24422 (N_24422,N_19838,N_20619);
nor U24423 (N_24423,N_20477,N_20191);
nand U24424 (N_24424,N_19582,N_21254);
nor U24425 (N_24425,N_19867,N_20189);
nand U24426 (N_24426,N_20162,N_19112);
xor U24427 (N_24427,N_21821,N_19530);
nor U24428 (N_24428,N_20380,N_21424);
or U24429 (N_24429,N_19859,N_19953);
nand U24430 (N_24430,N_18795,N_20994);
or U24431 (N_24431,N_19195,N_19279);
nor U24432 (N_24432,N_21399,N_21359);
xnor U24433 (N_24433,N_19050,N_21294);
or U24434 (N_24434,N_19373,N_20802);
and U24435 (N_24435,N_21442,N_18963);
xor U24436 (N_24436,N_18917,N_21653);
nor U24437 (N_24437,N_21401,N_20881);
and U24438 (N_24438,N_20752,N_18847);
xor U24439 (N_24439,N_21872,N_20780);
or U24440 (N_24440,N_19639,N_21263);
or U24441 (N_24441,N_19022,N_19842);
nor U24442 (N_24442,N_20790,N_21342);
or U24443 (N_24443,N_19947,N_20692);
xor U24444 (N_24444,N_20767,N_20873);
nor U24445 (N_24445,N_20816,N_21528);
or U24446 (N_24446,N_19462,N_20720);
xnor U24447 (N_24447,N_18963,N_21308);
or U24448 (N_24448,N_19932,N_20246);
xnor U24449 (N_24449,N_21421,N_20501);
and U24450 (N_24450,N_20366,N_18968);
nand U24451 (N_24451,N_21737,N_21516);
and U24452 (N_24452,N_20737,N_21497);
or U24453 (N_24453,N_20217,N_20548);
nor U24454 (N_24454,N_19241,N_19583);
and U24455 (N_24455,N_21282,N_21059);
nor U24456 (N_24456,N_21736,N_19003);
or U24457 (N_24457,N_19628,N_19231);
nor U24458 (N_24458,N_19191,N_21208);
nor U24459 (N_24459,N_19720,N_19617);
nand U24460 (N_24460,N_21637,N_20960);
xor U24461 (N_24461,N_21778,N_21131);
nand U24462 (N_24462,N_19695,N_18821);
and U24463 (N_24463,N_20080,N_21470);
nand U24464 (N_24464,N_20609,N_21151);
nor U24465 (N_24465,N_19396,N_21539);
or U24466 (N_24466,N_21513,N_20724);
or U24467 (N_24467,N_19644,N_19958);
nor U24468 (N_24468,N_20319,N_19502);
xor U24469 (N_24469,N_19508,N_21358);
and U24470 (N_24470,N_19351,N_21486);
nand U24471 (N_24471,N_20763,N_20343);
nand U24472 (N_24472,N_20631,N_21459);
nand U24473 (N_24473,N_21507,N_18979);
or U24474 (N_24474,N_21360,N_21610);
nor U24475 (N_24475,N_19556,N_19413);
nand U24476 (N_24476,N_20581,N_19776);
or U24477 (N_24477,N_21785,N_18972);
or U24478 (N_24478,N_19081,N_19457);
and U24479 (N_24479,N_21530,N_18822);
nor U24480 (N_24480,N_21720,N_19849);
nand U24481 (N_24481,N_19942,N_20202);
and U24482 (N_24482,N_20387,N_21625);
and U24483 (N_24483,N_19488,N_21177);
nor U24484 (N_24484,N_21593,N_21557);
or U24485 (N_24485,N_21306,N_21207);
xnor U24486 (N_24486,N_21505,N_19135);
nor U24487 (N_24487,N_20542,N_20598);
nand U24488 (N_24488,N_21608,N_21355);
xor U24489 (N_24489,N_19364,N_21838);
nand U24490 (N_24490,N_20689,N_20180);
or U24491 (N_24491,N_20628,N_19750);
and U24492 (N_24492,N_20889,N_19705);
or U24493 (N_24493,N_19971,N_21533);
xor U24494 (N_24494,N_21240,N_19070);
nand U24495 (N_24495,N_20516,N_19571);
or U24496 (N_24496,N_20789,N_20388);
or U24497 (N_24497,N_21516,N_19823);
nand U24498 (N_24498,N_21014,N_19734);
nor U24499 (N_24499,N_20610,N_20055);
and U24500 (N_24500,N_20778,N_19946);
nor U24501 (N_24501,N_21412,N_19194);
xnor U24502 (N_24502,N_21598,N_19539);
nand U24503 (N_24503,N_21513,N_21300);
xnor U24504 (N_24504,N_18858,N_21569);
and U24505 (N_24505,N_20216,N_20057);
nor U24506 (N_24506,N_21294,N_19938);
and U24507 (N_24507,N_18920,N_19558);
xor U24508 (N_24508,N_21069,N_19954);
nor U24509 (N_24509,N_21692,N_18765);
nand U24510 (N_24510,N_19036,N_19967);
xor U24511 (N_24511,N_19805,N_20661);
or U24512 (N_24512,N_20161,N_18771);
xnor U24513 (N_24513,N_19147,N_19174);
or U24514 (N_24514,N_19774,N_20622);
xnor U24515 (N_24515,N_19890,N_19822);
nor U24516 (N_24516,N_19997,N_21754);
nand U24517 (N_24517,N_19857,N_20237);
and U24518 (N_24518,N_18801,N_19766);
xnor U24519 (N_24519,N_19126,N_19035);
nor U24520 (N_24520,N_21022,N_18833);
nor U24521 (N_24521,N_21497,N_21189);
nor U24522 (N_24522,N_20525,N_19377);
xnor U24523 (N_24523,N_21516,N_19479);
nor U24524 (N_24524,N_18993,N_18884);
and U24525 (N_24525,N_20750,N_21626);
and U24526 (N_24526,N_21755,N_19242);
xnor U24527 (N_24527,N_19224,N_20820);
xor U24528 (N_24528,N_21405,N_20965);
or U24529 (N_24529,N_19880,N_18782);
nand U24530 (N_24530,N_20269,N_20620);
or U24531 (N_24531,N_20088,N_21682);
and U24532 (N_24532,N_21469,N_20602);
and U24533 (N_24533,N_21429,N_21589);
and U24534 (N_24534,N_21161,N_19638);
or U24535 (N_24535,N_20685,N_20155);
xnor U24536 (N_24536,N_20560,N_20004);
nor U24537 (N_24537,N_19479,N_21847);
xnor U24538 (N_24538,N_21811,N_18968);
and U24539 (N_24539,N_20314,N_21443);
nand U24540 (N_24540,N_21808,N_19491);
nand U24541 (N_24541,N_19052,N_19915);
and U24542 (N_24542,N_19349,N_20648);
nor U24543 (N_24543,N_21125,N_21142);
or U24544 (N_24544,N_19849,N_19447);
xnor U24545 (N_24545,N_19563,N_19543);
or U24546 (N_24546,N_18836,N_19891);
nor U24547 (N_24547,N_20748,N_20227);
nand U24548 (N_24548,N_21863,N_19760);
and U24549 (N_24549,N_21662,N_19087);
and U24550 (N_24550,N_21507,N_20317);
nand U24551 (N_24551,N_21010,N_20919);
nor U24552 (N_24552,N_19921,N_20832);
nor U24553 (N_24553,N_20409,N_19386);
nor U24554 (N_24554,N_18781,N_18894);
and U24555 (N_24555,N_18983,N_19138);
nor U24556 (N_24556,N_20781,N_21471);
and U24557 (N_24557,N_21344,N_19203);
or U24558 (N_24558,N_21356,N_19010);
xnor U24559 (N_24559,N_21303,N_21123);
or U24560 (N_24560,N_21293,N_21090);
or U24561 (N_24561,N_21862,N_20938);
or U24562 (N_24562,N_20398,N_21517);
and U24563 (N_24563,N_19536,N_21433);
and U24564 (N_24564,N_21621,N_21006);
nor U24565 (N_24565,N_21012,N_21260);
or U24566 (N_24566,N_20829,N_18998);
xnor U24567 (N_24567,N_20792,N_19134);
nand U24568 (N_24568,N_21287,N_21551);
nand U24569 (N_24569,N_21450,N_20281);
nand U24570 (N_24570,N_19865,N_19905);
xnor U24571 (N_24571,N_21383,N_20824);
and U24572 (N_24572,N_19092,N_19879);
nor U24573 (N_24573,N_20360,N_20649);
xor U24574 (N_24574,N_18992,N_19305);
or U24575 (N_24575,N_20066,N_19191);
and U24576 (N_24576,N_21803,N_19042);
nand U24577 (N_24577,N_21546,N_20136);
nand U24578 (N_24578,N_20599,N_21105);
nor U24579 (N_24579,N_20797,N_20350);
nor U24580 (N_24580,N_19186,N_21187);
nand U24581 (N_24581,N_20648,N_21030);
and U24582 (N_24582,N_21692,N_20525);
xnor U24583 (N_24583,N_21196,N_20052);
and U24584 (N_24584,N_21649,N_21173);
nand U24585 (N_24585,N_19897,N_21211);
xnor U24586 (N_24586,N_19844,N_19790);
or U24587 (N_24587,N_21465,N_19027);
nand U24588 (N_24588,N_19185,N_19353);
and U24589 (N_24589,N_21540,N_21115);
nor U24590 (N_24590,N_19937,N_19277);
nor U24591 (N_24591,N_19990,N_20002);
and U24592 (N_24592,N_19483,N_20630);
nand U24593 (N_24593,N_20487,N_20004);
or U24594 (N_24594,N_19700,N_19923);
or U24595 (N_24595,N_18762,N_20657);
nand U24596 (N_24596,N_20772,N_20250);
nor U24597 (N_24597,N_19519,N_19605);
nand U24598 (N_24598,N_20986,N_21538);
nor U24599 (N_24599,N_20387,N_19204);
nor U24600 (N_24600,N_20272,N_21535);
nand U24601 (N_24601,N_19698,N_20316);
nand U24602 (N_24602,N_20862,N_20991);
nand U24603 (N_24603,N_19104,N_19719);
and U24604 (N_24604,N_21520,N_19346);
nand U24605 (N_24605,N_19430,N_20024);
xor U24606 (N_24606,N_20287,N_19207);
or U24607 (N_24607,N_21086,N_18972);
nand U24608 (N_24608,N_20926,N_21271);
and U24609 (N_24609,N_20875,N_20395);
xnor U24610 (N_24610,N_20445,N_21776);
xor U24611 (N_24611,N_20478,N_19377);
or U24612 (N_24612,N_21828,N_21170);
nand U24613 (N_24613,N_21161,N_21152);
nor U24614 (N_24614,N_21299,N_21374);
xnor U24615 (N_24615,N_19975,N_18853);
xnor U24616 (N_24616,N_21844,N_20033);
nor U24617 (N_24617,N_19480,N_21210);
and U24618 (N_24618,N_20684,N_19825);
xnor U24619 (N_24619,N_20199,N_19144);
nor U24620 (N_24620,N_21049,N_18992);
and U24621 (N_24621,N_18803,N_19557);
and U24622 (N_24622,N_19525,N_20882);
nand U24623 (N_24623,N_20124,N_19892);
and U24624 (N_24624,N_18849,N_20352);
nor U24625 (N_24625,N_18951,N_21689);
nor U24626 (N_24626,N_18937,N_21488);
nor U24627 (N_24627,N_19638,N_18982);
nor U24628 (N_24628,N_19818,N_20785);
xor U24629 (N_24629,N_19210,N_19725);
and U24630 (N_24630,N_18899,N_19492);
and U24631 (N_24631,N_19106,N_20491);
or U24632 (N_24632,N_21385,N_21513);
nand U24633 (N_24633,N_19443,N_21826);
nor U24634 (N_24634,N_21688,N_21132);
xnor U24635 (N_24635,N_19182,N_21462);
and U24636 (N_24636,N_21026,N_20316);
nor U24637 (N_24637,N_19131,N_19792);
xnor U24638 (N_24638,N_20720,N_21397);
xor U24639 (N_24639,N_20655,N_19513);
nor U24640 (N_24640,N_18977,N_18892);
and U24641 (N_24641,N_18846,N_20945);
and U24642 (N_24642,N_19049,N_21584);
xnor U24643 (N_24643,N_21026,N_19691);
and U24644 (N_24644,N_18851,N_19925);
and U24645 (N_24645,N_21789,N_19485);
or U24646 (N_24646,N_21401,N_21408);
or U24647 (N_24647,N_21728,N_19383);
nand U24648 (N_24648,N_20986,N_21405);
or U24649 (N_24649,N_21362,N_18935);
xor U24650 (N_24650,N_18939,N_19886);
and U24651 (N_24651,N_19399,N_18923);
or U24652 (N_24652,N_20536,N_20563);
or U24653 (N_24653,N_21145,N_20411);
nand U24654 (N_24654,N_21370,N_19120);
or U24655 (N_24655,N_21527,N_20343);
xor U24656 (N_24656,N_21524,N_20617);
or U24657 (N_24657,N_19782,N_19212);
xnor U24658 (N_24658,N_21415,N_19228);
or U24659 (N_24659,N_19006,N_20759);
nand U24660 (N_24660,N_20660,N_20968);
or U24661 (N_24661,N_19651,N_20300);
nor U24662 (N_24662,N_21805,N_21302);
and U24663 (N_24663,N_19149,N_18763);
nor U24664 (N_24664,N_19888,N_20710);
nor U24665 (N_24665,N_19705,N_19481);
xnor U24666 (N_24666,N_18816,N_18803);
xnor U24667 (N_24667,N_21420,N_21352);
nand U24668 (N_24668,N_21231,N_21258);
nor U24669 (N_24669,N_21313,N_20847);
and U24670 (N_24670,N_19116,N_20786);
nor U24671 (N_24671,N_19306,N_19819);
or U24672 (N_24672,N_19534,N_20938);
or U24673 (N_24673,N_20987,N_20962);
xor U24674 (N_24674,N_20962,N_19073);
and U24675 (N_24675,N_19795,N_19381);
nand U24676 (N_24676,N_20437,N_20782);
and U24677 (N_24677,N_19391,N_19830);
and U24678 (N_24678,N_20016,N_20136);
nor U24679 (N_24679,N_19370,N_18888);
and U24680 (N_24680,N_21671,N_19552);
or U24681 (N_24681,N_20608,N_21640);
nor U24682 (N_24682,N_20372,N_21197);
xnor U24683 (N_24683,N_19333,N_21099);
nor U24684 (N_24684,N_19585,N_19437);
nand U24685 (N_24685,N_19727,N_20306);
nand U24686 (N_24686,N_19071,N_21113);
and U24687 (N_24687,N_19783,N_20105);
or U24688 (N_24688,N_20392,N_18820);
nor U24689 (N_24689,N_20058,N_21304);
xor U24690 (N_24690,N_20635,N_20004);
nor U24691 (N_24691,N_20297,N_19126);
nor U24692 (N_24692,N_18935,N_20997);
nor U24693 (N_24693,N_20026,N_20601);
nand U24694 (N_24694,N_20585,N_19969);
and U24695 (N_24695,N_21780,N_20011);
or U24696 (N_24696,N_21058,N_19248);
or U24697 (N_24697,N_18957,N_19874);
or U24698 (N_24698,N_20742,N_20541);
and U24699 (N_24699,N_18786,N_20425);
xnor U24700 (N_24700,N_19782,N_21420);
or U24701 (N_24701,N_19119,N_21618);
nor U24702 (N_24702,N_21236,N_19883);
or U24703 (N_24703,N_20932,N_18904);
xnor U24704 (N_24704,N_21670,N_20767);
and U24705 (N_24705,N_19308,N_19396);
xor U24706 (N_24706,N_19324,N_18889);
xor U24707 (N_24707,N_20173,N_20278);
nand U24708 (N_24708,N_20197,N_18840);
and U24709 (N_24709,N_20783,N_20041);
xor U24710 (N_24710,N_19379,N_19547);
and U24711 (N_24711,N_19331,N_20265);
xor U24712 (N_24712,N_18992,N_20648);
nor U24713 (N_24713,N_21684,N_19342);
xor U24714 (N_24714,N_21400,N_21599);
xor U24715 (N_24715,N_21257,N_21188);
and U24716 (N_24716,N_18806,N_19913);
xor U24717 (N_24717,N_20880,N_20440);
nor U24718 (N_24718,N_19912,N_19535);
xor U24719 (N_24719,N_21002,N_20075);
nand U24720 (N_24720,N_18801,N_20506);
and U24721 (N_24721,N_21840,N_19289);
nor U24722 (N_24722,N_21396,N_21631);
nand U24723 (N_24723,N_21489,N_20319);
nand U24724 (N_24724,N_19707,N_18789);
or U24725 (N_24725,N_21201,N_20509);
nor U24726 (N_24726,N_18807,N_20197);
nor U24727 (N_24727,N_20127,N_21269);
nand U24728 (N_24728,N_19993,N_21467);
xor U24729 (N_24729,N_20894,N_20670);
and U24730 (N_24730,N_20270,N_20540);
nand U24731 (N_24731,N_19823,N_19074);
nand U24732 (N_24732,N_19325,N_21248);
and U24733 (N_24733,N_20467,N_20718);
nor U24734 (N_24734,N_20360,N_18875);
nand U24735 (N_24735,N_20262,N_19839);
or U24736 (N_24736,N_20811,N_18892);
or U24737 (N_24737,N_21440,N_19966);
or U24738 (N_24738,N_20178,N_20283);
and U24739 (N_24739,N_20162,N_18831);
and U24740 (N_24740,N_21172,N_20493);
nand U24741 (N_24741,N_20479,N_20280);
nor U24742 (N_24742,N_19661,N_21084);
xnor U24743 (N_24743,N_20985,N_19731);
and U24744 (N_24744,N_19391,N_20806);
or U24745 (N_24745,N_20289,N_20758);
nor U24746 (N_24746,N_20745,N_21760);
nor U24747 (N_24747,N_18899,N_21262);
and U24748 (N_24748,N_19846,N_20188);
xnor U24749 (N_24749,N_21019,N_21809);
nor U24750 (N_24750,N_19264,N_19522);
nand U24751 (N_24751,N_20320,N_21605);
or U24752 (N_24752,N_19835,N_20735);
nand U24753 (N_24753,N_20948,N_21735);
nand U24754 (N_24754,N_20421,N_19220);
xor U24755 (N_24755,N_20180,N_19192);
xnor U24756 (N_24756,N_21373,N_20131);
or U24757 (N_24757,N_21191,N_20137);
nor U24758 (N_24758,N_19458,N_20942);
xor U24759 (N_24759,N_20389,N_19476);
and U24760 (N_24760,N_20076,N_20675);
nor U24761 (N_24761,N_19147,N_21437);
or U24762 (N_24762,N_21688,N_19941);
and U24763 (N_24763,N_21703,N_19451);
nand U24764 (N_24764,N_20232,N_19211);
or U24765 (N_24765,N_19836,N_20117);
nand U24766 (N_24766,N_21743,N_21071);
or U24767 (N_24767,N_20776,N_19784);
and U24768 (N_24768,N_20040,N_19870);
nand U24769 (N_24769,N_19363,N_19662);
nor U24770 (N_24770,N_21770,N_21081);
xor U24771 (N_24771,N_20702,N_19034);
or U24772 (N_24772,N_20561,N_20545);
nor U24773 (N_24773,N_21873,N_19361);
nand U24774 (N_24774,N_19161,N_20240);
nand U24775 (N_24775,N_21507,N_20506);
nand U24776 (N_24776,N_21329,N_21514);
nor U24777 (N_24777,N_20293,N_21413);
nor U24778 (N_24778,N_19441,N_19961);
and U24779 (N_24779,N_18776,N_19014);
and U24780 (N_24780,N_19393,N_19366);
nand U24781 (N_24781,N_21383,N_18779);
nor U24782 (N_24782,N_21452,N_20806);
nor U24783 (N_24783,N_19663,N_20885);
nand U24784 (N_24784,N_19590,N_21642);
nand U24785 (N_24785,N_20232,N_21477);
and U24786 (N_24786,N_21511,N_19382);
or U24787 (N_24787,N_20898,N_21712);
nand U24788 (N_24788,N_19786,N_20014);
and U24789 (N_24789,N_21704,N_19387);
or U24790 (N_24790,N_20342,N_21184);
and U24791 (N_24791,N_20198,N_21554);
nor U24792 (N_24792,N_20661,N_20190);
nand U24793 (N_24793,N_21204,N_20042);
or U24794 (N_24794,N_21783,N_19601);
nor U24795 (N_24795,N_19374,N_18971);
or U24796 (N_24796,N_21492,N_20359);
nor U24797 (N_24797,N_21672,N_20530);
nor U24798 (N_24798,N_18938,N_19352);
and U24799 (N_24799,N_18931,N_19751);
nand U24800 (N_24800,N_20368,N_20488);
or U24801 (N_24801,N_19114,N_21680);
nand U24802 (N_24802,N_20607,N_20785);
xor U24803 (N_24803,N_18802,N_20433);
and U24804 (N_24804,N_19000,N_21180);
or U24805 (N_24805,N_19198,N_20369);
nor U24806 (N_24806,N_21237,N_19200);
xnor U24807 (N_24807,N_20362,N_20809);
or U24808 (N_24808,N_20550,N_19878);
or U24809 (N_24809,N_19259,N_19154);
nand U24810 (N_24810,N_20843,N_19006);
and U24811 (N_24811,N_19919,N_18965);
and U24812 (N_24812,N_20847,N_19879);
or U24813 (N_24813,N_20770,N_19836);
nand U24814 (N_24814,N_19138,N_21602);
nand U24815 (N_24815,N_19374,N_19950);
or U24816 (N_24816,N_20167,N_20025);
xor U24817 (N_24817,N_21550,N_20689);
or U24818 (N_24818,N_19662,N_20073);
or U24819 (N_24819,N_19235,N_19823);
xor U24820 (N_24820,N_21543,N_19916);
and U24821 (N_24821,N_20261,N_20110);
and U24822 (N_24822,N_20206,N_20290);
nand U24823 (N_24823,N_20726,N_18812);
nor U24824 (N_24824,N_19419,N_20738);
and U24825 (N_24825,N_21456,N_19401);
nor U24826 (N_24826,N_20304,N_18890);
nand U24827 (N_24827,N_20743,N_20190);
nand U24828 (N_24828,N_18755,N_19817);
or U24829 (N_24829,N_21243,N_19865);
xor U24830 (N_24830,N_20552,N_19344);
or U24831 (N_24831,N_19259,N_21717);
or U24832 (N_24832,N_19590,N_19203);
or U24833 (N_24833,N_20120,N_20573);
nand U24834 (N_24834,N_21736,N_20211);
or U24835 (N_24835,N_19354,N_20267);
nor U24836 (N_24836,N_21382,N_19596);
xor U24837 (N_24837,N_19957,N_20611);
and U24838 (N_24838,N_18793,N_18794);
xor U24839 (N_24839,N_20859,N_19851);
nand U24840 (N_24840,N_19542,N_19096);
nand U24841 (N_24841,N_19994,N_19829);
nor U24842 (N_24842,N_20792,N_20198);
and U24843 (N_24843,N_21420,N_20492);
and U24844 (N_24844,N_21573,N_20155);
nand U24845 (N_24845,N_19761,N_21563);
and U24846 (N_24846,N_21649,N_21262);
or U24847 (N_24847,N_19036,N_20229);
or U24848 (N_24848,N_19836,N_19142);
nand U24849 (N_24849,N_21004,N_19258);
or U24850 (N_24850,N_21385,N_19505);
and U24851 (N_24851,N_19975,N_19560);
nand U24852 (N_24852,N_19064,N_21231);
nor U24853 (N_24853,N_20746,N_18758);
nor U24854 (N_24854,N_18976,N_20413);
nand U24855 (N_24855,N_20713,N_21232);
nand U24856 (N_24856,N_20188,N_20444);
and U24857 (N_24857,N_18884,N_20597);
xor U24858 (N_24858,N_21373,N_20514);
and U24859 (N_24859,N_20034,N_20498);
xnor U24860 (N_24860,N_20951,N_21190);
nor U24861 (N_24861,N_20792,N_19753);
nand U24862 (N_24862,N_21298,N_18944);
or U24863 (N_24863,N_19115,N_21005);
nor U24864 (N_24864,N_18863,N_21550);
xor U24865 (N_24865,N_20456,N_19231);
or U24866 (N_24866,N_20806,N_20319);
nand U24867 (N_24867,N_21570,N_21482);
and U24868 (N_24868,N_19381,N_20705);
and U24869 (N_24869,N_18830,N_20628);
nor U24870 (N_24870,N_20774,N_21610);
nor U24871 (N_24871,N_19434,N_20975);
nand U24872 (N_24872,N_20792,N_21159);
nor U24873 (N_24873,N_20626,N_21508);
xnor U24874 (N_24874,N_20151,N_21032);
nor U24875 (N_24875,N_20090,N_21725);
and U24876 (N_24876,N_20601,N_19544);
nor U24877 (N_24877,N_18756,N_20199);
and U24878 (N_24878,N_21473,N_19806);
nand U24879 (N_24879,N_21058,N_21405);
and U24880 (N_24880,N_20602,N_21582);
xor U24881 (N_24881,N_21391,N_18999);
xor U24882 (N_24882,N_20323,N_21758);
nand U24883 (N_24883,N_18966,N_21129);
or U24884 (N_24884,N_21107,N_20568);
xor U24885 (N_24885,N_21822,N_21250);
or U24886 (N_24886,N_20776,N_20998);
nand U24887 (N_24887,N_21829,N_19721);
and U24888 (N_24888,N_19620,N_19784);
or U24889 (N_24889,N_20988,N_19988);
or U24890 (N_24890,N_19935,N_20670);
and U24891 (N_24891,N_20436,N_21254);
nor U24892 (N_24892,N_20845,N_19248);
or U24893 (N_24893,N_21800,N_21133);
nor U24894 (N_24894,N_20984,N_19190);
nand U24895 (N_24895,N_21468,N_20177);
nor U24896 (N_24896,N_21399,N_21842);
or U24897 (N_24897,N_19027,N_20285);
nand U24898 (N_24898,N_21612,N_19014);
xnor U24899 (N_24899,N_21194,N_21088);
nor U24900 (N_24900,N_21611,N_19708);
and U24901 (N_24901,N_21309,N_20903);
nand U24902 (N_24902,N_20573,N_19299);
or U24903 (N_24903,N_19243,N_21731);
and U24904 (N_24904,N_21655,N_20238);
nand U24905 (N_24905,N_19506,N_21840);
nor U24906 (N_24906,N_20821,N_19555);
or U24907 (N_24907,N_21347,N_21823);
nor U24908 (N_24908,N_19637,N_20773);
or U24909 (N_24909,N_21588,N_21791);
nand U24910 (N_24910,N_19910,N_19416);
and U24911 (N_24911,N_19397,N_21840);
and U24912 (N_24912,N_19994,N_19196);
nand U24913 (N_24913,N_19228,N_21475);
and U24914 (N_24914,N_19040,N_19898);
nand U24915 (N_24915,N_18932,N_19965);
and U24916 (N_24916,N_20482,N_19090);
or U24917 (N_24917,N_19812,N_19071);
xor U24918 (N_24918,N_18944,N_19695);
or U24919 (N_24919,N_19620,N_18988);
and U24920 (N_24920,N_20093,N_20795);
and U24921 (N_24921,N_19809,N_19807);
and U24922 (N_24922,N_21817,N_18823);
and U24923 (N_24923,N_20963,N_21755);
nor U24924 (N_24924,N_20691,N_19552);
nand U24925 (N_24925,N_20611,N_19551);
nor U24926 (N_24926,N_19855,N_19040);
and U24927 (N_24927,N_20506,N_20209);
or U24928 (N_24928,N_21353,N_19865);
xor U24929 (N_24929,N_21485,N_19511);
xor U24930 (N_24930,N_20361,N_20927);
and U24931 (N_24931,N_21507,N_18939);
and U24932 (N_24932,N_19420,N_19935);
and U24933 (N_24933,N_18881,N_19494);
nor U24934 (N_24934,N_20660,N_21342);
nor U24935 (N_24935,N_20640,N_21281);
nor U24936 (N_24936,N_19843,N_21552);
or U24937 (N_24937,N_21677,N_21079);
xor U24938 (N_24938,N_20694,N_20099);
xnor U24939 (N_24939,N_21452,N_20596);
or U24940 (N_24940,N_21779,N_20393);
nand U24941 (N_24941,N_21866,N_18803);
xor U24942 (N_24942,N_19274,N_20524);
nand U24943 (N_24943,N_19100,N_21068);
nor U24944 (N_24944,N_19391,N_19153);
or U24945 (N_24945,N_19160,N_19057);
and U24946 (N_24946,N_20940,N_19292);
nor U24947 (N_24947,N_19329,N_20904);
nor U24948 (N_24948,N_19185,N_21209);
xor U24949 (N_24949,N_20816,N_21307);
or U24950 (N_24950,N_20106,N_19071);
nor U24951 (N_24951,N_20559,N_20839);
xnor U24952 (N_24952,N_19207,N_20478);
and U24953 (N_24953,N_18974,N_19075);
nor U24954 (N_24954,N_20532,N_20753);
or U24955 (N_24955,N_20588,N_19521);
or U24956 (N_24956,N_21621,N_21507);
xnor U24957 (N_24957,N_19495,N_21210);
nor U24958 (N_24958,N_19967,N_21271);
xnor U24959 (N_24959,N_21194,N_20769);
xor U24960 (N_24960,N_21848,N_21689);
or U24961 (N_24961,N_19121,N_18955);
nor U24962 (N_24962,N_20981,N_20315);
and U24963 (N_24963,N_21809,N_19932);
or U24964 (N_24964,N_19201,N_20376);
and U24965 (N_24965,N_20743,N_19086);
and U24966 (N_24966,N_20282,N_18940);
nor U24967 (N_24967,N_21466,N_21260);
xor U24968 (N_24968,N_20685,N_21194);
or U24969 (N_24969,N_19367,N_20037);
or U24970 (N_24970,N_20389,N_18912);
xnor U24971 (N_24971,N_20965,N_21279);
nor U24972 (N_24972,N_19542,N_20060);
or U24973 (N_24973,N_20395,N_19827);
nor U24974 (N_24974,N_20626,N_21384);
and U24975 (N_24975,N_19013,N_19465);
and U24976 (N_24976,N_19593,N_18807);
nor U24977 (N_24977,N_21193,N_19927);
xnor U24978 (N_24978,N_21590,N_21198);
or U24979 (N_24979,N_20178,N_20191);
or U24980 (N_24980,N_20444,N_20209);
nor U24981 (N_24981,N_20691,N_20847);
and U24982 (N_24982,N_21181,N_18797);
or U24983 (N_24983,N_21003,N_19130);
nand U24984 (N_24984,N_19562,N_20098);
nor U24985 (N_24985,N_20697,N_18879);
nand U24986 (N_24986,N_21373,N_19393);
or U24987 (N_24987,N_21316,N_21324);
nor U24988 (N_24988,N_21536,N_20525);
or U24989 (N_24989,N_19037,N_20497);
and U24990 (N_24990,N_18858,N_19894);
xor U24991 (N_24991,N_19669,N_21115);
and U24992 (N_24992,N_21744,N_21245);
and U24993 (N_24993,N_21758,N_19524);
or U24994 (N_24994,N_20431,N_18896);
and U24995 (N_24995,N_20343,N_18862);
or U24996 (N_24996,N_19535,N_21383);
nand U24997 (N_24997,N_21706,N_20200);
xor U24998 (N_24998,N_19402,N_20821);
nor U24999 (N_24999,N_18759,N_21073);
nor UO_0 (O_0,N_22308,N_22791);
xor UO_1 (O_1,N_24159,N_22919);
or UO_2 (O_2,N_23619,N_23846);
and UO_3 (O_3,N_22824,N_23652);
nor UO_4 (O_4,N_24344,N_23906);
xnor UO_5 (O_5,N_24503,N_24477);
and UO_6 (O_6,N_22306,N_23792);
xnor UO_7 (O_7,N_23279,N_23734);
nand UO_8 (O_8,N_22804,N_23845);
nand UO_9 (O_9,N_24686,N_23932);
xnor UO_10 (O_10,N_24571,N_23746);
xor UO_11 (O_11,N_24306,N_24094);
or UO_12 (O_12,N_22938,N_22632);
nand UO_13 (O_13,N_22433,N_22013);
or UO_14 (O_14,N_23120,N_23199);
or UO_15 (O_15,N_23991,N_23320);
xor UO_16 (O_16,N_24209,N_23851);
nand UO_17 (O_17,N_22134,N_23291);
and UO_18 (O_18,N_24546,N_23166);
and UO_19 (O_19,N_21877,N_22450);
nand UO_20 (O_20,N_22086,N_22878);
and UO_21 (O_21,N_23295,N_22302);
and UO_22 (O_22,N_23357,N_23569);
and UO_23 (O_23,N_24163,N_24877);
xor UO_24 (O_24,N_24239,N_21986);
nand UO_25 (O_25,N_24823,N_24088);
and UO_26 (O_26,N_23340,N_23171);
nand UO_27 (O_27,N_24573,N_23159);
xor UO_28 (O_28,N_22096,N_22376);
xnor UO_29 (O_29,N_24814,N_24966);
nor UO_30 (O_30,N_23406,N_22137);
xnor UO_31 (O_31,N_24915,N_22538);
and UO_32 (O_32,N_23049,N_24384);
nor UO_33 (O_33,N_23859,N_22975);
nand UO_34 (O_34,N_22158,N_24086);
nand UO_35 (O_35,N_21911,N_22546);
nor UO_36 (O_36,N_24023,N_24143);
nand UO_37 (O_37,N_22265,N_22423);
and UO_38 (O_38,N_21957,N_23980);
nor UO_39 (O_39,N_22602,N_22464);
nand UO_40 (O_40,N_22823,N_23894);
xnor UO_41 (O_41,N_22798,N_23333);
xor UO_42 (O_42,N_22976,N_24666);
nor UO_43 (O_43,N_22223,N_22643);
and UO_44 (O_44,N_24043,N_24372);
nor UO_45 (O_45,N_22569,N_24140);
or UO_46 (O_46,N_23163,N_24897);
or UO_47 (O_47,N_23415,N_22981);
and UO_48 (O_48,N_23133,N_24168);
xor UO_49 (O_49,N_24846,N_23312);
nor UO_50 (O_50,N_23399,N_23756);
or UO_51 (O_51,N_22204,N_22184);
and UO_52 (O_52,N_22552,N_22591);
nand UO_53 (O_53,N_23435,N_24544);
nand UO_54 (O_54,N_22753,N_22431);
nand UO_55 (O_55,N_23785,N_23254);
nand UO_56 (O_56,N_24407,N_22900);
and UO_57 (O_57,N_22192,N_24474);
or UO_58 (O_58,N_22787,N_23918);
xor UO_59 (O_59,N_24483,N_22326);
and UO_60 (O_60,N_24099,N_21950);
nor UO_61 (O_61,N_24702,N_24136);
and UO_62 (O_62,N_23390,N_24808);
or UO_63 (O_63,N_24624,N_21908);
or UO_64 (O_64,N_23974,N_23048);
nand UO_65 (O_65,N_24693,N_24183);
nor UO_66 (O_66,N_22053,N_24055);
xor UO_67 (O_67,N_22621,N_24764);
and UO_68 (O_68,N_21989,N_22066);
xor UO_69 (O_69,N_22110,N_24078);
or UO_70 (O_70,N_22662,N_22917);
nand UO_71 (O_71,N_23274,N_24881);
or UO_72 (O_72,N_21968,N_24780);
and UO_73 (O_73,N_24312,N_23492);
xor UO_74 (O_74,N_24371,N_24949);
nand UO_75 (O_75,N_23737,N_24001);
and UO_76 (O_76,N_24518,N_24021);
and UO_77 (O_77,N_24108,N_24600);
nor UO_78 (O_78,N_23451,N_23014);
nor UO_79 (O_79,N_23653,N_21960);
nand UO_80 (O_80,N_22183,N_22438);
nor UO_81 (O_81,N_22337,N_24633);
nor UO_82 (O_82,N_24012,N_24039);
or UO_83 (O_83,N_23332,N_22801);
xnor UO_84 (O_84,N_22967,N_23579);
and UO_85 (O_85,N_21914,N_22574);
nand UO_86 (O_86,N_22391,N_22076);
xnor UO_87 (O_87,N_22022,N_24064);
or UO_88 (O_88,N_21977,N_24022);
nor UO_89 (O_89,N_22694,N_22130);
nand UO_90 (O_90,N_22106,N_22898);
and UO_91 (O_91,N_22983,N_22522);
and UO_92 (O_92,N_21919,N_23498);
xnor UO_93 (O_93,N_22862,N_23947);
nor UO_94 (O_94,N_23531,N_22289);
nor UO_95 (O_95,N_23860,N_23700);
nor UO_96 (O_96,N_22924,N_24319);
xor UO_97 (O_97,N_22383,N_23468);
or UO_98 (O_98,N_24538,N_24998);
nor UO_99 (O_99,N_23681,N_23988);
and UO_100 (O_100,N_24013,N_23809);
nand UO_101 (O_101,N_23939,N_24036);
nand UO_102 (O_102,N_24029,N_23365);
xor UO_103 (O_103,N_24232,N_24382);
xor UO_104 (O_104,N_23857,N_22803);
or UO_105 (O_105,N_23488,N_22220);
and UO_106 (O_106,N_22839,N_22320);
or UO_107 (O_107,N_24848,N_24404);
nor UO_108 (O_108,N_22267,N_23814);
or UO_109 (O_109,N_24567,N_23367);
xor UO_110 (O_110,N_23346,N_23025);
nand UO_111 (O_111,N_23903,N_23280);
or UO_112 (O_112,N_23822,N_24931);
and UO_113 (O_113,N_23812,N_24575);
nand UO_114 (O_114,N_23398,N_23642);
and UO_115 (O_115,N_24880,N_23275);
xor UO_116 (O_116,N_24289,N_24855);
nor UO_117 (O_117,N_24913,N_24450);
nor UO_118 (O_118,N_24046,N_22208);
nor UO_119 (O_119,N_22042,N_24144);
nor UO_120 (O_120,N_24476,N_22825);
xor UO_121 (O_121,N_23339,N_23916);
and UO_122 (O_122,N_21965,N_22133);
or UO_123 (O_123,N_23364,N_21904);
nor UO_124 (O_124,N_22927,N_23200);
or UO_125 (O_125,N_24380,N_23058);
and UO_126 (O_126,N_23512,N_21881);
or UO_127 (O_127,N_24778,N_22470);
and UO_128 (O_128,N_24201,N_23998);
or UO_129 (O_129,N_24226,N_24215);
and UO_130 (O_130,N_22467,N_23331);
and UO_131 (O_131,N_22876,N_24228);
xor UO_132 (O_132,N_23808,N_22127);
or UO_133 (O_133,N_22612,N_24906);
xor UO_134 (O_134,N_23172,N_24956);
and UO_135 (O_135,N_22794,N_24646);
nor UO_136 (O_136,N_24616,N_23282);
nor UO_137 (O_137,N_23190,N_22889);
or UO_138 (O_138,N_24721,N_21903);
and UO_139 (O_139,N_23951,N_24333);
or UO_140 (O_140,N_22280,N_23348);
xor UO_141 (O_141,N_22985,N_22547);
xor UO_142 (O_142,N_22384,N_23949);
nand UO_143 (O_143,N_22125,N_23093);
xnor UO_144 (O_144,N_24851,N_24631);
nand UO_145 (O_145,N_24267,N_22865);
and UO_146 (O_146,N_22507,N_22962);
xnor UO_147 (O_147,N_23122,N_24082);
and UO_148 (O_148,N_23459,N_21887);
xnor UO_149 (O_149,N_22578,N_22519);
xnor UO_150 (O_150,N_22864,N_23185);
xnor UO_151 (O_151,N_23057,N_23237);
xnor UO_152 (O_152,N_23751,N_24914);
xnor UO_153 (O_153,N_21943,N_22230);
xor UO_154 (O_154,N_22997,N_22016);
and UO_155 (O_155,N_22888,N_23848);
and UO_156 (O_156,N_23626,N_22021);
or UO_157 (O_157,N_23002,N_22011);
nand UO_158 (O_158,N_24643,N_23052);
xor UO_159 (O_159,N_24759,N_23029);
nand UO_160 (O_160,N_23322,N_24153);
and UO_161 (O_161,N_24813,N_24845);
and UO_162 (O_162,N_22249,N_22398);
nor UO_163 (O_163,N_22647,N_23865);
nand UO_164 (O_164,N_24060,N_22421);
nand UO_165 (O_165,N_24155,N_24743);
or UO_166 (O_166,N_24423,N_24687);
nand UO_167 (O_167,N_23515,N_24004);
xor UO_168 (O_168,N_22189,N_22776);
xor UO_169 (O_169,N_23227,N_23729);
or UO_170 (O_170,N_23193,N_22290);
xor UO_171 (O_171,N_23382,N_24876);
and UO_172 (O_172,N_23880,N_22582);
nand UO_173 (O_173,N_22506,N_24963);
nand UO_174 (O_174,N_22113,N_24007);
xor UO_175 (O_175,N_22988,N_22868);
and UO_176 (O_176,N_23543,N_22543);
nand UO_177 (O_177,N_24104,N_23244);
nor UO_178 (O_178,N_23668,N_24254);
xor UO_179 (O_179,N_24385,N_23278);
or UO_180 (O_180,N_22681,N_23288);
nor UO_181 (O_181,N_23261,N_22599);
nor UO_182 (O_182,N_22564,N_23784);
or UO_183 (O_183,N_22327,N_24775);
nand UO_184 (O_184,N_23564,N_24577);
nor UO_185 (O_185,N_24773,N_24362);
and UO_186 (O_186,N_24718,N_23141);
or UO_187 (O_187,N_22394,N_22665);
nor UO_188 (O_188,N_23761,N_22529);
nand UO_189 (O_189,N_22119,N_22417);
or UO_190 (O_190,N_23044,N_24898);
and UO_191 (O_191,N_24047,N_22228);
or UO_192 (O_192,N_23197,N_22781);
xnor UO_193 (O_193,N_22994,N_24590);
nor UO_194 (O_194,N_24205,N_23300);
nand UO_195 (O_195,N_24954,N_24630);
and UO_196 (O_196,N_23082,N_22276);
xnor UO_197 (O_197,N_23968,N_22531);
or UO_198 (O_198,N_22309,N_22940);
nor UO_199 (O_199,N_24462,N_23240);
nor UO_200 (O_200,N_23591,N_24120);
nor UO_201 (O_201,N_24981,N_22572);
or UO_202 (O_202,N_24824,N_24310);
or UO_203 (O_203,N_24916,N_23999);
and UO_204 (O_204,N_24486,N_24042);
nand UO_205 (O_205,N_22872,N_22496);
nand UO_206 (O_206,N_24657,N_22233);
xor UO_207 (O_207,N_23752,N_22744);
and UO_208 (O_208,N_23107,N_23994);
nand UO_209 (O_209,N_22283,N_22424);
and UO_210 (O_210,N_24360,N_24996);
nand UO_211 (O_211,N_22114,N_23714);
or UO_212 (O_212,N_23375,N_23930);
and UO_213 (O_213,N_23369,N_22084);
nand UO_214 (O_214,N_23872,N_23730);
and UO_215 (O_215,N_23562,N_23595);
and UO_216 (O_216,N_23893,N_22587);
nand UO_217 (O_217,N_23632,N_23694);
or UO_218 (O_218,N_23264,N_22005);
or UO_219 (O_219,N_24519,N_24937);
or UO_220 (O_220,N_23495,N_23943);
xor UO_221 (O_221,N_23329,N_24134);
and UO_222 (O_222,N_24837,N_23189);
nand UO_223 (O_223,N_24110,N_23593);
or UO_224 (O_224,N_22343,N_24840);
or UO_225 (O_225,N_22474,N_23368);
nor UO_226 (O_226,N_23552,N_22369);
or UO_227 (O_227,N_24432,N_22949);
nor UO_228 (O_228,N_24599,N_23297);
nor UO_229 (O_229,N_24270,N_23783);
xnor UO_230 (O_230,N_22404,N_23613);
or UO_231 (O_231,N_23690,N_21953);
or UO_232 (O_232,N_24034,N_22622);
nand UO_233 (O_233,N_23328,N_24572);
nand UO_234 (O_234,N_24156,N_23313);
or UO_235 (O_235,N_22640,N_23478);
and UO_236 (O_236,N_24930,N_24634);
and UO_237 (O_237,N_24003,N_22762);
xor UO_238 (O_238,N_24160,N_23525);
or UO_239 (O_239,N_22484,N_22723);
xnor UO_240 (O_240,N_22627,N_22633);
nor UO_241 (O_241,N_24027,N_23376);
and UO_242 (O_242,N_24453,N_23750);
nand UO_243 (O_243,N_23127,N_22026);
and UO_244 (O_244,N_22333,N_22505);
nor UO_245 (O_245,N_24400,N_22715);
nand UO_246 (O_246,N_24279,N_24769);
and UO_247 (O_247,N_24944,N_24529);
and UO_248 (O_248,N_23753,N_24555);
xor UO_249 (O_249,N_23972,N_23769);
xor UO_250 (O_250,N_23699,N_23522);
nor UO_251 (O_251,N_22261,N_23231);
xnor UO_252 (O_252,N_22165,N_22416);
or UO_253 (O_253,N_24216,N_23105);
nand UO_254 (O_254,N_24604,N_24320);
and UO_255 (O_255,N_22434,N_22457);
nand UO_256 (O_256,N_23026,N_21878);
nor UO_257 (O_257,N_23780,N_23276);
xor UO_258 (O_258,N_23491,N_23534);
or UO_259 (O_259,N_24208,N_22169);
xnor UO_260 (O_260,N_22592,N_22501);
xor UO_261 (O_261,N_23220,N_23996);
or UO_262 (O_262,N_24669,N_24699);
nand UO_263 (O_263,N_21915,N_22686);
nor UO_264 (O_264,N_22006,N_24121);
nor UO_265 (O_265,N_24521,N_23663);
nor UO_266 (O_266,N_22335,N_22590);
nand UO_267 (O_267,N_23405,N_24838);
xnor UO_268 (O_268,N_24635,N_22048);
nand UO_269 (O_269,N_24191,N_24388);
and UO_270 (O_270,N_24127,N_23631);
or UO_271 (O_271,N_23315,N_23155);
and UO_272 (O_272,N_24223,N_24000);
xnor UO_273 (O_273,N_23889,N_24165);
and UO_274 (O_274,N_24069,N_22761);
or UO_275 (O_275,N_24999,N_23447);
nand UO_276 (O_276,N_23232,N_24879);
xnor UO_277 (O_277,N_23911,N_23176);
and UO_278 (O_278,N_22579,N_24660);
and UO_279 (O_279,N_22910,N_22254);
xor UO_280 (O_280,N_23841,N_23268);
nand UO_281 (O_281,N_22260,N_24324);
xnor UO_282 (O_282,N_22597,N_23651);
xor UO_283 (O_283,N_24866,N_22913);
or UO_284 (O_284,N_23024,N_22835);
nand UO_285 (O_285,N_24093,N_23854);
nand UO_286 (O_286,N_22773,N_24005);
nand UO_287 (O_287,N_22482,N_21993);
and UO_288 (O_288,N_24298,N_24977);
xnor UO_289 (O_289,N_22702,N_22933);
and UO_290 (O_290,N_24692,N_24656);
and UO_291 (O_291,N_24256,N_24435);
and UO_292 (O_292,N_24020,N_23378);
nor UO_293 (O_293,N_24974,N_22282);
nand UO_294 (O_294,N_22236,N_22925);
nor UO_295 (O_295,N_24429,N_24028);
nor UO_296 (O_296,N_23617,N_22705);
or UO_297 (O_297,N_22514,N_24861);
nor UO_298 (O_298,N_23047,N_24472);
nand UO_299 (O_299,N_22957,N_24091);
or UO_300 (O_300,N_23246,N_24713);
and UO_301 (O_301,N_23616,N_24826);
nor UO_302 (O_302,N_22142,N_23325);
or UO_303 (O_303,N_22441,N_22301);
or UO_304 (O_304,N_21951,N_22176);
or UO_305 (O_305,N_23799,N_23077);
nor UO_306 (O_306,N_24993,N_23828);
xnor UO_307 (O_307,N_23299,N_23990);
xor UO_308 (O_308,N_21980,N_22920);
nand UO_309 (O_309,N_23934,N_23766);
or UO_310 (O_310,N_24761,N_24961);
nor UO_311 (O_311,N_24264,N_22675);
or UO_312 (O_312,N_24141,N_24788);
nor UO_313 (O_313,N_22596,N_24524);
xnor UO_314 (O_314,N_24610,N_22747);
nand UO_315 (O_315,N_23762,N_23351);
xnor UO_316 (O_316,N_24950,N_23009);
nand UO_317 (O_317,N_22209,N_23412);
and UO_318 (O_318,N_22240,N_24077);
xnor UO_319 (O_319,N_24708,N_24283);
and UO_320 (O_320,N_22397,N_22348);
and UO_321 (O_321,N_24629,N_22754);
xor UO_322 (O_322,N_24909,N_24566);
nand UO_323 (O_323,N_22757,N_22748);
and UO_324 (O_324,N_22727,N_21937);
nor UO_325 (O_325,N_24300,N_24211);
xnor UO_326 (O_326,N_24089,N_22896);
xnor UO_327 (O_327,N_22834,N_22685);
xor UO_328 (O_328,N_24230,N_22832);
nand UO_329 (O_329,N_24337,N_22654);
nand UO_330 (O_330,N_22020,N_22674);
nand UO_331 (O_331,N_23864,N_22968);
xor UO_332 (O_332,N_24068,N_22526);
nor UO_333 (O_333,N_24128,N_24252);
and UO_334 (O_334,N_24419,N_24147);
xor UO_335 (O_335,N_23763,N_24361);
xor UO_336 (O_336,N_23843,N_24482);
xor UO_337 (O_337,N_22102,N_24691);
or UO_338 (O_338,N_22465,N_22846);
xor UO_339 (O_339,N_24864,N_22663);
xor UO_340 (O_340,N_22779,N_24569);
nand UO_341 (O_341,N_22078,N_24026);
and UO_342 (O_342,N_22577,N_22164);
or UO_343 (O_343,N_24053,N_23881);
xnor UO_344 (O_344,N_24819,N_22258);
nand UO_345 (O_345,N_23294,N_22163);
and UO_346 (O_346,N_23781,N_24679);
nor UO_347 (O_347,N_22677,N_23486);
or UO_348 (O_348,N_24238,N_22508);
or UO_349 (O_349,N_23735,N_23384);
or UO_350 (O_350,N_23188,N_22210);
nor UO_351 (O_351,N_22765,N_22936);
xor UO_352 (O_352,N_22718,N_23925);
or UO_353 (O_353,N_22027,N_22097);
or UO_354 (O_354,N_22373,N_23437);
xnor UO_355 (O_355,N_22775,N_24883);
and UO_356 (O_356,N_23053,N_22045);
or UO_357 (O_357,N_24222,N_22466);
nand UO_358 (O_358,N_23095,N_24146);
nor UO_359 (O_359,N_23475,N_22566);
nand UO_360 (O_360,N_23813,N_22444);
or UO_361 (O_361,N_22637,N_24303);
and UO_362 (O_362,N_23982,N_23732);
and UO_363 (O_363,N_24918,N_22907);
xnor UO_364 (O_364,N_22515,N_22653);
xor UO_365 (O_365,N_23606,N_24375);
nand UO_366 (O_366,N_23151,N_23938);
or UO_367 (O_367,N_24576,N_23380);
and UO_368 (O_368,N_23704,N_23560);
and UO_369 (O_369,N_23576,N_23902);
nor UO_370 (O_370,N_23920,N_24789);
nor UO_371 (O_371,N_23060,N_23234);
and UO_372 (O_372,N_23489,N_23508);
nand UO_373 (O_373,N_23302,N_22367);
nor UO_374 (O_374,N_22387,N_22960);
xor UO_375 (O_375,N_22472,N_22971);
or UO_376 (O_376,N_23271,N_24858);
nand UO_377 (O_377,N_24308,N_23655);
or UO_378 (O_378,N_24460,N_24085);
and UO_379 (O_379,N_23277,N_24101);
and UO_380 (O_380,N_23054,N_23403);
nor UO_381 (O_381,N_22171,N_22790);
xor UO_382 (O_382,N_23162,N_22729);
nand UO_383 (O_383,N_22201,N_22341);
and UO_384 (O_384,N_23010,N_22939);
and UO_385 (O_385,N_23801,N_23977);
or UO_386 (O_386,N_22334,N_24800);
or UO_387 (O_387,N_23180,N_24413);
and UO_388 (O_388,N_21906,N_23461);
and UO_389 (O_389,N_23957,N_22381);
nand UO_390 (O_390,N_24383,N_24499);
and UO_391 (O_391,N_23969,N_23381);
nor UO_392 (O_392,N_22418,N_24115);
nand UO_393 (O_393,N_22180,N_24843);
nor UO_394 (O_394,N_21905,N_23147);
or UO_395 (O_395,N_22372,N_23361);
nor UO_396 (O_396,N_24905,N_24889);
and UO_397 (O_397,N_22717,N_22279);
xnor UO_398 (O_398,N_22570,N_23472);
or UO_399 (O_399,N_23106,N_22512);
nand UO_400 (O_400,N_24366,N_23217);
xor UO_401 (O_401,N_22449,N_24626);
and UO_402 (O_402,N_22638,N_24979);
xor UO_403 (O_403,N_24116,N_23241);
xnor UO_404 (O_404,N_22439,N_22820);
nor UO_405 (O_405,N_24988,N_23612);
nand UO_406 (O_406,N_23929,N_24710);
xnor UO_407 (O_407,N_23572,N_24707);
xor UO_408 (O_408,N_24714,N_24059);
and UO_409 (O_409,N_22268,N_22523);
and UO_410 (O_410,N_22860,N_22237);
xor UO_411 (O_411,N_23948,N_24445);
xor UO_412 (O_412,N_24558,N_22074);
and UO_413 (O_413,N_23810,N_22610);
or UO_414 (O_414,N_22344,N_22168);
nand UO_415 (O_415,N_24340,N_23017);
or UO_416 (O_416,N_22366,N_22471);
or UO_417 (O_417,N_23109,N_22393);
xor UO_418 (O_418,N_23795,N_23896);
nand UO_419 (O_419,N_22105,N_23686);
nand UO_420 (O_420,N_23716,N_23794);
xor UO_421 (O_421,N_24126,N_23588);
xnor UO_422 (O_422,N_22710,N_23703);
xnor UO_423 (O_423,N_22986,N_23088);
nor UO_424 (O_424,N_24355,N_23236);
xor UO_425 (O_425,N_24545,N_23638);
and UO_426 (O_426,N_24345,N_22687);
and UO_427 (O_427,N_22154,N_24568);
and UO_428 (O_428,N_24595,N_21979);
nor UO_429 (O_429,N_22619,N_23520);
or UO_430 (O_430,N_24795,N_22539);
xnor UO_431 (O_431,N_23424,N_22764);
xnor UO_432 (O_432,N_24929,N_23118);
or UO_433 (O_433,N_24364,N_24900);
nor UO_434 (O_434,N_24682,N_22784);
nor UO_435 (O_435,N_22618,N_24010);
xnor UO_436 (O_436,N_23481,N_22585);
nor UO_437 (O_437,N_24446,N_24282);
nor UO_438 (O_438,N_23303,N_24427);
nor UO_439 (O_439,N_23111,N_22874);
xor UO_440 (O_440,N_22055,N_24016);
or UO_441 (O_441,N_23311,N_23772);
and UO_442 (O_442,N_22049,N_24615);
or UO_443 (O_443,N_24019,N_24031);
and UO_444 (O_444,N_24150,N_24741);
xor UO_445 (O_445,N_22842,N_24745);
and UO_446 (O_446,N_24739,N_23805);
nor UO_447 (O_447,N_24171,N_21884);
or UO_448 (O_448,N_23511,N_24389);
and UO_449 (O_449,N_24794,N_24451);
and UO_450 (O_450,N_22253,N_23353);
nor UO_451 (O_451,N_24071,N_23831);
or UO_452 (O_452,N_22533,N_24737);
xnor UO_453 (O_453,N_23316,N_22549);
xnor UO_454 (O_454,N_23228,N_22498);
and UO_455 (O_455,N_23542,N_23301);
nand UO_456 (O_456,N_23262,N_22486);
and UO_457 (O_457,N_24084,N_22175);
xnor UO_458 (O_458,N_22054,N_24640);
nand UO_459 (O_459,N_23207,N_24363);
and UO_460 (O_460,N_24970,N_23904);
nor UO_461 (O_461,N_22087,N_22931);
or UO_462 (O_462,N_24406,N_24170);
nand UO_463 (O_463,N_23862,N_23760);
nor UO_464 (O_464,N_24940,N_21910);
nand UO_465 (O_465,N_23961,N_22714);
and UO_466 (O_466,N_24671,N_23194);
xor UO_467 (O_467,N_21875,N_24111);
and UO_468 (O_468,N_23608,N_22789);
xor UO_469 (O_469,N_22942,N_22521);
nand UO_470 (O_470,N_24251,N_23091);
nor UO_471 (O_471,N_24987,N_23754);
nor UO_472 (O_472,N_24960,N_24703);
or UO_473 (O_473,N_24514,N_24976);
and UO_474 (O_474,N_23978,N_22490);
nand UO_475 (O_475,N_23659,N_22278);
xnor UO_476 (O_476,N_24917,N_21959);
xor UO_477 (O_477,N_22648,N_22356);
xnor UO_478 (O_478,N_24594,N_22060);
xnor UO_479 (O_479,N_24454,N_24964);
xnor UO_480 (O_480,N_23484,N_23391);
and UO_481 (O_481,N_24972,N_22758);
and UO_482 (O_482,N_24507,N_23414);
nor UO_483 (O_483,N_22453,N_24886);
and UO_484 (O_484,N_22721,N_24508);
and UO_485 (O_485,N_22436,N_22652);
or UO_486 (O_486,N_22146,N_23928);
nor UO_487 (O_487,N_22166,N_23360);
nand UO_488 (O_488,N_23379,N_23941);
and UO_489 (O_489,N_24755,N_21981);
xor UO_490 (O_490,N_22945,N_22520);
nand UO_491 (O_491,N_22600,N_23583);
nand UO_492 (O_492,N_24760,N_22826);
nor UO_493 (O_493,N_22015,N_24801);
or UO_494 (O_494,N_22118,N_22922);
xor UO_495 (O_495,N_24018,N_22903);
or UO_496 (O_496,N_24648,N_24169);
and UO_497 (O_497,N_24471,N_24618);
nand UO_498 (O_498,N_21916,N_23198);
xnor UO_499 (O_499,N_23099,N_23104);
nor UO_500 (O_500,N_22243,N_22304);
and UO_501 (O_501,N_23224,N_22688);
nor UO_502 (O_502,N_23210,N_24608);
nand UO_503 (O_503,N_24447,N_24044);
nand UO_504 (O_504,N_23950,N_23097);
xnor UO_505 (O_505,N_22285,N_22923);
nand UO_506 (O_506,N_23745,N_22838);
xnor UO_507 (O_507,N_24839,N_22990);
nor UO_508 (O_508,N_24652,N_22221);
or UO_509 (O_509,N_24871,N_24014);
or UO_510 (O_510,N_24066,N_24513);
and UO_511 (O_511,N_24247,N_22129);
or UO_512 (O_512,N_24732,N_24835);
xnor UO_513 (O_513,N_23506,N_22594);
and UO_514 (O_514,N_24784,N_24939);
or UO_515 (O_515,N_22937,N_22571);
nand UO_516 (O_516,N_23658,N_23952);
nand UO_517 (O_517,N_21985,N_22565);
or UO_518 (O_518,N_24154,N_24709);
xnor UO_519 (O_519,N_22788,N_22707);
and UO_520 (O_520,N_22312,N_24449);
nand UO_521 (O_521,N_23173,N_23290);
or UO_522 (O_522,N_22093,N_24325);
and UO_523 (O_523,N_23249,N_23233);
xor UO_524 (O_524,N_22395,N_21952);
nand UO_525 (O_525,N_23086,N_23102);
or UO_526 (O_526,N_23022,N_22270);
nor UO_527 (O_527,N_23863,N_24040);
and UO_528 (O_528,N_23117,N_23793);
nor UO_529 (O_529,N_23245,N_24402);
nor UO_530 (O_530,N_23533,N_22953);
nand UO_531 (O_531,N_24441,N_24517);
nor UO_532 (O_532,N_24935,N_23110);
or UO_533 (O_533,N_24017,N_23397);
xnor UO_534 (O_534,N_22476,N_24469);
or UO_535 (O_535,N_22461,N_24766);
xnor UO_536 (O_536,N_23087,N_23458);
and UO_537 (O_537,N_24309,N_23824);
nand UO_538 (O_538,N_24166,N_22242);
and UO_539 (O_539,N_24131,N_24338);
nand UO_540 (O_540,N_24680,N_24668);
xor UO_541 (O_541,N_24431,N_23976);
xnor UO_542 (O_542,N_23635,N_22310);
xnor UO_543 (O_543,N_22706,N_22080);
and UO_544 (O_544,N_23624,N_22305);
nand UO_545 (O_545,N_23089,N_22340);
or UO_546 (O_546,N_23387,N_23362);
xnor UO_547 (O_547,N_22683,N_24820);
and UO_548 (O_548,N_24772,N_23839);
or UO_549 (O_549,N_23697,N_24335);
or UO_550 (O_550,N_21944,N_22682);
nand UO_551 (O_551,N_23129,N_24161);
or UO_552 (O_552,N_22503,N_23283);
xnor UO_553 (O_553,N_24662,N_24505);
xor UO_554 (O_554,N_24504,N_22720);
xnor UO_555 (O_555,N_24727,N_23685);
nand UO_556 (O_556,N_22088,N_24313);
nand UO_557 (O_557,N_23423,N_22462);
and UO_558 (O_558,N_24611,N_24667);
and UO_559 (O_559,N_22793,N_23178);
xnor UO_560 (O_560,N_23112,N_22980);
or UO_561 (O_561,N_24908,N_24596);
nand UO_562 (O_562,N_24705,N_24684);
nor UO_563 (O_563,N_24736,N_24428);
xor UO_564 (O_564,N_22700,N_22414);
and UO_565 (O_565,N_24065,N_23570);
or UO_566 (O_566,N_24852,N_23433);
nand UO_567 (O_567,N_24198,N_22556);
and UO_568 (O_568,N_22778,N_24123);
and UO_569 (O_569,N_23923,N_22915);
nand UO_570 (O_570,N_24443,N_24578);
xnor UO_571 (O_571,N_24810,N_21954);
nor UO_572 (O_572,N_23568,N_21895);
nor UO_573 (O_573,N_23926,N_23208);
nor UO_574 (O_574,N_24809,N_21995);
or UO_575 (O_575,N_24465,N_22500);
xnor UO_576 (O_576,N_24132,N_22043);
nand UO_577 (O_577,N_24158,N_23269);
xnor UO_578 (O_578,N_23767,N_24526);
nand UO_579 (O_579,N_21928,N_24396);
nor UO_580 (O_580,N_24133,N_22298);
nand UO_581 (O_581,N_24951,N_24288);
xor UO_582 (O_582,N_24860,N_24369);
xor UO_583 (O_583,N_22092,N_24730);
nor UO_584 (O_584,N_23239,N_23046);
nand UO_585 (O_585,N_24081,N_23611);
nor UO_586 (O_586,N_23733,N_24329);
and UO_587 (O_587,N_22576,N_22403);
xor UO_588 (O_588,N_22932,N_23856);
nand UO_589 (O_589,N_23940,N_22064);
or UO_590 (O_590,N_22908,N_24791);
nand UO_591 (O_591,N_24367,N_23136);
xnor UO_592 (O_592,N_23586,N_24650);
nor UO_593 (O_593,N_23226,N_22003);
nor UO_594 (O_594,N_24532,N_22568);
and UO_595 (O_595,N_22513,N_24189);
nand UO_596 (O_596,N_23272,N_24415);
xor UO_597 (O_597,N_24096,N_22412);
nand UO_598 (O_598,N_23885,N_24376);
and UO_599 (O_599,N_23634,N_24782);
and UO_600 (O_600,N_24080,N_24214);
xor UO_601 (O_601,N_23242,N_24934);
and UO_602 (O_602,N_22691,N_22517);
nand UO_603 (O_603,N_24351,N_24927);
nand UO_604 (O_604,N_24754,N_23536);
and UO_605 (O_605,N_23630,N_23877);
or UO_606 (O_606,N_24480,N_22068);
xor UO_607 (O_607,N_23895,N_24162);
xor UO_608 (O_608,N_22382,N_24644);
nor UO_609 (O_609,N_22173,N_24893);
xnor UO_610 (O_610,N_23079,N_23620);
xor UO_611 (O_611,N_22774,N_24607);
or UO_612 (O_612,N_23598,N_24379);
nand UO_613 (O_613,N_24959,N_23201);
nand UO_614 (O_614,N_24688,N_23629);
or UO_615 (O_615,N_22284,N_22156);
nand UO_616 (O_616,N_24193,N_23050);
or UO_617 (O_617,N_23400,N_24103);
nand UO_618 (O_618,N_23186,N_22274);
nor UO_619 (O_619,N_23455,N_22331);
xnor UO_620 (O_620,N_22264,N_24548);
nand UO_621 (O_621,N_24067,N_24442);
or UO_622 (O_622,N_23284,N_21929);
xor UO_623 (O_623,N_23164,N_23321);
or UO_624 (O_624,N_22853,N_24048);
xnor UO_625 (O_625,N_21969,N_22121);
nor UO_626 (O_626,N_23971,N_23693);
or UO_627 (O_627,N_23582,N_24479);
and UO_628 (O_628,N_23566,N_24502);
xnor UO_629 (O_629,N_23460,N_23043);
or UO_630 (O_630,N_23654,N_24711);
nand UO_631 (O_631,N_22469,N_23623);
nand UO_632 (O_632,N_22160,N_22429);
or UO_633 (O_633,N_23680,N_24706);
and UO_634 (O_634,N_22639,N_22950);
nor UO_635 (O_635,N_22281,N_22996);
nor UO_636 (O_636,N_23251,N_24535);
and UO_637 (O_637,N_24129,N_23212);
and UO_638 (O_638,N_23355,N_22225);
nor UO_639 (O_639,N_23094,N_23778);
and UO_640 (O_640,N_23870,N_22593);
and UO_641 (O_641,N_24398,N_24817);
or UO_642 (O_642,N_24497,N_21898);
nand UO_643 (O_643,N_24796,N_22442);
or UO_644 (O_644,N_23526,N_23170);
or UO_645 (O_645,N_23773,N_23985);
or UO_646 (O_646,N_24639,N_23876);
xnor UO_647 (O_647,N_23135,N_23833);
xor UO_648 (O_648,N_23410,N_22786);
nand UO_649 (O_649,N_23519,N_22238);
xor UO_650 (O_650,N_24651,N_22277);
nand UO_651 (O_651,N_23633,N_24799);
nor UO_652 (O_652,N_24911,N_24051);
nor UO_653 (O_653,N_23074,N_24992);
xor UO_654 (O_654,N_24307,N_24536);
or UO_655 (O_655,N_23042,N_23408);
or UO_656 (O_656,N_23139,N_24062);
xor UO_657 (O_657,N_22328,N_22554);
xor UO_658 (O_658,N_22580,N_22679);
nor UO_659 (O_659,N_24627,N_24827);
nand UO_660 (O_660,N_22409,N_23023);
nor UO_661 (O_661,N_23051,N_24037);
or UO_662 (O_662,N_23959,N_24190);
or UO_663 (O_663,N_24887,N_24008);
nand UO_664 (O_664,N_24948,N_22629);
xnor UO_665 (O_665,N_22708,N_22458);
nor UO_666 (O_666,N_23479,N_23258);
nor UO_667 (O_667,N_22562,N_23907);
and UO_668 (O_668,N_24673,N_24694);
and UO_669 (O_669,N_23256,N_23080);
nand UO_670 (O_670,N_22992,N_23345);
and UO_671 (O_671,N_22430,N_24448);
xnor UO_672 (O_672,N_23748,N_22029);
and UO_673 (O_673,N_21924,N_23521);
or UO_674 (O_674,N_24530,N_23225);
nand UO_675 (O_675,N_22947,N_23741);
nor UO_676 (O_676,N_23973,N_24957);
or UO_677 (O_677,N_23363,N_24797);
nor UO_678 (O_678,N_23581,N_24206);
and UO_679 (O_679,N_23449,N_21889);
nand UO_680 (O_680,N_23518,N_23416);
and UO_681 (O_681,N_24343,N_24202);
nor UO_682 (O_682,N_24738,N_23956);
and UO_683 (O_683,N_22678,N_23395);
nand UO_684 (O_684,N_23558,N_24552);
or UO_685 (O_685,N_23609,N_23850);
xor UO_686 (O_686,N_23970,N_22135);
and UO_687 (O_687,N_23336,N_24882);
nor UO_688 (O_688,N_23837,N_21909);
or UO_689 (O_689,N_22560,N_23868);
nor UO_690 (O_690,N_23177,N_24924);
or UO_691 (O_691,N_24075,N_23771);
xnor UO_692 (O_692,N_23335,N_22432);
and UO_693 (O_693,N_21992,N_23168);
or UO_694 (O_694,N_23742,N_22091);
nor UO_695 (O_695,N_22695,N_22368);
nand UO_696 (O_696,N_22445,N_23547);
xor UO_697 (O_697,N_22364,N_23955);
xnor UO_698 (O_698,N_22071,N_23927);
and UO_699 (O_699,N_24112,N_24853);
and UO_700 (O_700,N_24174,N_23308);
xor UO_701 (O_701,N_24421,N_22407);
and UO_702 (O_702,N_23892,N_23419);
nor UO_703 (O_703,N_23064,N_24591);
and UO_704 (O_704,N_22711,N_23296);
xor UO_705 (O_705,N_22040,N_24776);
and UO_706 (O_706,N_24676,N_21935);
xnor UO_707 (O_707,N_22998,N_24833);
nand UO_708 (O_708,N_24765,N_22132);
nand UO_709 (O_709,N_22177,N_24100);
nor UO_710 (O_710,N_22357,N_24936);
or UO_711 (O_711,N_22495,N_23432);
and UO_712 (O_712,N_24978,N_22959);
or UO_713 (O_713,N_21893,N_23802);
xor UO_714 (O_714,N_23701,N_22329);
xor UO_715 (O_715,N_22336,N_23065);
and UO_716 (O_716,N_22489,N_22023);
nand UO_717 (O_717,N_23140,N_23255);
nor UO_718 (O_718,N_23448,N_24125);
and UO_719 (O_719,N_21940,N_23342);
and UO_720 (O_720,N_22524,N_24305);
and UO_721 (O_721,N_22036,N_22935);
or UO_722 (O_722,N_24563,N_22159);
nor UO_723 (O_723,N_22363,N_23888);
nor UO_724 (O_724,N_21907,N_23314);
or UO_725 (O_725,N_22207,N_22451);
and UO_726 (O_726,N_24515,N_22806);
xnor UO_727 (O_727,N_23470,N_22532);
xnor UO_728 (O_728,N_23673,N_24947);
nand UO_729 (O_729,N_23143,N_21958);
nor UO_730 (O_730,N_24461,N_23639);
xnor UO_731 (O_731,N_22887,N_23537);
xnor UO_732 (O_732,N_23252,N_22628);
or UO_733 (O_733,N_23317,N_23827);
nor UO_734 (O_734,N_22311,N_22018);
xnor UO_735 (O_735,N_24770,N_22000);
or UO_736 (O_736,N_22315,N_22607);
or UO_737 (O_737,N_22620,N_22645);
xnor UO_738 (O_738,N_23607,N_22245);
nor UO_739 (O_739,N_22699,N_23774);
nor UO_740 (O_740,N_24495,N_22559);
nor UO_741 (O_741,N_23965,N_22401);
or UO_742 (O_742,N_23401,N_22191);
or UO_743 (O_743,N_24557,N_24695);
and UO_744 (O_744,N_22415,N_22089);
nand UO_745 (O_745,N_24965,N_23096);
and UO_746 (O_746,N_22725,N_23157);
and UO_747 (O_747,N_23338,N_23440);
or UO_748 (O_748,N_22332,N_22325);
xnor UO_749 (O_749,N_24922,N_22440);
nand UO_750 (O_750,N_23986,N_22056);
and UO_751 (O_751,N_23869,N_24525);
nand UO_752 (O_752,N_21966,N_22007);
and UO_753 (O_753,N_22886,N_21956);
nand UO_754 (O_754,N_22051,N_24868);
nand UO_755 (O_755,N_22205,N_24186);
or UO_756 (O_756,N_23571,N_24393);
nor UO_757 (O_757,N_22731,N_23149);
nor UO_758 (O_758,N_23849,N_23235);
xor UO_759 (O_759,N_23175,N_22229);
nand UO_760 (O_760,N_24145,N_22073);
and UO_761 (O_761,N_24523,N_23603);
nor UO_762 (O_762,N_22252,N_22661);
xnor UO_763 (O_763,N_21933,N_23580);
nor UO_764 (O_764,N_24637,N_24152);
or UO_765 (O_765,N_23817,N_23788);
or UO_766 (O_766,N_24330,N_24352);
and UO_767 (O_767,N_24370,N_24818);
and UO_768 (O_768,N_23469,N_22463);
and UO_769 (O_769,N_23477,N_23466);
nand UO_770 (O_770,N_24587,N_23497);
nand UO_771 (O_771,N_23597,N_23016);
and UO_772 (O_772,N_24588,N_24804);
or UO_773 (O_773,N_24658,N_24856);
nor UO_774 (O_774,N_22603,N_24806);
and UO_775 (O_775,N_23354,N_23130);
xnor UO_776 (O_776,N_23281,N_23483);
or UO_777 (O_777,N_22977,N_22247);
nand UO_778 (O_778,N_23698,N_22669);
or UO_779 (O_779,N_24049,N_22286);
xor UO_780 (O_780,N_23306,N_22792);
nand UO_781 (O_781,N_23962,N_23004);
xnor UO_782 (O_782,N_24516,N_24244);
xor UO_783 (O_783,N_23055,N_22635);
nand UO_784 (O_784,N_24280,N_22079);
or UO_785 (O_785,N_23436,N_23637);
nand UO_786 (O_786,N_24953,N_22650);
xor UO_787 (O_787,N_23446,N_22812);
nor UO_788 (O_788,N_22181,N_23126);
or UO_789 (O_789,N_23487,N_22152);
or UO_790 (O_790,N_24933,N_22246);
or UO_791 (O_791,N_23890,N_23775);
nand UO_792 (O_792,N_22871,N_23905);
and UO_793 (O_793,N_23666,N_22730);
nand UO_794 (O_794,N_23967,N_24278);
or UO_795 (O_795,N_24980,N_22186);
nor UO_796 (O_796,N_23445,N_22606);
xnor UO_797 (O_797,N_24910,N_22144);
nor UO_798 (O_798,N_24438,N_22613);
or UO_799 (O_799,N_23720,N_22030);
or UO_800 (O_800,N_23549,N_22819);
nor UO_801 (O_801,N_24197,N_21912);
and UO_802 (O_802,N_23621,N_22318);
xor UO_803 (O_803,N_23187,N_22224);
xor UO_804 (O_804,N_24455,N_22300);
xnor UO_805 (O_805,N_22104,N_23656);
and UO_806 (O_806,N_23819,N_21883);
nor UO_807 (O_807,N_22234,N_22492);
xnor UO_808 (O_808,N_22269,N_23167);
nor UO_809 (O_809,N_23429,N_23021);
or UO_810 (O_810,N_24274,N_23692);
xor UO_811 (O_811,N_24386,N_23740);
nor UO_812 (O_812,N_22275,N_22353);
or UO_813 (O_813,N_24757,N_24038);
nor UO_814 (O_814,N_24522,N_24353);
xnor UO_815 (O_815,N_22841,N_22019);
or UO_816 (O_816,N_23535,N_23786);
xnor UO_817 (O_817,N_24716,N_22103);
nor UO_818 (O_818,N_23627,N_22170);
and UO_819 (O_819,N_22881,N_22598);
nor UO_820 (O_820,N_21891,N_22973);
and UO_821 (O_821,N_22724,N_22235);
or UO_822 (O_822,N_23909,N_24832);
nand UO_823 (O_823,N_24619,N_24593);
nand UO_824 (O_824,N_23005,N_22390);
and UO_825 (O_825,N_22836,N_22099);
nor UO_826 (O_826,N_22061,N_22032);
nand UO_827 (O_827,N_22009,N_22692);
or UO_828 (O_828,N_23257,N_22821);
xnor UO_829 (O_829,N_22767,N_23744);
or UO_830 (O_830,N_23359,N_24726);
xor UO_831 (O_831,N_23502,N_21990);
and UO_832 (O_832,N_24291,N_24296);
nor UO_833 (O_833,N_22709,N_22338);
nor UO_834 (O_834,N_24812,N_22689);
or UO_835 (O_835,N_22869,N_23218);
xor UO_836 (O_836,N_24734,N_24157);
and UO_837 (O_837,N_22307,N_24973);
xor UO_838 (O_838,N_23768,N_22358);
nand UO_839 (O_839,N_22319,N_24625);
nand UO_840 (O_840,N_24117,N_22676);
and UO_841 (O_841,N_23589,N_24907);
xor UO_842 (O_842,N_24381,N_23823);
nand UO_843 (O_843,N_23900,N_24943);
and UO_844 (O_844,N_22899,N_22611);
nand UO_845 (O_845,N_22856,N_23660);
xnor UO_846 (O_846,N_23601,N_24204);
xnor UO_847 (O_847,N_23203,N_24561);
xor UO_848 (O_848,N_23736,N_23090);
nand UO_849 (O_849,N_22605,N_21885);
nor UO_850 (O_850,N_24925,N_24350);
nand UO_851 (O_851,N_21894,N_21930);
and UO_852 (O_852,N_24277,N_22581);
or UO_853 (O_853,N_22615,N_22342);
or UO_854 (O_854,N_24746,N_22807);
xor UO_855 (O_855,N_23337,N_23238);
xnor UO_856 (O_856,N_23266,N_23471);
and UO_857 (O_857,N_22355,N_22227);
nand UO_858 (O_858,N_22601,N_24696);
xor UO_859 (O_859,N_22380,N_22805);
nor UO_860 (O_860,N_23538,N_23015);
xnor UO_861 (O_861,N_24243,N_23723);
nor UO_862 (O_862,N_24336,N_24468);
or UO_863 (O_863,N_23983,N_23946);
and UO_864 (O_864,N_22904,N_23293);
or UO_865 (O_865,N_24295,N_23584);
nand UO_866 (O_866,N_24901,N_23992);
nor UO_867 (O_867,N_23707,N_21971);
nor UO_868 (O_868,N_23545,N_24181);
or UO_869 (O_869,N_22017,N_22737);
nor UO_870 (O_870,N_24581,N_23829);
or UO_871 (O_871,N_24717,N_23935);
or UO_872 (O_872,N_24475,N_24276);
and UO_873 (O_873,N_23702,N_24751);
or UO_874 (O_874,N_22855,N_22575);
nand UO_875 (O_875,N_22759,N_23350);
nor UO_876 (O_876,N_22148,N_22742);
and UO_877 (O_877,N_24811,N_22345);
xor UO_878 (O_878,N_21994,N_24164);
or UO_879 (O_879,N_24467,N_24967);
and UO_880 (O_880,N_24417,N_23886);
xor UO_881 (O_881,N_22052,N_22115);
xnor UO_882 (O_882,N_23585,N_24377);
nor UO_883 (O_883,N_23267,N_23825);
or UO_884 (O_884,N_23709,N_24786);
or UO_885 (O_885,N_24237,N_23711);
nand UO_886 (O_886,N_22473,N_24173);
xnor UO_887 (O_887,N_22815,N_22634);
and UO_888 (O_888,N_22623,N_22058);
and UO_889 (O_889,N_22217,N_22646);
nor UO_890 (O_890,N_24715,N_22475);
xor UO_891 (O_891,N_22840,N_23347);
or UO_892 (O_892,N_24478,N_24492);
xnor UO_893 (O_893,N_24559,N_23791);
xor UO_894 (O_894,N_23643,N_23517);
nand UO_895 (O_895,N_23758,N_23573);
xnor UO_896 (O_896,N_24863,N_24114);
nor UO_897 (O_897,N_23457,N_23103);
or UO_898 (O_898,N_22548,N_24872);
nor UO_899 (O_899,N_22001,N_24087);
or UO_900 (O_900,N_23156,N_23085);
or UO_901 (O_901,N_23855,N_23779);
nand UO_902 (O_902,N_22843,N_22493);
nand UO_903 (O_903,N_24520,N_22460);
nand UO_904 (O_904,N_23020,N_22542);
nand UO_905 (O_905,N_22555,N_22481);
or UO_906 (O_906,N_24902,N_24253);
xnor UO_907 (O_907,N_22783,N_24236);
nor UO_908 (O_908,N_24946,N_22944);
xnor UO_909 (O_909,N_22894,N_22203);
or UO_910 (O_910,N_21913,N_24542);
or UO_911 (O_911,N_23715,N_22795);
nand UO_912 (O_912,N_22785,N_23073);
xor UO_913 (O_913,N_22583,N_21876);
xor UO_914 (O_914,N_21963,N_24490);
nand UO_915 (O_915,N_23452,N_23327);
xor UO_916 (O_916,N_23901,N_22374);
xor UO_917 (O_917,N_23356,N_22822);
xnor UO_918 (O_918,N_23555,N_24422);
nand UO_919 (O_919,N_21970,N_22350);
xnor UO_920 (O_920,N_24314,N_22339);
xor UO_921 (O_921,N_24240,N_22346);
and UO_922 (O_922,N_23679,N_24698);
and UO_923 (O_923,N_22046,N_23161);
nand UO_924 (O_924,N_22906,N_24425);
xnor UO_925 (O_925,N_22510,N_23386);
xor UO_926 (O_926,N_23500,N_22244);
nor UO_927 (O_927,N_24073,N_24903);
nor UO_928 (O_928,N_21886,N_23875);
and UO_929 (O_929,N_22361,N_22317);
and UO_930 (O_930,N_23119,N_24259);
and UO_931 (O_931,N_22755,N_23640);
nand UO_932 (O_932,N_22984,N_23039);
xnor UO_933 (O_933,N_23984,N_23567);
nor UO_934 (O_934,N_23385,N_24623);
and UO_935 (O_935,N_24430,N_24700);
and UO_936 (O_936,N_21973,N_22082);
and UO_937 (O_937,N_24592,N_22561);
nor UO_938 (O_938,N_22138,N_24653);
nor UO_939 (O_939,N_23078,N_22010);
xnor UO_940 (O_940,N_23038,N_23040);
and UO_941 (O_941,N_23858,N_21946);
xor UO_942 (O_942,N_24685,N_24321);
xor UO_943 (O_943,N_22226,N_23899);
and UO_944 (O_944,N_23202,N_23465);
or UO_945 (O_945,N_23032,N_23532);
and UO_946 (O_946,N_22713,N_23615);
and UO_947 (O_947,N_24647,N_24304);
xor UO_948 (O_948,N_23796,N_22239);
xnor UO_949 (O_949,N_24945,N_23878);
nand UO_950 (O_950,N_22454,N_24602);
nor UO_951 (O_951,N_22641,N_22625);
and UO_952 (O_952,N_24024,N_24399);
nor UO_953 (O_953,N_22085,N_22297);
and UO_954 (O_954,N_23574,N_23019);
and UO_955 (O_955,N_24052,N_21931);
or UO_956 (O_956,N_23285,N_23407);
or UO_957 (O_957,N_23196,N_22112);
nor UO_958 (O_958,N_24547,N_23259);
xor UO_959 (O_959,N_24785,N_24076);
and UO_960 (O_960,N_23719,N_23556);
and UO_961 (O_961,N_22405,N_22139);
nor UO_962 (O_962,N_24009,N_24601);
and UO_963 (O_963,N_23910,N_22892);
and UO_964 (O_964,N_23182,N_22200);
nand UO_965 (O_965,N_23012,N_22965);
or UO_966 (O_966,N_23430,N_24850);
or UO_967 (O_967,N_24712,N_23821);
or UO_968 (O_968,N_22716,N_22604);
nand UO_969 (O_969,N_23657,N_23373);
and UO_970 (O_970,N_24346,N_23334);
or UO_971 (O_971,N_21923,N_23966);
and UO_972 (O_972,N_21900,N_22188);
nor UO_973 (O_973,N_23551,N_21926);
nor UO_974 (O_974,N_22746,N_23524);
nand UO_975 (O_975,N_24932,N_23667);
or UO_976 (O_976,N_23153,N_23388);
nor UO_977 (O_977,N_22557,N_24210);
nand UO_978 (O_978,N_23816,N_24844);
and UO_979 (O_979,N_22033,N_23076);
and UO_980 (O_980,N_22693,N_23221);
xnor UO_981 (O_981,N_23247,N_22386);
nor UO_982 (O_982,N_23438,N_22970);
or UO_983 (O_983,N_23765,N_23614);
nand UO_984 (O_984,N_22145,N_24494);
nor UO_985 (O_985,N_23826,N_24724);
or UO_986 (O_986,N_22982,N_24119);
and UO_987 (O_987,N_24828,N_22854);
nor UO_988 (O_988,N_23485,N_22617);
nand UO_989 (O_989,N_22198,N_23250);
nor UO_990 (O_990,N_24318,N_23738);
nand UO_991 (O_991,N_22231,N_22763);
or UO_992 (O_992,N_24287,N_23454);
xnor UO_993 (O_993,N_24203,N_22291);
nand UO_994 (O_994,N_23645,N_23453);
or UO_995 (O_995,N_22614,N_23842);
nand UO_996 (O_996,N_21976,N_22150);
and UO_997 (O_997,N_24598,N_22796);
xor UO_998 (O_998,N_24227,N_23602);
or UO_999 (O_999,N_23041,N_22349);
xnor UO_1000 (O_1000,N_22667,N_23499);
nor UO_1001 (O_1001,N_22893,N_23008);
nor UO_1002 (O_1002,N_23169,N_24834);
or UO_1003 (O_1003,N_23473,N_24139);
nand UO_1004 (O_1004,N_24242,N_24670);
or UO_1005 (O_1005,N_23422,N_24148);
nor UO_1006 (O_1006,N_23191,N_22550);
nand UO_1007 (O_1007,N_24528,N_23979);
nor UO_1008 (O_1008,N_22497,N_24403);
nand UO_1009 (O_1009,N_22155,N_21892);
and UO_1010 (O_1010,N_24719,N_22499);
or UO_1011 (O_1011,N_24793,N_21901);
nor UO_1012 (O_1012,N_22584,N_24185);
xnor UO_1013 (O_1013,N_24539,N_23505);
and UO_1014 (O_1014,N_22882,N_24294);
nor UO_1015 (O_1015,N_24570,N_24672);
and UO_1016 (O_1016,N_21927,N_23664);
and UO_1017 (O_1017,N_23027,N_22324);
xnor UO_1018 (O_1018,N_22751,N_24968);
or UO_1019 (O_1019,N_22069,N_24070);
or UO_1020 (O_1020,N_22660,N_23439);
nor UO_1021 (O_1021,N_24356,N_23160);
nand UO_1022 (O_1022,N_24466,N_23037);
or UO_1023 (O_1023,N_22428,N_22802);
xnor UO_1024 (O_1024,N_22732,N_22420);
and UO_1025 (O_1025,N_22288,N_23944);
nand UO_1026 (O_1026,N_23987,N_22530);
xor UO_1027 (O_1027,N_22378,N_22359);
and UO_1028 (O_1028,N_23305,N_24899);
and UO_1029 (O_1029,N_24219,N_22848);
and UO_1030 (O_1030,N_24255,N_21972);
or UO_1031 (O_1031,N_24884,N_22673);
or UO_1032 (O_1032,N_24098,N_23393);
xnor UO_1033 (O_1033,N_24192,N_22636);
nand UO_1034 (O_1034,N_24873,N_23371);
nor UO_1035 (O_1035,N_24293,N_23442);
and UO_1036 (O_1036,N_23152,N_23853);
nand UO_1037 (O_1037,N_22743,N_23590);
nand UO_1038 (O_1038,N_23942,N_24678);
nor UO_1039 (O_1039,N_23206,N_21991);
or UO_1040 (O_1040,N_23209,N_24235);
nor UO_1041 (O_1041,N_24540,N_24962);
xnor UO_1042 (O_1042,N_24892,N_24744);
nand UO_1043 (O_1043,N_22151,N_23144);
or UO_1044 (O_1044,N_23137,N_22814);
nor UO_1045 (O_1045,N_23084,N_22863);
nor UO_1046 (O_1046,N_21880,N_23883);
and UO_1047 (O_1047,N_24790,N_22178);
nor UO_1048 (O_1048,N_24187,N_24920);
or UO_1049 (O_1049,N_22385,N_22248);
nand UO_1050 (O_1050,N_22259,N_22979);
xor UO_1051 (O_1051,N_22697,N_22722);
xor UO_1052 (O_1052,N_22870,N_24649);
and UO_1053 (O_1053,N_22070,N_24955);
nand UO_1054 (O_1054,N_24213,N_22528);
nor UO_1055 (O_1055,N_24481,N_22399);
or UO_1056 (O_1056,N_22511,N_24311);
nand UO_1057 (O_1057,N_22504,N_22294);
nand UO_1058 (O_1058,N_22895,N_23600);
nand UO_1059 (O_1059,N_23035,N_22766);
nor UO_1060 (O_1060,N_22659,N_24458);
nor UO_1061 (O_1061,N_22126,N_23389);
nor UO_1062 (O_1062,N_23464,N_23818);
nand UO_1063 (O_1063,N_24982,N_24763);
or UO_1064 (O_1064,N_23995,N_23650);
nand UO_1065 (O_1065,N_24609,N_24632);
nor UO_1066 (O_1066,N_23417,N_23229);
or UO_1067 (O_1067,N_24261,N_21978);
nor UO_1068 (O_1068,N_24035,N_22518);
xor UO_1069 (O_1069,N_24841,N_22455);
nor UO_1070 (O_1070,N_24919,N_22866);
nand UO_1071 (O_1071,N_23428,N_22194);
nor UO_1072 (O_1072,N_22921,N_24874);
xor UO_1073 (O_1073,N_23960,N_24975);
nor UO_1074 (O_1074,N_22197,N_24105);
xnor UO_1075 (O_1075,N_22419,N_21925);
or UO_1076 (O_1076,N_23443,N_22120);
nor UO_1077 (O_1077,N_24368,N_23691);
nor UO_1078 (O_1078,N_23425,N_23150);
or UO_1079 (O_1079,N_22738,N_22232);
nand UO_1080 (O_1080,N_22447,N_23674);
and UO_1081 (O_1081,N_23559,N_22772);
xor UO_1082 (O_1082,N_22479,N_22991);
or UO_1083 (O_1083,N_23804,N_24411);
nor UO_1084 (O_1084,N_23739,N_23604);
nand UO_1085 (O_1085,N_22902,N_22589);
nand UO_1086 (O_1086,N_22563,N_24271);
nor UO_1087 (O_1087,N_22065,N_22299);
nand UO_1088 (O_1088,N_24175,N_22062);
and UO_1089 (O_1089,N_23671,N_23592);
or UO_1090 (O_1090,N_24359,N_22941);
xor UO_1091 (O_1091,N_24527,N_23253);
nor UO_1092 (O_1092,N_24986,N_23649);
xnor UO_1093 (O_1093,N_21975,N_23033);
or UO_1094 (O_1094,N_22413,N_23213);
nand UO_1095 (O_1095,N_22370,N_23007);
nor UO_1096 (O_1096,N_23648,N_24985);
nand UO_1097 (O_1097,N_23179,N_23510);
or UO_1098 (O_1098,N_23309,N_22934);
nand UO_1099 (O_1099,N_23490,N_24501);
nor UO_1100 (O_1100,N_22141,N_22847);
nand UO_1101 (O_1101,N_23421,N_23131);
xnor UO_1102 (O_1102,N_22698,N_22655);
or UO_1103 (O_1103,N_24921,N_23830);
or UO_1104 (O_1104,N_23056,N_22885);
nor UO_1105 (O_1105,N_22187,N_23450);
nor UO_1106 (O_1106,N_22153,N_23230);
nand UO_1107 (O_1107,N_24493,N_23887);
nor UO_1108 (O_1108,N_24701,N_23145);
and UO_1109 (O_1109,N_22993,N_24323);
xor UO_1110 (O_1110,N_24867,N_22859);
or UO_1111 (O_1111,N_22219,N_24774);
or UO_1112 (O_1112,N_24416,N_22410);
or UO_1113 (O_1113,N_24257,N_23647);
or UO_1114 (O_1114,N_23128,N_24740);
nand UO_1115 (O_1115,N_24109,N_24286);
or UO_1116 (O_1116,N_23787,N_23071);
xnor UO_1117 (O_1117,N_24072,N_22534);
xor UO_1118 (O_1118,N_22002,N_22624);
nor UO_1119 (O_1119,N_22035,N_23181);
nand UO_1120 (O_1120,N_24802,N_24904);
or UO_1121 (O_1121,N_24895,N_24424);
nor UO_1122 (O_1122,N_23341,N_24348);
or UO_1123 (O_1123,N_24941,N_22262);
or UO_1124 (O_1124,N_24102,N_23575);
nor UO_1125 (O_1125,N_24258,N_24281);
or UO_1126 (O_1126,N_23507,N_22588);
and UO_1127 (O_1127,N_23873,N_23563);
or UO_1128 (O_1128,N_23142,N_23344);
and UO_1129 (O_1129,N_24130,N_24779);
and UO_1130 (O_1130,N_24327,N_22914);
or UO_1131 (O_1131,N_22077,N_24260);
or UO_1132 (O_1132,N_23662,N_24767);
or UO_1133 (O_1133,N_22031,N_22124);
nand UO_1134 (O_1134,N_24661,N_21920);
or UO_1135 (O_1135,N_24033,N_23898);
or UO_1136 (O_1136,N_24750,N_22389);
xor UO_1137 (O_1137,N_24556,N_24354);
and UO_1138 (O_1138,N_23061,N_22321);
nor UO_1139 (O_1139,N_22213,N_23777);
xnor UO_1140 (O_1140,N_23578,N_23108);
nor UO_1141 (O_1141,N_23501,N_24580);
nand UO_1142 (O_1142,N_22586,N_23993);
and UO_1143 (O_1143,N_24199,N_23463);
and UO_1144 (O_1144,N_24030,N_22371);
xor UO_1145 (O_1145,N_23712,N_24332);
nor UO_1146 (O_1146,N_23045,N_24815);
nor UO_1147 (O_1147,N_23836,N_23183);
nor UO_1148 (O_1148,N_24805,N_22488);
xor UO_1149 (O_1149,N_22083,N_22075);
or UO_1150 (O_1150,N_24349,N_23811);
nor UO_1151 (O_1151,N_24731,N_23370);
and UO_1152 (O_1152,N_23358,N_24890);
and UO_1153 (O_1153,N_23476,N_23480);
nor UO_1154 (O_1154,N_24728,N_23688);
xnor UO_1155 (O_1155,N_24584,N_24742);
xor UO_1156 (O_1156,N_21998,N_24488);
nor UO_1157 (O_1157,N_23963,N_22427);
nand UO_1158 (O_1158,N_24830,N_23937);
nand UO_1159 (O_1159,N_23326,N_23840);
xnor UO_1160 (O_1160,N_22541,N_23289);
nand UO_1161 (O_1161,N_23063,N_24409);
and UO_1162 (O_1162,N_23803,N_22174);
and UO_1163 (O_1163,N_24420,N_22964);
xnor UO_1164 (O_1164,N_24533,N_24220);
nor UO_1165 (O_1165,N_22012,N_22884);
or UO_1166 (O_1166,N_23912,N_22182);
or UO_1167 (O_1167,N_24317,N_23396);
or UO_1168 (O_1168,N_22459,N_23062);
nand UO_1169 (O_1169,N_21932,N_24912);
nor UO_1170 (O_1170,N_23724,N_24582);
nand UO_1171 (O_1171,N_24729,N_23764);
and UO_1172 (O_1172,N_22014,N_24869);
nor UO_1173 (O_1173,N_22948,N_21902);
nor UO_1174 (O_1174,N_22909,N_22485);
or UO_1175 (O_1175,N_24531,N_24341);
nand UO_1176 (O_1176,N_23684,N_24135);
nor UO_1177 (O_1177,N_22873,N_22354);
xor UO_1178 (O_1178,N_23184,N_22969);
nand UO_1179 (O_1179,N_21999,N_24233);
or UO_1180 (O_1180,N_24241,N_24050);
xor UO_1181 (O_1181,N_23372,N_24179);
or UO_1182 (O_1182,N_24512,N_22241);
or UO_1183 (O_1183,N_23101,N_23031);
nand UO_1184 (O_1184,N_22108,N_22041);
nand UO_1185 (O_1185,N_24248,N_23081);
or UO_1186 (O_1186,N_23731,N_23307);
xor UO_1187 (O_1187,N_24268,N_22850);
nand UO_1188 (O_1188,N_22494,N_23318);
or UO_1189 (O_1189,N_23075,N_23546);
nor UO_1190 (O_1190,N_24079,N_23550);
and UO_1191 (O_1191,N_23847,N_23444);
xor UO_1192 (O_1192,N_24063,N_23705);
xor UO_1193 (O_1193,N_24733,N_22149);
and UO_1194 (O_1194,N_24926,N_24122);
and UO_1195 (O_1195,N_24749,N_22901);
and UO_1196 (O_1196,N_22266,N_23527);
or UO_1197 (O_1197,N_22483,N_23509);
and UO_1198 (O_1198,N_24506,N_24436);
nor UO_1199 (O_1199,N_22406,N_22837);
and UO_1200 (O_1200,N_21922,N_21987);
nor UO_1201 (O_1201,N_24229,N_24118);
nand UO_1202 (O_1202,N_22351,N_24328);
and UO_1203 (O_1203,N_22123,N_23646);
or UO_1204 (O_1204,N_23513,N_23504);
and UO_1205 (O_1205,N_23981,N_24231);
and UO_1206 (O_1206,N_21938,N_23219);
nand UO_1207 (O_1207,N_24358,N_24885);
or UO_1208 (O_1208,N_24636,N_24825);
nand UO_1209 (O_1209,N_24177,N_23265);
and UO_1210 (O_1210,N_23072,N_22047);
nand UO_1211 (O_1211,N_23214,N_23964);
and UO_1212 (O_1212,N_24470,N_23815);
or UO_1213 (O_1213,N_23529,N_24645);
nor UO_1214 (O_1214,N_22330,N_24822);
or UO_1215 (O_1215,N_24217,N_24995);
and UO_1216 (O_1216,N_21945,N_22396);
xnor UO_1217 (O_1217,N_23800,N_22741);
nand UO_1218 (O_1218,N_24803,N_22448);
nand UO_1219 (O_1219,N_24056,N_24045);
xnor UO_1220 (O_1220,N_22912,N_22891);
nand UO_1221 (O_1221,N_24783,N_24015);
xor UO_1222 (O_1222,N_22987,N_21984);
nand UO_1223 (O_1223,N_23782,N_24554);
xor UO_1224 (O_1224,N_24989,N_22292);
nor UO_1225 (O_1225,N_23770,N_24275);
xnor UO_1226 (O_1226,N_23456,N_23539);
or UO_1227 (O_1227,N_23919,N_23917);
nor UO_1228 (O_1228,N_23997,N_23514);
and UO_1229 (O_1229,N_24326,N_23496);
or UO_1230 (O_1230,N_24551,N_22680);
or UO_1231 (O_1231,N_23011,N_22322);
or UO_1232 (O_1232,N_23434,N_21921);
or UO_1233 (O_1233,N_22883,N_22251);
or UO_1234 (O_1234,N_23165,N_22999);
nand UO_1235 (O_1235,N_21890,N_22651);
and UO_1236 (O_1236,N_23286,N_24357);
and UO_1237 (O_1237,N_22703,N_23100);
nor UO_1238 (O_1238,N_23070,N_24394);
nor UO_1239 (O_1239,N_24263,N_23710);
or UO_1240 (O_1240,N_24690,N_22456);
xor UO_1241 (O_1241,N_24249,N_21879);
nand UO_1242 (O_1242,N_23494,N_22098);
xnor UO_1243 (O_1243,N_23030,N_22314);
nand UO_1244 (O_1244,N_23125,N_22769);
nor UO_1245 (O_1245,N_23852,N_23721);
xnor UO_1246 (O_1246,N_21988,N_22028);
nor UO_1247 (O_1247,N_22034,N_24722);
and UO_1248 (O_1248,N_23287,N_23725);
or UO_1249 (O_1249,N_22816,N_24758);
nand UO_1250 (O_1250,N_24511,N_22024);
or UO_1251 (O_1251,N_24439,N_24269);
nand UO_1252 (O_1252,N_23124,N_22067);
or UO_1253 (O_1253,N_22540,N_23838);
nor UO_1254 (O_1254,N_23747,N_22136);
and UO_1255 (O_1255,N_22750,N_22956);
nand UO_1256 (O_1256,N_23523,N_23867);
xnor UO_1257 (O_1257,N_22179,N_24620);
and UO_1258 (O_1258,N_22609,N_21949);
nand UO_1259 (O_1259,N_22211,N_22446);
nand UO_1260 (O_1260,N_22362,N_23402);
and UO_1261 (O_1261,N_24074,N_23304);
xor UO_1262 (O_1262,N_23599,N_24302);
nor UO_1263 (O_1263,N_21983,N_22212);
xor UO_1264 (O_1264,N_22558,N_22905);
and UO_1265 (O_1265,N_22749,N_22752);
and UO_1266 (O_1266,N_24347,N_24456);
nand UO_1267 (O_1267,N_23577,N_24798);
xor UO_1268 (O_1268,N_22631,N_24621);
nor UO_1269 (O_1269,N_21996,N_22161);
and UO_1270 (O_1270,N_24991,N_24928);
and UO_1271 (O_1271,N_23034,N_22712);
nand UO_1272 (O_1272,N_22857,N_24704);
or UO_1273 (O_1273,N_24654,N_24095);
nor UO_1274 (O_1274,N_22063,N_24553);
and UO_1275 (O_1275,N_22365,N_24579);
xor UO_1276 (O_1276,N_22215,N_24697);
nor UO_1277 (O_1277,N_24560,N_24339);
and UO_1278 (O_1278,N_22880,N_22516);
nor UO_1279 (O_1279,N_24234,N_23708);
or UO_1280 (O_1280,N_24971,N_22216);
nor UO_1281 (O_1281,N_23352,N_23989);
and UO_1282 (O_1282,N_23915,N_22004);
and UO_1283 (O_1283,N_24952,N_22379);
or UO_1284 (O_1284,N_22400,N_22527);
and UO_1285 (O_1285,N_23661,N_22250);
nor UO_1286 (O_1286,N_23743,N_24777);
nor UO_1287 (O_1287,N_21955,N_24221);
xor UO_1288 (O_1288,N_24464,N_23374);
nand UO_1289 (O_1289,N_23755,N_24290);
xor UO_1290 (O_1290,N_23366,N_24176);
xor UO_1291 (O_1291,N_23540,N_22670);
or UO_1292 (O_1292,N_24178,N_22851);
xor UO_1293 (O_1293,N_23670,N_23215);
nor UO_1294 (O_1294,N_23832,N_23263);
nor UO_1295 (O_1295,N_23874,N_23913);
or UO_1296 (O_1296,N_22666,N_24888);
nand UO_1297 (O_1297,N_24137,N_24401);
or UO_1298 (O_1298,N_23158,N_22567);
nor UO_1299 (O_1299,N_22195,N_22911);
or UO_1300 (O_1300,N_22813,N_24225);
and UO_1301 (O_1301,N_23138,N_24969);
xnor UO_1302 (O_1302,N_22109,N_24997);
xnor UO_1303 (O_1303,N_24541,N_22044);
xor UO_1304 (O_1304,N_24200,N_21982);
and UO_1305 (O_1305,N_22273,N_23749);
and UO_1306 (O_1306,N_24792,N_21939);
or UO_1307 (O_1307,N_23806,N_21934);
xnor UO_1308 (O_1308,N_22800,N_24589);
nand UO_1309 (O_1309,N_23618,N_23797);
nand UO_1310 (O_1310,N_24301,N_22295);
and UO_1311 (O_1311,N_23790,N_24194);
nand UO_1312 (O_1312,N_22844,N_23420);
or UO_1313 (O_1313,N_22809,N_24444);
nor UO_1314 (O_1314,N_24297,N_21896);
nor UO_1315 (O_1315,N_22293,N_22739);
nand UO_1316 (O_1316,N_24334,N_23554);
or UO_1317 (O_1317,N_23544,N_22296);
and UO_1318 (O_1318,N_24831,N_22480);
or UO_1319 (O_1319,N_23223,N_22817);
or UO_1320 (O_1320,N_24316,N_24923);
nor UO_1321 (O_1321,N_24485,N_23404);
xnor UO_1322 (O_1322,N_23594,N_24655);
xnor UO_1323 (O_1323,N_24496,N_23083);
nand UO_1324 (O_1324,N_22966,N_24196);
and UO_1325 (O_1325,N_23503,N_22039);
xnor UO_1326 (O_1326,N_23211,N_24543);
nand UO_1327 (O_1327,N_24285,N_24748);
nor UO_1328 (O_1328,N_21948,N_21897);
nor UO_1329 (O_1329,N_24113,N_23059);
xnor UO_1330 (O_1330,N_22799,N_24057);
nand UO_1331 (O_1331,N_22672,N_22487);
and UO_1332 (O_1332,N_22740,N_23431);
and UO_1333 (O_1333,N_23561,N_22849);
nand UO_1334 (O_1334,N_22025,N_22701);
or UO_1335 (O_1335,N_22780,N_24207);
xor UO_1336 (O_1336,N_24659,N_24859);
nor UO_1337 (O_1337,N_21888,N_22388);
or UO_1338 (O_1338,N_22095,N_24836);
or UO_1339 (O_1339,N_23098,N_21967);
nor UO_1340 (O_1340,N_23759,N_23945);
or UO_1341 (O_1341,N_23820,N_22728);
or UO_1342 (O_1342,N_22926,N_22443);
and UO_1343 (O_1343,N_23718,N_23092);
xnor UO_1344 (O_1344,N_23975,N_24378);
or UO_1345 (O_1345,N_23411,N_23394);
nand UO_1346 (O_1346,N_22193,N_23726);
and UO_1347 (O_1347,N_24781,N_23669);
or UO_1348 (O_1348,N_23676,N_24641);
or UO_1349 (O_1349,N_24857,N_24984);
and UO_1350 (O_1350,N_22167,N_22360);
xor UO_1351 (O_1351,N_23067,N_22477);
nand UO_1352 (O_1352,N_22818,N_22111);
and UO_1353 (O_1353,N_22426,N_23677);
nor UO_1354 (O_1354,N_24614,N_24395);
nand UO_1355 (O_1355,N_24224,N_24195);
and UO_1356 (O_1356,N_23482,N_23882);
xnor UO_1357 (O_1357,N_23174,N_22316);
or UO_1358 (O_1358,N_23115,N_23757);
or UO_1359 (O_1359,N_22954,N_23683);
and UO_1360 (O_1360,N_22172,N_22608);
xor UO_1361 (O_1361,N_24172,N_23891);
xor UO_1362 (O_1362,N_24245,N_22117);
nor UO_1363 (O_1363,N_23897,N_23682);
and UO_1364 (O_1364,N_21899,N_24498);
or UO_1365 (O_1365,N_24138,N_23557);
or UO_1366 (O_1366,N_24854,N_24865);
or UO_1367 (O_1367,N_22946,N_24149);
nand UO_1368 (O_1368,N_24463,N_22287);
nand UO_1369 (O_1369,N_24994,N_24597);
nor UO_1370 (O_1370,N_23922,N_24092);
or UO_1371 (O_1371,N_23066,N_24983);
xor UO_1372 (O_1372,N_22852,N_22313);
nor UO_1373 (O_1373,N_24373,N_22072);
nor UO_1374 (O_1374,N_23528,N_22658);
or UO_1375 (O_1375,N_23467,N_22684);
and UO_1376 (O_1376,N_23672,N_23641);
or UO_1377 (O_1377,N_22955,N_24410);
or UO_1378 (O_1378,N_22897,N_21936);
xor UO_1379 (O_1379,N_21947,N_23134);
nand UO_1380 (O_1380,N_22649,N_24342);
or UO_1381 (O_1381,N_24642,N_24500);
nor UO_1382 (O_1382,N_22525,N_24054);
xnor UO_1383 (O_1383,N_22995,N_22303);
and UO_1384 (O_1384,N_24292,N_22943);
or UO_1385 (O_1385,N_24849,N_22877);
or UO_1386 (O_1386,N_24665,N_24151);
nand UO_1387 (O_1387,N_24272,N_23036);
xor UO_1388 (O_1388,N_22435,N_24184);
and UO_1389 (O_1389,N_22952,N_22989);
nor UO_1390 (O_1390,N_24107,N_22696);
nor UO_1391 (O_1391,N_23866,N_23687);
or UO_1392 (O_1392,N_22478,N_23377);
and UO_1393 (O_1393,N_22827,N_24720);
or UO_1394 (O_1394,N_23148,N_22768);
or UO_1395 (O_1395,N_23636,N_22038);
nor UO_1396 (O_1396,N_24771,N_22090);
nand UO_1397 (O_1397,N_24391,N_22375);
nor UO_1398 (O_1398,N_23689,N_24821);
nor UO_1399 (O_1399,N_22147,N_24752);
nor UO_1400 (O_1400,N_24025,N_24392);
nor UO_1401 (O_1401,N_23270,N_22263);
nor UO_1402 (O_1402,N_24562,N_22452);
xor UO_1403 (O_1403,N_21917,N_23427);
or UO_1404 (O_1404,N_22828,N_24674);
and UO_1405 (O_1405,N_21941,N_23835);
nor UO_1406 (O_1406,N_24246,N_22704);
nor UO_1407 (O_1407,N_23462,N_23000);
nor UO_1408 (O_1408,N_24894,N_23146);
or UO_1409 (O_1409,N_23493,N_22122);
xor UO_1410 (O_1410,N_22411,N_23516);
xnor UO_1411 (O_1411,N_24434,N_24106);
nor UO_1412 (O_1412,N_24331,N_22735);
nor UO_1413 (O_1413,N_23776,N_23298);
nor UO_1414 (O_1414,N_24564,N_22616);
nor UO_1415 (O_1415,N_23192,N_24426);
and UO_1416 (O_1416,N_22551,N_22916);
and UO_1417 (O_1417,N_24408,N_24617);
nor UO_1418 (O_1418,N_22509,N_24586);
xor UO_1419 (O_1419,N_23216,N_22642);
or UO_1420 (O_1420,N_23798,N_22094);
or UO_1421 (O_1421,N_22951,N_24762);
nor UO_1422 (O_1422,N_22595,N_22057);
nand UO_1423 (O_1423,N_21962,N_22734);
or UO_1424 (O_1424,N_24510,N_24387);
nand UO_1425 (O_1425,N_24606,N_22736);
nor UO_1426 (O_1426,N_21918,N_23727);
xnor UO_1427 (O_1427,N_24537,N_24574);
and UO_1428 (O_1428,N_23953,N_23678);
nor UO_1429 (O_1429,N_22257,N_23695);
xor UO_1430 (O_1430,N_24847,N_24058);
nand UO_1431 (O_1431,N_23013,N_23383);
xor UO_1432 (O_1432,N_22929,N_23195);
and UO_1433 (O_1433,N_22668,N_23605);
or UO_1434 (O_1434,N_22081,N_22202);
and UO_1435 (O_1435,N_24664,N_22271);
nand UO_1436 (O_1436,N_22974,N_22190);
xnor UO_1437 (O_1437,N_22199,N_22140);
nor UO_1438 (O_1438,N_24689,N_23884);
and UO_1439 (O_1439,N_22833,N_24683);
xnor UO_1440 (O_1440,N_22050,N_23628);
or UO_1441 (O_1441,N_22218,N_22256);
and UO_1442 (O_1442,N_23113,N_23713);
nor UO_1443 (O_1443,N_22861,N_24457);
or UO_1444 (O_1444,N_23324,N_22733);
nor UO_1445 (O_1445,N_23441,N_23003);
nor UO_1446 (O_1446,N_23861,N_24083);
or UO_1447 (O_1447,N_22196,N_22690);
xnor UO_1448 (O_1448,N_22214,N_22657);
xnor UO_1449 (O_1449,N_24534,N_21964);
xnor UO_1450 (O_1450,N_24250,N_24725);
nand UO_1451 (O_1451,N_24218,N_23908);
or UO_1452 (O_1452,N_22630,N_22131);
or UO_1453 (O_1453,N_23392,N_22664);
nand UO_1454 (O_1454,N_22059,N_23069);
xor UO_1455 (O_1455,N_24097,N_24322);
nor UO_1456 (O_1456,N_24829,N_22961);
nor UO_1457 (O_1457,N_24891,N_23154);
nand UO_1458 (O_1458,N_22502,N_22918);
nor UO_1459 (O_1459,N_24681,N_22468);
xor UO_1460 (O_1460,N_24875,N_24816);
nor UO_1461 (O_1461,N_24262,N_23844);
nor UO_1462 (O_1462,N_23914,N_24603);
nor UO_1463 (O_1463,N_22573,N_22008);
and UO_1464 (O_1464,N_22128,N_24677);
or UO_1465 (O_1465,N_22107,N_24167);
xor UO_1466 (O_1466,N_23696,N_24182);
and UO_1467 (O_1467,N_23001,N_23717);
or UO_1468 (O_1468,N_24180,N_24142);
or UO_1469 (O_1469,N_24612,N_23273);
xnor UO_1470 (O_1470,N_22810,N_22745);
nand UO_1471 (O_1471,N_23722,N_22879);
xor UO_1472 (O_1472,N_22782,N_23954);
nand UO_1473 (O_1473,N_23596,N_23323);
nand UO_1474 (O_1474,N_22626,N_21942);
nand UO_1475 (O_1475,N_24896,N_24583);
and UO_1476 (O_1476,N_24489,N_23625);
and UO_1477 (O_1477,N_22402,N_23834);
or UO_1478 (O_1478,N_23728,N_23116);
xnor UO_1479 (O_1479,N_22347,N_24315);
nand UO_1480 (O_1480,N_24374,N_23114);
xor UO_1481 (O_1481,N_23871,N_22408);
xor UO_1482 (O_1482,N_23924,N_22162);
nand UO_1483 (O_1483,N_24756,N_24124);
xnor UO_1484 (O_1484,N_22777,N_22845);
and UO_1485 (O_1485,N_22829,N_22760);
and UO_1486 (O_1486,N_24753,N_22831);
xor UO_1487 (O_1487,N_24365,N_22206);
nor UO_1488 (O_1488,N_24585,N_23330);
nor UO_1489 (O_1489,N_22719,N_22100);
and UO_1490 (O_1490,N_23222,N_23706);
xor UO_1491 (O_1491,N_23409,N_22535);
nand UO_1492 (O_1492,N_24433,N_22143);
nor UO_1493 (O_1493,N_22726,N_24188);
xor UO_1494 (O_1494,N_22972,N_24565);
nor UO_1495 (O_1495,N_24041,N_22930);
or UO_1496 (O_1496,N_22771,N_24452);
or UO_1497 (O_1497,N_23958,N_24990);
xnor UO_1498 (O_1498,N_24549,N_22867);
nor UO_1499 (O_1499,N_22858,N_22101);
nand UO_1500 (O_1500,N_23921,N_24273);
or UO_1501 (O_1501,N_23248,N_22352);
and UO_1502 (O_1502,N_22890,N_24842);
and UO_1503 (O_1503,N_24747,N_24418);
xor UO_1504 (O_1504,N_24006,N_24397);
or UO_1505 (O_1505,N_22808,N_23622);
or UO_1506 (O_1506,N_24484,N_24862);
or UO_1507 (O_1507,N_21961,N_24663);
and UO_1508 (O_1508,N_23936,N_22536);
or UO_1509 (O_1509,N_23541,N_22875);
and UO_1510 (O_1510,N_23243,N_24550);
or UO_1511 (O_1511,N_24787,N_24723);
nand UO_1512 (O_1512,N_22756,N_24405);
and UO_1513 (O_1513,N_23319,N_24266);
nor UO_1514 (O_1514,N_23349,N_22422);
nor UO_1515 (O_1515,N_24299,N_23260);
and UO_1516 (O_1516,N_22545,N_22811);
nand UO_1517 (O_1517,N_22157,N_22537);
and UO_1518 (O_1518,N_24605,N_24090);
xnor UO_1519 (O_1519,N_24011,N_23310);
xnor UO_1520 (O_1520,N_24212,N_22255);
nor UO_1521 (O_1521,N_21882,N_23530);
nand UO_1522 (O_1522,N_23006,N_24675);
and UO_1523 (O_1523,N_24473,N_23068);
nor UO_1524 (O_1524,N_23418,N_23879);
or UO_1525 (O_1525,N_22544,N_24491);
xnor UO_1526 (O_1526,N_23565,N_22797);
nor UO_1527 (O_1527,N_23553,N_22958);
or UO_1528 (O_1528,N_24942,N_24265);
nand UO_1529 (O_1529,N_24390,N_23132);
and UO_1530 (O_1530,N_23931,N_23292);
nand UO_1531 (O_1531,N_23426,N_23343);
and UO_1532 (O_1532,N_24613,N_24622);
nand UO_1533 (O_1533,N_23807,N_24412);
nor UO_1534 (O_1534,N_22553,N_22323);
nor UO_1535 (O_1535,N_22770,N_24807);
or UO_1536 (O_1536,N_22116,N_23587);
xor UO_1537 (O_1537,N_23644,N_24440);
or UO_1538 (O_1538,N_22671,N_24958);
nor UO_1539 (O_1539,N_23548,N_24628);
xnor UO_1540 (O_1540,N_22392,N_24414);
xnor UO_1541 (O_1541,N_23123,N_22644);
nor UO_1542 (O_1542,N_23204,N_23205);
nor UO_1543 (O_1543,N_22222,N_23675);
and UO_1544 (O_1544,N_22928,N_24032);
xor UO_1545 (O_1545,N_21974,N_22491);
nand UO_1546 (O_1546,N_22978,N_23474);
nor UO_1547 (O_1547,N_24061,N_22037);
nand UO_1548 (O_1548,N_24638,N_24878);
xnor UO_1549 (O_1549,N_24487,N_24735);
nand UO_1550 (O_1550,N_24459,N_24509);
nand UO_1551 (O_1551,N_23789,N_23018);
and UO_1552 (O_1552,N_22377,N_24870);
xnor UO_1553 (O_1553,N_22830,N_23413);
or UO_1554 (O_1554,N_22272,N_24768);
and UO_1555 (O_1555,N_22963,N_24284);
xor UO_1556 (O_1556,N_21997,N_23610);
nor UO_1557 (O_1557,N_22185,N_24938);
or UO_1558 (O_1558,N_23121,N_24437);
or UO_1559 (O_1559,N_22656,N_22425);
or UO_1560 (O_1560,N_23028,N_22437);
xor UO_1561 (O_1561,N_23933,N_23665);
xor UO_1562 (O_1562,N_24002,N_22295);
xnor UO_1563 (O_1563,N_24953,N_23371);
nor UO_1564 (O_1564,N_24461,N_22402);
xor UO_1565 (O_1565,N_22639,N_22001);
xnor UO_1566 (O_1566,N_22008,N_22526);
and UO_1567 (O_1567,N_22718,N_21923);
nor UO_1568 (O_1568,N_24403,N_22678);
and UO_1569 (O_1569,N_22560,N_22064);
and UO_1570 (O_1570,N_22470,N_24517);
nand UO_1571 (O_1571,N_24661,N_23123);
xor UO_1572 (O_1572,N_22068,N_22024);
and UO_1573 (O_1573,N_24089,N_22937);
and UO_1574 (O_1574,N_24243,N_23499);
and UO_1575 (O_1575,N_22292,N_24237);
and UO_1576 (O_1576,N_23957,N_22379);
or UO_1577 (O_1577,N_22214,N_23613);
nand UO_1578 (O_1578,N_23885,N_24742);
nand UO_1579 (O_1579,N_22077,N_22252);
nor UO_1580 (O_1580,N_22538,N_24210);
nand UO_1581 (O_1581,N_22944,N_24826);
nand UO_1582 (O_1582,N_24264,N_23445);
or UO_1583 (O_1583,N_24413,N_23751);
or UO_1584 (O_1584,N_22820,N_22391);
nand UO_1585 (O_1585,N_23940,N_24584);
nor UO_1586 (O_1586,N_22332,N_23681);
nor UO_1587 (O_1587,N_23472,N_22262);
nor UO_1588 (O_1588,N_24668,N_24994);
or UO_1589 (O_1589,N_23153,N_24180);
xor UO_1590 (O_1590,N_24751,N_23351);
and UO_1591 (O_1591,N_24748,N_24239);
nand UO_1592 (O_1592,N_23230,N_24484);
and UO_1593 (O_1593,N_23167,N_24995);
nand UO_1594 (O_1594,N_23783,N_23472);
xnor UO_1595 (O_1595,N_23213,N_24679);
nand UO_1596 (O_1596,N_23580,N_22343);
xnor UO_1597 (O_1597,N_23275,N_23854);
and UO_1598 (O_1598,N_24302,N_22249);
nor UO_1599 (O_1599,N_22456,N_23451);
and UO_1600 (O_1600,N_22133,N_24359);
and UO_1601 (O_1601,N_24348,N_23942);
and UO_1602 (O_1602,N_24213,N_22720);
nor UO_1603 (O_1603,N_24550,N_22009);
or UO_1604 (O_1604,N_23685,N_22889);
nor UO_1605 (O_1605,N_23505,N_23539);
nand UO_1606 (O_1606,N_24342,N_24913);
nor UO_1607 (O_1607,N_23038,N_23122);
nor UO_1608 (O_1608,N_22032,N_23742);
xnor UO_1609 (O_1609,N_24800,N_24273);
nor UO_1610 (O_1610,N_24240,N_22630);
and UO_1611 (O_1611,N_22017,N_22648);
nand UO_1612 (O_1612,N_23970,N_24377);
xnor UO_1613 (O_1613,N_21990,N_23736);
and UO_1614 (O_1614,N_24188,N_22000);
or UO_1615 (O_1615,N_23445,N_24636);
xnor UO_1616 (O_1616,N_22014,N_23629);
nand UO_1617 (O_1617,N_22029,N_24937);
and UO_1618 (O_1618,N_24948,N_24860);
nor UO_1619 (O_1619,N_23725,N_24537);
xor UO_1620 (O_1620,N_23886,N_23891);
nor UO_1621 (O_1621,N_24423,N_23540);
or UO_1622 (O_1622,N_24815,N_23102);
xor UO_1623 (O_1623,N_23306,N_24130);
nand UO_1624 (O_1624,N_23171,N_21913);
and UO_1625 (O_1625,N_24716,N_23364);
nor UO_1626 (O_1626,N_22214,N_23724);
xnor UO_1627 (O_1627,N_22940,N_22564);
xnor UO_1628 (O_1628,N_24804,N_24420);
nand UO_1629 (O_1629,N_23834,N_24828);
or UO_1630 (O_1630,N_23840,N_22029);
nand UO_1631 (O_1631,N_23029,N_24106);
nand UO_1632 (O_1632,N_23858,N_23054);
nor UO_1633 (O_1633,N_23611,N_23826);
nand UO_1634 (O_1634,N_22961,N_22156);
nand UO_1635 (O_1635,N_23499,N_22456);
nand UO_1636 (O_1636,N_22849,N_23643);
and UO_1637 (O_1637,N_22150,N_23780);
nand UO_1638 (O_1638,N_23629,N_24874);
or UO_1639 (O_1639,N_23984,N_24680);
and UO_1640 (O_1640,N_23265,N_23202);
and UO_1641 (O_1641,N_23957,N_22517);
nor UO_1642 (O_1642,N_24705,N_23755);
nor UO_1643 (O_1643,N_24813,N_23539);
and UO_1644 (O_1644,N_22102,N_23657);
xor UO_1645 (O_1645,N_24383,N_21895);
xnor UO_1646 (O_1646,N_24060,N_23838);
xnor UO_1647 (O_1647,N_23858,N_23089);
nand UO_1648 (O_1648,N_24535,N_24808);
nand UO_1649 (O_1649,N_24436,N_23881);
and UO_1650 (O_1650,N_24543,N_23981);
and UO_1651 (O_1651,N_23549,N_23849);
or UO_1652 (O_1652,N_24213,N_23788);
nand UO_1653 (O_1653,N_24553,N_23403);
or UO_1654 (O_1654,N_23689,N_23848);
xor UO_1655 (O_1655,N_24912,N_23665);
or UO_1656 (O_1656,N_23812,N_24047);
and UO_1657 (O_1657,N_24713,N_22175);
xor UO_1658 (O_1658,N_23150,N_22795);
xnor UO_1659 (O_1659,N_22510,N_24330);
nand UO_1660 (O_1660,N_23118,N_23963);
nor UO_1661 (O_1661,N_24763,N_23186);
nor UO_1662 (O_1662,N_24270,N_24362);
or UO_1663 (O_1663,N_24928,N_24662);
nand UO_1664 (O_1664,N_23740,N_23981);
xor UO_1665 (O_1665,N_22804,N_24078);
or UO_1666 (O_1666,N_23773,N_24200);
and UO_1667 (O_1667,N_23283,N_23801);
xor UO_1668 (O_1668,N_24481,N_24188);
nand UO_1669 (O_1669,N_22062,N_23316);
nor UO_1670 (O_1670,N_24277,N_23390);
nor UO_1671 (O_1671,N_23231,N_21889);
xnor UO_1672 (O_1672,N_22658,N_23870);
or UO_1673 (O_1673,N_22956,N_22259);
or UO_1674 (O_1674,N_22364,N_23037);
xor UO_1675 (O_1675,N_22014,N_23206);
xnor UO_1676 (O_1676,N_23424,N_23291);
and UO_1677 (O_1677,N_24534,N_24768);
nor UO_1678 (O_1678,N_24143,N_23356);
nand UO_1679 (O_1679,N_23899,N_22418);
nand UO_1680 (O_1680,N_22090,N_23232);
or UO_1681 (O_1681,N_23915,N_23953);
xor UO_1682 (O_1682,N_23462,N_22967);
xnor UO_1683 (O_1683,N_22160,N_22709);
xor UO_1684 (O_1684,N_22152,N_24758);
and UO_1685 (O_1685,N_21961,N_23729);
nor UO_1686 (O_1686,N_24446,N_22245);
or UO_1687 (O_1687,N_24901,N_24322);
nor UO_1688 (O_1688,N_23380,N_24241);
xor UO_1689 (O_1689,N_24202,N_23042);
nor UO_1690 (O_1690,N_23745,N_22230);
or UO_1691 (O_1691,N_23819,N_22750);
and UO_1692 (O_1692,N_22463,N_23795);
and UO_1693 (O_1693,N_24844,N_22970);
xnor UO_1694 (O_1694,N_22614,N_24703);
nor UO_1695 (O_1695,N_24628,N_23067);
xnor UO_1696 (O_1696,N_23318,N_23821);
or UO_1697 (O_1697,N_24703,N_23406);
or UO_1698 (O_1698,N_22440,N_21922);
xnor UO_1699 (O_1699,N_22510,N_22164);
or UO_1700 (O_1700,N_23779,N_23017);
nor UO_1701 (O_1701,N_23193,N_24008);
or UO_1702 (O_1702,N_24707,N_22912);
and UO_1703 (O_1703,N_24609,N_22132);
nand UO_1704 (O_1704,N_22404,N_22819);
or UO_1705 (O_1705,N_22861,N_22662);
nand UO_1706 (O_1706,N_23967,N_24433);
nand UO_1707 (O_1707,N_23722,N_23521);
nor UO_1708 (O_1708,N_22123,N_22255);
and UO_1709 (O_1709,N_24701,N_21883);
xnor UO_1710 (O_1710,N_22852,N_22353);
or UO_1711 (O_1711,N_24386,N_24944);
nor UO_1712 (O_1712,N_21966,N_24656);
nor UO_1713 (O_1713,N_22133,N_24971);
nand UO_1714 (O_1714,N_21967,N_22746);
nand UO_1715 (O_1715,N_24448,N_22409);
and UO_1716 (O_1716,N_24421,N_24098);
nor UO_1717 (O_1717,N_23302,N_24832);
nand UO_1718 (O_1718,N_24426,N_22125);
nor UO_1719 (O_1719,N_22787,N_23766);
and UO_1720 (O_1720,N_22219,N_24741);
xnor UO_1721 (O_1721,N_24394,N_22779);
nor UO_1722 (O_1722,N_22659,N_22435);
and UO_1723 (O_1723,N_23005,N_23104);
nor UO_1724 (O_1724,N_23695,N_24418);
xnor UO_1725 (O_1725,N_24663,N_22740);
nor UO_1726 (O_1726,N_24063,N_24760);
and UO_1727 (O_1727,N_24709,N_22526);
nand UO_1728 (O_1728,N_24540,N_22348);
nor UO_1729 (O_1729,N_23356,N_24523);
or UO_1730 (O_1730,N_23566,N_23032);
nand UO_1731 (O_1731,N_22078,N_23437);
and UO_1732 (O_1732,N_21931,N_23957);
and UO_1733 (O_1733,N_23115,N_23954);
xor UO_1734 (O_1734,N_22055,N_23023);
and UO_1735 (O_1735,N_23207,N_23195);
xnor UO_1736 (O_1736,N_24410,N_24172);
xnor UO_1737 (O_1737,N_24126,N_23721);
and UO_1738 (O_1738,N_24180,N_22475);
nor UO_1739 (O_1739,N_23395,N_22807);
and UO_1740 (O_1740,N_23429,N_22602);
and UO_1741 (O_1741,N_22990,N_23010);
nor UO_1742 (O_1742,N_22981,N_23037);
nor UO_1743 (O_1743,N_23344,N_24637);
xor UO_1744 (O_1744,N_22719,N_22684);
nor UO_1745 (O_1745,N_22945,N_23832);
and UO_1746 (O_1746,N_24245,N_24569);
xor UO_1747 (O_1747,N_24940,N_22178);
xnor UO_1748 (O_1748,N_23209,N_24913);
and UO_1749 (O_1749,N_22856,N_22592);
xor UO_1750 (O_1750,N_24385,N_24332);
nor UO_1751 (O_1751,N_22115,N_23835);
nor UO_1752 (O_1752,N_22377,N_24488);
xor UO_1753 (O_1753,N_22744,N_23745);
and UO_1754 (O_1754,N_22022,N_24990);
xnor UO_1755 (O_1755,N_24476,N_24022);
xnor UO_1756 (O_1756,N_22718,N_22697);
nor UO_1757 (O_1757,N_24870,N_22526);
and UO_1758 (O_1758,N_23872,N_22555);
xor UO_1759 (O_1759,N_23220,N_24782);
or UO_1760 (O_1760,N_22395,N_23914);
or UO_1761 (O_1761,N_22363,N_22720);
xnor UO_1762 (O_1762,N_22109,N_23650);
nor UO_1763 (O_1763,N_23747,N_22627);
and UO_1764 (O_1764,N_23574,N_24332);
nand UO_1765 (O_1765,N_22498,N_23820);
and UO_1766 (O_1766,N_22106,N_23610);
nand UO_1767 (O_1767,N_23303,N_23464);
nand UO_1768 (O_1768,N_23712,N_23572);
xnor UO_1769 (O_1769,N_23672,N_22895);
nor UO_1770 (O_1770,N_24053,N_24026);
nand UO_1771 (O_1771,N_22493,N_23686);
nor UO_1772 (O_1772,N_23750,N_22804);
xor UO_1773 (O_1773,N_23892,N_23125);
nor UO_1774 (O_1774,N_24529,N_24915);
nand UO_1775 (O_1775,N_23954,N_24707);
nand UO_1776 (O_1776,N_22641,N_24061);
xnor UO_1777 (O_1777,N_22920,N_24358);
xnor UO_1778 (O_1778,N_23843,N_23601);
nand UO_1779 (O_1779,N_22920,N_22881);
or UO_1780 (O_1780,N_23793,N_24763);
nand UO_1781 (O_1781,N_23223,N_24503);
nand UO_1782 (O_1782,N_23888,N_22238);
xor UO_1783 (O_1783,N_22696,N_21981);
nand UO_1784 (O_1784,N_23232,N_24517);
nand UO_1785 (O_1785,N_22486,N_23410);
or UO_1786 (O_1786,N_22053,N_23947);
nor UO_1787 (O_1787,N_23938,N_23399);
or UO_1788 (O_1788,N_23924,N_22157);
xnor UO_1789 (O_1789,N_22164,N_24608);
xor UO_1790 (O_1790,N_22496,N_23807);
nand UO_1791 (O_1791,N_24509,N_24546);
nand UO_1792 (O_1792,N_24895,N_22842);
xnor UO_1793 (O_1793,N_23434,N_24552);
xor UO_1794 (O_1794,N_23281,N_24539);
nor UO_1795 (O_1795,N_23306,N_23626);
nor UO_1796 (O_1796,N_24327,N_24574);
and UO_1797 (O_1797,N_22449,N_23638);
nor UO_1798 (O_1798,N_23179,N_22601);
and UO_1799 (O_1799,N_23977,N_23231);
xor UO_1800 (O_1800,N_22821,N_21954);
or UO_1801 (O_1801,N_23609,N_24194);
or UO_1802 (O_1802,N_24064,N_23445);
nand UO_1803 (O_1803,N_24222,N_22916);
or UO_1804 (O_1804,N_23988,N_24247);
or UO_1805 (O_1805,N_24826,N_22546);
or UO_1806 (O_1806,N_22077,N_24610);
xnor UO_1807 (O_1807,N_24447,N_22946);
nor UO_1808 (O_1808,N_24686,N_22241);
nand UO_1809 (O_1809,N_24512,N_23981);
and UO_1810 (O_1810,N_23016,N_23284);
and UO_1811 (O_1811,N_24499,N_24559);
nand UO_1812 (O_1812,N_24368,N_22797);
xnor UO_1813 (O_1813,N_22970,N_23708);
nor UO_1814 (O_1814,N_21961,N_23844);
nor UO_1815 (O_1815,N_22754,N_22011);
xor UO_1816 (O_1816,N_22754,N_23505);
xor UO_1817 (O_1817,N_23571,N_24170);
and UO_1818 (O_1818,N_23296,N_24135);
nor UO_1819 (O_1819,N_24362,N_22607);
or UO_1820 (O_1820,N_24629,N_24282);
nor UO_1821 (O_1821,N_24742,N_23438);
or UO_1822 (O_1822,N_22946,N_22327);
xor UO_1823 (O_1823,N_22558,N_24203);
nor UO_1824 (O_1824,N_22999,N_24441);
xor UO_1825 (O_1825,N_24062,N_24534);
and UO_1826 (O_1826,N_21995,N_24220);
xnor UO_1827 (O_1827,N_22366,N_23765);
xor UO_1828 (O_1828,N_23258,N_24025);
and UO_1829 (O_1829,N_24777,N_22890);
and UO_1830 (O_1830,N_24406,N_24033);
and UO_1831 (O_1831,N_21919,N_23707);
xor UO_1832 (O_1832,N_23663,N_24504);
xor UO_1833 (O_1833,N_24457,N_21994);
or UO_1834 (O_1834,N_23252,N_23038);
or UO_1835 (O_1835,N_24790,N_24000);
nand UO_1836 (O_1836,N_22232,N_23635);
nor UO_1837 (O_1837,N_21928,N_22655);
or UO_1838 (O_1838,N_22624,N_22917);
xnor UO_1839 (O_1839,N_22293,N_23561);
or UO_1840 (O_1840,N_22968,N_24367);
xnor UO_1841 (O_1841,N_22312,N_23994);
or UO_1842 (O_1842,N_24364,N_23008);
and UO_1843 (O_1843,N_24950,N_23285);
nor UO_1844 (O_1844,N_22096,N_24438);
nand UO_1845 (O_1845,N_24146,N_23821);
and UO_1846 (O_1846,N_22644,N_22214);
or UO_1847 (O_1847,N_22371,N_24831);
nand UO_1848 (O_1848,N_21884,N_24707);
or UO_1849 (O_1849,N_24130,N_24338);
or UO_1850 (O_1850,N_21931,N_23082);
nand UO_1851 (O_1851,N_22977,N_22059);
nand UO_1852 (O_1852,N_22407,N_22769);
nor UO_1853 (O_1853,N_24716,N_21943);
nor UO_1854 (O_1854,N_24338,N_22879);
nor UO_1855 (O_1855,N_24750,N_24201);
nand UO_1856 (O_1856,N_22660,N_23785);
or UO_1857 (O_1857,N_23162,N_23456);
xor UO_1858 (O_1858,N_24868,N_24505);
or UO_1859 (O_1859,N_22635,N_24250);
nor UO_1860 (O_1860,N_23692,N_24864);
xnor UO_1861 (O_1861,N_23118,N_23651);
nor UO_1862 (O_1862,N_23728,N_22270);
nand UO_1863 (O_1863,N_23931,N_24426);
or UO_1864 (O_1864,N_23111,N_23835);
nand UO_1865 (O_1865,N_23277,N_23070);
or UO_1866 (O_1866,N_23411,N_21921);
nand UO_1867 (O_1867,N_22068,N_23927);
nor UO_1868 (O_1868,N_22332,N_23445);
nor UO_1869 (O_1869,N_24684,N_22141);
or UO_1870 (O_1870,N_21884,N_24795);
nand UO_1871 (O_1871,N_23541,N_23938);
or UO_1872 (O_1872,N_22085,N_22060);
or UO_1873 (O_1873,N_23111,N_22317);
nor UO_1874 (O_1874,N_24920,N_23157);
and UO_1875 (O_1875,N_23333,N_24711);
and UO_1876 (O_1876,N_21879,N_23236);
nand UO_1877 (O_1877,N_22727,N_24819);
or UO_1878 (O_1878,N_24603,N_23979);
nand UO_1879 (O_1879,N_21921,N_24417);
and UO_1880 (O_1880,N_24144,N_23467);
or UO_1881 (O_1881,N_23006,N_22002);
nand UO_1882 (O_1882,N_23968,N_23522);
nor UO_1883 (O_1883,N_22002,N_24740);
and UO_1884 (O_1884,N_23011,N_24141);
or UO_1885 (O_1885,N_22122,N_24096);
xnor UO_1886 (O_1886,N_22981,N_22657);
nor UO_1887 (O_1887,N_22903,N_23021);
nand UO_1888 (O_1888,N_22097,N_23388);
or UO_1889 (O_1889,N_23060,N_24933);
nor UO_1890 (O_1890,N_24322,N_23412);
or UO_1891 (O_1891,N_22068,N_23007);
and UO_1892 (O_1892,N_24010,N_22792);
xor UO_1893 (O_1893,N_23055,N_23966);
xor UO_1894 (O_1894,N_24864,N_24185);
and UO_1895 (O_1895,N_23179,N_24568);
xnor UO_1896 (O_1896,N_24139,N_24224);
nand UO_1897 (O_1897,N_23763,N_24339);
xor UO_1898 (O_1898,N_23695,N_21924);
and UO_1899 (O_1899,N_22151,N_24423);
nor UO_1900 (O_1900,N_23529,N_24388);
nand UO_1901 (O_1901,N_23015,N_22047);
and UO_1902 (O_1902,N_23167,N_22649);
or UO_1903 (O_1903,N_23208,N_24408);
nor UO_1904 (O_1904,N_24001,N_24692);
and UO_1905 (O_1905,N_23743,N_23575);
nor UO_1906 (O_1906,N_23906,N_23359);
nor UO_1907 (O_1907,N_22297,N_24570);
xnor UO_1908 (O_1908,N_22465,N_22485);
xnor UO_1909 (O_1909,N_22792,N_23588);
xor UO_1910 (O_1910,N_24078,N_23005);
nand UO_1911 (O_1911,N_23787,N_22700);
nor UO_1912 (O_1912,N_23490,N_23901);
and UO_1913 (O_1913,N_24619,N_22402);
xnor UO_1914 (O_1914,N_24791,N_23364);
nand UO_1915 (O_1915,N_22416,N_24480);
nor UO_1916 (O_1916,N_24614,N_23227);
nor UO_1917 (O_1917,N_24109,N_24869);
xor UO_1918 (O_1918,N_23552,N_24905);
or UO_1919 (O_1919,N_22923,N_24278);
xor UO_1920 (O_1920,N_24885,N_23566);
or UO_1921 (O_1921,N_22513,N_23637);
and UO_1922 (O_1922,N_22946,N_22308);
xnor UO_1923 (O_1923,N_23526,N_22552);
or UO_1924 (O_1924,N_22833,N_24054);
and UO_1925 (O_1925,N_24167,N_24185);
and UO_1926 (O_1926,N_23741,N_22408);
xor UO_1927 (O_1927,N_22528,N_23792);
nand UO_1928 (O_1928,N_23947,N_21903);
and UO_1929 (O_1929,N_23651,N_24863);
and UO_1930 (O_1930,N_24334,N_24053);
xnor UO_1931 (O_1931,N_21988,N_23279);
and UO_1932 (O_1932,N_23737,N_24780);
or UO_1933 (O_1933,N_22427,N_22969);
or UO_1934 (O_1934,N_22791,N_24664);
or UO_1935 (O_1935,N_23416,N_22181);
nand UO_1936 (O_1936,N_22449,N_23262);
xnor UO_1937 (O_1937,N_24358,N_24543);
nand UO_1938 (O_1938,N_22488,N_23614);
xor UO_1939 (O_1939,N_24823,N_24194);
nand UO_1940 (O_1940,N_24997,N_23011);
xnor UO_1941 (O_1941,N_22159,N_24887);
nor UO_1942 (O_1942,N_24301,N_23888);
and UO_1943 (O_1943,N_24785,N_22770);
nand UO_1944 (O_1944,N_22347,N_22918);
xor UO_1945 (O_1945,N_22349,N_23555);
xor UO_1946 (O_1946,N_21968,N_22120);
or UO_1947 (O_1947,N_24590,N_23899);
nor UO_1948 (O_1948,N_22210,N_23348);
and UO_1949 (O_1949,N_22708,N_24026);
or UO_1950 (O_1950,N_24501,N_22286);
nor UO_1951 (O_1951,N_24024,N_22137);
or UO_1952 (O_1952,N_22665,N_23224);
or UO_1953 (O_1953,N_22947,N_22556);
and UO_1954 (O_1954,N_22964,N_23893);
nor UO_1955 (O_1955,N_23011,N_24439);
xnor UO_1956 (O_1956,N_22510,N_23580);
xor UO_1957 (O_1957,N_23281,N_24570);
nand UO_1958 (O_1958,N_23162,N_22086);
or UO_1959 (O_1959,N_23059,N_23633);
or UO_1960 (O_1960,N_24083,N_23838);
nor UO_1961 (O_1961,N_22172,N_23833);
xnor UO_1962 (O_1962,N_22258,N_23891);
or UO_1963 (O_1963,N_22159,N_22103);
xor UO_1964 (O_1964,N_24784,N_23517);
or UO_1965 (O_1965,N_23076,N_24306);
and UO_1966 (O_1966,N_22282,N_24614);
nand UO_1967 (O_1967,N_22599,N_24897);
xnor UO_1968 (O_1968,N_23037,N_24867);
nand UO_1969 (O_1969,N_22677,N_23582);
xor UO_1970 (O_1970,N_24126,N_23996);
and UO_1971 (O_1971,N_22592,N_24949);
and UO_1972 (O_1972,N_21960,N_24347);
nand UO_1973 (O_1973,N_22468,N_22776);
nor UO_1974 (O_1974,N_23845,N_22037);
nand UO_1975 (O_1975,N_23165,N_24041);
xnor UO_1976 (O_1976,N_21879,N_22865);
nor UO_1977 (O_1977,N_23527,N_24850);
xnor UO_1978 (O_1978,N_22340,N_24718);
nand UO_1979 (O_1979,N_21977,N_22531);
nand UO_1980 (O_1980,N_23155,N_23821);
and UO_1981 (O_1981,N_23507,N_24808);
and UO_1982 (O_1982,N_22977,N_22770);
nand UO_1983 (O_1983,N_24471,N_24507);
nor UO_1984 (O_1984,N_23828,N_23505);
or UO_1985 (O_1985,N_22710,N_22451);
or UO_1986 (O_1986,N_22421,N_23739);
or UO_1987 (O_1987,N_22708,N_22382);
nor UO_1988 (O_1988,N_23104,N_24239);
nor UO_1989 (O_1989,N_22397,N_24668);
nand UO_1990 (O_1990,N_22949,N_23701);
nor UO_1991 (O_1991,N_23623,N_23908);
and UO_1992 (O_1992,N_22412,N_24232);
and UO_1993 (O_1993,N_22530,N_22958);
and UO_1994 (O_1994,N_23655,N_24642);
nand UO_1995 (O_1995,N_22641,N_23433);
xnor UO_1996 (O_1996,N_22218,N_22760);
or UO_1997 (O_1997,N_22625,N_22287);
nand UO_1998 (O_1998,N_22271,N_22410);
or UO_1999 (O_1999,N_23669,N_24096);
nor UO_2000 (O_2000,N_22726,N_22900);
xor UO_2001 (O_2001,N_21964,N_24516);
or UO_2002 (O_2002,N_23959,N_22812);
and UO_2003 (O_2003,N_23118,N_24212);
nor UO_2004 (O_2004,N_23188,N_22427);
xor UO_2005 (O_2005,N_22022,N_24908);
or UO_2006 (O_2006,N_23287,N_23317);
nand UO_2007 (O_2007,N_23631,N_24566);
nor UO_2008 (O_2008,N_22641,N_24851);
or UO_2009 (O_2009,N_22044,N_23238);
nor UO_2010 (O_2010,N_24859,N_22570);
and UO_2011 (O_2011,N_24067,N_23704);
nor UO_2012 (O_2012,N_23541,N_23596);
xor UO_2013 (O_2013,N_24621,N_24327);
xnor UO_2014 (O_2014,N_23235,N_24670);
or UO_2015 (O_2015,N_23971,N_24941);
xor UO_2016 (O_2016,N_24551,N_22239);
and UO_2017 (O_2017,N_24105,N_24536);
or UO_2018 (O_2018,N_24908,N_22949);
nand UO_2019 (O_2019,N_24884,N_23095);
nor UO_2020 (O_2020,N_24198,N_24270);
nor UO_2021 (O_2021,N_24888,N_21914);
and UO_2022 (O_2022,N_23878,N_24813);
or UO_2023 (O_2023,N_24410,N_24645);
nand UO_2024 (O_2024,N_23525,N_24719);
nand UO_2025 (O_2025,N_22663,N_22680);
or UO_2026 (O_2026,N_24050,N_24864);
xnor UO_2027 (O_2027,N_23886,N_24343);
and UO_2028 (O_2028,N_24245,N_23637);
nand UO_2029 (O_2029,N_23311,N_23838);
or UO_2030 (O_2030,N_24150,N_23274);
nand UO_2031 (O_2031,N_24457,N_22647);
or UO_2032 (O_2032,N_24695,N_23333);
xnor UO_2033 (O_2033,N_21980,N_24692);
nand UO_2034 (O_2034,N_24927,N_21986);
nand UO_2035 (O_2035,N_23558,N_24890);
xor UO_2036 (O_2036,N_22317,N_24798);
and UO_2037 (O_2037,N_23441,N_24999);
xor UO_2038 (O_2038,N_23067,N_24684);
xor UO_2039 (O_2039,N_22030,N_23537);
nor UO_2040 (O_2040,N_22477,N_22512);
and UO_2041 (O_2041,N_22218,N_23201);
nor UO_2042 (O_2042,N_23505,N_24460);
or UO_2043 (O_2043,N_22774,N_23570);
xor UO_2044 (O_2044,N_24256,N_22050);
nand UO_2045 (O_2045,N_24090,N_23491);
and UO_2046 (O_2046,N_24898,N_23036);
or UO_2047 (O_2047,N_24393,N_24496);
or UO_2048 (O_2048,N_22423,N_24610);
xor UO_2049 (O_2049,N_22277,N_22436);
nand UO_2050 (O_2050,N_23386,N_24810);
xnor UO_2051 (O_2051,N_24558,N_24389);
and UO_2052 (O_2052,N_24915,N_24240);
nand UO_2053 (O_2053,N_22689,N_22929);
and UO_2054 (O_2054,N_24980,N_24434);
nor UO_2055 (O_2055,N_24791,N_24951);
nand UO_2056 (O_2056,N_22311,N_23822);
or UO_2057 (O_2057,N_24242,N_23487);
or UO_2058 (O_2058,N_22567,N_24411);
nand UO_2059 (O_2059,N_23702,N_24989);
nand UO_2060 (O_2060,N_22904,N_21950);
nand UO_2061 (O_2061,N_24626,N_24700);
nand UO_2062 (O_2062,N_23120,N_22187);
and UO_2063 (O_2063,N_24160,N_23665);
nor UO_2064 (O_2064,N_22496,N_22586);
nand UO_2065 (O_2065,N_23386,N_24957);
nor UO_2066 (O_2066,N_24128,N_24035);
or UO_2067 (O_2067,N_23189,N_24151);
nor UO_2068 (O_2068,N_22539,N_22541);
or UO_2069 (O_2069,N_22552,N_23295);
or UO_2070 (O_2070,N_24022,N_23798);
nand UO_2071 (O_2071,N_23053,N_23980);
or UO_2072 (O_2072,N_23148,N_24901);
and UO_2073 (O_2073,N_23658,N_23265);
or UO_2074 (O_2074,N_22005,N_24054);
nand UO_2075 (O_2075,N_23657,N_22132);
nand UO_2076 (O_2076,N_24033,N_22615);
or UO_2077 (O_2077,N_24471,N_23733);
or UO_2078 (O_2078,N_22751,N_22371);
nor UO_2079 (O_2079,N_23791,N_24431);
nand UO_2080 (O_2080,N_23795,N_24036);
or UO_2081 (O_2081,N_24834,N_22924);
and UO_2082 (O_2082,N_24466,N_22075);
or UO_2083 (O_2083,N_22477,N_24052);
or UO_2084 (O_2084,N_23616,N_22492);
or UO_2085 (O_2085,N_24839,N_24270);
xnor UO_2086 (O_2086,N_22413,N_22379);
and UO_2087 (O_2087,N_23030,N_21934);
or UO_2088 (O_2088,N_24290,N_24236);
nor UO_2089 (O_2089,N_24642,N_23630);
or UO_2090 (O_2090,N_23320,N_22709);
or UO_2091 (O_2091,N_24267,N_22783);
nand UO_2092 (O_2092,N_23144,N_22884);
xor UO_2093 (O_2093,N_23816,N_24593);
or UO_2094 (O_2094,N_23019,N_22401);
nand UO_2095 (O_2095,N_22503,N_24888);
or UO_2096 (O_2096,N_22632,N_24031);
nand UO_2097 (O_2097,N_24289,N_23016);
nand UO_2098 (O_2098,N_23855,N_24167);
xor UO_2099 (O_2099,N_24518,N_24261);
or UO_2100 (O_2100,N_24928,N_24428);
nand UO_2101 (O_2101,N_24712,N_21969);
and UO_2102 (O_2102,N_23544,N_22811);
and UO_2103 (O_2103,N_23931,N_24380);
nand UO_2104 (O_2104,N_22470,N_24851);
nor UO_2105 (O_2105,N_24409,N_23351);
or UO_2106 (O_2106,N_22656,N_24236);
and UO_2107 (O_2107,N_24029,N_23001);
xnor UO_2108 (O_2108,N_23346,N_23484);
and UO_2109 (O_2109,N_23159,N_23351);
xnor UO_2110 (O_2110,N_23909,N_21979);
and UO_2111 (O_2111,N_24547,N_23247);
nand UO_2112 (O_2112,N_21958,N_24149);
xnor UO_2113 (O_2113,N_23233,N_23583);
nor UO_2114 (O_2114,N_23910,N_22022);
and UO_2115 (O_2115,N_24247,N_24427);
nor UO_2116 (O_2116,N_21923,N_22477);
nor UO_2117 (O_2117,N_24847,N_23977);
or UO_2118 (O_2118,N_22329,N_24379);
nor UO_2119 (O_2119,N_22998,N_22919);
xnor UO_2120 (O_2120,N_23604,N_22096);
and UO_2121 (O_2121,N_22360,N_24000);
nand UO_2122 (O_2122,N_24988,N_22974);
or UO_2123 (O_2123,N_21939,N_21959);
nor UO_2124 (O_2124,N_24247,N_24445);
and UO_2125 (O_2125,N_21877,N_22430);
xor UO_2126 (O_2126,N_23296,N_22335);
nor UO_2127 (O_2127,N_22693,N_23121);
or UO_2128 (O_2128,N_24419,N_23069);
and UO_2129 (O_2129,N_24076,N_23763);
and UO_2130 (O_2130,N_22707,N_24047);
xor UO_2131 (O_2131,N_22856,N_22699);
nand UO_2132 (O_2132,N_22092,N_23683);
or UO_2133 (O_2133,N_24056,N_22146);
nand UO_2134 (O_2134,N_23176,N_24744);
nor UO_2135 (O_2135,N_22589,N_24690);
nand UO_2136 (O_2136,N_23224,N_24588);
xnor UO_2137 (O_2137,N_23895,N_22567);
nor UO_2138 (O_2138,N_23953,N_23023);
nor UO_2139 (O_2139,N_22465,N_22452);
nor UO_2140 (O_2140,N_24703,N_23087);
nand UO_2141 (O_2141,N_24843,N_22063);
nor UO_2142 (O_2142,N_23118,N_24901);
nor UO_2143 (O_2143,N_23061,N_23520);
or UO_2144 (O_2144,N_22719,N_21969);
nor UO_2145 (O_2145,N_24656,N_23281);
xor UO_2146 (O_2146,N_22400,N_24906);
nor UO_2147 (O_2147,N_24377,N_22272);
or UO_2148 (O_2148,N_24755,N_24298);
nor UO_2149 (O_2149,N_24700,N_23387);
nor UO_2150 (O_2150,N_22504,N_23970);
xor UO_2151 (O_2151,N_21990,N_24224);
nand UO_2152 (O_2152,N_23240,N_24676);
nand UO_2153 (O_2153,N_23991,N_22003);
nand UO_2154 (O_2154,N_23775,N_23604);
and UO_2155 (O_2155,N_24256,N_21896);
xnor UO_2156 (O_2156,N_24247,N_24963);
nand UO_2157 (O_2157,N_23603,N_21976);
and UO_2158 (O_2158,N_23956,N_24654);
or UO_2159 (O_2159,N_24602,N_24284);
and UO_2160 (O_2160,N_22684,N_23525);
nand UO_2161 (O_2161,N_24491,N_24230);
xnor UO_2162 (O_2162,N_22723,N_22856);
or UO_2163 (O_2163,N_24673,N_22975);
xnor UO_2164 (O_2164,N_24966,N_22649);
nand UO_2165 (O_2165,N_22347,N_23687);
nand UO_2166 (O_2166,N_23712,N_22498);
nor UO_2167 (O_2167,N_23863,N_24130);
nand UO_2168 (O_2168,N_24844,N_22623);
xnor UO_2169 (O_2169,N_23114,N_22015);
and UO_2170 (O_2170,N_22193,N_23763);
and UO_2171 (O_2171,N_24647,N_24391);
and UO_2172 (O_2172,N_23449,N_24032);
nand UO_2173 (O_2173,N_24260,N_24524);
or UO_2174 (O_2174,N_23948,N_23165);
xor UO_2175 (O_2175,N_22785,N_23941);
nor UO_2176 (O_2176,N_23093,N_22006);
nor UO_2177 (O_2177,N_23593,N_21981);
or UO_2178 (O_2178,N_23267,N_22750);
and UO_2179 (O_2179,N_24012,N_24041);
or UO_2180 (O_2180,N_22541,N_24649);
nand UO_2181 (O_2181,N_23600,N_23503);
nand UO_2182 (O_2182,N_23796,N_21938);
or UO_2183 (O_2183,N_24977,N_22521);
and UO_2184 (O_2184,N_24713,N_23998);
or UO_2185 (O_2185,N_21894,N_22810);
and UO_2186 (O_2186,N_23448,N_22473);
xnor UO_2187 (O_2187,N_23756,N_24953);
and UO_2188 (O_2188,N_23955,N_22576);
or UO_2189 (O_2189,N_24081,N_24053);
and UO_2190 (O_2190,N_24449,N_24922);
and UO_2191 (O_2191,N_24575,N_24773);
nand UO_2192 (O_2192,N_22043,N_22012);
and UO_2193 (O_2193,N_22997,N_23941);
or UO_2194 (O_2194,N_24656,N_24366);
and UO_2195 (O_2195,N_24424,N_24516);
xnor UO_2196 (O_2196,N_24308,N_21934);
and UO_2197 (O_2197,N_24204,N_22705);
nor UO_2198 (O_2198,N_23648,N_23844);
and UO_2199 (O_2199,N_22759,N_24656);
xor UO_2200 (O_2200,N_24661,N_24303);
xor UO_2201 (O_2201,N_23931,N_23562);
or UO_2202 (O_2202,N_24517,N_24950);
or UO_2203 (O_2203,N_24037,N_22636);
xor UO_2204 (O_2204,N_24198,N_22186);
and UO_2205 (O_2205,N_22164,N_23557);
xnor UO_2206 (O_2206,N_22094,N_23490);
and UO_2207 (O_2207,N_23993,N_24239);
nand UO_2208 (O_2208,N_21908,N_24575);
nor UO_2209 (O_2209,N_24268,N_23414);
nand UO_2210 (O_2210,N_23022,N_22456);
and UO_2211 (O_2211,N_23367,N_24588);
nor UO_2212 (O_2212,N_24936,N_23232);
xnor UO_2213 (O_2213,N_24487,N_24144);
xor UO_2214 (O_2214,N_22982,N_23106);
and UO_2215 (O_2215,N_22434,N_24760);
nand UO_2216 (O_2216,N_22074,N_24093);
nand UO_2217 (O_2217,N_23378,N_21966);
xnor UO_2218 (O_2218,N_23008,N_22439);
or UO_2219 (O_2219,N_24103,N_22446);
or UO_2220 (O_2220,N_22997,N_23222);
and UO_2221 (O_2221,N_22015,N_23060);
nor UO_2222 (O_2222,N_24083,N_24181);
xor UO_2223 (O_2223,N_23791,N_24006);
nor UO_2224 (O_2224,N_23806,N_23150);
and UO_2225 (O_2225,N_23892,N_23104);
or UO_2226 (O_2226,N_22540,N_23720);
and UO_2227 (O_2227,N_24563,N_23214);
nand UO_2228 (O_2228,N_24884,N_22580);
or UO_2229 (O_2229,N_24744,N_22921);
xnor UO_2230 (O_2230,N_24327,N_23198);
nor UO_2231 (O_2231,N_24901,N_23876);
nand UO_2232 (O_2232,N_23203,N_22055);
or UO_2233 (O_2233,N_23990,N_23180);
nand UO_2234 (O_2234,N_23161,N_23669);
or UO_2235 (O_2235,N_22294,N_24054);
xnor UO_2236 (O_2236,N_22176,N_23722);
xor UO_2237 (O_2237,N_22322,N_22593);
xor UO_2238 (O_2238,N_24337,N_22104);
nor UO_2239 (O_2239,N_24714,N_22158);
and UO_2240 (O_2240,N_23319,N_22755);
or UO_2241 (O_2241,N_24645,N_24057);
nand UO_2242 (O_2242,N_23320,N_24238);
or UO_2243 (O_2243,N_24357,N_24744);
and UO_2244 (O_2244,N_24425,N_22815);
xor UO_2245 (O_2245,N_24475,N_22471);
nor UO_2246 (O_2246,N_23351,N_24458);
and UO_2247 (O_2247,N_24266,N_22184);
or UO_2248 (O_2248,N_22306,N_24425);
nand UO_2249 (O_2249,N_23957,N_22124);
xnor UO_2250 (O_2250,N_22980,N_22317);
xnor UO_2251 (O_2251,N_24235,N_22123);
or UO_2252 (O_2252,N_24669,N_22434);
and UO_2253 (O_2253,N_23726,N_22428);
or UO_2254 (O_2254,N_23965,N_22603);
and UO_2255 (O_2255,N_23807,N_24446);
nor UO_2256 (O_2256,N_23379,N_22395);
nor UO_2257 (O_2257,N_24832,N_23326);
and UO_2258 (O_2258,N_22497,N_22786);
xnor UO_2259 (O_2259,N_24339,N_24627);
nor UO_2260 (O_2260,N_22742,N_23509);
nand UO_2261 (O_2261,N_22420,N_24679);
nand UO_2262 (O_2262,N_24575,N_24662);
xor UO_2263 (O_2263,N_22415,N_22829);
nand UO_2264 (O_2264,N_24318,N_23870);
nand UO_2265 (O_2265,N_24909,N_24637);
xnor UO_2266 (O_2266,N_23696,N_23748);
nor UO_2267 (O_2267,N_22655,N_23177);
and UO_2268 (O_2268,N_23854,N_22391);
nor UO_2269 (O_2269,N_24675,N_24386);
nor UO_2270 (O_2270,N_24061,N_22684);
xor UO_2271 (O_2271,N_23537,N_23955);
nor UO_2272 (O_2272,N_24939,N_24539);
or UO_2273 (O_2273,N_23028,N_22772);
or UO_2274 (O_2274,N_22624,N_24719);
or UO_2275 (O_2275,N_24020,N_24014);
or UO_2276 (O_2276,N_24651,N_24092);
or UO_2277 (O_2277,N_22990,N_23412);
and UO_2278 (O_2278,N_23226,N_22072);
and UO_2279 (O_2279,N_23714,N_24872);
and UO_2280 (O_2280,N_24415,N_23536);
and UO_2281 (O_2281,N_22310,N_23284);
or UO_2282 (O_2282,N_24616,N_22797);
xor UO_2283 (O_2283,N_22597,N_23412);
or UO_2284 (O_2284,N_23532,N_21941);
nand UO_2285 (O_2285,N_23351,N_22193);
xnor UO_2286 (O_2286,N_23607,N_24537);
or UO_2287 (O_2287,N_24208,N_23941);
nor UO_2288 (O_2288,N_22358,N_22328);
or UO_2289 (O_2289,N_24724,N_22154);
or UO_2290 (O_2290,N_24452,N_22412);
and UO_2291 (O_2291,N_21940,N_22993);
or UO_2292 (O_2292,N_24581,N_23423);
or UO_2293 (O_2293,N_24795,N_24779);
or UO_2294 (O_2294,N_24537,N_22626);
nand UO_2295 (O_2295,N_24514,N_23606);
nand UO_2296 (O_2296,N_22222,N_24136);
nor UO_2297 (O_2297,N_23220,N_22134);
nor UO_2298 (O_2298,N_22563,N_23149);
nand UO_2299 (O_2299,N_22368,N_24447);
and UO_2300 (O_2300,N_23059,N_23488);
nand UO_2301 (O_2301,N_24243,N_22961);
nor UO_2302 (O_2302,N_22063,N_24248);
nand UO_2303 (O_2303,N_23497,N_24097);
xor UO_2304 (O_2304,N_22892,N_22898);
nor UO_2305 (O_2305,N_23715,N_23813);
xor UO_2306 (O_2306,N_24776,N_22666);
nor UO_2307 (O_2307,N_24823,N_22532);
or UO_2308 (O_2308,N_23140,N_24165);
xnor UO_2309 (O_2309,N_23128,N_22676);
or UO_2310 (O_2310,N_24717,N_24460);
and UO_2311 (O_2311,N_23421,N_24773);
nand UO_2312 (O_2312,N_24807,N_24502);
or UO_2313 (O_2313,N_21901,N_24279);
or UO_2314 (O_2314,N_23048,N_22972);
nor UO_2315 (O_2315,N_22498,N_23793);
and UO_2316 (O_2316,N_23259,N_21963);
and UO_2317 (O_2317,N_23898,N_22709);
and UO_2318 (O_2318,N_24751,N_23657);
nand UO_2319 (O_2319,N_23539,N_24396);
xor UO_2320 (O_2320,N_24100,N_24634);
xnor UO_2321 (O_2321,N_22566,N_22483);
xnor UO_2322 (O_2322,N_24492,N_23378);
or UO_2323 (O_2323,N_22157,N_24177);
nor UO_2324 (O_2324,N_21962,N_24361);
nor UO_2325 (O_2325,N_24292,N_24327);
and UO_2326 (O_2326,N_24326,N_21917);
and UO_2327 (O_2327,N_22283,N_22916);
or UO_2328 (O_2328,N_24834,N_23610);
nor UO_2329 (O_2329,N_24037,N_22788);
and UO_2330 (O_2330,N_24733,N_24429);
xor UO_2331 (O_2331,N_24853,N_23888);
nand UO_2332 (O_2332,N_23764,N_21940);
and UO_2333 (O_2333,N_22895,N_23272);
nor UO_2334 (O_2334,N_23395,N_22458);
and UO_2335 (O_2335,N_23341,N_24169);
and UO_2336 (O_2336,N_24010,N_23499);
and UO_2337 (O_2337,N_23357,N_23207);
nor UO_2338 (O_2338,N_22791,N_23956);
xnor UO_2339 (O_2339,N_23312,N_23601);
or UO_2340 (O_2340,N_24540,N_22300);
and UO_2341 (O_2341,N_22000,N_23161);
or UO_2342 (O_2342,N_22250,N_23435);
nand UO_2343 (O_2343,N_23185,N_24388);
xor UO_2344 (O_2344,N_24869,N_24994);
nor UO_2345 (O_2345,N_22739,N_21976);
xnor UO_2346 (O_2346,N_24957,N_23372);
nor UO_2347 (O_2347,N_24566,N_24495);
and UO_2348 (O_2348,N_24136,N_24375);
xnor UO_2349 (O_2349,N_24757,N_24501);
nor UO_2350 (O_2350,N_22570,N_22535);
and UO_2351 (O_2351,N_23545,N_23701);
nor UO_2352 (O_2352,N_22365,N_23835);
nor UO_2353 (O_2353,N_23559,N_22800);
and UO_2354 (O_2354,N_23492,N_24472);
xor UO_2355 (O_2355,N_21964,N_22006);
nand UO_2356 (O_2356,N_22510,N_24572);
xnor UO_2357 (O_2357,N_23722,N_22825);
xnor UO_2358 (O_2358,N_22677,N_23107);
xnor UO_2359 (O_2359,N_24706,N_22134);
nor UO_2360 (O_2360,N_24172,N_22911);
nor UO_2361 (O_2361,N_24416,N_24298);
or UO_2362 (O_2362,N_23326,N_22834);
xnor UO_2363 (O_2363,N_23900,N_23588);
and UO_2364 (O_2364,N_23388,N_22787);
or UO_2365 (O_2365,N_22709,N_24667);
nor UO_2366 (O_2366,N_23468,N_24755);
nand UO_2367 (O_2367,N_22213,N_22339);
nand UO_2368 (O_2368,N_24943,N_22398);
nor UO_2369 (O_2369,N_22112,N_22624);
nor UO_2370 (O_2370,N_23095,N_23751);
or UO_2371 (O_2371,N_21902,N_22367);
and UO_2372 (O_2372,N_22954,N_24529);
or UO_2373 (O_2373,N_22950,N_22277);
xor UO_2374 (O_2374,N_24170,N_23649);
nor UO_2375 (O_2375,N_24427,N_23931);
xor UO_2376 (O_2376,N_22453,N_22737);
xnor UO_2377 (O_2377,N_23304,N_23585);
nor UO_2378 (O_2378,N_23287,N_22882);
xnor UO_2379 (O_2379,N_22659,N_22161);
nor UO_2380 (O_2380,N_22176,N_23295);
nor UO_2381 (O_2381,N_23387,N_22047);
and UO_2382 (O_2382,N_24083,N_24678);
and UO_2383 (O_2383,N_23946,N_22562);
or UO_2384 (O_2384,N_23842,N_22373);
xor UO_2385 (O_2385,N_23802,N_22475);
nor UO_2386 (O_2386,N_22945,N_24980);
nand UO_2387 (O_2387,N_22905,N_22541);
and UO_2388 (O_2388,N_24041,N_22964);
nor UO_2389 (O_2389,N_23058,N_23656);
nor UO_2390 (O_2390,N_23824,N_24570);
xor UO_2391 (O_2391,N_23096,N_23511);
nor UO_2392 (O_2392,N_22562,N_22537);
nand UO_2393 (O_2393,N_24673,N_24935);
nor UO_2394 (O_2394,N_24271,N_23124);
or UO_2395 (O_2395,N_23480,N_23792);
nor UO_2396 (O_2396,N_24480,N_21888);
nor UO_2397 (O_2397,N_24485,N_23137);
nand UO_2398 (O_2398,N_24561,N_23399);
xor UO_2399 (O_2399,N_22592,N_23205);
xor UO_2400 (O_2400,N_24185,N_23515);
and UO_2401 (O_2401,N_23553,N_22656);
xor UO_2402 (O_2402,N_23253,N_24604);
or UO_2403 (O_2403,N_23058,N_24262);
and UO_2404 (O_2404,N_23771,N_22420);
and UO_2405 (O_2405,N_24499,N_23832);
nor UO_2406 (O_2406,N_22088,N_22005);
xnor UO_2407 (O_2407,N_22162,N_23523);
xor UO_2408 (O_2408,N_23710,N_23041);
xor UO_2409 (O_2409,N_24605,N_23815);
or UO_2410 (O_2410,N_24903,N_22672);
xor UO_2411 (O_2411,N_22872,N_22615);
or UO_2412 (O_2412,N_23404,N_22360);
nor UO_2413 (O_2413,N_23695,N_24596);
or UO_2414 (O_2414,N_24657,N_23826);
xor UO_2415 (O_2415,N_22922,N_23023);
nor UO_2416 (O_2416,N_22010,N_24902);
and UO_2417 (O_2417,N_23260,N_24026);
nand UO_2418 (O_2418,N_24803,N_22559);
xor UO_2419 (O_2419,N_24527,N_22652);
or UO_2420 (O_2420,N_21976,N_22064);
xor UO_2421 (O_2421,N_24168,N_23532);
nand UO_2422 (O_2422,N_23611,N_24862);
or UO_2423 (O_2423,N_22508,N_24869);
xor UO_2424 (O_2424,N_23404,N_23883);
nor UO_2425 (O_2425,N_23652,N_23043);
and UO_2426 (O_2426,N_23914,N_21930);
and UO_2427 (O_2427,N_24669,N_22256);
xnor UO_2428 (O_2428,N_21918,N_22830);
and UO_2429 (O_2429,N_21981,N_23988);
and UO_2430 (O_2430,N_22820,N_22084);
nor UO_2431 (O_2431,N_22448,N_22167);
or UO_2432 (O_2432,N_22282,N_22217);
nand UO_2433 (O_2433,N_24528,N_24576);
xor UO_2434 (O_2434,N_23872,N_22767);
nand UO_2435 (O_2435,N_23328,N_21936);
nor UO_2436 (O_2436,N_24456,N_24892);
nor UO_2437 (O_2437,N_24877,N_22066);
and UO_2438 (O_2438,N_21919,N_23580);
or UO_2439 (O_2439,N_23652,N_22548);
nor UO_2440 (O_2440,N_22532,N_24435);
and UO_2441 (O_2441,N_22493,N_24275);
nor UO_2442 (O_2442,N_24395,N_23333);
or UO_2443 (O_2443,N_24998,N_24925);
nor UO_2444 (O_2444,N_22763,N_24127);
xnor UO_2445 (O_2445,N_23557,N_22726);
nand UO_2446 (O_2446,N_24810,N_22795);
xor UO_2447 (O_2447,N_24325,N_22874);
or UO_2448 (O_2448,N_24143,N_24969);
and UO_2449 (O_2449,N_22498,N_24451);
and UO_2450 (O_2450,N_24082,N_23662);
and UO_2451 (O_2451,N_23883,N_21914);
xnor UO_2452 (O_2452,N_23553,N_23941);
or UO_2453 (O_2453,N_23593,N_23653);
nor UO_2454 (O_2454,N_24045,N_22379);
xor UO_2455 (O_2455,N_24693,N_23304);
and UO_2456 (O_2456,N_24585,N_23036);
nor UO_2457 (O_2457,N_24427,N_22496);
nand UO_2458 (O_2458,N_21931,N_22452);
nor UO_2459 (O_2459,N_24320,N_24300);
or UO_2460 (O_2460,N_24404,N_24628);
xor UO_2461 (O_2461,N_22538,N_24838);
or UO_2462 (O_2462,N_24695,N_23098);
or UO_2463 (O_2463,N_24971,N_24377);
nand UO_2464 (O_2464,N_22635,N_24272);
xor UO_2465 (O_2465,N_22336,N_24572);
nor UO_2466 (O_2466,N_22401,N_24907);
xnor UO_2467 (O_2467,N_23429,N_23745);
nand UO_2468 (O_2468,N_23134,N_24942);
and UO_2469 (O_2469,N_23420,N_23760);
xor UO_2470 (O_2470,N_23590,N_24386);
xnor UO_2471 (O_2471,N_22333,N_24598);
or UO_2472 (O_2472,N_23412,N_24139);
xnor UO_2473 (O_2473,N_22667,N_22822);
xor UO_2474 (O_2474,N_22980,N_22617);
xnor UO_2475 (O_2475,N_24989,N_23231);
nor UO_2476 (O_2476,N_23281,N_22299);
nand UO_2477 (O_2477,N_23081,N_24692);
and UO_2478 (O_2478,N_22277,N_24469);
xnor UO_2479 (O_2479,N_24277,N_23354);
or UO_2480 (O_2480,N_24885,N_22122);
and UO_2481 (O_2481,N_23159,N_23281);
and UO_2482 (O_2482,N_24285,N_22505);
nor UO_2483 (O_2483,N_23329,N_23047);
and UO_2484 (O_2484,N_24467,N_24208);
nand UO_2485 (O_2485,N_22277,N_21966);
xnor UO_2486 (O_2486,N_21961,N_23313);
nand UO_2487 (O_2487,N_21900,N_22595);
and UO_2488 (O_2488,N_24273,N_22196);
nand UO_2489 (O_2489,N_23551,N_22251);
or UO_2490 (O_2490,N_24649,N_23539);
or UO_2491 (O_2491,N_22784,N_24314);
or UO_2492 (O_2492,N_24638,N_21906);
nor UO_2493 (O_2493,N_22944,N_23133);
xnor UO_2494 (O_2494,N_24752,N_23657);
xor UO_2495 (O_2495,N_22536,N_22127);
nand UO_2496 (O_2496,N_23052,N_24280);
or UO_2497 (O_2497,N_22264,N_24955);
nor UO_2498 (O_2498,N_22755,N_24702);
xor UO_2499 (O_2499,N_22097,N_22575);
or UO_2500 (O_2500,N_23795,N_23281);
or UO_2501 (O_2501,N_24587,N_22635);
or UO_2502 (O_2502,N_23415,N_23059);
xnor UO_2503 (O_2503,N_22326,N_24013);
nand UO_2504 (O_2504,N_23457,N_22943);
and UO_2505 (O_2505,N_22858,N_24078);
or UO_2506 (O_2506,N_22141,N_24464);
nor UO_2507 (O_2507,N_23756,N_22909);
nor UO_2508 (O_2508,N_24916,N_22883);
and UO_2509 (O_2509,N_22952,N_24909);
xor UO_2510 (O_2510,N_24734,N_23348);
or UO_2511 (O_2511,N_24991,N_23581);
and UO_2512 (O_2512,N_22716,N_23359);
nand UO_2513 (O_2513,N_24134,N_23755);
or UO_2514 (O_2514,N_24330,N_23361);
or UO_2515 (O_2515,N_21898,N_22207);
and UO_2516 (O_2516,N_23035,N_22972);
or UO_2517 (O_2517,N_22267,N_23416);
and UO_2518 (O_2518,N_22679,N_24839);
nor UO_2519 (O_2519,N_22719,N_22730);
and UO_2520 (O_2520,N_22758,N_24507);
and UO_2521 (O_2521,N_23524,N_22251);
or UO_2522 (O_2522,N_23276,N_22375);
nand UO_2523 (O_2523,N_24741,N_24210);
nand UO_2524 (O_2524,N_23874,N_23110);
nand UO_2525 (O_2525,N_24969,N_24109);
and UO_2526 (O_2526,N_23856,N_22797);
and UO_2527 (O_2527,N_22533,N_22906);
xnor UO_2528 (O_2528,N_24785,N_24181);
nand UO_2529 (O_2529,N_24008,N_24537);
or UO_2530 (O_2530,N_24196,N_23666);
nor UO_2531 (O_2531,N_22198,N_24874);
xor UO_2532 (O_2532,N_21911,N_24455);
nand UO_2533 (O_2533,N_24552,N_23887);
or UO_2534 (O_2534,N_22273,N_23696);
or UO_2535 (O_2535,N_23852,N_22404);
nand UO_2536 (O_2536,N_24294,N_23113);
nor UO_2537 (O_2537,N_24247,N_24447);
nor UO_2538 (O_2538,N_23973,N_23246);
nand UO_2539 (O_2539,N_24996,N_23875);
nor UO_2540 (O_2540,N_23010,N_24500);
and UO_2541 (O_2541,N_23555,N_23212);
nand UO_2542 (O_2542,N_24972,N_22866);
and UO_2543 (O_2543,N_23031,N_22127);
and UO_2544 (O_2544,N_22756,N_24757);
or UO_2545 (O_2545,N_24049,N_24403);
or UO_2546 (O_2546,N_24203,N_22884);
nor UO_2547 (O_2547,N_22857,N_23666);
xor UO_2548 (O_2548,N_21991,N_23907);
nand UO_2549 (O_2549,N_23407,N_24218);
or UO_2550 (O_2550,N_23362,N_22233);
nand UO_2551 (O_2551,N_23344,N_24287);
nand UO_2552 (O_2552,N_22892,N_24570);
nor UO_2553 (O_2553,N_24054,N_23068);
or UO_2554 (O_2554,N_23097,N_24131);
or UO_2555 (O_2555,N_22122,N_22531);
xor UO_2556 (O_2556,N_22661,N_22156);
nor UO_2557 (O_2557,N_24361,N_22179);
xnor UO_2558 (O_2558,N_22513,N_22806);
nand UO_2559 (O_2559,N_22694,N_22949);
xnor UO_2560 (O_2560,N_23490,N_23246);
xor UO_2561 (O_2561,N_23910,N_22941);
nor UO_2562 (O_2562,N_22766,N_24242);
and UO_2563 (O_2563,N_22961,N_24464);
or UO_2564 (O_2564,N_22000,N_23873);
xor UO_2565 (O_2565,N_23356,N_22831);
and UO_2566 (O_2566,N_22040,N_23817);
xor UO_2567 (O_2567,N_22012,N_22839);
or UO_2568 (O_2568,N_24975,N_23592);
xor UO_2569 (O_2569,N_23375,N_23468);
nor UO_2570 (O_2570,N_23348,N_23516);
nor UO_2571 (O_2571,N_23220,N_24561);
nor UO_2572 (O_2572,N_22555,N_21964);
nor UO_2573 (O_2573,N_24541,N_24434);
nor UO_2574 (O_2574,N_23700,N_23254);
or UO_2575 (O_2575,N_22770,N_24291);
nor UO_2576 (O_2576,N_22736,N_24045);
xor UO_2577 (O_2577,N_24166,N_22870);
xor UO_2578 (O_2578,N_23268,N_22452);
and UO_2579 (O_2579,N_24677,N_24783);
nor UO_2580 (O_2580,N_22227,N_22904);
nor UO_2581 (O_2581,N_22785,N_23531);
xnor UO_2582 (O_2582,N_24079,N_22833);
nor UO_2583 (O_2583,N_24047,N_24050);
and UO_2584 (O_2584,N_23054,N_24200);
nand UO_2585 (O_2585,N_23240,N_24530);
nand UO_2586 (O_2586,N_23371,N_22667);
xor UO_2587 (O_2587,N_22896,N_23964);
xor UO_2588 (O_2588,N_22022,N_24228);
and UO_2589 (O_2589,N_22601,N_22299);
or UO_2590 (O_2590,N_23638,N_23645);
xor UO_2591 (O_2591,N_24672,N_23613);
nand UO_2592 (O_2592,N_23850,N_24321);
nor UO_2593 (O_2593,N_24725,N_24853);
xnor UO_2594 (O_2594,N_23508,N_23853);
or UO_2595 (O_2595,N_23119,N_24646);
or UO_2596 (O_2596,N_24737,N_24684);
xnor UO_2597 (O_2597,N_22546,N_23667);
nand UO_2598 (O_2598,N_22725,N_23618);
or UO_2599 (O_2599,N_22243,N_21998);
nor UO_2600 (O_2600,N_22606,N_23093);
and UO_2601 (O_2601,N_23329,N_22740);
xnor UO_2602 (O_2602,N_24524,N_23471);
and UO_2603 (O_2603,N_22295,N_22108);
xnor UO_2604 (O_2604,N_23352,N_22428);
or UO_2605 (O_2605,N_24869,N_22650);
nor UO_2606 (O_2606,N_23172,N_23397);
nand UO_2607 (O_2607,N_23811,N_24088);
nand UO_2608 (O_2608,N_21919,N_23397);
nor UO_2609 (O_2609,N_23696,N_23816);
xor UO_2610 (O_2610,N_22706,N_24246);
or UO_2611 (O_2611,N_22616,N_21913);
nand UO_2612 (O_2612,N_23060,N_24025);
or UO_2613 (O_2613,N_24853,N_22811);
and UO_2614 (O_2614,N_23161,N_22092);
or UO_2615 (O_2615,N_23012,N_23497);
and UO_2616 (O_2616,N_23610,N_23488);
nor UO_2617 (O_2617,N_22972,N_23185);
nand UO_2618 (O_2618,N_23246,N_24474);
or UO_2619 (O_2619,N_23810,N_24472);
or UO_2620 (O_2620,N_22670,N_23207);
or UO_2621 (O_2621,N_22949,N_23706);
or UO_2622 (O_2622,N_23514,N_24000);
xor UO_2623 (O_2623,N_24906,N_22499);
nor UO_2624 (O_2624,N_24560,N_23048);
or UO_2625 (O_2625,N_23739,N_22335);
nor UO_2626 (O_2626,N_22357,N_23341);
and UO_2627 (O_2627,N_22325,N_23636);
or UO_2628 (O_2628,N_22871,N_24121);
nand UO_2629 (O_2629,N_23235,N_22814);
nand UO_2630 (O_2630,N_22285,N_23533);
nor UO_2631 (O_2631,N_23160,N_23115);
and UO_2632 (O_2632,N_23831,N_23261);
xor UO_2633 (O_2633,N_24799,N_24697);
or UO_2634 (O_2634,N_22377,N_24674);
and UO_2635 (O_2635,N_22207,N_22084);
xnor UO_2636 (O_2636,N_24864,N_24568);
and UO_2637 (O_2637,N_22540,N_22252);
xor UO_2638 (O_2638,N_22857,N_24686);
nor UO_2639 (O_2639,N_24787,N_24103);
nor UO_2640 (O_2640,N_23395,N_22137);
and UO_2641 (O_2641,N_21887,N_21877);
nor UO_2642 (O_2642,N_24716,N_24928);
and UO_2643 (O_2643,N_22966,N_22181);
and UO_2644 (O_2644,N_22402,N_22684);
and UO_2645 (O_2645,N_22254,N_23833);
nor UO_2646 (O_2646,N_22383,N_23003);
nor UO_2647 (O_2647,N_23723,N_24458);
and UO_2648 (O_2648,N_21940,N_24810);
nand UO_2649 (O_2649,N_23856,N_24948);
nor UO_2650 (O_2650,N_22629,N_23019);
or UO_2651 (O_2651,N_23664,N_22855);
xnor UO_2652 (O_2652,N_22107,N_24143);
or UO_2653 (O_2653,N_22527,N_22884);
xnor UO_2654 (O_2654,N_22951,N_23095);
nor UO_2655 (O_2655,N_22082,N_23281);
and UO_2656 (O_2656,N_22265,N_22814);
nand UO_2657 (O_2657,N_24371,N_24281);
and UO_2658 (O_2658,N_24913,N_21901);
xor UO_2659 (O_2659,N_23341,N_22080);
nor UO_2660 (O_2660,N_23992,N_24026);
nand UO_2661 (O_2661,N_24562,N_22505);
nand UO_2662 (O_2662,N_23947,N_23434);
and UO_2663 (O_2663,N_23797,N_23028);
xor UO_2664 (O_2664,N_23357,N_22103);
or UO_2665 (O_2665,N_23109,N_23702);
nor UO_2666 (O_2666,N_22930,N_22450);
nor UO_2667 (O_2667,N_23691,N_24540);
and UO_2668 (O_2668,N_23807,N_22151);
or UO_2669 (O_2669,N_23194,N_24735);
or UO_2670 (O_2670,N_22798,N_24520);
nand UO_2671 (O_2671,N_23147,N_21880);
nor UO_2672 (O_2672,N_24279,N_24665);
nor UO_2673 (O_2673,N_24229,N_22960);
and UO_2674 (O_2674,N_22848,N_24381);
nand UO_2675 (O_2675,N_22467,N_23727);
and UO_2676 (O_2676,N_24939,N_23397);
nand UO_2677 (O_2677,N_23868,N_24817);
xnor UO_2678 (O_2678,N_24585,N_23961);
or UO_2679 (O_2679,N_23063,N_21965);
nor UO_2680 (O_2680,N_23289,N_22274);
or UO_2681 (O_2681,N_24151,N_21876);
nor UO_2682 (O_2682,N_23535,N_24963);
nor UO_2683 (O_2683,N_23807,N_22774);
and UO_2684 (O_2684,N_22121,N_24127);
and UO_2685 (O_2685,N_22114,N_24015);
or UO_2686 (O_2686,N_22220,N_23167);
nor UO_2687 (O_2687,N_24725,N_22412);
xnor UO_2688 (O_2688,N_23358,N_24267);
nor UO_2689 (O_2689,N_24583,N_23524);
or UO_2690 (O_2690,N_23537,N_24906);
nor UO_2691 (O_2691,N_23088,N_23182);
xnor UO_2692 (O_2692,N_23294,N_22422);
xnor UO_2693 (O_2693,N_23851,N_23969);
and UO_2694 (O_2694,N_23471,N_23815);
nand UO_2695 (O_2695,N_22675,N_24328);
xor UO_2696 (O_2696,N_24969,N_23910);
or UO_2697 (O_2697,N_24254,N_24656);
nand UO_2698 (O_2698,N_22399,N_22694);
or UO_2699 (O_2699,N_21996,N_22624);
and UO_2700 (O_2700,N_22089,N_22736);
or UO_2701 (O_2701,N_24629,N_23640);
xor UO_2702 (O_2702,N_22307,N_24223);
xor UO_2703 (O_2703,N_24051,N_23761);
and UO_2704 (O_2704,N_24515,N_23591);
or UO_2705 (O_2705,N_24233,N_24415);
nor UO_2706 (O_2706,N_23871,N_22091);
xnor UO_2707 (O_2707,N_24543,N_23826);
xor UO_2708 (O_2708,N_24350,N_24660);
xor UO_2709 (O_2709,N_22294,N_24848);
nor UO_2710 (O_2710,N_23382,N_24626);
xnor UO_2711 (O_2711,N_22924,N_24996);
or UO_2712 (O_2712,N_22336,N_24372);
nand UO_2713 (O_2713,N_23460,N_23807);
xnor UO_2714 (O_2714,N_24014,N_23093);
nor UO_2715 (O_2715,N_23582,N_23418);
and UO_2716 (O_2716,N_23103,N_23181);
and UO_2717 (O_2717,N_24877,N_23670);
xnor UO_2718 (O_2718,N_24810,N_23589);
nor UO_2719 (O_2719,N_22465,N_23788);
and UO_2720 (O_2720,N_22157,N_23967);
nor UO_2721 (O_2721,N_23347,N_22515);
nand UO_2722 (O_2722,N_22573,N_22807);
xor UO_2723 (O_2723,N_22049,N_24462);
or UO_2724 (O_2724,N_22830,N_24567);
and UO_2725 (O_2725,N_22953,N_22482);
or UO_2726 (O_2726,N_24983,N_22133);
and UO_2727 (O_2727,N_22599,N_23201);
xnor UO_2728 (O_2728,N_24044,N_22404);
nand UO_2729 (O_2729,N_24262,N_21878);
or UO_2730 (O_2730,N_23329,N_23871);
nor UO_2731 (O_2731,N_22633,N_22736);
or UO_2732 (O_2732,N_21878,N_23452);
nor UO_2733 (O_2733,N_22779,N_24656);
nand UO_2734 (O_2734,N_22988,N_22001);
and UO_2735 (O_2735,N_24886,N_24262);
and UO_2736 (O_2736,N_23722,N_24019);
and UO_2737 (O_2737,N_23103,N_23117);
nand UO_2738 (O_2738,N_23956,N_24981);
or UO_2739 (O_2739,N_23623,N_23777);
xor UO_2740 (O_2740,N_23135,N_23492);
nor UO_2741 (O_2741,N_22478,N_22329);
or UO_2742 (O_2742,N_23260,N_22253);
and UO_2743 (O_2743,N_23748,N_23022);
or UO_2744 (O_2744,N_22588,N_23489);
and UO_2745 (O_2745,N_22703,N_24227);
or UO_2746 (O_2746,N_23220,N_24485);
nand UO_2747 (O_2747,N_22383,N_22739);
nor UO_2748 (O_2748,N_22048,N_24352);
nor UO_2749 (O_2749,N_24938,N_24529);
nand UO_2750 (O_2750,N_23032,N_24043);
nor UO_2751 (O_2751,N_23514,N_23978);
nor UO_2752 (O_2752,N_22892,N_22786);
or UO_2753 (O_2753,N_24520,N_24550);
and UO_2754 (O_2754,N_23837,N_22527);
or UO_2755 (O_2755,N_24174,N_24077);
nor UO_2756 (O_2756,N_22240,N_22161);
and UO_2757 (O_2757,N_21983,N_23938);
nand UO_2758 (O_2758,N_24215,N_23782);
and UO_2759 (O_2759,N_23563,N_24441);
nand UO_2760 (O_2760,N_24344,N_22532);
or UO_2761 (O_2761,N_24172,N_22034);
nand UO_2762 (O_2762,N_24624,N_23560);
or UO_2763 (O_2763,N_24401,N_23953);
xor UO_2764 (O_2764,N_24759,N_24336);
xnor UO_2765 (O_2765,N_23682,N_22944);
nor UO_2766 (O_2766,N_22040,N_24307);
nor UO_2767 (O_2767,N_23960,N_22545);
nor UO_2768 (O_2768,N_22148,N_23212);
nor UO_2769 (O_2769,N_24947,N_23532);
and UO_2770 (O_2770,N_22247,N_23649);
nor UO_2771 (O_2771,N_21904,N_23807);
nor UO_2772 (O_2772,N_22656,N_24142);
and UO_2773 (O_2773,N_24655,N_24393);
and UO_2774 (O_2774,N_23997,N_22668);
nor UO_2775 (O_2775,N_23532,N_23477);
nor UO_2776 (O_2776,N_21944,N_22643);
or UO_2777 (O_2777,N_23423,N_24438);
xor UO_2778 (O_2778,N_23139,N_22589);
nand UO_2779 (O_2779,N_24580,N_22408);
nand UO_2780 (O_2780,N_22013,N_24244);
xor UO_2781 (O_2781,N_24290,N_22059);
nand UO_2782 (O_2782,N_22384,N_22482);
nand UO_2783 (O_2783,N_23437,N_23917);
and UO_2784 (O_2784,N_24276,N_24362);
xor UO_2785 (O_2785,N_22756,N_23394);
xor UO_2786 (O_2786,N_24957,N_23464);
xnor UO_2787 (O_2787,N_23865,N_21925);
and UO_2788 (O_2788,N_21957,N_24373);
or UO_2789 (O_2789,N_23430,N_22281);
xor UO_2790 (O_2790,N_23726,N_23279);
nand UO_2791 (O_2791,N_22273,N_22678);
nand UO_2792 (O_2792,N_24696,N_24060);
nor UO_2793 (O_2793,N_23287,N_22225);
xor UO_2794 (O_2794,N_22925,N_24698);
or UO_2795 (O_2795,N_23856,N_22396);
or UO_2796 (O_2796,N_24632,N_23583);
nor UO_2797 (O_2797,N_21975,N_24232);
xor UO_2798 (O_2798,N_22252,N_22352);
nor UO_2799 (O_2799,N_24128,N_23586);
xnor UO_2800 (O_2800,N_23209,N_24296);
nor UO_2801 (O_2801,N_24569,N_22397);
nor UO_2802 (O_2802,N_24939,N_22657);
or UO_2803 (O_2803,N_22983,N_24210);
and UO_2804 (O_2804,N_24227,N_23245);
nor UO_2805 (O_2805,N_22617,N_24636);
nor UO_2806 (O_2806,N_23978,N_22374);
xnor UO_2807 (O_2807,N_24044,N_24379);
nor UO_2808 (O_2808,N_22810,N_23461);
or UO_2809 (O_2809,N_23428,N_23617);
nor UO_2810 (O_2810,N_24018,N_22110);
and UO_2811 (O_2811,N_22741,N_23069);
nand UO_2812 (O_2812,N_24386,N_22645);
nand UO_2813 (O_2813,N_23126,N_24213);
or UO_2814 (O_2814,N_22914,N_22182);
xnor UO_2815 (O_2815,N_21934,N_24702);
and UO_2816 (O_2816,N_24106,N_22691);
and UO_2817 (O_2817,N_22753,N_24216);
and UO_2818 (O_2818,N_22539,N_22386);
or UO_2819 (O_2819,N_24053,N_22300);
nand UO_2820 (O_2820,N_24429,N_22223);
xnor UO_2821 (O_2821,N_24538,N_24889);
or UO_2822 (O_2822,N_23306,N_23182);
nand UO_2823 (O_2823,N_22449,N_24606);
or UO_2824 (O_2824,N_22132,N_22655);
nor UO_2825 (O_2825,N_22057,N_24252);
or UO_2826 (O_2826,N_22089,N_23797);
xnor UO_2827 (O_2827,N_22264,N_23721);
and UO_2828 (O_2828,N_23390,N_22914);
nand UO_2829 (O_2829,N_22704,N_23058);
nand UO_2830 (O_2830,N_24040,N_24685);
nand UO_2831 (O_2831,N_22535,N_24352);
or UO_2832 (O_2832,N_24947,N_24292);
and UO_2833 (O_2833,N_22363,N_22629);
nand UO_2834 (O_2834,N_23060,N_24084);
or UO_2835 (O_2835,N_22934,N_24797);
nor UO_2836 (O_2836,N_22118,N_23147);
xor UO_2837 (O_2837,N_24764,N_23232);
nor UO_2838 (O_2838,N_23465,N_24224);
and UO_2839 (O_2839,N_22030,N_23938);
nand UO_2840 (O_2840,N_23478,N_22548);
and UO_2841 (O_2841,N_22581,N_22156);
and UO_2842 (O_2842,N_22774,N_23938);
nand UO_2843 (O_2843,N_22444,N_22092);
or UO_2844 (O_2844,N_22491,N_24965);
nand UO_2845 (O_2845,N_24938,N_22619);
xor UO_2846 (O_2846,N_24298,N_22346);
or UO_2847 (O_2847,N_24945,N_23845);
nor UO_2848 (O_2848,N_22715,N_23222);
and UO_2849 (O_2849,N_24886,N_22707);
xnor UO_2850 (O_2850,N_23628,N_23638);
and UO_2851 (O_2851,N_23197,N_23725);
and UO_2852 (O_2852,N_23008,N_23261);
or UO_2853 (O_2853,N_24636,N_22651);
or UO_2854 (O_2854,N_24251,N_22770);
nand UO_2855 (O_2855,N_24407,N_22179);
or UO_2856 (O_2856,N_23891,N_24617);
or UO_2857 (O_2857,N_21910,N_22913);
or UO_2858 (O_2858,N_22601,N_24093);
or UO_2859 (O_2859,N_24923,N_24610);
nand UO_2860 (O_2860,N_23779,N_22600);
nor UO_2861 (O_2861,N_23393,N_22815);
nor UO_2862 (O_2862,N_24834,N_24813);
and UO_2863 (O_2863,N_24322,N_24027);
nand UO_2864 (O_2864,N_23894,N_24624);
xor UO_2865 (O_2865,N_24189,N_23438);
or UO_2866 (O_2866,N_24625,N_22301);
nor UO_2867 (O_2867,N_24914,N_23983);
or UO_2868 (O_2868,N_24726,N_22687);
xnor UO_2869 (O_2869,N_22961,N_21979);
or UO_2870 (O_2870,N_22245,N_23242);
or UO_2871 (O_2871,N_22363,N_22228);
xor UO_2872 (O_2872,N_23862,N_24592);
xor UO_2873 (O_2873,N_24028,N_22738);
or UO_2874 (O_2874,N_21946,N_22768);
nand UO_2875 (O_2875,N_22323,N_22943);
or UO_2876 (O_2876,N_23971,N_22772);
nor UO_2877 (O_2877,N_24489,N_22950);
and UO_2878 (O_2878,N_22670,N_23679);
xnor UO_2879 (O_2879,N_24682,N_23994);
nand UO_2880 (O_2880,N_23217,N_22855);
nand UO_2881 (O_2881,N_21933,N_22334);
xnor UO_2882 (O_2882,N_22001,N_24845);
nor UO_2883 (O_2883,N_23366,N_23669);
xnor UO_2884 (O_2884,N_24852,N_23226);
and UO_2885 (O_2885,N_23398,N_22477);
or UO_2886 (O_2886,N_22503,N_22134);
nand UO_2887 (O_2887,N_22003,N_24302);
or UO_2888 (O_2888,N_24448,N_24902);
nor UO_2889 (O_2889,N_23229,N_24665);
nor UO_2890 (O_2890,N_24583,N_22829);
or UO_2891 (O_2891,N_23827,N_23439);
xor UO_2892 (O_2892,N_24706,N_24730);
nor UO_2893 (O_2893,N_22154,N_22789);
xor UO_2894 (O_2894,N_23802,N_24737);
nand UO_2895 (O_2895,N_24191,N_23488);
or UO_2896 (O_2896,N_24477,N_24959);
nand UO_2897 (O_2897,N_22677,N_22973);
and UO_2898 (O_2898,N_22559,N_21996);
nand UO_2899 (O_2899,N_22540,N_23484);
or UO_2900 (O_2900,N_24782,N_23407);
or UO_2901 (O_2901,N_23082,N_24831);
nand UO_2902 (O_2902,N_24320,N_22883);
nor UO_2903 (O_2903,N_23670,N_24633);
or UO_2904 (O_2904,N_24836,N_22918);
xor UO_2905 (O_2905,N_23524,N_23547);
and UO_2906 (O_2906,N_23411,N_23302);
xor UO_2907 (O_2907,N_23238,N_24363);
or UO_2908 (O_2908,N_24814,N_23447);
nand UO_2909 (O_2909,N_24664,N_23527);
and UO_2910 (O_2910,N_24371,N_24116);
or UO_2911 (O_2911,N_24116,N_23536);
xnor UO_2912 (O_2912,N_22358,N_23140);
xor UO_2913 (O_2913,N_24444,N_23791);
and UO_2914 (O_2914,N_23777,N_22093);
or UO_2915 (O_2915,N_22952,N_22157);
nor UO_2916 (O_2916,N_22671,N_24163);
or UO_2917 (O_2917,N_23010,N_22058);
nand UO_2918 (O_2918,N_23029,N_24664);
and UO_2919 (O_2919,N_23160,N_22040);
nor UO_2920 (O_2920,N_23855,N_22862);
nor UO_2921 (O_2921,N_22126,N_22300);
nor UO_2922 (O_2922,N_23057,N_23437);
and UO_2923 (O_2923,N_23687,N_24817);
nor UO_2924 (O_2924,N_22612,N_21894);
or UO_2925 (O_2925,N_22950,N_22982);
nand UO_2926 (O_2926,N_22992,N_24644);
and UO_2927 (O_2927,N_23968,N_24920);
nor UO_2928 (O_2928,N_24798,N_23353);
nor UO_2929 (O_2929,N_24403,N_23784);
nand UO_2930 (O_2930,N_22191,N_22580);
and UO_2931 (O_2931,N_22859,N_24724);
nor UO_2932 (O_2932,N_22705,N_24954);
nand UO_2933 (O_2933,N_23144,N_24699);
nand UO_2934 (O_2934,N_22924,N_22261);
xnor UO_2935 (O_2935,N_24044,N_23257);
xnor UO_2936 (O_2936,N_23039,N_23359);
or UO_2937 (O_2937,N_22359,N_23987);
and UO_2938 (O_2938,N_22193,N_22126);
and UO_2939 (O_2939,N_23097,N_23823);
xnor UO_2940 (O_2940,N_24044,N_24153);
and UO_2941 (O_2941,N_24321,N_22990);
xor UO_2942 (O_2942,N_23021,N_23857);
and UO_2943 (O_2943,N_24661,N_23620);
nor UO_2944 (O_2944,N_23214,N_24614);
nand UO_2945 (O_2945,N_23407,N_22861);
nand UO_2946 (O_2946,N_24430,N_22049);
nand UO_2947 (O_2947,N_22260,N_22274);
or UO_2948 (O_2948,N_22156,N_23030);
xor UO_2949 (O_2949,N_22266,N_24431);
nand UO_2950 (O_2950,N_24839,N_24167);
and UO_2951 (O_2951,N_24111,N_24421);
nor UO_2952 (O_2952,N_22878,N_24029);
or UO_2953 (O_2953,N_24627,N_22533);
xor UO_2954 (O_2954,N_23633,N_23196);
and UO_2955 (O_2955,N_22470,N_24608);
nand UO_2956 (O_2956,N_22106,N_23705);
and UO_2957 (O_2957,N_24586,N_22344);
and UO_2958 (O_2958,N_22177,N_22403);
and UO_2959 (O_2959,N_22168,N_24112);
or UO_2960 (O_2960,N_22522,N_22549);
and UO_2961 (O_2961,N_22415,N_24470);
xnor UO_2962 (O_2962,N_21967,N_23873);
or UO_2963 (O_2963,N_24142,N_23441);
nand UO_2964 (O_2964,N_22062,N_22306);
or UO_2965 (O_2965,N_24103,N_23414);
or UO_2966 (O_2966,N_22298,N_23221);
xor UO_2967 (O_2967,N_24810,N_23975);
xnor UO_2968 (O_2968,N_23706,N_24819);
nand UO_2969 (O_2969,N_24255,N_22164);
xnor UO_2970 (O_2970,N_22591,N_24527);
or UO_2971 (O_2971,N_24476,N_23187);
and UO_2972 (O_2972,N_22000,N_22369);
or UO_2973 (O_2973,N_22274,N_23716);
nor UO_2974 (O_2974,N_22515,N_22163);
nor UO_2975 (O_2975,N_22105,N_23137);
or UO_2976 (O_2976,N_22924,N_22506);
nor UO_2977 (O_2977,N_24219,N_22192);
nand UO_2978 (O_2978,N_23517,N_23916);
xor UO_2979 (O_2979,N_23242,N_22947);
or UO_2980 (O_2980,N_23046,N_23459);
or UO_2981 (O_2981,N_22232,N_22086);
and UO_2982 (O_2982,N_22463,N_24953);
nand UO_2983 (O_2983,N_23316,N_22869);
nor UO_2984 (O_2984,N_23626,N_23069);
nor UO_2985 (O_2985,N_21956,N_23206);
or UO_2986 (O_2986,N_22169,N_23399);
and UO_2987 (O_2987,N_24175,N_22039);
or UO_2988 (O_2988,N_22478,N_21991);
or UO_2989 (O_2989,N_23811,N_22538);
or UO_2990 (O_2990,N_23939,N_22538);
nand UO_2991 (O_2991,N_24178,N_24185);
xor UO_2992 (O_2992,N_23938,N_24738);
xor UO_2993 (O_2993,N_23444,N_22273);
nand UO_2994 (O_2994,N_22408,N_24828);
nand UO_2995 (O_2995,N_24332,N_23370);
xnor UO_2996 (O_2996,N_23455,N_24875);
nor UO_2997 (O_2997,N_24175,N_24036);
and UO_2998 (O_2998,N_24827,N_23826);
nor UO_2999 (O_2999,N_24227,N_23926);
endmodule