module basic_1000_10000_1500_50_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_265,In_410);
nand U1 (N_1,In_968,In_286);
nor U2 (N_2,In_485,In_693);
or U3 (N_3,In_345,In_582);
nand U4 (N_4,In_852,In_718);
nand U5 (N_5,In_184,In_720);
and U6 (N_6,In_525,In_200);
or U7 (N_7,In_935,In_608);
nor U8 (N_8,In_375,In_181);
nor U9 (N_9,In_120,In_289);
nand U10 (N_10,In_668,In_16);
and U11 (N_11,In_229,In_431);
and U12 (N_12,In_857,In_727);
or U13 (N_13,In_666,In_340);
and U14 (N_14,In_58,In_700);
nor U15 (N_15,In_712,In_356);
nor U16 (N_16,In_490,In_80);
or U17 (N_17,In_257,In_94);
nand U18 (N_18,In_263,In_391);
nor U19 (N_19,In_427,In_556);
nand U20 (N_20,In_237,In_385);
or U21 (N_21,In_282,In_602);
nor U22 (N_22,In_551,In_238);
and U23 (N_23,In_69,In_818);
nor U24 (N_24,In_805,In_692);
nand U25 (N_25,In_631,In_25);
and U26 (N_26,In_248,In_308);
nand U27 (N_27,In_285,In_126);
and U28 (N_28,In_507,In_275);
nand U29 (N_29,In_27,In_167);
or U30 (N_30,In_520,In_449);
nor U31 (N_31,In_847,In_998);
or U32 (N_32,In_813,In_611);
nand U33 (N_33,In_639,In_757);
nand U34 (N_34,In_500,In_158);
nor U35 (N_35,In_305,In_7);
or U36 (N_36,In_481,In_251);
nor U37 (N_37,In_130,In_258);
or U38 (N_38,In_399,In_785);
and U39 (N_39,In_961,In_11);
or U40 (N_40,In_203,In_766);
nand U41 (N_41,In_734,In_295);
nand U42 (N_42,In_91,In_176);
or U43 (N_43,In_966,In_657);
and U44 (N_44,In_676,In_661);
and U45 (N_45,In_883,In_597);
nor U46 (N_46,In_950,In_911);
and U47 (N_47,In_916,In_194);
and U48 (N_48,In_561,In_665);
or U49 (N_49,In_509,In_791);
or U50 (N_50,In_495,In_637);
or U51 (N_51,In_68,In_836);
or U52 (N_52,In_817,In_421);
nor U53 (N_53,In_952,In_922);
xor U54 (N_54,In_779,In_435);
nand U55 (N_55,In_843,In_686);
or U56 (N_56,In_749,In_359);
and U57 (N_57,In_18,In_706);
nor U58 (N_58,In_644,In_521);
nand U59 (N_59,In_863,In_554);
and U60 (N_60,In_636,In_302);
nor U61 (N_61,In_654,In_951);
and U62 (N_62,In_400,In_216);
or U63 (N_63,In_423,In_211);
nand U64 (N_64,In_862,In_990);
or U65 (N_65,In_771,In_47);
nor U66 (N_66,In_957,In_136);
and U67 (N_67,In_792,In_955);
nand U68 (N_68,In_812,In_746);
nand U69 (N_69,In_220,In_317);
nor U70 (N_70,In_536,In_867);
xnor U71 (N_71,In_174,In_103);
nand U72 (N_72,In_591,In_336);
and U73 (N_73,In_568,In_988);
or U74 (N_74,In_616,In_938);
and U75 (N_75,In_982,In_772);
or U76 (N_76,In_747,In_563);
or U77 (N_77,In_182,In_972);
nand U78 (N_78,In_905,In_230);
and U79 (N_79,In_815,In_439);
nand U80 (N_80,In_801,In_104);
and U81 (N_81,In_398,In_774);
or U82 (N_82,In_992,In_527);
or U83 (N_83,In_458,In_963);
nor U84 (N_84,In_226,In_477);
or U85 (N_85,In_309,In_729);
nor U86 (N_86,In_735,In_235);
or U87 (N_87,In_869,In_380);
and U88 (N_88,In_41,In_778);
or U89 (N_89,In_594,In_113);
nor U90 (N_90,In_151,In_111);
or U91 (N_91,In_853,In_583);
or U92 (N_92,In_733,In_546);
nor U93 (N_93,In_386,In_150);
or U94 (N_94,In_180,In_555);
xnor U95 (N_95,In_986,In_259);
and U96 (N_96,In_910,In_267);
nand U97 (N_97,In_190,In_760);
or U98 (N_98,In_981,In_378);
or U99 (N_99,In_848,In_252);
nand U100 (N_100,In_465,In_417);
nand U101 (N_101,In_924,In_13);
nand U102 (N_102,In_985,In_586);
and U103 (N_103,In_165,In_467);
nor U104 (N_104,In_511,In_626);
nand U105 (N_105,In_73,In_839);
nand U106 (N_106,In_761,In_728);
nand U107 (N_107,In_365,In_669);
nand U108 (N_108,In_680,In_156);
xor U109 (N_109,In_708,In_962);
or U110 (N_110,In_830,In_494);
or U111 (N_111,In_379,In_393);
nand U112 (N_112,In_914,In_559);
or U113 (N_113,In_756,In_217);
nor U114 (N_114,In_307,In_428);
and U115 (N_115,In_195,In_925);
or U116 (N_116,In_4,In_339);
or U117 (N_117,In_810,In_675);
nor U118 (N_118,In_371,In_19);
nand U119 (N_119,In_625,In_939);
nand U120 (N_120,In_662,In_519);
and U121 (N_121,In_983,In_711);
nand U122 (N_122,In_683,In_247);
nor U123 (N_123,In_321,In_60);
or U124 (N_124,In_102,In_415);
nor U125 (N_125,In_806,In_108);
nand U126 (N_126,In_530,In_553);
and U127 (N_127,In_945,In_456);
or U128 (N_128,In_717,In_407);
and U129 (N_129,In_638,In_516);
and U130 (N_130,In_976,In_890);
or U131 (N_131,In_278,In_442);
or U132 (N_132,In_763,In_508);
nor U133 (N_133,In_991,In_946);
nand U134 (N_134,In_587,In_658);
and U135 (N_135,In_893,In_566);
or U136 (N_136,In_34,In_441);
or U137 (N_137,In_45,In_462);
and U138 (N_138,In_739,In_802);
and U139 (N_139,In_725,In_560);
and U140 (N_140,In_172,In_383);
or U141 (N_141,In_470,In_189);
nand U142 (N_142,In_798,In_506);
nand U143 (N_143,In_213,In_118);
and U144 (N_144,In_876,In_463);
xor U145 (N_145,In_8,In_777);
xnor U146 (N_146,In_532,In_138);
or U147 (N_147,In_851,In_592);
and U148 (N_148,In_613,In_89);
nor U149 (N_149,In_87,In_472);
nor U150 (N_150,In_811,In_129);
or U151 (N_151,In_672,In_759);
nand U152 (N_152,In_628,In_92);
and U153 (N_153,In_589,In_653);
nor U154 (N_154,In_845,In_394);
nand U155 (N_155,In_748,In_833);
nand U156 (N_156,In_565,In_361);
nand U157 (N_157,In_534,In_970);
or U158 (N_158,In_856,In_457);
and U159 (N_159,In_884,In_943);
and U160 (N_160,In_166,In_816);
and U161 (N_161,In_178,In_20);
nand U162 (N_162,In_9,In_24);
nor U163 (N_163,In_350,In_231);
or U164 (N_164,In_842,In_736);
nor U165 (N_165,In_603,In_898);
nand U166 (N_166,In_599,In_871);
and U167 (N_167,In_438,In_796);
nor U168 (N_168,In_29,In_934);
and U169 (N_169,In_996,In_742);
nor U170 (N_170,In_635,In_335);
and U171 (N_171,In_809,In_406);
and U172 (N_172,In_897,In_93);
nand U173 (N_173,In_786,In_142);
xnor U174 (N_174,In_242,In_948);
nor U175 (N_175,In_436,In_59);
nor U176 (N_176,In_496,In_177);
nor U177 (N_177,In_510,In_368);
and U178 (N_178,In_429,In_139);
nand U179 (N_179,In_243,In_980);
and U180 (N_180,In_425,In_12);
nor U181 (N_181,In_959,In_38);
or U182 (N_182,In_873,In_146);
nand U183 (N_183,In_926,In_362);
nor U184 (N_184,In_899,In_67);
and U185 (N_185,In_670,In_419);
or U186 (N_186,In_402,In_620);
nand U187 (N_187,In_54,In_570);
nor U188 (N_188,In_186,In_524);
or U189 (N_189,In_901,In_491);
or U190 (N_190,In_206,In_701);
nand U191 (N_191,In_74,In_426);
or U192 (N_192,In_0,In_77);
nand U193 (N_193,In_316,In_170);
and U194 (N_194,In_900,In_753);
nand U195 (N_195,In_420,In_413);
and U196 (N_196,In_659,In_674);
nand U197 (N_197,In_831,In_794);
nor U198 (N_198,In_598,In_78);
nor U199 (N_199,In_502,In_124);
nand U200 (N_200,In_100,In_412);
and U201 (N_201,N_70,In_523);
and U202 (N_202,In_72,In_175);
nand U203 (N_203,In_82,In_55);
nand U204 (N_204,In_121,In_197);
nor U205 (N_205,In_341,N_10);
nor U206 (N_206,In_478,In_453);
nand U207 (N_207,In_714,N_109);
nand U208 (N_208,In_304,In_334);
nand U209 (N_209,In_125,In_515);
and U210 (N_210,In_906,N_12);
and U211 (N_211,In_106,In_609);
nand U212 (N_212,In_548,N_118);
nand U213 (N_213,In_40,In_593);
nor U214 (N_214,In_770,In_253);
nor U215 (N_215,In_223,N_106);
or U216 (N_216,In_214,N_169);
or U217 (N_217,N_103,In_488);
nand U218 (N_218,N_51,In_758);
and U219 (N_219,N_191,N_72);
and U220 (N_220,N_89,N_102);
and U221 (N_221,In_141,In_21);
or U222 (N_222,In_671,In_244);
and U223 (N_223,In_128,N_138);
or U224 (N_224,N_38,In_347);
or U225 (N_225,In_787,N_88);
and U226 (N_226,In_221,In_315);
nor U227 (N_227,N_45,In_88);
nand U228 (N_228,In_941,In_820);
nand U229 (N_229,In_192,In_373);
or U230 (N_230,In_932,In_65);
nand U231 (N_231,In_617,In_468);
nand U232 (N_232,In_891,In_877);
or U233 (N_233,In_287,In_246);
nand U234 (N_234,In_858,N_163);
and U235 (N_235,N_137,In_808);
and U236 (N_236,N_160,In_49);
or U237 (N_237,In_483,In_894);
nand U238 (N_238,In_314,In_155);
nor U239 (N_239,In_140,In_401);
nand U240 (N_240,In_629,In_754);
and U241 (N_241,In_726,N_8);
and U242 (N_242,N_162,N_195);
and U243 (N_243,In_942,In_552);
nor U244 (N_244,In_698,In_606);
nand U245 (N_245,In_164,In_37);
or U246 (N_246,N_76,In_461);
nand U247 (N_247,In_994,N_18);
nand U248 (N_248,In_260,In_50);
nor U249 (N_249,In_967,N_166);
nor U250 (N_250,In_76,In_547);
and U251 (N_251,In_349,In_96);
nor U252 (N_252,N_129,In_585);
nor U253 (N_253,In_395,In_651);
and U254 (N_254,N_39,In_997);
nor U255 (N_255,In_149,In_936);
and U256 (N_256,In_240,N_75);
and U257 (N_257,In_646,In_580);
nor U258 (N_258,In_973,In_381);
and U259 (N_259,N_150,In_117);
nand U260 (N_260,In_537,In_793);
and U261 (N_261,In_294,In_332);
nand U262 (N_262,In_346,In_404);
nor U263 (N_263,In_323,In_663);
nand U264 (N_264,In_239,N_32);
or U265 (N_265,N_120,N_167);
and U266 (N_266,In_414,N_54);
and U267 (N_267,In_43,In_882);
or U268 (N_268,In_917,In_42);
and U269 (N_269,N_24,In_473);
nand U270 (N_270,N_9,N_48);
and U271 (N_271,In_277,N_50);
nor U272 (N_272,In_266,In_288);
or U273 (N_273,In_437,In_673);
nand U274 (N_274,In_360,In_526);
and U275 (N_275,In_46,In_62);
or U276 (N_276,N_186,N_119);
nand U277 (N_277,In_964,In_861);
nand U278 (N_278,In_270,In_612);
and U279 (N_279,In_448,N_174);
and U280 (N_280,In_835,N_152);
and U281 (N_281,In_601,In_97);
nand U282 (N_282,In_969,In_784);
nand U283 (N_283,In_374,In_623);
nand U284 (N_284,In_800,N_151);
and U285 (N_285,In_716,In_469);
nor U286 (N_286,In_262,In_357);
nand U287 (N_287,In_342,N_187);
or U288 (N_288,In_829,N_176);
and U289 (N_289,N_41,N_170);
and U290 (N_290,In_826,N_101);
and U291 (N_291,N_55,N_154);
and U292 (N_292,In_782,N_115);
nand U293 (N_293,In_499,In_17);
and U294 (N_294,In_51,N_0);
and U295 (N_295,In_908,In_471);
nor U296 (N_296,In_630,In_965);
nor U297 (N_297,In_367,In_643);
and U298 (N_298,In_127,N_123);
nand U299 (N_299,In_540,In_572);
and U300 (N_300,N_146,In_44);
or U301 (N_301,In_528,In_834);
and U302 (N_302,N_142,In_434);
nor U303 (N_303,In_614,In_298);
nor U304 (N_304,N_122,In_227);
and U305 (N_305,In_256,In_879);
or U306 (N_306,N_17,In_878);
and U307 (N_307,N_165,In_387);
and U308 (N_308,In_397,In_274);
nand U309 (N_309,N_29,In_354);
and U310 (N_310,In_392,N_69);
or U311 (N_311,In_133,N_5);
and U312 (N_312,In_2,In_198);
or U313 (N_313,In_930,In_529);
and U314 (N_314,In_956,In_578);
and U315 (N_315,N_190,In_476);
or U316 (N_316,In_215,N_86);
and U317 (N_317,In_390,In_987);
and U318 (N_318,N_93,In_655);
nor U319 (N_319,In_228,N_61);
and U320 (N_320,In_685,In_797);
and U321 (N_321,N_168,N_49);
or U322 (N_322,In_807,N_56);
nor U323 (N_323,In_909,In_875);
and U324 (N_324,In_915,N_87);
and U325 (N_325,In_619,In_755);
nand U326 (N_326,In_697,In_940);
and U327 (N_327,In_416,In_588);
and U328 (N_328,In_144,N_113);
nand U329 (N_329,In_39,In_489);
or U330 (N_330,In_63,In_460);
and U331 (N_331,N_132,In_193);
nand U332 (N_332,In_333,N_149);
or U333 (N_333,N_73,In_781);
nor U334 (N_334,N_53,In_98);
nand U335 (N_335,In_650,In_740);
nor U336 (N_336,In_649,In_541);
nand U337 (N_337,In_607,N_15);
nand U338 (N_338,In_501,N_116);
and U339 (N_339,N_117,In_191);
nand U340 (N_340,N_197,In_695);
nor U341 (N_341,In_880,N_177);
nor U342 (N_342,In_32,N_35);
nand U343 (N_343,N_80,In_690);
nor U344 (N_344,In_595,In_574);
nor U345 (N_345,In_539,In_888);
nand U346 (N_346,In_902,N_127);
and U347 (N_347,In_372,In_874);
nor U348 (N_348,N_192,In_621);
or U349 (N_349,N_37,N_33);
or U350 (N_350,In_280,In_571);
or U351 (N_351,N_141,In_569);
or U352 (N_352,In_169,N_31);
or U353 (N_353,N_16,In_750);
nor U354 (N_354,In_79,N_159);
or U355 (N_355,N_13,In_290);
and U356 (N_356,In_53,N_7);
nand U357 (N_357,In_86,In_101);
or U358 (N_358,In_408,N_148);
nor U359 (N_359,In_804,In_642);
or U360 (N_360,In_161,In_493);
or U361 (N_361,In_31,In_919);
or U362 (N_362,In_162,In_85);
nand U363 (N_363,In_788,In_210);
and U364 (N_364,In_75,In_907);
nand U365 (N_365,In_648,In_738);
or U366 (N_366,In_388,In_208);
nand U367 (N_367,In_518,In_984);
and U368 (N_368,In_769,In_15);
and U369 (N_369,In_445,In_209);
or U370 (N_370,In_232,N_64);
and U371 (N_371,N_180,In_411);
nor U372 (N_372,In_652,In_821);
nor U373 (N_373,N_175,N_22);
nand U374 (N_374,In_558,In_705);
and U375 (N_375,In_115,In_730);
nand U376 (N_376,In_694,In_225);
nor U377 (N_377,In_250,In_199);
nand U378 (N_378,In_713,In_95);
and U379 (N_379,N_6,N_126);
nor U380 (N_380,In_660,N_94);
nand U381 (N_381,In_306,In_931);
nor U382 (N_382,In_864,In_36);
nor U383 (N_383,In_768,In_1);
nand U384 (N_384,In_179,In_691);
nand U385 (N_385,In_928,In_475);
and U386 (N_386,In_56,In_775);
and U387 (N_387,In_183,In_283);
nand U388 (N_388,In_291,In_377);
or U389 (N_389,In_107,In_443);
nor U390 (N_390,In_205,In_3);
nor U391 (N_391,In_269,In_824);
or U392 (N_392,N_164,In_327);
xnor U393 (N_393,N_91,N_193);
nand U394 (N_394,In_366,In_823);
nor U395 (N_395,In_732,In_866);
nor U396 (N_396,N_135,In_918);
and U397 (N_397,In_236,In_254);
and U398 (N_398,In_33,In_783);
nand U399 (N_399,In_480,N_182);
nor U400 (N_400,N_384,In_892);
and U401 (N_401,N_68,In_479);
nor U402 (N_402,In_234,In_249);
nor U403 (N_403,In_313,N_288);
nor U404 (N_404,In_550,In_825);
nor U405 (N_405,In_110,In_224);
nor U406 (N_406,N_333,In_573);
or U407 (N_407,In_474,N_171);
and U408 (N_408,N_353,In_696);
nand U409 (N_409,In_311,N_292);
nor U410 (N_410,In_143,In_531);
nor U411 (N_411,N_329,In_322);
nand U412 (N_412,In_767,N_248);
or U413 (N_413,N_1,N_234);
nor U414 (N_414,N_319,In_576);
and U415 (N_415,N_28,In_81);
or U416 (N_416,In_929,In_6);
nand U417 (N_417,In_678,In_722);
nor U418 (N_418,N_78,N_267);
and U419 (N_419,In_71,N_240);
nor U420 (N_420,N_315,In_505);
nor U421 (N_421,In_48,In_913);
nor U422 (N_422,N_107,In_123);
or U423 (N_423,N_275,In_447);
nor U424 (N_424,In_99,N_351);
or U425 (N_425,N_40,N_304);
and U426 (N_426,N_362,In_881);
or U427 (N_427,In_464,In_14);
and U428 (N_428,N_136,In_590);
nand U429 (N_429,N_259,In_549);
or U430 (N_430,N_383,N_381);
nand U431 (N_431,In_656,In_430);
nand U432 (N_432,In_131,N_380);
nand U433 (N_433,N_235,In_301);
nand U434 (N_434,In_610,In_105);
and U435 (N_435,In_188,N_134);
and U436 (N_436,In_22,In_187);
nand U437 (N_437,N_188,In_268);
or U438 (N_438,N_231,N_324);
or U439 (N_439,In_854,In_403);
nand U440 (N_440,In_715,N_373);
nand U441 (N_441,In_352,In_264);
and U442 (N_442,N_358,In_604);
nand U443 (N_443,N_222,In_358);
nor U444 (N_444,N_305,N_90);
or U445 (N_445,In_709,N_338);
and U446 (N_446,In_557,In_789);
or U447 (N_447,N_85,N_133);
or U448 (N_448,In_112,N_392);
nand U449 (N_449,N_228,In_535);
nor U450 (N_450,N_377,In_627);
nand U451 (N_451,In_564,In_795);
nand U452 (N_452,In_999,In_544);
and U453 (N_453,In_903,In_513);
nand U454 (N_454,N_249,In_364);
nor U455 (N_455,N_243,In_119);
nor U456 (N_456,N_251,N_318);
nor U457 (N_457,N_74,In_452);
or U458 (N_458,N_289,N_232);
nand U459 (N_459,N_343,N_286);
and U460 (N_460,N_349,N_140);
or U461 (N_461,In_896,In_844);
nand U462 (N_462,N_208,In_832);
and U463 (N_463,In_272,In_450);
nand U464 (N_464,In_562,In_859);
nor U465 (N_465,In_159,N_378);
or U466 (N_466,In_328,In_865);
nand U467 (N_467,In_433,In_887);
nand U468 (N_468,N_328,N_344);
nor U469 (N_469,In_752,N_214);
nand U470 (N_470,In_135,In_324);
nor U471 (N_471,N_246,In_382);
nor U472 (N_472,N_375,In_376);
nor U473 (N_473,In_522,N_198);
nor U474 (N_474,In_764,In_533);
or U475 (N_475,In_773,N_299);
and U476 (N_476,In_741,N_340);
nor U477 (N_477,N_282,N_96);
or U478 (N_478,N_312,In_482);
or U479 (N_479,In_702,N_67);
or U480 (N_480,N_30,In_35);
nand U481 (N_481,N_369,N_345);
and U482 (N_482,In_827,N_217);
or U483 (N_483,In_201,In_667);
and U484 (N_484,N_347,N_331);
nor U485 (N_485,In_171,N_43);
nand U486 (N_486,In_960,N_280);
nor U487 (N_487,In_276,In_765);
or U488 (N_488,N_211,In_618);
or U489 (N_489,In_822,In_634);
nor U490 (N_490,N_194,N_326);
nand U491 (N_491,N_58,In_581);
nand U492 (N_492,N_114,In_737);
or U493 (N_493,N_95,N_252);
nor U494 (N_494,N_396,N_274);
or U495 (N_495,N_11,In_641);
nor U496 (N_496,In_543,N_325);
nand U497 (N_497,In_369,N_223);
nand U498 (N_498,In_677,N_253);
nand U499 (N_499,In_596,In_424);
nor U500 (N_500,N_279,N_399);
and U501 (N_501,In_137,In_814);
nand U502 (N_502,In_271,In_664);
nand U503 (N_503,N_320,N_356);
xor U504 (N_504,In_933,In_446);
and U505 (N_505,In_319,In_575);
or U506 (N_506,N_110,N_44);
or U507 (N_507,N_161,In_744);
nor U508 (N_508,In_790,N_268);
or U509 (N_509,N_23,In_920);
nand U510 (N_510,N_153,N_111);
nor U511 (N_511,In_320,N_309);
nor U512 (N_512,In_745,In_297);
nor U513 (N_513,In_154,In_422);
or U514 (N_514,N_233,In_923);
and U515 (N_515,N_4,N_291);
nor U516 (N_516,In_868,In_325);
or U517 (N_517,In_204,N_297);
and U518 (N_518,In_219,N_365);
and U519 (N_519,In_870,In_348);
or U520 (N_520,N_302,In_724);
nand U521 (N_521,In_954,N_360);
nand U522 (N_522,In_330,N_155);
nand U523 (N_523,N_212,N_2);
nand U524 (N_524,N_368,In_344);
nor U525 (N_525,N_306,In_921);
and U526 (N_526,N_363,N_397);
nor U527 (N_527,N_284,N_62);
or U528 (N_528,N_265,N_81);
nor U529 (N_529,N_173,In_303);
and U530 (N_530,In_995,In_498);
nand U531 (N_531,In_504,In_633);
nor U532 (N_532,N_355,N_341);
and U533 (N_533,N_157,In_409);
nand U534 (N_534,In_370,N_372);
nor U535 (N_535,In_484,In_83);
nor U536 (N_536,In_872,N_247);
or U537 (N_537,N_322,N_82);
or U538 (N_538,N_112,N_236);
and U539 (N_539,In_584,In_567);
or U540 (N_540,In_837,N_391);
and U541 (N_541,In_632,N_60);
or U542 (N_542,In_279,In_148);
nand U543 (N_543,In_979,N_389);
or U544 (N_544,N_336,In_699);
or U545 (N_545,N_213,In_114);
xor U546 (N_546,In_23,In_904);
nor U547 (N_547,In_647,In_538);
or U548 (N_548,N_218,In_731);
nand U549 (N_549,In_26,N_144);
or U550 (N_550,N_323,In_776);
and U551 (N_551,In_273,In_487);
or U552 (N_552,In_689,N_348);
and U553 (N_553,N_14,In_296);
and U554 (N_554,N_346,In_255);
or U555 (N_555,In_222,In_704);
xnor U556 (N_556,In_207,In_840);
and U557 (N_557,In_418,N_287);
nor U558 (N_558,N_370,N_376);
nand U559 (N_559,N_63,N_385);
nand U560 (N_560,In_202,N_172);
nor U561 (N_561,In_66,In_343);
nand U562 (N_562,In_212,N_394);
or U563 (N_563,In_944,N_276);
and U564 (N_564,In_440,In_885);
nand U565 (N_565,In_293,N_335);
nand U566 (N_566,N_178,In_389);
and U567 (N_567,In_134,In_318);
and U568 (N_568,In_721,In_28);
and U569 (N_569,N_386,N_256);
or U570 (N_570,In_886,N_221);
nand U571 (N_571,In_860,N_334);
nand U572 (N_572,N_364,N_311);
or U573 (N_573,N_34,N_390);
nand U574 (N_574,N_65,N_205);
or U575 (N_575,N_238,In_743);
nand U576 (N_576,N_379,In_299);
or U577 (N_577,In_338,N_330);
and U578 (N_578,N_342,In_90);
nand U579 (N_579,In_281,N_321);
nand U580 (N_580,In_444,N_183);
or U581 (N_581,N_313,In_600);
or U582 (N_582,N_52,In_803);
or U583 (N_583,N_229,In_218);
nand U584 (N_584,In_492,In_889);
nor U585 (N_585,In_846,N_254);
nand U586 (N_586,N_296,In_310);
nor U587 (N_587,N_66,N_219);
nand U588 (N_588,In_850,N_79);
or U589 (N_589,N_388,N_21);
or U590 (N_590,In_454,N_272);
nor U591 (N_591,N_147,In_989);
nand U592 (N_592,N_260,In_622);
and U593 (N_593,In_615,In_196);
nand U594 (N_594,In_503,In_971);
nor U595 (N_595,N_202,N_283);
nor U596 (N_596,N_184,In_624);
nand U597 (N_597,N_124,N_209);
nand U598 (N_598,N_245,N_203);
and U599 (N_599,N_263,N_354);
nor U600 (N_600,N_493,In_703);
nor U601 (N_601,N_524,In_895);
and U602 (N_602,N_255,N_526);
nand U603 (N_603,N_507,N_71);
or U604 (N_604,In_451,N_224);
and U605 (N_605,N_206,N_216);
and U606 (N_606,N_542,N_121);
nand U607 (N_607,N_513,N_501);
nor U608 (N_608,N_307,N_465);
and U609 (N_609,In_326,In_109);
or U610 (N_610,In_855,N_512);
and U611 (N_611,In_185,N_100);
nand U612 (N_612,In_512,N_584);
nand U613 (N_613,N_540,In_828);
nor U614 (N_614,N_432,In_160);
or U615 (N_615,N_410,N_156);
or U616 (N_616,N_592,In_497);
and U617 (N_617,In_684,N_595);
and U618 (N_618,N_359,N_332);
or U619 (N_619,In_799,In_681);
nor U620 (N_620,N_552,N_487);
nor U621 (N_621,N_445,N_498);
and U622 (N_622,N_572,N_277);
or U623 (N_623,N_586,N_424);
and U624 (N_624,N_201,N_92);
or U625 (N_625,N_564,N_447);
or U626 (N_626,N_494,N_455);
and U627 (N_627,N_478,N_339);
nand U628 (N_628,N_371,N_588);
nor U629 (N_629,N_489,N_538);
nand U630 (N_630,In_70,N_409);
or U631 (N_631,N_463,N_430);
and U632 (N_632,In_517,N_543);
nor U633 (N_633,N_528,N_303);
nand U634 (N_634,N_495,N_143);
or U635 (N_635,N_468,N_527);
and U636 (N_636,N_200,N_20);
or U637 (N_637,In_384,N_273);
nand U638 (N_638,N_19,N_428);
and U639 (N_639,N_290,N_460);
nand U640 (N_640,N_416,In_947);
and U641 (N_641,N_502,N_529);
nor U642 (N_642,N_475,N_486);
nor U643 (N_643,N_565,In_261);
or U644 (N_644,N_587,N_374);
and U645 (N_645,N_361,N_443);
nand U646 (N_646,N_417,N_559);
nand U647 (N_647,N_453,N_497);
and U648 (N_648,N_293,N_450);
nor U649 (N_649,N_471,N_539);
or U650 (N_650,N_47,N_480);
or U651 (N_651,In_153,N_418);
nand U652 (N_652,In_10,N_519);
nand U653 (N_653,N_499,N_400);
nand U654 (N_654,In_64,N_131);
nor U655 (N_655,In_605,N_215);
nand U656 (N_656,N_549,In_173);
nor U657 (N_657,N_239,N_570);
or U658 (N_658,N_444,In_710);
or U659 (N_659,In_147,N_199);
and U660 (N_660,N_27,N_436);
nor U661 (N_661,In_486,N_36);
nor U662 (N_662,In_707,N_401);
or U663 (N_663,N_108,In_579);
or U664 (N_664,N_433,N_518);
nand U665 (N_665,N_503,In_353);
and U666 (N_666,N_598,N_461);
or U667 (N_667,In_762,N_207);
nor U668 (N_668,N_506,N_555);
nor U669 (N_669,In_157,N_533);
and U670 (N_670,In_331,N_594);
and U671 (N_671,N_230,N_250);
and U672 (N_672,N_300,N_181);
or U673 (N_673,N_504,In_396);
and U674 (N_674,In_679,In_351);
or U675 (N_675,N_553,N_3);
nor U676 (N_676,In_958,N_484);
nor U677 (N_677,N_479,N_422);
nand U678 (N_678,N_357,N_566);
nand U679 (N_679,N_412,N_281);
and U680 (N_680,N_337,N_568);
and U681 (N_681,N_597,N_99);
nor U682 (N_682,N_295,N_57);
or U683 (N_683,In_163,N_420);
nor U684 (N_684,N_278,In_355);
and U685 (N_685,N_407,N_84);
or U686 (N_686,In_61,N_352);
nor U687 (N_687,N_561,N_578);
nor U688 (N_688,N_467,N_474);
or U689 (N_689,N_558,N_548);
and U690 (N_690,N_261,N_556);
nand U691 (N_691,N_488,N_242);
nand U692 (N_692,N_257,N_546);
nor U693 (N_693,N_393,N_419);
nand U694 (N_694,N_589,N_258);
nor U695 (N_695,N_435,N_413);
or U696 (N_696,N_569,N_511);
and U697 (N_697,In_937,N_145);
nor U698 (N_698,In_145,N_462);
nor U699 (N_699,N_541,N_59);
or U700 (N_700,N_490,In_363);
nand U701 (N_701,In_780,N_226);
or U702 (N_702,N_196,In_168);
nand U703 (N_703,N_508,N_457);
or U704 (N_704,N_439,N_408);
or U705 (N_705,In_723,N_425);
nor U706 (N_706,N_220,N_492);
nand U707 (N_707,In_542,In_132);
nor U708 (N_708,N_314,N_25);
nand U709 (N_709,N_241,N_532);
and U710 (N_710,N_237,N_500);
or U711 (N_711,N_599,In_577);
nand U712 (N_712,N_262,N_464);
nand U713 (N_713,N_442,N_404);
or U714 (N_714,N_438,N_210);
nor U715 (N_715,N_105,In_640);
and U716 (N_716,In_841,N_515);
or U717 (N_717,N_459,N_316);
and U718 (N_718,In_978,N_411);
nand U719 (N_719,N_130,In_57);
or U720 (N_720,N_562,In_5);
and U721 (N_721,N_421,N_225);
nor U722 (N_722,In_949,N_466);
or U723 (N_723,In_975,N_366);
or U724 (N_724,N_590,N_530);
nor U725 (N_725,N_270,N_441);
and U726 (N_726,N_454,In_466);
nand U727 (N_727,In_719,N_579);
and U728 (N_728,N_525,N_535);
or U729 (N_729,N_405,N_536);
nand U730 (N_730,N_576,N_496);
and U731 (N_731,N_406,In_300);
nor U732 (N_732,N_98,N_310);
or U733 (N_733,In_241,N_327);
nand U734 (N_734,In_245,N_423);
nand U735 (N_735,N_550,N_317);
nor U736 (N_736,N_510,N_398);
nor U737 (N_737,In_819,N_573);
nor U738 (N_738,N_298,N_426);
or U739 (N_739,N_264,N_158);
or U740 (N_740,N_469,In_292);
nand U741 (N_741,In_849,N_477);
and U742 (N_742,N_308,N_476);
nor U743 (N_743,N_367,N_571);
or U744 (N_744,N_414,N_544);
nand U745 (N_745,N_128,N_350);
or U746 (N_746,N_522,In_30);
nand U747 (N_747,In_284,N_46);
nand U748 (N_748,N_179,In_645);
or U749 (N_749,In_329,In_405);
and U750 (N_750,N_514,In_233);
and U751 (N_751,N_591,N_382);
and U752 (N_752,In_993,N_554);
and U753 (N_753,N_26,N_563);
or U754 (N_754,N_545,N_271);
or U755 (N_755,In_974,In_838);
nor U756 (N_756,N_593,N_557);
and U757 (N_757,In_52,N_266);
nand U758 (N_758,In_432,In_912);
nor U759 (N_759,N_575,N_583);
nor U760 (N_760,N_403,N_451);
nand U761 (N_761,N_104,N_458);
nor U762 (N_762,N_547,In_751);
nand U763 (N_763,N_427,N_482);
nand U764 (N_764,In_682,In_337);
and U765 (N_765,N_585,N_431);
and U766 (N_766,N_83,In_545);
and U767 (N_767,N_537,N_440);
and U768 (N_768,N_531,N_227);
and U769 (N_769,In_84,N_185);
nand U770 (N_770,N_473,N_395);
or U771 (N_771,N_301,N_294);
and U772 (N_772,In_687,N_551);
or U773 (N_773,N_125,N_481);
or U774 (N_774,N_42,N_448);
and U775 (N_775,N_77,N_596);
nand U776 (N_776,In_152,N_567);
nand U777 (N_777,N_505,N_189);
nand U778 (N_778,N_523,In_455);
nand U779 (N_779,N_574,N_434);
nor U780 (N_780,N_517,N_429);
and U781 (N_781,N_437,In_514);
nor U782 (N_782,N_520,N_582);
nand U783 (N_783,N_581,N_402);
nand U784 (N_784,N_446,In_116);
nand U785 (N_785,In_688,N_452);
nand U786 (N_786,In_312,N_449);
or U787 (N_787,In_122,N_491);
nand U788 (N_788,N_204,N_483);
and U789 (N_789,N_97,N_387);
and U790 (N_790,N_456,In_977);
or U791 (N_791,In_927,N_509);
and U792 (N_792,N_580,N_244);
nor U793 (N_793,N_269,N_560);
nor U794 (N_794,N_415,N_285);
nor U795 (N_795,N_472,N_534);
or U796 (N_796,N_521,N_516);
and U797 (N_797,In_953,In_459);
nand U798 (N_798,N_470,N_577);
or U799 (N_799,N_139,N_485);
nand U800 (N_800,N_755,N_757);
nor U801 (N_801,N_708,N_785);
nand U802 (N_802,N_695,N_746);
nand U803 (N_803,N_783,N_779);
nor U804 (N_804,N_717,N_658);
nor U805 (N_805,N_628,N_644);
and U806 (N_806,N_676,N_633);
nor U807 (N_807,N_603,N_721);
or U808 (N_808,N_669,N_731);
or U809 (N_809,N_769,N_724);
nand U810 (N_810,N_601,N_743);
nand U811 (N_811,N_700,N_740);
nor U812 (N_812,N_733,N_610);
and U813 (N_813,N_798,N_795);
nand U814 (N_814,N_667,N_775);
nand U815 (N_815,N_675,N_638);
nor U816 (N_816,N_789,N_753);
or U817 (N_817,N_694,N_696);
or U818 (N_818,N_673,N_651);
or U819 (N_819,N_650,N_759);
and U820 (N_820,N_701,N_647);
nand U821 (N_821,N_776,N_698);
or U822 (N_822,N_631,N_712);
nor U823 (N_823,N_615,N_674);
or U824 (N_824,N_713,N_773);
nor U825 (N_825,N_774,N_672);
or U826 (N_826,N_679,N_691);
nand U827 (N_827,N_758,N_699);
or U828 (N_828,N_745,N_756);
or U829 (N_829,N_632,N_639);
and U830 (N_830,N_709,N_702);
nand U831 (N_831,N_682,N_749);
and U832 (N_832,N_778,N_792);
nor U833 (N_833,N_715,N_652);
or U834 (N_834,N_722,N_705);
nand U835 (N_835,N_787,N_747);
and U836 (N_836,N_616,N_767);
nor U837 (N_837,N_752,N_671);
nand U838 (N_838,N_666,N_681);
or U839 (N_839,N_734,N_687);
and U840 (N_840,N_661,N_780);
and U841 (N_841,N_744,N_623);
nor U842 (N_842,N_654,N_684);
or U843 (N_843,N_608,N_727);
and U844 (N_844,N_765,N_643);
nor U845 (N_845,N_604,N_613);
nand U846 (N_846,N_649,N_646);
nand U847 (N_847,N_737,N_750);
or U848 (N_848,N_609,N_707);
nand U849 (N_849,N_685,N_723);
and U850 (N_850,N_791,N_751);
nand U851 (N_851,N_635,N_636);
nand U852 (N_852,N_678,N_606);
nand U853 (N_853,N_720,N_600);
nand U854 (N_854,N_692,N_686);
and U855 (N_855,N_710,N_714);
or U856 (N_856,N_653,N_716);
nor U857 (N_857,N_732,N_602);
and U858 (N_858,N_784,N_683);
or U859 (N_859,N_624,N_754);
xor U860 (N_860,N_728,N_656);
or U861 (N_861,N_642,N_697);
nor U862 (N_862,N_761,N_660);
nor U863 (N_863,N_771,N_607);
nand U864 (N_864,N_766,N_663);
and U865 (N_865,N_781,N_680);
or U866 (N_866,N_736,N_620);
and U867 (N_867,N_772,N_763);
nor U868 (N_868,N_611,N_618);
and U869 (N_869,N_668,N_725);
or U870 (N_870,N_617,N_612);
nand U871 (N_871,N_782,N_645);
nor U872 (N_872,N_625,N_786);
nor U873 (N_873,N_735,N_762);
xor U874 (N_874,N_630,N_655);
nor U875 (N_875,N_796,N_648);
nor U876 (N_876,N_793,N_711);
or U877 (N_877,N_693,N_739);
nand U878 (N_878,N_622,N_690);
or U879 (N_879,N_794,N_788);
nand U880 (N_880,N_718,N_677);
nand U881 (N_881,N_777,N_659);
or U882 (N_882,N_726,N_605);
or U883 (N_883,N_729,N_738);
nand U884 (N_884,N_760,N_799);
nand U885 (N_885,N_742,N_790);
nand U886 (N_886,N_614,N_703);
and U887 (N_887,N_719,N_665);
nor U888 (N_888,N_662,N_704);
or U889 (N_889,N_627,N_619);
nor U890 (N_890,N_689,N_706);
nor U891 (N_891,N_640,N_629);
and U892 (N_892,N_657,N_626);
nand U893 (N_893,N_748,N_688);
nand U894 (N_894,N_797,N_664);
xor U895 (N_895,N_770,N_730);
or U896 (N_896,N_621,N_768);
nand U897 (N_897,N_741,N_641);
or U898 (N_898,N_670,N_637);
and U899 (N_899,N_764,N_634);
nor U900 (N_900,N_760,N_656);
nand U901 (N_901,N_757,N_780);
and U902 (N_902,N_747,N_689);
nand U903 (N_903,N_613,N_797);
nand U904 (N_904,N_784,N_770);
nor U905 (N_905,N_725,N_746);
nor U906 (N_906,N_661,N_745);
and U907 (N_907,N_626,N_694);
or U908 (N_908,N_750,N_741);
or U909 (N_909,N_754,N_744);
nor U910 (N_910,N_752,N_738);
nand U911 (N_911,N_656,N_676);
nand U912 (N_912,N_701,N_775);
nor U913 (N_913,N_703,N_688);
nand U914 (N_914,N_729,N_776);
and U915 (N_915,N_771,N_676);
and U916 (N_916,N_778,N_655);
nor U917 (N_917,N_716,N_692);
nor U918 (N_918,N_623,N_706);
nand U919 (N_919,N_787,N_616);
nand U920 (N_920,N_730,N_668);
and U921 (N_921,N_785,N_773);
and U922 (N_922,N_630,N_620);
or U923 (N_923,N_638,N_793);
nor U924 (N_924,N_605,N_770);
and U925 (N_925,N_648,N_778);
and U926 (N_926,N_776,N_749);
nor U927 (N_927,N_684,N_627);
nand U928 (N_928,N_671,N_600);
or U929 (N_929,N_769,N_657);
and U930 (N_930,N_655,N_672);
nor U931 (N_931,N_771,N_635);
nand U932 (N_932,N_640,N_648);
and U933 (N_933,N_679,N_607);
nor U934 (N_934,N_790,N_631);
or U935 (N_935,N_653,N_738);
or U936 (N_936,N_762,N_731);
and U937 (N_937,N_747,N_793);
nand U938 (N_938,N_610,N_698);
nor U939 (N_939,N_600,N_740);
or U940 (N_940,N_781,N_791);
nor U941 (N_941,N_658,N_689);
nor U942 (N_942,N_717,N_738);
and U943 (N_943,N_777,N_641);
nor U944 (N_944,N_668,N_639);
nand U945 (N_945,N_678,N_719);
nor U946 (N_946,N_740,N_706);
or U947 (N_947,N_715,N_687);
and U948 (N_948,N_747,N_656);
nand U949 (N_949,N_797,N_740);
or U950 (N_950,N_776,N_601);
or U951 (N_951,N_624,N_712);
or U952 (N_952,N_693,N_632);
nor U953 (N_953,N_652,N_702);
and U954 (N_954,N_603,N_605);
and U955 (N_955,N_717,N_740);
nand U956 (N_956,N_601,N_733);
nor U957 (N_957,N_701,N_769);
nor U958 (N_958,N_721,N_771);
nand U959 (N_959,N_635,N_678);
or U960 (N_960,N_615,N_798);
and U961 (N_961,N_767,N_764);
and U962 (N_962,N_612,N_642);
nor U963 (N_963,N_689,N_754);
and U964 (N_964,N_786,N_622);
or U965 (N_965,N_615,N_646);
and U966 (N_966,N_711,N_761);
or U967 (N_967,N_633,N_658);
nor U968 (N_968,N_678,N_661);
nor U969 (N_969,N_783,N_603);
nor U970 (N_970,N_758,N_742);
nor U971 (N_971,N_767,N_675);
nand U972 (N_972,N_766,N_775);
nand U973 (N_973,N_649,N_633);
and U974 (N_974,N_628,N_764);
or U975 (N_975,N_775,N_789);
nor U976 (N_976,N_629,N_792);
and U977 (N_977,N_707,N_698);
nor U978 (N_978,N_730,N_768);
nand U979 (N_979,N_630,N_757);
nor U980 (N_980,N_673,N_614);
and U981 (N_981,N_646,N_725);
or U982 (N_982,N_786,N_603);
nand U983 (N_983,N_662,N_663);
nand U984 (N_984,N_683,N_704);
and U985 (N_985,N_738,N_719);
nor U986 (N_986,N_767,N_758);
and U987 (N_987,N_634,N_771);
nor U988 (N_988,N_732,N_715);
and U989 (N_989,N_784,N_690);
and U990 (N_990,N_729,N_788);
and U991 (N_991,N_762,N_748);
and U992 (N_992,N_783,N_606);
nand U993 (N_993,N_777,N_694);
nand U994 (N_994,N_680,N_673);
nand U995 (N_995,N_736,N_767);
and U996 (N_996,N_682,N_605);
nand U997 (N_997,N_658,N_725);
nand U998 (N_998,N_686,N_629);
and U999 (N_999,N_760,N_704);
and U1000 (N_1000,N_917,N_949);
nor U1001 (N_1001,N_945,N_852);
nor U1002 (N_1002,N_976,N_872);
nand U1003 (N_1003,N_902,N_865);
and U1004 (N_1004,N_828,N_842);
or U1005 (N_1005,N_815,N_996);
nand U1006 (N_1006,N_812,N_894);
nor U1007 (N_1007,N_994,N_823);
nand U1008 (N_1008,N_809,N_911);
nor U1009 (N_1009,N_983,N_855);
nor U1010 (N_1010,N_951,N_824);
nor U1011 (N_1011,N_924,N_856);
nor U1012 (N_1012,N_849,N_891);
nand U1013 (N_1013,N_825,N_800);
xor U1014 (N_1014,N_999,N_897);
nor U1015 (N_1015,N_948,N_990);
or U1016 (N_1016,N_882,N_942);
nor U1017 (N_1017,N_975,N_862);
nor U1018 (N_1018,N_916,N_946);
or U1019 (N_1019,N_811,N_851);
or U1020 (N_1020,N_907,N_866);
nor U1021 (N_1021,N_845,N_914);
or U1022 (N_1022,N_889,N_892);
or U1023 (N_1023,N_805,N_879);
nand U1024 (N_1024,N_909,N_989);
or U1025 (N_1025,N_933,N_880);
nor U1026 (N_1026,N_972,N_884);
nand U1027 (N_1027,N_968,N_806);
and U1028 (N_1028,N_804,N_912);
and U1029 (N_1029,N_817,N_858);
nand U1030 (N_1030,N_992,N_934);
nand U1031 (N_1031,N_887,N_843);
nand U1032 (N_1032,N_844,N_985);
or U1033 (N_1033,N_939,N_931);
nand U1034 (N_1034,N_877,N_910);
nand U1035 (N_1035,N_860,N_839);
nand U1036 (N_1036,N_923,N_873);
nand U1037 (N_1037,N_955,N_921);
nor U1038 (N_1038,N_875,N_871);
nand U1039 (N_1039,N_928,N_957);
or U1040 (N_1040,N_970,N_926);
nand U1041 (N_1041,N_956,N_941);
nand U1042 (N_1042,N_920,N_995);
nor U1043 (N_1043,N_965,N_922);
and U1044 (N_1044,N_973,N_846);
or U1045 (N_1045,N_859,N_867);
nor U1046 (N_1046,N_803,N_881);
or U1047 (N_1047,N_818,N_937);
nand U1048 (N_1048,N_890,N_982);
or U1049 (N_1049,N_962,N_930);
or U1050 (N_1050,N_953,N_961);
nor U1051 (N_1051,N_807,N_906);
nand U1052 (N_1052,N_997,N_898);
and U1053 (N_1053,N_834,N_993);
or U1054 (N_1054,N_896,N_838);
nand U1055 (N_1055,N_952,N_827);
or U1056 (N_1056,N_940,N_905);
or U1057 (N_1057,N_863,N_984);
nand U1058 (N_1058,N_904,N_981);
nand U1059 (N_1059,N_813,N_848);
nor U1060 (N_1060,N_814,N_980);
or U1061 (N_1061,N_927,N_963);
nand U1062 (N_1062,N_850,N_954);
nor U1063 (N_1063,N_998,N_895);
nor U1064 (N_1064,N_893,N_925);
nand U1065 (N_1065,N_801,N_883);
nor U1066 (N_1066,N_938,N_836);
and U1067 (N_1067,N_829,N_853);
or U1068 (N_1068,N_874,N_903);
and U1069 (N_1069,N_857,N_950);
or U1070 (N_1070,N_988,N_919);
or U1071 (N_1071,N_932,N_847);
nor U1072 (N_1072,N_802,N_822);
and U1073 (N_1073,N_900,N_915);
nand U1074 (N_1074,N_830,N_826);
or U1075 (N_1075,N_816,N_835);
nand U1076 (N_1076,N_885,N_959);
nand U1077 (N_1077,N_918,N_958);
or U1078 (N_1078,N_854,N_929);
and U1079 (N_1079,N_870,N_947);
or U1080 (N_1080,N_978,N_966);
or U1081 (N_1081,N_837,N_841);
and U1082 (N_1082,N_964,N_840);
nand U1083 (N_1083,N_832,N_886);
or U1084 (N_1084,N_908,N_868);
and U1085 (N_1085,N_820,N_913);
nor U1086 (N_1086,N_831,N_878);
or U1087 (N_1087,N_969,N_899);
and U1088 (N_1088,N_869,N_986);
and U1089 (N_1089,N_974,N_808);
or U1090 (N_1090,N_810,N_833);
nor U1091 (N_1091,N_936,N_967);
or U1092 (N_1092,N_876,N_821);
nor U1093 (N_1093,N_819,N_979);
nand U1094 (N_1094,N_943,N_888);
nand U1095 (N_1095,N_960,N_901);
or U1096 (N_1096,N_971,N_864);
and U1097 (N_1097,N_944,N_987);
nor U1098 (N_1098,N_991,N_935);
and U1099 (N_1099,N_977,N_861);
and U1100 (N_1100,N_860,N_994);
or U1101 (N_1101,N_881,N_935);
and U1102 (N_1102,N_866,N_990);
or U1103 (N_1103,N_941,N_979);
nand U1104 (N_1104,N_916,N_880);
or U1105 (N_1105,N_969,N_941);
xor U1106 (N_1106,N_949,N_807);
nand U1107 (N_1107,N_992,N_849);
nor U1108 (N_1108,N_951,N_981);
nor U1109 (N_1109,N_999,N_853);
nor U1110 (N_1110,N_873,N_943);
and U1111 (N_1111,N_922,N_944);
or U1112 (N_1112,N_862,N_825);
nand U1113 (N_1113,N_974,N_951);
or U1114 (N_1114,N_850,N_857);
nand U1115 (N_1115,N_874,N_804);
nand U1116 (N_1116,N_886,N_889);
and U1117 (N_1117,N_825,N_804);
nor U1118 (N_1118,N_868,N_849);
nor U1119 (N_1119,N_929,N_862);
or U1120 (N_1120,N_981,N_992);
nor U1121 (N_1121,N_927,N_944);
nor U1122 (N_1122,N_996,N_847);
and U1123 (N_1123,N_853,N_870);
and U1124 (N_1124,N_811,N_947);
nor U1125 (N_1125,N_959,N_859);
nand U1126 (N_1126,N_840,N_955);
or U1127 (N_1127,N_841,N_933);
or U1128 (N_1128,N_839,N_900);
nor U1129 (N_1129,N_830,N_963);
nor U1130 (N_1130,N_926,N_933);
nor U1131 (N_1131,N_803,N_827);
and U1132 (N_1132,N_852,N_813);
nor U1133 (N_1133,N_911,N_931);
nand U1134 (N_1134,N_850,N_941);
nand U1135 (N_1135,N_845,N_818);
nand U1136 (N_1136,N_910,N_941);
nor U1137 (N_1137,N_984,N_867);
or U1138 (N_1138,N_982,N_870);
and U1139 (N_1139,N_960,N_968);
nor U1140 (N_1140,N_880,N_889);
and U1141 (N_1141,N_827,N_891);
nor U1142 (N_1142,N_857,N_803);
and U1143 (N_1143,N_979,N_913);
or U1144 (N_1144,N_911,N_999);
nor U1145 (N_1145,N_829,N_885);
nand U1146 (N_1146,N_833,N_883);
nor U1147 (N_1147,N_904,N_828);
or U1148 (N_1148,N_907,N_881);
and U1149 (N_1149,N_803,N_840);
nor U1150 (N_1150,N_933,N_932);
nand U1151 (N_1151,N_980,N_975);
nor U1152 (N_1152,N_865,N_889);
and U1153 (N_1153,N_978,N_935);
nand U1154 (N_1154,N_915,N_825);
and U1155 (N_1155,N_947,N_888);
nand U1156 (N_1156,N_989,N_833);
and U1157 (N_1157,N_978,N_963);
nor U1158 (N_1158,N_851,N_954);
or U1159 (N_1159,N_973,N_917);
and U1160 (N_1160,N_937,N_961);
and U1161 (N_1161,N_836,N_962);
or U1162 (N_1162,N_820,N_945);
nand U1163 (N_1163,N_963,N_899);
and U1164 (N_1164,N_809,N_920);
nor U1165 (N_1165,N_986,N_832);
nand U1166 (N_1166,N_818,N_913);
and U1167 (N_1167,N_984,N_904);
xnor U1168 (N_1168,N_816,N_958);
or U1169 (N_1169,N_889,N_806);
nor U1170 (N_1170,N_803,N_934);
nor U1171 (N_1171,N_906,N_868);
and U1172 (N_1172,N_818,N_879);
or U1173 (N_1173,N_862,N_838);
or U1174 (N_1174,N_819,N_929);
nand U1175 (N_1175,N_842,N_914);
and U1176 (N_1176,N_919,N_818);
nor U1177 (N_1177,N_949,N_837);
and U1178 (N_1178,N_817,N_857);
and U1179 (N_1179,N_959,N_999);
nand U1180 (N_1180,N_855,N_853);
and U1181 (N_1181,N_839,N_865);
nand U1182 (N_1182,N_908,N_941);
nor U1183 (N_1183,N_876,N_850);
nor U1184 (N_1184,N_827,N_937);
nand U1185 (N_1185,N_971,N_892);
nor U1186 (N_1186,N_838,N_987);
or U1187 (N_1187,N_911,N_935);
and U1188 (N_1188,N_819,N_881);
nand U1189 (N_1189,N_887,N_821);
nor U1190 (N_1190,N_871,N_805);
and U1191 (N_1191,N_988,N_941);
and U1192 (N_1192,N_807,N_845);
nor U1193 (N_1193,N_952,N_895);
nor U1194 (N_1194,N_839,N_854);
or U1195 (N_1195,N_892,N_880);
nand U1196 (N_1196,N_888,N_885);
or U1197 (N_1197,N_873,N_907);
and U1198 (N_1198,N_926,N_978);
or U1199 (N_1199,N_972,N_845);
nor U1200 (N_1200,N_1038,N_1034);
and U1201 (N_1201,N_1195,N_1010);
or U1202 (N_1202,N_1063,N_1095);
and U1203 (N_1203,N_1125,N_1190);
or U1204 (N_1204,N_1120,N_1102);
nand U1205 (N_1205,N_1033,N_1153);
and U1206 (N_1206,N_1019,N_1179);
nor U1207 (N_1207,N_1029,N_1178);
and U1208 (N_1208,N_1139,N_1154);
or U1209 (N_1209,N_1087,N_1091);
nand U1210 (N_1210,N_1057,N_1182);
nand U1211 (N_1211,N_1148,N_1072);
or U1212 (N_1212,N_1162,N_1198);
and U1213 (N_1213,N_1022,N_1068);
and U1214 (N_1214,N_1160,N_1174);
and U1215 (N_1215,N_1150,N_1168);
nor U1216 (N_1216,N_1058,N_1144);
or U1217 (N_1217,N_1074,N_1082);
or U1218 (N_1218,N_1056,N_1170);
nand U1219 (N_1219,N_1166,N_1042);
and U1220 (N_1220,N_1151,N_1081);
nor U1221 (N_1221,N_1061,N_1023);
nor U1222 (N_1222,N_1096,N_1141);
nor U1223 (N_1223,N_1027,N_1066);
and U1224 (N_1224,N_1197,N_1191);
nor U1225 (N_1225,N_1110,N_1075);
nand U1226 (N_1226,N_1051,N_1052);
nor U1227 (N_1227,N_1124,N_1009);
nor U1228 (N_1228,N_1177,N_1156);
or U1229 (N_1229,N_1099,N_1085);
or U1230 (N_1230,N_1136,N_1123);
nand U1231 (N_1231,N_1172,N_1006);
nand U1232 (N_1232,N_1107,N_1089);
and U1233 (N_1233,N_1180,N_1014);
nand U1234 (N_1234,N_1069,N_1059);
or U1235 (N_1235,N_1186,N_1181);
nor U1236 (N_1236,N_1005,N_1055);
and U1237 (N_1237,N_1012,N_1094);
or U1238 (N_1238,N_1024,N_1127);
or U1239 (N_1239,N_1113,N_1163);
and U1240 (N_1240,N_1106,N_1031);
nor U1241 (N_1241,N_1115,N_1088);
nand U1242 (N_1242,N_1011,N_1043);
or U1243 (N_1243,N_1128,N_1000);
nor U1244 (N_1244,N_1002,N_1070);
and U1245 (N_1245,N_1134,N_1001);
nor U1246 (N_1246,N_1013,N_1086);
nor U1247 (N_1247,N_1080,N_1194);
nand U1248 (N_1248,N_1126,N_1041);
nor U1249 (N_1249,N_1103,N_1093);
nor U1250 (N_1250,N_1114,N_1155);
and U1251 (N_1251,N_1003,N_1129);
or U1252 (N_1252,N_1049,N_1111);
or U1253 (N_1253,N_1077,N_1193);
and U1254 (N_1254,N_1036,N_1108);
and U1255 (N_1255,N_1025,N_1116);
nand U1256 (N_1256,N_1045,N_1092);
and U1257 (N_1257,N_1135,N_1062);
nand U1258 (N_1258,N_1083,N_1021);
nand U1259 (N_1259,N_1164,N_1140);
or U1260 (N_1260,N_1100,N_1048);
and U1261 (N_1261,N_1132,N_1188);
or U1262 (N_1262,N_1053,N_1112);
nand U1263 (N_1263,N_1071,N_1078);
nor U1264 (N_1264,N_1101,N_1020);
nor U1265 (N_1265,N_1050,N_1187);
nor U1266 (N_1266,N_1165,N_1054);
or U1267 (N_1267,N_1184,N_1143);
nand U1268 (N_1268,N_1098,N_1146);
or U1269 (N_1269,N_1035,N_1161);
nand U1270 (N_1270,N_1133,N_1064);
nor U1271 (N_1271,N_1142,N_1131);
nor U1272 (N_1272,N_1137,N_1199);
and U1273 (N_1273,N_1007,N_1105);
or U1274 (N_1274,N_1147,N_1060);
or U1275 (N_1275,N_1040,N_1037);
or U1276 (N_1276,N_1145,N_1118);
or U1277 (N_1277,N_1167,N_1183);
nand U1278 (N_1278,N_1169,N_1104);
or U1279 (N_1279,N_1196,N_1032);
and U1280 (N_1280,N_1175,N_1073);
and U1281 (N_1281,N_1015,N_1192);
or U1282 (N_1282,N_1030,N_1084);
or U1283 (N_1283,N_1026,N_1138);
nand U1284 (N_1284,N_1067,N_1157);
nor U1285 (N_1285,N_1189,N_1008);
nand U1286 (N_1286,N_1028,N_1079);
nand U1287 (N_1287,N_1185,N_1018);
nor U1288 (N_1288,N_1016,N_1039);
nor U1289 (N_1289,N_1117,N_1159);
nor U1290 (N_1290,N_1173,N_1122);
and U1291 (N_1291,N_1158,N_1047);
and U1292 (N_1292,N_1121,N_1149);
nand U1293 (N_1293,N_1046,N_1109);
or U1294 (N_1294,N_1017,N_1065);
or U1295 (N_1295,N_1090,N_1004);
and U1296 (N_1296,N_1119,N_1176);
and U1297 (N_1297,N_1044,N_1076);
nand U1298 (N_1298,N_1130,N_1152);
or U1299 (N_1299,N_1097,N_1171);
nor U1300 (N_1300,N_1107,N_1037);
and U1301 (N_1301,N_1042,N_1101);
or U1302 (N_1302,N_1167,N_1152);
or U1303 (N_1303,N_1058,N_1103);
or U1304 (N_1304,N_1085,N_1002);
or U1305 (N_1305,N_1147,N_1092);
or U1306 (N_1306,N_1141,N_1102);
nand U1307 (N_1307,N_1100,N_1047);
nand U1308 (N_1308,N_1179,N_1089);
and U1309 (N_1309,N_1034,N_1153);
nand U1310 (N_1310,N_1031,N_1123);
and U1311 (N_1311,N_1025,N_1161);
nand U1312 (N_1312,N_1149,N_1058);
nand U1313 (N_1313,N_1084,N_1022);
and U1314 (N_1314,N_1138,N_1040);
or U1315 (N_1315,N_1061,N_1118);
nand U1316 (N_1316,N_1010,N_1095);
nor U1317 (N_1317,N_1002,N_1072);
or U1318 (N_1318,N_1004,N_1038);
or U1319 (N_1319,N_1154,N_1169);
and U1320 (N_1320,N_1096,N_1170);
or U1321 (N_1321,N_1180,N_1018);
and U1322 (N_1322,N_1176,N_1180);
and U1323 (N_1323,N_1071,N_1009);
and U1324 (N_1324,N_1131,N_1103);
nor U1325 (N_1325,N_1066,N_1042);
and U1326 (N_1326,N_1181,N_1184);
nand U1327 (N_1327,N_1043,N_1073);
or U1328 (N_1328,N_1102,N_1015);
nor U1329 (N_1329,N_1071,N_1194);
nand U1330 (N_1330,N_1014,N_1023);
and U1331 (N_1331,N_1162,N_1177);
and U1332 (N_1332,N_1085,N_1075);
nand U1333 (N_1333,N_1046,N_1074);
nand U1334 (N_1334,N_1058,N_1069);
and U1335 (N_1335,N_1060,N_1042);
nand U1336 (N_1336,N_1094,N_1186);
or U1337 (N_1337,N_1112,N_1030);
nor U1338 (N_1338,N_1116,N_1153);
and U1339 (N_1339,N_1108,N_1188);
nor U1340 (N_1340,N_1038,N_1084);
nand U1341 (N_1341,N_1162,N_1081);
or U1342 (N_1342,N_1153,N_1022);
nand U1343 (N_1343,N_1191,N_1033);
and U1344 (N_1344,N_1063,N_1131);
nor U1345 (N_1345,N_1000,N_1054);
and U1346 (N_1346,N_1196,N_1136);
or U1347 (N_1347,N_1015,N_1084);
nand U1348 (N_1348,N_1133,N_1127);
and U1349 (N_1349,N_1065,N_1177);
and U1350 (N_1350,N_1099,N_1121);
or U1351 (N_1351,N_1043,N_1156);
nor U1352 (N_1352,N_1103,N_1156);
and U1353 (N_1353,N_1120,N_1123);
nand U1354 (N_1354,N_1038,N_1079);
nor U1355 (N_1355,N_1083,N_1139);
nand U1356 (N_1356,N_1140,N_1009);
and U1357 (N_1357,N_1039,N_1024);
and U1358 (N_1358,N_1089,N_1133);
nand U1359 (N_1359,N_1101,N_1032);
or U1360 (N_1360,N_1181,N_1001);
nand U1361 (N_1361,N_1094,N_1095);
nand U1362 (N_1362,N_1135,N_1080);
nor U1363 (N_1363,N_1016,N_1102);
nor U1364 (N_1364,N_1100,N_1164);
nor U1365 (N_1365,N_1059,N_1147);
nor U1366 (N_1366,N_1198,N_1194);
nand U1367 (N_1367,N_1052,N_1183);
and U1368 (N_1368,N_1021,N_1191);
or U1369 (N_1369,N_1064,N_1181);
or U1370 (N_1370,N_1067,N_1140);
or U1371 (N_1371,N_1073,N_1091);
nand U1372 (N_1372,N_1133,N_1020);
or U1373 (N_1373,N_1052,N_1134);
nor U1374 (N_1374,N_1049,N_1053);
nand U1375 (N_1375,N_1125,N_1179);
nand U1376 (N_1376,N_1138,N_1029);
and U1377 (N_1377,N_1073,N_1190);
nand U1378 (N_1378,N_1157,N_1184);
and U1379 (N_1379,N_1066,N_1192);
and U1380 (N_1380,N_1099,N_1054);
or U1381 (N_1381,N_1165,N_1024);
or U1382 (N_1382,N_1157,N_1081);
or U1383 (N_1383,N_1153,N_1037);
or U1384 (N_1384,N_1140,N_1077);
or U1385 (N_1385,N_1140,N_1158);
and U1386 (N_1386,N_1041,N_1101);
nand U1387 (N_1387,N_1181,N_1166);
nand U1388 (N_1388,N_1171,N_1192);
nor U1389 (N_1389,N_1019,N_1018);
nor U1390 (N_1390,N_1138,N_1038);
and U1391 (N_1391,N_1010,N_1067);
and U1392 (N_1392,N_1025,N_1098);
and U1393 (N_1393,N_1100,N_1074);
and U1394 (N_1394,N_1160,N_1029);
nor U1395 (N_1395,N_1157,N_1009);
nor U1396 (N_1396,N_1006,N_1060);
and U1397 (N_1397,N_1147,N_1139);
nand U1398 (N_1398,N_1119,N_1014);
and U1399 (N_1399,N_1150,N_1058);
and U1400 (N_1400,N_1352,N_1263);
or U1401 (N_1401,N_1284,N_1222);
and U1402 (N_1402,N_1340,N_1304);
nand U1403 (N_1403,N_1314,N_1216);
and U1404 (N_1404,N_1242,N_1296);
nand U1405 (N_1405,N_1337,N_1321);
or U1406 (N_1406,N_1245,N_1240);
or U1407 (N_1407,N_1287,N_1206);
or U1408 (N_1408,N_1346,N_1388);
or U1409 (N_1409,N_1248,N_1289);
or U1410 (N_1410,N_1210,N_1246);
nor U1411 (N_1411,N_1267,N_1244);
and U1412 (N_1412,N_1286,N_1344);
and U1413 (N_1413,N_1350,N_1367);
nor U1414 (N_1414,N_1227,N_1396);
nor U1415 (N_1415,N_1270,N_1279);
nor U1416 (N_1416,N_1241,N_1376);
and U1417 (N_1417,N_1306,N_1207);
nor U1418 (N_1418,N_1260,N_1282);
nand U1419 (N_1419,N_1293,N_1272);
and U1420 (N_1420,N_1239,N_1379);
nand U1421 (N_1421,N_1274,N_1230);
nand U1422 (N_1422,N_1370,N_1257);
or U1423 (N_1423,N_1285,N_1372);
nor U1424 (N_1424,N_1330,N_1301);
and U1425 (N_1425,N_1250,N_1358);
or U1426 (N_1426,N_1317,N_1366);
and U1427 (N_1427,N_1312,N_1364);
nor U1428 (N_1428,N_1353,N_1271);
nand U1429 (N_1429,N_1217,N_1223);
or U1430 (N_1430,N_1323,N_1343);
and U1431 (N_1431,N_1234,N_1215);
nand U1432 (N_1432,N_1313,N_1386);
nor U1433 (N_1433,N_1324,N_1292);
nand U1434 (N_1434,N_1318,N_1235);
or U1435 (N_1435,N_1208,N_1373);
nor U1436 (N_1436,N_1236,N_1209);
and U1437 (N_1437,N_1362,N_1225);
nor U1438 (N_1438,N_1204,N_1348);
or U1439 (N_1439,N_1275,N_1345);
and U1440 (N_1440,N_1331,N_1398);
or U1441 (N_1441,N_1214,N_1221);
nor U1442 (N_1442,N_1395,N_1202);
nor U1443 (N_1443,N_1384,N_1276);
and U1444 (N_1444,N_1299,N_1392);
and U1445 (N_1445,N_1322,N_1375);
and U1446 (N_1446,N_1300,N_1297);
or U1447 (N_1447,N_1360,N_1336);
and U1448 (N_1448,N_1365,N_1291);
and U1449 (N_1449,N_1211,N_1254);
xnor U1450 (N_1450,N_1247,N_1233);
nor U1451 (N_1451,N_1231,N_1377);
nor U1452 (N_1452,N_1309,N_1264);
or U1453 (N_1453,N_1385,N_1203);
nor U1454 (N_1454,N_1213,N_1268);
nand U1455 (N_1455,N_1391,N_1361);
and U1456 (N_1456,N_1371,N_1277);
or U1457 (N_1457,N_1338,N_1351);
nand U1458 (N_1458,N_1243,N_1315);
nand U1459 (N_1459,N_1394,N_1229);
and U1460 (N_1460,N_1320,N_1380);
nor U1461 (N_1461,N_1387,N_1238);
and U1462 (N_1462,N_1294,N_1355);
and U1463 (N_1463,N_1265,N_1278);
nand U1464 (N_1464,N_1266,N_1326);
nand U1465 (N_1465,N_1383,N_1381);
nand U1466 (N_1466,N_1325,N_1232);
and U1467 (N_1467,N_1332,N_1224);
and U1468 (N_1468,N_1220,N_1339);
nand U1469 (N_1469,N_1356,N_1354);
nand U1470 (N_1470,N_1281,N_1359);
and U1471 (N_1471,N_1251,N_1218);
or U1472 (N_1472,N_1261,N_1393);
xnor U1473 (N_1473,N_1305,N_1335);
and U1474 (N_1474,N_1295,N_1347);
and U1475 (N_1475,N_1200,N_1328);
nor U1476 (N_1476,N_1357,N_1226);
nor U1477 (N_1477,N_1397,N_1298);
and U1478 (N_1478,N_1237,N_1333);
nand U1479 (N_1479,N_1389,N_1368);
nand U1480 (N_1480,N_1349,N_1283);
nand U1481 (N_1481,N_1253,N_1273);
or U1482 (N_1482,N_1262,N_1363);
or U1483 (N_1483,N_1342,N_1399);
nand U1484 (N_1484,N_1319,N_1205);
nor U1485 (N_1485,N_1327,N_1269);
or U1486 (N_1486,N_1219,N_1307);
and U1487 (N_1487,N_1259,N_1310);
nor U1488 (N_1488,N_1378,N_1302);
nand U1489 (N_1489,N_1382,N_1290);
and U1490 (N_1490,N_1308,N_1334);
and U1491 (N_1491,N_1369,N_1374);
or U1492 (N_1492,N_1311,N_1329);
nand U1493 (N_1493,N_1255,N_1228);
and U1494 (N_1494,N_1288,N_1316);
and U1495 (N_1495,N_1252,N_1256);
nand U1496 (N_1496,N_1249,N_1341);
nor U1497 (N_1497,N_1280,N_1212);
or U1498 (N_1498,N_1258,N_1390);
nand U1499 (N_1499,N_1201,N_1303);
and U1500 (N_1500,N_1368,N_1393);
or U1501 (N_1501,N_1240,N_1324);
nor U1502 (N_1502,N_1201,N_1327);
nor U1503 (N_1503,N_1233,N_1264);
and U1504 (N_1504,N_1324,N_1396);
nor U1505 (N_1505,N_1352,N_1310);
nor U1506 (N_1506,N_1375,N_1235);
and U1507 (N_1507,N_1352,N_1295);
nand U1508 (N_1508,N_1327,N_1207);
nand U1509 (N_1509,N_1348,N_1379);
nor U1510 (N_1510,N_1369,N_1356);
or U1511 (N_1511,N_1384,N_1275);
nor U1512 (N_1512,N_1312,N_1317);
nor U1513 (N_1513,N_1269,N_1296);
or U1514 (N_1514,N_1352,N_1383);
or U1515 (N_1515,N_1309,N_1260);
nand U1516 (N_1516,N_1218,N_1214);
nor U1517 (N_1517,N_1239,N_1221);
nand U1518 (N_1518,N_1253,N_1360);
or U1519 (N_1519,N_1339,N_1310);
or U1520 (N_1520,N_1235,N_1211);
or U1521 (N_1521,N_1289,N_1371);
nor U1522 (N_1522,N_1377,N_1327);
nor U1523 (N_1523,N_1247,N_1287);
and U1524 (N_1524,N_1272,N_1203);
or U1525 (N_1525,N_1237,N_1287);
nand U1526 (N_1526,N_1324,N_1304);
nand U1527 (N_1527,N_1286,N_1358);
and U1528 (N_1528,N_1259,N_1356);
nor U1529 (N_1529,N_1235,N_1236);
nand U1530 (N_1530,N_1389,N_1396);
or U1531 (N_1531,N_1276,N_1365);
xnor U1532 (N_1532,N_1310,N_1306);
and U1533 (N_1533,N_1382,N_1381);
nor U1534 (N_1534,N_1265,N_1295);
nor U1535 (N_1535,N_1395,N_1353);
or U1536 (N_1536,N_1326,N_1207);
nand U1537 (N_1537,N_1312,N_1308);
and U1538 (N_1538,N_1239,N_1299);
nor U1539 (N_1539,N_1213,N_1282);
or U1540 (N_1540,N_1354,N_1314);
nor U1541 (N_1541,N_1379,N_1298);
or U1542 (N_1542,N_1311,N_1297);
nand U1543 (N_1543,N_1388,N_1289);
nor U1544 (N_1544,N_1353,N_1301);
nor U1545 (N_1545,N_1226,N_1249);
or U1546 (N_1546,N_1213,N_1245);
nor U1547 (N_1547,N_1251,N_1219);
nor U1548 (N_1548,N_1272,N_1229);
nor U1549 (N_1549,N_1341,N_1213);
or U1550 (N_1550,N_1399,N_1237);
and U1551 (N_1551,N_1322,N_1366);
nor U1552 (N_1552,N_1321,N_1386);
nand U1553 (N_1553,N_1396,N_1322);
nor U1554 (N_1554,N_1291,N_1316);
and U1555 (N_1555,N_1324,N_1362);
nand U1556 (N_1556,N_1229,N_1232);
nand U1557 (N_1557,N_1302,N_1392);
nand U1558 (N_1558,N_1366,N_1292);
nand U1559 (N_1559,N_1214,N_1293);
nand U1560 (N_1560,N_1219,N_1367);
or U1561 (N_1561,N_1368,N_1383);
nand U1562 (N_1562,N_1330,N_1351);
nor U1563 (N_1563,N_1396,N_1230);
and U1564 (N_1564,N_1236,N_1205);
or U1565 (N_1565,N_1392,N_1313);
nand U1566 (N_1566,N_1230,N_1213);
or U1567 (N_1567,N_1294,N_1306);
or U1568 (N_1568,N_1200,N_1276);
and U1569 (N_1569,N_1201,N_1386);
nor U1570 (N_1570,N_1216,N_1225);
and U1571 (N_1571,N_1222,N_1333);
nand U1572 (N_1572,N_1398,N_1283);
nand U1573 (N_1573,N_1239,N_1274);
and U1574 (N_1574,N_1333,N_1289);
or U1575 (N_1575,N_1213,N_1296);
nand U1576 (N_1576,N_1280,N_1259);
and U1577 (N_1577,N_1363,N_1254);
or U1578 (N_1578,N_1331,N_1289);
nor U1579 (N_1579,N_1290,N_1327);
or U1580 (N_1580,N_1228,N_1289);
nor U1581 (N_1581,N_1390,N_1347);
nand U1582 (N_1582,N_1391,N_1318);
xnor U1583 (N_1583,N_1377,N_1289);
or U1584 (N_1584,N_1367,N_1262);
nor U1585 (N_1585,N_1220,N_1200);
nand U1586 (N_1586,N_1233,N_1236);
nor U1587 (N_1587,N_1338,N_1322);
nor U1588 (N_1588,N_1211,N_1290);
or U1589 (N_1589,N_1355,N_1312);
or U1590 (N_1590,N_1327,N_1380);
nor U1591 (N_1591,N_1339,N_1236);
nor U1592 (N_1592,N_1267,N_1305);
nor U1593 (N_1593,N_1275,N_1390);
nand U1594 (N_1594,N_1212,N_1248);
and U1595 (N_1595,N_1327,N_1250);
nor U1596 (N_1596,N_1354,N_1286);
or U1597 (N_1597,N_1337,N_1225);
nor U1598 (N_1598,N_1213,N_1379);
nor U1599 (N_1599,N_1342,N_1213);
or U1600 (N_1600,N_1461,N_1400);
and U1601 (N_1601,N_1562,N_1507);
or U1602 (N_1602,N_1471,N_1596);
and U1603 (N_1603,N_1545,N_1550);
nor U1604 (N_1604,N_1558,N_1598);
and U1605 (N_1605,N_1428,N_1429);
nand U1606 (N_1606,N_1439,N_1520);
nand U1607 (N_1607,N_1423,N_1552);
or U1608 (N_1608,N_1515,N_1519);
and U1609 (N_1609,N_1453,N_1452);
nand U1610 (N_1610,N_1442,N_1402);
and U1611 (N_1611,N_1445,N_1522);
or U1612 (N_1612,N_1415,N_1409);
or U1613 (N_1613,N_1424,N_1455);
nand U1614 (N_1614,N_1525,N_1509);
and U1615 (N_1615,N_1593,N_1472);
and U1616 (N_1616,N_1494,N_1516);
and U1617 (N_1617,N_1579,N_1436);
nand U1618 (N_1618,N_1440,N_1510);
and U1619 (N_1619,N_1529,N_1430);
and U1620 (N_1620,N_1556,N_1444);
nor U1621 (N_1621,N_1569,N_1457);
nand U1622 (N_1622,N_1501,N_1567);
nor U1623 (N_1623,N_1403,N_1481);
or U1624 (N_1624,N_1437,N_1483);
nand U1625 (N_1625,N_1546,N_1575);
and U1626 (N_1626,N_1554,N_1419);
or U1627 (N_1627,N_1580,N_1502);
nand U1628 (N_1628,N_1486,N_1576);
nand U1629 (N_1629,N_1599,N_1406);
nor U1630 (N_1630,N_1427,N_1506);
nand U1631 (N_1631,N_1548,N_1584);
nand U1632 (N_1632,N_1412,N_1587);
nand U1633 (N_1633,N_1496,N_1553);
or U1634 (N_1634,N_1564,N_1470);
nand U1635 (N_1635,N_1531,N_1467);
nor U1636 (N_1636,N_1574,N_1493);
nor U1637 (N_1637,N_1508,N_1446);
or U1638 (N_1638,N_1527,N_1523);
nand U1639 (N_1639,N_1497,N_1417);
or U1640 (N_1640,N_1517,N_1513);
and U1641 (N_1641,N_1521,N_1504);
and U1642 (N_1642,N_1475,N_1434);
nand U1643 (N_1643,N_1410,N_1416);
nand U1644 (N_1644,N_1482,N_1414);
nand U1645 (N_1645,N_1592,N_1466);
nor U1646 (N_1646,N_1568,N_1500);
or U1647 (N_1647,N_1578,N_1407);
nor U1648 (N_1648,N_1449,N_1570);
and U1649 (N_1649,N_1591,N_1408);
nand U1650 (N_1650,N_1528,N_1425);
or U1651 (N_1651,N_1476,N_1418);
nand U1652 (N_1652,N_1539,N_1582);
or U1653 (N_1653,N_1480,N_1588);
and U1654 (N_1654,N_1514,N_1534);
or U1655 (N_1655,N_1478,N_1581);
and U1656 (N_1656,N_1435,N_1563);
nand U1657 (N_1657,N_1573,N_1572);
nor U1658 (N_1658,N_1485,N_1571);
nor U1659 (N_1659,N_1477,N_1469);
and U1660 (N_1660,N_1491,N_1511);
and U1661 (N_1661,N_1565,N_1538);
nor U1662 (N_1662,N_1489,N_1441);
or U1663 (N_1663,N_1464,N_1492);
nand U1664 (N_1664,N_1474,N_1585);
or U1665 (N_1665,N_1433,N_1541);
nand U1666 (N_1666,N_1454,N_1518);
and U1667 (N_1667,N_1451,N_1503);
or U1668 (N_1668,N_1560,N_1411);
nor U1669 (N_1669,N_1555,N_1490);
nand U1670 (N_1670,N_1530,N_1594);
nand U1671 (N_1671,N_1597,N_1512);
nor U1672 (N_1672,N_1577,N_1532);
nand U1673 (N_1673,N_1463,N_1404);
nand U1674 (N_1674,N_1479,N_1420);
nor U1675 (N_1675,N_1566,N_1499);
and U1676 (N_1676,N_1590,N_1465);
or U1677 (N_1677,N_1498,N_1432);
nor U1678 (N_1678,N_1450,N_1583);
and U1679 (N_1679,N_1438,N_1487);
or U1680 (N_1680,N_1524,N_1543);
nor U1681 (N_1681,N_1533,N_1405);
nand U1682 (N_1682,N_1448,N_1421);
or U1683 (N_1683,N_1413,N_1456);
and U1684 (N_1684,N_1595,N_1589);
nand U1685 (N_1685,N_1557,N_1505);
or U1686 (N_1686,N_1447,N_1458);
or U1687 (N_1687,N_1547,N_1459);
nor U1688 (N_1688,N_1422,N_1526);
and U1689 (N_1689,N_1561,N_1426);
nor U1690 (N_1690,N_1549,N_1401);
and U1691 (N_1691,N_1473,N_1535);
nand U1692 (N_1692,N_1559,N_1462);
and U1693 (N_1693,N_1537,N_1460);
nand U1694 (N_1694,N_1536,N_1586);
nor U1695 (N_1695,N_1551,N_1484);
or U1696 (N_1696,N_1443,N_1488);
or U1697 (N_1697,N_1544,N_1540);
nand U1698 (N_1698,N_1495,N_1542);
nand U1699 (N_1699,N_1468,N_1431);
nand U1700 (N_1700,N_1488,N_1571);
or U1701 (N_1701,N_1524,N_1541);
or U1702 (N_1702,N_1432,N_1534);
or U1703 (N_1703,N_1503,N_1483);
or U1704 (N_1704,N_1491,N_1400);
nor U1705 (N_1705,N_1539,N_1531);
or U1706 (N_1706,N_1470,N_1538);
and U1707 (N_1707,N_1458,N_1495);
nand U1708 (N_1708,N_1453,N_1451);
and U1709 (N_1709,N_1416,N_1456);
nand U1710 (N_1710,N_1578,N_1542);
nor U1711 (N_1711,N_1532,N_1575);
or U1712 (N_1712,N_1440,N_1590);
nor U1713 (N_1713,N_1494,N_1582);
nand U1714 (N_1714,N_1430,N_1488);
nand U1715 (N_1715,N_1442,N_1432);
nand U1716 (N_1716,N_1543,N_1408);
and U1717 (N_1717,N_1488,N_1558);
or U1718 (N_1718,N_1553,N_1513);
nand U1719 (N_1719,N_1539,N_1445);
and U1720 (N_1720,N_1512,N_1491);
and U1721 (N_1721,N_1545,N_1506);
nand U1722 (N_1722,N_1537,N_1455);
or U1723 (N_1723,N_1420,N_1591);
nand U1724 (N_1724,N_1442,N_1533);
nand U1725 (N_1725,N_1460,N_1520);
or U1726 (N_1726,N_1458,N_1570);
nor U1727 (N_1727,N_1522,N_1429);
nand U1728 (N_1728,N_1428,N_1532);
nand U1729 (N_1729,N_1406,N_1508);
nor U1730 (N_1730,N_1426,N_1493);
nand U1731 (N_1731,N_1594,N_1476);
and U1732 (N_1732,N_1474,N_1467);
nor U1733 (N_1733,N_1507,N_1423);
nand U1734 (N_1734,N_1444,N_1524);
or U1735 (N_1735,N_1453,N_1425);
or U1736 (N_1736,N_1587,N_1473);
or U1737 (N_1737,N_1405,N_1590);
and U1738 (N_1738,N_1518,N_1423);
nand U1739 (N_1739,N_1429,N_1555);
or U1740 (N_1740,N_1412,N_1526);
nor U1741 (N_1741,N_1438,N_1544);
and U1742 (N_1742,N_1504,N_1529);
and U1743 (N_1743,N_1530,N_1432);
nor U1744 (N_1744,N_1454,N_1567);
and U1745 (N_1745,N_1589,N_1482);
nand U1746 (N_1746,N_1469,N_1516);
nor U1747 (N_1747,N_1437,N_1415);
nor U1748 (N_1748,N_1447,N_1500);
or U1749 (N_1749,N_1588,N_1530);
or U1750 (N_1750,N_1579,N_1527);
nor U1751 (N_1751,N_1425,N_1581);
nor U1752 (N_1752,N_1455,N_1412);
nor U1753 (N_1753,N_1559,N_1407);
nand U1754 (N_1754,N_1582,N_1458);
nor U1755 (N_1755,N_1420,N_1423);
and U1756 (N_1756,N_1488,N_1438);
nand U1757 (N_1757,N_1565,N_1568);
or U1758 (N_1758,N_1558,N_1546);
nand U1759 (N_1759,N_1585,N_1481);
or U1760 (N_1760,N_1405,N_1443);
nand U1761 (N_1761,N_1490,N_1432);
or U1762 (N_1762,N_1414,N_1529);
nor U1763 (N_1763,N_1526,N_1507);
or U1764 (N_1764,N_1551,N_1561);
xnor U1765 (N_1765,N_1513,N_1437);
or U1766 (N_1766,N_1431,N_1420);
nand U1767 (N_1767,N_1463,N_1579);
nor U1768 (N_1768,N_1433,N_1477);
nand U1769 (N_1769,N_1551,N_1583);
and U1770 (N_1770,N_1414,N_1437);
or U1771 (N_1771,N_1544,N_1488);
or U1772 (N_1772,N_1406,N_1581);
nand U1773 (N_1773,N_1551,N_1518);
nand U1774 (N_1774,N_1545,N_1553);
and U1775 (N_1775,N_1424,N_1574);
nand U1776 (N_1776,N_1456,N_1469);
or U1777 (N_1777,N_1449,N_1460);
and U1778 (N_1778,N_1521,N_1422);
nand U1779 (N_1779,N_1553,N_1466);
xor U1780 (N_1780,N_1411,N_1444);
and U1781 (N_1781,N_1445,N_1408);
or U1782 (N_1782,N_1455,N_1540);
or U1783 (N_1783,N_1542,N_1455);
nand U1784 (N_1784,N_1508,N_1466);
nand U1785 (N_1785,N_1476,N_1539);
nand U1786 (N_1786,N_1517,N_1508);
nand U1787 (N_1787,N_1595,N_1446);
nand U1788 (N_1788,N_1543,N_1442);
nand U1789 (N_1789,N_1440,N_1428);
nor U1790 (N_1790,N_1561,N_1593);
nor U1791 (N_1791,N_1596,N_1588);
and U1792 (N_1792,N_1520,N_1425);
or U1793 (N_1793,N_1505,N_1498);
nand U1794 (N_1794,N_1422,N_1555);
and U1795 (N_1795,N_1540,N_1500);
nand U1796 (N_1796,N_1571,N_1526);
or U1797 (N_1797,N_1409,N_1438);
nand U1798 (N_1798,N_1576,N_1567);
nand U1799 (N_1799,N_1507,N_1469);
nor U1800 (N_1800,N_1771,N_1780);
nand U1801 (N_1801,N_1653,N_1714);
and U1802 (N_1802,N_1718,N_1630);
xnor U1803 (N_1803,N_1710,N_1699);
or U1804 (N_1804,N_1613,N_1761);
nand U1805 (N_1805,N_1729,N_1661);
nand U1806 (N_1806,N_1728,N_1736);
nor U1807 (N_1807,N_1788,N_1600);
nand U1808 (N_1808,N_1732,N_1787);
nor U1809 (N_1809,N_1617,N_1626);
nor U1810 (N_1810,N_1752,N_1712);
nand U1811 (N_1811,N_1755,N_1707);
nand U1812 (N_1812,N_1622,N_1620);
nor U1813 (N_1813,N_1649,N_1705);
and U1814 (N_1814,N_1621,N_1616);
or U1815 (N_1815,N_1618,N_1765);
and U1816 (N_1816,N_1686,N_1751);
nor U1817 (N_1817,N_1681,N_1656);
nor U1818 (N_1818,N_1724,N_1623);
and U1819 (N_1819,N_1773,N_1744);
nor U1820 (N_1820,N_1657,N_1655);
and U1821 (N_1821,N_1760,N_1645);
or U1822 (N_1822,N_1766,N_1665);
nand U1823 (N_1823,N_1637,N_1646);
and U1824 (N_1824,N_1745,N_1636);
or U1825 (N_1825,N_1759,N_1739);
nand U1826 (N_1826,N_1647,N_1627);
and U1827 (N_1827,N_1775,N_1722);
nand U1828 (N_1828,N_1619,N_1783);
nor U1829 (N_1829,N_1650,N_1667);
or U1830 (N_1830,N_1635,N_1682);
or U1831 (N_1831,N_1651,N_1721);
xor U1832 (N_1832,N_1689,N_1659);
or U1833 (N_1833,N_1735,N_1716);
and U1834 (N_1834,N_1691,N_1777);
nor U1835 (N_1835,N_1789,N_1678);
and U1836 (N_1836,N_1737,N_1762);
nand U1837 (N_1837,N_1606,N_1668);
or U1838 (N_1838,N_1713,N_1634);
or U1839 (N_1839,N_1676,N_1781);
or U1840 (N_1840,N_1706,N_1671);
nand U1841 (N_1841,N_1719,N_1604);
or U1842 (N_1842,N_1631,N_1612);
nand U1843 (N_1843,N_1741,N_1685);
or U1844 (N_1844,N_1652,N_1654);
nor U1845 (N_1845,N_1614,N_1750);
and U1846 (N_1846,N_1795,N_1730);
nand U1847 (N_1847,N_1723,N_1727);
nor U1848 (N_1848,N_1709,N_1605);
or U1849 (N_1849,N_1639,N_1748);
and U1850 (N_1850,N_1763,N_1694);
or U1851 (N_1851,N_1674,N_1731);
nand U1852 (N_1852,N_1749,N_1738);
and U1853 (N_1853,N_1670,N_1677);
and U1854 (N_1854,N_1640,N_1711);
nand U1855 (N_1855,N_1767,N_1740);
or U1856 (N_1856,N_1704,N_1797);
nor U1857 (N_1857,N_1798,N_1708);
or U1858 (N_1858,N_1779,N_1733);
nor U1859 (N_1859,N_1725,N_1610);
or U1860 (N_1860,N_1642,N_1663);
nand U1861 (N_1861,N_1796,N_1633);
or U1862 (N_1862,N_1785,N_1603);
nand U1863 (N_1863,N_1680,N_1611);
nor U1864 (N_1864,N_1792,N_1658);
or U1865 (N_1865,N_1743,N_1715);
nand U1866 (N_1866,N_1687,N_1764);
nand U1867 (N_1867,N_1734,N_1742);
and U1868 (N_1868,N_1688,N_1615);
nand U1869 (N_1869,N_1675,N_1754);
nor U1870 (N_1870,N_1660,N_1664);
nor U1871 (N_1871,N_1608,N_1769);
nor U1872 (N_1872,N_1628,N_1644);
and U1873 (N_1873,N_1698,N_1669);
or U1874 (N_1874,N_1692,N_1673);
nand U1875 (N_1875,N_1602,N_1747);
nand U1876 (N_1876,N_1643,N_1697);
nand U1877 (N_1877,N_1776,N_1648);
nor U1878 (N_1878,N_1786,N_1757);
and U1879 (N_1879,N_1703,N_1782);
nor U1880 (N_1880,N_1726,N_1701);
nor U1881 (N_1881,N_1629,N_1695);
or U1882 (N_1882,N_1700,N_1696);
nor U1883 (N_1883,N_1662,N_1756);
and U1884 (N_1884,N_1601,N_1632);
and U1885 (N_1885,N_1625,N_1790);
nand U1886 (N_1886,N_1638,N_1607);
and U1887 (N_1887,N_1672,N_1772);
nand U1888 (N_1888,N_1768,N_1684);
nor U1889 (N_1889,N_1784,N_1753);
nor U1890 (N_1890,N_1693,N_1758);
nor U1891 (N_1891,N_1683,N_1794);
nor U1892 (N_1892,N_1799,N_1690);
and U1893 (N_1893,N_1702,N_1770);
or U1894 (N_1894,N_1778,N_1791);
and U1895 (N_1895,N_1717,N_1666);
nor U1896 (N_1896,N_1624,N_1774);
or U1897 (N_1897,N_1641,N_1679);
nand U1898 (N_1898,N_1793,N_1609);
and U1899 (N_1899,N_1746,N_1720);
nor U1900 (N_1900,N_1779,N_1776);
nor U1901 (N_1901,N_1782,N_1629);
and U1902 (N_1902,N_1637,N_1714);
nand U1903 (N_1903,N_1665,N_1792);
nor U1904 (N_1904,N_1643,N_1645);
nor U1905 (N_1905,N_1793,N_1695);
nor U1906 (N_1906,N_1757,N_1694);
and U1907 (N_1907,N_1623,N_1683);
nand U1908 (N_1908,N_1615,N_1679);
and U1909 (N_1909,N_1668,N_1793);
or U1910 (N_1910,N_1682,N_1600);
xor U1911 (N_1911,N_1721,N_1664);
xor U1912 (N_1912,N_1729,N_1664);
or U1913 (N_1913,N_1674,N_1642);
nand U1914 (N_1914,N_1620,N_1683);
nor U1915 (N_1915,N_1753,N_1604);
nand U1916 (N_1916,N_1621,N_1768);
nand U1917 (N_1917,N_1612,N_1635);
nand U1918 (N_1918,N_1701,N_1716);
nand U1919 (N_1919,N_1769,N_1787);
and U1920 (N_1920,N_1638,N_1796);
or U1921 (N_1921,N_1666,N_1799);
nand U1922 (N_1922,N_1700,N_1662);
and U1923 (N_1923,N_1687,N_1766);
or U1924 (N_1924,N_1792,N_1661);
nor U1925 (N_1925,N_1763,N_1603);
or U1926 (N_1926,N_1616,N_1685);
nor U1927 (N_1927,N_1667,N_1793);
nand U1928 (N_1928,N_1738,N_1786);
or U1929 (N_1929,N_1623,N_1660);
and U1930 (N_1930,N_1753,N_1668);
and U1931 (N_1931,N_1693,N_1686);
nor U1932 (N_1932,N_1606,N_1730);
nor U1933 (N_1933,N_1763,N_1686);
nor U1934 (N_1934,N_1612,N_1694);
nand U1935 (N_1935,N_1666,N_1626);
xor U1936 (N_1936,N_1702,N_1736);
and U1937 (N_1937,N_1602,N_1689);
nor U1938 (N_1938,N_1659,N_1739);
and U1939 (N_1939,N_1794,N_1626);
nor U1940 (N_1940,N_1722,N_1681);
or U1941 (N_1941,N_1733,N_1681);
or U1942 (N_1942,N_1731,N_1740);
nor U1943 (N_1943,N_1630,N_1717);
or U1944 (N_1944,N_1662,N_1741);
nor U1945 (N_1945,N_1645,N_1795);
nor U1946 (N_1946,N_1623,N_1763);
or U1947 (N_1947,N_1707,N_1628);
nand U1948 (N_1948,N_1763,N_1699);
nor U1949 (N_1949,N_1611,N_1785);
or U1950 (N_1950,N_1764,N_1766);
or U1951 (N_1951,N_1788,N_1746);
or U1952 (N_1952,N_1739,N_1748);
nor U1953 (N_1953,N_1649,N_1612);
xnor U1954 (N_1954,N_1648,N_1712);
and U1955 (N_1955,N_1661,N_1659);
or U1956 (N_1956,N_1632,N_1600);
nand U1957 (N_1957,N_1678,N_1736);
nand U1958 (N_1958,N_1614,N_1782);
nor U1959 (N_1959,N_1664,N_1781);
or U1960 (N_1960,N_1689,N_1661);
nor U1961 (N_1961,N_1781,N_1752);
nand U1962 (N_1962,N_1688,N_1716);
or U1963 (N_1963,N_1654,N_1647);
nand U1964 (N_1964,N_1786,N_1645);
and U1965 (N_1965,N_1638,N_1669);
and U1966 (N_1966,N_1660,N_1765);
nor U1967 (N_1967,N_1724,N_1782);
nor U1968 (N_1968,N_1699,N_1666);
and U1969 (N_1969,N_1615,N_1721);
nand U1970 (N_1970,N_1689,N_1645);
nand U1971 (N_1971,N_1764,N_1762);
nor U1972 (N_1972,N_1783,N_1711);
nand U1973 (N_1973,N_1743,N_1777);
nand U1974 (N_1974,N_1716,N_1675);
nand U1975 (N_1975,N_1674,N_1636);
or U1976 (N_1976,N_1701,N_1689);
or U1977 (N_1977,N_1717,N_1623);
and U1978 (N_1978,N_1799,N_1727);
or U1979 (N_1979,N_1675,N_1798);
nor U1980 (N_1980,N_1628,N_1620);
or U1981 (N_1981,N_1762,N_1773);
nor U1982 (N_1982,N_1651,N_1675);
or U1983 (N_1983,N_1704,N_1798);
nor U1984 (N_1984,N_1643,N_1781);
and U1985 (N_1985,N_1764,N_1736);
and U1986 (N_1986,N_1709,N_1603);
nand U1987 (N_1987,N_1656,N_1641);
and U1988 (N_1988,N_1721,N_1717);
or U1989 (N_1989,N_1718,N_1704);
and U1990 (N_1990,N_1707,N_1702);
nor U1991 (N_1991,N_1693,N_1600);
and U1992 (N_1992,N_1743,N_1754);
and U1993 (N_1993,N_1648,N_1671);
or U1994 (N_1994,N_1718,N_1633);
nor U1995 (N_1995,N_1773,N_1622);
nor U1996 (N_1996,N_1742,N_1767);
and U1997 (N_1997,N_1627,N_1724);
nand U1998 (N_1998,N_1623,N_1732);
or U1999 (N_1999,N_1661,N_1769);
or U2000 (N_2000,N_1827,N_1900);
nand U2001 (N_2001,N_1994,N_1931);
or U2002 (N_2002,N_1853,N_1846);
nor U2003 (N_2003,N_1875,N_1842);
nor U2004 (N_2004,N_1993,N_1834);
or U2005 (N_2005,N_1992,N_1920);
or U2006 (N_2006,N_1851,N_1991);
nand U2007 (N_2007,N_1883,N_1837);
or U2008 (N_2008,N_1958,N_1823);
and U2009 (N_2009,N_1917,N_1923);
nand U2010 (N_2010,N_1813,N_1828);
xnor U2011 (N_2011,N_1873,N_1985);
nand U2012 (N_2012,N_1830,N_1806);
or U2013 (N_2013,N_1808,N_1911);
nand U2014 (N_2014,N_1858,N_1980);
nand U2015 (N_2015,N_1836,N_1871);
nand U2016 (N_2016,N_1848,N_1819);
nor U2017 (N_2017,N_1935,N_1949);
nor U2018 (N_2018,N_1930,N_1999);
or U2019 (N_2019,N_1857,N_1989);
nand U2020 (N_2020,N_1976,N_1816);
or U2021 (N_2021,N_1845,N_1972);
nor U2022 (N_2022,N_1925,N_1898);
or U2023 (N_2023,N_1805,N_1986);
nand U2024 (N_2024,N_1987,N_1859);
or U2025 (N_2025,N_1961,N_1988);
nand U2026 (N_2026,N_1855,N_1901);
or U2027 (N_2027,N_1952,N_1905);
and U2028 (N_2028,N_1894,N_1821);
or U2029 (N_2029,N_1908,N_1940);
and U2030 (N_2030,N_1983,N_1850);
or U2031 (N_2031,N_1943,N_1835);
nor U2032 (N_2032,N_1929,N_1843);
nor U2033 (N_2033,N_1945,N_1876);
nand U2034 (N_2034,N_1967,N_1918);
and U2035 (N_2035,N_1953,N_1887);
nor U2036 (N_2036,N_1960,N_1870);
nor U2037 (N_2037,N_1990,N_1979);
nor U2038 (N_2038,N_1915,N_1914);
nor U2039 (N_2039,N_1880,N_1965);
and U2040 (N_2040,N_1888,N_1825);
or U2041 (N_2041,N_1934,N_1877);
or U2042 (N_2042,N_1959,N_1854);
nand U2043 (N_2043,N_1907,N_1868);
nand U2044 (N_2044,N_1838,N_1937);
or U2045 (N_2045,N_1939,N_1897);
and U2046 (N_2046,N_1982,N_1942);
and U2047 (N_2047,N_1802,N_1924);
nand U2048 (N_2048,N_1938,N_1909);
or U2049 (N_2049,N_1866,N_1969);
nand U2050 (N_2050,N_1807,N_1973);
or U2051 (N_2051,N_1861,N_1804);
and U2052 (N_2052,N_1862,N_1885);
nand U2053 (N_2053,N_1849,N_1839);
nand U2054 (N_2054,N_1817,N_1831);
nand U2055 (N_2055,N_1893,N_1964);
or U2056 (N_2056,N_1912,N_1881);
and U2057 (N_2057,N_1882,N_1956);
nand U2058 (N_2058,N_1803,N_1978);
or U2059 (N_2059,N_1891,N_1902);
nor U2060 (N_2060,N_1832,N_1874);
and U2061 (N_2061,N_1878,N_1975);
or U2062 (N_2062,N_1998,N_1867);
and U2063 (N_2063,N_1957,N_1933);
nor U2064 (N_2064,N_1995,N_1815);
or U2065 (N_2065,N_1981,N_1922);
nand U2066 (N_2066,N_1890,N_1812);
or U2067 (N_2067,N_1904,N_1944);
or U2068 (N_2068,N_1946,N_1974);
or U2069 (N_2069,N_1954,N_1856);
and U2070 (N_2070,N_1968,N_1962);
nor U2071 (N_2071,N_1899,N_1928);
and U2072 (N_2072,N_1984,N_1970);
and U2073 (N_2073,N_1977,N_1841);
nor U2074 (N_2074,N_1864,N_1844);
nand U2075 (N_2075,N_1941,N_1936);
nand U2076 (N_2076,N_1895,N_1919);
and U2077 (N_2077,N_1860,N_1800);
or U2078 (N_2078,N_1955,N_1932);
or U2079 (N_2079,N_1996,N_1809);
nor U2080 (N_2080,N_1824,N_1829);
or U2081 (N_2081,N_1810,N_1818);
nand U2082 (N_2082,N_1801,N_1872);
and U2083 (N_2083,N_1833,N_1840);
nor U2084 (N_2084,N_1863,N_1879);
and U2085 (N_2085,N_1921,N_1910);
nor U2086 (N_2086,N_1820,N_1847);
nor U2087 (N_2087,N_1906,N_1948);
nand U2088 (N_2088,N_1826,N_1869);
and U2089 (N_2089,N_1814,N_1951);
nor U2090 (N_2090,N_1896,N_1947);
nor U2091 (N_2091,N_1926,N_1892);
nand U2092 (N_2092,N_1889,N_1884);
and U2093 (N_2093,N_1916,N_1963);
nand U2094 (N_2094,N_1822,N_1886);
and U2095 (N_2095,N_1950,N_1903);
nor U2096 (N_2096,N_1971,N_1927);
and U2097 (N_2097,N_1865,N_1811);
or U2098 (N_2098,N_1913,N_1997);
or U2099 (N_2099,N_1852,N_1966);
nand U2100 (N_2100,N_1836,N_1842);
nand U2101 (N_2101,N_1897,N_1810);
xor U2102 (N_2102,N_1971,N_1873);
or U2103 (N_2103,N_1926,N_1966);
and U2104 (N_2104,N_1806,N_1990);
nand U2105 (N_2105,N_1913,N_1839);
nor U2106 (N_2106,N_1844,N_1982);
and U2107 (N_2107,N_1961,N_1986);
and U2108 (N_2108,N_1828,N_1886);
nor U2109 (N_2109,N_1885,N_1827);
and U2110 (N_2110,N_1945,N_1993);
nor U2111 (N_2111,N_1936,N_1976);
and U2112 (N_2112,N_1867,N_1973);
nand U2113 (N_2113,N_1959,N_1953);
nand U2114 (N_2114,N_1811,N_1956);
nor U2115 (N_2115,N_1899,N_1863);
or U2116 (N_2116,N_1897,N_1969);
nand U2117 (N_2117,N_1838,N_1803);
nand U2118 (N_2118,N_1867,N_1886);
and U2119 (N_2119,N_1870,N_1935);
or U2120 (N_2120,N_1811,N_1899);
or U2121 (N_2121,N_1927,N_1963);
nor U2122 (N_2122,N_1846,N_1870);
or U2123 (N_2123,N_1859,N_1886);
nor U2124 (N_2124,N_1915,N_1868);
nand U2125 (N_2125,N_1808,N_1854);
nand U2126 (N_2126,N_1841,N_1914);
or U2127 (N_2127,N_1896,N_1900);
nand U2128 (N_2128,N_1970,N_1817);
and U2129 (N_2129,N_1982,N_1884);
nor U2130 (N_2130,N_1996,N_1984);
and U2131 (N_2131,N_1801,N_1891);
or U2132 (N_2132,N_1859,N_1835);
and U2133 (N_2133,N_1911,N_1966);
or U2134 (N_2134,N_1953,N_1983);
or U2135 (N_2135,N_1961,N_1823);
nand U2136 (N_2136,N_1846,N_1857);
and U2137 (N_2137,N_1802,N_1881);
or U2138 (N_2138,N_1843,N_1835);
and U2139 (N_2139,N_1997,N_1909);
nor U2140 (N_2140,N_1860,N_1965);
or U2141 (N_2141,N_1919,N_1974);
nand U2142 (N_2142,N_1978,N_1964);
nand U2143 (N_2143,N_1850,N_1930);
and U2144 (N_2144,N_1944,N_1892);
or U2145 (N_2145,N_1922,N_1912);
and U2146 (N_2146,N_1846,N_1877);
or U2147 (N_2147,N_1903,N_1909);
nor U2148 (N_2148,N_1829,N_1933);
nand U2149 (N_2149,N_1973,N_1910);
nand U2150 (N_2150,N_1916,N_1827);
and U2151 (N_2151,N_1813,N_1946);
or U2152 (N_2152,N_1878,N_1955);
or U2153 (N_2153,N_1952,N_1818);
nand U2154 (N_2154,N_1970,N_1916);
and U2155 (N_2155,N_1843,N_1988);
nand U2156 (N_2156,N_1868,N_1836);
and U2157 (N_2157,N_1984,N_1924);
nand U2158 (N_2158,N_1960,N_1907);
nand U2159 (N_2159,N_1917,N_1919);
nor U2160 (N_2160,N_1985,N_1910);
or U2161 (N_2161,N_1858,N_1916);
nor U2162 (N_2162,N_1815,N_1977);
nor U2163 (N_2163,N_1978,N_1868);
and U2164 (N_2164,N_1871,N_1869);
nand U2165 (N_2165,N_1949,N_1934);
nand U2166 (N_2166,N_1805,N_1994);
nand U2167 (N_2167,N_1837,N_1864);
or U2168 (N_2168,N_1887,N_1821);
nor U2169 (N_2169,N_1821,N_1923);
nor U2170 (N_2170,N_1930,N_1813);
or U2171 (N_2171,N_1876,N_1847);
and U2172 (N_2172,N_1860,N_1966);
nand U2173 (N_2173,N_1814,N_1954);
and U2174 (N_2174,N_1826,N_1955);
nand U2175 (N_2175,N_1969,N_1864);
or U2176 (N_2176,N_1808,N_1869);
or U2177 (N_2177,N_1905,N_1818);
nand U2178 (N_2178,N_1846,N_1844);
or U2179 (N_2179,N_1875,N_1996);
and U2180 (N_2180,N_1985,N_1994);
nand U2181 (N_2181,N_1823,N_1881);
or U2182 (N_2182,N_1947,N_1974);
nor U2183 (N_2183,N_1856,N_1943);
and U2184 (N_2184,N_1810,N_1830);
and U2185 (N_2185,N_1850,N_1813);
and U2186 (N_2186,N_1981,N_1976);
nand U2187 (N_2187,N_1898,N_1883);
or U2188 (N_2188,N_1988,N_1870);
and U2189 (N_2189,N_1830,N_1917);
or U2190 (N_2190,N_1944,N_1865);
or U2191 (N_2191,N_1883,N_1941);
and U2192 (N_2192,N_1894,N_1819);
and U2193 (N_2193,N_1900,N_1868);
nor U2194 (N_2194,N_1890,N_1831);
nand U2195 (N_2195,N_1985,N_1947);
nor U2196 (N_2196,N_1863,N_1819);
or U2197 (N_2197,N_1972,N_1855);
nor U2198 (N_2198,N_1898,N_1814);
and U2199 (N_2199,N_1957,N_1967);
nor U2200 (N_2200,N_2071,N_2052);
nand U2201 (N_2201,N_2032,N_2134);
nor U2202 (N_2202,N_2049,N_2054);
and U2203 (N_2203,N_2077,N_2162);
or U2204 (N_2204,N_2115,N_2069);
and U2205 (N_2205,N_2072,N_2155);
nor U2206 (N_2206,N_2031,N_2012);
nor U2207 (N_2207,N_2166,N_2004);
and U2208 (N_2208,N_2075,N_2175);
or U2209 (N_2209,N_2195,N_2177);
nor U2210 (N_2210,N_2006,N_2065);
nand U2211 (N_2211,N_2027,N_2002);
nand U2212 (N_2212,N_2157,N_2010);
nand U2213 (N_2213,N_2017,N_2122);
or U2214 (N_2214,N_2000,N_2124);
nand U2215 (N_2215,N_2185,N_2060);
nand U2216 (N_2216,N_2007,N_2139);
nand U2217 (N_2217,N_2014,N_2187);
or U2218 (N_2218,N_2154,N_2085);
and U2219 (N_2219,N_2074,N_2116);
or U2220 (N_2220,N_2148,N_2117);
nor U2221 (N_2221,N_2136,N_2090);
nor U2222 (N_2222,N_2126,N_2053);
nor U2223 (N_2223,N_2009,N_2094);
nand U2224 (N_2224,N_2184,N_2183);
nor U2225 (N_2225,N_2102,N_2013);
or U2226 (N_2226,N_2064,N_2040);
nor U2227 (N_2227,N_2062,N_2045);
nor U2228 (N_2228,N_2152,N_2035);
or U2229 (N_2229,N_2180,N_2028);
nand U2230 (N_2230,N_2005,N_2068);
nor U2231 (N_2231,N_2104,N_2147);
and U2232 (N_2232,N_2100,N_2140);
or U2233 (N_2233,N_2114,N_2137);
or U2234 (N_2234,N_2083,N_2063);
nand U2235 (N_2235,N_2112,N_2024);
or U2236 (N_2236,N_2170,N_2055);
or U2237 (N_2237,N_2101,N_2034);
nor U2238 (N_2238,N_2087,N_2194);
nand U2239 (N_2239,N_2119,N_2108);
or U2240 (N_2240,N_2086,N_2120);
nor U2241 (N_2241,N_2179,N_2176);
and U2242 (N_2242,N_2097,N_2111);
nor U2243 (N_2243,N_2172,N_2105);
and U2244 (N_2244,N_2079,N_2098);
or U2245 (N_2245,N_2149,N_2089);
nand U2246 (N_2246,N_2048,N_2159);
nor U2247 (N_2247,N_2164,N_2003);
and U2248 (N_2248,N_2036,N_2151);
or U2249 (N_2249,N_2123,N_2167);
or U2250 (N_2250,N_2093,N_2130);
and U2251 (N_2251,N_2145,N_2129);
nor U2252 (N_2252,N_2131,N_2153);
or U2253 (N_2253,N_2037,N_2171);
xor U2254 (N_2254,N_2178,N_2039);
nand U2255 (N_2255,N_2186,N_2110);
or U2256 (N_2256,N_2047,N_2189);
or U2257 (N_2257,N_2197,N_2044);
or U2258 (N_2258,N_2196,N_2011);
and U2259 (N_2259,N_2135,N_2109);
or U2260 (N_2260,N_2125,N_2141);
and U2261 (N_2261,N_2199,N_2046);
and U2262 (N_2262,N_2080,N_2160);
nand U2263 (N_2263,N_2144,N_2023);
and U2264 (N_2264,N_2066,N_2192);
and U2265 (N_2265,N_2132,N_2146);
nor U2266 (N_2266,N_2073,N_2042);
nor U2267 (N_2267,N_2051,N_2161);
or U2268 (N_2268,N_2138,N_2096);
nand U2269 (N_2269,N_2182,N_2001);
xor U2270 (N_2270,N_2084,N_2059);
nand U2271 (N_2271,N_2070,N_2067);
nand U2272 (N_2272,N_2082,N_2058);
nor U2273 (N_2273,N_2033,N_2025);
or U2274 (N_2274,N_2018,N_2015);
nand U2275 (N_2275,N_2088,N_2019);
xnor U2276 (N_2276,N_2026,N_2127);
nor U2277 (N_2277,N_2078,N_2143);
nor U2278 (N_2278,N_2165,N_2043);
nand U2279 (N_2279,N_2103,N_2022);
or U2280 (N_2280,N_2113,N_2008);
or U2281 (N_2281,N_2099,N_2188);
nor U2282 (N_2282,N_2128,N_2169);
or U2283 (N_2283,N_2163,N_2030);
nand U2284 (N_2284,N_2091,N_2156);
and U2285 (N_2285,N_2076,N_2016);
nand U2286 (N_2286,N_2158,N_2173);
and U2287 (N_2287,N_2193,N_2029);
nor U2288 (N_2288,N_2057,N_2191);
or U2289 (N_2289,N_2095,N_2118);
nor U2290 (N_2290,N_2107,N_2133);
and U2291 (N_2291,N_2061,N_2181);
nor U2292 (N_2292,N_2106,N_2038);
nand U2293 (N_2293,N_2021,N_2092);
and U2294 (N_2294,N_2198,N_2020);
nor U2295 (N_2295,N_2190,N_2121);
and U2296 (N_2296,N_2150,N_2081);
nand U2297 (N_2297,N_2050,N_2168);
nand U2298 (N_2298,N_2142,N_2174);
nand U2299 (N_2299,N_2056,N_2041);
and U2300 (N_2300,N_2095,N_2198);
and U2301 (N_2301,N_2102,N_2043);
nand U2302 (N_2302,N_2057,N_2023);
or U2303 (N_2303,N_2158,N_2136);
nor U2304 (N_2304,N_2146,N_2017);
or U2305 (N_2305,N_2001,N_2101);
nor U2306 (N_2306,N_2091,N_2041);
nand U2307 (N_2307,N_2137,N_2107);
or U2308 (N_2308,N_2065,N_2108);
and U2309 (N_2309,N_2006,N_2165);
nor U2310 (N_2310,N_2116,N_2004);
nor U2311 (N_2311,N_2037,N_2170);
nor U2312 (N_2312,N_2132,N_2030);
nand U2313 (N_2313,N_2173,N_2011);
and U2314 (N_2314,N_2148,N_2091);
or U2315 (N_2315,N_2090,N_2012);
nor U2316 (N_2316,N_2110,N_2099);
and U2317 (N_2317,N_2130,N_2097);
and U2318 (N_2318,N_2060,N_2172);
or U2319 (N_2319,N_2061,N_2008);
and U2320 (N_2320,N_2152,N_2108);
and U2321 (N_2321,N_2051,N_2180);
nand U2322 (N_2322,N_2149,N_2139);
nor U2323 (N_2323,N_2090,N_2193);
or U2324 (N_2324,N_2065,N_2083);
and U2325 (N_2325,N_2019,N_2152);
or U2326 (N_2326,N_2078,N_2135);
nand U2327 (N_2327,N_2002,N_2143);
nor U2328 (N_2328,N_2199,N_2125);
nand U2329 (N_2329,N_2198,N_2175);
nor U2330 (N_2330,N_2065,N_2070);
or U2331 (N_2331,N_2168,N_2081);
and U2332 (N_2332,N_2035,N_2018);
nand U2333 (N_2333,N_2000,N_2138);
nand U2334 (N_2334,N_2051,N_2159);
nor U2335 (N_2335,N_2140,N_2089);
nand U2336 (N_2336,N_2023,N_2139);
and U2337 (N_2337,N_2095,N_2138);
and U2338 (N_2338,N_2064,N_2098);
nor U2339 (N_2339,N_2169,N_2153);
nor U2340 (N_2340,N_2153,N_2098);
and U2341 (N_2341,N_2012,N_2057);
and U2342 (N_2342,N_2152,N_2007);
nor U2343 (N_2343,N_2151,N_2008);
or U2344 (N_2344,N_2040,N_2092);
or U2345 (N_2345,N_2049,N_2056);
and U2346 (N_2346,N_2071,N_2159);
or U2347 (N_2347,N_2148,N_2006);
nand U2348 (N_2348,N_2177,N_2080);
nand U2349 (N_2349,N_2089,N_2121);
xnor U2350 (N_2350,N_2195,N_2004);
or U2351 (N_2351,N_2131,N_2098);
and U2352 (N_2352,N_2098,N_2017);
or U2353 (N_2353,N_2080,N_2026);
nor U2354 (N_2354,N_2129,N_2103);
nor U2355 (N_2355,N_2032,N_2177);
nor U2356 (N_2356,N_2016,N_2114);
nand U2357 (N_2357,N_2021,N_2089);
nand U2358 (N_2358,N_2192,N_2136);
nor U2359 (N_2359,N_2197,N_2150);
and U2360 (N_2360,N_2141,N_2147);
or U2361 (N_2361,N_2092,N_2190);
and U2362 (N_2362,N_2102,N_2114);
and U2363 (N_2363,N_2186,N_2109);
nor U2364 (N_2364,N_2013,N_2169);
or U2365 (N_2365,N_2158,N_2111);
or U2366 (N_2366,N_2176,N_2144);
nand U2367 (N_2367,N_2104,N_2090);
and U2368 (N_2368,N_2026,N_2082);
nand U2369 (N_2369,N_2065,N_2074);
nand U2370 (N_2370,N_2161,N_2091);
nor U2371 (N_2371,N_2120,N_2154);
or U2372 (N_2372,N_2197,N_2148);
nor U2373 (N_2373,N_2032,N_2172);
nor U2374 (N_2374,N_2145,N_2086);
and U2375 (N_2375,N_2168,N_2054);
nor U2376 (N_2376,N_2050,N_2045);
or U2377 (N_2377,N_2123,N_2194);
and U2378 (N_2378,N_2174,N_2075);
and U2379 (N_2379,N_2033,N_2133);
nand U2380 (N_2380,N_2102,N_2147);
nand U2381 (N_2381,N_2009,N_2135);
nand U2382 (N_2382,N_2126,N_2035);
and U2383 (N_2383,N_2180,N_2022);
and U2384 (N_2384,N_2119,N_2127);
nand U2385 (N_2385,N_2126,N_2014);
nor U2386 (N_2386,N_2066,N_2095);
nor U2387 (N_2387,N_2019,N_2136);
or U2388 (N_2388,N_2130,N_2182);
nand U2389 (N_2389,N_2026,N_2153);
or U2390 (N_2390,N_2196,N_2155);
nor U2391 (N_2391,N_2081,N_2076);
nand U2392 (N_2392,N_2006,N_2007);
nor U2393 (N_2393,N_2170,N_2088);
nand U2394 (N_2394,N_2141,N_2026);
nor U2395 (N_2395,N_2056,N_2030);
or U2396 (N_2396,N_2163,N_2189);
nand U2397 (N_2397,N_2180,N_2191);
nand U2398 (N_2398,N_2054,N_2106);
nand U2399 (N_2399,N_2025,N_2149);
and U2400 (N_2400,N_2219,N_2375);
nand U2401 (N_2401,N_2334,N_2317);
and U2402 (N_2402,N_2276,N_2283);
nor U2403 (N_2403,N_2301,N_2343);
nand U2404 (N_2404,N_2262,N_2252);
nand U2405 (N_2405,N_2218,N_2347);
nand U2406 (N_2406,N_2309,N_2292);
nand U2407 (N_2407,N_2315,N_2399);
nand U2408 (N_2408,N_2373,N_2266);
and U2409 (N_2409,N_2378,N_2244);
nor U2410 (N_2410,N_2287,N_2392);
nand U2411 (N_2411,N_2390,N_2337);
or U2412 (N_2412,N_2277,N_2257);
and U2413 (N_2413,N_2371,N_2323);
nor U2414 (N_2414,N_2365,N_2366);
nand U2415 (N_2415,N_2318,N_2286);
and U2416 (N_2416,N_2232,N_2220);
and U2417 (N_2417,N_2224,N_2293);
nand U2418 (N_2418,N_2340,N_2226);
nor U2419 (N_2419,N_2302,N_2258);
nand U2420 (N_2420,N_2304,N_2387);
or U2421 (N_2421,N_2351,N_2289);
and U2422 (N_2422,N_2386,N_2377);
or U2423 (N_2423,N_2200,N_2327);
and U2424 (N_2424,N_2321,N_2324);
nor U2425 (N_2425,N_2269,N_2357);
or U2426 (N_2426,N_2238,N_2290);
or U2427 (N_2427,N_2355,N_2295);
nor U2428 (N_2428,N_2299,N_2354);
nor U2429 (N_2429,N_2349,N_2298);
and U2430 (N_2430,N_2336,N_2228);
or U2431 (N_2431,N_2331,N_2256);
and U2432 (N_2432,N_2381,N_2245);
nor U2433 (N_2433,N_2329,N_2367);
or U2434 (N_2434,N_2243,N_2234);
or U2435 (N_2435,N_2393,N_2388);
nor U2436 (N_2436,N_2255,N_2284);
nor U2437 (N_2437,N_2271,N_2307);
nand U2438 (N_2438,N_2344,N_2312);
nand U2439 (N_2439,N_2397,N_2207);
and U2440 (N_2440,N_2239,N_2382);
nand U2441 (N_2441,N_2254,N_2310);
xor U2442 (N_2442,N_2341,N_2303);
nor U2443 (N_2443,N_2332,N_2227);
nand U2444 (N_2444,N_2364,N_2359);
or U2445 (N_2445,N_2260,N_2396);
or U2446 (N_2446,N_2251,N_2384);
or U2447 (N_2447,N_2209,N_2350);
nand U2448 (N_2448,N_2353,N_2217);
nand U2449 (N_2449,N_2368,N_2215);
or U2450 (N_2450,N_2325,N_2230);
nor U2451 (N_2451,N_2370,N_2265);
or U2452 (N_2452,N_2237,N_2259);
nand U2453 (N_2453,N_2297,N_2389);
and U2454 (N_2454,N_2272,N_2248);
nor U2455 (N_2455,N_2246,N_2278);
nand U2456 (N_2456,N_2328,N_2316);
nand U2457 (N_2457,N_2208,N_2270);
nor U2458 (N_2458,N_2242,N_2291);
nand U2459 (N_2459,N_2204,N_2326);
or U2460 (N_2460,N_2273,N_2210);
nand U2461 (N_2461,N_2358,N_2398);
or U2462 (N_2462,N_2305,N_2372);
and U2463 (N_2463,N_2335,N_2360);
nand U2464 (N_2464,N_2300,N_2313);
nor U2465 (N_2465,N_2352,N_2333);
nor U2466 (N_2466,N_2320,N_2383);
and U2467 (N_2467,N_2342,N_2233);
and U2468 (N_2468,N_2395,N_2314);
or U2469 (N_2469,N_2240,N_2345);
or U2470 (N_2470,N_2282,N_2274);
nand U2471 (N_2471,N_2319,N_2247);
nor U2472 (N_2472,N_2202,N_2308);
xor U2473 (N_2473,N_2263,N_2213);
or U2474 (N_2474,N_2261,N_2348);
nor U2475 (N_2475,N_2267,N_2253);
nor U2476 (N_2476,N_2296,N_2264);
and U2477 (N_2477,N_2221,N_2338);
and U2478 (N_2478,N_2214,N_2369);
nor U2479 (N_2479,N_2339,N_2206);
and U2480 (N_2480,N_2288,N_2280);
nor U2481 (N_2481,N_2363,N_2212);
nor U2482 (N_2482,N_2249,N_2306);
nor U2483 (N_2483,N_2235,N_2241);
and U2484 (N_2484,N_2281,N_2391);
nor U2485 (N_2485,N_2275,N_2356);
and U2486 (N_2486,N_2361,N_2201);
nand U2487 (N_2487,N_2279,N_2379);
nor U2488 (N_2488,N_2330,N_2346);
nor U2489 (N_2489,N_2229,N_2225);
nor U2490 (N_2490,N_2216,N_2222);
nand U2491 (N_2491,N_2322,N_2362);
nand U2492 (N_2492,N_2211,N_2250);
nand U2493 (N_2493,N_2223,N_2231);
nor U2494 (N_2494,N_2236,N_2203);
and U2495 (N_2495,N_2311,N_2205);
and U2496 (N_2496,N_2380,N_2385);
nor U2497 (N_2497,N_2376,N_2374);
or U2498 (N_2498,N_2285,N_2268);
nand U2499 (N_2499,N_2394,N_2294);
or U2500 (N_2500,N_2255,N_2292);
and U2501 (N_2501,N_2257,N_2256);
nor U2502 (N_2502,N_2281,N_2353);
or U2503 (N_2503,N_2345,N_2249);
nand U2504 (N_2504,N_2205,N_2377);
nor U2505 (N_2505,N_2233,N_2399);
and U2506 (N_2506,N_2368,N_2345);
nand U2507 (N_2507,N_2349,N_2226);
and U2508 (N_2508,N_2283,N_2396);
and U2509 (N_2509,N_2243,N_2263);
nor U2510 (N_2510,N_2210,N_2395);
nand U2511 (N_2511,N_2220,N_2202);
and U2512 (N_2512,N_2359,N_2335);
or U2513 (N_2513,N_2239,N_2331);
nand U2514 (N_2514,N_2225,N_2290);
and U2515 (N_2515,N_2252,N_2214);
nand U2516 (N_2516,N_2214,N_2320);
nand U2517 (N_2517,N_2256,N_2393);
or U2518 (N_2518,N_2261,N_2286);
and U2519 (N_2519,N_2296,N_2335);
or U2520 (N_2520,N_2222,N_2368);
or U2521 (N_2521,N_2300,N_2373);
nor U2522 (N_2522,N_2275,N_2326);
nand U2523 (N_2523,N_2309,N_2382);
and U2524 (N_2524,N_2218,N_2289);
nand U2525 (N_2525,N_2302,N_2299);
nand U2526 (N_2526,N_2345,N_2372);
and U2527 (N_2527,N_2208,N_2367);
and U2528 (N_2528,N_2392,N_2250);
nor U2529 (N_2529,N_2221,N_2228);
nand U2530 (N_2530,N_2300,N_2375);
or U2531 (N_2531,N_2299,N_2233);
and U2532 (N_2532,N_2351,N_2226);
and U2533 (N_2533,N_2290,N_2276);
and U2534 (N_2534,N_2264,N_2396);
xnor U2535 (N_2535,N_2319,N_2260);
and U2536 (N_2536,N_2348,N_2383);
or U2537 (N_2537,N_2278,N_2232);
or U2538 (N_2538,N_2207,N_2218);
nor U2539 (N_2539,N_2266,N_2384);
and U2540 (N_2540,N_2366,N_2234);
nand U2541 (N_2541,N_2374,N_2266);
nor U2542 (N_2542,N_2259,N_2339);
nor U2543 (N_2543,N_2394,N_2310);
nor U2544 (N_2544,N_2200,N_2394);
or U2545 (N_2545,N_2259,N_2213);
and U2546 (N_2546,N_2318,N_2383);
or U2547 (N_2547,N_2258,N_2371);
nand U2548 (N_2548,N_2282,N_2243);
nor U2549 (N_2549,N_2258,N_2279);
nand U2550 (N_2550,N_2296,N_2237);
or U2551 (N_2551,N_2270,N_2287);
nand U2552 (N_2552,N_2313,N_2217);
xnor U2553 (N_2553,N_2314,N_2323);
and U2554 (N_2554,N_2393,N_2288);
nor U2555 (N_2555,N_2253,N_2293);
and U2556 (N_2556,N_2208,N_2218);
nor U2557 (N_2557,N_2366,N_2289);
nor U2558 (N_2558,N_2302,N_2349);
or U2559 (N_2559,N_2267,N_2207);
and U2560 (N_2560,N_2319,N_2337);
nand U2561 (N_2561,N_2226,N_2344);
or U2562 (N_2562,N_2203,N_2368);
or U2563 (N_2563,N_2245,N_2390);
nand U2564 (N_2564,N_2283,N_2240);
and U2565 (N_2565,N_2298,N_2301);
and U2566 (N_2566,N_2256,N_2341);
or U2567 (N_2567,N_2273,N_2281);
nand U2568 (N_2568,N_2203,N_2215);
or U2569 (N_2569,N_2373,N_2356);
nand U2570 (N_2570,N_2319,N_2200);
or U2571 (N_2571,N_2362,N_2252);
nand U2572 (N_2572,N_2354,N_2329);
and U2573 (N_2573,N_2252,N_2374);
nand U2574 (N_2574,N_2308,N_2312);
nor U2575 (N_2575,N_2242,N_2301);
nand U2576 (N_2576,N_2212,N_2315);
nand U2577 (N_2577,N_2204,N_2256);
nor U2578 (N_2578,N_2387,N_2282);
or U2579 (N_2579,N_2396,N_2289);
or U2580 (N_2580,N_2280,N_2245);
nor U2581 (N_2581,N_2253,N_2218);
or U2582 (N_2582,N_2367,N_2345);
or U2583 (N_2583,N_2226,N_2325);
nand U2584 (N_2584,N_2393,N_2378);
nand U2585 (N_2585,N_2374,N_2305);
nand U2586 (N_2586,N_2208,N_2220);
and U2587 (N_2587,N_2261,N_2276);
nor U2588 (N_2588,N_2291,N_2351);
and U2589 (N_2589,N_2232,N_2250);
or U2590 (N_2590,N_2244,N_2314);
and U2591 (N_2591,N_2322,N_2240);
nor U2592 (N_2592,N_2313,N_2355);
nand U2593 (N_2593,N_2303,N_2305);
nand U2594 (N_2594,N_2346,N_2303);
and U2595 (N_2595,N_2300,N_2218);
nand U2596 (N_2596,N_2356,N_2279);
and U2597 (N_2597,N_2338,N_2354);
nand U2598 (N_2598,N_2361,N_2363);
nand U2599 (N_2599,N_2315,N_2232);
nand U2600 (N_2600,N_2466,N_2502);
or U2601 (N_2601,N_2591,N_2454);
and U2602 (N_2602,N_2423,N_2575);
and U2603 (N_2603,N_2557,N_2459);
nor U2604 (N_2604,N_2536,N_2586);
nor U2605 (N_2605,N_2499,N_2553);
or U2606 (N_2606,N_2419,N_2456);
nor U2607 (N_2607,N_2426,N_2442);
nand U2608 (N_2608,N_2522,N_2547);
xor U2609 (N_2609,N_2573,N_2483);
or U2610 (N_2610,N_2560,N_2517);
nor U2611 (N_2611,N_2492,N_2519);
nor U2612 (N_2612,N_2535,N_2475);
nand U2613 (N_2613,N_2574,N_2425);
or U2614 (N_2614,N_2491,N_2411);
nor U2615 (N_2615,N_2427,N_2581);
and U2616 (N_2616,N_2452,N_2428);
nor U2617 (N_2617,N_2494,N_2448);
and U2618 (N_2618,N_2416,N_2524);
nor U2619 (N_2619,N_2417,N_2495);
nand U2620 (N_2620,N_2540,N_2430);
nor U2621 (N_2621,N_2403,N_2541);
and U2622 (N_2622,N_2420,N_2464);
or U2623 (N_2623,N_2577,N_2409);
and U2624 (N_2624,N_2538,N_2444);
or U2625 (N_2625,N_2438,N_2434);
and U2626 (N_2626,N_2482,N_2479);
xnor U2627 (N_2627,N_2408,N_2572);
nand U2628 (N_2628,N_2570,N_2555);
nor U2629 (N_2629,N_2595,N_2503);
nor U2630 (N_2630,N_2500,N_2432);
or U2631 (N_2631,N_2558,N_2515);
or U2632 (N_2632,N_2497,N_2583);
and U2633 (N_2633,N_2437,N_2549);
and U2634 (N_2634,N_2514,N_2410);
or U2635 (N_2635,N_2512,N_2488);
nand U2636 (N_2636,N_2468,N_2490);
and U2637 (N_2637,N_2436,N_2480);
and U2638 (N_2638,N_2518,N_2548);
and U2639 (N_2639,N_2477,N_2412);
nand U2640 (N_2640,N_2565,N_2506);
nand U2641 (N_2641,N_2415,N_2443);
xor U2642 (N_2642,N_2435,N_2487);
and U2643 (N_2643,N_2465,N_2441);
nand U2644 (N_2644,N_2453,N_2505);
xor U2645 (N_2645,N_2470,N_2467);
nand U2646 (N_2646,N_2401,N_2546);
and U2647 (N_2647,N_2578,N_2592);
or U2648 (N_2648,N_2478,N_2413);
and U2649 (N_2649,N_2520,N_2474);
or U2650 (N_2650,N_2461,N_2593);
nor U2651 (N_2651,N_2596,N_2588);
and U2652 (N_2652,N_2579,N_2460);
nand U2653 (N_2653,N_2537,N_2567);
and U2654 (N_2654,N_2552,N_2424);
nor U2655 (N_2655,N_2433,N_2405);
nor U2656 (N_2656,N_2406,N_2476);
nor U2657 (N_2657,N_2473,N_2599);
and U2658 (N_2658,N_2523,N_2446);
nand U2659 (N_2659,N_2559,N_2526);
nor U2660 (N_2660,N_2462,N_2528);
nor U2661 (N_2661,N_2533,N_2509);
nor U2662 (N_2662,N_2404,N_2472);
and U2663 (N_2663,N_2440,N_2511);
nand U2664 (N_2664,N_2498,N_2463);
nand U2665 (N_2665,N_2493,N_2590);
and U2666 (N_2666,N_2457,N_2584);
and U2667 (N_2667,N_2534,N_2429);
nand U2668 (N_2668,N_2585,N_2568);
nor U2669 (N_2669,N_2513,N_2484);
nand U2670 (N_2670,N_2598,N_2532);
or U2671 (N_2671,N_2407,N_2531);
or U2672 (N_2672,N_2471,N_2582);
nor U2673 (N_2673,N_2550,N_2485);
nand U2674 (N_2674,N_2496,N_2594);
and U2675 (N_2675,N_2431,N_2551);
or U2676 (N_2676,N_2402,N_2563);
nor U2677 (N_2677,N_2529,N_2580);
nor U2678 (N_2678,N_2562,N_2561);
and U2679 (N_2679,N_2508,N_2589);
nor U2680 (N_2680,N_2414,N_2489);
and U2681 (N_2681,N_2501,N_2481);
and U2682 (N_2682,N_2510,N_2544);
or U2683 (N_2683,N_2458,N_2418);
nand U2684 (N_2684,N_2525,N_2451);
nand U2685 (N_2685,N_2597,N_2554);
or U2686 (N_2686,N_2521,N_2530);
and U2687 (N_2687,N_2450,N_2587);
and U2688 (N_2688,N_2422,N_2400);
xnor U2689 (N_2689,N_2545,N_2421);
and U2690 (N_2690,N_2516,N_2449);
nand U2691 (N_2691,N_2539,N_2543);
nand U2692 (N_2692,N_2564,N_2542);
xnor U2693 (N_2693,N_2447,N_2527);
or U2694 (N_2694,N_2507,N_2445);
nand U2695 (N_2695,N_2576,N_2455);
and U2696 (N_2696,N_2439,N_2569);
and U2697 (N_2697,N_2469,N_2504);
nand U2698 (N_2698,N_2566,N_2571);
nand U2699 (N_2699,N_2556,N_2486);
nor U2700 (N_2700,N_2417,N_2472);
or U2701 (N_2701,N_2405,N_2499);
and U2702 (N_2702,N_2408,N_2516);
and U2703 (N_2703,N_2419,N_2498);
nand U2704 (N_2704,N_2482,N_2531);
xor U2705 (N_2705,N_2433,N_2596);
xnor U2706 (N_2706,N_2483,N_2499);
and U2707 (N_2707,N_2490,N_2558);
and U2708 (N_2708,N_2550,N_2522);
nand U2709 (N_2709,N_2557,N_2405);
and U2710 (N_2710,N_2449,N_2557);
and U2711 (N_2711,N_2500,N_2556);
nand U2712 (N_2712,N_2482,N_2529);
nand U2713 (N_2713,N_2491,N_2536);
nor U2714 (N_2714,N_2588,N_2556);
or U2715 (N_2715,N_2578,N_2486);
and U2716 (N_2716,N_2484,N_2540);
xnor U2717 (N_2717,N_2501,N_2559);
or U2718 (N_2718,N_2455,N_2493);
and U2719 (N_2719,N_2474,N_2504);
and U2720 (N_2720,N_2578,N_2498);
nor U2721 (N_2721,N_2500,N_2483);
nand U2722 (N_2722,N_2504,N_2412);
nand U2723 (N_2723,N_2495,N_2537);
nand U2724 (N_2724,N_2506,N_2423);
nor U2725 (N_2725,N_2513,N_2595);
nand U2726 (N_2726,N_2425,N_2575);
nand U2727 (N_2727,N_2582,N_2458);
nor U2728 (N_2728,N_2566,N_2530);
and U2729 (N_2729,N_2557,N_2453);
nor U2730 (N_2730,N_2492,N_2418);
xnor U2731 (N_2731,N_2587,N_2456);
nor U2732 (N_2732,N_2460,N_2438);
nor U2733 (N_2733,N_2539,N_2459);
nor U2734 (N_2734,N_2572,N_2414);
nand U2735 (N_2735,N_2511,N_2489);
and U2736 (N_2736,N_2446,N_2500);
nand U2737 (N_2737,N_2591,N_2471);
nand U2738 (N_2738,N_2582,N_2492);
nor U2739 (N_2739,N_2536,N_2482);
nand U2740 (N_2740,N_2460,N_2513);
nand U2741 (N_2741,N_2403,N_2408);
and U2742 (N_2742,N_2402,N_2406);
nor U2743 (N_2743,N_2525,N_2499);
or U2744 (N_2744,N_2451,N_2426);
or U2745 (N_2745,N_2552,N_2530);
nor U2746 (N_2746,N_2548,N_2457);
and U2747 (N_2747,N_2520,N_2427);
nand U2748 (N_2748,N_2539,N_2534);
or U2749 (N_2749,N_2539,N_2430);
nor U2750 (N_2750,N_2430,N_2535);
or U2751 (N_2751,N_2522,N_2444);
nand U2752 (N_2752,N_2440,N_2555);
nand U2753 (N_2753,N_2535,N_2574);
or U2754 (N_2754,N_2523,N_2558);
or U2755 (N_2755,N_2598,N_2400);
or U2756 (N_2756,N_2544,N_2445);
and U2757 (N_2757,N_2546,N_2464);
or U2758 (N_2758,N_2573,N_2531);
or U2759 (N_2759,N_2496,N_2444);
or U2760 (N_2760,N_2508,N_2497);
nor U2761 (N_2761,N_2515,N_2486);
and U2762 (N_2762,N_2439,N_2480);
and U2763 (N_2763,N_2540,N_2461);
nor U2764 (N_2764,N_2411,N_2515);
and U2765 (N_2765,N_2535,N_2488);
nor U2766 (N_2766,N_2498,N_2443);
or U2767 (N_2767,N_2403,N_2423);
or U2768 (N_2768,N_2444,N_2478);
nor U2769 (N_2769,N_2588,N_2452);
and U2770 (N_2770,N_2588,N_2413);
or U2771 (N_2771,N_2484,N_2538);
or U2772 (N_2772,N_2538,N_2498);
nand U2773 (N_2773,N_2571,N_2461);
xnor U2774 (N_2774,N_2413,N_2599);
and U2775 (N_2775,N_2564,N_2457);
nand U2776 (N_2776,N_2407,N_2446);
nor U2777 (N_2777,N_2405,N_2548);
and U2778 (N_2778,N_2463,N_2536);
or U2779 (N_2779,N_2403,N_2424);
and U2780 (N_2780,N_2518,N_2511);
nand U2781 (N_2781,N_2597,N_2568);
and U2782 (N_2782,N_2534,N_2554);
xor U2783 (N_2783,N_2507,N_2426);
nand U2784 (N_2784,N_2561,N_2596);
nand U2785 (N_2785,N_2542,N_2562);
nor U2786 (N_2786,N_2402,N_2573);
and U2787 (N_2787,N_2449,N_2456);
and U2788 (N_2788,N_2580,N_2431);
nor U2789 (N_2789,N_2408,N_2503);
nand U2790 (N_2790,N_2553,N_2564);
or U2791 (N_2791,N_2524,N_2424);
nor U2792 (N_2792,N_2440,N_2553);
and U2793 (N_2793,N_2402,N_2501);
nand U2794 (N_2794,N_2408,N_2566);
nand U2795 (N_2795,N_2494,N_2477);
nand U2796 (N_2796,N_2453,N_2419);
and U2797 (N_2797,N_2405,N_2419);
nor U2798 (N_2798,N_2547,N_2479);
nor U2799 (N_2799,N_2530,N_2562);
or U2800 (N_2800,N_2705,N_2780);
or U2801 (N_2801,N_2735,N_2785);
nand U2802 (N_2802,N_2667,N_2614);
and U2803 (N_2803,N_2606,N_2791);
nand U2804 (N_2804,N_2696,N_2744);
or U2805 (N_2805,N_2708,N_2688);
nor U2806 (N_2806,N_2710,N_2750);
or U2807 (N_2807,N_2730,N_2722);
and U2808 (N_2808,N_2761,N_2691);
nor U2809 (N_2809,N_2798,N_2641);
nand U2810 (N_2810,N_2733,N_2674);
nor U2811 (N_2811,N_2719,N_2713);
nor U2812 (N_2812,N_2771,N_2736);
and U2813 (N_2813,N_2671,N_2753);
nand U2814 (N_2814,N_2602,N_2652);
nor U2815 (N_2815,N_2712,N_2699);
and U2816 (N_2816,N_2680,N_2615);
nand U2817 (N_2817,N_2788,N_2651);
and U2818 (N_2818,N_2789,N_2677);
nor U2819 (N_2819,N_2665,N_2716);
or U2820 (N_2820,N_2635,N_2778);
nor U2821 (N_2821,N_2703,N_2768);
nor U2822 (N_2822,N_2668,N_2628);
or U2823 (N_2823,N_2757,N_2681);
nor U2824 (N_2824,N_2676,N_2756);
nand U2825 (N_2825,N_2729,N_2773);
nor U2826 (N_2826,N_2620,N_2786);
nor U2827 (N_2827,N_2654,N_2687);
or U2828 (N_2828,N_2790,N_2617);
nand U2829 (N_2829,N_2767,N_2657);
or U2830 (N_2830,N_2700,N_2772);
nor U2831 (N_2831,N_2720,N_2618);
nor U2832 (N_2832,N_2776,N_2721);
and U2833 (N_2833,N_2686,N_2679);
nor U2834 (N_2834,N_2734,N_2658);
or U2835 (N_2835,N_2707,N_2644);
nand U2836 (N_2836,N_2726,N_2782);
nand U2837 (N_2837,N_2683,N_2723);
nand U2838 (N_2838,N_2648,N_2670);
nor U2839 (N_2839,N_2653,N_2682);
nor U2840 (N_2840,N_2612,N_2797);
and U2841 (N_2841,N_2619,N_2638);
and U2842 (N_2842,N_2689,N_2784);
or U2843 (N_2843,N_2613,N_2601);
or U2844 (N_2844,N_2746,N_2792);
nor U2845 (N_2845,N_2752,N_2675);
nor U2846 (N_2846,N_2745,N_2775);
nand U2847 (N_2847,N_2603,N_2759);
or U2848 (N_2848,N_2695,N_2765);
nor U2849 (N_2849,N_2702,N_2639);
nand U2850 (N_2850,N_2728,N_2781);
nand U2851 (N_2851,N_2714,N_2770);
and U2852 (N_2852,N_2666,N_2793);
and U2853 (N_2853,N_2739,N_2701);
or U2854 (N_2854,N_2634,N_2711);
or U2855 (N_2855,N_2616,N_2685);
nor U2856 (N_2856,N_2631,N_2626);
nor U2857 (N_2857,N_2625,N_2777);
and U2858 (N_2858,N_2600,N_2662);
nor U2859 (N_2859,N_2795,N_2660);
nor U2860 (N_2860,N_2650,N_2643);
or U2861 (N_2861,N_2611,N_2632);
or U2862 (N_2862,N_2754,N_2718);
nand U2863 (N_2863,N_2655,N_2740);
or U2864 (N_2864,N_2610,N_2684);
nor U2865 (N_2865,N_2725,N_2672);
or U2866 (N_2866,N_2715,N_2694);
and U2867 (N_2867,N_2659,N_2787);
or U2868 (N_2868,N_2678,N_2697);
or U2869 (N_2869,N_2607,N_2656);
and U2870 (N_2870,N_2742,N_2647);
nor U2871 (N_2871,N_2743,N_2623);
nor U2872 (N_2872,N_2760,N_2763);
nor U2873 (N_2873,N_2766,N_2724);
nand U2874 (N_2874,N_2774,N_2755);
and U2875 (N_2875,N_2764,N_2669);
nand U2876 (N_2876,N_2796,N_2779);
nor U2877 (N_2877,N_2706,N_2629);
nand U2878 (N_2878,N_2621,N_2627);
or U2879 (N_2879,N_2633,N_2624);
nand U2880 (N_2880,N_2622,N_2642);
nor U2881 (N_2881,N_2604,N_2758);
nor U2882 (N_2882,N_2747,N_2609);
nand U2883 (N_2883,N_2762,N_2799);
nor U2884 (N_2884,N_2608,N_2645);
and U2885 (N_2885,N_2748,N_2640);
nand U2886 (N_2886,N_2646,N_2692);
nor U2887 (N_2887,N_2690,N_2704);
and U2888 (N_2888,N_2649,N_2605);
or U2889 (N_2889,N_2749,N_2741);
or U2890 (N_2890,N_2661,N_2737);
nor U2891 (N_2891,N_2717,N_2738);
nand U2892 (N_2892,N_2637,N_2731);
nand U2893 (N_2893,N_2698,N_2783);
or U2894 (N_2894,N_2636,N_2664);
nand U2895 (N_2895,N_2794,N_2663);
nor U2896 (N_2896,N_2769,N_2732);
nand U2897 (N_2897,N_2673,N_2709);
nor U2898 (N_2898,N_2751,N_2630);
and U2899 (N_2899,N_2693,N_2727);
nand U2900 (N_2900,N_2718,N_2706);
or U2901 (N_2901,N_2757,N_2645);
and U2902 (N_2902,N_2725,N_2650);
nand U2903 (N_2903,N_2764,N_2701);
and U2904 (N_2904,N_2610,N_2602);
nand U2905 (N_2905,N_2706,N_2783);
nor U2906 (N_2906,N_2715,N_2713);
nor U2907 (N_2907,N_2776,N_2727);
or U2908 (N_2908,N_2643,N_2669);
or U2909 (N_2909,N_2706,N_2716);
or U2910 (N_2910,N_2753,N_2778);
nand U2911 (N_2911,N_2625,N_2759);
nand U2912 (N_2912,N_2707,N_2608);
nand U2913 (N_2913,N_2653,N_2657);
nor U2914 (N_2914,N_2720,N_2647);
or U2915 (N_2915,N_2676,N_2746);
nor U2916 (N_2916,N_2657,N_2654);
and U2917 (N_2917,N_2794,N_2753);
and U2918 (N_2918,N_2675,N_2676);
nor U2919 (N_2919,N_2603,N_2643);
nand U2920 (N_2920,N_2767,N_2771);
nor U2921 (N_2921,N_2793,N_2696);
or U2922 (N_2922,N_2763,N_2650);
nor U2923 (N_2923,N_2776,N_2760);
nor U2924 (N_2924,N_2707,N_2795);
or U2925 (N_2925,N_2683,N_2706);
and U2926 (N_2926,N_2734,N_2748);
and U2927 (N_2927,N_2772,N_2648);
or U2928 (N_2928,N_2771,N_2703);
nand U2929 (N_2929,N_2640,N_2744);
and U2930 (N_2930,N_2706,N_2744);
nor U2931 (N_2931,N_2766,N_2709);
nand U2932 (N_2932,N_2610,N_2686);
nand U2933 (N_2933,N_2776,N_2781);
nand U2934 (N_2934,N_2642,N_2709);
or U2935 (N_2935,N_2713,N_2703);
nand U2936 (N_2936,N_2601,N_2608);
nor U2937 (N_2937,N_2687,N_2677);
and U2938 (N_2938,N_2770,N_2731);
and U2939 (N_2939,N_2663,N_2617);
or U2940 (N_2940,N_2694,N_2696);
or U2941 (N_2941,N_2678,N_2657);
nand U2942 (N_2942,N_2793,N_2769);
nor U2943 (N_2943,N_2641,N_2638);
xnor U2944 (N_2944,N_2737,N_2768);
nor U2945 (N_2945,N_2657,N_2744);
nor U2946 (N_2946,N_2693,N_2679);
or U2947 (N_2947,N_2680,N_2676);
nor U2948 (N_2948,N_2691,N_2622);
and U2949 (N_2949,N_2652,N_2604);
and U2950 (N_2950,N_2706,N_2620);
nor U2951 (N_2951,N_2793,N_2795);
nand U2952 (N_2952,N_2604,N_2686);
and U2953 (N_2953,N_2663,N_2675);
nand U2954 (N_2954,N_2647,N_2660);
nand U2955 (N_2955,N_2755,N_2791);
nand U2956 (N_2956,N_2654,N_2653);
or U2957 (N_2957,N_2722,N_2689);
nor U2958 (N_2958,N_2797,N_2715);
nor U2959 (N_2959,N_2680,N_2728);
nand U2960 (N_2960,N_2683,N_2695);
or U2961 (N_2961,N_2648,N_2693);
and U2962 (N_2962,N_2678,N_2791);
nand U2963 (N_2963,N_2797,N_2723);
nand U2964 (N_2964,N_2732,N_2621);
nor U2965 (N_2965,N_2671,N_2690);
nor U2966 (N_2966,N_2601,N_2712);
and U2967 (N_2967,N_2779,N_2616);
or U2968 (N_2968,N_2644,N_2648);
and U2969 (N_2969,N_2614,N_2631);
and U2970 (N_2970,N_2672,N_2680);
and U2971 (N_2971,N_2711,N_2620);
nand U2972 (N_2972,N_2685,N_2722);
and U2973 (N_2973,N_2745,N_2644);
nor U2974 (N_2974,N_2674,N_2644);
xor U2975 (N_2975,N_2733,N_2668);
or U2976 (N_2976,N_2679,N_2641);
and U2977 (N_2977,N_2786,N_2613);
nand U2978 (N_2978,N_2671,N_2652);
and U2979 (N_2979,N_2643,N_2756);
nor U2980 (N_2980,N_2644,N_2661);
nand U2981 (N_2981,N_2754,N_2776);
or U2982 (N_2982,N_2664,N_2735);
nand U2983 (N_2983,N_2610,N_2712);
and U2984 (N_2984,N_2723,N_2785);
nor U2985 (N_2985,N_2769,N_2643);
and U2986 (N_2986,N_2654,N_2748);
nor U2987 (N_2987,N_2783,N_2617);
nor U2988 (N_2988,N_2795,N_2724);
and U2989 (N_2989,N_2768,N_2683);
nand U2990 (N_2990,N_2727,N_2611);
or U2991 (N_2991,N_2713,N_2720);
nand U2992 (N_2992,N_2608,N_2771);
nor U2993 (N_2993,N_2743,N_2762);
nand U2994 (N_2994,N_2663,N_2768);
and U2995 (N_2995,N_2644,N_2647);
nand U2996 (N_2996,N_2694,N_2626);
nor U2997 (N_2997,N_2737,N_2784);
or U2998 (N_2998,N_2626,N_2703);
and U2999 (N_2999,N_2724,N_2698);
or U3000 (N_3000,N_2878,N_2913);
and U3001 (N_3001,N_2967,N_2999);
or U3002 (N_3002,N_2945,N_2804);
or U3003 (N_3003,N_2819,N_2901);
or U3004 (N_3004,N_2946,N_2834);
and U3005 (N_3005,N_2998,N_2889);
and U3006 (N_3006,N_2994,N_2846);
nand U3007 (N_3007,N_2848,N_2839);
and U3008 (N_3008,N_2921,N_2900);
and U3009 (N_3009,N_2873,N_2805);
nand U3010 (N_3010,N_2924,N_2898);
nand U3011 (N_3011,N_2934,N_2990);
and U3012 (N_3012,N_2983,N_2938);
or U3013 (N_3013,N_2871,N_2920);
nand U3014 (N_3014,N_2884,N_2831);
or U3015 (N_3015,N_2970,N_2858);
nor U3016 (N_3016,N_2874,N_2899);
nand U3017 (N_3017,N_2903,N_2929);
and U3018 (N_3018,N_2853,N_2830);
nand U3019 (N_3019,N_2895,N_2928);
and U3020 (N_3020,N_2815,N_2933);
and U3021 (N_3021,N_2997,N_2849);
or U3022 (N_3022,N_2947,N_2811);
nand U3023 (N_3023,N_2948,N_2965);
nor U3024 (N_3024,N_2865,N_2914);
nand U3025 (N_3025,N_2837,N_2963);
and U3026 (N_3026,N_2802,N_2918);
nor U3027 (N_3027,N_2880,N_2808);
or U3028 (N_3028,N_2940,N_2863);
or U3029 (N_3029,N_2957,N_2915);
nand U3030 (N_3030,N_2887,N_2992);
nor U3031 (N_3031,N_2866,N_2961);
nor U3032 (N_3032,N_2845,N_2800);
and U3033 (N_3033,N_2801,N_2881);
and U3034 (N_3034,N_2809,N_2959);
and U3035 (N_3035,N_2879,N_2814);
nor U3036 (N_3036,N_2876,N_2986);
and U3037 (N_3037,N_2972,N_2890);
nor U3038 (N_3038,N_2906,N_2868);
and U3039 (N_3039,N_2841,N_2955);
or U3040 (N_3040,N_2984,N_2989);
or U3041 (N_3041,N_2976,N_2888);
nor U3042 (N_3042,N_2995,N_2893);
nor U3043 (N_3043,N_2843,N_2850);
and U3044 (N_3044,N_2923,N_2882);
and U3045 (N_3045,N_2960,N_2939);
and U3046 (N_3046,N_2968,N_2877);
nor U3047 (N_3047,N_2833,N_2954);
or U3048 (N_3048,N_2859,N_2860);
or U3049 (N_3049,N_2836,N_2854);
nand U3050 (N_3050,N_2993,N_2932);
or U3051 (N_3051,N_2907,N_2813);
nand U3052 (N_3052,N_2935,N_2870);
and U3053 (N_3053,N_2991,N_2980);
nand U3054 (N_3054,N_2810,N_2971);
nand U3055 (N_3055,N_2926,N_2949);
or U3056 (N_3056,N_2807,N_2872);
and U3057 (N_3057,N_2964,N_2861);
nand U3058 (N_3058,N_2936,N_2896);
and U3059 (N_3059,N_2987,N_2827);
nor U3060 (N_3060,N_2973,N_2816);
nor U3061 (N_3061,N_2909,N_2985);
or U3062 (N_3062,N_2817,N_2996);
and U3063 (N_3063,N_2812,N_2826);
nor U3064 (N_3064,N_2922,N_2883);
nand U3065 (N_3065,N_2952,N_2891);
or U3066 (N_3066,N_2842,N_2988);
nor U3067 (N_3067,N_2803,N_2917);
nor U3068 (N_3068,N_2956,N_2885);
or U3069 (N_3069,N_2981,N_2916);
nand U3070 (N_3070,N_2902,N_2847);
nand U3071 (N_3071,N_2867,N_2840);
nor U3072 (N_3072,N_2978,N_2897);
or U3073 (N_3073,N_2886,N_2912);
nand U3074 (N_3074,N_2977,N_2966);
or U3075 (N_3075,N_2835,N_2822);
and U3076 (N_3076,N_2975,N_2828);
nor U3077 (N_3077,N_2864,N_2962);
nand U3078 (N_3078,N_2838,N_2908);
or U3079 (N_3079,N_2806,N_2910);
or U3080 (N_3080,N_2821,N_2927);
and U3081 (N_3081,N_2857,N_2911);
and U3082 (N_3082,N_2829,N_2974);
nor U3083 (N_3083,N_2925,N_2820);
nor U3084 (N_3084,N_2950,N_2937);
and U3085 (N_3085,N_2982,N_2958);
and U3086 (N_3086,N_2852,N_2851);
nand U3087 (N_3087,N_2856,N_2855);
nor U3088 (N_3088,N_2892,N_2942);
nand U3089 (N_3089,N_2943,N_2904);
and U3090 (N_3090,N_2919,N_2951);
and U3091 (N_3091,N_2862,N_2869);
and U3092 (N_3092,N_2941,N_2823);
nor U3093 (N_3093,N_2944,N_2953);
or U3094 (N_3094,N_2894,N_2832);
or U3095 (N_3095,N_2875,N_2930);
and U3096 (N_3096,N_2844,N_2818);
nor U3097 (N_3097,N_2824,N_2969);
nor U3098 (N_3098,N_2979,N_2931);
and U3099 (N_3099,N_2825,N_2905);
and U3100 (N_3100,N_2946,N_2948);
nand U3101 (N_3101,N_2939,N_2845);
and U3102 (N_3102,N_2898,N_2906);
and U3103 (N_3103,N_2824,N_2915);
nand U3104 (N_3104,N_2905,N_2971);
nand U3105 (N_3105,N_2977,N_2997);
and U3106 (N_3106,N_2857,N_2818);
nor U3107 (N_3107,N_2887,N_2980);
nand U3108 (N_3108,N_2863,N_2941);
nor U3109 (N_3109,N_2846,N_2854);
or U3110 (N_3110,N_2864,N_2800);
nand U3111 (N_3111,N_2939,N_2889);
or U3112 (N_3112,N_2938,N_2920);
or U3113 (N_3113,N_2856,N_2972);
or U3114 (N_3114,N_2835,N_2965);
or U3115 (N_3115,N_2957,N_2993);
and U3116 (N_3116,N_2992,N_2807);
nand U3117 (N_3117,N_2901,N_2842);
or U3118 (N_3118,N_2936,N_2909);
nor U3119 (N_3119,N_2872,N_2885);
nand U3120 (N_3120,N_2911,N_2979);
nor U3121 (N_3121,N_2906,N_2975);
or U3122 (N_3122,N_2907,N_2823);
nor U3123 (N_3123,N_2816,N_2852);
and U3124 (N_3124,N_2902,N_2998);
and U3125 (N_3125,N_2851,N_2857);
nor U3126 (N_3126,N_2859,N_2977);
nand U3127 (N_3127,N_2946,N_2991);
or U3128 (N_3128,N_2901,N_2923);
nor U3129 (N_3129,N_2914,N_2922);
or U3130 (N_3130,N_2985,N_2870);
and U3131 (N_3131,N_2968,N_2903);
nand U3132 (N_3132,N_2828,N_2972);
or U3133 (N_3133,N_2951,N_2895);
nand U3134 (N_3134,N_2880,N_2926);
nor U3135 (N_3135,N_2903,N_2808);
and U3136 (N_3136,N_2830,N_2937);
nor U3137 (N_3137,N_2980,N_2842);
nor U3138 (N_3138,N_2814,N_2857);
or U3139 (N_3139,N_2884,N_2969);
nand U3140 (N_3140,N_2895,N_2836);
nor U3141 (N_3141,N_2947,N_2877);
and U3142 (N_3142,N_2917,N_2925);
nand U3143 (N_3143,N_2872,N_2821);
or U3144 (N_3144,N_2889,N_2990);
and U3145 (N_3145,N_2893,N_2861);
or U3146 (N_3146,N_2984,N_2812);
nand U3147 (N_3147,N_2859,N_2995);
and U3148 (N_3148,N_2905,N_2943);
nand U3149 (N_3149,N_2861,N_2919);
and U3150 (N_3150,N_2880,N_2862);
and U3151 (N_3151,N_2903,N_2956);
and U3152 (N_3152,N_2823,N_2867);
nor U3153 (N_3153,N_2939,N_2922);
nand U3154 (N_3154,N_2986,N_2843);
and U3155 (N_3155,N_2945,N_2974);
and U3156 (N_3156,N_2868,N_2954);
and U3157 (N_3157,N_2936,N_2845);
nor U3158 (N_3158,N_2849,N_2859);
or U3159 (N_3159,N_2874,N_2971);
and U3160 (N_3160,N_2888,N_2988);
nand U3161 (N_3161,N_2983,N_2852);
nor U3162 (N_3162,N_2849,N_2893);
nand U3163 (N_3163,N_2987,N_2804);
nor U3164 (N_3164,N_2944,N_2815);
nor U3165 (N_3165,N_2942,N_2958);
and U3166 (N_3166,N_2808,N_2915);
or U3167 (N_3167,N_2874,N_2822);
nor U3168 (N_3168,N_2814,N_2846);
and U3169 (N_3169,N_2842,N_2822);
nor U3170 (N_3170,N_2968,N_2933);
nand U3171 (N_3171,N_2827,N_2894);
and U3172 (N_3172,N_2880,N_2844);
nor U3173 (N_3173,N_2897,N_2947);
and U3174 (N_3174,N_2977,N_2819);
or U3175 (N_3175,N_2918,N_2805);
and U3176 (N_3176,N_2959,N_2836);
and U3177 (N_3177,N_2879,N_2863);
nand U3178 (N_3178,N_2867,N_2934);
nand U3179 (N_3179,N_2812,N_2862);
and U3180 (N_3180,N_2812,N_2997);
and U3181 (N_3181,N_2870,N_2897);
nor U3182 (N_3182,N_2917,N_2866);
nand U3183 (N_3183,N_2947,N_2805);
or U3184 (N_3184,N_2916,N_2940);
nand U3185 (N_3185,N_2916,N_2954);
or U3186 (N_3186,N_2937,N_2817);
nand U3187 (N_3187,N_2922,N_2957);
nor U3188 (N_3188,N_2884,N_2970);
or U3189 (N_3189,N_2966,N_2847);
nor U3190 (N_3190,N_2873,N_2831);
nor U3191 (N_3191,N_2977,N_2842);
nand U3192 (N_3192,N_2917,N_2883);
and U3193 (N_3193,N_2909,N_2856);
or U3194 (N_3194,N_2971,N_2934);
or U3195 (N_3195,N_2971,N_2858);
and U3196 (N_3196,N_2970,N_2850);
nand U3197 (N_3197,N_2988,N_2953);
nand U3198 (N_3198,N_2889,N_2904);
nor U3199 (N_3199,N_2945,N_2896);
and U3200 (N_3200,N_3139,N_3005);
or U3201 (N_3201,N_3153,N_3137);
and U3202 (N_3202,N_3091,N_3051);
or U3203 (N_3203,N_3183,N_3193);
or U3204 (N_3204,N_3086,N_3092);
or U3205 (N_3205,N_3038,N_3127);
nor U3206 (N_3206,N_3022,N_3138);
nand U3207 (N_3207,N_3040,N_3088);
and U3208 (N_3208,N_3121,N_3012);
nand U3209 (N_3209,N_3105,N_3049);
or U3210 (N_3210,N_3182,N_3077);
or U3211 (N_3211,N_3039,N_3120);
nand U3212 (N_3212,N_3132,N_3177);
and U3213 (N_3213,N_3172,N_3047);
and U3214 (N_3214,N_3003,N_3028);
nand U3215 (N_3215,N_3165,N_3050);
or U3216 (N_3216,N_3016,N_3112);
or U3217 (N_3217,N_3184,N_3150);
or U3218 (N_3218,N_3128,N_3114);
nor U3219 (N_3219,N_3191,N_3011);
nand U3220 (N_3220,N_3009,N_3106);
and U3221 (N_3221,N_3111,N_3076);
or U3222 (N_3222,N_3029,N_3180);
or U3223 (N_3223,N_3010,N_3136);
or U3224 (N_3224,N_3064,N_3037);
nor U3225 (N_3225,N_3056,N_3052);
or U3226 (N_3226,N_3046,N_3164);
nand U3227 (N_3227,N_3024,N_3041);
nand U3228 (N_3228,N_3142,N_3099);
or U3229 (N_3229,N_3166,N_3162);
and U3230 (N_3230,N_3109,N_3079);
nand U3231 (N_3231,N_3084,N_3149);
or U3232 (N_3232,N_3098,N_3090);
and U3233 (N_3233,N_3093,N_3185);
and U3234 (N_3234,N_3133,N_3078);
and U3235 (N_3235,N_3071,N_3021);
nand U3236 (N_3236,N_3067,N_3030);
nand U3237 (N_3237,N_3196,N_3116);
or U3238 (N_3238,N_3036,N_3168);
and U3239 (N_3239,N_3035,N_3181);
nand U3240 (N_3240,N_3148,N_3107);
and U3241 (N_3241,N_3123,N_3042);
or U3242 (N_3242,N_3174,N_3082);
or U3243 (N_3243,N_3062,N_3134);
nor U3244 (N_3244,N_3140,N_3008);
and U3245 (N_3245,N_3048,N_3169);
nand U3246 (N_3246,N_3190,N_3043);
or U3247 (N_3247,N_3125,N_3000);
and U3248 (N_3248,N_3073,N_3130);
or U3249 (N_3249,N_3158,N_3060);
nand U3250 (N_3250,N_3186,N_3033);
nand U3251 (N_3251,N_3178,N_3108);
nor U3252 (N_3252,N_3083,N_3007);
nor U3253 (N_3253,N_3004,N_3061);
or U3254 (N_3254,N_3198,N_3194);
xor U3255 (N_3255,N_3100,N_3075);
nand U3256 (N_3256,N_3192,N_3147);
nor U3257 (N_3257,N_3163,N_3069);
and U3258 (N_3258,N_3026,N_3096);
or U3259 (N_3259,N_3159,N_3059);
and U3260 (N_3260,N_3014,N_3032);
or U3261 (N_3261,N_3188,N_3034);
and U3262 (N_3262,N_3131,N_3146);
nor U3263 (N_3263,N_3023,N_3013);
or U3264 (N_3264,N_3145,N_3101);
nor U3265 (N_3265,N_3081,N_3006);
or U3266 (N_3266,N_3160,N_3104);
nand U3267 (N_3267,N_3045,N_3066);
nor U3268 (N_3268,N_3151,N_3072);
nor U3269 (N_3269,N_3058,N_3063);
nand U3270 (N_3270,N_3141,N_3126);
or U3271 (N_3271,N_3129,N_3068);
or U3272 (N_3272,N_3017,N_3171);
nand U3273 (N_3273,N_3020,N_3094);
or U3274 (N_3274,N_3095,N_3179);
and U3275 (N_3275,N_3156,N_3117);
nand U3276 (N_3276,N_3065,N_3119);
nor U3277 (N_3277,N_3113,N_3057);
and U3278 (N_3278,N_3167,N_3176);
and U3279 (N_3279,N_3002,N_3070);
nand U3280 (N_3280,N_3097,N_3154);
nor U3281 (N_3281,N_3155,N_3025);
or U3282 (N_3282,N_3031,N_3015);
or U3283 (N_3283,N_3118,N_3199);
nand U3284 (N_3284,N_3143,N_3115);
nand U3285 (N_3285,N_3027,N_3195);
and U3286 (N_3286,N_3157,N_3124);
and U3287 (N_3287,N_3144,N_3089);
or U3288 (N_3288,N_3170,N_3074);
or U3289 (N_3289,N_3080,N_3173);
nor U3290 (N_3290,N_3018,N_3175);
or U3291 (N_3291,N_3197,N_3189);
or U3292 (N_3292,N_3087,N_3054);
and U3293 (N_3293,N_3053,N_3187);
and U3294 (N_3294,N_3103,N_3135);
or U3295 (N_3295,N_3152,N_3110);
and U3296 (N_3296,N_3085,N_3019);
nor U3297 (N_3297,N_3044,N_3122);
and U3298 (N_3298,N_3161,N_3055);
nor U3299 (N_3299,N_3001,N_3102);
nor U3300 (N_3300,N_3016,N_3170);
and U3301 (N_3301,N_3012,N_3065);
or U3302 (N_3302,N_3064,N_3130);
and U3303 (N_3303,N_3000,N_3057);
nand U3304 (N_3304,N_3146,N_3046);
and U3305 (N_3305,N_3003,N_3020);
nand U3306 (N_3306,N_3111,N_3181);
nor U3307 (N_3307,N_3096,N_3133);
and U3308 (N_3308,N_3168,N_3015);
nor U3309 (N_3309,N_3007,N_3001);
nor U3310 (N_3310,N_3037,N_3023);
or U3311 (N_3311,N_3097,N_3162);
or U3312 (N_3312,N_3105,N_3057);
or U3313 (N_3313,N_3180,N_3068);
nor U3314 (N_3314,N_3167,N_3098);
or U3315 (N_3315,N_3190,N_3114);
nor U3316 (N_3316,N_3104,N_3131);
or U3317 (N_3317,N_3002,N_3037);
nor U3318 (N_3318,N_3012,N_3006);
or U3319 (N_3319,N_3163,N_3102);
or U3320 (N_3320,N_3043,N_3052);
nor U3321 (N_3321,N_3197,N_3039);
or U3322 (N_3322,N_3018,N_3128);
and U3323 (N_3323,N_3148,N_3162);
nand U3324 (N_3324,N_3176,N_3148);
nor U3325 (N_3325,N_3158,N_3036);
and U3326 (N_3326,N_3170,N_3158);
nor U3327 (N_3327,N_3152,N_3039);
nand U3328 (N_3328,N_3137,N_3173);
and U3329 (N_3329,N_3166,N_3098);
nor U3330 (N_3330,N_3008,N_3152);
nand U3331 (N_3331,N_3151,N_3037);
and U3332 (N_3332,N_3036,N_3050);
and U3333 (N_3333,N_3105,N_3098);
or U3334 (N_3334,N_3148,N_3138);
nor U3335 (N_3335,N_3078,N_3108);
nor U3336 (N_3336,N_3181,N_3017);
nor U3337 (N_3337,N_3114,N_3055);
and U3338 (N_3338,N_3030,N_3118);
or U3339 (N_3339,N_3198,N_3019);
nand U3340 (N_3340,N_3192,N_3106);
nor U3341 (N_3341,N_3001,N_3129);
nor U3342 (N_3342,N_3002,N_3092);
nand U3343 (N_3343,N_3176,N_3073);
nor U3344 (N_3344,N_3146,N_3001);
nor U3345 (N_3345,N_3097,N_3064);
or U3346 (N_3346,N_3105,N_3028);
or U3347 (N_3347,N_3021,N_3111);
nand U3348 (N_3348,N_3115,N_3030);
and U3349 (N_3349,N_3038,N_3174);
nor U3350 (N_3350,N_3182,N_3038);
nor U3351 (N_3351,N_3056,N_3111);
and U3352 (N_3352,N_3106,N_3173);
and U3353 (N_3353,N_3176,N_3138);
nand U3354 (N_3354,N_3056,N_3151);
and U3355 (N_3355,N_3193,N_3090);
nand U3356 (N_3356,N_3022,N_3196);
nand U3357 (N_3357,N_3109,N_3029);
nand U3358 (N_3358,N_3140,N_3053);
nand U3359 (N_3359,N_3098,N_3067);
nor U3360 (N_3360,N_3169,N_3163);
and U3361 (N_3361,N_3156,N_3136);
nand U3362 (N_3362,N_3047,N_3004);
nor U3363 (N_3363,N_3139,N_3172);
nor U3364 (N_3364,N_3133,N_3153);
and U3365 (N_3365,N_3068,N_3128);
and U3366 (N_3366,N_3150,N_3019);
and U3367 (N_3367,N_3081,N_3117);
nand U3368 (N_3368,N_3197,N_3108);
nand U3369 (N_3369,N_3171,N_3151);
nand U3370 (N_3370,N_3084,N_3136);
or U3371 (N_3371,N_3060,N_3073);
or U3372 (N_3372,N_3185,N_3029);
or U3373 (N_3373,N_3136,N_3122);
nor U3374 (N_3374,N_3099,N_3063);
and U3375 (N_3375,N_3133,N_3108);
nor U3376 (N_3376,N_3163,N_3143);
nand U3377 (N_3377,N_3198,N_3148);
nand U3378 (N_3378,N_3007,N_3079);
or U3379 (N_3379,N_3189,N_3062);
nor U3380 (N_3380,N_3110,N_3083);
nand U3381 (N_3381,N_3175,N_3161);
or U3382 (N_3382,N_3124,N_3071);
or U3383 (N_3383,N_3020,N_3165);
or U3384 (N_3384,N_3163,N_3188);
nand U3385 (N_3385,N_3099,N_3122);
nand U3386 (N_3386,N_3139,N_3114);
or U3387 (N_3387,N_3115,N_3085);
nand U3388 (N_3388,N_3174,N_3052);
nand U3389 (N_3389,N_3130,N_3188);
nor U3390 (N_3390,N_3014,N_3095);
nor U3391 (N_3391,N_3141,N_3020);
or U3392 (N_3392,N_3122,N_3028);
or U3393 (N_3393,N_3151,N_3086);
or U3394 (N_3394,N_3066,N_3105);
or U3395 (N_3395,N_3130,N_3104);
nand U3396 (N_3396,N_3045,N_3026);
nand U3397 (N_3397,N_3103,N_3128);
or U3398 (N_3398,N_3073,N_3134);
nor U3399 (N_3399,N_3042,N_3031);
or U3400 (N_3400,N_3234,N_3299);
nand U3401 (N_3401,N_3227,N_3397);
and U3402 (N_3402,N_3367,N_3292);
nor U3403 (N_3403,N_3326,N_3283);
and U3404 (N_3404,N_3322,N_3310);
nor U3405 (N_3405,N_3341,N_3390);
xnor U3406 (N_3406,N_3399,N_3363);
nor U3407 (N_3407,N_3284,N_3281);
nand U3408 (N_3408,N_3383,N_3300);
nor U3409 (N_3409,N_3221,N_3231);
and U3410 (N_3410,N_3238,N_3220);
or U3411 (N_3411,N_3216,N_3286);
nand U3412 (N_3412,N_3364,N_3260);
nand U3413 (N_3413,N_3241,N_3378);
nand U3414 (N_3414,N_3393,N_3249);
nand U3415 (N_3415,N_3388,N_3314);
nor U3416 (N_3416,N_3273,N_3285);
nor U3417 (N_3417,N_3362,N_3348);
and U3418 (N_3418,N_3261,N_3291);
and U3419 (N_3419,N_3370,N_3275);
nand U3420 (N_3420,N_3208,N_3213);
and U3421 (N_3421,N_3282,N_3312);
and U3422 (N_3422,N_3204,N_3209);
and U3423 (N_3423,N_3205,N_3369);
nand U3424 (N_3424,N_3232,N_3344);
or U3425 (N_3425,N_3360,N_3379);
or U3426 (N_3426,N_3337,N_3368);
nor U3427 (N_3427,N_3254,N_3385);
or U3428 (N_3428,N_3288,N_3373);
or U3429 (N_3429,N_3214,N_3391);
or U3430 (N_3430,N_3233,N_3347);
nand U3431 (N_3431,N_3380,N_3287);
or U3432 (N_3432,N_3256,N_3382);
or U3433 (N_3433,N_3280,N_3243);
or U3434 (N_3434,N_3351,N_3219);
nand U3435 (N_3435,N_3253,N_3338);
nor U3436 (N_3436,N_3377,N_3218);
and U3437 (N_3437,N_3236,N_3257);
nand U3438 (N_3438,N_3332,N_3250);
or U3439 (N_3439,N_3255,N_3237);
nand U3440 (N_3440,N_3316,N_3398);
nand U3441 (N_3441,N_3268,N_3349);
or U3442 (N_3442,N_3251,N_3361);
nor U3443 (N_3443,N_3357,N_3392);
nand U3444 (N_3444,N_3319,N_3343);
and U3445 (N_3445,N_3200,N_3272);
nor U3446 (N_3446,N_3225,N_3230);
nor U3447 (N_3447,N_3203,N_3289);
or U3448 (N_3448,N_3323,N_3331);
nor U3449 (N_3449,N_3387,N_3222);
and U3450 (N_3450,N_3324,N_3274);
or U3451 (N_3451,N_3269,N_3226);
and U3452 (N_3452,N_3327,N_3389);
nand U3453 (N_3453,N_3352,N_3333);
or U3454 (N_3454,N_3202,N_3258);
nand U3455 (N_3455,N_3290,N_3215);
nand U3456 (N_3456,N_3358,N_3229);
and U3457 (N_3457,N_3212,N_3295);
or U3458 (N_3458,N_3293,N_3305);
nand U3459 (N_3459,N_3307,N_3320);
xor U3460 (N_3460,N_3270,N_3371);
nor U3461 (N_3461,N_3353,N_3340);
nand U3462 (N_3462,N_3223,N_3317);
or U3463 (N_3463,N_3354,N_3303);
or U3464 (N_3464,N_3381,N_3315);
and U3465 (N_3465,N_3356,N_3262);
nor U3466 (N_3466,N_3259,N_3308);
nand U3467 (N_3467,N_3395,N_3244);
nand U3468 (N_3468,N_3248,N_3345);
nand U3469 (N_3469,N_3266,N_3302);
or U3470 (N_3470,N_3365,N_3366);
or U3471 (N_3471,N_3330,N_3246);
nor U3472 (N_3472,N_3394,N_3384);
and U3473 (N_3473,N_3375,N_3206);
or U3474 (N_3474,N_3240,N_3386);
and U3475 (N_3475,N_3247,N_3328);
or U3476 (N_3476,N_3396,N_3334);
and U3477 (N_3477,N_3355,N_3325);
or U3478 (N_3478,N_3207,N_3374);
or U3479 (N_3479,N_3271,N_3228);
nor U3480 (N_3480,N_3279,N_3372);
or U3481 (N_3481,N_3306,N_3217);
or U3482 (N_3482,N_3339,N_3336);
or U3483 (N_3483,N_3294,N_3264);
nor U3484 (N_3484,N_3252,N_3263);
nand U3485 (N_3485,N_3298,N_3201);
nand U3486 (N_3486,N_3296,N_3318);
or U3487 (N_3487,N_3276,N_3342);
and U3488 (N_3488,N_3235,N_3297);
or U3489 (N_3489,N_3210,N_3304);
or U3490 (N_3490,N_3224,N_3346);
nand U3491 (N_3491,N_3350,N_3311);
or U3492 (N_3492,N_3313,N_3309);
nand U3493 (N_3493,N_3335,N_3277);
xnor U3494 (N_3494,N_3239,N_3301);
or U3495 (N_3495,N_3329,N_3211);
or U3496 (N_3496,N_3245,N_3278);
or U3497 (N_3497,N_3265,N_3359);
nor U3498 (N_3498,N_3321,N_3376);
or U3499 (N_3499,N_3242,N_3267);
and U3500 (N_3500,N_3392,N_3257);
and U3501 (N_3501,N_3303,N_3232);
and U3502 (N_3502,N_3271,N_3236);
or U3503 (N_3503,N_3310,N_3264);
nor U3504 (N_3504,N_3385,N_3259);
nor U3505 (N_3505,N_3242,N_3237);
nor U3506 (N_3506,N_3281,N_3237);
nand U3507 (N_3507,N_3320,N_3269);
nor U3508 (N_3508,N_3229,N_3363);
nor U3509 (N_3509,N_3241,N_3243);
and U3510 (N_3510,N_3380,N_3365);
nand U3511 (N_3511,N_3396,N_3257);
or U3512 (N_3512,N_3341,N_3207);
nand U3513 (N_3513,N_3397,N_3265);
nand U3514 (N_3514,N_3238,N_3305);
and U3515 (N_3515,N_3381,N_3224);
nor U3516 (N_3516,N_3325,N_3337);
nand U3517 (N_3517,N_3341,N_3365);
or U3518 (N_3518,N_3269,N_3239);
nand U3519 (N_3519,N_3312,N_3256);
nor U3520 (N_3520,N_3234,N_3276);
or U3521 (N_3521,N_3306,N_3252);
nor U3522 (N_3522,N_3235,N_3358);
and U3523 (N_3523,N_3344,N_3358);
or U3524 (N_3524,N_3304,N_3390);
and U3525 (N_3525,N_3253,N_3305);
or U3526 (N_3526,N_3306,N_3305);
and U3527 (N_3527,N_3222,N_3265);
nor U3528 (N_3528,N_3336,N_3346);
and U3529 (N_3529,N_3316,N_3308);
and U3530 (N_3530,N_3388,N_3335);
and U3531 (N_3531,N_3395,N_3316);
nor U3532 (N_3532,N_3346,N_3302);
nor U3533 (N_3533,N_3241,N_3211);
nand U3534 (N_3534,N_3287,N_3376);
and U3535 (N_3535,N_3361,N_3368);
or U3536 (N_3536,N_3323,N_3286);
nand U3537 (N_3537,N_3243,N_3317);
or U3538 (N_3538,N_3306,N_3363);
nand U3539 (N_3539,N_3294,N_3278);
or U3540 (N_3540,N_3292,N_3360);
nand U3541 (N_3541,N_3266,N_3227);
and U3542 (N_3542,N_3228,N_3247);
nand U3543 (N_3543,N_3385,N_3246);
and U3544 (N_3544,N_3380,N_3288);
and U3545 (N_3545,N_3341,N_3226);
nor U3546 (N_3546,N_3350,N_3201);
and U3547 (N_3547,N_3368,N_3349);
or U3548 (N_3548,N_3294,N_3367);
nor U3549 (N_3549,N_3340,N_3211);
nand U3550 (N_3550,N_3309,N_3266);
or U3551 (N_3551,N_3262,N_3205);
or U3552 (N_3552,N_3381,N_3333);
nand U3553 (N_3553,N_3295,N_3370);
or U3554 (N_3554,N_3272,N_3351);
and U3555 (N_3555,N_3360,N_3369);
nand U3556 (N_3556,N_3343,N_3246);
and U3557 (N_3557,N_3278,N_3220);
and U3558 (N_3558,N_3276,N_3322);
or U3559 (N_3559,N_3301,N_3204);
nor U3560 (N_3560,N_3372,N_3389);
or U3561 (N_3561,N_3258,N_3290);
nand U3562 (N_3562,N_3232,N_3397);
nand U3563 (N_3563,N_3300,N_3336);
nor U3564 (N_3564,N_3346,N_3241);
and U3565 (N_3565,N_3321,N_3237);
and U3566 (N_3566,N_3253,N_3352);
and U3567 (N_3567,N_3202,N_3237);
nor U3568 (N_3568,N_3298,N_3245);
and U3569 (N_3569,N_3308,N_3283);
nand U3570 (N_3570,N_3242,N_3286);
nand U3571 (N_3571,N_3319,N_3371);
nor U3572 (N_3572,N_3269,N_3220);
nor U3573 (N_3573,N_3225,N_3252);
nand U3574 (N_3574,N_3237,N_3315);
and U3575 (N_3575,N_3354,N_3250);
or U3576 (N_3576,N_3310,N_3375);
or U3577 (N_3577,N_3349,N_3322);
and U3578 (N_3578,N_3276,N_3317);
or U3579 (N_3579,N_3218,N_3286);
or U3580 (N_3580,N_3319,N_3375);
and U3581 (N_3581,N_3241,N_3236);
nand U3582 (N_3582,N_3246,N_3383);
and U3583 (N_3583,N_3318,N_3280);
nand U3584 (N_3584,N_3267,N_3291);
nor U3585 (N_3585,N_3204,N_3325);
nand U3586 (N_3586,N_3317,N_3389);
and U3587 (N_3587,N_3275,N_3364);
or U3588 (N_3588,N_3248,N_3237);
or U3589 (N_3589,N_3369,N_3313);
and U3590 (N_3590,N_3206,N_3347);
nor U3591 (N_3591,N_3378,N_3302);
nor U3592 (N_3592,N_3362,N_3259);
or U3593 (N_3593,N_3267,N_3215);
or U3594 (N_3594,N_3346,N_3395);
nor U3595 (N_3595,N_3348,N_3327);
nor U3596 (N_3596,N_3274,N_3353);
and U3597 (N_3597,N_3240,N_3292);
nand U3598 (N_3598,N_3329,N_3281);
or U3599 (N_3599,N_3312,N_3384);
xor U3600 (N_3600,N_3524,N_3480);
nand U3601 (N_3601,N_3527,N_3432);
and U3602 (N_3602,N_3553,N_3570);
nor U3603 (N_3603,N_3563,N_3560);
nor U3604 (N_3604,N_3405,N_3500);
xnor U3605 (N_3605,N_3593,N_3583);
and U3606 (N_3606,N_3596,N_3521);
or U3607 (N_3607,N_3562,N_3410);
or U3608 (N_3608,N_3454,N_3558);
and U3609 (N_3609,N_3417,N_3569);
nor U3610 (N_3610,N_3556,N_3574);
and U3611 (N_3611,N_3506,N_3551);
and U3612 (N_3612,N_3437,N_3494);
and U3613 (N_3613,N_3406,N_3595);
nand U3614 (N_3614,N_3585,N_3435);
or U3615 (N_3615,N_3516,N_3580);
nor U3616 (N_3616,N_3597,N_3420);
and U3617 (N_3617,N_3415,N_3490);
and U3618 (N_3618,N_3492,N_3515);
and U3619 (N_3619,N_3479,N_3470);
nand U3620 (N_3620,N_3409,N_3428);
nor U3621 (N_3621,N_3486,N_3444);
nand U3622 (N_3622,N_3443,N_3462);
nand U3623 (N_3623,N_3468,N_3557);
nand U3624 (N_3624,N_3511,N_3481);
and U3625 (N_3625,N_3588,N_3540);
nand U3626 (N_3626,N_3517,N_3416);
or U3627 (N_3627,N_3446,N_3598);
nor U3628 (N_3628,N_3451,N_3425);
nand U3629 (N_3629,N_3413,N_3449);
nor U3630 (N_3630,N_3478,N_3427);
nor U3631 (N_3631,N_3594,N_3418);
nand U3632 (N_3632,N_3421,N_3431);
nand U3633 (N_3633,N_3545,N_3441);
nor U3634 (N_3634,N_3550,N_3402);
nor U3635 (N_3635,N_3568,N_3485);
or U3636 (N_3636,N_3461,N_3457);
nand U3637 (N_3637,N_3471,N_3467);
and U3638 (N_3638,N_3549,N_3499);
or U3639 (N_3639,N_3555,N_3572);
or U3640 (N_3640,N_3571,N_3447);
or U3641 (N_3641,N_3591,N_3532);
and U3642 (N_3642,N_3534,N_3528);
nand U3643 (N_3643,N_3455,N_3541);
and U3644 (N_3644,N_3491,N_3590);
and U3645 (N_3645,N_3531,N_3484);
or U3646 (N_3646,N_3510,N_3577);
nor U3647 (N_3647,N_3452,N_3426);
nor U3648 (N_3648,N_3450,N_3404);
or U3649 (N_3649,N_3439,N_3463);
nor U3650 (N_3650,N_3448,N_3548);
nand U3651 (N_3651,N_3400,N_3543);
nor U3652 (N_3652,N_3414,N_3465);
nand U3653 (N_3653,N_3552,N_3436);
nand U3654 (N_3654,N_3561,N_3505);
and U3655 (N_3655,N_3592,N_3411);
or U3656 (N_3656,N_3483,N_3582);
nand U3657 (N_3657,N_3566,N_3498);
and U3658 (N_3658,N_3547,N_3469);
or U3659 (N_3659,N_3564,N_3488);
nor U3660 (N_3660,N_3542,N_3496);
nand U3661 (N_3661,N_3403,N_3530);
nor U3662 (N_3662,N_3520,N_3407);
nand U3663 (N_3663,N_3581,N_3523);
and U3664 (N_3664,N_3474,N_3423);
nand U3665 (N_3665,N_3573,N_3579);
or U3666 (N_3666,N_3424,N_3419);
and U3667 (N_3667,N_3473,N_3538);
and U3668 (N_3668,N_3502,N_3460);
and U3669 (N_3669,N_3578,N_3475);
nand U3670 (N_3670,N_3442,N_3453);
or U3671 (N_3671,N_3544,N_3584);
nor U3672 (N_3672,N_3476,N_3586);
nand U3673 (N_3673,N_3565,N_3587);
and U3674 (N_3674,N_3575,N_3433);
nand U3675 (N_3675,N_3599,N_3539);
nand U3676 (N_3676,N_3472,N_3493);
nor U3677 (N_3677,N_3513,N_3430);
and U3678 (N_3678,N_3401,N_3514);
or U3679 (N_3679,N_3434,N_3495);
nor U3680 (N_3680,N_3477,N_3533);
nor U3681 (N_3681,N_3466,N_3482);
or U3682 (N_3682,N_3464,N_3559);
and U3683 (N_3683,N_3489,N_3508);
nor U3684 (N_3684,N_3445,N_3509);
xnor U3685 (N_3685,N_3487,N_3567);
nand U3686 (N_3686,N_3519,N_3529);
and U3687 (N_3687,N_3507,N_3518);
or U3688 (N_3688,N_3459,N_3512);
nand U3689 (N_3689,N_3503,N_3526);
or U3690 (N_3690,N_3440,N_3501);
or U3691 (N_3691,N_3422,N_3438);
and U3692 (N_3692,N_3412,N_3497);
or U3693 (N_3693,N_3456,N_3535);
or U3694 (N_3694,N_3522,N_3576);
and U3695 (N_3695,N_3458,N_3537);
or U3696 (N_3696,N_3525,N_3408);
nand U3697 (N_3697,N_3536,N_3546);
and U3698 (N_3698,N_3589,N_3554);
nand U3699 (N_3699,N_3429,N_3504);
or U3700 (N_3700,N_3569,N_3461);
and U3701 (N_3701,N_3432,N_3474);
nand U3702 (N_3702,N_3499,N_3435);
nand U3703 (N_3703,N_3477,N_3415);
nor U3704 (N_3704,N_3446,N_3581);
nor U3705 (N_3705,N_3587,N_3454);
and U3706 (N_3706,N_3463,N_3405);
nor U3707 (N_3707,N_3556,N_3504);
and U3708 (N_3708,N_3508,N_3552);
nand U3709 (N_3709,N_3477,N_3595);
nor U3710 (N_3710,N_3482,N_3434);
and U3711 (N_3711,N_3450,N_3581);
or U3712 (N_3712,N_3500,N_3554);
or U3713 (N_3713,N_3436,N_3461);
nand U3714 (N_3714,N_3573,N_3557);
or U3715 (N_3715,N_3491,N_3563);
or U3716 (N_3716,N_3576,N_3437);
and U3717 (N_3717,N_3593,N_3465);
nor U3718 (N_3718,N_3425,N_3565);
nand U3719 (N_3719,N_3440,N_3415);
or U3720 (N_3720,N_3541,N_3596);
and U3721 (N_3721,N_3505,N_3535);
and U3722 (N_3722,N_3429,N_3572);
or U3723 (N_3723,N_3599,N_3481);
nor U3724 (N_3724,N_3506,N_3411);
and U3725 (N_3725,N_3471,N_3457);
and U3726 (N_3726,N_3541,N_3577);
nor U3727 (N_3727,N_3489,N_3444);
nor U3728 (N_3728,N_3422,N_3542);
and U3729 (N_3729,N_3424,N_3536);
and U3730 (N_3730,N_3418,N_3541);
and U3731 (N_3731,N_3488,N_3462);
and U3732 (N_3732,N_3401,N_3567);
or U3733 (N_3733,N_3517,N_3515);
nand U3734 (N_3734,N_3581,N_3448);
or U3735 (N_3735,N_3476,N_3402);
nor U3736 (N_3736,N_3599,N_3468);
or U3737 (N_3737,N_3502,N_3418);
nor U3738 (N_3738,N_3556,N_3537);
nor U3739 (N_3739,N_3596,N_3438);
or U3740 (N_3740,N_3402,N_3533);
nand U3741 (N_3741,N_3569,N_3408);
or U3742 (N_3742,N_3568,N_3403);
nor U3743 (N_3743,N_3453,N_3575);
and U3744 (N_3744,N_3588,N_3566);
or U3745 (N_3745,N_3534,N_3440);
and U3746 (N_3746,N_3404,N_3540);
and U3747 (N_3747,N_3483,N_3586);
or U3748 (N_3748,N_3528,N_3460);
or U3749 (N_3749,N_3575,N_3558);
nor U3750 (N_3750,N_3525,N_3522);
nor U3751 (N_3751,N_3486,N_3580);
nor U3752 (N_3752,N_3556,N_3596);
nor U3753 (N_3753,N_3494,N_3469);
nand U3754 (N_3754,N_3563,N_3473);
or U3755 (N_3755,N_3529,N_3575);
or U3756 (N_3756,N_3587,N_3541);
nand U3757 (N_3757,N_3438,N_3581);
or U3758 (N_3758,N_3418,N_3425);
nor U3759 (N_3759,N_3550,N_3506);
nand U3760 (N_3760,N_3567,N_3568);
or U3761 (N_3761,N_3577,N_3431);
nand U3762 (N_3762,N_3413,N_3528);
and U3763 (N_3763,N_3417,N_3412);
nand U3764 (N_3764,N_3557,N_3470);
nor U3765 (N_3765,N_3534,N_3563);
nor U3766 (N_3766,N_3490,N_3467);
nand U3767 (N_3767,N_3414,N_3501);
nand U3768 (N_3768,N_3439,N_3443);
and U3769 (N_3769,N_3570,N_3567);
or U3770 (N_3770,N_3468,N_3537);
or U3771 (N_3771,N_3456,N_3450);
nand U3772 (N_3772,N_3422,N_3423);
nor U3773 (N_3773,N_3489,N_3541);
and U3774 (N_3774,N_3548,N_3511);
nor U3775 (N_3775,N_3573,N_3495);
nand U3776 (N_3776,N_3476,N_3487);
and U3777 (N_3777,N_3403,N_3560);
or U3778 (N_3778,N_3586,N_3447);
and U3779 (N_3779,N_3550,N_3567);
nor U3780 (N_3780,N_3409,N_3478);
nor U3781 (N_3781,N_3528,N_3488);
and U3782 (N_3782,N_3430,N_3503);
or U3783 (N_3783,N_3422,N_3499);
nand U3784 (N_3784,N_3533,N_3459);
nor U3785 (N_3785,N_3441,N_3464);
nor U3786 (N_3786,N_3525,N_3419);
or U3787 (N_3787,N_3562,N_3592);
or U3788 (N_3788,N_3436,N_3468);
nor U3789 (N_3789,N_3565,N_3402);
nand U3790 (N_3790,N_3477,N_3515);
nor U3791 (N_3791,N_3515,N_3530);
xnor U3792 (N_3792,N_3502,N_3486);
nand U3793 (N_3793,N_3534,N_3465);
nor U3794 (N_3794,N_3449,N_3594);
or U3795 (N_3795,N_3588,N_3595);
nand U3796 (N_3796,N_3536,N_3472);
and U3797 (N_3797,N_3599,N_3447);
and U3798 (N_3798,N_3453,N_3464);
nor U3799 (N_3799,N_3576,N_3475);
or U3800 (N_3800,N_3626,N_3789);
and U3801 (N_3801,N_3775,N_3651);
nor U3802 (N_3802,N_3780,N_3616);
nand U3803 (N_3803,N_3613,N_3719);
and U3804 (N_3804,N_3608,N_3742);
nand U3805 (N_3805,N_3791,N_3604);
or U3806 (N_3806,N_3680,N_3729);
nand U3807 (N_3807,N_3758,N_3612);
or U3808 (N_3808,N_3618,N_3706);
nand U3809 (N_3809,N_3649,N_3761);
and U3810 (N_3810,N_3668,N_3796);
or U3811 (N_3811,N_3747,N_3624);
or U3812 (N_3812,N_3707,N_3666);
and U3813 (N_3813,N_3799,N_3783);
or U3814 (N_3814,N_3715,N_3732);
nor U3815 (N_3815,N_3756,N_3751);
or U3816 (N_3816,N_3671,N_3643);
or U3817 (N_3817,N_3743,N_3772);
and U3818 (N_3818,N_3660,N_3678);
and U3819 (N_3819,N_3632,N_3689);
or U3820 (N_3820,N_3736,N_3638);
and U3821 (N_3821,N_3645,N_3697);
and U3822 (N_3822,N_3718,N_3781);
or U3823 (N_3823,N_3641,N_3788);
or U3824 (N_3824,N_3746,N_3766);
nor U3825 (N_3825,N_3712,N_3670);
xor U3826 (N_3826,N_3723,N_3713);
nor U3827 (N_3827,N_3691,N_3739);
and U3828 (N_3828,N_3681,N_3771);
nor U3829 (N_3829,N_3669,N_3754);
or U3830 (N_3830,N_3606,N_3731);
and U3831 (N_3831,N_3720,N_3726);
or U3832 (N_3832,N_3619,N_3655);
and U3833 (N_3833,N_3777,N_3621);
nand U3834 (N_3834,N_3635,N_3665);
or U3835 (N_3835,N_3629,N_3633);
nor U3836 (N_3836,N_3711,N_3701);
or U3837 (N_3837,N_3611,N_3644);
and U3838 (N_3838,N_3709,N_3702);
nand U3839 (N_3839,N_3674,N_3762);
and U3840 (N_3840,N_3748,N_3603);
and U3841 (N_3841,N_3693,N_3763);
and U3842 (N_3842,N_3647,N_3770);
or U3843 (N_3843,N_3675,N_3708);
nand U3844 (N_3844,N_3741,N_3614);
and U3845 (N_3845,N_3740,N_3600);
or U3846 (N_3846,N_3677,N_3656);
nor U3847 (N_3847,N_3631,N_3636);
or U3848 (N_3848,N_3757,N_3653);
and U3849 (N_3849,N_3714,N_3664);
nor U3850 (N_3850,N_3735,N_3725);
xor U3851 (N_3851,N_3710,N_3690);
and U3852 (N_3852,N_3755,N_3676);
or U3853 (N_3853,N_3768,N_3778);
and U3854 (N_3854,N_3730,N_3767);
nor U3855 (N_3855,N_3695,N_3662);
or U3856 (N_3856,N_3779,N_3682);
nand U3857 (N_3857,N_3773,N_3717);
nor U3858 (N_3858,N_3672,N_3673);
or U3859 (N_3859,N_3769,N_3704);
and U3860 (N_3860,N_3745,N_3692);
nand U3861 (N_3861,N_3776,N_3721);
or U3862 (N_3862,N_3663,N_3688);
xor U3863 (N_3863,N_3733,N_3786);
nor U3864 (N_3864,N_3699,N_3684);
nor U3865 (N_3865,N_3630,N_3620);
nor U3866 (N_3866,N_3787,N_3646);
xor U3867 (N_3867,N_3795,N_3752);
or U3868 (N_3868,N_3615,N_3700);
or U3869 (N_3869,N_3683,N_3750);
or U3870 (N_3870,N_3634,N_3628);
and U3871 (N_3871,N_3765,N_3698);
or U3872 (N_3872,N_3760,N_3602);
nor U3873 (N_3873,N_3694,N_3648);
or U3874 (N_3874,N_3764,N_3744);
nor U3875 (N_3875,N_3601,N_3685);
nor U3876 (N_3876,N_3716,N_3782);
or U3877 (N_3877,N_3659,N_3790);
nand U3878 (N_3878,N_3722,N_3774);
or U3879 (N_3879,N_3679,N_3609);
or U3880 (N_3880,N_3753,N_3749);
or U3881 (N_3881,N_3797,N_3687);
or U3882 (N_3882,N_3724,N_3737);
nand U3883 (N_3883,N_3652,N_3728);
and U3884 (N_3884,N_3610,N_3658);
or U3885 (N_3885,N_3617,N_3627);
nor U3886 (N_3886,N_3759,N_3667);
nand U3887 (N_3887,N_3794,N_3640);
and U3888 (N_3888,N_3639,N_3607);
nor U3889 (N_3889,N_3661,N_3703);
nor U3890 (N_3890,N_3622,N_3727);
or U3891 (N_3891,N_3793,N_3705);
nand U3892 (N_3892,N_3792,N_3734);
nand U3893 (N_3893,N_3650,N_3605);
nor U3894 (N_3894,N_3785,N_3642);
and U3895 (N_3895,N_3784,N_3686);
and U3896 (N_3896,N_3798,N_3623);
and U3897 (N_3897,N_3625,N_3738);
or U3898 (N_3898,N_3696,N_3657);
or U3899 (N_3899,N_3637,N_3654);
nor U3900 (N_3900,N_3687,N_3762);
nor U3901 (N_3901,N_3645,N_3633);
nand U3902 (N_3902,N_3781,N_3702);
nand U3903 (N_3903,N_3720,N_3646);
and U3904 (N_3904,N_3674,N_3694);
and U3905 (N_3905,N_3710,N_3629);
nand U3906 (N_3906,N_3775,N_3612);
or U3907 (N_3907,N_3611,N_3723);
and U3908 (N_3908,N_3785,N_3658);
nor U3909 (N_3909,N_3790,N_3602);
or U3910 (N_3910,N_3607,N_3677);
and U3911 (N_3911,N_3729,N_3694);
or U3912 (N_3912,N_3660,N_3605);
nor U3913 (N_3913,N_3770,N_3652);
or U3914 (N_3914,N_3614,N_3615);
or U3915 (N_3915,N_3740,N_3657);
nand U3916 (N_3916,N_3650,N_3657);
nor U3917 (N_3917,N_3723,N_3656);
and U3918 (N_3918,N_3604,N_3615);
nand U3919 (N_3919,N_3666,N_3685);
or U3920 (N_3920,N_3749,N_3746);
or U3921 (N_3921,N_3778,N_3655);
nand U3922 (N_3922,N_3719,N_3789);
and U3923 (N_3923,N_3655,N_3613);
and U3924 (N_3924,N_3644,N_3760);
nand U3925 (N_3925,N_3620,N_3611);
and U3926 (N_3926,N_3754,N_3772);
nand U3927 (N_3927,N_3604,N_3620);
or U3928 (N_3928,N_3619,N_3688);
nor U3929 (N_3929,N_3787,N_3759);
nor U3930 (N_3930,N_3723,N_3674);
nor U3931 (N_3931,N_3655,N_3700);
nor U3932 (N_3932,N_3675,N_3663);
nand U3933 (N_3933,N_3671,N_3734);
or U3934 (N_3934,N_3661,N_3632);
and U3935 (N_3935,N_3780,N_3663);
nand U3936 (N_3936,N_3755,N_3689);
nor U3937 (N_3937,N_3631,N_3672);
and U3938 (N_3938,N_3793,N_3687);
nor U3939 (N_3939,N_3780,N_3665);
nor U3940 (N_3940,N_3743,N_3684);
and U3941 (N_3941,N_3784,N_3789);
or U3942 (N_3942,N_3743,N_3775);
and U3943 (N_3943,N_3780,N_3737);
and U3944 (N_3944,N_3642,N_3609);
or U3945 (N_3945,N_3776,N_3794);
nand U3946 (N_3946,N_3687,N_3739);
or U3947 (N_3947,N_3662,N_3663);
nand U3948 (N_3948,N_3792,N_3785);
or U3949 (N_3949,N_3693,N_3798);
nand U3950 (N_3950,N_3702,N_3608);
nor U3951 (N_3951,N_3664,N_3694);
nor U3952 (N_3952,N_3677,N_3661);
nor U3953 (N_3953,N_3718,N_3678);
nor U3954 (N_3954,N_3675,N_3672);
or U3955 (N_3955,N_3610,N_3624);
or U3956 (N_3956,N_3670,N_3757);
nor U3957 (N_3957,N_3687,N_3702);
nand U3958 (N_3958,N_3683,N_3672);
and U3959 (N_3959,N_3713,N_3621);
or U3960 (N_3960,N_3745,N_3701);
nand U3961 (N_3961,N_3764,N_3734);
nand U3962 (N_3962,N_3680,N_3688);
nor U3963 (N_3963,N_3621,N_3781);
or U3964 (N_3964,N_3603,N_3694);
or U3965 (N_3965,N_3743,N_3728);
nor U3966 (N_3966,N_3671,N_3603);
or U3967 (N_3967,N_3666,N_3739);
and U3968 (N_3968,N_3635,N_3745);
and U3969 (N_3969,N_3743,N_3742);
nand U3970 (N_3970,N_3684,N_3658);
nor U3971 (N_3971,N_3752,N_3614);
nand U3972 (N_3972,N_3673,N_3693);
nor U3973 (N_3973,N_3749,N_3725);
or U3974 (N_3974,N_3721,N_3677);
and U3975 (N_3975,N_3656,N_3716);
and U3976 (N_3976,N_3602,N_3628);
and U3977 (N_3977,N_3636,N_3628);
or U3978 (N_3978,N_3637,N_3792);
and U3979 (N_3979,N_3614,N_3700);
and U3980 (N_3980,N_3610,N_3788);
or U3981 (N_3981,N_3601,N_3705);
nor U3982 (N_3982,N_3696,N_3705);
nor U3983 (N_3983,N_3779,N_3711);
or U3984 (N_3984,N_3648,N_3701);
nand U3985 (N_3985,N_3723,N_3686);
nand U3986 (N_3986,N_3708,N_3630);
nand U3987 (N_3987,N_3622,N_3681);
or U3988 (N_3988,N_3769,N_3607);
nor U3989 (N_3989,N_3628,N_3710);
nor U3990 (N_3990,N_3725,N_3770);
nor U3991 (N_3991,N_3779,N_3628);
or U3992 (N_3992,N_3720,N_3719);
nand U3993 (N_3993,N_3693,N_3680);
nor U3994 (N_3994,N_3679,N_3766);
and U3995 (N_3995,N_3636,N_3728);
or U3996 (N_3996,N_3729,N_3754);
or U3997 (N_3997,N_3703,N_3757);
and U3998 (N_3998,N_3668,N_3679);
nor U3999 (N_3999,N_3723,N_3710);
or U4000 (N_4000,N_3979,N_3823);
and U4001 (N_4001,N_3859,N_3948);
nor U4002 (N_4002,N_3940,N_3969);
or U4003 (N_4003,N_3816,N_3885);
or U4004 (N_4004,N_3960,N_3879);
nor U4005 (N_4005,N_3873,N_3909);
nor U4006 (N_4006,N_3970,N_3901);
nand U4007 (N_4007,N_3981,N_3853);
nand U4008 (N_4008,N_3809,N_3943);
nor U4009 (N_4009,N_3972,N_3838);
or U4010 (N_4010,N_3910,N_3955);
nand U4011 (N_4011,N_3976,N_3835);
and U4012 (N_4012,N_3840,N_3937);
nand U4013 (N_4013,N_3876,N_3830);
nand U4014 (N_4014,N_3810,N_3966);
nand U4015 (N_4015,N_3867,N_3927);
nand U4016 (N_4016,N_3825,N_3914);
nor U4017 (N_4017,N_3820,N_3986);
or U4018 (N_4018,N_3984,N_3837);
or U4019 (N_4019,N_3990,N_3847);
nor U4020 (N_4020,N_3900,N_3958);
and U4021 (N_4021,N_3964,N_3921);
nor U4022 (N_4022,N_3922,N_3854);
and U4023 (N_4023,N_3860,N_3822);
nor U4024 (N_4024,N_3868,N_3991);
nor U4025 (N_4025,N_3913,N_3965);
nor U4026 (N_4026,N_3925,N_3996);
nand U4027 (N_4027,N_3973,N_3829);
nand U4028 (N_4028,N_3931,N_3875);
nand U4029 (N_4029,N_3803,N_3915);
or U4030 (N_4030,N_3999,N_3952);
nand U4031 (N_4031,N_3827,N_3811);
nand U4032 (N_4032,N_3818,N_3924);
and U4033 (N_4033,N_3890,N_3911);
nor U4034 (N_4034,N_3907,N_3850);
nor U4035 (N_4035,N_3848,N_3896);
and U4036 (N_4036,N_3845,N_3834);
and U4037 (N_4037,N_3912,N_3956);
nand U4038 (N_4038,N_3828,N_3800);
or U4039 (N_4039,N_3898,N_3985);
and U4040 (N_4040,N_3852,N_3871);
and U4041 (N_4041,N_3904,N_3886);
nor U4042 (N_4042,N_3938,N_3826);
or U4043 (N_4043,N_3814,N_3947);
or U4044 (N_4044,N_3849,N_3963);
nand U4045 (N_4045,N_3987,N_3872);
nor U4046 (N_4046,N_3950,N_3870);
nand U4047 (N_4047,N_3928,N_3988);
or U4048 (N_4048,N_3923,N_3980);
and U4049 (N_4049,N_3930,N_3968);
nor U4050 (N_4050,N_3831,N_3841);
nand U4051 (N_4051,N_3884,N_3807);
nor U4052 (N_4052,N_3926,N_3839);
nor U4053 (N_4053,N_3891,N_3864);
nor U4054 (N_4054,N_3992,N_3878);
or U4055 (N_4055,N_3869,N_3805);
nand U4056 (N_4056,N_3908,N_3857);
or U4057 (N_4057,N_3812,N_3945);
or U4058 (N_4058,N_3959,N_3978);
nand U4059 (N_4059,N_3817,N_3902);
or U4060 (N_4060,N_3865,N_3806);
nor U4061 (N_4061,N_3932,N_3842);
nor U4062 (N_4062,N_3967,N_3939);
and U4063 (N_4063,N_3974,N_3874);
nor U4064 (N_4064,N_3851,N_3862);
nand U4065 (N_4065,N_3946,N_3888);
nor U4066 (N_4066,N_3920,N_3855);
nor U4067 (N_4067,N_3929,N_3881);
nand U4068 (N_4068,N_3894,N_3905);
and U4069 (N_4069,N_3889,N_3919);
and U4070 (N_4070,N_3962,N_3802);
or U4071 (N_4071,N_3861,N_3993);
or U4072 (N_4072,N_3903,N_3844);
nand U4073 (N_4073,N_3843,N_3892);
or U4074 (N_4074,N_3877,N_3821);
nand U4075 (N_4075,N_3998,N_3935);
nor U4076 (N_4076,N_3863,N_3887);
nand U4077 (N_4077,N_3977,N_3953);
or U4078 (N_4078,N_3989,N_3858);
and U4079 (N_4079,N_3997,N_3899);
or U4080 (N_4080,N_3897,N_3895);
nand U4081 (N_4081,N_3995,N_3808);
nand U4082 (N_4082,N_3934,N_3941);
or U4083 (N_4083,N_3961,N_3880);
and U4084 (N_4084,N_3833,N_3846);
and U4085 (N_4085,N_3824,N_3975);
nor U4086 (N_4086,N_3893,N_3971);
and U4087 (N_4087,N_3856,N_3983);
or U4088 (N_4088,N_3883,N_3866);
and U4089 (N_4089,N_3949,N_3944);
nor U4090 (N_4090,N_3917,N_3957);
or U4091 (N_4091,N_3994,N_3918);
nor U4092 (N_4092,N_3804,N_3936);
nor U4093 (N_4093,N_3801,N_3951);
nand U4094 (N_4094,N_3836,N_3954);
nor U4095 (N_4095,N_3815,N_3882);
nor U4096 (N_4096,N_3942,N_3819);
nand U4097 (N_4097,N_3933,N_3906);
or U4098 (N_4098,N_3832,N_3916);
and U4099 (N_4099,N_3813,N_3982);
nor U4100 (N_4100,N_3997,N_3825);
or U4101 (N_4101,N_3883,N_3959);
nand U4102 (N_4102,N_3942,N_3883);
and U4103 (N_4103,N_3972,N_3872);
nor U4104 (N_4104,N_3980,N_3876);
nor U4105 (N_4105,N_3850,N_3909);
nor U4106 (N_4106,N_3920,N_3928);
nand U4107 (N_4107,N_3878,N_3808);
nand U4108 (N_4108,N_3881,N_3862);
nand U4109 (N_4109,N_3858,N_3840);
nor U4110 (N_4110,N_3853,N_3874);
or U4111 (N_4111,N_3970,N_3852);
nand U4112 (N_4112,N_3974,N_3906);
nand U4113 (N_4113,N_3905,N_3988);
nor U4114 (N_4114,N_3865,N_3973);
or U4115 (N_4115,N_3837,N_3951);
nor U4116 (N_4116,N_3838,N_3863);
nand U4117 (N_4117,N_3944,N_3979);
nor U4118 (N_4118,N_3970,N_3952);
nand U4119 (N_4119,N_3981,N_3868);
or U4120 (N_4120,N_3859,N_3944);
or U4121 (N_4121,N_3804,N_3923);
and U4122 (N_4122,N_3908,N_3830);
or U4123 (N_4123,N_3945,N_3883);
nand U4124 (N_4124,N_3892,N_3967);
and U4125 (N_4125,N_3850,N_3851);
nand U4126 (N_4126,N_3893,N_3866);
nand U4127 (N_4127,N_3872,N_3852);
nand U4128 (N_4128,N_3950,N_3906);
and U4129 (N_4129,N_3938,N_3835);
or U4130 (N_4130,N_3897,N_3870);
and U4131 (N_4131,N_3826,N_3967);
or U4132 (N_4132,N_3961,N_3819);
or U4133 (N_4133,N_3948,N_3997);
nor U4134 (N_4134,N_3815,N_3952);
and U4135 (N_4135,N_3827,N_3890);
or U4136 (N_4136,N_3972,N_3869);
or U4137 (N_4137,N_3816,N_3958);
nand U4138 (N_4138,N_3912,N_3892);
and U4139 (N_4139,N_3930,N_3960);
or U4140 (N_4140,N_3899,N_3946);
nor U4141 (N_4141,N_3943,N_3933);
or U4142 (N_4142,N_3880,N_3869);
and U4143 (N_4143,N_3814,N_3820);
nor U4144 (N_4144,N_3963,N_3848);
nor U4145 (N_4145,N_3947,N_3839);
or U4146 (N_4146,N_3984,N_3862);
or U4147 (N_4147,N_3985,N_3855);
or U4148 (N_4148,N_3828,N_3832);
nand U4149 (N_4149,N_3900,N_3804);
or U4150 (N_4150,N_3835,N_3940);
nor U4151 (N_4151,N_3956,N_3944);
or U4152 (N_4152,N_3867,N_3803);
and U4153 (N_4153,N_3924,N_3917);
nand U4154 (N_4154,N_3844,N_3873);
nand U4155 (N_4155,N_3918,N_3839);
nand U4156 (N_4156,N_3913,N_3993);
and U4157 (N_4157,N_3982,N_3930);
nand U4158 (N_4158,N_3980,N_3868);
nor U4159 (N_4159,N_3846,N_3931);
nand U4160 (N_4160,N_3855,N_3947);
nor U4161 (N_4161,N_3972,N_3997);
and U4162 (N_4162,N_3842,N_3821);
nor U4163 (N_4163,N_3972,N_3904);
and U4164 (N_4164,N_3896,N_3814);
nand U4165 (N_4165,N_3978,N_3852);
nand U4166 (N_4166,N_3963,N_3807);
nor U4167 (N_4167,N_3937,N_3964);
or U4168 (N_4168,N_3908,N_3823);
nor U4169 (N_4169,N_3977,N_3817);
or U4170 (N_4170,N_3873,N_3849);
nor U4171 (N_4171,N_3868,N_3946);
nor U4172 (N_4172,N_3825,N_3872);
nand U4173 (N_4173,N_3830,N_3870);
and U4174 (N_4174,N_3934,N_3833);
nor U4175 (N_4175,N_3801,N_3800);
or U4176 (N_4176,N_3931,N_3993);
or U4177 (N_4177,N_3916,N_3882);
and U4178 (N_4178,N_3948,N_3888);
and U4179 (N_4179,N_3866,N_3834);
nand U4180 (N_4180,N_3878,N_3930);
nand U4181 (N_4181,N_3915,N_3983);
nor U4182 (N_4182,N_3832,N_3837);
nor U4183 (N_4183,N_3912,N_3993);
nand U4184 (N_4184,N_3968,N_3986);
and U4185 (N_4185,N_3810,N_3814);
nor U4186 (N_4186,N_3985,N_3938);
nand U4187 (N_4187,N_3930,N_3860);
and U4188 (N_4188,N_3869,N_3930);
nor U4189 (N_4189,N_3946,N_3852);
or U4190 (N_4190,N_3843,N_3997);
or U4191 (N_4191,N_3817,N_3863);
and U4192 (N_4192,N_3958,N_3835);
or U4193 (N_4193,N_3930,N_3996);
nor U4194 (N_4194,N_3816,N_3897);
and U4195 (N_4195,N_3957,N_3843);
and U4196 (N_4196,N_3997,N_3815);
nor U4197 (N_4197,N_3944,N_3933);
nand U4198 (N_4198,N_3892,N_3822);
and U4199 (N_4199,N_3948,N_3850);
nand U4200 (N_4200,N_4183,N_4153);
nor U4201 (N_4201,N_4036,N_4107);
and U4202 (N_4202,N_4021,N_4101);
or U4203 (N_4203,N_4134,N_4074);
and U4204 (N_4204,N_4009,N_4067);
nor U4205 (N_4205,N_4185,N_4022);
nand U4206 (N_4206,N_4156,N_4033);
or U4207 (N_4207,N_4092,N_4015);
and U4208 (N_4208,N_4179,N_4146);
or U4209 (N_4209,N_4094,N_4106);
and U4210 (N_4210,N_4041,N_4042);
or U4211 (N_4211,N_4023,N_4173);
nor U4212 (N_4212,N_4068,N_4006);
nand U4213 (N_4213,N_4091,N_4027);
or U4214 (N_4214,N_4145,N_4010);
nand U4215 (N_4215,N_4054,N_4029);
and U4216 (N_4216,N_4181,N_4082);
nor U4217 (N_4217,N_4063,N_4051);
and U4218 (N_4218,N_4114,N_4062);
nand U4219 (N_4219,N_4127,N_4165);
or U4220 (N_4220,N_4119,N_4017);
and U4221 (N_4221,N_4157,N_4047);
nor U4222 (N_4222,N_4132,N_4138);
nor U4223 (N_4223,N_4144,N_4086);
nor U4224 (N_4224,N_4169,N_4171);
or U4225 (N_4225,N_4123,N_4085);
or U4226 (N_4226,N_4131,N_4161);
nand U4227 (N_4227,N_4105,N_4071);
nor U4228 (N_4228,N_4170,N_4053);
nand U4229 (N_4229,N_4172,N_4155);
nor U4230 (N_4230,N_4058,N_4007);
and U4231 (N_4231,N_4166,N_4037);
nor U4232 (N_4232,N_4180,N_4003);
nand U4233 (N_4233,N_4059,N_4126);
nor U4234 (N_4234,N_4141,N_4028);
and U4235 (N_4235,N_4096,N_4040);
and U4236 (N_4236,N_4133,N_4100);
and U4237 (N_4237,N_4113,N_4046);
nand U4238 (N_4238,N_4081,N_4176);
nor U4239 (N_4239,N_4137,N_4075);
nor U4240 (N_4240,N_4044,N_4135);
and U4241 (N_4241,N_4110,N_4035);
nor U4242 (N_4242,N_4108,N_4178);
nor U4243 (N_4243,N_4103,N_4012);
and U4244 (N_4244,N_4192,N_4056);
and U4245 (N_4245,N_4025,N_4060);
or U4246 (N_4246,N_4152,N_4089);
or U4247 (N_4247,N_4147,N_4043);
or U4248 (N_4248,N_4158,N_4194);
nand U4249 (N_4249,N_4079,N_4013);
and U4250 (N_4250,N_4039,N_4129);
nor U4251 (N_4251,N_4118,N_4032);
or U4252 (N_4252,N_4088,N_4014);
nand U4253 (N_4253,N_4130,N_4049);
or U4254 (N_4254,N_4045,N_4050);
or U4255 (N_4255,N_4143,N_4177);
or U4256 (N_4256,N_4190,N_4154);
or U4257 (N_4257,N_4084,N_4182);
nand U4258 (N_4258,N_4034,N_4184);
and U4259 (N_4259,N_4159,N_4095);
xor U4260 (N_4260,N_4191,N_4073);
nand U4261 (N_4261,N_4164,N_4199);
and U4262 (N_4262,N_4112,N_4188);
and U4263 (N_4263,N_4055,N_4160);
or U4264 (N_4264,N_4030,N_4061);
or U4265 (N_4265,N_4000,N_4162);
nor U4266 (N_4266,N_4052,N_4139);
or U4267 (N_4267,N_4142,N_4186);
nor U4268 (N_4268,N_4002,N_4115);
or U4269 (N_4269,N_4093,N_4168);
and U4270 (N_4270,N_4163,N_4128);
and U4271 (N_4271,N_4109,N_4175);
nor U4272 (N_4272,N_4198,N_4140);
and U4273 (N_4273,N_4064,N_4196);
or U4274 (N_4274,N_4066,N_4011);
nand U4275 (N_4275,N_4018,N_4149);
nor U4276 (N_4276,N_4065,N_4001);
or U4277 (N_4277,N_4102,N_4098);
nor U4278 (N_4278,N_4057,N_4125);
nor U4279 (N_4279,N_4077,N_4016);
and U4280 (N_4280,N_4189,N_4004);
nand U4281 (N_4281,N_4070,N_4122);
nor U4282 (N_4282,N_4117,N_4005);
nor U4283 (N_4283,N_4019,N_4080);
and U4284 (N_4284,N_4104,N_4150);
and U4285 (N_4285,N_4038,N_4072);
or U4286 (N_4286,N_4008,N_4124);
or U4287 (N_4287,N_4116,N_4087);
nor U4288 (N_4288,N_4136,N_4090);
and U4289 (N_4289,N_4148,N_4167);
nand U4290 (N_4290,N_4024,N_4187);
nor U4291 (N_4291,N_4097,N_4111);
or U4292 (N_4292,N_4193,N_4151);
nor U4293 (N_4293,N_4121,N_4099);
or U4294 (N_4294,N_4069,N_4026);
and U4295 (N_4295,N_4195,N_4031);
nor U4296 (N_4296,N_4120,N_4078);
or U4297 (N_4297,N_4197,N_4020);
and U4298 (N_4298,N_4048,N_4076);
nor U4299 (N_4299,N_4083,N_4174);
or U4300 (N_4300,N_4057,N_4020);
nand U4301 (N_4301,N_4018,N_4029);
or U4302 (N_4302,N_4136,N_4138);
nand U4303 (N_4303,N_4129,N_4053);
nand U4304 (N_4304,N_4019,N_4105);
and U4305 (N_4305,N_4076,N_4138);
and U4306 (N_4306,N_4145,N_4045);
nor U4307 (N_4307,N_4199,N_4056);
nand U4308 (N_4308,N_4016,N_4133);
nand U4309 (N_4309,N_4112,N_4027);
nor U4310 (N_4310,N_4170,N_4101);
or U4311 (N_4311,N_4195,N_4000);
and U4312 (N_4312,N_4071,N_4097);
or U4313 (N_4313,N_4172,N_4116);
and U4314 (N_4314,N_4106,N_4112);
and U4315 (N_4315,N_4094,N_4040);
or U4316 (N_4316,N_4015,N_4007);
and U4317 (N_4317,N_4134,N_4038);
nor U4318 (N_4318,N_4081,N_4118);
or U4319 (N_4319,N_4173,N_4049);
and U4320 (N_4320,N_4189,N_4159);
nand U4321 (N_4321,N_4055,N_4068);
nor U4322 (N_4322,N_4023,N_4019);
nor U4323 (N_4323,N_4162,N_4025);
or U4324 (N_4324,N_4006,N_4198);
and U4325 (N_4325,N_4004,N_4001);
nor U4326 (N_4326,N_4167,N_4114);
nor U4327 (N_4327,N_4139,N_4072);
or U4328 (N_4328,N_4119,N_4195);
or U4329 (N_4329,N_4088,N_4190);
and U4330 (N_4330,N_4127,N_4090);
and U4331 (N_4331,N_4174,N_4186);
nand U4332 (N_4332,N_4017,N_4034);
nand U4333 (N_4333,N_4135,N_4173);
nor U4334 (N_4334,N_4039,N_4038);
and U4335 (N_4335,N_4178,N_4191);
and U4336 (N_4336,N_4199,N_4110);
or U4337 (N_4337,N_4193,N_4074);
nand U4338 (N_4338,N_4124,N_4112);
and U4339 (N_4339,N_4010,N_4098);
or U4340 (N_4340,N_4132,N_4179);
or U4341 (N_4341,N_4174,N_4188);
nand U4342 (N_4342,N_4186,N_4124);
or U4343 (N_4343,N_4154,N_4049);
nor U4344 (N_4344,N_4180,N_4112);
or U4345 (N_4345,N_4180,N_4029);
nand U4346 (N_4346,N_4176,N_4187);
nand U4347 (N_4347,N_4072,N_4050);
and U4348 (N_4348,N_4069,N_4084);
nor U4349 (N_4349,N_4145,N_4187);
nor U4350 (N_4350,N_4078,N_4169);
and U4351 (N_4351,N_4089,N_4006);
or U4352 (N_4352,N_4108,N_4070);
nor U4353 (N_4353,N_4156,N_4138);
nor U4354 (N_4354,N_4035,N_4017);
and U4355 (N_4355,N_4019,N_4004);
and U4356 (N_4356,N_4117,N_4086);
and U4357 (N_4357,N_4045,N_4132);
or U4358 (N_4358,N_4002,N_4180);
nand U4359 (N_4359,N_4045,N_4137);
or U4360 (N_4360,N_4092,N_4016);
and U4361 (N_4361,N_4084,N_4095);
nand U4362 (N_4362,N_4034,N_4057);
nand U4363 (N_4363,N_4178,N_4041);
nor U4364 (N_4364,N_4062,N_4065);
and U4365 (N_4365,N_4132,N_4170);
and U4366 (N_4366,N_4098,N_4002);
nor U4367 (N_4367,N_4143,N_4146);
or U4368 (N_4368,N_4013,N_4189);
nor U4369 (N_4369,N_4128,N_4109);
or U4370 (N_4370,N_4063,N_4137);
nand U4371 (N_4371,N_4102,N_4139);
nand U4372 (N_4372,N_4103,N_4026);
or U4373 (N_4373,N_4153,N_4019);
nand U4374 (N_4374,N_4136,N_4195);
or U4375 (N_4375,N_4148,N_4145);
or U4376 (N_4376,N_4028,N_4123);
nor U4377 (N_4377,N_4127,N_4003);
xnor U4378 (N_4378,N_4160,N_4099);
nand U4379 (N_4379,N_4068,N_4024);
and U4380 (N_4380,N_4028,N_4102);
nor U4381 (N_4381,N_4017,N_4169);
nand U4382 (N_4382,N_4077,N_4145);
nand U4383 (N_4383,N_4187,N_4074);
or U4384 (N_4384,N_4058,N_4052);
nand U4385 (N_4385,N_4108,N_4035);
and U4386 (N_4386,N_4061,N_4001);
or U4387 (N_4387,N_4052,N_4167);
xor U4388 (N_4388,N_4076,N_4069);
nor U4389 (N_4389,N_4136,N_4179);
nand U4390 (N_4390,N_4176,N_4149);
and U4391 (N_4391,N_4005,N_4173);
nor U4392 (N_4392,N_4108,N_4050);
nand U4393 (N_4393,N_4063,N_4009);
nand U4394 (N_4394,N_4039,N_4060);
nor U4395 (N_4395,N_4165,N_4172);
nor U4396 (N_4396,N_4190,N_4035);
nor U4397 (N_4397,N_4136,N_4170);
nor U4398 (N_4398,N_4018,N_4073);
or U4399 (N_4399,N_4021,N_4153);
and U4400 (N_4400,N_4346,N_4321);
nor U4401 (N_4401,N_4310,N_4223);
nor U4402 (N_4402,N_4314,N_4340);
or U4403 (N_4403,N_4390,N_4356);
nand U4404 (N_4404,N_4202,N_4301);
nor U4405 (N_4405,N_4316,N_4203);
or U4406 (N_4406,N_4277,N_4327);
or U4407 (N_4407,N_4315,N_4278);
nor U4408 (N_4408,N_4395,N_4216);
nand U4409 (N_4409,N_4292,N_4399);
or U4410 (N_4410,N_4344,N_4259);
nand U4411 (N_4411,N_4322,N_4373);
and U4412 (N_4412,N_4359,N_4355);
nor U4413 (N_4413,N_4253,N_4298);
nand U4414 (N_4414,N_4367,N_4200);
nand U4415 (N_4415,N_4381,N_4217);
nor U4416 (N_4416,N_4204,N_4362);
or U4417 (N_4417,N_4352,N_4371);
nand U4418 (N_4418,N_4267,N_4319);
nand U4419 (N_4419,N_4323,N_4242);
nor U4420 (N_4420,N_4258,N_4342);
nand U4421 (N_4421,N_4254,N_4376);
or U4422 (N_4422,N_4308,N_4363);
and U4423 (N_4423,N_4256,N_4343);
nand U4424 (N_4424,N_4304,N_4279);
or U4425 (N_4425,N_4320,N_4350);
nand U4426 (N_4426,N_4326,N_4330);
nand U4427 (N_4427,N_4288,N_4234);
and U4428 (N_4428,N_4365,N_4271);
and U4429 (N_4429,N_4303,N_4375);
and U4430 (N_4430,N_4299,N_4382);
and U4431 (N_4431,N_4353,N_4392);
nor U4432 (N_4432,N_4348,N_4374);
or U4433 (N_4433,N_4361,N_4351);
nand U4434 (N_4434,N_4296,N_4295);
and U4435 (N_4435,N_4214,N_4269);
nor U4436 (N_4436,N_4290,N_4249);
nor U4437 (N_4437,N_4397,N_4265);
or U4438 (N_4438,N_4387,N_4246);
and U4439 (N_4439,N_4218,N_4307);
or U4440 (N_4440,N_4283,N_4385);
and U4441 (N_4441,N_4324,N_4360);
nand U4442 (N_4442,N_4391,N_4239);
and U4443 (N_4443,N_4238,N_4335);
nand U4444 (N_4444,N_4305,N_4241);
nor U4445 (N_4445,N_4255,N_4222);
or U4446 (N_4446,N_4328,N_4225);
nand U4447 (N_4447,N_4380,N_4229);
nand U4448 (N_4448,N_4325,N_4369);
nand U4449 (N_4449,N_4302,N_4289);
nand U4450 (N_4450,N_4284,N_4370);
nand U4451 (N_4451,N_4224,N_4354);
nand U4452 (N_4452,N_4245,N_4336);
or U4453 (N_4453,N_4273,N_4262);
or U4454 (N_4454,N_4268,N_4215);
or U4455 (N_4455,N_4383,N_4398);
xnor U4456 (N_4456,N_4338,N_4266);
nand U4457 (N_4457,N_4263,N_4227);
and U4458 (N_4458,N_4368,N_4280);
nor U4459 (N_4459,N_4209,N_4233);
nor U4460 (N_4460,N_4331,N_4388);
and U4461 (N_4461,N_4219,N_4384);
nor U4462 (N_4462,N_4261,N_4358);
and U4463 (N_4463,N_4309,N_4275);
nand U4464 (N_4464,N_4339,N_4201);
and U4465 (N_4465,N_4250,N_4294);
nand U4466 (N_4466,N_4240,N_4377);
nor U4467 (N_4467,N_4291,N_4394);
or U4468 (N_4468,N_4270,N_4226);
nand U4469 (N_4469,N_4286,N_4282);
or U4470 (N_4470,N_4287,N_4332);
or U4471 (N_4471,N_4386,N_4396);
nor U4472 (N_4472,N_4237,N_4379);
nand U4473 (N_4473,N_4341,N_4297);
nand U4474 (N_4474,N_4235,N_4207);
nand U4475 (N_4475,N_4329,N_4393);
nor U4476 (N_4476,N_4347,N_4272);
nand U4477 (N_4477,N_4378,N_4236);
nor U4478 (N_4478,N_4276,N_4274);
or U4479 (N_4479,N_4252,N_4345);
nor U4480 (N_4480,N_4349,N_4206);
or U4481 (N_4481,N_4317,N_4306);
nor U4482 (N_4482,N_4281,N_4260);
nor U4483 (N_4483,N_4285,N_4231);
and U4484 (N_4484,N_4228,N_4372);
or U4485 (N_4485,N_4230,N_4205);
and U4486 (N_4486,N_4334,N_4220);
or U4487 (N_4487,N_4333,N_4337);
nor U4488 (N_4488,N_4364,N_4357);
or U4489 (N_4489,N_4243,N_4210);
nand U4490 (N_4490,N_4212,N_4221);
nand U4491 (N_4491,N_4211,N_4264);
and U4492 (N_4492,N_4312,N_4366);
nand U4493 (N_4493,N_4389,N_4213);
or U4494 (N_4494,N_4248,N_4313);
nand U4495 (N_4495,N_4318,N_4300);
nor U4496 (N_4496,N_4244,N_4232);
or U4497 (N_4497,N_4251,N_4257);
or U4498 (N_4498,N_4293,N_4311);
or U4499 (N_4499,N_4247,N_4208);
and U4500 (N_4500,N_4372,N_4276);
nor U4501 (N_4501,N_4318,N_4391);
and U4502 (N_4502,N_4241,N_4261);
nand U4503 (N_4503,N_4246,N_4353);
nor U4504 (N_4504,N_4269,N_4396);
nor U4505 (N_4505,N_4349,N_4379);
nor U4506 (N_4506,N_4233,N_4264);
nor U4507 (N_4507,N_4371,N_4265);
or U4508 (N_4508,N_4287,N_4220);
nor U4509 (N_4509,N_4248,N_4276);
and U4510 (N_4510,N_4364,N_4320);
nor U4511 (N_4511,N_4375,N_4249);
nand U4512 (N_4512,N_4299,N_4364);
nor U4513 (N_4513,N_4338,N_4274);
or U4514 (N_4514,N_4377,N_4385);
and U4515 (N_4515,N_4371,N_4330);
nand U4516 (N_4516,N_4310,N_4339);
and U4517 (N_4517,N_4347,N_4323);
and U4518 (N_4518,N_4294,N_4331);
nand U4519 (N_4519,N_4222,N_4395);
nor U4520 (N_4520,N_4383,N_4399);
nand U4521 (N_4521,N_4246,N_4293);
nor U4522 (N_4522,N_4281,N_4353);
or U4523 (N_4523,N_4381,N_4318);
xnor U4524 (N_4524,N_4286,N_4219);
nand U4525 (N_4525,N_4216,N_4343);
or U4526 (N_4526,N_4308,N_4369);
and U4527 (N_4527,N_4307,N_4346);
or U4528 (N_4528,N_4398,N_4285);
or U4529 (N_4529,N_4346,N_4387);
or U4530 (N_4530,N_4288,N_4215);
nor U4531 (N_4531,N_4312,N_4214);
or U4532 (N_4532,N_4343,N_4326);
nand U4533 (N_4533,N_4227,N_4379);
and U4534 (N_4534,N_4299,N_4318);
or U4535 (N_4535,N_4259,N_4218);
nand U4536 (N_4536,N_4351,N_4202);
nor U4537 (N_4537,N_4260,N_4368);
or U4538 (N_4538,N_4343,N_4238);
and U4539 (N_4539,N_4298,N_4384);
and U4540 (N_4540,N_4233,N_4305);
and U4541 (N_4541,N_4341,N_4369);
and U4542 (N_4542,N_4231,N_4331);
nand U4543 (N_4543,N_4377,N_4288);
nor U4544 (N_4544,N_4282,N_4294);
nand U4545 (N_4545,N_4239,N_4289);
or U4546 (N_4546,N_4298,N_4265);
and U4547 (N_4547,N_4302,N_4205);
xnor U4548 (N_4548,N_4353,N_4371);
or U4549 (N_4549,N_4317,N_4269);
nand U4550 (N_4550,N_4307,N_4296);
and U4551 (N_4551,N_4202,N_4366);
or U4552 (N_4552,N_4273,N_4257);
nor U4553 (N_4553,N_4247,N_4243);
or U4554 (N_4554,N_4322,N_4292);
and U4555 (N_4555,N_4237,N_4365);
nor U4556 (N_4556,N_4293,N_4269);
nor U4557 (N_4557,N_4393,N_4398);
and U4558 (N_4558,N_4383,N_4209);
nand U4559 (N_4559,N_4361,N_4226);
nor U4560 (N_4560,N_4399,N_4284);
xnor U4561 (N_4561,N_4354,N_4226);
nand U4562 (N_4562,N_4256,N_4254);
nor U4563 (N_4563,N_4347,N_4341);
or U4564 (N_4564,N_4259,N_4337);
or U4565 (N_4565,N_4352,N_4254);
nor U4566 (N_4566,N_4223,N_4255);
nand U4567 (N_4567,N_4340,N_4367);
nand U4568 (N_4568,N_4360,N_4338);
and U4569 (N_4569,N_4228,N_4289);
or U4570 (N_4570,N_4267,N_4320);
xnor U4571 (N_4571,N_4340,N_4257);
nor U4572 (N_4572,N_4218,N_4369);
or U4573 (N_4573,N_4327,N_4376);
nand U4574 (N_4574,N_4204,N_4299);
nor U4575 (N_4575,N_4280,N_4208);
nand U4576 (N_4576,N_4237,N_4249);
nor U4577 (N_4577,N_4358,N_4392);
and U4578 (N_4578,N_4311,N_4330);
nand U4579 (N_4579,N_4285,N_4330);
or U4580 (N_4580,N_4223,N_4391);
or U4581 (N_4581,N_4256,N_4266);
nand U4582 (N_4582,N_4223,N_4201);
nor U4583 (N_4583,N_4230,N_4340);
nand U4584 (N_4584,N_4383,N_4370);
and U4585 (N_4585,N_4273,N_4377);
nand U4586 (N_4586,N_4246,N_4334);
nor U4587 (N_4587,N_4302,N_4268);
nor U4588 (N_4588,N_4324,N_4363);
and U4589 (N_4589,N_4349,N_4233);
or U4590 (N_4590,N_4304,N_4302);
and U4591 (N_4591,N_4303,N_4313);
nand U4592 (N_4592,N_4235,N_4326);
nand U4593 (N_4593,N_4335,N_4315);
nand U4594 (N_4594,N_4294,N_4244);
and U4595 (N_4595,N_4313,N_4227);
nand U4596 (N_4596,N_4320,N_4376);
and U4597 (N_4597,N_4309,N_4218);
nand U4598 (N_4598,N_4287,N_4216);
or U4599 (N_4599,N_4227,N_4315);
nand U4600 (N_4600,N_4520,N_4478);
nor U4601 (N_4601,N_4521,N_4519);
nor U4602 (N_4602,N_4425,N_4448);
and U4603 (N_4603,N_4569,N_4412);
and U4604 (N_4604,N_4536,N_4576);
nor U4605 (N_4605,N_4582,N_4565);
or U4606 (N_4606,N_4441,N_4431);
and U4607 (N_4607,N_4575,N_4434);
nand U4608 (N_4608,N_4413,N_4444);
nand U4609 (N_4609,N_4513,N_4421);
and U4610 (N_4610,N_4417,N_4447);
nand U4611 (N_4611,N_4564,N_4499);
or U4612 (N_4612,N_4526,N_4462);
nor U4613 (N_4613,N_4436,N_4454);
and U4614 (N_4614,N_4491,N_4430);
nor U4615 (N_4615,N_4405,N_4533);
nand U4616 (N_4616,N_4556,N_4545);
or U4617 (N_4617,N_4594,N_4498);
nand U4618 (N_4618,N_4581,N_4407);
nand U4619 (N_4619,N_4470,N_4461);
nand U4620 (N_4620,N_4518,N_4563);
or U4621 (N_4621,N_4449,N_4488);
nand U4622 (N_4622,N_4437,N_4466);
nand U4623 (N_4623,N_4524,N_4535);
or U4624 (N_4624,N_4540,N_4450);
nand U4625 (N_4625,N_4503,N_4458);
nand U4626 (N_4626,N_4426,N_4493);
nor U4627 (N_4627,N_4473,N_4501);
nand U4628 (N_4628,N_4428,N_4577);
nand U4629 (N_4629,N_4588,N_4476);
xnor U4630 (N_4630,N_4538,N_4487);
nand U4631 (N_4631,N_4459,N_4525);
nor U4632 (N_4632,N_4490,N_4500);
or U4633 (N_4633,N_4504,N_4512);
or U4634 (N_4634,N_4591,N_4422);
or U4635 (N_4635,N_4557,N_4481);
nor U4636 (N_4636,N_4570,N_4541);
nor U4637 (N_4637,N_4592,N_4406);
and U4638 (N_4638,N_4559,N_4584);
and U4639 (N_4639,N_4420,N_4401);
or U4640 (N_4640,N_4483,N_4497);
and U4641 (N_4641,N_4587,N_4502);
or U4642 (N_4642,N_4469,N_4403);
nand U4643 (N_4643,N_4456,N_4457);
nand U4644 (N_4644,N_4530,N_4414);
nand U4645 (N_4645,N_4567,N_4475);
nand U4646 (N_4646,N_4534,N_4463);
nor U4647 (N_4647,N_4558,N_4451);
nand U4648 (N_4648,N_4548,N_4589);
or U4649 (N_4649,N_4593,N_4400);
or U4650 (N_4650,N_4508,N_4532);
nor U4651 (N_4651,N_4544,N_4560);
nor U4652 (N_4652,N_4566,N_4554);
nor U4653 (N_4653,N_4585,N_4439);
nand U4654 (N_4654,N_4598,N_4552);
or U4655 (N_4655,N_4510,N_4409);
or U4656 (N_4656,N_4489,N_4468);
and U4657 (N_4657,N_4402,N_4527);
nand U4658 (N_4658,N_4419,N_4474);
nor U4659 (N_4659,N_4543,N_4590);
or U4660 (N_4660,N_4486,N_4446);
nor U4661 (N_4661,N_4432,N_4416);
or U4662 (N_4662,N_4578,N_4484);
nand U4663 (N_4663,N_4410,N_4443);
or U4664 (N_4664,N_4507,N_4442);
nor U4665 (N_4665,N_4597,N_4472);
or U4666 (N_4666,N_4572,N_4531);
and U4667 (N_4667,N_4579,N_4408);
nor U4668 (N_4668,N_4523,N_4528);
nor U4669 (N_4669,N_4539,N_4452);
and U4670 (N_4670,N_4511,N_4551);
nand U4671 (N_4671,N_4516,N_4573);
or U4672 (N_4672,N_4514,N_4440);
or U4673 (N_4673,N_4477,N_4479);
nor U4674 (N_4674,N_4429,N_4537);
nor U4675 (N_4675,N_4415,N_4404);
or U4676 (N_4676,N_4492,N_4424);
and U4677 (N_4677,N_4427,N_4561);
nand U4678 (N_4678,N_4480,N_4571);
or U4679 (N_4679,N_4550,N_4494);
or U4680 (N_4680,N_4485,N_4465);
or U4681 (N_4681,N_4586,N_4574);
nor U4682 (N_4682,N_4453,N_4505);
nand U4683 (N_4683,N_4595,N_4555);
or U4684 (N_4684,N_4568,N_4517);
nand U4685 (N_4685,N_4509,N_4562);
or U4686 (N_4686,N_4471,N_4542);
nor U4687 (N_4687,N_4460,N_4553);
or U4688 (N_4688,N_4495,N_4418);
nor U4689 (N_4689,N_4599,N_4515);
and U4690 (N_4690,N_4455,N_4433);
and U4691 (N_4691,N_4506,N_4549);
or U4692 (N_4692,N_4445,N_4435);
or U4693 (N_4693,N_4423,N_4546);
nor U4694 (N_4694,N_4496,N_4438);
nand U4695 (N_4695,N_4580,N_4464);
and U4696 (N_4696,N_4411,N_4482);
and U4697 (N_4697,N_4467,N_4547);
or U4698 (N_4698,N_4583,N_4522);
and U4699 (N_4699,N_4596,N_4529);
nor U4700 (N_4700,N_4493,N_4402);
nand U4701 (N_4701,N_4410,N_4490);
nor U4702 (N_4702,N_4568,N_4412);
xnor U4703 (N_4703,N_4557,N_4543);
nor U4704 (N_4704,N_4459,N_4431);
and U4705 (N_4705,N_4484,N_4405);
or U4706 (N_4706,N_4532,N_4492);
and U4707 (N_4707,N_4489,N_4561);
nand U4708 (N_4708,N_4517,N_4497);
nand U4709 (N_4709,N_4540,N_4578);
and U4710 (N_4710,N_4547,N_4506);
and U4711 (N_4711,N_4526,N_4592);
nor U4712 (N_4712,N_4565,N_4517);
and U4713 (N_4713,N_4483,N_4412);
nand U4714 (N_4714,N_4556,N_4567);
nor U4715 (N_4715,N_4483,N_4476);
or U4716 (N_4716,N_4469,N_4451);
or U4717 (N_4717,N_4592,N_4453);
and U4718 (N_4718,N_4498,N_4591);
or U4719 (N_4719,N_4569,N_4521);
or U4720 (N_4720,N_4558,N_4559);
nand U4721 (N_4721,N_4462,N_4426);
nor U4722 (N_4722,N_4582,N_4451);
or U4723 (N_4723,N_4579,N_4550);
or U4724 (N_4724,N_4512,N_4419);
and U4725 (N_4725,N_4519,N_4553);
or U4726 (N_4726,N_4468,N_4578);
and U4727 (N_4727,N_4545,N_4559);
nor U4728 (N_4728,N_4475,N_4534);
and U4729 (N_4729,N_4593,N_4418);
nor U4730 (N_4730,N_4421,N_4584);
nor U4731 (N_4731,N_4588,N_4590);
or U4732 (N_4732,N_4466,N_4584);
or U4733 (N_4733,N_4533,N_4474);
or U4734 (N_4734,N_4564,N_4558);
nor U4735 (N_4735,N_4523,N_4485);
nor U4736 (N_4736,N_4491,N_4550);
nor U4737 (N_4737,N_4474,N_4546);
nand U4738 (N_4738,N_4471,N_4509);
nand U4739 (N_4739,N_4580,N_4597);
nand U4740 (N_4740,N_4442,N_4574);
or U4741 (N_4741,N_4452,N_4533);
or U4742 (N_4742,N_4520,N_4595);
nor U4743 (N_4743,N_4521,N_4579);
or U4744 (N_4744,N_4549,N_4482);
or U4745 (N_4745,N_4493,N_4512);
or U4746 (N_4746,N_4431,N_4416);
or U4747 (N_4747,N_4409,N_4528);
and U4748 (N_4748,N_4556,N_4528);
and U4749 (N_4749,N_4520,N_4517);
nor U4750 (N_4750,N_4490,N_4458);
xor U4751 (N_4751,N_4535,N_4495);
nor U4752 (N_4752,N_4570,N_4418);
nand U4753 (N_4753,N_4408,N_4404);
or U4754 (N_4754,N_4416,N_4426);
nor U4755 (N_4755,N_4543,N_4466);
or U4756 (N_4756,N_4505,N_4503);
nor U4757 (N_4757,N_4450,N_4464);
and U4758 (N_4758,N_4548,N_4413);
and U4759 (N_4759,N_4436,N_4559);
or U4760 (N_4760,N_4443,N_4424);
nand U4761 (N_4761,N_4403,N_4461);
or U4762 (N_4762,N_4401,N_4572);
nor U4763 (N_4763,N_4433,N_4590);
and U4764 (N_4764,N_4597,N_4508);
nand U4765 (N_4765,N_4430,N_4539);
nand U4766 (N_4766,N_4531,N_4510);
or U4767 (N_4767,N_4585,N_4547);
or U4768 (N_4768,N_4542,N_4484);
and U4769 (N_4769,N_4559,N_4431);
nor U4770 (N_4770,N_4520,N_4436);
and U4771 (N_4771,N_4544,N_4486);
nor U4772 (N_4772,N_4449,N_4587);
nor U4773 (N_4773,N_4579,N_4502);
and U4774 (N_4774,N_4427,N_4586);
and U4775 (N_4775,N_4444,N_4576);
nor U4776 (N_4776,N_4555,N_4579);
nor U4777 (N_4777,N_4476,N_4403);
nor U4778 (N_4778,N_4449,N_4450);
nor U4779 (N_4779,N_4494,N_4594);
nand U4780 (N_4780,N_4422,N_4496);
or U4781 (N_4781,N_4484,N_4435);
or U4782 (N_4782,N_4578,N_4466);
nor U4783 (N_4783,N_4572,N_4569);
or U4784 (N_4784,N_4518,N_4478);
or U4785 (N_4785,N_4431,N_4512);
and U4786 (N_4786,N_4475,N_4580);
and U4787 (N_4787,N_4478,N_4563);
or U4788 (N_4788,N_4570,N_4442);
nor U4789 (N_4789,N_4467,N_4465);
nand U4790 (N_4790,N_4578,N_4559);
nor U4791 (N_4791,N_4480,N_4555);
or U4792 (N_4792,N_4473,N_4448);
or U4793 (N_4793,N_4550,N_4594);
nand U4794 (N_4794,N_4540,N_4483);
or U4795 (N_4795,N_4560,N_4461);
nor U4796 (N_4796,N_4444,N_4532);
and U4797 (N_4797,N_4408,N_4528);
and U4798 (N_4798,N_4473,N_4552);
nand U4799 (N_4799,N_4491,N_4498);
nand U4800 (N_4800,N_4642,N_4630);
and U4801 (N_4801,N_4649,N_4720);
nand U4802 (N_4802,N_4656,N_4635);
and U4803 (N_4803,N_4640,N_4637);
nor U4804 (N_4804,N_4758,N_4616);
nor U4805 (N_4805,N_4783,N_4683);
nand U4806 (N_4806,N_4704,N_4661);
and U4807 (N_4807,N_4620,N_4615);
nand U4808 (N_4808,N_4751,N_4770);
nand U4809 (N_4809,N_4673,N_4768);
nand U4810 (N_4810,N_4767,N_4716);
and U4811 (N_4811,N_4714,N_4709);
nand U4812 (N_4812,N_4687,N_4762);
or U4813 (N_4813,N_4644,N_4662);
nand U4814 (N_4814,N_4652,N_4638);
or U4815 (N_4815,N_4625,N_4645);
or U4816 (N_4816,N_4746,N_4753);
nand U4817 (N_4817,N_4633,N_4749);
nand U4818 (N_4818,N_4786,N_4735);
nand U4819 (N_4819,N_4611,N_4691);
nand U4820 (N_4820,N_4732,N_4699);
nand U4821 (N_4821,N_4692,N_4772);
and U4822 (N_4822,N_4680,N_4710);
or U4823 (N_4823,N_4679,N_4648);
and U4824 (N_4824,N_4670,N_4621);
or U4825 (N_4825,N_4723,N_4764);
nand U4826 (N_4826,N_4756,N_4612);
nand U4827 (N_4827,N_4696,N_4654);
and U4828 (N_4828,N_4726,N_4602);
or U4829 (N_4829,N_4658,N_4702);
nand U4830 (N_4830,N_4603,N_4632);
nor U4831 (N_4831,N_4655,N_4799);
nand U4832 (N_4832,N_4643,N_4610);
xnor U4833 (N_4833,N_4766,N_4759);
or U4834 (N_4834,N_4761,N_4733);
or U4835 (N_4835,N_4698,N_4697);
nor U4836 (N_4836,N_4790,N_4779);
and U4837 (N_4837,N_4719,N_4795);
and U4838 (N_4838,N_4787,N_4774);
nor U4839 (N_4839,N_4685,N_4659);
and U4840 (N_4840,N_4639,N_4744);
and U4841 (N_4841,N_4600,N_4700);
nand U4842 (N_4842,N_4788,N_4628);
or U4843 (N_4843,N_4796,N_4717);
nand U4844 (N_4844,N_4688,N_4686);
and U4845 (N_4845,N_4609,N_4728);
nor U4846 (N_4846,N_4678,N_4782);
and U4847 (N_4847,N_4624,N_4693);
and U4848 (N_4848,N_4608,N_4619);
nor U4849 (N_4849,N_4684,N_4739);
nand U4850 (N_4850,N_4731,N_4669);
and U4851 (N_4851,N_4727,N_4706);
nor U4852 (N_4852,N_4765,N_4657);
and U4853 (N_4853,N_4613,N_4694);
nor U4854 (N_4854,N_4614,N_4789);
xnor U4855 (N_4855,N_4622,N_4734);
and U4856 (N_4856,N_4682,N_4660);
nor U4857 (N_4857,N_4650,N_4791);
nor U4858 (N_4858,N_4607,N_4776);
and U4859 (N_4859,N_4745,N_4631);
nand U4860 (N_4860,N_4646,N_4778);
nand U4861 (N_4861,N_4663,N_4736);
nand U4862 (N_4862,N_4703,N_4653);
nor U4863 (N_4863,N_4771,N_4741);
nand U4864 (N_4864,N_4623,N_4668);
nor U4865 (N_4865,N_4618,N_4626);
and U4866 (N_4866,N_4636,N_4627);
nor U4867 (N_4867,N_4634,N_4674);
and U4868 (N_4868,N_4737,N_4705);
or U4869 (N_4869,N_4711,N_4675);
or U4870 (N_4870,N_4690,N_4740);
nor U4871 (N_4871,N_4665,N_4672);
nand U4872 (N_4872,N_4677,N_4689);
or U4873 (N_4873,N_4721,N_4777);
and U4874 (N_4874,N_4666,N_4747);
nand U4875 (N_4875,N_4738,N_4664);
and U4876 (N_4876,N_4629,N_4617);
or U4877 (N_4877,N_4792,N_4671);
and U4878 (N_4878,N_4724,N_4647);
nand U4879 (N_4879,N_4712,N_4773);
and U4880 (N_4880,N_4651,N_4794);
nand U4881 (N_4881,N_4763,N_4730);
or U4882 (N_4882,N_4785,N_4729);
nor U4883 (N_4883,N_4604,N_4641);
or U4884 (N_4884,N_4775,N_4754);
and U4885 (N_4885,N_4797,N_4718);
and U4886 (N_4886,N_4798,N_4667);
nor U4887 (N_4887,N_4707,N_4713);
and U4888 (N_4888,N_4752,N_4750);
nor U4889 (N_4889,N_4725,N_4701);
nand U4890 (N_4890,N_4601,N_4757);
nor U4891 (N_4891,N_4695,N_4743);
and U4892 (N_4892,N_4681,N_4676);
nor U4893 (N_4893,N_4760,N_4748);
nor U4894 (N_4894,N_4793,N_4769);
nand U4895 (N_4895,N_4780,N_4742);
or U4896 (N_4896,N_4722,N_4708);
nor U4897 (N_4897,N_4755,N_4784);
or U4898 (N_4898,N_4606,N_4781);
nand U4899 (N_4899,N_4715,N_4605);
and U4900 (N_4900,N_4659,N_4751);
nor U4901 (N_4901,N_4782,N_4728);
nor U4902 (N_4902,N_4646,N_4658);
and U4903 (N_4903,N_4667,N_4604);
nand U4904 (N_4904,N_4648,N_4735);
xnor U4905 (N_4905,N_4786,N_4660);
nor U4906 (N_4906,N_4700,N_4636);
nand U4907 (N_4907,N_4640,N_4744);
and U4908 (N_4908,N_4685,N_4660);
or U4909 (N_4909,N_4608,N_4771);
nor U4910 (N_4910,N_4793,N_4772);
nand U4911 (N_4911,N_4743,N_4757);
or U4912 (N_4912,N_4612,N_4723);
nor U4913 (N_4913,N_4667,N_4676);
nand U4914 (N_4914,N_4689,N_4717);
or U4915 (N_4915,N_4773,N_4633);
and U4916 (N_4916,N_4640,N_4740);
xnor U4917 (N_4917,N_4644,N_4693);
nand U4918 (N_4918,N_4602,N_4784);
nand U4919 (N_4919,N_4727,N_4677);
nor U4920 (N_4920,N_4608,N_4775);
or U4921 (N_4921,N_4729,N_4797);
and U4922 (N_4922,N_4773,N_4769);
and U4923 (N_4923,N_4748,N_4744);
or U4924 (N_4924,N_4703,N_4721);
or U4925 (N_4925,N_4716,N_4694);
or U4926 (N_4926,N_4652,N_4763);
nor U4927 (N_4927,N_4778,N_4785);
nor U4928 (N_4928,N_4779,N_4675);
nor U4929 (N_4929,N_4691,N_4634);
nand U4930 (N_4930,N_4798,N_4684);
or U4931 (N_4931,N_4797,N_4615);
or U4932 (N_4932,N_4791,N_4663);
nand U4933 (N_4933,N_4610,N_4684);
and U4934 (N_4934,N_4693,N_4628);
nor U4935 (N_4935,N_4791,N_4639);
nor U4936 (N_4936,N_4791,N_4653);
and U4937 (N_4937,N_4763,N_4690);
nor U4938 (N_4938,N_4648,N_4777);
and U4939 (N_4939,N_4720,N_4643);
or U4940 (N_4940,N_4650,N_4689);
and U4941 (N_4941,N_4608,N_4652);
nor U4942 (N_4942,N_4767,N_4607);
and U4943 (N_4943,N_4745,N_4691);
or U4944 (N_4944,N_4794,N_4690);
and U4945 (N_4945,N_4643,N_4657);
nand U4946 (N_4946,N_4601,N_4652);
nand U4947 (N_4947,N_4694,N_4675);
nor U4948 (N_4948,N_4630,N_4636);
nand U4949 (N_4949,N_4774,N_4698);
nand U4950 (N_4950,N_4749,N_4663);
nand U4951 (N_4951,N_4790,N_4643);
and U4952 (N_4952,N_4782,N_4784);
nand U4953 (N_4953,N_4723,N_4749);
or U4954 (N_4954,N_4742,N_4638);
and U4955 (N_4955,N_4726,N_4798);
nand U4956 (N_4956,N_4738,N_4725);
and U4957 (N_4957,N_4666,N_4797);
or U4958 (N_4958,N_4625,N_4671);
or U4959 (N_4959,N_4732,N_4768);
nand U4960 (N_4960,N_4681,N_4734);
nand U4961 (N_4961,N_4740,N_4636);
and U4962 (N_4962,N_4683,N_4630);
and U4963 (N_4963,N_4771,N_4750);
or U4964 (N_4964,N_4636,N_4691);
or U4965 (N_4965,N_4773,N_4755);
and U4966 (N_4966,N_4607,N_4649);
or U4967 (N_4967,N_4799,N_4782);
or U4968 (N_4968,N_4721,N_4602);
and U4969 (N_4969,N_4741,N_4791);
nor U4970 (N_4970,N_4759,N_4773);
nor U4971 (N_4971,N_4641,N_4691);
and U4972 (N_4972,N_4601,N_4733);
and U4973 (N_4973,N_4603,N_4728);
nor U4974 (N_4974,N_4736,N_4783);
nand U4975 (N_4975,N_4782,N_4720);
or U4976 (N_4976,N_4752,N_4786);
nand U4977 (N_4977,N_4695,N_4704);
nor U4978 (N_4978,N_4692,N_4605);
nor U4979 (N_4979,N_4777,N_4656);
or U4980 (N_4980,N_4712,N_4678);
or U4981 (N_4981,N_4713,N_4769);
nor U4982 (N_4982,N_4663,N_4643);
nand U4983 (N_4983,N_4723,N_4639);
nand U4984 (N_4984,N_4631,N_4608);
nand U4985 (N_4985,N_4706,N_4647);
nand U4986 (N_4986,N_4796,N_4649);
or U4987 (N_4987,N_4780,N_4619);
and U4988 (N_4988,N_4748,N_4609);
and U4989 (N_4989,N_4703,N_4631);
and U4990 (N_4990,N_4664,N_4720);
or U4991 (N_4991,N_4748,N_4796);
and U4992 (N_4992,N_4696,N_4721);
nand U4993 (N_4993,N_4787,N_4649);
and U4994 (N_4994,N_4727,N_4616);
or U4995 (N_4995,N_4614,N_4689);
or U4996 (N_4996,N_4697,N_4787);
nor U4997 (N_4997,N_4622,N_4607);
nand U4998 (N_4998,N_4644,N_4615);
or U4999 (N_4999,N_4676,N_4741);
nand U5000 (N_5000,N_4931,N_4999);
and U5001 (N_5001,N_4920,N_4893);
and U5002 (N_5002,N_4800,N_4868);
nand U5003 (N_5003,N_4903,N_4938);
nor U5004 (N_5004,N_4873,N_4930);
and U5005 (N_5005,N_4841,N_4862);
nand U5006 (N_5006,N_4969,N_4855);
nor U5007 (N_5007,N_4933,N_4832);
nand U5008 (N_5008,N_4911,N_4808);
nand U5009 (N_5009,N_4945,N_4954);
or U5010 (N_5010,N_4995,N_4972);
or U5011 (N_5011,N_4924,N_4913);
or U5012 (N_5012,N_4927,N_4974);
nor U5013 (N_5013,N_4856,N_4882);
nand U5014 (N_5014,N_4964,N_4850);
or U5015 (N_5015,N_4942,N_4990);
or U5016 (N_5016,N_4848,N_4846);
or U5017 (N_5017,N_4949,N_4963);
nand U5018 (N_5018,N_4810,N_4912);
nand U5019 (N_5019,N_4943,N_4894);
and U5020 (N_5020,N_4910,N_4830);
xnor U5021 (N_5021,N_4859,N_4857);
nand U5022 (N_5022,N_4971,N_4858);
nor U5023 (N_5023,N_4998,N_4831);
and U5024 (N_5024,N_4878,N_4803);
nand U5025 (N_5025,N_4922,N_4989);
and U5026 (N_5026,N_4881,N_4839);
or U5027 (N_5027,N_4946,N_4853);
nand U5028 (N_5028,N_4840,N_4937);
nor U5029 (N_5029,N_4960,N_4934);
or U5030 (N_5030,N_4861,N_4854);
nor U5031 (N_5031,N_4864,N_4898);
or U5032 (N_5032,N_4996,N_4897);
nor U5033 (N_5033,N_4895,N_4885);
or U5034 (N_5034,N_4968,N_4829);
nand U5035 (N_5035,N_4994,N_4825);
and U5036 (N_5036,N_4886,N_4980);
or U5037 (N_5037,N_4965,N_4958);
and U5038 (N_5038,N_4879,N_4953);
and U5039 (N_5039,N_4932,N_4973);
and U5040 (N_5040,N_4872,N_4802);
or U5041 (N_5041,N_4834,N_4904);
or U5042 (N_5042,N_4816,N_4884);
and U5043 (N_5043,N_4935,N_4818);
nor U5044 (N_5044,N_4941,N_4806);
nor U5045 (N_5045,N_4906,N_4915);
nor U5046 (N_5046,N_4837,N_4993);
or U5047 (N_5047,N_4842,N_4908);
and U5048 (N_5048,N_4871,N_4813);
xnor U5049 (N_5049,N_4838,N_4950);
or U5050 (N_5050,N_4822,N_4992);
or U5051 (N_5051,N_4807,N_4940);
nor U5052 (N_5052,N_4966,N_4833);
and U5053 (N_5053,N_4919,N_4959);
nand U5054 (N_5054,N_4918,N_4890);
nand U5055 (N_5055,N_4978,N_4819);
and U5056 (N_5056,N_4815,N_4985);
nor U5057 (N_5057,N_4902,N_4983);
or U5058 (N_5058,N_4962,N_4847);
nor U5059 (N_5059,N_4923,N_4899);
nor U5060 (N_5060,N_4811,N_4874);
nor U5061 (N_5061,N_4970,N_4827);
nand U5062 (N_5062,N_4892,N_4976);
and U5063 (N_5063,N_4948,N_4952);
nand U5064 (N_5064,N_4977,N_4896);
nor U5065 (N_5065,N_4988,N_4925);
nor U5066 (N_5066,N_4826,N_4801);
or U5067 (N_5067,N_4835,N_4814);
and U5068 (N_5068,N_4891,N_4986);
and U5069 (N_5069,N_4867,N_4984);
and U5070 (N_5070,N_4851,N_4957);
or U5071 (N_5071,N_4870,N_4843);
or U5072 (N_5072,N_4875,N_4956);
and U5073 (N_5073,N_4929,N_4887);
and U5074 (N_5074,N_4967,N_4975);
nand U5075 (N_5075,N_4888,N_4914);
nor U5076 (N_5076,N_4804,N_4844);
nor U5077 (N_5077,N_4828,N_4823);
nand U5078 (N_5078,N_4909,N_4820);
nand U5079 (N_5079,N_4997,N_4947);
nand U5080 (N_5080,N_4936,N_4812);
nor U5081 (N_5081,N_4824,N_4880);
nand U5082 (N_5082,N_4901,N_4979);
and U5083 (N_5083,N_4866,N_4921);
or U5084 (N_5084,N_4852,N_4951);
nor U5085 (N_5085,N_4907,N_4928);
and U5086 (N_5086,N_4860,N_4805);
nor U5087 (N_5087,N_4981,N_4917);
or U5088 (N_5088,N_4987,N_4849);
nand U5089 (N_5089,N_4900,N_4876);
or U5090 (N_5090,N_4821,N_4991);
nand U5091 (N_5091,N_4877,N_4863);
nand U5092 (N_5092,N_4961,N_4869);
xor U5093 (N_5093,N_4955,N_4817);
or U5094 (N_5094,N_4916,N_4939);
nand U5095 (N_5095,N_4836,N_4865);
and U5096 (N_5096,N_4905,N_4926);
or U5097 (N_5097,N_4845,N_4889);
and U5098 (N_5098,N_4982,N_4883);
or U5099 (N_5099,N_4809,N_4944);
and U5100 (N_5100,N_4967,N_4981);
or U5101 (N_5101,N_4947,N_4814);
or U5102 (N_5102,N_4980,N_4882);
and U5103 (N_5103,N_4888,N_4867);
nand U5104 (N_5104,N_4915,N_4944);
or U5105 (N_5105,N_4883,N_4804);
or U5106 (N_5106,N_4900,N_4980);
nand U5107 (N_5107,N_4901,N_4991);
nor U5108 (N_5108,N_4830,N_4862);
or U5109 (N_5109,N_4853,N_4966);
nand U5110 (N_5110,N_4865,N_4942);
nand U5111 (N_5111,N_4828,N_4950);
nand U5112 (N_5112,N_4954,N_4813);
nand U5113 (N_5113,N_4941,N_4858);
and U5114 (N_5114,N_4844,N_4821);
nor U5115 (N_5115,N_4862,N_4822);
or U5116 (N_5116,N_4871,N_4836);
nand U5117 (N_5117,N_4899,N_4802);
nor U5118 (N_5118,N_4912,N_4993);
or U5119 (N_5119,N_4852,N_4814);
nor U5120 (N_5120,N_4802,N_4928);
and U5121 (N_5121,N_4932,N_4976);
nand U5122 (N_5122,N_4828,N_4974);
nor U5123 (N_5123,N_4922,N_4833);
xor U5124 (N_5124,N_4960,N_4932);
nor U5125 (N_5125,N_4814,N_4925);
nor U5126 (N_5126,N_4844,N_4932);
nand U5127 (N_5127,N_4952,N_4930);
or U5128 (N_5128,N_4801,N_4845);
nor U5129 (N_5129,N_4940,N_4860);
nor U5130 (N_5130,N_4812,N_4931);
nand U5131 (N_5131,N_4894,N_4875);
nor U5132 (N_5132,N_4937,N_4897);
nor U5133 (N_5133,N_4911,N_4881);
nor U5134 (N_5134,N_4959,N_4848);
nor U5135 (N_5135,N_4861,N_4946);
nand U5136 (N_5136,N_4837,N_4976);
or U5137 (N_5137,N_4987,N_4819);
nor U5138 (N_5138,N_4950,N_4881);
nand U5139 (N_5139,N_4954,N_4888);
or U5140 (N_5140,N_4948,N_4807);
nor U5141 (N_5141,N_4960,N_4887);
nor U5142 (N_5142,N_4932,N_4876);
nor U5143 (N_5143,N_4960,N_4833);
or U5144 (N_5144,N_4942,N_4867);
and U5145 (N_5145,N_4935,N_4978);
nor U5146 (N_5146,N_4871,N_4905);
or U5147 (N_5147,N_4820,N_4800);
nor U5148 (N_5148,N_4941,N_4969);
nor U5149 (N_5149,N_4811,N_4960);
and U5150 (N_5150,N_4855,N_4955);
nand U5151 (N_5151,N_4995,N_4960);
nand U5152 (N_5152,N_4969,N_4983);
or U5153 (N_5153,N_4953,N_4974);
or U5154 (N_5154,N_4870,N_4893);
nor U5155 (N_5155,N_4997,N_4941);
and U5156 (N_5156,N_4958,N_4886);
nand U5157 (N_5157,N_4959,N_4943);
nand U5158 (N_5158,N_4838,N_4913);
nor U5159 (N_5159,N_4998,N_4872);
nor U5160 (N_5160,N_4837,N_4805);
nand U5161 (N_5161,N_4812,N_4838);
nor U5162 (N_5162,N_4831,N_4855);
or U5163 (N_5163,N_4823,N_4969);
or U5164 (N_5164,N_4834,N_4967);
nor U5165 (N_5165,N_4938,N_4986);
and U5166 (N_5166,N_4893,N_4867);
or U5167 (N_5167,N_4906,N_4965);
or U5168 (N_5168,N_4865,N_4830);
and U5169 (N_5169,N_4899,N_4931);
and U5170 (N_5170,N_4818,N_4898);
or U5171 (N_5171,N_4983,N_4936);
nor U5172 (N_5172,N_4993,N_4925);
nor U5173 (N_5173,N_4981,N_4919);
and U5174 (N_5174,N_4936,N_4819);
nor U5175 (N_5175,N_4972,N_4922);
nor U5176 (N_5176,N_4906,N_4895);
nor U5177 (N_5177,N_4990,N_4888);
nor U5178 (N_5178,N_4963,N_4883);
nor U5179 (N_5179,N_4884,N_4912);
nor U5180 (N_5180,N_4953,N_4823);
and U5181 (N_5181,N_4962,N_4816);
or U5182 (N_5182,N_4924,N_4975);
and U5183 (N_5183,N_4973,N_4831);
xnor U5184 (N_5184,N_4832,N_4942);
and U5185 (N_5185,N_4842,N_4914);
nor U5186 (N_5186,N_4825,N_4870);
nor U5187 (N_5187,N_4927,N_4825);
and U5188 (N_5188,N_4824,N_4978);
nor U5189 (N_5189,N_4846,N_4993);
nor U5190 (N_5190,N_4838,N_4910);
or U5191 (N_5191,N_4902,N_4928);
nor U5192 (N_5192,N_4854,N_4969);
or U5193 (N_5193,N_4962,N_4850);
or U5194 (N_5194,N_4918,N_4855);
nor U5195 (N_5195,N_4965,N_4929);
nand U5196 (N_5196,N_4939,N_4858);
and U5197 (N_5197,N_4880,N_4973);
or U5198 (N_5198,N_4992,N_4969);
and U5199 (N_5199,N_4962,N_4956);
nor U5200 (N_5200,N_5171,N_5109);
nor U5201 (N_5201,N_5154,N_5048);
nor U5202 (N_5202,N_5167,N_5172);
nor U5203 (N_5203,N_5168,N_5044);
or U5204 (N_5204,N_5005,N_5142);
nor U5205 (N_5205,N_5121,N_5170);
or U5206 (N_5206,N_5122,N_5021);
nor U5207 (N_5207,N_5059,N_5194);
nor U5208 (N_5208,N_5066,N_5153);
and U5209 (N_5209,N_5099,N_5141);
nor U5210 (N_5210,N_5051,N_5174);
nor U5211 (N_5211,N_5057,N_5054);
and U5212 (N_5212,N_5037,N_5101);
and U5213 (N_5213,N_5079,N_5187);
and U5214 (N_5214,N_5163,N_5190);
nand U5215 (N_5215,N_5148,N_5095);
nor U5216 (N_5216,N_5151,N_5127);
nand U5217 (N_5217,N_5150,N_5160);
or U5218 (N_5218,N_5115,N_5126);
nor U5219 (N_5219,N_5182,N_5119);
nor U5220 (N_5220,N_5158,N_5178);
or U5221 (N_5221,N_5123,N_5047);
nand U5222 (N_5222,N_5164,N_5030);
or U5223 (N_5223,N_5087,N_5009);
nand U5224 (N_5224,N_5188,N_5149);
or U5225 (N_5225,N_5189,N_5091);
and U5226 (N_5226,N_5117,N_5084);
nor U5227 (N_5227,N_5036,N_5092);
and U5228 (N_5228,N_5019,N_5027);
or U5229 (N_5229,N_5146,N_5103);
nand U5230 (N_5230,N_5139,N_5152);
nand U5231 (N_5231,N_5007,N_5014);
nand U5232 (N_5232,N_5008,N_5157);
or U5233 (N_5233,N_5096,N_5025);
or U5234 (N_5234,N_5055,N_5105);
or U5235 (N_5235,N_5018,N_5068);
nor U5236 (N_5236,N_5196,N_5015);
or U5237 (N_5237,N_5063,N_5069);
nor U5238 (N_5238,N_5062,N_5088);
and U5239 (N_5239,N_5137,N_5041);
nor U5240 (N_5240,N_5026,N_5089);
nand U5241 (N_5241,N_5046,N_5045);
nand U5242 (N_5242,N_5136,N_5012);
nor U5243 (N_5243,N_5024,N_5118);
nand U5244 (N_5244,N_5074,N_5011);
xnor U5245 (N_5245,N_5097,N_5071);
and U5246 (N_5246,N_5112,N_5052);
nand U5247 (N_5247,N_5114,N_5078);
or U5248 (N_5248,N_5085,N_5162);
nor U5249 (N_5249,N_5191,N_5001);
nand U5250 (N_5250,N_5133,N_5077);
or U5251 (N_5251,N_5013,N_5080);
and U5252 (N_5252,N_5017,N_5042);
nor U5253 (N_5253,N_5140,N_5199);
nor U5254 (N_5254,N_5006,N_5145);
nand U5255 (N_5255,N_5143,N_5072);
and U5256 (N_5256,N_5111,N_5049);
nor U5257 (N_5257,N_5020,N_5093);
and U5258 (N_5258,N_5169,N_5147);
and U5259 (N_5259,N_5124,N_5193);
nor U5260 (N_5260,N_5022,N_5129);
nor U5261 (N_5261,N_5086,N_5198);
nor U5262 (N_5262,N_5156,N_5065);
or U5263 (N_5263,N_5083,N_5107);
nor U5264 (N_5264,N_5179,N_5100);
or U5265 (N_5265,N_5132,N_5184);
and U5266 (N_5266,N_5023,N_5177);
nand U5267 (N_5267,N_5050,N_5134);
and U5268 (N_5268,N_5186,N_5035);
nand U5269 (N_5269,N_5128,N_5192);
nor U5270 (N_5270,N_5038,N_5028);
or U5271 (N_5271,N_5061,N_5081);
or U5272 (N_5272,N_5098,N_5183);
and U5273 (N_5273,N_5004,N_5120);
or U5274 (N_5274,N_5175,N_5135);
nand U5275 (N_5275,N_5029,N_5075);
or U5276 (N_5276,N_5060,N_5166);
and U5277 (N_5277,N_5144,N_5040);
nand U5278 (N_5278,N_5104,N_5033);
or U5279 (N_5279,N_5161,N_5173);
nor U5280 (N_5280,N_5106,N_5180);
and U5281 (N_5281,N_5056,N_5116);
and U5282 (N_5282,N_5064,N_5053);
and U5283 (N_5283,N_5016,N_5031);
nor U5284 (N_5284,N_5197,N_5165);
nor U5285 (N_5285,N_5058,N_5003);
nor U5286 (N_5286,N_5076,N_5113);
nor U5287 (N_5287,N_5108,N_5090);
or U5288 (N_5288,N_5002,N_5110);
and U5289 (N_5289,N_5130,N_5070);
nor U5290 (N_5290,N_5032,N_5125);
nor U5291 (N_5291,N_5195,N_5185);
nand U5292 (N_5292,N_5082,N_5176);
or U5293 (N_5293,N_5067,N_5094);
nand U5294 (N_5294,N_5043,N_5010);
nand U5295 (N_5295,N_5039,N_5102);
nand U5296 (N_5296,N_5000,N_5155);
or U5297 (N_5297,N_5131,N_5034);
nor U5298 (N_5298,N_5073,N_5181);
nor U5299 (N_5299,N_5159,N_5138);
nor U5300 (N_5300,N_5082,N_5168);
nand U5301 (N_5301,N_5133,N_5180);
and U5302 (N_5302,N_5019,N_5130);
nand U5303 (N_5303,N_5018,N_5022);
nand U5304 (N_5304,N_5039,N_5133);
or U5305 (N_5305,N_5005,N_5194);
or U5306 (N_5306,N_5095,N_5010);
nor U5307 (N_5307,N_5042,N_5122);
nand U5308 (N_5308,N_5131,N_5132);
nor U5309 (N_5309,N_5145,N_5077);
nand U5310 (N_5310,N_5151,N_5100);
nand U5311 (N_5311,N_5128,N_5178);
and U5312 (N_5312,N_5196,N_5186);
nand U5313 (N_5313,N_5014,N_5015);
nand U5314 (N_5314,N_5111,N_5075);
or U5315 (N_5315,N_5045,N_5074);
and U5316 (N_5316,N_5188,N_5071);
nand U5317 (N_5317,N_5124,N_5179);
and U5318 (N_5318,N_5149,N_5115);
nor U5319 (N_5319,N_5188,N_5077);
nand U5320 (N_5320,N_5195,N_5198);
nor U5321 (N_5321,N_5060,N_5078);
and U5322 (N_5322,N_5014,N_5077);
nand U5323 (N_5323,N_5170,N_5158);
nand U5324 (N_5324,N_5168,N_5134);
nand U5325 (N_5325,N_5077,N_5118);
or U5326 (N_5326,N_5138,N_5190);
or U5327 (N_5327,N_5122,N_5032);
nor U5328 (N_5328,N_5147,N_5181);
and U5329 (N_5329,N_5079,N_5032);
and U5330 (N_5330,N_5099,N_5049);
and U5331 (N_5331,N_5020,N_5133);
and U5332 (N_5332,N_5115,N_5102);
nand U5333 (N_5333,N_5182,N_5092);
and U5334 (N_5334,N_5175,N_5074);
nor U5335 (N_5335,N_5164,N_5053);
nand U5336 (N_5336,N_5016,N_5123);
nor U5337 (N_5337,N_5192,N_5086);
or U5338 (N_5338,N_5003,N_5071);
nand U5339 (N_5339,N_5109,N_5067);
nand U5340 (N_5340,N_5032,N_5147);
or U5341 (N_5341,N_5184,N_5112);
and U5342 (N_5342,N_5151,N_5054);
and U5343 (N_5343,N_5074,N_5162);
nand U5344 (N_5344,N_5066,N_5040);
nor U5345 (N_5345,N_5184,N_5134);
nor U5346 (N_5346,N_5090,N_5064);
or U5347 (N_5347,N_5082,N_5120);
nor U5348 (N_5348,N_5184,N_5011);
nor U5349 (N_5349,N_5144,N_5112);
and U5350 (N_5350,N_5177,N_5182);
or U5351 (N_5351,N_5188,N_5175);
nor U5352 (N_5352,N_5194,N_5076);
nand U5353 (N_5353,N_5160,N_5004);
and U5354 (N_5354,N_5098,N_5008);
nor U5355 (N_5355,N_5026,N_5103);
nand U5356 (N_5356,N_5125,N_5052);
nand U5357 (N_5357,N_5147,N_5078);
and U5358 (N_5358,N_5134,N_5091);
nand U5359 (N_5359,N_5046,N_5104);
nand U5360 (N_5360,N_5046,N_5184);
and U5361 (N_5361,N_5040,N_5192);
and U5362 (N_5362,N_5103,N_5085);
or U5363 (N_5363,N_5132,N_5035);
nand U5364 (N_5364,N_5195,N_5044);
nand U5365 (N_5365,N_5041,N_5198);
nand U5366 (N_5366,N_5091,N_5133);
nor U5367 (N_5367,N_5099,N_5081);
nand U5368 (N_5368,N_5104,N_5188);
and U5369 (N_5369,N_5107,N_5060);
nor U5370 (N_5370,N_5008,N_5164);
nor U5371 (N_5371,N_5143,N_5167);
or U5372 (N_5372,N_5123,N_5030);
nand U5373 (N_5373,N_5088,N_5165);
nand U5374 (N_5374,N_5136,N_5129);
nand U5375 (N_5375,N_5165,N_5091);
nor U5376 (N_5376,N_5060,N_5034);
nand U5377 (N_5377,N_5001,N_5139);
or U5378 (N_5378,N_5042,N_5031);
and U5379 (N_5379,N_5087,N_5076);
nor U5380 (N_5380,N_5133,N_5189);
nand U5381 (N_5381,N_5129,N_5197);
nor U5382 (N_5382,N_5001,N_5019);
nor U5383 (N_5383,N_5046,N_5042);
nand U5384 (N_5384,N_5046,N_5194);
or U5385 (N_5385,N_5090,N_5026);
nor U5386 (N_5386,N_5120,N_5118);
and U5387 (N_5387,N_5003,N_5098);
and U5388 (N_5388,N_5143,N_5096);
or U5389 (N_5389,N_5078,N_5143);
nand U5390 (N_5390,N_5174,N_5141);
and U5391 (N_5391,N_5061,N_5050);
and U5392 (N_5392,N_5065,N_5076);
or U5393 (N_5393,N_5041,N_5012);
and U5394 (N_5394,N_5023,N_5076);
nor U5395 (N_5395,N_5011,N_5094);
or U5396 (N_5396,N_5122,N_5098);
nor U5397 (N_5397,N_5007,N_5055);
xor U5398 (N_5398,N_5009,N_5052);
nor U5399 (N_5399,N_5123,N_5006);
and U5400 (N_5400,N_5250,N_5306);
nand U5401 (N_5401,N_5256,N_5384);
or U5402 (N_5402,N_5357,N_5288);
nor U5403 (N_5403,N_5302,N_5351);
and U5404 (N_5404,N_5371,N_5322);
nor U5405 (N_5405,N_5380,N_5280);
and U5406 (N_5406,N_5221,N_5205);
nor U5407 (N_5407,N_5346,N_5273);
nor U5408 (N_5408,N_5212,N_5318);
or U5409 (N_5409,N_5342,N_5233);
xnor U5410 (N_5410,N_5382,N_5214);
nand U5411 (N_5411,N_5276,N_5309);
nor U5412 (N_5412,N_5366,N_5249);
or U5413 (N_5413,N_5210,N_5348);
nor U5414 (N_5414,N_5218,N_5230);
nor U5415 (N_5415,N_5264,N_5278);
and U5416 (N_5416,N_5245,N_5202);
nand U5417 (N_5417,N_5364,N_5231);
and U5418 (N_5418,N_5332,N_5270);
and U5419 (N_5419,N_5227,N_5326);
or U5420 (N_5420,N_5283,N_5294);
and U5421 (N_5421,N_5395,N_5329);
nor U5422 (N_5422,N_5299,N_5258);
or U5423 (N_5423,N_5379,N_5293);
nor U5424 (N_5424,N_5338,N_5385);
or U5425 (N_5425,N_5307,N_5285);
and U5426 (N_5426,N_5207,N_5327);
or U5427 (N_5427,N_5303,N_5372);
or U5428 (N_5428,N_5263,N_5208);
or U5429 (N_5429,N_5229,N_5314);
nand U5430 (N_5430,N_5335,N_5315);
nand U5431 (N_5431,N_5267,N_5370);
nor U5432 (N_5432,N_5339,N_5203);
and U5433 (N_5433,N_5253,N_5320);
nor U5434 (N_5434,N_5246,N_5271);
nand U5435 (N_5435,N_5344,N_5397);
or U5436 (N_5436,N_5393,N_5305);
or U5437 (N_5437,N_5240,N_5247);
or U5438 (N_5438,N_5204,N_5308);
nand U5439 (N_5439,N_5312,N_5244);
nand U5440 (N_5440,N_5301,N_5228);
nand U5441 (N_5441,N_5289,N_5343);
or U5442 (N_5442,N_5238,N_5209);
nand U5443 (N_5443,N_5324,N_5296);
or U5444 (N_5444,N_5224,N_5388);
nor U5445 (N_5445,N_5259,N_5260);
nor U5446 (N_5446,N_5255,N_5359);
nand U5447 (N_5447,N_5376,N_5358);
nor U5448 (N_5448,N_5292,N_5341);
nor U5449 (N_5449,N_5236,N_5252);
and U5450 (N_5450,N_5353,N_5281);
or U5451 (N_5451,N_5323,N_5352);
and U5452 (N_5452,N_5396,N_5362);
or U5453 (N_5453,N_5356,N_5219);
or U5454 (N_5454,N_5297,N_5391);
xnor U5455 (N_5455,N_5257,N_5206);
nand U5456 (N_5456,N_5217,N_5389);
and U5457 (N_5457,N_5321,N_5331);
nor U5458 (N_5458,N_5235,N_5347);
or U5459 (N_5459,N_5242,N_5268);
and U5460 (N_5460,N_5334,N_5248);
and U5461 (N_5461,N_5355,N_5354);
and U5462 (N_5462,N_5226,N_5232);
and U5463 (N_5463,N_5274,N_5237);
nand U5464 (N_5464,N_5298,N_5216);
nor U5465 (N_5465,N_5361,N_5386);
and U5466 (N_5466,N_5375,N_5313);
nand U5467 (N_5467,N_5241,N_5215);
or U5468 (N_5468,N_5265,N_5310);
nand U5469 (N_5469,N_5201,N_5377);
nor U5470 (N_5470,N_5390,N_5374);
or U5471 (N_5471,N_5287,N_5398);
or U5472 (N_5472,N_5381,N_5319);
nand U5473 (N_5473,N_5211,N_5261);
nor U5474 (N_5474,N_5311,N_5330);
and U5475 (N_5475,N_5222,N_5392);
and U5476 (N_5476,N_5394,N_5360);
nand U5477 (N_5477,N_5291,N_5269);
nor U5478 (N_5478,N_5282,N_5387);
nand U5479 (N_5479,N_5378,N_5266);
and U5480 (N_5480,N_5213,N_5363);
or U5481 (N_5481,N_5345,N_5223);
or U5482 (N_5482,N_5349,N_5239);
and U5483 (N_5483,N_5304,N_5383);
and U5484 (N_5484,N_5336,N_5275);
nor U5485 (N_5485,N_5369,N_5316);
and U5486 (N_5486,N_5251,N_5317);
nand U5487 (N_5487,N_5340,N_5290);
and U5488 (N_5488,N_5328,N_5262);
and U5489 (N_5489,N_5295,N_5367);
or U5490 (N_5490,N_5337,N_5243);
nand U5491 (N_5491,N_5254,N_5277);
or U5492 (N_5492,N_5373,N_5365);
and U5493 (N_5493,N_5279,N_5325);
nand U5494 (N_5494,N_5300,N_5286);
nor U5495 (N_5495,N_5333,N_5200);
and U5496 (N_5496,N_5399,N_5234);
nand U5497 (N_5497,N_5284,N_5225);
nor U5498 (N_5498,N_5220,N_5272);
nor U5499 (N_5499,N_5368,N_5350);
nor U5500 (N_5500,N_5364,N_5327);
or U5501 (N_5501,N_5258,N_5322);
or U5502 (N_5502,N_5348,N_5316);
or U5503 (N_5503,N_5267,N_5315);
nand U5504 (N_5504,N_5280,N_5231);
nor U5505 (N_5505,N_5333,N_5224);
and U5506 (N_5506,N_5214,N_5330);
and U5507 (N_5507,N_5338,N_5365);
nor U5508 (N_5508,N_5379,N_5263);
or U5509 (N_5509,N_5367,N_5218);
and U5510 (N_5510,N_5294,N_5335);
or U5511 (N_5511,N_5265,N_5248);
or U5512 (N_5512,N_5227,N_5211);
nand U5513 (N_5513,N_5230,N_5332);
and U5514 (N_5514,N_5225,N_5221);
nand U5515 (N_5515,N_5343,N_5380);
and U5516 (N_5516,N_5342,N_5217);
or U5517 (N_5517,N_5264,N_5325);
nand U5518 (N_5518,N_5374,N_5245);
nor U5519 (N_5519,N_5291,N_5348);
and U5520 (N_5520,N_5204,N_5246);
nor U5521 (N_5521,N_5308,N_5290);
nand U5522 (N_5522,N_5355,N_5379);
and U5523 (N_5523,N_5323,N_5312);
nor U5524 (N_5524,N_5320,N_5219);
or U5525 (N_5525,N_5392,N_5219);
nand U5526 (N_5526,N_5393,N_5334);
nor U5527 (N_5527,N_5376,N_5316);
and U5528 (N_5528,N_5209,N_5251);
or U5529 (N_5529,N_5372,N_5254);
nand U5530 (N_5530,N_5282,N_5211);
nand U5531 (N_5531,N_5337,N_5216);
and U5532 (N_5532,N_5346,N_5374);
nand U5533 (N_5533,N_5258,N_5289);
nor U5534 (N_5534,N_5300,N_5397);
and U5535 (N_5535,N_5243,N_5319);
or U5536 (N_5536,N_5369,N_5333);
or U5537 (N_5537,N_5274,N_5344);
and U5538 (N_5538,N_5279,N_5383);
nor U5539 (N_5539,N_5298,N_5251);
and U5540 (N_5540,N_5390,N_5267);
nor U5541 (N_5541,N_5200,N_5394);
nand U5542 (N_5542,N_5369,N_5224);
nor U5543 (N_5543,N_5254,N_5215);
or U5544 (N_5544,N_5200,N_5268);
or U5545 (N_5545,N_5319,N_5358);
or U5546 (N_5546,N_5374,N_5215);
nor U5547 (N_5547,N_5314,N_5235);
nor U5548 (N_5548,N_5385,N_5280);
or U5549 (N_5549,N_5288,N_5389);
and U5550 (N_5550,N_5297,N_5226);
and U5551 (N_5551,N_5339,N_5271);
xor U5552 (N_5552,N_5396,N_5202);
and U5553 (N_5553,N_5316,N_5258);
or U5554 (N_5554,N_5280,N_5319);
nand U5555 (N_5555,N_5264,N_5241);
nor U5556 (N_5556,N_5370,N_5357);
nor U5557 (N_5557,N_5377,N_5229);
and U5558 (N_5558,N_5398,N_5376);
nand U5559 (N_5559,N_5345,N_5279);
nand U5560 (N_5560,N_5208,N_5392);
or U5561 (N_5561,N_5217,N_5209);
nand U5562 (N_5562,N_5331,N_5296);
nor U5563 (N_5563,N_5317,N_5315);
and U5564 (N_5564,N_5277,N_5283);
nand U5565 (N_5565,N_5293,N_5364);
nor U5566 (N_5566,N_5270,N_5230);
nand U5567 (N_5567,N_5269,N_5319);
nand U5568 (N_5568,N_5390,N_5254);
nor U5569 (N_5569,N_5398,N_5297);
and U5570 (N_5570,N_5318,N_5374);
nand U5571 (N_5571,N_5386,N_5314);
and U5572 (N_5572,N_5212,N_5247);
nand U5573 (N_5573,N_5308,N_5222);
nor U5574 (N_5574,N_5328,N_5207);
nand U5575 (N_5575,N_5367,N_5200);
nor U5576 (N_5576,N_5287,N_5314);
nand U5577 (N_5577,N_5265,N_5364);
or U5578 (N_5578,N_5318,N_5280);
nand U5579 (N_5579,N_5330,N_5290);
or U5580 (N_5580,N_5348,N_5387);
or U5581 (N_5581,N_5321,N_5386);
and U5582 (N_5582,N_5395,N_5204);
nand U5583 (N_5583,N_5345,N_5315);
and U5584 (N_5584,N_5315,N_5356);
nand U5585 (N_5585,N_5376,N_5229);
nor U5586 (N_5586,N_5356,N_5343);
xnor U5587 (N_5587,N_5245,N_5333);
nor U5588 (N_5588,N_5281,N_5375);
nand U5589 (N_5589,N_5333,N_5308);
and U5590 (N_5590,N_5202,N_5222);
nand U5591 (N_5591,N_5322,N_5270);
or U5592 (N_5592,N_5264,N_5280);
nand U5593 (N_5593,N_5280,N_5246);
or U5594 (N_5594,N_5224,N_5268);
nand U5595 (N_5595,N_5329,N_5353);
or U5596 (N_5596,N_5283,N_5329);
xnor U5597 (N_5597,N_5365,N_5309);
nand U5598 (N_5598,N_5207,N_5393);
nor U5599 (N_5599,N_5380,N_5224);
and U5600 (N_5600,N_5473,N_5442);
nor U5601 (N_5601,N_5434,N_5500);
or U5602 (N_5602,N_5475,N_5440);
or U5603 (N_5603,N_5496,N_5418);
or U5604 (N_5604,N_5493,N_5443);
nor U5605 (N_5605,N_5487,N_5590);
nand U5606 (N_5606,N_5447,N_5489);
or U5607 (N_5607,N_5520,N_5563);
nor U5608 (N_5608,N_5510,N_5547);
or U5609 (N_5609,N_5429,N_5458);
or U5610 (N_5610,N_5462,N_5559);
nand U5611 (N_5611,N_5457,N_5412);
or U5612 (N_5612,N_5555,N_5421);
nand U5613 (N_5613,N_5596,N_5595);
and U5614 (N_5614,N_5504,N_5545);
or U5615 (N_5615,N_5461,N_5539);
nand U5616 (N_5616,N_5594,N_5400);
xnor U5617 (N_5617,N_5542,N_5406);
nand U5618 (N_5618,N_5576,N_5466);
or U5619 (N_5619,N_5561,N_5407);
and U5620 (N_5620,N_5567,N_5578);
nand U5621 (N_5621,N_5544,N_5557);
and U5622 (N_5622,N_5509,N_5568);
nor U5623 (N_5623,N_5571,N_5413);
and U5624 (N_5624,N_5454,N_5591);
nor U5625 (N_5625,N_5404,N_5512);
nand U5626 (N_5626,N_5599,N_5564);
nand U5627 (N_5627,N_5452,N_5543);
xnor U5628 (N_5628,N_5515,N_5477);
nor U5629 (N_5629,N_5538,N_5472);
nor U5630 (N_5630,N_5436,N_5433);
or U5631 (N_5631,N_5451,N_5551);
nor U5632 (N_5632,N_5572,N_5587);
xor U5633 (N_5633,N_5536,N_5581);
nor U5634 (N_5634,N_5588,N_5492);
nor U5635 (N_5635,N_5507,N_5597);
or U5636 (N_5636,N_5584,N_5486);
nand U5637 (N_5637,N_5592,N_5468);
and U5638 (N_5638,N_5414,N_5476);
nor U5639 (N_5639,N_5502,N_5415);
or U5640 (N_5640,N_5430,N_5431);
nand U5641 (N_5641,N_5401,N_5582);
nor U5642 (N_5642,N_5437,N_5422);
and U5643 (N_5643,N_5419,N_5499);
nand U5644 (N_5644,N_5537,N_5425);
or U5645 (N_5645,N_5416,N_5549);
nor U5646 (N_5646,N_5426,N_5501);
or U5647 (N_5647,N_5575,N_5478);
and U5648 (N_5648,N_5491,N_5585);
and U5649 (N_5649,N_5448,N_5459);
or U5650 (N_5650,N_5471,N_5573);
nand U5651 (N_5651,N_5565,N_5410);
xnor U5652 (N_5652,N_5488,N_5562);
nor U5653 (N_5653,N_5424,N_5463);
nor U5654 (N_5654,N_5497,N_5558);
nand U5655 (N_5655,N_5552,N_5574);
or U5656 (N_5656,N_5479,N_5521);
nand U5657 (N_5657,N_5528,N_5405);
or U5658 (N_5658,N_5460,N_5534);
nor U5659 (N_5659,N_5540,N_5583);
or U5660 (N_5660,N_5550,N_5593);
nand U5661 (N_5661,N_5484,N_5456);
xnor U5662 (N_5662,N_5403,N_5511);
xor U5663 (N_5663,N_5439,N_5438);
nand U5664 (N_5664,N_5546,N_5522);
or U5665 (N_5665,N_5598,N_5560);
nor U5666 (N_5666,N_5481,N_5483);
nand U5667 (N_5667,N_5579,N_5408);
and U5668 (N_5668,N_5455,N_5519);
and U5669 (N_5669,N_5498,N_5427);
nand U5670 (N_5670,N_5589,N_5420);
nor U5671 (N_5671,N_5495,N_5432);
nand U5672 (N_5672,N_5535,N_5541);
and U5673 (N_5673,N_5465,N_5532);
or U5674 (N_5674,N_5554,N_5548);
and U5675 (N_5675,N_5469,N_5428);
nand U5676 (N_5676,N_5474,N_5523);
nand U5677 (N_5677,N_5417,N_5518);
and U5678 (N_5678,N_5530,N_5490);
or U5679 (N_5679,N_5508,N_5445);
nor U5680 (N_5680,N_5577,N_5525);
or U5681 (N_5681,N_5516,N_5450);
nand U5682 (N_5682,N_5506,N_5449);
or U5683 (N_5683,N_5529,N_5517);
nor U5684 (N_5684,N_5553,N_5435);
or U5685 (N_5685,N_5569,N_5467);
nand U5686 (N_5686,N_5453,N_5570);
nand U5687 (N_5687,N_5423,N_5446);
or U5688 (N_5688,N_5494,N_5411);
or U5689 (N_5689,N_5480,N_5527);
and U5690 (N_5690,N_5524,N_5556);
and U5691 (N_5691,N_5464,N_5514);
nor U5692 (N_5692,N_5444,N_5513);
and U5693 (N_5693,N_5441,N_5485);
xor U5694 (N_5694,N_5409,N_5531);
and U5695 (N_5695,N_5533,N_5586);
or U5696 (N_5696,N_5505,N_5580);
and U5697 (N_5697,N_5470,N_5566);
or U5698 (N_5698,N_5402,N_5482);
nor U5699 (N_5699,N_5526,N_5503);
nand U5700 (N_5700,N_5482,N_5420);
or U5701 (N_5701,N_5540,N_5539);
nand U5702 (N_5702,N_5413,N_5444);
nor U5703 (N_5703,N_5456,N_5594);
and U5704 (N_5704,N_5543,N_5440);
nor U5705 (N_5705,N_5535,N_5487);
nor U5706 (N_5706,N_5538,N_5550);
and U5707 (N_5707,N_5570,N_5491);
nor U5708 (N_5708,N_5597,N_5485);
and U5709 (N_5709,N_5522,N_5524);
or U5710 (N_5710,N_5492,N_5476);
and U5711 (N_5711,N_5418,N_5525);
nor U5712 (N_5712,N_5573,N_5549);
nand U5713 (N_5713,N_5596,N_5510);
nor U5714 (N_5714,N_5414,N_5528);
nand U5715 (N_5715,N_5557,N_5488);
or U5716 (N_5716,N_5463,N_5531);
nand U5717 (N_5717,N_5455,N_5430);
nor U5718 (N_5718,N_5558,N_5406);
or U5719 (N_5719,N_5567,N_5561);
nand U5720 (N_5720,N_5578,N_5446);
nand U5721 (N_5721,N_5485,N_5411);
nor U5722 (N_5722,N_5458,N_5553);
xnor U5723 (N_5723,N_5492,N_5599);
nor U5724 (N_5724,N_5442,N_5578);
or U5725 (N_5725,N_5572,N_5489);
nand U5726 (N_5726,N_5597,N_5590);
nor U5727 (N_5727,N_5416,N_5432);
nand U5728 (N_5728,N_5522,N_5412);
nor U5729 (N_5729,N_5589,N_5468);
or U5730 (N_5730,N_5549,N_5522);
nor U5731 (N_5731,N_5545,N_5534);
nor U5732 (N_5732,N_5483,N_5443);
nand U5733 (N_5733,N_5446,N_5591);
and U5734 (N_5734,N_5430,N_5451);
and U5735 (N_5735,N_5584,N_5407);
and U5736 (N_5736,N_5428,N_5409);
nor U5737 (N_5737,N_5414,N_5598);
nor U5738 (N_5738,N_5588,N_5559);
xor U5739 (N_5739,N_5520,N_5590);
and U5740 (N_5740,N_5493,N_5568);
nor U5741 (N_5741,N_5501,N_5545);
or U5742 (N_5742,N_5457,N_5442);
nor U5743 (N_5743,N_5421,N_5437);
and U5744 (N_5744,N_5528,N_5416);
nor U5745 (N_5745,N_5478,N_5453);
nand U5746 (N_5746,N_5445,N_5550);
or U5747 (N_5747,N_5464,N_5559);
and U5748 (N_5748,N_5422,N_5463);
nor U5749 (N_5749,N_5569,N_5454);
nand U5750 (N_5750,N_5576,N_5575);
nor U5751 (N_5751,N_5514,N_5505);
nand U5752 (N_5752,N_5468,N_5544);
and U5753 (N_5753,N_5594,N_5526);
and U5754 (N_5754,N_5462,N_5494);
or U5755 (N_5755,N_5514,N_5498);
or U5756 (N_5756,N_5599,N_5525);
and U5757 (N_5757,N_5579,N_5492);
nor U5758 (N_5758,N_5456,N_5567);
or U5759 (N_5759,N_5448,N_5436);
nor U5760 (N_5760,N_5572,N_5451);
or U5761 (N_5761,N_5438,N_5520);
and U5762 (N_5762,N_5478,N_5402);
or U5763 (N_5763,N_5435,N_5517);
and U5764 (N_5764,N_5451,N_5522);
and U5765 (N_5765,N_5476,N_5493);
and U5766 (N_5766,N_5454,N_5444);
and U5767 (N_5767,N_5518,N_5556);
or U5768 (N_5768,N_5417,N_5413);
nand U5769 (N_5769,N_5450,N_5460);
and U5770 (N_5770,N_5550,N_5476);
and U5771 (N_5771,N_5519,N_5473);
or U5772 (N_5772,N_5485,N_5536);
or U5773 (N_5773,N_5479,N_5599);
nand U5774 (N_5774,N_5417,N_5460);
and U5775 (N_5775,N_5548,N_5526);
and U5776 (N_5776,N_5494,N_5471);
nor U5777 (N_5777,N_5448,N_5524);
nor U5778 (N_5778,N_5406,N_5581);
nand U5779 (N_5779,N_5448,N_5570);
and U5780 (N_5780,N_5470,N_5576);
or U5781 (N_5781,N_5561,N_5511);
nand U5782 (N_5782,N_5415,N_5576);
nor U5783 (N_5783,N_5556,N_5585);
or U5784 (N_5784,N_5537,N_5449);
nor U5785 (N_5785,N_5523,N_5433);
nand U5786 (N_5786,N_5514,N_5556);
or U5787 (N_5787,N_5527,N_5497);
nand U5788 (N_5788,N_5496,N_5424);
and U5789 (N_5789,N_5410,N_5529);
nor U5790 (N_5790,N_5510,N_5421);
or U5791 (N_5791,N_5424,N_5493);
nor U5792 (N_5792,N_5545,N_5569);
or U5793 (N_5793,N_5416,N_5443);
or U5794 (N_5794,N_5492,N_5520);
nand U5795 (N_5795,N_5461,N_5521);
nand U5796 (N_5796,N_5584,N_5585);
nor U5797 (N_5797,N_5414,N_5595);
and U5798 (N_5798,N_5515,N_5590);
nor U5799 (N_5799,N_5584,N_5401);
and U5800 (N_5800,N_5690,N_5785);
xnor U5801 (N_5801,N_5645,N_5724);
or U5802 (N_5802,N_5654,N_5725);
and U5803 (N_5803,N_5699,N_5707);
and U5804 (N_5804,N_5795,N_5761);
or U5805 (N_5805,N_5762,N_5766);
and U5806 (N_5806,N_5744,N_5636);
nor U5807 (N_5807,N_5756,N_5774);
or U5808 (N_5808,N_5688,N_5771);
or U5809 (N_5809,N_5642,N_5747);
nand U5810 (N_5810,N_5748,N_5779);
nor U5811 (N_5811,N_5664,N_5663);
nor U5812 (N_5812,N_5709,N_5608);
or U5813 (N_5813,N_5635,N_5655);
and U5814 (N_5814,N_5691,N_5714);
nor U5815 (N_5815,N_5644,N_5629);
nor U5816 (N_5816,N_5799,N_5626);
or U5817 (N_5817,N_5677,N_5742);
and U5818 (N_5818,N_5759,N_5722);
nor U5819 (N_5819,N_5778,N_5648);
nor U5820 (N_5820,N_5777,N_5676);
or U5821 (N_5821,N_5702,N_5620);
nand U5822 (N_5822,N_5755,N_5773);
nor U5823 (N_5823,N_5662,N_5685);
nor U5824 (N_5824,N_5752,N_5751);
and U5825 (N_5825,N_5682,N_5753);
or U5826 (N_5826,N_5658,N_5730);
nor U5827 (N_5827,N_5765,N_5618);
nand U5828 (N_5828,N_5609,N_5772);
nor U5829 (N_5829,N_5704,N_5711);
nor U5830 (N_5830,N_5768,N_5652);
or U5831 (N_5831,N_5735,N_5729);
and U5832 (N_5832,N_5713,N_5697);
nand U5833 (N_5833,N_5604,N_5671);
and U5834 (N_5834,N_5675,N_5615);
and U5835 (N_5835,N_5775,N_5616);
nand U5836 (N_5836,N_5602,N_5625);
nand U5837 (N_5837,N_5732,N_5781);
or U5838 (N_5838,N_5605,N_5703);
nand U5839 (N_5839,N_5763,N_5784);
nand U5840 (N_5840,N_5670,N_5736);
or U5841 (N_5841,N_5681,N_5695);
or U5842 (N_5842,N_5678,N_5706);
and U5843 (N_5843,N_5617,N_5737);
and U5844 (N_5844,N_5760,N_5694);
nor U5845 (N_5845,N_5684,N_5791);
and U5846 (N_5846,N_5767,N_5728);
nor U5847 (N_5847,N_5666,N_5627);
nor U5848 (N_5848,N_5754,N_5749);
nand U5849 (N_5849,N_5698,N_5740);
or U5850 (N_5850,N_5672,N_5758);
nor U5851 (N_5851,N_5661,N_5628);
and U5852 (N_5852,N_5659,N_5668);
nand U5853 (N_5853,N_5601,N_5679);
and U5854 (N_5854,N_5794,N_5614);
nand U5855 (N_5855,N_5673,N_5712);
nor U5856 (N_5856,N_5798,N_5792);
nor U5857 (N_5857,N_5710,N_5610);
and U5858 (N_5858,N_5631,N_5633);
and U5859 (N_5859,N_5623,N_5776);
nand U5860 (N_5860,N_5669,N_5787);
nor U5861 (N_5861,N_5797,N_5632);
or U5862 (N_5862,N_5793,N_5640);
nand U5863 (N_5863,N_5733,N_5716);
nor U5864 (N_5864,N_5790,N_5650);
nand U5865 (N_5865,N_5750,N_5731);
nor U5866 (N_5866,N_5783,N_5700);
or U5867 (N_5867,N_5622,N_5674);
nand U5868 (N_5868,N_5660,N_5789);
nor U5869 (N_5869,N_5680,N_5746);
nor U5870 (N_5870,N_5739,N_5769);
nand U5871 (N_5871,N_5600,N_5721);
nand U5872 (N_5872,N_5653,N_5720);
nand U5873 (N_5873,N_5630,N_5646);
nand U5874 (N_5874,N_5612,N_5786);
nand U5875 (N_5875,N_5667,N_5613);
or U5876 (N_5876,N_5723,N_5656);
and U5877 (N_5877,N_5782,N_5649);
nand U5878 (N_5878,N_5726,N_5764);
nand U5879 (N_5879,N_5692,N_5686);
nor U5880 (N_5880,N_5718,N_5705);
nor U5881 (N_5881,N_5780,N_5745);
nor U5882 (N_5882,N_5641,N_5619);
or U5883 (N_5883,N_5611,N_5643);
nand U5884 (N_5884,N_5624,N_5743);
or U5885 (N_5885,N_5701,N_5606);
or U5886 (N_5886,N_5741,N_5715);
and U5887 (N_5887,N_5693,N_5757);
or U5888 (N_5888,N_5717,N_5770);
nand U5889 (N_5889,N_5665,N_5708);
and U5890 (N_5890,N_5796,N_5657);
nand U5891 (N_5891,N_5621,N_5603);
nor U5892 (N_5892,N_5638,N_5687);
or U5893 (N_5893,N_5683,N_5719);
nand U5894 (N_5894,N_5738,N_5647);
and U5895 (N_5895,N_5696,N_5651);
and U5896 (N_5896,N_5634,N_5788);
nor U5897 (N_5897,N_5637,N_5607);
and U5898 (N_5898,N_5689,N_5734);
nand U5899 (N_5899,N_5727,N_5639);
or U5900 (N_5900,N_5681,N_5655);
nor U5901 (N_5901,N_5665,N_5762);
and U5902 (N_5902,N_5752,N_5614);
nor U5903 (N_5903,N_5708,N_5641);
nor U5904 (N_5904,N_5635,N_5662);
nand U5905 (N_5905,N_5676,N_5718);
or U5906 (N_5906,N_5698,N_5739);
or U5907 (N_5907,N_5756,N_5761);
and U5908 (N_5908,N_5692,N_5780);
nand U5909 (N_5909,N_5799,N_5616);
or U5910 (N_5910,N_5762,N_5654);
and U5911 (N_5911,N_5614,N_5637);
or U5912 (N_5912,N_5643,N_5616);
or U5913 (N_5913,N_5639,N_5689);
nand U5914 (N_5914,N_5753,N_5717);
nand U5915 (N_5915,N_5603,N_5704);
or U5916 (N_5916,N_5727,N_5603);
nand U5917 (N_5917,N_5640,N_5714);
and U5918 (N_5918,N_5793,N_5620);
nor U5919 (N_5919,N_5730,N_5768);
and U5920 (N_5920,N_5785,N_5794);
nand U5921 (N_5921,N_5675,N_5745);
nor U5922 (N_5922,N_5696,N_5781);
nor U5923 (N_5923,N_5630,N_5772);
or U5924 (N_5924,N_5665,N_5615);
nand U5925 (N_5925,N_5791,N_5630);
or U5926 (N_5926,N_5737,N_5702);
or U5927 (N_5927,N_5682,N_5673);
nor U5928 (N_5928,N_5734,N_5776);
nand U5929 (N_5929,N_5792,N_5750);
or U5930 (N_5930,N_5633,N_5626);
nand U5931 (N_5931,N_5717,N_5642);
nand U5932 (N_5932,N_5710,N_5773);
nand U5933 (N_5933,N_5784,N_5632);
or U5934 (N_5934,N_5787,N_5789);
and U5935 (N_5935,N_5665,N_5673);
nor U5936 (N_5936,N_5666,N_5616);
nand U5937 (N_5937,N_5746,N_5639);
and U5938 (N_5938,N_5654,N_5624);
or U5939 (N_5939,N_5617,N_5756);
nand U5940 (N_5940,N_5760,N_5665);
nand U5941 (N_5941,N_5636,N_5758);
and U5942 (N_5942,N_5672,N_5707);
nand U5943 (N_5943,N_5638,N_5718);
nand U5944 (N_5944,N_5743,N_5686);
nand U5945 (N_5945,N_5766,N_5792);
or U5946 (N_5946,N_5632,N_5711);
nand U5947 (N_5947,N_5702,N_5685);
and U5948 (N_5948,N_5602,N_5777);
and U5949 (N_5949,N_5631,N_5640);
nor U5950 (N_5950,N_5722,N_5746);
or U5951 (N_5951,N_5656,N_5756);
nand U5952 (N_5952,N_5604,N_5780);
nand U5953 (N_5953,N_5779,N_5623);
nor U5954 (N_5954,N_5743,N_5729);
nor U5955 (N_5955,N_5716,N_5705);
nor U5956 (N_5956,N_5722,N_5777);
or U5957 (N_5957,N_5748,N_5736);
and U5958 (N_5958,N_5707,N_5724);
and U5959 (N_5959,N_5726,N_5794);
nor U5960 (N_5960,N_5687,N_5701);
and U5961 (N_5961,N_5605,N_5658);
nand U5962 (N_5962,N_5742,N_5799);
and U5963 (N_5963,N_5758,N_5623);
nand U5964 (N_5964,N_5778,N_5634);
nand U5965 (N_5965,N_5613,N_5726);
nand U5966 (N_5966,N_5728,N_5669);
or U5967 (N_5967,N_5715,N_5764);
or U5968 (N_5968,N_5770,N_5629);
xnor U5969 (N_5969,N_5727,N_5707);
nand U5970 (N_5970,N_5637,N_5695);
nor U5971 (N_5971,N_5755,N_5682);
nand U5972 (N_5972,N_5617,N_5749);
and U5973 (N_5973,N_5711,N_5772);
nand U5974 (N_5974,N_5748,N_5640);
nor U5975 (N_5975,N_5783,N_5773);
nor U5976 (N_5976,N_5756,N_5697);
nand U5977 (N_5977,N_5680,N_5726);
or U5978 (N_5978,N_5762,N_5700);
nor U5979 (N_5979,N_5606,N_5671);
nor U5980 (N_5980,N_5741,N_5726);
or U5981 (N_5981,N_5655,N_5676);
nand U5982 (N_5982,N_5685,N_5790);
or U5983 (N_5983,N_5643,N_5618);
and U5984 (N_5984,N_5671,N_5633);
xnor U5985 (N_5985,N_5630,N_5750);
nor U5986 (N_5986,N_5606,N_5608);
and U5987 (N_5987,N_5621,N_5715);
or U5988 (N_5988,N_5766,N_5625);
or U5989 (N_5989,N_5632,N_5719);
and U5990 (N_5990,N_5770,N_5748);
or U5991 (N_5991,N_5733,N_5616);
nor U5992 (N_5992,N_5614,N_5796);
and U5993 (N_5993,N_5693,N_5623);
nor U5994 (N_5994,N_5613,N_5778);
nand U5995 (N_5995,N_5731,N_5696);
nor U5996 (N_5996,N_5654,N_5630);
nor U5997 (N_5997,N_5714,N_5681);
or U5998 (N_5998,N_5759,N_5703);
nor U5999 (N_5999,N_5605,N_5756);
and U6000 (N_6000,N_5887,N_5968);
or U6001 (N_6001,N_5970,N_5830);
or U6002 (N_6002,N_5950,N_5923);
nand U6003 (N_6003,N_5946,N_5891);
nor U6004 (N_6004,N_5910,N_5945);
nor U6005 (N_6005,N_5850,N_5875);
or U6006 (N_6006,N_5938,N_5909);
nor U6007 (N_6007,N_5904,N_5852);
nor U6008 (N_6008,N_5930,N_5984);
or U6009 (N_6009,N_5884,N_5965);
nor U6010 (N_6010,N_5944,N_5870);
nor U6011 (N_6011,N_5882,N_5975);
nor U6012 (N_6012,N_5974,N_5892);
nand U6013 (N_6013,N_5841,N_5952);
nor U6014 (N_6014,N_5802,N_5929);
and U6015 (N_6015,N_5993,N_5804);
and U6016 (N_6016,N_5819,N_5885);
or U6017 (N_6017,N_5988,N_5898);
nand U6018 (N_6018,N_5911,N_5996);
and U6019 (N_6019,N_5880,N_5848);
or U6020 (N_6020,N_5955,N_5964);
and U6021 (N_6021,N_5801,N_5971);
and U6022 (N_6022,N_5847,N_5916);
or U6023 (N_6023,N_5833,N_5845);
nor U6024 (N_6024,N_5810,N_5991);
or U6025 (N_6025,N_5808,N_5969);
nor U6026 (N_6026,N_5978,N_5973);
nand U6027 (N_6027,N_5829,N_5824);
or U6028 (N_6028,N_5901,N_5919);
or U6029 (N_6029,N_5933,N_5865);
nor U6030 (N_6030,N_5989,N_5997);
nand U6031 (N_6031,N_5890,N_5921);
xor U6032 (N_6032,N_5873,N_5888);
nor U6033 (N_6033,N_5878,N_5920);
nand U6034 (N_6034,N_5867,N_5839);
and U6035 (N_6035,N_5939,N_5815);
nand U6036 (N_6036,N_5800,N_5995);
nor U6037 (N_6037,N_5924,N_5836);
nand U6038 (N_6038,N_5994,N_5877);
nor U6039 (N_6039,N_5931,N_5853);
nand U6040 (N_6040,N_5992,N_5840);
or U6041 (N_6041,N_5807,N_5897);
and U6042 (N_6042,N_5906,N_5863);
nor U6043 (N_6043,N_5983,N_5822);
nor U6044 (N_6044,N_5854,N_5941);
nand U6045 (N_6045,N_5957,N_5862);
nand U6046 (N_6046,N_5874,N_5951);
nor U6047 (N_6047,N_5861,N_5935);
or U6048 (N_6048,N_5954,N_5917);
nand U6049 (N_6049,N_5851,N_5826);
nor U6050 (N_6050,N_5817,N_5963);
nor U6051 (N_6051,N_5858,N_5942);
nand U6052 (N_6052,N_5979,N_5903);
nor U6053 (N_6053,N_5828,N_5816);
nor U6054 (N_6054,N_5895,N_5827);
and U6055 (N_6055,N_5925,N_5976);
nor U6056 (N_6056,N_5859,N_5820);
and U6057 (N_6057,N_5837,N_5985);
nand U6058 (N_6058,N_5868,N_5881);
nor U6059 (N_6059,N_5948,N_5928);
or U6060 (N_6060,N_5962,N_5855);
nand U6061 (N_6061,N_5894,N_5966);
and U6062 (N_6062,N_5932,N_5812);
and U6063 (N_6063,N_5835,N_5922);
or U6064 (N_6064,N_5866,N_5899);
and U6065 (N_6065,N_5960,N_5915);
nand U6066 (N_6066,N_5857,N_5846);
and U6067 (N_6067,N_5821,N_5918);
and U6068 (N_6068,N_5832,N_5981);
nand U6069 (N_6069,N_5889,N_5805);
and U6070 (N_6070,N_5907,N_5806);
nor U6071 (N_6071,N_5823,N_5914);
or U6072 (N_6072,N_5986,N_5809);
or U6073 (N_6073,N_5831,N_5912);
nand U6074 (N_6074,N_5956,N_5818);
or U6075 (N_6075,N_5825,N_5849);
or U6076 (N_6076,N_5813,N_5936);
or U6077 (N_6077,N_5959,N_5893);
nand U6078 (N_6078,N_5967,N_5998);
and U6079 (N_6079,N_5937,N_5872);
nand U6080 (N_6080,N_5977,N_5940);
and U6081 (N_6081,N_5902,N_5990);
nand U6082 (N_6082,N_5844,N_5908);
or U6083 (N_6083,N_5943,N_5814);
or U6084 (N_6084,N_5972,N_5860);
or U6085 (N_6085,N_5876,N_5838);
and U6086 (N_6086,N_5953,N_5834);
nor U6087 (N_6087,N_5913,N_5864);
nor U6088 (N_6088,N_5900,N_5926);
nor U6089 (N_6089,N_5947,N_5961);
or U6090 (N_6090,N_5842,N_5843);
nor U6091 (N_6091,N_5883,N_5999);
nor U6092 (N_6092,N_5980,N_5927);
nor U6093 (N_6093,N_5987,N_5949);
xor U6094 (N_6094,N_5803,N_5896);
nand U6095 (N_6095,N_5934,N_5869);
nor U6096 (N_6096,N_5871,N_5886);
or U6097 (N_6097,N_5879,N_5811);
nor U6098 (N_6098,N_5982,N_5856);
nor U6099 (N_6099,N_5905,N_5958);
or U6100 (N_6100,N_5813,N_5851);
nor U6101 (N_6101,N_5929,N_5884);
nor U6102 (N_6102,N_5943,N_5884);
and U6103 (N_6103,N_5971,N_5836);
nor U6104 (N_6104,N_5846,N_5914);
or U6105 (N_6105,N_5811,N_5926);
or U6106 (N_6106,N_5996,N_5986);
nand U6107 (N_6107,N_5812,N_5948);
or U6108 (N_6108,N_5867,N_5899);
and U6109 (N_6109,N_5938,N_5831);
nor U6110 (N_6110,N_5820,N_5937);
or U6111 (N_6111,N_5916,N_5859);
nor U6112 (N_6112,N_5804,N_5999);
nor U6113 (N_6113,N_5888,N_5938);
nand U6114 (N_6114,N_5838,N_5886);
or U6115 (N_6115,N_5940,N_5961);
and U6116 (N_6116,N_5861,N_5800);
and U6117 (N_6117,N_5848,N_5806);
or U6118 (N_6118,N_5845,N_5925);
nand U6119 (N_6119,N_5813,N_5815);
and U6120 (N_6120,N_5920,N_5916);
and U6121 (N_6121,N_5986,N_5850);
nor U6122 (N_6122,N_5945,N_5879);
nand U6123 (N_6123,N_5892,N_5823);
and U6124 (N_6124,N_5864,N_5856);
nand U6125 (N_6125,N_5824,N_5880);
and U6126 (N_6126,N_5929,N_5833);
and U6127 (N_6127,N_5968,N_5834);
and U6128 (N_6128,N_5805,N_5988);
and U6129 (N_6129,N_5832,N_5906);
nor U6130 (N_6130,N_5914,N_5989);
or U6131 (N_6131,N_5943,N_5955);
and U6132 (N_6132,N_5807,N_5962);
nand U6133 (N_6133,N_5936,N_5942);
and U6134 (N_6134,N_5913,N_5825);
nand U6135 (N_6135,N_5995,N_5971);
or U6136 (N_6136,N_5898,N_5943);
nor U6137 (N_6137,N_5827,N_5998);
nand U6138 (N_6138,N_5824,N_5896);
nand U6139 (N_6139,N_5906,N_5834);
nand U6140 (N_6140,N_5913,N_5892);
nor U6141 (N_6141,N_5800,N_5987);
nand U6142 (N_6142,N_5994,N_5899);
or U6143 (N_6143,N_5840,N_5901);
nor U6144 (N_6144,N_5976,N_5951);
and U6145 (N_6145,N_5853,N_5980);
nand U6146 (N_6146,N_5829,N_5925);
or U6147 (N_6147,N_5982,N_5821);
and U6148 (N_6148,N_5828,N_5916);
nand U6149 (N_6149,N_5940,N_5879);
or U6150 (N_6150,N_5902,N_5879);
or U6151 (N_6151,N_5816,N_5915);
nand U6152 (N_6152,N_5956,N_5844);
nor U6153 (N_6153,N_5916,N_5931);
nand U6154 (N_6154,N_5908,N_5930);
or U6155 (N_6155,N_5851,N_5936);
nand U6156 (N_6156,N_5915,N_5872);
or U6157 (N_6157,N_5906,N_5823);
nand U6158 (N_6158,N_5859,N_5944);
nor U6159 (N_6159,N_5977,N_5830);
and U6160 (N_6160,N_5808,N_5984);
and U6161 (N_6161,N_5984,N_5890);
nand U6162 (N_6162,N_5877,N_5919);
or U6163 (N_6163,N_5927,N_5823);
and U6164 (N_6164,N_5922,N_5926);
nor U6165 (N_6165,N_5845,N_5905);
and U6166 (N_6166,N_5864,N_5915);
and U6167 (N_6167,N_5846,N_5804);
nor U6168 (N_6168,N_5830,N_5912);
or U6169 (N_6169,N_5999,N_5909);
nand U6170 (N_6170,N_5971,N_5846);
nand U6171 (N_6171,N_5992,N_5868);
or U6172 (N_6172,N_5902,N_5873);
nor U6173 (N_6173,N_5874,N_5930);
and U6174 (N_6174,N_5973,N_5957);
or U6175 (N_6175,N_5877,N_5832);
nand U6176 (N_6176,N_5959,N_5980);
and U6177 (N_6177,N_5906,N_5888);
or U6178 (N_6178,N_5962,N_5933);
and U6179 (N_6179,N_5943,N_5912);
nor U6180 (N_6180,N_5918,N_5924);
xnor U6181 (N_6181,N_5981,N_5904);
nand U6182 (N_6182,N_5947,N_5949);
nor U6183 (N_6183,N_5896,N_5840);
nor U6184 (N_6184,N_5862,N_5815);
or U6185 (N_6185,N_5801,N_5869);
nor U6186 (N_6186,N_5972,N_5983);
nand U6187 (N_6187,N_5918,N_5859);
and U6188 (N_6188,N_5978,N_5867);
or U6189 (N_6189,N_5805,N_5915);
or U6190 (N_6190,N_5970,N_5928);
or U6191 (N_6191,N_5952,N_5804);
and U6192 (N_6192,N_5886,N_5876);
nor U6193 (N_6193,N_5892,N_5878);
or U6194 (N_6194,N_5851,N_5870);
and U6195 (N_6195,N_5871,N_5815);
or U6196 (N_6196,N_5856,N_5880);
or U6197 (N_6197,N_5831,N_5952);
nor U6198 (N_6198,N_5974,N_5824);
nor U6199 (N_6199,N_5885,N_5810);
or U6200 (N_6200,N_6149,N_6147);
nand U6201 (N_6201,N_6168,N_6085);
or U6202 (N_6202,N_6008,N_6089);
nor U6203 (N_6203,N_6025,N_6030);
nor U6204 (N_6204,N_6127,N_6121);
and U6205 (N_6205,N_6065,N_6022);
or U6206 (N_6206,N_6074,N_6036);
and U6207 (N_6207,N_6176,N_6175);
or U6208 (N_6208,N_6139,N_6100);
nor U6209 (N_6209,N_6161,N_6131);
and U6210 (N_6210,N_6106,N_6033);
nor U6211 (N_6211,N_6099,N_6152);
nand U6212 (N_6212,N_6086,N_6172);
or U6213 (N_6213,N_6058,N_6037);
or U6214 (N_6214,N_6108,N_6042);
and U6215 (N_6215,N_6116,N_6028);
nand U6216 (N_6216,N_6132,N_6047);
or U6217 (N_6217,N_6141,N_6120);
nand U6218 (N_6218,N_6077,N_6186);
nand U6219 (N_6219,N_6069,N_6024);
or U6220 (N_6220,N_6157,N_6073);
nand U6221 (N_6221,N_6000,N_6050);
nand U6222 (N_6222,N_6061,N_6193);
and U6223 (N_6223,N_6129,N_6166);
and U6224 (N_6224,N_6197,N_6124);
or U6225 (N_6225,N_6104,N_6144);
and U6226 (N_6226,N_6081,N_6192);
and U6227 (N_6227,N_6173,N_6079);
and U6228 (N_6228,N_6001,N_6041);
nand U6229 (N_6229,N_6184,N_6179);
nor U6230 (N_6230,N_6023,N_6138);
nand U6231 (N_6231,N_6133,N_6196);
nor U6232 (N_6232,N_6191,N_6169);
nor U6233 (N_6233,N_6002,N_6091);
nand U6234 (N_6234,N_6095,N_6060);
or U6235 (N_6235,N_6187,N_6031);
nor U6236 (N_6236,N_6123,N_6185);
nor U6237 (N_6237,N_6093,N_6087);
nor U6238 (N_6238,N_6017,N_6051);
nor U6239 (N_6239,N_6170,N_6150);
or U6240 (N_6240,N_6004,N_6083);
and U6241 (N_6241,N_6126,N_6135);
nand U6242 (N_6242,N_6034,N_6143);
and U6243 (N_6243,N_6071,N_6125);
or U6244 (N_6244,N_6199,N_6122);
nor U6245 (N_6245,N_6182,N_6183);
nand U6246 (N_6246,N_6165,N_6153);
nor U6247 (N_6247,N_6102,N_6059);
nor U6248 (N_6248,N_6067,N_6040);
nand U6249 (N_6249,N_6181,N_6090);
nand U6250 (N_6250,N_6076,N_6180);
or U6251 (N_6251,N_6020,N_6068);
and U6252 (N_6252,N_6109,N_6015);
or U6253 (N_6253,N_6174,N_6009);
nand U6254 (N_6254,N_6026,N_6107);
or U6255 (N_6255,N_6156,N_6136);
nor U6256 (N_6256,N_6029,N_6078);
and U6257 (N_6257,N_6048,N_6057);
xor U6258 (N_6258,N_6140,N_6103);
nand U6259 (N_6259,N_6072,N_6101);
or U6260 (N_6260,N_6055,N_6075);
or U6261 (N_6261,N_6084,N_6164);
or U6262 (N_6262,N_6114,N_6052);
nor U6263 (N_6263,N_6049,N_6011);
nor U6264 (N_6264,N_6092,N_6012);
nand U6265 (N_6265,N_6178,N_6006);
or U6266 (N_6266,N_6110,N_6162);
and U6267 (N_6267,N_6056,N_6128);
or U6268 (N_6268,N_6198,N_6188);
or U6269 (N_6269,N_6190,N_6044);
nand U6270 (N_6270,N_6046,N_6159);
and U6271 (N_6271,N_6054,N_6080);
or U6272 (N_6272,N_6007,N_6021);
or U6273 (N_6273,N_6115,N_6134);
or U6274 (N_6274,N_6154,N_6146);
nor U6275 (N_6275,N_6171,N_6119);
nand U6276 (N_6276,N_6113,N_6195);
nor U6277 (N_6277,N_6194,N_6066);
nand U6278 (N_6278,N_6094,N_6003);
or U6279 (N_6279,N_6151,N_6097);
nand U6280 (N_6280,N_6177,N_6105);
nand U6281 (N_6281,N_6160,N_6010);
nor U6282 (N_6282,N_6035,N_6148);
and U6283 (N_6283,N_6005,N_6142);
nand U6284 (N_6284,N_6043,N_6063);
xnor U6285 (N_6285,N_6112,N_6082);
nor U6286 (N_6286,N_6098,N_6070);
and U6287 (N_6287,N_6189,N_6062);
nand U6288 (N_6288,N_6032,N_6016);
and U6289 (N_6289,N_6027,N_6137);
or U6290 (N_6290,N_6038,N_6053);
or U6291 (N_6291,N_6111,N_6155);
nand U6292 (N_6292,N_6039,N_6013);
and U6293 (N_6293,N_6064,N_6019);
and U6294 (N_6294,N_6118,N_6167);
or U6295 (N_6295,N_6018,N_6145);
nand U6296 (N_6296,N_6158,N_6045);
and U6297 (N_6297,N_6130,N_6088);
or U6298 (N_6298,N_6163,N_6096);
nand U6299 (N_6299,N_6117,N_6014);
and U6300 (N_6300,N_6018,N_6056);
and U6301 (N_6301,N_6164,N_6186);
nor U6302 (N_6302,N_6123,N_6118);
and U6303 (N_6303,N_6182,N_6030);
nor U6304 (N_6304,N_6085,N_6005);
or U6305 (N_6305,N_6100,N_6021);
and U6306 (N_6306,N_6172,N_6106);
nand U6307 (N_6307,N_6151,N_6095);
and U6308 (N_6308,N_6046,N_6001);
or U6309 (N_6309,N_6100,N_6178);
nand U6310 (N_6310,N_6071,N_6122);
or U6311 (N_6311,N_6153,N_6175);
nor U6312 (N_6312,N_6145,N_6048);
nand U6313 (N_6313,N_6183,N_6134);
or U6314 (N_6314,N_6041,N_6072);
and U6315 (N_6315,N_6063,N_6049);
and U6316 (N_6316,N_6192,N_6078);
and U6317 (N_6317,N_6082,N_6053);
xor U6318 (N_6318,N_6117,N_6079);
nor U6319 (N_6319,N_6082,N_6105);
or U6320 (N_6320,N_6119,N_6043);
or U6321 (N_6321,N_6026,N_6113);
and U6322 (N_6322,N_6138,N_6095);
nand U6323 (N_6323,N_6031,N_6083);
nor U6324 (N_6324,N_6112,N_6152);
and U6325 (N_6325,N_6013,N_6122);
or U6326 (N_6326,N_6075,N_6094);
and U6327 (N_6327,N_6003,N_6182);
or U6328 (N_6328,N_6112,N_6143);
nor U6329 (N_6329,N_6036,N_6190);
or U6330 (N_6330,N_6143,N_6019);
nand U6331 (N_6331,N_6169,N_6020);
or U6332 (N_6332,N_6129,N_6157);
nand U6333 (N_6333,N_6124,N_6068);
and U6334 (N_6334,N_6179,N_6127);
and U6335 (N_6335,N_6026,N_6007);
nand U6336 (N_6336,N_6022,N_6170);
or U6337 (N_6337,N_6123,N_6040);
nand U6338 (N_6338,N_6143,N_6127);
nor U6339 (N_6339,N_6163,N_6168);
and U6340 (N_6340,N_6193,N_6171);
or U6341 (N_6341,N_6190,N_6140);
or U6342 (N_6342,N_6097,N_6158);
or U6343 (N_6343,N_6027,N_6155);
nor U6344 (N_6344,N_6120,N_6088);
or U6345 (N_6345,N_6056,N_6017);
nand U6346 (N_6346,N_6144,N_6102);
or U6347 (N_6347,N_6044,N_6013);
nand U6348 (N_6348,N_6139,N_6131);
nor U6349 (N_6349,N_6187,N_6138);
and U6350 (N_6350,N_6175,N_6065);
or U6351 (N_6351,N_6088,N_6107);
nor U6352 (N_6352,N_6151,N_6161);
nor U6353 (N_6353,N_6029,N_6071);
and U6354 (N_6354,N_6199,N_6028);
or U6355 (N_6355,N_6119,N_6049);
nor U6356 (N_6356,N_6106,N_6157);
and U6357 (N_6357,N_6050,N_6137);
and U6358 (N_6358,N_6140,N_6066);
and U6359 (N_6359,N_6145,N_6159);
nand U6360 (N_6360,N_6181,N_6116);
nor U6361 (N_6361,N_6082,N_6019);
or U6362 (N_6362,N_6147,N_6164);
or U6363 (N_6363,N_6153,N_6180);
nand U6364 (N_6364,N_6087,N_6085);
nand U6365 (N_6365,N_6024,N_6136);
or U6366 (N_6366,N_6111,N_6056);
or U6367 (N_6367,N_6051,N_6185);
nor U6368 (N_6368,N_6077,N_6044);
nand U6369 (N_6369,N_6054,N_6154);
and U6370 (N_6370,N_6123,N_6080);
nand U6371 (N_6371,N_6141,N_6088);
and U6372 (N_6372,N_6188,N_6041);
nand U6373 (N_6373,N_6017,N_6049);
nor U6374 (N_6374,N_6020,N_6132);
nand U6375 (N_6375,N_6049,N_6084);
nor U6376 (N_6376,N_6039,N_6001);
nor U6377 (N_6377,N_6004,N_6149);
nor U6378 (N_6378,N_6131,N_6003);
or U6379 (N_6379,N_6050,N_6080);
nand U6380 (N_6380,N_6144,N_6147);
nand U6381 (N_6381,N_6041,N_6156);
nand U6382 (N_6382,N_6141,N_6054);
and U6383 (N_6383,N_6131,N_6022);
or U6384 (N_6384,N_6015,N_6192);
nand U6385 (N_6385,N_6103,N_6189);
and U6386 (N_6386,N_6145,N_6054);
or U6387 (N_6387,N_6174,N_6082);
and U6388 (N_6388,N_6157,N_6051);
and U6389 (N_6389,N_6197,N_6027);
and U6390 (N_6390,N_6009,N_6185);
or U6391 (N_6391,N_6025,N_6044);
nor U6392 (N_6392,N_6188,N_6064);
or U6393 (N_6393,N_6121,N_6132);
nor U6394 (N_6394,N_6096,N_6057);
or U6395 (N_6395,N_6053,N_6080);
nor U6396 (N_6396,N_6091,N_6127);
and U6397 (N_6397,N_6052,N_6195);
and U6398 (N_6398,N_6016,N_6194);
nor U6399 (N_6399,N_6010,N_6011);
or U6400 (N_6400,N_6288,N_6206);
and U6401 (N_6401,N_6259,N_6325);
nor U6402 (N_6402,N_6349,N_6376);
or U6403 (N_6403,N_6204,N_6341);
nand U6404 (N_6404,N_6324,N_6332);
nor U6405 (N_6405,N_6342,N_6298);
nand U6406 (N_6406,N_6269,N_6382);
and U6407 (N_6407,N_6265,N_6356);
nand U6408 (N_6408,N_6303,N_6292);
or U6409 (N_6409,N_6366,N_6337);
nand U6410 (N_6410,N_6367,N_6217);
nand U6411 (N_6411,N_6363,N_6320);
and U6412 (N_6412,N_6245,N_6257);
and U6413 (N_6413,N_6392,N_6227);
or U6414 (N_6414,N_6237,N_6306);
nor U6415 (N_6415,N_6388,N_6314);
and U6416 (N_6416,N_6283,N_6358);
and U6417 (N_6417,N_6308,N_6322);
nor U6418 (N_6418,N_6290,N_6244);
and U6419 (N_6419,N_6255,N_6271);
or U6420 (N_6420,N_6397,N_6262);
or U6421 (N_6421,N_6264,N_6398);
nor U6422 (N_6422,N_6222,N_6246);
or U6423 (N_6423,N_6330,N_6256);
and U6424 (N_6424,N_6348,N_6225);
nor U6425 (N_6425,N_6234,N_6395);
or U6426 (N_6426,N_6281,N_6365);
nand U6427 (N_6427,N_6258,N_6364);
or U6428 (N_6428,N_6309,N_6353);
nor U6429 (N_6429,N_6241,N_6377);
or U6430 (N_6430,N_6384,N_6205);
nand U6431 (N_6431,N_6285,N_6385);
or U6432 (N_6432,N_6305,N_6374);
nand U6433 (N_6433,N_6310,N_6389);
nand U6434 (N_6434,N_6380,N_6360);
or U6435 (N_6435,N_6381,N_6211);
or U6436 (N_6436,N_6313,N_6216);
and U6437 (N_6437,N_6391,N_6201);
nand U6438 (N_6438,N_6316,N_6295);
or U6439 (N_6439,N_6243,N_6287);
nor U6440 (N_6440,N_6327,N_6253);
nand U6441 (N_6441,N_6239,N_6296);
nor U6442 (N_6442,N_6312,N_6268);
or U6443 (N_6443,N_6247,N_6351);
nand U6444 (N_6444,N_6266,N_6352);
or U6445 (N_6445,N_6319,N_6361);
or U6446 (N_6446,N_6307,N_6371);
and U6447 (N_6447,N_6236,N_6372);
nand U6448 (N_6448,N_6345,N_6209);
and U6449 (N_6449,N_6267,N_6386);
or U6450 (N_6450,N_6375,N_6242);
and U6451 (N_6451,N_6311,N_6362);
and U6452 (N_6452,N_6286,N_6354);
nor U6453 (N_6453,N_6214,N_6383);
nor U6454 (N_6454,N_6218,N_6202);
and U6455 (N_6455,N_6220,N_6334);
or U6456 (N_6456,N_6280,N_6219);
nand U6457 (N_6457,N_6321,N_6275);
nor U6458 (N_6458,N_6250,N_6333);
and U6459 (N_6459,N_6331,N_6291);
nor U6460 (N_6460,N_6323,N_6369);
nand U6461 (N_6461,N_6370,N_6347);
nor U6462 (N_6462,N_6273,N_6357);
nor U6463 (N_6463,N_6226,N_6221);
nor U6464 (N_6464,N_6252,N_6223);
nand U6465 (N_6465,N_6203,N_6260);
or U6466 (N_6466,N_6293,N_6289);
or U6467 (N_6467,N_6379,N_6329);
or U6468 (N_6468,N_6336,N_6317);
or U6469 (N_6469,N_6393,N_6278);
nor U6470 (N_6470,N_6390,N_6233);
or U6471 (N_6471,N_6373,N_6207);
and U6472 (N_6472,N_6208,N_6343);
or U6473 (N_6473,N_6378,N_6318);
nor U6474 (N_6474,N_6213,N_6344);
nand U6475 (N_6475,N_6228,N_6261);
nor U6476 (N_6476,N_6272,N_6279);
nor U6477 (N_6477,N_6224,N_6263);
or U6478 (N_6478,N_6210,N_6238);
and U6479 (N_6479,N_6282,N_6254);
nor U6480 (N_6480,N_6339,N_6368);
and U6481 (N_6481,N_6231,N_6215);
and U6482 (N_6482,N_6302,N_6230);
nor U6483 (N_6483,N_6249,N_6212);
nand U6484 (N_6484,N_6350,N_6251);
and U6485 (N_6485,N_6297,N_6355);
nor U6486 (N_6486,N_6346,N_6326);
or U6487 (N_6487,N_6232,N_6200);
and U6488 (N_6488,N_6248,N_6340);
nor U6489 (N_6489,N_6277,N_6338);
or U6490 (N_6490,N_6276,N_6299);
or U6491 (N_6491,N_6300,N_6335);
nor U6492 (N_6492,N_6315,N_6294);
and U6493 (N_6493,N_6328,N_6304);
or U6494 (N_6494,N_6387,N_6359);
or U6495 (N_6495,N_6235,N_6229);
and U6496 (N_6496,N_6270,N_6240);
nor U6497 (N_6497,N_6301,N_6394);
or U6498 (N_6498,N_6284,N_6274);
nor U6499 (N_6499,N_6396,N_6399);
nand U6500 (N_6500,N_6288,N_6289);
and U6501 (N_6501,N_6399,N_6297);
or U6502 (N_6502,N_6386,N_6226);
nor U6503 (N_6503,N_6380,N_6385);
nand U6504 (N_6504,N_6339,N_6253);
or U6505 (N_6505,N_6397,N_6275);
or U6506 (N_6506,N_6260,N_6242);
and U6507 (N_6507,N_6216,N_6242);
nor U6508 (N_6508,N_6263,N_6243);
nor U6509 (N_6509,N_6252,N_6321);
nand U6510 (N_6510,N_6245,N_6225);
or U6511 (N_6511,N_6365,N_6373);
or U6512 (N_6512,N_6389,N_6271);
or U6513 (N_6513,N_6273,N_6214);
nand U6514 (N_6514,N_6281,N_6317);
nand U6515 (N_6515,N_6240,N_6243);
xnor U6516 (N_6516,N_6265,N_6358);
and U6517 (N_6517,N_6355,N_6381);
or U6518 (N_6518,N_6347,N_6248);
nor U6519 (N_6519,N_6203,N_6206);
nand U6520 (N_6520,N_6238,N_6276);
nand U6521 (N_6521,N_6260,N_6280);
and U6522 (N_6522,N_6356,N_6390);
or U6523 (N_6523,N_6318,N_6205);
nand U6524 (N_6524,N_6248,N_6220);
and U6525 (N_6525,N_6385,N_6397);
or U6526 (N_6526,N_6321,N_6347);
nand U6527 (N_6527,N_6339,N_6223);
nand U6528 (N_6528,N_6297,N_6319);
nand U6529 (N_6529,N_6306,N_6394);
or U6530 (N_6530,N_6366,N_6358);
or U6531 (N_6531,N_6363,N_6303);
nand U6532 (N_6532,N_6230,N_6353);
nand U6533 (N_6533,N_6241,N_6385);
or U6534 (N_6534,N_6325,N_6306);
nand U6535 (N_6535,N_6285,N_6228);
nand U6536 (N_6536,N_6210,N_6314);
or U6537 (N_6537,N_6348,N_6388);
or U6538 (N_6538,N_6358,N_6213);
and U6539 (N_6539,N_6364,N_6301);
or U6540 (N_6540,N_6391,N_6361);
and U6541 (N_6541,N_6211,N_6286);
nand U6542 (N_6542,N_6313,N_6382);
nor U6543 (N_6543,N_6395,N_6309);
nor U6544 (N_6544,N_6202,N_6224);
nand U6545 (N_6545,N_6239,N_6353);
nor U6546 (N_6546,N_6276,N_6304);
nand U6547 (N_6547,N_6355,N_6367);
nor U6548 (N_6548,N_6316,N_6200);
nand U6549 (N_6549,N_6267,N_6253);
nand U6550 (N_6550,N_6358,N_6394);
nor U6551 (N_6551,N_6244,N_6220);
or U6552 (N_6552,N_6362,N_6216);
and U6553 (N_6553,N_6267,N_6227);
or U6554 (N_6554,N_6254,N_6283);
nor U6555 (N_6555,N_6296,N_6258);
nor U6556 (N_6556,N_6366,N_6288);
nor U6557 (N_6557,N_6383,N_6312);
or U6558 (N_6558,N_6216,N_6271);
nor U6559 (N_6559,N_6213,N_6345);
nor U6560 (N_6560,N_6260,N_6363);
nor U6561 (N_6561,N_6379,N_6361);
or U6562 (N_6562,N_6241,N_6226);
xnor U6563 (N_6563,N_6244,N_6213);
and U6564 (N_6564,N_6283,N_6318);
nand U6565 (N_6565,N_6219,N_6213);
nand U6566 (N_6566,N_6301,N_6240);
nand U6567 (N_6567,N_6360,N_6226);
nor U6568 (N_6568,N_6351,N_6279);
or U6569 (N_6569,N_6255,N_6312);
nand U6570 (N_6570,N_6382,N_6265);
nor U6571 (N_6571,N_6330,N_6274);
nor U6572 (N_6572,N_6298,N_6287);
nand U6573 (N_6573,N_6330,N_6310);
or U6574 (N_6574,N_6347,N_6254);
nand U6575 (N_6575,N_6318,N_6395);
nor U6576 (N_6576,N_6332,N_6231);
or U6577 (N_6577,N_6397,N_6290);
or U6578 (N_6578,N_6210,N_6329);
or U6579 (N_6579,N_6215,N_6350);
nor U6580 (N_6580,N_6300,N_6217);
nand U6581 (N_6581,N_6277,N_6256);
and U6582 (N_6582,N_6285,N_6245);
nand U6583 (N_6583,N_6354,N_6219);
nand U6584 (N_6584,N_6248,N_6292);
or U6585 (N_6585,N_6208,N_6391);
nand U6586 (N_6586,N_6341,N_6344);
nand U6587 (N_6587,N_6222,N_6347);
or U6588 (N_6588,N_6346,N_6344);
nand U6589 (N_6589,N_6301,N_6342);
and U6590 (N_6590,N_6213,N_6251);
or U6591 (N_6591,N_6231,N_6317);
nor U6592 (N_6592,N_6218,N_6336);
and U6593 (N_6593,N_6246,N_6339);
nor U6594 (N_6594,N_6386,N_6284);
nand U6595 (N_6595,N_6304,N_6391);
nand U6596 (N_6596,N_6202,N_6216);
nor U6597 (N_6597,N_6278,N_6385);
nand U6598 (N_6598,N_6282,N_6310);
nand U6599 (N_6599,N_6221,N_6335);
nor U6600 (N_6600,N_6488,N_6595);
and U6601 (N_6601,N_6556,N_6563);
nor U6602 (N_6602,N_6504,N_6494);
and U6603 (N_6603,N_6502,N_6468);
nand U6604 (N_6604,N_6485,N_6562);
nor U6605 (N_6605,N_6586,N_6406);
nand U6606 (N_6606,N_6497,N_6466);
and U6607 (N_6607,N_6549,N_6589);
nor U6608 (N_6608,N_6479,N_6525);
or U6609 (N_6609,N_6454,N_6545);
and U6610 (N_6610,N_6583,N_6420);
and U6611 (N_6611,N_6492,N_6418);
nand U6612 (N_6612,N_6574,N_6421);
or U6613 (N_6613,N_6408,N_6426);
or U6614 (N_6614,N_6489,N_6433);
and U6615 (N_6615,N_6431,N_6592);
xnor U6616 (N_6616,N_6453,N_6473);
and U6617 (N_6617,N_6417,N_6498);
and U6618 (N_6618,N_6540,N_6535);
and U6619 (N_6619,N_6512,N_6523);
or U6620 (N_6620,N_6532,N_6510);
nor U6621 (N_6621,N_6566,N_6461);
nand U6622 (N_6622,N_6518,N_6500);
nor U6623 (N_6623,N_6544,N_6425);
and U6624 (N_6624,N_6564,N_6531);
or U6625 (N_6625,N_6596,N_6437);
nor U6626 (N_6626,N_6438,N_6499);
nand U6627 (N_6627,N_6520,N_6591);
nor U6628 (N_6628,N_6590,N_6519);
and U6629 (N_6629,N_6597,N_6588);
nand U6630 (N_6630,N_6474,N_6599);
nor U6631 (N_6631,N_6422,N_6580);
and U6632 (N_6632,N_6475,N_6542);
nand U6633 (N_6633,N_6427,N_6491);
or U6634 (N_6634,N_6471,N_6515);
or U6635 (N_6635,N_6561,N_6430);
and U6636 (N_6636,N_6446,N_6546);
or U6637 (N_6637,N_6465,N_6441);
nand U6638 (N_6638,N_6521,N_6411);
nand U6639 (N_6639,N_6402,N_6528);
or U6640 (N_6640,N_6577,N_6505);
nor U6641 (N_6641,N_6413,N_6449);
or U6642 (N_6642,N_6559,N_6529);
and U6643 (N_6643,N_6587,N_6524);
or U6644 (N_6644,N_6442,N_6568);
or U6645 (N_6645,N_6536,N_6469);
nor U6646 (N_6646,N_6552,N_6533);
or U6647 (N_6647,N_6456,N_6572);
and U6648 (N_6648,N_6560,N_6578);
and U6649 (N_6649,N_6455,N_6506);
nor U6650 (N_6650,N_6548,N_6554);
nor U6651 (N_6651,N_6557,N_6571);
nand U6652 (N_6652,N_6565,N_6434);
or U6653 (N_6653,N_6405,N_6407);
or U6654 (N_6654,N_6403,N_6569);
nand U6655 (N_6655,N_6443,N_6470);
or U6656 (N_6656,N_6503,N_6447);
or U6657 (N_6657,N_6493,N_6436);
and U6658 (N_6658,N_6480,N_6401);
and U6659 (N_6659,N_6487,N_6584);
and U6660 (N_6660,N_6526,N_6541);
or U6661 (N_6661,N_6472,N_6409);
or U6662 (N_6662,N_6484,N_6508);
or U6663 (N_6663,N_6432,N_6483);
and U6664 (N_6664,N_6573,N_6452);
or U6665 (N_6665,N_6404,N_6478);
or U6666 (N_6666,N_6415,N_6598);
or U6667 (N_6667,N_6550,N_6464);
or U6668 (N_6668,N_6517,N_6576);
nand U6669 (N_6669,N_6440,N_6527);
and U6670 (N_6670,N_6410,N_6537);
or U6671 (N_6671,N_6495,N_6594);
and U6672 (N_6672,N_6593,N_6579);
and U6673 (N_6673,N_6585,N_6486);
and U6674 (N_6674,N_6513,N_6424);
nor U6675 (N_6675,N_6400,N_6511);
and U6676 (N_6676,N_6463,N_6582);
and U6677 (N_6677,N_6575,N_6496);
nand U6678 (N_6678,N_6539,N_6439);
or U6679 (N_6679,N_6460,N_6558);
and U6680 (N_6680,N_6428,N_6514);
or U6681 (N_6681,N_6522,N_6481);
or U6682 (N_6682,N_6412,N_6458);
nor U6683 (N_6683,N_6457,N_6435);
nor U6684 (N_6684,N_6451,N_6553);
and U6685 (N_6685,N_6462,N_6476);
nor U6686 (N_6686,N_6477,N_6467);
nand U6687 (N_6687,N_6534,N_6490);
nor U6688 (N_6688,N_6538,N_6423);
or U6689 (N_6689,N_6543,N_6501);
nor U6690 (N_6690,N_6507,N_6509);
nor U6691 (N_6691,N_6570,N_6448);
nor U6692 (N_6692,N_6530,N_6419);
nand U6693 (N_6693,N_6567,N_6414);
nand U6694 (N_6694,N_6445,N_6482);
and U6695 (N_6695,N_6450,N_6555);
or U6696 (N_6696,N_6416,N_6429);
nand U6697 (N_6697,N_6551,N_6516);
and U6698 (N_6698,N_6459,N_6444);
and U6699 (N_6699,N_6547,N_6581);
nand U6700 (N_6700,N_6472,N_6445);
nand U6701 (N_6701,N_6530,N_6444);
and U6702 (N_6702,N_6439,N_6411);
nor U6703 (N_6703,N_6472,N_6518);
or U6704 (N_6704,N_6459,N_6529);
or U6705 (N_6705,N_6492,N_6495);
or U6706 (N_6706,N_6519,N_6573);
nor U6707 (N_6707,N_6423,N_6567);
nand U6708 (N_6708,N_6403,N_6465);
or U6709 (N_6709,N_6434,N_6538);
or U6710 (N_6710,N_6583,N_6494);
and U6711 (N_6711,N_6483,N_6473);
and U6712 (N_6712,N_6435,N_6419);
or U6713 (N_6713,N_6448,N_6466);
or U6714 (N_6714,N_6506,N_6452);
or U6715 (N_6715,N_6420,N_6537);
nor U6716 (N_6716,N_6465,N_6461);
nand U6717 (N_6717,N_6550,N_6401);
nor U6718 (N_6718,N_6543,N_6589);
or U6719 (N_6719,N_6468,N_6429);
nor U6720 (N_6720,N_6594,N_6567);
and U6721 (N_6721,N_6413,N_6448);
nand U6722 (N_6722,N_6441,N_6545);
nor U6723 (N_6723,N_6521,N_6501);
or U6724 (N_6724,N_6405,N_6546);
nand U6725 (N_6725,N_6522,N_6447);
or U6726 (N_6726,N_6562,N_6526);
nor U6727 (N_6727,N_6581,N_6553);
or U6728 (N_6728,N_6583,N_6424);
nor U6729 (N_6729,N_6578,N_6458);
and U6730 (N_6730,N_6402,N_6465);
nand U6731 (N_6731,N_6540,N_6593);
nor U6732 (N_6732,N_6562,N_6575);
or U6733 (N_6733,N_6462,N_6580);
nand U6734 (N_6734,N_6480,N_6477);
and U6735 (N_6735,N_6533,N_6415);
or U6736 (N_6736,N_6416,N_6577);
or U6737 (N_6737,N_6512,N_6475);
nor U6738 (N_6738,N_6562,N_6594);
and U6739 (N_6739,N_6595,N_6568);
nor U6740 (N_6740,N_6596,N_6493);
nor U6741 (N_6741,N_6524,N_6503);
nor U6742 (N_6742,N_6587,N_6506);
nor U6743 (N_6743,N_6588,N_6493);
nand U6744 (N_6744,N_6537,N_6400);
nand U6745 (N_6745,N_6402,N_6538);
or U6746 (N_6746,N_6598,N_6518);
nand U6747 (N_6747,N_6547,N_6525);
and U6748 (N_6748,N_6474,N_6496);
or U6749 (N_6749,N_6499,N_6505);
nand U6750 (N_6750,N_6586,N_6428);
nand U6751 (N_6751,N_6422,N_6520);
and U6752 (N_6752,N_6539,N_6408);
nor U6753 (N_6753,N_6575,N_6476);
nor U6754 (N_6754,N_6442,N_6479);
nand U6755 (N_6755,N_6455,N_6452);
or U6756 (N_6756,N_6589,N_6567);
nor U6757 (N_6757,N_6473,N_6517);
or U6758 (N_6758,N_6593,N_6514);
nor U6759 (N_6759,N_6543,N_6427);
and U6760 (N_6760,N_6582,N_6541);
nor U6761 (N_6761,N_6443,N_6490);
nor U6762 (N_6762,N_6419,N_6404);
and U6763 (N_6763,N_6584,N_6400);
nor U6764 (N_6764,N_6564,N_6573);
and U6765 (N_6765,N_6517,N_6516);
nand U6766 (N_6766,N_6578,N_6404);
nand U6767 (N_6767,N_6456,N_6402);
nand U6768 (N_6768,N_6487,N_6588);
nor U6769 (N_6769,N_6547,N_6543);
nor U6770 (N_6770,N_6454,N_6533);
nand U6771 (N_6771,N_6553,N_6454);
or U6772 (N_6772,N_6412,N_6588);
and U6773 (N_6773,N_6473,N_6475);
and U6774 (N_6774,N_6487,N_6514);
nand U6775 (N_6775,N_6579,N_6434);
and U6776 (N_6776,N_6471,N_6438);
or U6777 (N_6777,N_6452,N_6582);
nor U6778 (N_6778,N_6527,N_6497);
nand U6779 (N_6779,N_6401,N_6440);
nor U6780 (N_6780,N_6488,N_6541);
or U6781 (N_6781,N_6548,N_6441);
nor U6782 (N_6782,N_6407,N_6416);
nor U6783 (N_6783,N_6447,N_6415);
nand U6784 (N_6784,N_6525,N_6403);
and U6785 (N_6785,N_6537,N_6593);
or U6786 (N_6786,N_6419,N_6484);
nor U6787 (N_6787,N_6558,N_6409);
and U6788 (N_6788,N_6599,N_6547);
or U6789 (N_6789,N_6464,N_6527);
nor U6790 (N_6790,N_6552,N_6572);
nor U6791 (N_6791,N_6585,N_6419);
and U6792 (N_6792,N_6451,N_6575);
xor U6793 (N_6793,N_6465,N_6562);
and U6794 (N_6794,N_6500,N_6449);
or U6795 (N_6795,N_6402,N_6454);
xnor U6796 (N_6796,N_6572,N_6517);
or U6797 (N_6797,N_6494,N_6557);
and U6798 (N_6798,N_6582,N_6465);
and U6799 (N_6799,N_6460,N_6476);
and U6800 (N_6800,N_6761,N_6747);
nand U6801 (N_6801,N_6710,N_6624);
nand U6802 (N_6802,N_6734,N_6793);
nor U6803 (N_6803,N_6713,N_6601);
nand U6804 (N_6804,N_6714,N_6704);
nand U6805 (N_6805,N_6623,N_6662);
or U6806 (N_6806,N_6667,N_6759);
nor U6807 (N_6807,N_6612,N_6751);
nand U6808 (N_6808,N_6649,N_6725);
and U6809 (N_6809,N_6782,N_6634);
nand U6810 (N_6810,N_6772,N_6702);
nor U6811 (N_6811,N_6669,N_6622);
nand U6812 (N_6812,N_6658,N_6693);
nand U6813 (N_6813,N_6722,N_6605);
nor U6814 (N_6814,N_6754,N_6645);
nand U6815 (N_6815,N_6686,N_6672);
and U6816 (N_6816,N_6684,N_6688);
and U6817 (N_6817,N_6746,N_6659);
and U6818 (N_6818,N_6703,N_6735);
and U6819 (N_6819,N_6680,N_6660);
nand U6820 (N_6820,N_6661,N_6687);
or U6821 (N_6821,N_6653,N_6603);
nor U6822 (N_6822,N_6628,N_6600);
and U6823 (N_6823,N_6699,N_6633);
nor U6824 (N_6824,N_6609,N_6642);
and U6825 (N_6825,N_6651,N_6666);
and U6826 (N_6826,N_6696,N_6729);
and U6827 (N_6827,N_6723,N_6654);
nor U6828 (N_6828,N_6656,N_6743);
nand U6829 (N_6829,N_6787,N_6630);
nand U6830 (N_6830,N_6671,N_6705);
nor U6831 (N_6831,N_6727,N_6640);
nand U6832 (N_6832,N_6773,N_6758);
or U6833 (N_6833,N_6790,N_6708);
nand U6834 (N_6834,N_6732,N_6785);
nor U6835 (N_6835,N_6730,N_6742);
xor U6836 (N_6836,N_6698,N_6607);
nand U6837 (N_6837,N_6768,N_6786);
nand U6838 (N_6838,N_6738,N_6736);
and U6839 (N_6839,N_6779,N_6744);
nand U6840 (N_6840,N_6748,N_6720);
and U6841 (N_6841,N_6652,N_6631);
nand U6842 (N_6842,N_6692,N_6755);
nor U6843 (N_6843,N_6778,N_6641);
or U6844 (N_6844,N_6724,N_6602);
and U6845 (N_6845,N_6739,N_6663);
nor U6846 (N_6846,N_6611,N_6769);
nand U6847 (N_6847,N_6616,N_6648);
or U6848 (N_6848,N_6719,N_6753);
nor U6849 (N_6849,N_6615,N_6789);
or U6850 (N_6850,N_6783,N_6689);
and U6851 (N_6851,N_6617,N_6749);
or U6852 (N_6852,N_6668,N_6670);
and U6853 (N_6853,N_6681,N_6695);
nor U6854 (N_6854,N_6780,N_6610);
and U6855 (N_6855,N_6756,N_6774);
nor U6856 (N_6856,N_6618,N_6608);
nor U6857 (N_6857,N_6614,N_6657);
nor U6858 (N_6858,N_6792,N_6781);
nand U6859 (N_6859,N_6635,N_6664);
or U6860 (N_6860,N_6752,N_6637);
nor U6861 (N_6861,N_6683,N_6665);
nand U6862 (N_6862,N_6626,N_6647);
nand U6863 (N_6863,N_6685,N_6726);
nand U6864 (N_6864,N_6798,N_6682);
nor U6865 (N_6865,N_6679,N_6766);
nor U6866 (N_6866,N_6740,N_6717);
nand U6867 (N_6867,N_6795,N_6697);
and U6868 (N_6868,N_6784,N_6643);
or U6869 (N_6869,N_6797,N_6604);
nand U6870 (N_6870,N_6655,N_6775);
or U6871 (N_6871,N_6788,N_6745);
nand U6872 (N_6872,N_6690,N_6777);
or U6873 (N_6873,N_6644,N_6776);
and U6874 (N_6874,N_6712,N_6613);
xor U6875 (N_6875,N_6731,N_6718);
and U6876 (N_6876,N_6706,N_6733);
or U6877 (N_6877,N_6636,N_6638);
or U6878 (N_6878,N_6757,N_6691);
or U6879 (N_6879,N_6621,N_6764);
and U6880 (N_6880,N_6762,N_6675);
and U6881 (N_6881,N_6673,N_6737);
and U6882 (N_6882,N_6767,N_6763);
or U6883 (N_6883,N_6701,N_6629);
xor U6884 (N_6884,N_6700,N_6650);
and U6885 (N_6885,N_6760,N_6728);
nor U6886 (N_6886,N_6709,N_6677);
and U6887 (N_6887,N_6771,N_6646);
nor U6888 (N_6888,N_6765,N_6715);
nor U6889 (N_6889,N_6639,N_6606);
or U6890 (N_6890,N_6627,N_6750);
and U6891 (N_6891,N_6770,N_6619);
nand U6892 (N_6892,N_6678,N_6796);
or U6893 (N_6893,N_6799,N_6716);
nor U6894 (N_6894,N_6791,N_6674);
nor U6895 (N_6895,N_6741,N_6794);
nor U6896 (N_6896,N_6711,N_6632);
nand U6897 (N_6897,N_6707,N_6694);
or U6898 (N_6898,N_6721,N_6676);
or U6899 (N_6899,N_6620,N_6625);
and U6900 (N_6900,N_6655,N_6657);
or U6901 (N_6901,N_6608,N_6622);
nand U6902 (N_6902,N_6775,N_6696);
or U6903 (N_6903,N_6604,N_6772);
or U6904 (N_6904,N_6622,N_6706);
and U6905 (N_6905,N_6693,N_6797);
nor U6906 (N_6906,N_6676,N_6735);
and U6907 (N_6907,N_6779,N_6714);
nand U6908 (N_6908,N_6638,N_6610);
or U6909 (N_6909,N_6667,N_6625);
and U6910 (N_6910,N_6701,N_6783);
or U6911 (N_6911,N_6642,N_6691);
nor U6912 (N_6912,N_6663,N_6638);
or U6913 (N_6913,N_6772,N_6603);
and U6914 (N_6914,N_6664,N_6742);
and U6915 (N_6915,N_6794,N_6654);
and U6916 (N_6916,N_6757,N_6679);
nand U6917 (N_6917,N_6678,N_6778);
nand U6918 (N_6918,N_6635,N_6678);
nor U6919 (N_6919,N_6653,N_6761);
nor U6920 (N_6920,N_6708,N_6653);
and U6921 (N_6921,N_6748,N_6681);
and U6922 (N_6922,N_6657,N_6778);
nand U6923 (N_6923,N_6649,N_6601);
or U6924 (N_6924,N_6601,N_6719);
nor U6925 (N_6925,N_6664,N_6795);
or U6926 (N_6926,N_6722,N_6762);
and U6927 (N_6927,N_6783,N_6798);
or U6928 (N_6928,N_6761,N_6621);
and U6929 (N_6929,N_6688,N_6771);
nor U6930 (N_6930,N_6759,N_6763);
nor U6931 (N_6931,N_6618,N_6604);
or U6932 (N_6932,N_6775,N_6609);
or U6933 (N_6933,N_6602,N_6676);
nand U6934 (N_6934,N_6637,N_6677);
and U6935 (N_6935,N_6604,N_6605);
nor U6936 (N_6936,N_6772,N_6755);
or U6937 (N_6937,N_6729,N_6649);
nand U6938 (N_6938,N_6767,N_6778);
or U6939 (N_6939,N_6696,N_6715);
nand U6940 (N_6940,N_6611,N_6716);
nor U6941 (N_6941,N_6706,N_6630);
nand U6942 (N_6942,N_6699,N_6791);
and U6943 (N_6943,N_6761,N_6667);
or U6944 (N_6944,N_6723,N_6694);
nor U6945 (N_6945,N_6693,N_6629);
and U6946 (N_6946,N_6699,N_6603);
or U6947 (N_6947,N_6784,N_6704);
or U6948 (N_6948,N_6727,N_6753);
nand U6949 (N_6949,N_6764,N_6669);
nor U6950 (N_6950,N_6758,N_6652);
or U6951 (N_6951,N_6688,N_6661);
nor U6952 (N_6952,N_6720,N_6751);
nand U6953 (N_6953,N_6795,N_6634);
and U6954 (N_6954,N_6693,N_6679);
nand U6955 (N_6955,N_6622,N_6606);
and U6956 (N_6956,N_6773,N_6747);
or U6957 (N_6957,N_6721,N_6613);
nor U6958 (N_6958,N_6612,N_6607);
nand U6959 (N_6959,N_6641,N_6789);
or U6960 (N_6960,N_6684,N_6632);
nand U6961 (N_6961,N_6684,N_6704);
or U6962 (N_6962,N_6781,N_6719);
nor U6963 (N_6963,N_6738,N_6714);
or U6964 (N_6964,N_6708,N_6656);
and U6965 (N_6965,N_6610,N_6611);
nor U6966 (N_6966,N_6761,N_6640);
and U6967 (N_6967,N_6612,N_6621);
or U6968 (N_6968,N_6671,N_6641);
nor U6969 (N_6969,N_6785,N_6743);
and U6970 (N_6970,N_6680,N_6693);
nor U6971 (N_6971,N_6775,N_6657);
and U6972 (N_6972,N_6734,N_6786);
nand U6973 (N_6973,N_6721,N_6620);
nand U6974 (N_6974,N_6692,N_6642);
nand U6975 (N_6975,N_6696,N_6654);
or U6976 (N_6976,N_6653,N_6660);
nor U6977 (N_6977,N_6761,N_6704);
nand U6978 (N_6978,N_6711,N_6616);
nand U6979 (N_6979,N_6624,N_6794);
nor U6980 (N_6980,N_6681,N_6797);
nand U6981 (N_6981,N_6626,N_6762);
nor U6982 (N_6982,N_6713,N_6603);
or U6983 (N_6983,N_6756,N_6670);
nor U6984 (N_6984,N_6623,N_6637);
and U6985 (N_6985,N_6752,N_6672);
and U6986 (N_6986,N_6651,N_6739);
nor U6987 (N_6987,N_6719,N_6700);
nor U6988 (N_6988,N_6628,N_6607);
or U6989 (N_6989,N_6695,N_6721);
and U6990 (N_6990,N_6715,N_6759);
and U6991 (N_6991,N_6727,N_6674);
nor U6992 (N_6992,N_6770,N_6673);
nor U6993 (N_6993,N_6792,N_6780);
and U6994 (N_6994,N_6674,N_6787);
and U6995 (N_6995,N_6708,N_6762);
or U6996 (N_6996,N_6659,N_6794);
and U6997 (N_6997,N_6713,N_6771);
or U6998 (N_6998,N_6753,N_6667);
and U6999 (N_6999,N_6615,N_6653);
and U7000 (N_7000,N_6906,N_6960);
and U7001 (N_7001,N_6934,N_6956);
nor U7002 (N_7002,N_6899,N_6829);
or U7003 (N_7003,N_6913,N_6871);
nand U7004 (N_7004,N_6907,N_6955);
or U7005 (N_7005,N_6833,N_6809);
nor U7006 (N_7006,N_6982,N_6888);
nand U7007 (N_7007,N_6842,N_6971);
nand U7008 (N_7008,N_6917,N_6890);
and U7009 (N_7009,N_6848,N_6900);
nor U7010 (N_7010,N_6841,N_6922);
nor U7011 (N_7011,N_6948,N_6814);
nor U7012 (N_7012,N_6976,N_6817);
nor U7013 (N_7013,N_6927,N_6930);
or U7014 (N_7014,N_6962,N_6891);
nor U7015 (N_7015,N_6920,N_6808);
nor U7016 (N_7016,N_6911,N_6884);
and U7017 (N_7017,N_6897,N_6925);
and U7018 (N_7018,N_6981,N_6855);
nor U7019 (N_7019,N_6880,N_6802);
or U7020 (N_7020,N_6827,N_6926);
and U7021 (N_7021,N_6861,N_6912);
nor U7022 (N_7022,N_6994,N_6983);
or U7023 (N_7023,N_6835,N_6815);
nand U7024 (N_7024,N_6810,N_6873);
nor U7025 (N_7025,N_6980,N_6850);
and U7026 (N_7026,N_6995,N_6967);
or U7027 (N_7027,N_6964,N_6919);
and U7028 (N_7028,N_6915,N_6844);
nor U7029 (N_7029,N_6941,N_6921);
and U7030 (N_7030,N_6826,N_6818);
nand U7031 (N_7031,N_6977,N_6837);
or U7032 (N_7032,N_6940,N_6851);
and U7033 (N_7033,N_6916,N_6867);
nand U7034 (N_7034,N_6840,N_6988);
and U7035 (N_7035,N_6979,N_6951);
nor U7036 (N_7036,N_6975,N_6885);
nand U7037 (N_7037,N_6957,N_6847);
nand U7038 (N_7038,N_6811,N_6932);
nand U7039 (N_7039,N_6801,N_6965);
or U7040 (N_7040,N_6918,N_6836);
or U7041 (N_7041,N_6992,N_6883);
and U7042 (N_7042,N_6999,N_6806);
nor U7043 (N_7043,N_6984,N_6901);
and U7044 (N_7044,N_6966,N_6838);
or U7045 (N_7045,N_6902,N_6931);
and U7046 (N_7046,N_6893,N_6824);
nand U7047 (N_7047,N_6936,N_6896);
nand U7048 (N_7048,N_6822,N_6996);
and U7049 (N_7049,N_6989,N_6942);
or U7050 (N_7050,N_6895,N_6990);
or U7051 (N_7051,N_6875,N_6991);
and U7052 (N_7052,N_6857,N_6892);
and U7053 (N_7053,N_6929,N_6886);
and U7054 (N_7054,N_6914,N_6972);
or U7055 (N_7055,N_6856,N_6908);
or U7056 (N_7056,N_6963,N_6974);
nand U7057 (N_7057,N_6993,N_6862);
nand U7058 (N_7058,N_6820,N_6816);
nor U7059 (N_7059,N_6952,N_6866);
nand U7060 (N_7060,N_6909,N_6953);
nand U7061 (N_7061,N_6878,N_6830);
or U7062 (N_7062,N_6938,N_6954);
nor U7063 (N_7063,N_6870,N_6877);
nor U7064 (N_7064,N_6823,N_6803);
or U7065 (N_7065,N_6998,N_6959);
or U7066 (N_7066,N_6946,N_6874);
and U7067 (N_7067,N_6939,N_6968);
and U7068 (N_7068,N_6872,N_6904);
nand U7069 (N_7069,N_6813,N_6839);
and U7070 (N_7070,N_6947,N_6882);
nor U7071 (N_7071,N_6804,N_6935);
or U7072 (N_7072,N_6910,N_6961);
and U7073 (N_7073,N_6843,N_6978);
nand U7074 (N_7074,N_6854,N_6944);
nor U7075 (N_7075,N_6969,N_6831);
or U7076 (N_7076,N_6898,N_6986);
nand U7077 (N_7077,N_6943,N_6849);
and U7078 (N_7078,N_6846,N_6865);
nor U7079 (N_7079,N_6869,N_6800);
nand U7080 (N_7080,N_6923,N_6807);
or U7081 (N_7081,N_6845,N_6973);
nand U7082 (N_7082,N_6859,N_6834);
nor U7083 (N_7083,N_6903,N_6832);
nand U7084 (N_7084,N_6949,N_6987);
and U7085 (N_7085,N_6933,N_6864);
or U7086 (N_7086,N_6805,N_6858);
nor U7087 (N_7087,N_6876,N_6985);
xor U7088 (N_7088,N_6828,N_6881);
nand U7089 (N_7089,N_6970,N_6889);
and U7090 (N_7090,N_6819,N_6825);
or U7091 (N_7091,N_6937,N_6821);
nand U7092 (N_7092,N_6945,N_6997);
nor U7093 (N_7093,N_6868,N_6879);
nor U7094 (N_7094,N_6905,N_6958);
nor U7095 (N_7095,N_6894,N_6887);
nor U7096 (N_7096,N_6853,N_6863);
nor U7097 (N_7097,N_6924,N_6812);
or U7098 (N_7098,N_6928,N_6860);
or U7099 (N_7099,N_6852,N_6950);
or U7100 (N_7100,N_6915,N_6966);
or U7101 (N_7101,N_6800,N_6890);
nand U7102 (N_7102,N_6845,N_6898);
or U7103 (N_7103,N_6820,N_6885);
nand U7104 (N_7104,N_6869,N_6843);
or U7105 (N_7105,N_6828,N_6835);
nor U7106 (N_7106,N_6844,N_6804);
or U7107 (N_7107,N_6979,N_6949);
nand U7108 (N_7108,N_6955,N_6888);
nand U7109 (N_7109,N_6819,N_6915);
nand U7110 (N_7110,N_6808,N_6845);
nor U7111 (N_7111,N_6899,N_6919);
nand U7112 (N_7112,N_6890,N_6871);
nand U7113 (N_7113,N_6872,N_6888);
nand U7114 (N_7114,N_6944,N_6924);
and U7115 (N_7115,N_6977,N_6910);
nand U7116 (N_7116,N_6956,N_6985);
or U7117 (N_7117,N_6823,N_6938);
nor U7118 (N_7118,N_6896,N_6995);
nor U7119 (N_7119,N_6955,N_6995);
and U7120 (N_7120,N_6808,N_6858);
and U7121 (N_7121,N_6916,N_6802);
or U7122 (N_7122,N_6950,N_6873);
and U7123 (N_7123,N_6998,N_6933);
and U7124 (N_7124,N_6803,N_6923);
nand U7125 (N_7125,N_6901,N_6992);
and U7126 (N_7126,N_6969,N_6966);
or U7127 (N_7127,N_6969,N_6930);
nor U7128 (N_7128,N_6825,N_6954);
nor U7129 (N_7129,N_6912,N_6817);
xor U7130 (N_7130,N_6926,N_6824);
nand U7131 (N_7131,N_6923,N_6924);
or U7132 (N_7132,N_6844,N_6977);
or U7133 (N_7133,N_6835,N_6810);
and U7134 (N_7134,N_6955,N_6871);
nand U7135 (N_7135,N_6800,N_6857);
or U7136 (N_7136,N_6967,N_6969);
nor U7137 (N_7137,N_6913,N_6916);
nor U7138 (N_7138,N_6847,N_6850);
nand U7139 (N_7139,N_6938,N_6877);
nor U7140 (N_7140,N_6928,N_6849);
xor U7141 (N_7141,N_6860,N_6847);
or U7142 (N_7142,N_6924,N_6920);
nor U7143 (N_7143,N_6852,N_6954);
or U7144 (N_7144,N_6933,N_6912);
nand U7145 (N_7145,N_6800,N_6974);
nand U7146 (N_7146,N_6912,N_6858);
or U7147 (N_7147,N_6906,N_6821);
or U7148 (N_7148,N_6955,N_6862);
and U7149 (N_7149,N_6927,N_6919);
or U7150 (N_7150,N_6859,N_6818);
and U7151 (N_7151,N_6995,N_6804);
nor U7152 (N_7152,N_6987,N_6945);
nor U7153 (N_7153,N_6828,N_6962);
xnor U7154 (N_7154,N_6887,N_6837);
nor U7155 (N_7155,N_6953,N_6971);
nor U7156 (N_7156,N_6866,N_6805);
nor U7157 (N_7157,N_6896,N_6898);
nor U7158 (N_7158,N_6803,N_6810);
and U7159 (N_7159,N_6900,N_6879);
nor U7160 (N_7160,N_6807,N_6805);
nor U7161 (N_7161,N_6907,N_6951);
nand U7162 (N_7162,N_6871,N_6954);
and U7163 (N_7163,N_6866,N_6984);
or U7164 (N_7164,N_6978,N_6891);
nand U7165 (N_7165,N_6971,N_6950);
nor U7166 (N_7166,N_6802,N_6981);
nand U7167 (N_7167,N_6814,N_6842);
and U7168 (N_7168,N_6972,N_6918);
nand U7169 (N_7169,N_6809,N_6997);
nor U7170 (N_7170,N_6960,N_6925);
nor U7171 (N_7171,N_6995,N_6867);
nand U7172 (N_7172,N_6896,N_6859);
or U7173 (N_7173,N_6830,N_6901);
or U7174 (N_7174,N_6946,N_6880);
nor U7175 (N_7175,N_6964,N_6877);
nand U7176 (N_7176,N_6892,N_6883);
or U7177 (N_7177,N_6835,N_6834);
nand U7178 (N_7178,N_6842,N_6908);
or U7179 (N_7179,N_6880,N_6950);
or U7180 (N_7180,N_6871,N_6881);
and U7181 (N_7181,N_6833,N_6931);
nand U7182 (N_7182,N_6801,N_6907);
nand U7183 (N_7183,N_6922,N_6879);
and U7184 (N_7184,N_6845,N_6944);
and U7185 (N_7185,N_6980,N_6872);
or U7186 (N_7186,N_6818,N_6825);
nand U7187 (N_7187,N_6802,N_6922);
and U7188 (N_7188,N_6807,N_6995);
and U7189 (N_7189,N_6842,N_6898);
or U7190 (N_7190,N_6853,N_6977);
or U7191 (N_7191,N_6921,N_6875);
nor U7192 (N_7192,N_6995,N_6991);
and U7193 (N_7193,N_6847,N_6982);
nor U7194 (N_7194,N_6895,N_6880);
nand U7195 (N_7195,N_6889,N_6954);
nand U7196 (N_7196,N_6813,N_6876);
or U7197 (N_7197,N_6881,N_6945);
nor U7198 (N_7198,N_6973,N_6994);
or U7199 (N_7199,N_6993,N_6982);
or U7200 (N_7200,N_7031,N_7113);
or U7201 (N_7201,N_7103,N_7096);
nand U7202 (N_7202,N_7115,N_7048);
nand U7203 (N_7203,N_7030,N_7035);
and U7204 (N_7204,N_7047,N_7154);
or U7205 (N_7205,N_7078,N_7184);
nor U7206 (N_7206,N_7053,N_7063);
or U7207 (N_7207,N_7094,N_7043);
and U7208 (N_7208,N_7017,N_7083);
and U7209 (N_7209,N_7138,N_7098);
or U7210 (N_7210,N_7158,N_7197);
nor U7211 (N_7211,N_7165,N_7022);
and U7212 (N_7212,N_7146,N_7037);
or U7213 (N_7213,N_7012,N_7044);
nand U7214 (N_7214,N_7157,N_7075);
and U7215 (N_7215,N_7172,N_7149);
nor U7216 (N_7216,N_7198,N_7010);
nand U7217 (N_7217,N_7191,N_7056);
nor U7218 (N_7218,N_7170,N_7135);
or U7219 (N_7219,N_7190,N_7189);
nand U7220 (N_7220,N_7153,N_7059);
or U7221 (N_7221,N_7093,N_7061);
nor U7222 (N_7222,N_7106,N_7007);
xor U7223 (N_7223,N_7069,N_7133);
or U7224 (N_7224,N_7193,N_7101);
and U7225 (N_7225,N_7100,N_7084);
nand U7226 (N_7226,N_7001,N_7112);
nor U7227 (N_7227,N_7156,N_7058);
and U7228 (N_7228,N_7178,N_7004);
and U7229 (N_7229,N_7182,N_7041);
and U7230 (N_7230,N_7039,N_7130);
or U7231 (N_7231,N_7161,N_7033);
nor U7232 (N_7232,N_7076,N_7159);
or U7233 (N_7233,N_7183,N_7023);
nand U7234 (N_7234,N_7181,N_7049);
and U7235 (N_7235,N_7095,N_7167);
nand U7236 (N_7236,N_7051,N_7176);
nand U7237 (N_7237,N_7088,N_7145);
or U7238 (N_7238,N_7060,N_7029);
nor U7239 (N_7239,N_7124,N_7092);
nor U7240 (N_7240,N_7068,N_7097);
nor U7241 (N_7241,N_7090,N_7117);
nor U7242 (N_7242,N_7186,N_7034);
and U7243 (N_7243,N_7091,N_7136);
xnor U7244 (N_7244,N_7114,N_7195);
and U7245 (N_7245,N_7099,N_7109);
nor U7246 (N_7246,N_7110,N_7026);
or U7247 (N_7247,N_7028,N_7074);
nor U7248 (N_7248,N_7143,N_7024);
or U7249 (N_7249,N_7127,N_7042);
and U7250 (N_7250,N_7105,N_7150);
or U7251 (N_7251,N_7122,N_7192);
or U7252 (N_7252,N_7177,N_7046);
nand U7253 (N_7253,N_7005,N_7123);
and U7254 (N_7254,N_7164,N_7000);
and U7255 (N_7255,N_7072,N_7008);
or U7256 (N_7256,N_7139,N_7196);
and U7257 (N_7257,N_7065,N_7020);
or U7258 (N_7258,N_7032,N_7108);
or U7259 (N_7259,N_7129,N_7018);
nand U7260 (N_7260,N_7073,N_7116);
nand U7261 (N_7261,N_7188,N_7055);
and U7262 (N_7262,N_7070,N_7134);
or U7263 (N_7263,N_7045,N_7187);
or U7264 (N_7264,N_7057,N_7185);
nor U7265 (N_7265,N_7111,N_7118);
nand U7266 (N_7266,N_7141,N_7140);
and U7267 (N_7267,N_7040,N_7163);
and U7268 (N_7268,N_7168,N_7171);
and U7269 (N_7269,N_7194,N_7086);
and U7270 (N_7270,N_7152,N_7160);
nand U7271 (N_7271,N_7011,N_7064);
nor U7272 (N_7272,N_7137,N_7013);
nand U7273 (N_7273,N_7104,N_7066);
and U7274 (N_7274,N_7175,N_7085);
and U7275 (N_7275,N_7006,N_7071);
or U7276 (N_7276,N_7180,N_7148);
and U7277 (N_7277,N_7079,N_7125);
nand U7278 (N_7278,N_7082,N_7128);
nand U7279 (N_7279,N_7132,N_7036);
nor U7280 (N_7280,N_7166,N_7102);
nor U7281 (N_7281,N_7162,N_7151);
or U7282 (N_7282,N_7016,N_7009);
nand U7283 (N_7283,N_7173,N_7174);
or U7284 (N_7284,N_7107,N_7003);
nand U7285 (N_7285,N_7054,N_7019);
or U7286 (N_7286,N_7080,N_7131);
or U7287 (N_7287,N_7050,N_7002);
or U7288 (N_7288,N_7199,N_7144);
nand U7289 (N_7289,N_7120,N_7038);
or U7290 (N_7290,N_7081,N_7121);
nand U7291 (N_7291,N_7014,N_7142);
or U7292 (N_7292,N_7077,N_7052);
nand U7293 (N_7293,N_7025,N_7021);
nor U7294 (N_7294,N_7067,N_7169);
nand U7295 (N_7295,N_7147,N_7179);
and U7296 (N_7296,N_7119,N_7089);
nor U7297 (N_7297,N_7015,N_7087);
nor U7298 (N_7298,N_7155,N_7126);
and U7299 (N_7299,N_7027,N_7062);
or U7300 (N_7300,N_7048,N_7074);
xor U7301 (N_7301,N_7168,N_7135);
or U7302 (N_7302,N_7162,N_7118);
and U7303 (N_7303,N_7054,N_7117);
nand U7304 (N_7304,N_7003,N_7169);
nor U7305 (N_7305,N_7165,N_7070);
nor U7306 (N_7306,N_7088,N_7110);
or U7307 (N_7307,N_7192,N_7006);
or U7308 (N_7308,N_7081,N_7163);
nand U7309 (N_7309,N_7082,N_7074);
or U7310 (N_7310,N_7109,N_7152);
nor U7311 (N_7311,N_7065,N_7043);
nor U7312 (N_7312,N_7055,N_7074);
nor U7313 (N_7313,N_7158,N_7024);
xnor U7314 (N_7314,N_7020,N_7086);
nand U7315 (N_7315,N_7161,N_7002);
or U7316 (N_7316,N_7089,N_7166);
nor U7317 (N_7317,N_7050,N_7145);
or U7318 (N_7318,N_7126,N_7069);
nand U7319 (N_7319,N_7174,N_7008);
and U7320 (N_7320,N_7046,N_7034);
nand U7321 (N_7321,N_7007,N_7027);
and U7322 (N_7322,N_7169,N_7113);
or U7323 (N_7323,N_7076,N_7192);
nand U7324 (N_7324,N_7083,N_7109);
nand U7325 (N_7325,N_7075,N_7101);
nor U7326 (N_7326,N_7079,N_7118);
or U7327 (N_7327,N_7035,N_7089);
or U7328 (N_7328,N_7121,N_7119);
or U7329 (N_7329,N_7157,N_7060);
and U7330 (N_7330,N_7096,N_7023);
nor U7331 (N_7331,N_7164,N_7079);
nor U7332 (N_7332,N_7192,N_7009);
nor U7333 (N_7333,N_7048,N_7184);
and U7334 (N_7334,N_7067,N_7120);
or U7335 (N_7335,N_7096,N_7031);
or U7336 (N_7336,N_7182,N_7113);
or U7337 (N_7337,N_7035,N_7053);
nand U7338 (N_7338,N_7088,N_7150);
nand U7339 (N_7339,N_7062,N_7025);
and U7340 (N_7340,N_7025,N_7099);
nor U7341 (N_7341,N_7121,N_7183);
and U7342 (N_7342,N_7003,N_7097);
or U7343 (N_7343,N_7043,N_7078);
nand U7344 (N_7344,N_7083,N_7041);
nand U7345 (N_7345,N_7040,N_7008);
nor U7346 (N_7346,N_7160,N_7016);
nand U7347 (N_7347,N_7109,N_7051);
nand U7348 (N_7348,N_7199,N_7109);
and U7349 (N_7349,N_7073,N_7133);
nor U7350 (N_7350,N_7038,N_7177);
or U7351 (N_7351,N_7148,N_7109);
or U7352 (N_7352,N_7051,N_7153);
nor U7353 (N_7353,N_7021,N_7057);
and U7354 (N_7354,N_7063,N_7059);
xnor U7355 (N_7355,N_7126,N_7107);
or U7356 (N_7356,N_7010,N_7011);
or U7357 (N_7357,N_7195,N_7026);
and U7358 (N_7358,N_7157,N_7130);
or U7359 (N_7359,N_7122,N_7027);
or U7360 (N_7360,N_7053,N_7185);
nor U7361 (N_7361,N_7139,N_7095);
nand U7362 (N_7362,N_7010,N_7051);
and U7363 (N_7363,N_7097,N_7038);
and U7364 (N_7364,N_7174,N_7134);
or U7365 (N_7365,N_7156,N_7123);
or U7366 (N_7366,N_7100,N_7187);
nand U7367 (N_7367,N_7008,N_7010);
nor U7368 (N_7368,N_7053,N_7092);
or U7369 (N_7369,N_7155,N_7051);
or U7370 (N_7370,N_7145,N_7128);
or U7371 (N_7371,N_7148,N_7084);
and U7372 (N_7372,N_7074,N_7161);
nand U7373 (N_7373,N_7035,N_7109);
nor U7374 (N_7374,N_7123,N_7031);
and U7375 (N_7375,N_7085,N_7026);
or U7376 (N_7376,N_7025,N_7010);
or U7377 (N_7377,N_7039,N_7045);
nand U7378 (N_7378,N_7183,N_7131);
and U7379 (N_7379,N_7061,N_7014);
or U7380 (N_7380,N_7044,N_7181);
or U7381 (N_7381,N_7169,N_7180);
nor U7382 (N_7382,N_7157,N_7191);
xor U7383 (N_7383,N_7182,N_7111);
nand U7384 (N_7384,N_7046,N_7196);
nand U7385 (N_7385,N_7146,N_7158);
or U7386 (N_7386,N_7194,N_7166);
nand U7387 (N_7387,N_7106,N_7034);
nor U7388 (N_7388,N_7073,N_7022);
or U7389 (N_7389,N_7008,N_7058);
and U7390 (N_7390,N_7147,N_7031);
nand U7391 (N_7391,N_7190,N_7092);
nor U7392 (N_7392,N_7112,N_7065);
and U7393 (N_7393,N_7042,N_7048);
or U7394 (N_7394,N_7142,N_7105);
and U7395 (N_7395,N_7071,N_7166);
or U7396 (N_7396,N_7126,N_7184);
or U7397 (N_7397,N_7117,N_7071);
or U7398 (N_7398,N_7087,N_7061);
nand U7399 (N_7399,N_7025,N_7170);
nor U7400 (N_7400,N_7344,N_7250);
nor U7401 (N_7401,N_7395,N_7249);
nand U7402 (N_7402,N_7383,N_7259);
nand U7403 (N_7403,N_7293,N_7372);
and U7404 (N_7404,N_7260,N_7346);
or U7405 (N_7405,N_7313,N_7345);
nor U7406 (N_7406,N_7377,N_7357);
or U7407 (N_7407,N_7333,N_7360);
nand U7408 (N_7408,N_7353,N_7285);
or U7409 (N_7409,N_7298,N_7247);
nand U7410 (N_7410,N_7299,N_7233);
or U7411 (N_7411,N_7314,N_7244);
nor U7412 (N_7412,N_7365,N_7374);
and U7413 (N_7413,N_7327,N_7253);
and U7414 (N_7414,N_7217,N_7339);
nor U7415 (N_7415,N_7282,N_7231);
or U7416 (N_7416,N_7286,N_7207);
and U7417 (N_7417,N_7397,N_7255);
and U7418 (N_7418,N_7200,N_7274);
nor U7419 (N_7419,N_7238,N_7328);
and U7420 (N_7420,N_7213,N_7246);
and U7421 (N_7421,N_7348,N_7373);
or U7422 (N_7422,N_7394,N_7292);
and U7423 (N_7423,N_7214,N_7354);
nand U7424 (N_7424,N_7218,N_7316);
and U7425 (N_7425,N_7295,N_7368);
or U7426 (N_7426,N_7257,N_7245);
and U7427 (N_7427,N_7399,N_7370);
or U7428 (N_7428,N_7202,N_7273);
or U7429 (N_7429,N_7223,N_7270);
nand U7430 (N_7430,N_7387,N_7204);
nor U7431 (N_7431,N_7227,N_7385);
nor U7432 (N_7432,N_7330,N_7389);
nand U7433 (N_7433,N_7358,N_7258);
or U7434 (N_7434,N_7284,N_7243);
nor U7435 (N_7435,N_7278,N_7288);
nor U7436 (N_7436,N_7239,N_7291);
or U7437 (N_7437,N_7275,N_7268);
nor U7438 (N_7438,N_7281,N_7396);
nand U7439 (N_7439,N_7392,N_7210);
nand U7440 (N_7440,N_7359,N_7341);
or U7441 (N_7441,N_7376,N_7312);
or U7442 (N_7442,N_7232,N_7332);
and U7443 (N_7443,N_7271,N_7325);
nor U7444 (N_7444,N_7221,N_7201);
and U7445 (N_7445,N_7315,N_7300);
nor U7446 (N_7446,N_7351,N_7267);
nand U7447 (N_7447,N_7265,N_7350);
or U7448 (N_7448,N_7296,N_7248);
nor U7449 (N_7449,N_7352,N_7229);
nand U7450 (N_7450,N_7256,N_7317);
or U7451 (N_7451,N_7215,N_7382);
or U7452 (N_7452,N_7277,N_7356);
xor U7453 (N_7453,N_7326,N_7391);
and U7454 (N_7454,N_7363,N_7225);
and U7455 (N_7455,N_7371,N_7216);
or U7456 (N_7456,N_7219,N_7224);
or U7457 (N_7457,N_7289,N_7254);
nand U7458 (N_7458,N_7355,N_7369);
nand U7459 (N_7459,N_7307,N_7336);
and U7460 (N_7460,N_7302,N_7261);
nor U7461 (N_7461,N_7308,N_7220);
or U7462 (N_7462,N_7390,N_7319);
nand U7463 (N_7463,N_7375,N_7340);
nor U7464 (N_7464,N_7335,N_7251);
nand U7465 (N_7465,N_7342,N_7311);
nand U7466 (N_7466,N_7309,N_7209);
nand U7467 (N_7467,N_7303,N_7310);
and U7468 (N_7468,N_7320,N_7280);
and U7469 (N_7469,N_7305,N_7306);
nor U7470 (N_7470,N_7321,N_7331);
nand U7471 (N_7471,N_7235,N_7240);
nand U7472 (N_7472,N_7337,N_7301);
nand U7473 (N_7473,N_7241,N_7228);
nor U7474 (N_7474,N_7329,N_7206);
and U7475 (N_7475,N_7347,N_7324);
and U7476 (N_7476,N_7242,N_7290);
nor U7477 (N_7477,N_7367,N_7236);
nor U7478 (N_7478,N_7361,N_7283);
or U7479 (N_7479,N_7266,N_7205);
nor U7480 (N_7480,N_7222,N_7323);
nor U7481 (N_7481,N_7203,N_7338);
and U7482 (N_7482,N_7264,N_7208);
nor U7483 (N_7483,N_7234,N_7380);
nor U7484 (N_7484,N_7262,N_7386);
nand U7485 (N_7485,N_7226,N_7322);
and U7486 (N_7486,N_7212,N_7378);
and U7487 (N_7487,N_7381,N_7279);
nor U7488 (N_7488,N_7318,N_7388);
or U7489 (N_7489,N_7276,N_7269);
nand U7490 (N_7490,N_7272,N_7230);
nand U7491 (N_7491,N_7349,N_7304);
nand U7492 (N_7492,N_7364,N_7393);
nor U7493 (N_7493,N_7297,N_7287);
and U7494 (N_7494,N_7343,N_7294);
and U7495 (N_7495,N_7362,N_7398);
or U7496 (N_7496,N_7379,N_7334);
or U7497 (N_7497,N_7384,N_7366);
and U7498 (N_7498,N_7237,N_7263);
nor U7499 (N_7499,N_7211,N_7252);
or U7500 (N_7500,N_7284,N_7210);
or U7501 (N_7501,N_7204,N_7305);
and U7502 (N_7502,N_7239,N_7218);
nor U7503 (N_7503,N_7270,N_7304);
and U7504 (N_7504,N_7278,N_7391);
nor U7505 (N_7505,N_7200,N_7367);
and U7506 (N_7506,N_7234,N_7392);
or U7507 (N_7507,N_7356,N_7366);
or U7508 (N_7508,N_7300,N_7297);
and U7509 (N_7509,N_7313,N_7217);
or U7510 (N_7510,N_7295,N_7276);
xor U7511 (N_7511,N_7271,N_7221);
or U7512 (N_7512,N_7334,N_7268);
nand U7513 (N_7513,N_7344,N_7258);
nand U7514 (N_7514,N_7321,N_7260);
nand U7515 (N_7515,N_7342,N_7291);
and U7516 (N_7516,N_7359,N_7248);
and U7517 (N_7517,N_7319,N_7204);
and U7518 (N_7518,N_7346,N_7357);
and U7519 (N_7519,N_7268,N_7211);
or U7520 (N_7520,N_7213,N_7265);
and U7521 (N_7521,N_7366,N_7320);
nand U7522 (N_7522,N_7357,N_7328);
and U7523 (N_7523,N_7332,N_7206);
nor U7524 (N_7524,N_7218,N_7279);
or U7525 (N_7525,N_7222,N_7295);
or U7526 (N_7526,N_7252,N_7277);
nand U7527 (N_7527,N_7298,N_7209);
and U7528 (N_7528,N_7319,N_7265);
and U7529 (N_7529,N_7386,N_7345);
nand U7530 (N_7530,N_7243,N_7244);
nand U7531 (N_7531,N_7353,N_7328);
and U7532 (N_7532,N_7275,N_7265);
or U7533 (N_7533,N_7208,N_7226);
and U7534 (N_7534,N_7335,N_7283);
or U7535 (N_7535,N_7273,N_7256);
nand U7536 (N_7536,N_7389,N_7242);
and U7537 (N_7537,N_7273,N_7272);
nor U7538 (N_7538,N_7345,N_7285);
or U7539 (N_7539,N_7395,N_7362);
nor U7540 (N_7540,N_7321,N_7268);
nand U7541 (N_7541,N_7328,N_7230);
nand U7542 (N_7542,N_7230,N_7358);
nand U7543 (N_7543,N_7260,N_7216);
nor U7544 (N_7544,N_7287,N_7216);
nand U7545 (N_7545,N_7214,N_7217);
nand U7546 (N_7546,N_7346,N_7291);
nand U7547 (N_7547,N_7313,N_7399);
nor U7548 (N_7548,N_7243,N_7398);
nor U7549 (N_7549,N_7307,N_7247);
nand U7550 (N_7550,N_7397,N_7295);
nand U7551 (N_7551,N_7397,N_7298);
or U7552 (N_7552,N_7332,N_7359);
nand U7553 (N_7553,N_7272,N_7292);
nor U7554 (N_7554,N_7300,N_7278);
nand U7555 (N_7555,N_7263,N_7261);
or U7556 (N_7556,N_7223,N_7337);
or U7557 (N_7557,N_7287,N_7298);
nor U7558 (N_7558,N_7260,N_7254);
nor U7559 (N_7559,N_7252,N_7217);
nor U7560 (N_7560,N_7381,N_7227);
and U7561 (N_7561,N_7379,N_7314);
and U7562 (N_7562,N_7347,N_7230);
nand U7563 (N_7563,N_7344,N_7330);
nand U7564 (N_7564,N_7281,N_7388);
nor U7565 (N_7565,N_7397,N_7288);
or U7566 (N_7566,N_7318,N_7260);
nor U7567 (N_7567,N_7381,N_7260);
and U7568 (N_7568,N_7321,N_7294);
nor U7569 (N_7569,N_7274,N_7319);
and U7570 (N_7570,N_7204,N_7367);
nand U7571 (N_7571,N_7326,N_7338);
nor U7572 (N_7572,N_7314,N_7359);
nand U7573 (N_7573,N_7389,N_7203);
and U7574 (N_7574,N_7236,N_7249);
nand U7575 (N_7575,N_7227,N_7246);
and U7576 (N_7576,N_7317,N_7227);
or U7577 (N_7577,N_7275,N_7296);
or U7578 (N_7578,N_7252,N_7201);
or U7579 (N_7579,N_7238,N_7230);
and U7580 (N_7580,N_7265,N_7386);
nand U7581 (N_7581,N_7304,N_7226);
or U7582 (N_7582,N_7340,N_7251);
or U7583 (N_7583,N_7214,N_7340);
or U7584 (N_7584,N_7280,N_7224);
nand U7585 (N_7585,N_7251,N_7388);
nand U7586 (N_7586,N_7268,N_7377);
or U7587 (N_7587,N_7380,N_7282);
or U7588 (N_7588,N_7384,N_7308);
nand U7589 (N_7589,N_7353,N_7208);
or U7590 (N_7590,N_7368,N_7282);
and U7591 (N_7591,N_7252,N_7244);
and U7592 (N_7592,N_7202,N_7392);
or U7593 (N_7593,N_7347,N_7312);
and U7594 (N_7594,N_7267,N_7234);
nor U7595 (N_7595,N_7279,N_7265);
nor U7596 (N_7596,N_7349,N_7346);
or U7597 (N_7597,N_7277,N_7355);
and U7598 (N_7598,N_7376,N_7227);
or U7599 (N_7599,N_7290,N_7356);
nand U7600 (N_7600,N_7537,N_7459);
or U7601 (N_7601,N_7415,N_7560);
nor U7602 (N_7602,N_7576,N_7559);
and U7603 (N_7603,N_7588,N_7512);
and U7604 (N_7604,N_7461,N_7578);
and U7605 (N_7605,N_7476,N_7465);
nand U7606 (N_7606,N_7555,N_7421);
or U7607 (N_7607,N_7529,N_7460);
nor U7608 (N_7608,N_7458,N_7597);
and U7609 (N_7609,N_7478,N_7556);
nor U7610 (N_7610,N_7433,N_7434);
or U7611 (N_7611,N_7590,N_7429);
nor U7612 (N_7612,N_7515,N_7492);
and U7613 (N_7613,N_7532,N_7577);
nand U7614 (N_7614,N_7466,N_7565);
or U7615 (N_7615,N_7518,N_7424);
nand U7616 (N_7616,N_7468,N_7447);
nor U7617 (N_7617,N_7451,N_7589);
or U7618 (N_7618,N_7536,N_7439);
nor U7619 (N_7619,N_7490,N_7413);
nor U7620 (N_7620,N_7475,N_7463);
nor U7621 (N_7621,N_7527,N_7551);
nand U7622 (N_7622,N_7530,N_7594);
and U7623 (N_7623,N_7405,N_7561);
nor U7624 (N_7624,N_7423,N_7418);
and U7625 (N_7625,N_7541,N_7535);
nor U7626 (N_7626,N_7484,N_7487);
and U7627 (N_7627,N_7571,N_7438);
or U7628 (N_7628,N_7514,N_7474);
nand U7629 (N_7629,N_7472,N_7402);
nand U7630 (N_7630,N_7428,N_7573);
and U7631 (N_7631,N_7443,N_7548);
nor U7632 (N_7632,N_7572,N_7400);
or U7633 (N_7633,N_7441,N_7470);
and U7634 (N_7634,N_7408,N_7549);
nand U7635 (N_7635,N_7403,N_7471);
or U7636 (N_7636,N_7473,N_7440);
nand U7637 (N_7637,N_7510,N_7483);
and U7638 (N_7638,N_7546,N_7427);
xor U7639 (N_7639,N_7509,N_7534);
or U7640 (N_7640,N_7455,N_7580);
or U7641 (N_7641,N_7505,N_7432);
nand U7642 (N_7642,N_7502,N_7584);
or U7643 (N_7643,N_7528,N_7491);
nor U7644 (N_7644,N_7442,N_7419);
nand U7645 (N_7645,N_7511,N_7416);
nand U7646 (N_7646,N_7596,N_7554);
nor U7647 (N_7647,N_7486,N_7569);
nor U7648 (N_7648,N_7482,N_7407);
or U7649 (N_7649,N_7409,N_7457);
or U7650 (N_7650,N_7498,N_7524);
and U7651 (N_7651,N_7422,N_7553);
nand U7652 (N_7652,N_7598,N_7489);
and U7653 (N_7653,N_7550,N_7480);
nand U7654 (N_7654,N_7464,N_7507);
or U7655 (N_7655,N_7496,N_7531);
and U7656 (N_7656,N_7436,N_7401);
nor U7657 (N_7657,N_7445,N_7404);
or U7658 (N_7658,N_7410,N_7493);
or U7659 (N_7659,N_7583,N_7599);
nand U7660 (N_7660,N_7503,N_7574);
nor U7661 (N_7661,N_7522,N_7513);
nand U7662 (N_7662,N_7446,N_7435);
nor U7663 (N_7663,N_7499,N_7414);
or U7664 (N_7664,N_7444,N_7456);
or U7665 (N_7665,N_7570,N_7595);
and U7666 (N_7666,N_7519,N_7430);
and U7667 (N_7667,N_7477,N_7431);
or U7668 (N_7668,N_7479,N_7517);
nand U7669 (N_7669,N_7540,N_7542);
or U7670 (N_7670,N_7591,N_7450);
and U7671 (N_7671,N_7582,N_7544);
nor U7672 (N_7672,N_7533,N_7547);
xnor U7673 (N_7673,N_7462,N_7425);
and U7674 (N_7674,N_7504,N_7500);
nor U7675 (N_7675,N_7501,N_7566);
nand U7676 (N_7676,N_7587,N_7545);
or U7677 (N_7677,N_7406,N_7526);
and U7678 (N_7678,N_7452,N_7467);
and U7679 (N_7679,N_7523,N_7568);
and U7680 (N_7680,N_7538,N_7506);
nor U7681 (N_7681,N_7411,N_7412);
and U7682 (N_7682,N_7495,N_7585);
and U7683 (N_7683,N_7567,N_7593);
and U7684 (N_7684,N_7437,N_7557);
or U7685 (N_7685,N_7485,N_7539);
nand U7686 (N_7686,N_7586,N_7488);
nand U7687 (N_7687,N_7417,N_7481);
nand U7688 (N_7688,N_7469,N_7449);
and U7689 (N_7689,N_7592,N_7453);
nand U7690 (N_7690,N_7520,N_7508);
nand U7691 (N_7691,N_7581,N_7575);
or U7692 (N_7692,N_7454,N_7494);
nor U7693 (N_7693,N_7497,N_7426);
and U7694 (N_7694,N_7525,N_7552);
and U7695 (N_7695,N_7420,N_7558);
or U7696 (N_7696,N_7516,N_7564);
nand U7697 (N_7697,N_7521,N_7543);
and U7698 (N_7698,N_7448,N_7579);
or U7699 (N_7699,N_7562,N_7563);
and U7700 (N_7700,N_7477,N_7452);
and U7701 (N_7701,N_7550,N_7475);
and U7702 (N_7702,N_7572,N_7544);
and U7703 (N_7703,N_7579,N_7484);
and U7704 (N_7704,N_7539,N_7455);
nor U7705 (N_7705,N_7512,N_7403);
nand U7706 (N_7706,N_7442,N_7441);
or U7707 (N_7707,N_7564,N_7404);
nor U7708 (N_7708,N_7527,N_7508);
or U7709 (N_7709,N_7552,N_7515);
or U7710 (N_7710,N_7587,N_7506);
and U7711 (N_7711,N_7434,N_7594);
nand U7712 (N_7712,N_7583,N_7440);
nand U7713 (N_7713,N_7466,N_7576);
and U7714 (N_7714,N_7405,N_7557);
nor U7715 (N_7715,N_7509,N_7403);
and U7716 (N_7716,N_7460,N_7550);
nor U7717 (N_7717,N_7585,N_7509);
or U7718 (N_7718,N_7540,N_7595);
or U7719 (N_7719,N_7518,N_7530);
or U7720 (N_7720,N_7464,N_7508);
or U7721 (N_7721,N_7485,N_7542);
and U7722 (N_7722,N_7547,N_7569);
nand U7723 (N_7723,N_7554,N_7417);
nor U7724 (N_7724,N_7560,N_7454);
nand U7725 (N_7725,N_7580,N_7575);
and U7726 (N_7726,N_7417,N_7499);
nand U7727 (N_7727,N_7474,N_7560);
and U7728 (N_7728,N_7584,N_7555);
nor U7729 (N_7729,N_7448,N_7525);
and U7730 (N_7730,N_7590,N_7554);
nand U7731 (N_7731,N_7514,N_7428);
and U7732 (N_7732,N_7421,N_7570);
nand U7733 (N_7733,N_7518,N_7431);
nand U7734 (N_7734,N_7592,N_7578);
nor U7735 (N_7735,N_7555,N_7414);
and U7736 (N_7736,N_7528,N_7597);
or U7737 (N_7737,N_7439,N_7411);
nor U7738 (N_7738,N_7443,N_7520);
and U7739 (N_7739,N_7440,N_7590);
or U7740 (N_7740,N_7562,N_7514);
nor U7741 (N_7741,N_7470,N_7497);
or U7742 (N_7742,N_7554,N_7499);
nand U7743 (N_7743,N_7562,N_7437);
and U7744 (N_7744,N_7551,N_7578);
nor U7745 (N_7745,N_7551,N_7488);
and U7746 (N_7746,N_7486,N_7558);
or U7747 (N_7747,N_7441,N_7447);
and U7748 (N_7748,N_7573,N_7547);
nor U7749 (N_7749,N_7414,N_7433);
and U7750 (N_7750,N_7562,N_7571);
nor U7751 (N_7751,N_7453,N_7498);
nand U7752 (N_7752,N_7457,N_7406);
and U7753 (N_7753,N_7591,N_7404);
nand U7754 (N_7754,N_7435,N_7471);
nand U7755 (N_7755,N_7462,N_7514);
or U7756 (N_7756,N_7456,N_7461);
nand U7757 (N_7757,N_7451,N_7516);
nand U7758 (N_7758,N_7437,N_7424);
or U7759 (N_7759,N_7572,N_7488);
nand U7760 (N_7760,N_7549,N_7492);
or U7761 (N_7761,N_7525,N_7533);
nand U7762 (N_7762,N_7488,N_7591);
xor U7763 (N_7763,N_7474,N_7481);
and U7764 (N_7764,N_7596,N_7439);
and U7765 (N_7765,N_7423,N_7571);
or U7766 (N_7766,N_7422,N_7524);
nor U7767 (N_7767,N_7528,N_7589);
or U7768 (N_7768,N_7461,N_7519);
or U7769 (N_7769,N_7454,N_7510);
nor U7770 (N_7770,N_7510,N_7402);
nand U7771 (N_7771,N_7574,N_7426);
nor U7772 (N_7772,N_7526,N_7591);
or U7773 (N_7773,N_7497,N_7435);
nor U7774 (N_7774,N_7592,N_7518);
nand U7775 (N_7775,N_7532,N_7420);
or U7776 (N_7776,N_7538,N_7403);
or U7777 (N_7777,N_7519,N_7537);
nor U7778 (N_7778,N_7444,N_7519);
nand U7779 (N_7779,N_7562,N_7443);
and U7780 (N_7780,N_7457,N_7547);
nand U7781 (N_7781,N_7520,N_7484);
or U7782 (N_7782,N_7551,N_7475);
and U7783 (N_7783,N_7537,N_7587);
nor U7784 (N_7784,N_7429,N_7419);
nor U7785 (N_7785,N_7480,N_7430);
and U7786 (N_7786,N_7460,N_7566);
nor U7787 (N_7787,N_7418,N_7545);
nor U7788 (N_7788,N_7551,N_7435);
or U7789 (N_7789,N_7491,N_7574);
and U7790 (N_7790,N_7537,N_7480);
and U7791 (N_7791,N_7505,N_7523);
or U7792 (N_7792,N_7487,N_7540);
or U7793 (N_7793,N_7526,N_7479);
nand U7794 (N_7794,N_7593,N_7523);
nor U7795 (N_7795,N_7499,N_7593);
nor U7796 (N_7796,N_7488,N_7509);
and U7797 (N_7797,N_7415,N_7427);
nand U7798 (N_7798,N_7570,N_7543);
nand U7799 (N_7799,N_7485,N_7533);
or U7800 (N_7800,N_7691,N_7697);
and U7801 (N_7801,N_7706,N_7789);
nand U7802 (N_7802,N_7748,N_7749);
or U7803 (N_7803,N_7687,N_7678);
and U7804 (N_7804,N_7710,N_7665);
nor U7805 (N_7805,N_7776,N_7640);
and U7806 (N_7806,N_7635,N_7680);
nand U7807 (N_7807,N_7699,N_7690);
nand U7808 (N_7808,N_7734,N_7775);
or U7809 (N_7809,N_7607,N_7617);
nor U7810 (N_7810,N_7661,N_7608);
nor U7811 (N_7811,N_7686,N_7646);
nand U7812 (N_7812,N_7703,N_7673);
nor U7813 (N_7813,N_7781,N_7630);
and U7814 (N_7814,N_7753,N_7747);
and U7815 (N_7815,N_7724,N_7723);
nor U7816 (N_7816,N_7681,N_7752);
nand U7817 (N_7817,N_7656,N_7799);
or U7818 (N_7818,N_7766,N_7797);
nor U7819 (N_7819,N_7662,N_7733);
or U7820 (N_7820,N_7639,N_7778);
nand U7821 (N_7821,N_7663,N_7725);
nand U7822 (N_7822,N_7658,N_7742);
nor U7823 (N_7823,N_7652,N_7705);
nor U7824 (N_7824,N_7768,N_7793);
or U7825 (N_7825,N_7784,N_7709);
nand U7826 (N_7826,N_7614,N_7738);
and U7827 (N_7827,N_7759,N_7745);
nor U7828 (N_7828,N_7667,N_7692);
nor U7829 (N_7829,N_7669,N_7717);
nor U7830 (N_7830,N_7758,N_7782);
nand U7831 (N_7831,N_7739,N_7712);
or U7832 (N_7832,N_7675,N_7715);
nor U7833 (N_7833,N_7701,N_7603);
or U7834 (N_7834,N_7610,N_7732);
and U7835 (N_7835,N_7679,N_7772);
nand U7836 (N_7836,N_7790,N_7633);
or U7837 (N_7837,N_7609,N_7666);
nor U7838 (N_7838,N_7629,N_7627);
nor U7839 (N_7839,N_7744,N_7693);
nand U7840 (N_7840,N_7743,N_7716);
and U7841 (N_7841,N_7719,N_7761);
or U7842 (N_7842,N_7769,N_7619);
nand U7843 (N_7843,N_7626,N_7688);
and U7844 (N_7844,N_7721,N_7726);
nor U7845 (N_7845,N_7700,N_7787);
and U7846 (N_7846,N_7774,N_7735);
and U7847 (N_7847,N_7668,N_7644);
and U7848 (N_7848,N_7720,N_7750);
nand U7849 (N_7849,N_7740,N_7685);
or U7850 (N_7850,N_7605,N_7643);
or U7851 (N_7851,N_7695,N_7730);
or U7852 (N_7852,N_7624,N_7677);
or U7853 (N_7853,N_7796,N_7674);
or U7854 (N_7854,N_7670,N_7648);
nor U7855 (N_7855,N_7751,N_7601);
or U7856 (N_7856,N_7762,N_7764);
nor U7857 (N_7857,N_7786,N_7671);
nand U7858 (N_7858,N_7754,N_7613);
or U7859 (N_7859,N_7647,N_7711);
nor U7860 (N_7860,N_7757,N_7632);
or U7861 (N_7861,N_7765,N_7637);
nand U7862 (N_7862,N_7713,N_7767);
and U7863 (N_7863,N_7746,N_7794);
nor U7864 (N_7864,N_7696,N_7631);
or U7865 (N_7865,N_7798,N_7783);
nand U7866 (N_7866,N_7650,N_7623);
and U7867 (N_7867,N_7756,N_7682);
nor U7868 (N_7868,N_7618,N_7676);
nor U7869 (N_7869,N_7620,N_7777);
nand U7870 (N_7870,N_7655,N_7628);
or U7871 (N_7871,N_7788,N_7763);
or U7872 (N_7872,N_7741,N_7651);
nor U7873 (N_7873,N_7664,N_7604);
or U7874 (N_7874,N_7642,N_7660);
or U7875 (N_7875,N_7731,N_7714);
nor U7876 (N_7876,N_7736,N_7616);
or U7877 (N_7877,N_7791,N_7636);
and U7878 (N_7878,N_7602,N_7773);
nor U7879 (N_7879,N_7785,N_7708);
or U7880 (N_7880,N_7702,N_7684);
or U7881 (N_7881,N_7760,N_7729);
or U7882 (N_7882,N_7645,N_7770);
and U7883 (N_7883,N_7649,N_7653);
and U7884 (N_7884,N_7718,N_7606);
nand U7885 (N_7885,N_7625,N_7722);
nand U7886 (N_7886,N_7792,N_7780);
nor U7887 (N_7887,N_7704,N_7615);
and U7888 (N_7888,N_7771,N_7728);
or U7889 (N_7889,N_7683,N_7698);
or U7890 (N_7890,N_7779,N_7641);
or U7891 (N_7891,N_7634,N_7612);
nand U7892 (N_7892,N_7621,N_7672);
nor U7893 (N_7893,N_7755,N_7694);
nor U7894 (N_7894,N_7600,N_7638);
and U7895 (N_7895,N_7737,N_7654);
nand U7896 (N_7896,N_7727,N_7659);
and U7897 (N_7897,N_7657,N_7795);
and U7898 (N_7898,N_7707,N_7689);
nor U7899 (N_7899,N_7611,N_7622);
or U7900 (N_7900,N_7763,N_7643);
nor U7901 (N_7901,N_7789,N_7600);
nor U7902 (N_7902,N_7673,N_7640);
nand U7903 (N_7903,N_7636,N_7681);
nand U7904 (N_7904,N_7613,N_7652);
and U7905 (N_7905,N_7692,N_7614);
nand U7906 (N_7906,N_7748,N_7702);
nand U7907 (N_7907,N_7750,N_7659);
and U7908 (N_7908,N_7693,N_7730);
nor U7909 (N_7909,N_7641,N_7618);
nor U7910 (N_7910,N_7627,N_7709);
nor U7911 (N_7911,N_7661,N_7711);
or U7912 (N_7912,N_7777,N_7675);
and U7913 (N_7913,N_7731,N_7664);
nand U7914 (N_7914,N_7675,N_7758);
nand U7915 (N_7915,N_7675,N_7770);
and U7916 (N_7916,N_7784,N_7662);
or U7917 (N_7917,N_7654,N_7645);
or U7918 (N_7918,N_7792,N_7671);
nand U7919 (N_7919,N_7695,N_7686);
nand U7920 (N_7920,N_7674,N_7678);
or U7921 (N_7921,N_7680,N_7684);
nand U7922 (N_7922,N_7769,N_7712);
nand U7923 (N_7923,N_7769,N_7650);
nor U7924 (N_7924,N_7676,N_7773);
nor U7925 (N_7925,N_7756,N_7783);
nor U7926 (N_7926,N_7758,N_7619);
or U7927 (N_7927,N_7796,N_7684);
or U7928 (N_7928,N_7606,N_7664);
nand U7929 (N_7929,N_7725,N_7737);
or U7930 (N_7930,N_7702,N_7765);
nand U7931 (N_7931,N_7682,N_7658);
nand U7932 (N_7932,N_7604,N_7759);
nor U7933 (N_7933,N_7739,N_7757);
nand U7934 (N_7934,N_7756,N_7672);
nor U7935 (N_7935,N_7736,N_7730);
nor U7936 (N_7936,N_7656,N_7733);
or U7937 (N_7937,N_7649,N_7640);
nand U7938 (N_7938,N_7610,N_7728);
or U7939 (N_7939,N_7608,N_7603);
or U7940 (N_7940,N_7629,N_7731);
or U7941 (N_7941,N_7675,N_7689);
nand U7942 (N_7942,N_7697,N_7619);
or U7943 (N_7943,N_7661,N_7725);
nor U7944 (N_7944,N_7721,N_7768);
xnor U7945 (N_7945,N_7756,N_7762);
nand U7946 (N_7946,N_7787,N_7751);
nor U7947 (N_7947,N_7648,N_7618);
and U7948 (N_7948,N_7755,N_7721);
nand U7949 (N_7949,N_7761,N_7775);
nand U7950 (N_7950,N_7742,N_7768);
nand U7951 (N_7951,N_7672,N_7648);
and U7952 (N_7952,N_7654,N_7605);
and U7953 (N_7953,N_7713,N_7611);
nand U7954 (N_7954,N_7738,N_7796);
nand U7955 (N_7955,N_7674,N_7701);
or U7956 (N_7956,N_7671,N_7637);
or U7957 (N_7957,N_7643,N_7775);
and U7958 (N_7958,N_7606,N_7647);
or U7959 (N_7959,N_7695,N_7676);
or U7960 (N_7960,N_7749,N_7760);
nor U7961 (N_7961,N_7716,N_7623);
and U7962 (N_7962,N_7608,N_7633);
nand U7963 (N_7963,N_7623,N_7606);
nand U7964 (N_7964,N_7617,N_7796);
or U7965 (N_7965,N_7707,N_7672);
and U7966 (N_7966,N_7643,N_7783);
nor U7967 (N_7967,N_7731,N_7728);
nand U7968 (N_7968,N_7707,N_7720);
nor U7969 (N_7969,N_7729,N_7611);
or U7970 (N_7970,N_7778,N_7786);
nand U7971 (N_7971,N_7719,N_7789);
or U7972 (N_7972,N_7750,N_7746);
or U7973 (N_7973,N_7626,N_7756);
nand U7974 (N_7974,N_7799,N_7735);
or U7975 (N_7975,N_7752,N_7754);
or U7976 (N_7976,N_7692,N_7606);
nor U7977 (N_7977,N_7680,N_7668);
and U7978 (N_7978,N_7739,N_7680);
and U7979 (N_7979,N_7642,N_7766);
and U7980 (N_7980,N_7704,N_7675);
or U7981 (N_7981,N_7626,N_7696);
nand U7982 (N_7982,N_7662,N_7664);
nand U7983 (N_7983,N_7662,N_7726);
nand U7984 (N_7984,N_7631,N_7716);
nand U7985 (N_7985,N_7689,N_7643);
nand U7986 (N_7986,N_7657,N_7783);
nand U7987 (N_7987,N_7698,N_7722);
nand U7988 (N_7988,N_7790,N_7647);
nor U7989 (N_7989,N_7708,N_7787);
or U7990 (N_7990,N_7647,N_7756);
nor U7991 (N_7991,N_7759,N_7741);
nor U7992 (N_7992,N_7797,N_7785);
and U7993 (N_7993,N_7608,N_7705);
or U7994 (N_7994,N_7614,N_7785);
and U7995 (N_7995,N_7672,N_7791);
nor U7996 (N_7996,N_7678,N_7785);
nand U7997 (N_7997,N_7661,N_7693);
nand U7998 (N_7998,N_7631,N_7751);
nor U7999 (N_7999,N_7725,N_7796);
and U8000 (N_8000,N_7843,N_7810);
nand U8001 (N_8001,N_7896,N_7935);
or U8002 (N_8002,N_7819,N_7900);
and U8003 (N_8003,N_7828,N_7844);
or U8004 (N_8004,N_7877,N_7841);
or U8005 (N_8005,N_7992,N_7822);
nand U8006 (N_8006,N_7874,N_7945);
nor U8007 (N_8007,N_7865,N_7805);
and U8008 (N_8008,N_7940,N_7813);
nor U8009 (N_8009,N_7821,N_7881);
nor U8010 (N_8010,N_7826,N_7839);
nand U8011 (N_8011,N_7946,N_7955);
and U8012 (N_8012,N_7908,N_7978);
nand U8013 (N_8013,N_7860,N_7985);
or U8014 (N_8014,N_7927,N_7885);
nand U8015 (N_8015,N_7818,N_7995);
and U8016 (N_8016,N_7933,N_7897);
nand U8017 (N_8017,N_7996,N_7975);
or U8018 (N_8018,N_7884,N_7876);
and U8019 (N_8019,N_7838,N_7820);
and U8020 (N_8020,N_7970,N_7943);
nand U8021 (N_8021,N_7903,N_7976);
or U8022 (N_8022,N_7949,N_7960);
and U8023 (N_8023,N_7859,N_7834);
and U8024 (N_8024,N_7981,N_7909);
nand U8025 (N_8025,N_7901,N_7952);
or U8026 (N_8026,N_7837,N_7921);
and U8027 (N_8027,N_7950,N_7801);
nand U8028 (N_8028,N_7845,N_7871);
and U8029 (N_8029,N_7967,N_7984);
or U8030 (N_8030,N_7962,N_7811);
and U8031 (N_8031,N_7961,N_7889);
nand U8032 (N_8032,N_7920,N_7808);
nand U8033 (N_8033,N_7911,N_7847);
or U8034 (N_8034,N_7895,N_7906);
or U8035 (N_8035,N_7938,N_7925);
nor U8036 (N_8036,N_7954,N_7868);
nor U8037 (N_8037,N_7890,N_7999);
or U8038 (N_8038,N_7983,N_7886);
nand U8039 (N_8039,N_7947,N_7833);
nor U8040 (N_8040,N_7831,N_7918);
and U8041 (N_8041,N_7968,N_7923);
nand U8042 (N_8042,N_7861,N_7836);
nor U8043 (N_8043,N_7803,N_7870);
nand U8044 (N_8044,N_7963,N_7817);
nor U8045 (N_8045,N_7806,N_7825);
or U8046 (N_8046,N_7892,N_7977);
nor U8047 (N_8047,N_7936,N_7849);
or U8048 (N_8048,N_7913,N_7807);
or U8049 (N_8049,N_7829,N_7934);
nand U8050 (N_8050,N_7848,N_7948);
and U8051 (N_8051,N_7815,N_7875);
and U8052 (N_8052,N_7854,N_7941);
nor U8053 (N_8053,N_7898,N_7907);
nor U8054 (N_8054,N_7855,N_7917);
and U8055 (N_8055,N_7988,N_7997);
or U8056 (N_8056,N_7846,N_7823);
nor U8057 (N_8057,N_7882,N_7969);
nand U8058 (N_8058,N_7851,N_7893);
nand U8059 (N_8059,N_7872,N_7878);
and U8060 (N_8060,N_7956,N_7850);
nor U8061 (N_8061,N_7916,N_7804);
or U8062 (N_8062,N_7816,N_7939);
nand U8063 (N_8063,N_7902,N_7899);
or U8064 (N_8064,N_7928,N_7842);
nand U8065 (N_8065,N_7852,N_7915);
nand U8066 (N_8066,N_7814,N_7991);
or U8067 (N_8067,N_7887,N_7986);
nor U8068 (N_8068,N_7924,N_7994);
or U8069 (N_8069,N_7971,N_7800);
nor U8070 (N_8070,N_7830,N_7922);
nor U8071 (N_8071,N_7951,N_7857);
or U8072 (N_8072,N_7926,N_7929);
and U8073 (N_8073,N_7891,N_7989);
nand U8074 (N_8074,N_7856,N_7932);
and U8075 (N_8075,N_7888,N_7824);
nor U8076 (N_8076,N_7862,N_7953);
or U8077 (N_8077,N_7979,N_7883);
or U8078 (N_8078,N_7993,N_7958);
and U8079 (N_8079,N_7864,N_7858);
or U8080 (N_8080,N_7937,N_7957);
or U8081 (N_8081,N_7980,N_7910);
nor U8082 (N_8082,N_7867,N_7990);
or U8083 (N_8083,N_7894,N_7944);
nand U8084 (N_8084,N_7840,N_7812);
or U8085 (N_8085,N_7879,N_7998);
nor U8086 (N_8086,N_7853,N_7904);
and U8087 (N_8087,N_7930,N_7942);
nor U8088 (N_8088,N_7919,N_7873);
nand U8089 (N_8089,N_7959,N_7974);
and U8090 (N_8090,N_7802,N_7931);
or U8091 (N_8091,N_7912,N_7972);
or U8092 (N_8092,N_7832,N_7905);
or U8093 (N_8093,N_7966,N_7880);
xor U8094 (N_8094,N_7863,N_7869);
or U8095 (N_8095,N_7973,N_7866);
and U8096 (N_8096,N_7964,N_7965);
or U8097 (N_8097,N_7914,N_7809);
nor U8098 (N_8098,N_7982,N_7987);
nor U8099 (N_8099,N_7835,N_7827);
nor U8100 (N_8100,N_7842,N_7944);
nor U8101 (N_8101,N_7964,N_7936);
nand U8102 (N_8102,N_7917,N_7874);
nand U8103 (N_8103,N_7986,N_7814);
and U8104 (N_8104,N_7901,N_7804);
nand U8105 (N_8105,N_7954,N_7953);
nor U8106 (N_8106,N_7948,N_7992);
nand U8107 (N_8107,N_7894,N_7803);
nand U8108 (N_8108,N_7966,N_7915);
nor U8109 (N_8109,N_7983,N_7829);
nand U8110 (N_8110,N_7970,N_7897);
or U8111 (N_8111,N_7871,N_7978);
nor U8112 (N_8112,N_7987,N_7812);
or U8113 (N_8113,N_7911,N_7828);
nor U8114 (N_8114,N_7867,N_7835);
or U8115 (N_8115,N_7885,N_7811);
and U8116 (N_8116,N_7888,N_7932);
and U8117 (N_8117,N_7949,N_7822);
nor U8118 (N_8118,N_7872,N_7959);
and U8119 (N_8119,N_7914,N_7951);
and U8120 (N_8120,N_7832,N_7955);
nand U8121 (N_8121,N_7828,N_7880);
nand U8122 (N_8122,N_7808,N_7885);
and U8123 (N_8123,N_7862,N_7979);
and U8124 (N_8124,N_7944,N_7982);
nor U8125 (N_8125,N_7924,N_7847);
or U8126 (N_8126,N_7870,N_7852);
nand U8127 (N_8127,N_7871,N_7908);
nor U8128 (N_8128,N_7918,N_7824);
nor U8129 (N_8129,N_7880,N_7829);
or U8130 (N_8130,N_7977,N_7985);
nor U8131 (N_8131,N_7931,N_7979);
and U8132 (N_8132,N_7940,N_7923);
and U8133 (N_8133,N_7899,N_7878);
or U8134 (N_8134,N_7985,N_7803);
or U8135 (N_8135,N_7987,N_7981);
nand U8136 (N_8136,N_7975,N_7847);
or U8137 (N_8137,N_7848,N_7952);
nor U8138 (N_8138,N_7909,N_7921);
or U8139 (N_8139,N_7953,N_7822);
nand U8140 (N_8140,N_7949,N_7902);
or U8141 (N_8141,N_7860,N_7937);
and U8142 (N_8142,N_7918,N_7830);
and U8143 (N_8143,N_7806,N_7845);
nor U8144 (N_8144,N_7921,N_7997);
or U8145 (N_8145,N_7989,N_7980);
or U8146 (N_8146,N_7850,N_7857);
and U8147 (N_8147,N_7904,N_7989);
or U8148 (N_8148,N_7870,N_7942);
or U8149 (N_8149,N_7815,N_7895);
nor U8150 (N_8150,N_7995,N_7998);
nand U8151 (N_8151,N_7864,N_7828);
nand U8152 (N_8152,N_7861,N_7915);
or U8153 (N_8153,N_7945,N_7849);
nand U8154 (N_8154,N_7986,N_7920);
nor U8155 (N_8155,N_7949,N_7995);
xor U8156 (N_8156,N_7934,N_7859);
or U8157 (N_8157,N_7852,N_7848);
nor U8158 (N_8158,N_7981,N_7952);
and U8159 (N_8159,N_7886,N_7966);
nor U8160 (N_8160,N_7948,N_7994);
nand U8161 (N_8161,N_7937,N_7978);
or U8162 (N_8162,N_7862,N_7824);
nand U8163 (N_8163,N_7976,N_7876);
nor U8164 (N_8164,N_7859,N_7899);
or U8165 (N_8165,N_7956,N_7892);
and U8166 (N_8166,N_7959,N_7915);
nor U8167 (N_8167,N_7875,N_7887);
nor U8168 (N_8168,N_7809,N_7884);
and U8169 (N_8169,N_7932,N_7939);
and U8170 (N_8170,N_7900,N_7802);
or U8171 (N_8171,N_7992,N_7801);
and U8172 (N_8172,N_7932,N_7852);
or U8173 (N_8173,N_7946,N_7972);
nor U8174 (N_8174,N_7840,N_7885);
nor U8175 (N_8175,N_7819,N_7954);
and U8176 (N_8176,N_7964,N_7904);
nor U8177 (N_8177,N_7870,N_7941);
nand U8178 (N_8178,N_7950,N_7911);
nor U8179 (N_8179,N_7819,N_7907);
or U8180 (N_8180,N_7887,N_7806);
and U8181 (N_8181,N_7875,N_7884);
nand U8182 (N_8182,N_7968,N_7862);
nor U8183 (N_8183,N_7973,N_7889);
or U8184 (N_8184,N_7826,N_7814);
or U8185 (N_8185,N_7812,N_7887);
nor U8186 (N_8186,N_7829,N_7847);
and U8187 (N_8187,N_7977,N_7912);
or U8188 (N_8188,N_7806,N_7871);
or U8189 (N_8189,N_7891,N_7978);
nor U8190 (N_8190,N_7865,N_7812);
and U8191 (N_8191,N_7814,N_7989);
nand U8192 (N_8192,N_7864,N_7955);
nand U8193 (N_8193,N_7846,N_7975);
nor U8194 (N_8194,N_7844,N_7832);
or U8195 (N_8195,N_7972,N_7862);
nand U8196 (N_8196,N_7888,N_7809);
nor U8197 (N_8197,N_7984,N_7835);
or U8198 (N_8198,N_7971,N_7984);
or U8199 (N_8199,N_7800,N_7877);
and U8200 (N_8200,N_8174,N_8156);
and U8201 (N_8201,N_8050,N_8008);
or U8202 (N_8202,N_8163,N_8171);
or U8203 (N_8203,N_8124,N_8067);
nand U8204 (N_8204,N_8136,N_8196);
and U8205 (N_8205,N_8164,N_8035);
or U8206 (N_8206,N_8023,N_8009);
nor U8207 (N_8207,N_8143,N_8028);
nand U8208 (N_8208,N_8186,N_8061);
and U8209 (N_8209,N_8178,N_8165);
or U8210 (N_8210,N_8104,N_8056);
or U8211 (N_8211,N_8007,N_8134);
nor U8212 (N_8212,N_8103,N_8059);
nand U8213 (N_8213,N_8013,N_8139);
nor U8214 (N_8214,N_8058,N_8072);
nor U8215 (N_8215,N_8005,N_8141);
nand U8216 (N_8216,N_8181,N_8096);
or U8217 (N_8217,N_8167,N_8112);
nand U8218 (N_8218,N_8052,N_8199);
and U8219 (N_8219,N_8049,N_8102);
or U8220 (N_8220,N_8019,N_8033);
nand U8221 (N_8221,N_8119,N_8173);
and U8222 (N_8222,N_8155,N_8159);
nand U8223 (N_8223,N_8114,N_8083);
and U8224 (N_8224,N_8168,N_8099);
and U8225 (N_8225,N_8182,N_8197);
or U8226 (N_8226,N_8161,N_8047);
nor U8227 (N_8227,N_8020,N_8079);
and U8228 (N_8228,N_8026,N_8138);
nand U8229 (N_8229,N_8110,N_8031);
or U8230 (N_8230,N_8145,N_8169);
nor U8231 (N_8231,N_8085,N_8120);
or U8232 (N_8232,N_8027,N_8045);
and U8233 (N_8233,N_8063,N_8011);
or U8234 (N_8234,N_8021,N_8041);
or U8235 (N_8235,N_8188,N_8088);
and U8236 (N_8236,N_8093,N_8038);
and U8237 (N_8237,N_8122,N_8060);
and U8238 (N_8238,N_8131,N_8001);
nand U8239 (N_8239,N_8068,N_8195);
nor U8240 (N_8240,N_8091,N_8098);
or U8241 (N_8241,N_8046,N_8125);
nor U8242 (N_8242,N_8109,N_8087);
nor U8243 (N_8243,N_8121,N_8025);
or U8244 (N_8244,N_8128,N_8132);
nor U8245 (N_8245,N_8166,N_8123);
nand U8246 (N_8246,N_8017,N_8014);
nor U8247 (N_8247,N_8151,N_8185);
and U8248 (N_8248,N_8157,N_8016);
and U8249 (N_8249,N_8154,N_8127);
and U8250 (N_8250,N_8111,N_8012);
nand U8251 (N_8251,N_8160,N_8010);
and U8252 (N_8252,N_8090,N_8042);
nor U8253 (N_8253,N_8133,N_8053);
and U8254 (N_8254,N_8004,N_8153);
nor U8255 (N_8255,N_8094,N_8177);
nand U8256 (N_8256,N_8101,N_8022);
nand U8257 (N_8257,N_8000,N_8149);
or U8258 (N_8258,N_8064,N_8106);
nor U8259 (N_8259,N_8066,N_8089);
nor U8260 (N_8260,N_8002,N_8076);
nor U8261 (N_8261,N_8162,N_8032);
nand U8262 (N_8262,N_8084,N_8180);
nor U8263 (N_8263,N_8176,N_8054);
nor U8264 (N_8264,N_8148,N_8191);
or U8265 (N_8265,N_8034,N_8092);
nand U8266 (N_8266,N_8116,N_8187);
or U8267 (N_8267,N_8043,N_8140);
or U8268 (N_8268,N_8040,N_8044);
nor U8269 (N_8269,N_8172,N_8147);
and U8270 (N_8270,N_8105,N_8073);
and U8271 (N_8271,N_8137,N_8108);
and U8272 (N_8272,N_8184,N_8158);
nor U8273 (N_8273,N_8037,N_8082);
or U8274 (N_8274,N_8036,N_8065);
or U8275 (N_8275,N_8057,N_8095);
nor U8276 (N_8276,N_8077,N_8150);
and U8277 (N_8277,N_8080,N_8029);
nor U8278 (N_8278,N_8100,N_8117);
or U8279 (N_8279,N_8051,N_8135);
nand U8280 (N_8280,N_8189,N_8048);
or U8281 (N_8281,N_8015,N_8193);
nand U8282 (N_8282,N_8144,N_8194);
or U8283 (N_8283,N_8107,N_8097);
and U8284 (N_8284,N_8086,N_8146);
or U8285 (N_8285,N_8115,N_8183);
and U8286 (N_8286,N_8190,N_8081);
nor U8287 (N_8287,N_8113,N_8070);
nor U8288 (N_8288,N_8179,N_8030);
and U8289 (N_8289,N_8192,N_8130);
or U8290 (N_8290,N_8074,N_8075);
or U8291 (N_8291,N_8069,N_8170);
nor U8292 (N_8292,N_8039,N_8118);
nand U8293 (N_8293,N_8129,N_8006);
nand U8294 (N_8294,N_8024,N_8003);
nor U8295 (N_8295,N_8198,N_8078);
nand U8296 (N_8296,N_8175,N_8018);
nand U8297 (N_8297,N_8062,N_8152);
nor U8298 (N_8298,N_8055,N_8126);
or U8299 (N_8299,N_8071,N_8142);
nor U8300 (N_8300,N_8130,N_8132);
nand U8301 (N_8301,N_8124,N_8050);
or U8302 (N_8302,N_8108,N_8161);
nand U8303 (N_8303,N_8020,N_8031);
nand U8304 (N_8304,N_8135,N_8155);
nor U8305 (N_8305,N_8009,N_8187);
or U8306 (N_8306,N_8075,N_8015);
and U8307 (N_8307,N_8169,N_8119);
or U8308 (N_8308,N_8176,N_8081);
nand U8309 (N_8309,N_8133,N_8187);
and U8310 (N_8310,N_8182,N_8163);
nor U8311 (N_8311,N_8058,N_8013);
nor U8312 (N_8312,N_8079,N_8016);
and U8313 (N_8313,N_8088,N_8014);
nand U8314 (N_8314,N_8057,N_8163);
nor U8315 (N_8315,N_8100,N_8004);
or U8316 (N_8316,N_8035,N_8159);
and U8317 (N_8317,N_8136,N_8109);
and U8318 (N_8318,N_8197,N_8045);
and U8319 (N_8319,N_8095,N_8168);
or U8320 (N_8320,N_8149,N_8065);
or U8321 (N_8321,N_8039,N_8090);
or U8322 (N_8322,N_8167,N_8001);
and U8323 (N_8323,N_8014,N_8022);
and U8324 (N_8324,N_8158,N_8126);
or U8325 (N_8325,N_8114,N_8007);
or U8326 (N_8326,N_8153,N_8178);
nor U8327 (N_8327,N_8031,N_8170);
and U8328 (N_8328,N_8087,N_8078);
and U8329 (N_8329,N_8022,N_8131);
or U8330 (N_8330,N_8116,N_8096);
and U8331 (N_8331,N_8096,N_8163);
or U8332 (N_8332,N_8188,N_8026);
nand U8333 (N_8333,N_8011,N_8110);
nand U8334 (N_8334,N_8133,N_8003);
nor U8335 (N_8335,N_8138,N_8100);
or U8336 (N_8336,N_8036,N_8024);
and U8337 (N_8337,N_8161,N_8136);
and U8338 (N_8338,N_8165,N_8175);
and U8339 (N_8339,N_8145,N_8035);
nand U8340 (N_8340,N_8100,N_8180);
and U8341 (N_8341,N_8008,N_8042);
nor U8342 (N_8342,N_8012,N_8093);
or U8343 (N_8343,N_8086,N_8014);
nor U8344 (N_8344,N_8097,N_8130);
nor U8345 (N_8345,N_8133,N_8102);
nor U8346 (N_8346,N_8183,N_8192);
nor U8347 (N_8347,N_8092,N_8098);
nand U8348 (N_8348,N_8160,N_8029);
or U8349 (N_8349,N_8181,N_8108);
and U8350 (N_8350,N_8064,N_8177);
nand U8351 (N_8351,N_8055,N_8085);
nor U8352 (N_8352,N_8001,N_8030);
nor U8353 (N_8353,N_8102,N_8183);
or U8354 (N_8354,N_8021,N_8068);
and U8355 (N_8355,N_8093,N_8054);
nor U8356 (N_8356,N_8060,N_8138);
or U8357 (N_8357,N_8069,N_8137);
nor U8358 (N_8358,N_8179,N_8079);
nor U8359 (N_8359,N_8061,N_8060);
and U8360 (N_8360,N_8050,N_8098);
nor U8361 (N_8361,N_8096,N_8135);
nand U8362 (N_8362,N_8103,N_8147);
nand U8363 (N_8363,N_8053,N_8061);
nor U8364 (N_8364,N_8043,N_8177);
nand U8365 (N_8365,N_8142,N_8043);
and U8366 (N_8366,N_8147,N_8036);
and U8367 (N_8367,N_8141,N_8015);
nand U8368 (N_8368,N_8161,N_8186);
nor U8369 (N_8369,N_8125,N_8083);
nor U8370 (N_8370,N_8006,N_8117);
or U8371 (N_8371,N_8043,N_8158);
or U8372 (N_8372,N_8102,N_8180);
nand U8373 (N_8373,N_8136,N_8056);
nand U8374 (N_8374,N_8175,N_8016);
nor U8375 (N_8375,N_8169,N_8115);
and U8376 (N_8376,N_8170,N_8160);
nand U8377 (N_8377,N_8153,N_8075);
nand U8378 (N_8378,N_8136,N_8028);
or U8379 (N_8379,N_8013,N_8120);
or U8380 (N_8380,N_8072,N_8001);
nand U8381 (N_8381,N_8071,N_8178);
nor U8382 (N_8382,N_8041,N_8068);
and U8383 (N_8383,N_8170,N_8050);
nand U8384 (N_8384,N_8095,N_8038);
and U8385 (N_8385,N_8027,N_8089);
or U8386 (N_8386,N_8000,N_8051);
nand U8387 (N_8387,N_8047,N_8080);
nor U8388 (N_8388,N_8007,N_8087);
or U8389 (N_8389,N_8193,N_8112);
nor U8390 (N_8390,N_8148,N_8130);
or U8391 (N_8391,N_8000,N_8083);
or U8392 (N_8392,N_8077,N_8175);
or U8393 (N_8393,N_8126,N_8191);
nor U8394 (N_8394,N_8184,N_8037);
nand U8395 (N_8395,N_8183,N_8030);
nor U8396 (N_8396,N_8172,N_8134);
and U8397 (N_8397,N_8110,N_8016);
or U8398 (N_8398,N_8142,N_8129);
nor U8399 (N_8399,N_8054,N_8056);
nor U8400 (N_8400,N_8267,N_8388);
or U8401 (N_8401,N_8234,N_8231);
nand U8402 (N_8402,N_8366,N_8376);
and U8403 (N_8403,N_8212,N_8389);
or U8404 (N_8404,N_8299,N_8256);
nor U8405 (N_8405,N_8217,N_8393);
nor U8406 (N_8406,N_8283,N_8312);
or U8407 (N_8407,N_8352,N_8247);
nor U8408 (N_8408,N_8249,N_8361);
or U8409 (N_8409,N_8271,N_8258);
nand U8410 (N_8410,N_8297,N_8300);
nand U8411 (N_8411,N_8296,N_8244);
nand U8412 (N_8412,N_8208,N_8282);
nor U8413 (N_8413,N_8224,N_8370);
nor U8414 (N_8414,N_8209,N_8240);
or U8415 (N_8415,N_8202,N_8276);
nor U8416 (N_8416,N_8291,N_8230);
and U8417 (N_8417,N_8223,N_8353);
nand U8418 (N_8418,N_8338,N_8242);
or U8419 (N_8419,N_8371,N_8394);
or U8420 (N_8420,N_8266,N_8399);
and U8421 (N_8421,N_8205,N_8243);
nand U8422 (N_8422,N_8285,N_8301);
nand U8423 (N_8423,N_8257,N_8277);
nand U8424 (N_8424,N_8313,N_8226);
nor U8425 (N_8425,N_8211,N_8375);
nand U8426 (N_8426,N_8236,N_8333);
nand U8427 (N_8427,N_8324,N_8325);
nor U8428 (N_8428,N_8263,N_8303);
and U8429 (N_8429,N_8369,N_8397);
nor U8430 (N_8430,N_8377,N_8354);
nor U8431 (N_8431,N_8311,N_8289);
and U8432 (N_8432,N_8274,N_8248);
nor U8433 (N_8433,N_8329,N_8278);
xnor U8434 (N_8434,N_8265,N_8279);
nand U8435 (N_8435,N_8384,N_8293);
and U8436 (N_8436,N_8382,N_8241);
and U8437 (N_8437,N_8239,N_8385);
or U8438 (N_8438,N_8328,N_8395);
nand U8439 (N_8439,N_8339,N_8229);
or U8440 (N_8440,N_8367,N_8356);
nor U8441 (N_8441,N_8380,N_8306);
or U8442 (N_8442,N_8343,N_8259);
nor U8443 (N_8443,N_8372,N_8348);
or U8444 (N_8444,N_8355,N_8294);
and U8445 (N_8445,N_8310,N_8307);
xnor U8446 (N_8446,N_8268,N_8316);
nand U8447 (N_8447,N_8270,N_8336);
or U8448 (N_8448,N_8201,N_8213);
nor U8449 (N_8449,N_8381,N_8308);
or U8450 (N_8450,N_8320,N_8281);
nand U8451 (N_8451,N_8292,N_8323);
and U8452 (N_8452,N_8326,N_8390);
and U8453 (N_8453,N_8254,N_8344);
xor U8454 (N_8454,N_8346,N_8261);
nor U8455 (N_8455,N_8221,N_8364);
or U8456 (N_8456,N_8318,N_8387);
nand U8457 (N_8457,N_8347,N_8215);
or U8458 (N_8458,N_8284,N_8246);
nor U8459 (N_8459,N_8272,N_8349);
nand U8460 (N_8460,N_8360,N_8218);
and U8461 (N_8461,N_8396,N_8332);
nand U8462 (N_8462,N_8378,N_8327);
or U8463 (N_8463,N_8341,N_8335);
nand U8464 (N_8464,N_8262,N_8351);
nor U8465 (N_8465,N_8309,N_8363);
or U8466 (N_8466,N_8200,N_8379);
nor U8467 (N_8467,N_8286,N_8368);
or U8468 (N_8468,N_8227,N_8322);
or U8469 (N_8469,N_8304,N_8255);
or U8470 (N_8470,N_8359,N_8222);
nand U8471 (N_8471,N_8383,N_8275);
nor U8472 (N_8472,N_8362,N_8340);
or U8473 (N_8473,N_8319,N_8225);
nor U8474 (N_8474,N_8251,N_8305);
or U8475 (N_8475,N_8295,N_8330);
nand U8476 (N_8476,N_8302,N_8391);
nor U8477 (N_8477,N_8264,N_8214);
nand U8478 (N_8478,N_8238,N_8334);
nand U8479 (N_8479,N_8337,N_8210);
or U8480 (N_8480,N_8216,N_8252);
and U8481 (N_8481,N_8287,N_8220);
or U8482 (N_8482,N_8253,N_8269);
nand U8483 (N_8483,N_8373,N_8398);
nand U8484 (N_8484,N_8290,N_8206);
or U8485 (N_8485,N_8315,N_8260);
nand U8486 (N_8486,N_8321,N_8237);
nand U8487 (N_8487,N_8374,N_8207);
or U8488 (N_8488,N_8288,N_8314);
or U8489 (N_8489,N_8204,N_8350);
nand U8490 (N_8490,N_8317,N_8280);
nand U8491 (N_8491,N_8228,N_8235);
and U8492 (N_8492,N_8358,N_8203);
or U8493 (N_8493,N_8219,N_8245);
or U8494 (N_8494,N_8298,N_8386);
or U8495 (N_8495,N_8250,N_8232);
or U8496 (N_8496,N_8331,N_8342);
or U8497 (N_8497,N_8365,N_8273);
or U8498 (N_8498,N_8345,N_8357);
and U8499 (N_8499,N_8392,N_8233);
nand U8500 (N_8500,N_8256,N_8213);
nor U8501 (N_8501,N_8375,N_8350);
nand U8502 (N_8502,N_8285,N_8399);
or U8503 (N_8503,N_8215,N_8308);
or U8504 (N_8504,N_8362,N_8367);
and U8505 (N_8505,N_8295,N_8299);
or U8506 (N_8506,N_8336,N_8321);
nand U8507 (N_8507,N_8290,N_8386);
and U8508 (N_8508,N_8367,N_8325);
nand U8509 (N_8509,N_8242,N_8216);
nor U8510 (N_8510,N_8360,N_8381);
nand U8511 (N_8511,N_8227,N_8202);
nor U8512 (N_8512,N_8377,N_8319);
and U8513 (N_8513,N_8326,N_8296);
and U8514 (N_8514,N_8235,N_8299);
nand U8515 (N_8515,N_8389,N_8335);
nand U8516 (N_8516,N_8265,N_8341);
or U8517 (N_8517,N_8353,N_8398);
nor U8518 (N_8518,N_8213,N_8317);
xor U8519 (N_8519,N_8239,N_8295);
and U8520 (N_8520,N_8286,N_8283);
and U8521 (N_8521,N_8376,N_8266);
nand U8522 (N_8522,N_8226,N_8333);
nand U8523 (N_8523,N_8388,N_8244);
nand U8524 (N_8524,N_8268,N_8396);
or U8525 (N_8525,N_8278,N_8275);
or U8526 (N_8526,N_8398,N_8396);
and U8527 (N_8527,N_8394,N_8285);
or U8528 (N_8528,N_8358,N_8264);
nor U8529 (N_8529,N_8299,N_8317);
and U8530 (N_8530,N_8219,N_8217);
and U8531 (N_8531,N_8316,N_8208);
and U8532 (N_8532,N_8294,N_8234);
or U8533 (N_8533,N_8392,N_8340);
nand U8534 (N_8534,N_8380,N_8203);
or U8535 (N_8535,N_8304,N_8306);
nor U8536 (N_8536,N_8255,N_8250);
nand U8537 (N_8537,N_8388,N_8309);
nor U8538 (N_8538,N_8341,N_8295);
nand U8539 (N_8539,N_8232,N_8328);
and U8540 (N_8540,N_8273,N_8341);
nor U8541 (N_8541,N_8283,N_8293);
and U8542 (N_8542,N_8367,N_8274);
and U8543 (N_8543,N_8327,N_8354);
and U8544 (N_8544,N_8315,N_8362);
and U8545 (N_8545,N_8288,N_8226);
and U8546 (N_8546,N_8277,N_8348);
and U8547 (N_8547,N_8223,N_8344);
or U8548 (N_8548,N_8288,N_8263);
or U8549 (N_8549,N_8343,N_8302);
nor U8550 (N_8550,N_8279,N_8361);
and U8551 (N_8551,N_8386,N_8353);
nand U8552 (N_8552,N_8241,N_8274);
or U8553 (N_8553,N_8246,N_8256);
and U8554 (N_8554,N_8329,N_8357);
nand U8555 (N_8555,N_8319,N_8349);
or U8556 (N_8556,N_8238,N_8273);
nor U8557 (N_8557,N_8228,N_8329);
nor U8558 (N_8558,N_8254,N_8392);
nand U8559 (N_8559,N_8258,N_8241);
nor U8560 (N_8560,N_8337,N_8360);
and U8561 (N_8561,N_8292,N_8389);
nand U8562 (N_8562,N_8343,N_8360);
nand U8563 (N_8563,N_8332,N_8380);
nor U8564 (N_8564,N_8361,N_8387);
and U8565 (N_8565,N_8292,N_8296);
nor U8566 (N_8566,N_8241,N_8378);
nor U8567 (N_8567,N_8299,N_8298);
xnor U8568 (N_8568,N_8382,N_8383);
or U8569 (N_8569,N_8233,N_8313);
and U8570 (N_8570,N_8370,N_8275);
nand U8571 (N_8571,N_8337,N_8248);
nor U8572 (N_8572,N_8379,N_8375);
xor U8573 (N_8573,N_8211,N_8248);
nand U8574 (N_8574,N_8237,N_8370);
and U8575 (N_8575,N_8225,N_8277);
nor U8576 (N_8576,N_8355,N_8316);
and U8577 (N_8577,N_8253,N_8239);
nand U8578 (N_8578,N_8323,N_8346);
and U8579 (N_8579,N_8236,N_8256);
nand U8580 (N_8580,N_8359,N_8361);
nor U8581 (N_8581,N_8288,N_8205);
nor U8582 (N_8582,N_8355,N_8377);
and U8583 (N_8583,N_8263,N_8356);
nor U8584 (N_8584,N_8253,N_8360);
nand U8585 (N_8585,N_8259,N_8220);
nand U8586 (N_8586,N_8368,N_8275);
nor U8587 (N_8587,N_8355,N_8312);
xnor U8588 (N_8588,N_8380,N_8365);
nor U8589 (N_8589,N_8372,N_8367);
nor U8590 (N_8590,N_8366,N_8330);
nand U8591 (N_8591,N_8224,N_8290);
nand U8592 (N_8592,N_8396,N_8393);
nor U8593 (N_8593,N_8295,N_8225);
and U8594 (N_8594,N_8302,N_8292);
and U8595 (N_8595,N_8383,N_8243);
nor U8596 (N_8596,N_8247,N_8277);
nand U8597 (N_8597,N_8384,N_8271);
or U8598 (N_8598,N_8279,N_8242);
or U8599 (N_8599,N_8225,N_8392);
and U8600 (N_8600,N_8434,N_8500);
xor U8601 (N_8601,N_8591,N_8425);
and U8602 (N_8602,N_8578,N_8439);
and U8603 (N_8603,N_8420,N_8543);
or U8604 (N_8604,N_8482,N_8505);
and U8605 (N_8605,N_8414,N_8501);
or U8606 (N_8606,N_8597,N_8528);
and U8607 (N_8607,N_8585,N_8484);
nor U8608 (N_8608,N_8407,N_8475);
and U8609 (N_8609,N_8447,N_8523);
nor U8610 (N_8610,N_8530,N_8562);
nand U8611 (N_8611,N_8461,N_8454);
nor U8612 (N_8612,N_8552,N_8557);
nand U8613 (N_8613,N_8438,N_8563);
nor U8614 (N_8614,N_8512,N_8419);
and U8615 (N_8615,N_8479,N_8429);
nor U8616 (N_8616,N_8506,N_8508);
nor U8617 (N_8617,N_8430,N_8404);
and U8618 (N_8618,N_8464,N_8435);
and U8619 (N_8619,N_8402,N_8558);
and U8620 (N_8620,N_8589,N_8415);
nand U8621 (N_8621,N_8426,N_8443);
and U8622 (N_8622,N_8445,N_8536);
and U8623 (N_8623,N_8599,N_8514);
nor U8624 (N_8624,N_8452,N_8521);
nand U8625 (N_8625,N_8564,N_8453);
or U8626 (N_8626,N_8499,N_8551);
or U8627 (N_8627,N_8590,N_8569);
or U8628 (N_8628,N_8567,N_8527);
nand U8629 (N_8629,N_8574,N_8579);
and U8630 (N_8630,N_8568,N_8587);
nor U8631 (N_8631,N_8525,N_8565);
nand U8632 (N_8632,N_8465,N_8549);
nand U8633 (N_8633,N_8532,N_8483);
nand U8634 (N_8634,N_8513,N_8497);
nand U8635 (N_8635,N_8400,N_8517);
nand U8636 (N_8636,N_8441,N_8580);
nand U8637 (N_8637,N_8442,N_8494);
or U8638 (N_8638,N_8553,N_8518);
or U8639 (N_8639,N_8486,N_8418);
nor U8640 (N_8640,N_8531,N_8421);
and U8641 (N_8641,N_8493,N_8432);
or U8642 (N_8642,N_8411,N_8490);
or U8643 (N_8643,N_8408,N_8427);
or U8644 (N_8644,N_8509,N_8598);
nand U8645 (N_8645,N_8462,N_8582);
nor U8646 (N_8646,N_8594,N_8540);
nand U8647 (N_8647,N_8586,N_8539);
nand U8648 (N_8648,N_8477,N_8417);
or U8649 (N_8649,N_8476,N_8480);
or U8650 (N_8650,N_8529,N_8489);
nor U8651 (N_8651,N_8538,N_8547);
and U8652 (N_8652,N_8511,N_8572);
nor U8653 (N_8653,N_8466,N_8588);
and U8654 (N_8654,N_8533,N_8428);
or U8655 (N_8655,N_8449,N_8584);
nor U8656 (N_8656,N_8592,N_8503);
nand U8657 (N_8657,N_8405,N_8556);
nor U8658 (N_8658,N_8502,N_8422);
or U8659 (N_8659,N_8423,N_8520);
or U8660 (N_8660,N_8581,N_8444);
nand U8661 (N_8661,N_8491,N_8460);
or U8662 (N_8662,N_8577,N_8575);
and U8663 (N_8663,N_8555,N_8488);
or U8664 (N_8664,N_8560,N_8535);
or U8665 (N_8665,N_8515,N_8448);
and U8666 (N_8666,N_8596,N_8576);
or U8667 (N_8667,N_8450,N_8406);
nand U8668 (N_8668,N_8537,N_8478);
nand U8669 (N_8669,N_8534,N_8456);
nor U8670 (N_8670,N_8595,N_8496);
or U8671 (N_8671,N_8548,N_8455);
and U8672 (N_8672,N_8433,N_8492);
and U8673 (N_8673,N_8545,N_8473);
nor U8674 (N_8674,N_8472,N_8554);
nand U8675 (N_8675,N_8424,N_8573);
or U8676 (N_8676,N_8437,N_8459);
and U8677 (N_8677,N_8458,N_8436);
or U8678 (N_8678,N_8504,N_8446);
nand U8679 (N_8679,N_8481,N_8566);
nor U8680 (N_8680,N_8487,N_8468);
nor U8681 (N_8681,N_8559,N_8469);
and U8682 (N_8682,N_8413,N_8516);
or U8683 (N_8683,N_8416,N_8463);
xnor U8684 (N_8684,N_8471,N_8403);
and U8685 (N_8685,N_8550,N_8495);
or U8686 (N_8686,N_8410,N_8474);
nor U8687 (N_8687,N_8544,N_8526);
nor U8688 (N_8688,N_8457,N_8561);
nand U8689 (N_8689,N_8507,N_8467);
and U8690 (N_8690,N_8522,N_8451);
nor U8691 (N_8691,N_8412,N_8519);
or U8692 (N_8692,N_8510,N_8431);
and U8693 (N_8693,N_8583,N_8470);
nand U8694 (N_8694,N_8440,N_8571);
nand U8695 (N_8695,N_8498,N_8409);
nand U8696 (N_8696,N_8541,N_8570);
or U8697 (N_8697,N_8546,N_8485);
and U8698 (N_8698,N_8542,N_8401);
or U8699 (N_8699,N_8524,N_8593);
and U8700 (N_8700,N_8537,N_8458);
and U8701 (N_8701,N_8497,N_8448);
and U8702 (N_8702,N_8572,N_8543);
or U8703 (N_8703,N_8537,N_8588);
nand U8704 (N_8704,N_8438,N_8538);
nand U8705 (N_8705,N_8445,N_8443);
nand U8706 (N_8706,N_8574,N_8517);
nor U8707 (N_8707,N_8420,N_8567);
nor U8708 (N_8708,N_8549,N_8529);
nand U8709 (N_8709,N_8593,N_8498);
and U8710 (N_8710,N_8411,N_8457);
or U8711 (N_8711,N_8401,N_8450);
nor U8712 (N_8712,N_8588,N_8541);
nand U8713 (N_8713,N_8461,N_8450);
or U8714 (N_8714,N_8429,N_8457);
or U8715 (N_8715,N_8505,N_8499);
and U8716 (N_8716,N_8497,N_8482);
nor U8717 (N_8717,N_8483,N_8442);
nor U8718 (N_8718,N_8452,N_8596);
and U8719 (N_8719,N_8423,N_8454);
or U8720 (N_8720,N_8444,N_8499);
nor U8721 (N_8721,N_8441,N_8438);
and U8722 (N_8722,N_8410,N_8579);
nand U8723 (N_8723,N_8480,N_8549);
nor U8724 (N_8724,N_8480,N_8564);
or U8725 (N_8725,N_8422,N_8455);
or U8726 (N_8726,N_8580,N_8579);
or U8727 (N_8727,N_8400,N_8420);
nand U8728 (N_8728,N_8414,N_8485);
nor U8729 (N_8729,N_8501,N_8594);
nor U8730 (N_8730,N_8562,N_8555);
nor U8731 (N_8731,N_8549,N_8583);
nand U8732 (N_8732,N_8558,N_8469);
nand U8733 (N_8733,N_8432,N_8558);
nand U8734 (N_8734,N_8472,N_8526);
and U8735 (N_8735,N_8447,N_8594);
and U8736 (N_8736,N_8496,N_8560);
or U8737 (N_8737,N_8524,N_8460);
nor U8738 (N_8738,N_8465,N_8571);
nand U8739 (N_8739,N_8572,N_8490);
and U8740 (N_8740,N_8460,N_8526);
or U8741 (N_8741,N_8444,N_8575);
and U8742 (N_8742,N_8499,N_8562);
nor U8743 (N_8743,N_8428,N_8486);
nand U8744 (N_8744,N_8585,N_8575);
nand U8745 (N_8745,N_8527,N_8518);
and U8746 (N_8746,N_8515,N_8503);
and U8747 (N_8747,N_8500,N_8564);
or U8748 (N_8748,N_8498,N_8490);
and U8749 (N_8749,N_8446,N_8595);
nor U8750 (N_8750,N_8430,N_8547);
nor U8751 (N_8751,N_8519,N_8597);
or U8752 (N_8752,N_8450,N_8419);
and U8753 (N_8753,N_8428,N_8497);
or U8754 (N_8754,N_8487,N_8433);
nor U8755 (N_8755,N_8597,N_8442);
or U8756 (N_8756,N_8480,N_8547);
nor U8757 (N_8757,N_8419,N_8485);
and U8758 (N_8758,N_8429,N_8423);
nor U8759 (N_8759,N_8456,N_8524);
nor U8760 (N_8760,N_8517,N_8449);
nand U8761 (N_8761,N_8442,N_8535);
nor U8762 (N_8762,N_8481,N_8553);
nand U8763 (N_8763,N_8527,N_8498);
and U8764 (N_8764,N_8563,N_8508);
and U8765 (N_8765,N_8562,N_8470);
nor U8766 (N_8766,N_8587,N_8517);
and U8767 (N_8767,N_8474,N_8524);
nand U8768 (N_8768,N_8491,N_8561);
or U8769 (N_8769,N_8595,N_8559);
or U8770 (N_8770,N_8467,N_8571);
or U8771 (N_8771,N_8581,N_8580);
xor U8772 (N_8772,N_8407,N_8451);
nor U8773 (N_8773,N_8407,N_8541);
and U8774 (N_8774,N_8408,N_8409);
and U8775 (N_8775,N_8401,N_8549);
or U8776 (N_8776,N_8580,N_8588);
and U8777 (N_8777,N_8587,N_8573);
nor U8778 (N_8778,N_8441,N_8516);
or U8779 (N_8779,N_8423,N_8586);
nand U8780 (N_8780,N_8532,N_8589);
and U8781 (N_8781,N_8595,N_8581);
nor U8782 (N_8782,N_8496,N_8434);
nor U8783 (N_8783,N_8526,N_8468);
or U8784 (N_8784,N_8427,N_8431);
or U8785 (N_8785,N_8593,N_8448);
nand U8786 (N_8786,N_8520,N_8482);
and U8787 (N_8787,N_8492,N_8491);
and U8788 (N_8788,N_8493,N_8536);
nand U8789 (N_8789,N_8471,N_8505);
nor U8790 (N_8790,N_8493,N_8526);
or U8791 (N_8791,N_8594,N_8584);
and U8792 (N_8792,N_8586,N_8499);
nor U8793 (N_8793,N_8562,N_8446);
and U8794 (N_8794,N_8438,N_8463);
nor U8795 (N_8795,N_8484,N_8477);
nand U8796 (N_8796,N_8518,N_8588);
and U8797 (N_8797,N_8559,N_8592);
or U8798 (N_8798,N_8437,N_8521);
nor U8799 (N_8799,N_8484,N_8521);
nor U8800 (N_8800,N_8623,N_8695);
nand U8801 (N_8801,N_8659,N_8674);
nand U8802 (N_8802,N_8709,N_8795);
nor U8803 (N_8803,N_8693,N_8756);
nor U8804 (N_8804,N_8616,N_8730);
or U8805 (N_8805,N_8612,N_8654);
or U8806 (N_8806,N_8707,N_8712);
and U8807 (N_8807,N_8717,N_8656);
nor U8808 (N_8808,N_8648,N_8711);
or U8809 (N_8809,N_8615,N_8749);
or U8810 (N_8810,N_8607,N_8672);
nor U8811 (N_8811,N_8742,N_8755);
nand U8812 (N_8812,N_8671,N_8767);
nand U8813 (N_8813,N_8690,N_8737);
xnor U8814 (N_8814,N_8724,N_8747);
and U8815 (N_8815,N_8633,N_8748);
nor U8816 (N_8816,N_8618,N_8630);
or U8817 (N_8817,N_8669,N_8641);
or U8818 (N_8818,N_8699,N_8744);
nand U8819 (N_8819,N_8774,N_8652);
and U8820 (N_8820,N_8664,N_8777);
and U8821 (N_8821,N_8610,N_8752);
nand U8822 (N_8822,N_8697,N_8673);
nor U8823 (N_8823,N_8644,N_8703);
or U8824 (N_8824,N_8613,N_8708);
nand U8825 (N_8825,N_8791,N_8725);
nand U8826 (N_8826,N_8772,N_8685);
or U8827 (N_8827,N_8776,N_8735);
nor U8828 (N_8828,N_8705,N_8625);
nand U8829 (N_8829,N_8770,N_8682);
or U8830 (N_8830,N_8784,N_8793);
nor U8831 (N_8831,N_8720,N_8646);
or U8832 (N_8832,N_8786,N_8734);
nor U8833 (N_8833,N_8759,N_8754);
nand U8834 (N_8834,N_8726,N_8773);
and U8835 (N_8835,N_8740,N_8617);
nor U8836 (N_8836,N_8691,N_8728);
nand U8837 (N_8837,N_8614,N_8663);
and U8838 (N_8838,N_8796,N_8713);
and U8839 (N_8839,N_8788,N_8622);
or U8840 (N_8840,N_8653,N_8736);
nand U8841 (N_8841,N_8718,N_8769);
nor U8842 (N_8842,N_8761,N_8743);
or U8843 (N_8843,N_8687,N_8620);
nor U8844 (N_8844,N_8739,N_8775);
and U8845 (N_8845,N_8636,N_8643);
nand U8846 (N_8846,N_8624,N_8781);
nand U8847 (N_8847,N_8689,N_8765);
nand U8848 (N_8848,N_8619,N_8745);
and U8849 (N_8849,N_8670,N_8727);
nor U8850 (N_8850,N_8721,N_8602);
nor U8851 (N_8851,N_8797,N_8680);
nand U8852 (N_8852,N_8655,N_8760);
or U8853 (N_8853,N_8683,N_8686);
or U8854 (N_8854,N_8787,N_8746);
and U8855 (N_8855,N_8783,N_8668);
nand U8856 (N_8856,N_8764,N_8660);
nor U8857 (N_8857,N_8782,N_8661);
and U8858 (N_8858,N_8738,N_8722);
nor U8859 (N_8859,N_8716,N_8635);
nand U8860 (N_8860,N_8799,N_8688);
or U8861 (N_8861,N_8601,N_8676);
nor U8862 (N_8862,N_8640,N_8649);
and U8863 (N_8863,N_8753,N_8665);
nor U8864 (N_8864,N_8667,N_8758);
nand U8865 (N_8865,N_8605,N_8651);
nor U8866 (N_8866,N_8666,N_8762);
nand U8867 (N_8867,N_8627,N_8692);
or U8868 (N_8868,N_8751,N_8710);
nand U8869 (N_8869,N_8662,N_8731);
or U8870 (N_8870,N_8647,N_8609);
nand U8871 (N_8871,N_8629,N_8696);
and U8872 (N_8872,N_8790,N_8768);
or U8873 (N_8873,N_8681,N_8637);
or U8874 (N_8874,N_8789,N_8657);
and U8875 (N_8875,N_8785,N_8704);
or U8876 (N_8876,N_8732,N_8714);
or U8877 (N_8877,N_8715,N_8634);
nand U8878 (N_8878,N_8611,N_8679);
nand U8879 (N_8879,N_8706,N_8658);
or U8880 (N_8880,N_8639,N_8779);
and U8881 (N_8881,N_8600,N_8763);
nand U8882 (N_8882,N_8642,N_8792);
and U8883 (N_8883,N_8645,N_8694);
nand U8884 (N_8884,N_8794,N_8698);
nor U8885 (N_8885,N_8604,N_8723);
nor U8886 (N_8886,N_8608,N_8606);
nor U8887 (N_8887,N_8632,N_8701);
or U8888 (N_8888,N_8702,N_8766);
or U8889 (N_8889,N_8628,N_8733);
or U8890 (N_8890,N_8741,N_8798);
and U8891 (N_8891,N_8678,N_8778);
and U8892 (N_8892,N_8626,N_8621);
and U8893 (N_8893,N_8729,N_8684);
nor U8894 (N_8894,N_8677,N_8757);
nand U8895 (N_8895,N_8780,N_8675);
or U8896 (N_8896,N_8750,N_8603);
or U8897 (N_8897,N_8650,N_8771);
nand U8898 (N_8898,N_8631,N_8638);
nor U8899 (N_8899,N_8719,N_8700);
nor U8900 (N_8900,N_8665,N_8639);
and U8901 (N_8901,N_8651,N_8642);
and U8902 (N_8902,N_8712,N_8768);
nand U8903 (N_8903,N_8632,N_8786);
nor U8904 (N_8904,N_8691,N_8696);
nor U8905 (N_8905,N_8720,N_8763);
nand U8906 (N_8906,N_8794,N_8710);
nand U8907 (N_8907,N_8760,N_8610);
and U8908 (N_8908,N_8782,N_8702);
or U8909 (N_8909,N_8710,N_8789);
nor U8910 (N_8910,N_8705,N_8748);
and U8911 (N_8911,N_8691,N_8693);
nor U8912 (N_8912,N_8637,N_8668);
or U8913 (N_8913,N_8706,N_8714);
or U8914 (N_8914,N_8671,N_8633);
nand U8915 (N_8915,N_8646,N_8750);
and U8916 (N_8916,N_8727,N_8711);
nand U8917 (N_8917,N_8795,N_8688);
nor U8918 (N_8918,N_8641,N_8714);
nand U8919 (N_8919,N_8600,N_8646);
nand U8920 (N_8920,N_8725,N_8788);
or U8921 (N_8921,N_8749,N_8757);
or U8922 (N_8922,N_8717,N_8712);
and U8923 (N_8923,N_8725,N_8692);
xnor U8924 (N_8924,N_8745,N_8695);
or U8925 (N_8925,N_8720,N_8619);
or U8926 (N_8926,N_8690,N_8652);
or U8927 (N_8927,N_8622,N_8777);
or U8928 (N_8928,N_8676,N_8696);
nor U8929 (N_8929,N_8657,N_8648);
nand U8930 (N_8930,N_8681,N_8779);
xor U8931 (N_8931,N_8794,N_8607);
or U8932 (N_8932,N_8791,N_8715);
and U8933 (N_8933,N_8693,N_8618);
and U8934 (N_8934,N_8662,N_8738);
or U8935 (N_8935,N_8760,N_8651);
nand U8936 (N_8936,N_8603,N_8782);
and U8937 (N_8937,N_8705,N_8613);
nand U8938 (N_8938,N_8680,N_8758);
nand U8939 (N_8939,N_8720,N_8786);
or U8940 (N_8940,N_8611,N_8603);
nand U8941 (N_8941,N_8619,N_8649);
and U8942 (N_8942,N_8737,N_8710);
nor U8943 (N_8943,N_8703,N_8663);
nand U8944 (N_8944,N_8712,N_8704);
nand U8945 (N_8945,N_8620,N_8615);
and U8946 (N_8946,N_8607,N_8670);
nor U8947 (N_8947,N_8739,N_8768);
nand U8948 (N_8948,N_8624,N_8656);
or U8949 (N_8949,N_8685,N_8780);
or U8950 (N_8950,N_8714,N_8696);
nand U8951 (N_8951,N_8619,N_8796);
and U8952 (N_8952,N_8764,N_8784);
nor U8953 (N_8953,N_8715,N_8784);
nand U8954 (N_8954,N_8763,N_8619);
nor U8955 (N_8955,N_8707,N_8666);
or U8956 (N_8956,N_8693,N_8666);
nor U8957 (N_8957,N_8709,N_8746);
or U8958 (N_8958,N_8748,N_8615);
and U8959 (N_8959,N_8668,N_8686);
or U8960 (N_8960,N_8665,N_8798);
or U8961 (N_8961,N_8754,N_8762);
nand U8962 (N_8962,N_8608,N_8682);
or U8963 (N_8963,N_8727,N_8757);
nor U8964 (N_8964,N_8788,N_8742);
nand U8965 (N_8965,N_8608,N_8693);
nor U8966 (N_8966,N_8623,N_8619);
nor U8967 (N_8967,N_8779,N_8608);
or U8968 (N_8968,N_8710,N_8774);
and U8969 (N_8969,N_8706,N_8650);
and U8970 (N_8970,N_8655,N_8603);
or U8971 (N_8971,N_8694,N_8735);
or U8972 (N_8972,N_8684,N_8672);
nand U8973 (N_8973,N_8786,N_8784);
or U8974 (N_8974,N_8760,N_8733);
nor U8975 (N_8975,N_8607,N_8779);
and U8976 (N_8976,N_8708,N_8727);
nand U8977 (N_8977,N_8648,N_8781);
nor U8978 (N_8978,N_8761,N_8610);
or U8979 (N_8979,N_8796,N_8762);
nand U8980 (N_8980,N_8621,N_8692);
and U8981 (N_8981,N_8754,N_8771);
nor U8982 (N_8982,N_8648,N_8675);
nand U8983 (N_8983,N_8665,N_8768);
nor U8984 (N_8984,N_8696,N_8757);
xnor U8985 (N_8985,N_8611,N_8785);
nor U8986 (N_8986,N_8676,N_8728);
and U8987 (N_8987,N_8645,N_8665);
nand U8988 (N_8988,N_8786,N_8767);
and U8989 (N_8989,N_8641,N_8634);
or U8990 (N_8990,N_8659,N_8741);
nand U8991 (N_8991,N_8710,N_8744);
nor U8992 (N_8992,N_8764,N_8738);
or U8993 (N_8993,N_8778,N_8687);
and U8994 (N_8994,N_8644,N_8603);
nor U8995 (N_8995,N_8778,N_8677);
nand U8996 (N_8996,N_8706,N_8620);
nor U8997 (N_8997,N_8793,N_8667);
nand U8998 (N_8998,N_8734,N_8649);
nand U8999 (N_8999,N_8630,N_8648);
and U9000 (N_9000,N_8872,N_8898);
nand U9001 (N_9001,N_8943,N_8950);
or U9002 (N_9002,N_8836,N_8972);
nand U9003 (N_9003,N_8983,N_8881);
nand U9004 (N_9004,N_8861,N_8859);
or U9005 (N_9005,N_8833,N_8849);
or U9006 (N_9006,N_8944,N_8933);
nor U9007 (N_9007,N_8902,N_8949);
nand U9008 (N_9008,N_8989,N_8886);
nor U9009 (N_9009,N_8918,N_8807);
or U9010 (N_9010,N_8848,N_8904);
or U9011 (N_9011,N_8862,N_8815);
and U9012 (N_9012,N_8830,N_8938);
nand U9013 (N_9013,N_8941,N_8867);
and U9014 (N_9014,N_8915,N_8877);
nor U9015 (N_9015,N_8884,N_8976);
nor U9016 (N_9016,N_8926,N_8817);
nor U9017 (N_9017,N_8835,N_8810);
nor U9018 (N_9018,N_8963,N_8857);
nand U9019 (N_9019,N_8843,N_8945);
nand U9020 (N_9020,N_8931,N_8865);
nand U9021 (N_9021,N_8912,N_8992);
and U9022 (N_9022,N_8828,N_8984);
and U9023 (N_9023,N_8850,N_8934);
nor U9024 (N_9024,N_8812,N_8970);
nand U9025 (N_9025,N_8855,N_8973);
and U9026 (N_9026,N_8840,N_8889);
or U9027 (N_9027,N_8883,N_8996);
nor U9028 (N_9028,N_8925,N_8837);
or U9029 (N_9029,N_8927,N_8910);
and U9030 (N_9030,N_8977,N_8980);
nand U9031 (N_9031,N_8894,N_8824);
or U9032 (N_9032,N_8986,N_8863);
nor U9033 (N_9033,N_8952,N_8826);
or U9034 (N_9034,N_8900,N_8831);
nor U9035 (N_9035,N_8960,N_8813);
or U9036 (N_9036,N_8935,N_8821);
or U9037 (N_9037,N_8866,N_8800);
and U9038 (N_9038,N_8806,N_8921);
nor U9039 (N_9039,N_8899,N_8887);
or U9040 (N_9040,N_8852,N_8804);
or U9041 (N_9041,N_8802,N_8805);
and U9042 (N_9042,N_8868,N_8879);
or U9043 (N_9043,N_8873,N_8864);
nand U9044 (N_9044,N_8909,N_8966);
nor U9045 (N_9045,N_8911,N_8839);
or U9046 (N_9046,N_8814,N_8841);
nor U9047 (N_9047,N_8954,N_8961);
and U9048 (N_9048,N_8946,N_8939);
and U9049 (N_9049,N_8834,N_8892);
and U9050 (N_9050,N_8875,N_8844);
nor U9051 (N_9051,N_8846,N_8908);
and U9052 (N_9052,N_8885,N_8975);
or U9053 (N_9053,N_8968,N_8985);
and U9054 (N_9054,N_8922,N_8890);
or U9055 (N_9055,N_8818,N_8832);
nand U9056 (N_9056,N_8823,N_8953);
nand U9057 (N_9057,N_8993,N_8988);
and U9058 (N_9058,N_8854,N_8947);
and U9059 (N_9059,N_8842,N_8856);
and U9060 (N_9060,N_8891,N_8995);
and U9061 (N_9061,N_8959,N_8917);
nand U9062 (N_9062,N_8858,N_8907);
or U9063 (N_9063,N_8870,N_8990);
and U9064 (N_9064,N_8853,N_8999);
xor U9065 (N_9065,N_8940,N_8895);
and U9066 (N_9066,N_8974,N_8882);
and U9067 (N_9067,N_8829,N_8903);
nor U9068 (N_9068,N_8978,N_8965);
nand U9069 (N_9069,N_8820,N_8956);
or U9070 (N_9070,N_8811,N_8860);
or U9071 (N_9071,N_8878,N_8967);
or U9072 (N_9072,N_8951,N_8809);
and U9073 (N_9073,N_8964,N_8801);
and U9074 (N_9074,N_8876,N_8957);
nor U9075 (N_9075,N_8979,N_8913);
nor U9076 (N_9076,N_8825,N_8920);
nor U9077 (N_9077,N_8803,N_8948);
nor U9078 (N_9078,N_8888,N_8924);
and U9079 (N_9079,N_8822,N_8919);
or U9080 (N_9080,N_8982,N_8981);
and U9081 (N_9081,N_8962,N_8914);
nor U9082 (N_9082,N_8906,N_8893);
and U9083 (N_9083,N_8997,N_8871);
nand U9084 (N_9084,N_8880,N_8958);
nand U9085 (N_9085,N_8897,N_8955);
nor U9086 (N_9086,N_8905,N_8896);
and U9087 (N_9087,N_8816,N_8847);
nand U9088 (N_9088,N_8987,N_8928);
nand U9089 (N_9089,N_8923,N_8930);
and U9090 (N_9090,N_8937,N_8851);
and U9091 (N_9091,N_8838,N_8808);
and U9092 (N_9092,N_8969,N_8901);
or U9093 (N_9093,N_8942,N_8936);
and U9094 (N_9094,N_8874,N_8916);
nor U9095 (N_9095,N_8971,N_8994);
or U9096 (N_9096,N_8819,N_8998);
or U9097 (N_9097,N_8827,N_8929);
and U9098 (N_9098,N_8932,N_8845);
or U9099 (N_9099,N_8991,N_8869);
and U9100 (N_9100,N_8846,N_8921);
and U9101 (N_9101,N_8869,N_8940);
nor U9102 (N_9102,N_8933,N_8989);
or U9103 (N_9103,N_8846,N_8958);
nand U9104 (N_9104,N_8858,N_8886);
nand U9105 (N_9105,N_8861,N_8936);
nor U9106 (N_9106,N_8998,N_8834);
and U9107 (N_9107,N_8827,N_8988);
nand U9108 (N_9108,N_8910,N_8979);
or U9109 (N_9109,N_8843,N_8935);
and U9110 (N_9110,N_8945,N_8998);
or U9111 (N_9111,N_8823,N_8962);
nor U9112 (N_9112,N_8825,N_8966);
and U9113 (N_9113,N_8871,N_8969);
nor U9114 (N_9114,N_8928,N_8829);
or U9115 (N_9115,N_8840,N_8805);
or U9116 (N_9116,N_8852,N_8854);
nor U9117 (N_9117,N_8979,N_8987);
nor U9118 (N_9118,N_8953,N_8982);
and U9119 (N_9119,N_8873,N_8943);
and U9120 (N_9120,N_8858,N_8807);
nand U9121 (N_9121,N_8989,N_8826);
and U9122 (N_9122,N_8993,N_8833);
or U9123 (N_9123,N_8929,N_8887);
or U9124 (N_9124,N_8951,N_8949);
nor U9125 (N_9125,N_8962,N_8970);
nor U9126 (N_9126,N_8932,N_8859);
nand U9127 (N_9127,N_8896,N_8834);
or U9128 (N_9128,N_8844,N_8952);
nand U9129 (N_9129,N_8995,N_8960);
and U9130 (N_9130,N_8959,N_8906);
nand U9131 (N_9131,N_8880,N_8803);
nand U9132 (N_9132,N_8879,N_8839);
or U9133 (N_9133,N_8917,N_8876);
and U9134 (N_9134,N_8882,N_8844);
nor U9135 (N_9135,N_8834,N_8804);
nand U9136 (N_9136,N_8976,N_8926);
and U9137 (N_9137,N_8853,N_8861);
nor U9138 (N_9138,N_8832,N_8878);
and U9139 (N_9139,N_8889,N_8937);
or U9140 (N_9140,N_8995,N_8881);
and U9141 (N_9141,N_8898,N_8908);
and U9142 (N_9142,N_8896,N_8850);
and U9143 (N_9143,N_8943,N_8886);
nor U9144 (N_9144,N_8809,N_8921);
and U9145 (N_9145,N_8860,N_8901);
nor U9146 (N_9146,N_8974,N_8924);
and U9147 (N_9147,N_8899,N_8848);
or U9148 (N_9148,N_8868,N_8946);
nor U9149 (N_9149,N_8955,N_8936);
and U9150 (N_9150,N_8871,N_8971);
and U9151 (N_9151,N_8964,N_8834);
nand U9152 (N_9152,N_8834,N_8830);
and U9153 (N_9153,N_8830,N_8825);
and U9154 (N_9154,N_8806,N_8847);
nand U9155 (N_9155,N_8866,N_8811);
or U9156 (N_9156,N_8840,N_8968);
nor U9157 (N_9157,N_8938,N_8956);
nand U9158 (N_9158,N_8941,N_8972);
nand U9159 (N_9159,N_8846,N_8967);
and U9160 (N_9160,N_8886,N_8808);
and U9161 (N_9161,N_8916,N_8838);
nand U9162 (N_9162,N_8968,N_8901);
or U9163 (N_9163,N_8981,N_8866);
nand U9164 (N_9164,N_8921,N_8948);
and U9165 (N_9165,N_8927,N_8999);
nor U9166 (N_9166,N_8872,N_8920);
or U9167 (N_9167,N_8880,N_8940);
and U9168 (N_9168,N_8992,N_8898);
nor U9169 (N_9169,N_8998,N_8986);
nor U9170 (N_9170,N_8860,N_8879);
nor U9171 (N_9171,N_8857,N_8854);
and U9172 (N_9172,N_8938,N_8972);
nand U9173 (N_9173,N_8803,N_8960);
nand U9174 (N_9174,N_8903,N_8848);
or U9175 (N_9175,N_8957,N_8964);
nor U9176 (N_9176,N_8861,N_8883);
and U9177 (N_9177,N_8901,N_8850);
and U9178 (N_9178,N_8860,N_8817);
nand U9179 (N_9179,N_8886,N_8890);
nor U9180 (N_9180,N_8946,N_8835);
and U9181 (N_9181,N_8802,N_8844);
and U9182 (N_9182,N_8809,N_8862);
nor U9183 (N_9183,N_8959,N_8854);
nor U9184 (N_9184,N_8810,N_8868);
and U9185 (N_9185,N_8814,N_8862);
nor U9186 (N_9186,N_8832,N_8819);
and U9187 (N_9187,N_8818,N_8811);
or U9188 (N_9188,N_8833,N_8966);
or U9189 (N_9189,N_8887,N_8990);
or U9190 (N_9190,N_8906,N_8922);
nand U9191 (N_9191,N_8806,N_8992);
nand U9192 (N_9192,N_8988,N_8828);
nor U9193 (N_9193,N_8878,N_8906);
nor U9194 (N_9194,N_8841,N_8953);
or U9195 (N_9195,N_8949,N_8977);
nand U9196 (N_9196,N_8978,N_8990);
or U9197 (N_9197,N_8845,N_8936);
nand U9198 (N_9198,N_8862,N_8928);
nor U9199 (N_9199,N_8869,N_8879);
and U9200 (N_9200,N_9172,N_9137);
and U9201 (N_9201,N_9042,N_9190);
or U9202 (N_9202,N_9009,N_9171);
nor U9203 (N_9203,N_9158,N_9151);
nor U9204 (N_9204,N_9110,N_9125);
nor U9205 (N_9205,N_9085,N_9186);
and U9206 (N_9206,N_9078,N_9038);
or U9207 (N_9207,N_9057,N_9103);
nor U9208 (N_9208,N_9126,N_9083);
or U9209 (N_9209,N_9066,N_9022);
and U9210 (N_9210,N_9161,N_9142);
or U9211 (N_9211,N_9132,N_9153);
and U9212 (N_9212,N_9055,N_9024);
and U9213 (N_9213,N_9069,N_9053);
and U9214 (N_9214,N_9101,N_9168);
and U9215 (N_9215,N_9154,N_9033);
nand U9216 (N_9216,N_9164,N_9105);
or U9217 (N_9217,N_9084,N_9138);
nor U9218 (N_9218,N_9188,N_9109);
or U9219 (N_9219,N_9170,N_9149);
and U9220 (N_9220,N_9124,N_9061);
nor U9221 (N_9221,N_9043,N_9015);
and U9222 (N_9222,N_9178,N_9064);
or U9223 (N_9223,N_9058,N_9095);
nor U9224 (N_9224,N_9060,N_9011);
nand U9225 (N_9225,N_9037,N_9191);
or U9226 (N_9226,N_9004,N_9006);
and U9227 (N_9227,N_9116,N_9050);
and U9228 (N_9228,N_9147,N_9123);
nand U9229 (N_9229,N_9150,N_9143);
nand U9230 (N_9230,N_9096,N_9081);
nand U9231 (N_9231,N_9065,N_9157);
nor U9232 (N_9232,N_9062,N_9160);
nor U9233 (N_9233,N_9165,N_9148);
xnor U9234 (N_9234,N_9187,N_9045);
and U9235 (N_9235,N_9029,N_9021);
nand U9236 (N_9236,N_9005,N_9199);
nor U9237 (N_9237,N_9087,N_9007);
and U9238 (N_9238,N_9012,N_9048);
or U9239 (N_9239,N_9195,N_9008);
nand U9240 (N_9240,N_9102,N_9185);
and U9241 (N_9241,N_9175,N_9093);
nand U9242 (N_9242,N_9121,N_9119);
or U9243 (N_9243,N_9063,N_9054);
and U9244 (N_9244,N_9040,N_9117);
and U9245 (N_9245,N_9014,N_9086);
nor U9246 (N_9246,N_9136,N_9155);
and U9247 (N_9247,N_9193,N_9047);
and U9248 (N_9248,N_9099,N_9166);
and U9249 (N_9249,N_9162,N_9002);
and U9250 (N_9250,N_9189,N_9156);
nor U9251 (N_9251,N_9131,N_9122);
and U9252 (N_9252,N_9044,N_9074);
and U9253 (N_9253,N_9183,N_9113);
nand U9254 (N_9254,N_9134,N_9039);
nand U9255 (N_9255,N_9091,N_9067);
nand U9256 (N_9256,N_9127,N_9115);
nand U9257 (N_9257,N_9144,N_9167);
and U9258 (N_9258,N_9010,N_9090);
or U9259 (N_9259,N_9194,N_9097);
nand U9260 (N_9260,N_9088,N_9013);
nor U9261 (N_9261,N_9094,N_9025);
nand U9262 (N_9262,N_9071,N_9114);
nor U9263 (N_9263,N_9129,N_9003);
or U9264 (N_9264,N_9177,N_9020);
and U9265 (N_9265,N_9089,N_9184);
nor U9266 (N_9266,N_9041,N_9016);
nor U9267 (N_9267,N_9035,N_9070);
and U9268 (N_9268,N_9111,N_9192);
nand U9269 (N_9269,N_9076,N_9174);
nor U9270 (N_9270,N_9073,N_9028);
or U9271 (N_9271,N_9072,N_9169);
nand U9272 (N_9272,N_9163,N_9128);
nand U9273 (N_9273,N_9026,N_9106);
nor U9274 (N_9274,N_9180,N_9052);
and U9275 (N_9275,N_9118,N_9141);
or U9276 (N_9276,N_9140,N_9017);
nor U9277 (N_9277,N_9098,N_9159);
nor U9278 (N_9278,N_9056,N_9100);
nor U9279 (N_9279,N_9032,N_9000);
nand U9280 (N_9280,N_9176,N_9051);
nor U9281 (N_9281,N_9068,N_9107);
or U9282 (N_9282,N_9059,N_9198);
or U9283 (N_9283,N_9120,N_9197);
nor U9284 (N_9284,N_9079,N_9077);
nor U9285 (N_9285,N_9075,N_9046);
nor U9286 (N_9286,N_9182,N_9108);
or U9287 (N_9287,N_9133,N_9018);
nand U9288 (N_9288,N_9179,N_9130);
and U9289 (N_9289,N_9023,N_9036);
and U9290 (N_9290,N_9145,N_9082);
or U9291 (N_9291,N_9139,N_9031);
nor U9292 (N_9292,N_9092,N_9034);
nand U9293 (N_9293,N_9135,N_9001);
or U9294 (N_9294,N_9104,N_9049);
or U9295 (N_9295,N_9146,N_9173);
or U9296 (N_9296,N_9027,N_9019);
nor U9297 (N_9297,N_9152,N_9030);
nor U9298 (N_9298,N_9196,N_9080);
and U9299 (N_9299,N_9181,N_9112);
and U9300 (N_9300,N_9123,N_9148);
nor U9301 (N_9301,N_9196,N_9070);
and U9302 (N_9302,N_9169,N_9091);
nor U9303 (N_9303,N_9091,N_9009);
and U9304 (N_9304,N_9134,N_9113);
nand U9305 (N_9305,N_9177,N_9066);
nand U9306 (N_9306,N_9089,N_9096);
or U9307 (N_9307,N_9095,N_9021);
and U9308 (N_9308,N_9139,N_9173);
nor U9309 (N_9309,N_9169,N_9064);
or U9310 (N_9310,N_9091,N_9117);
or U9311 (N_9311,N_9136,N_9104);
and U9312 (N_9312,N_9177,N_9144);
or U9313 (N_9313,N_9111,N_9061);
nand U9314 (N_9314,N_9076,N_9049);
or U9315 (N_9315,N_9156,N_9155);
and U9316 (N_9316,N_9148,N_9087);
nor U9317 (N_9317,N_9010,N_9156);
and U9318 (N_9318,N_9052,N_9190);
or U9319 (N_9319,N_9197,N_9025);
and U9320 (N_9320,N_9105,N_9006);
nor U9321 (N_9321,N_9090,N_9106);
nand U9322 (N_9322,N_9197,N_9138);
nand U9323 (N_9323,N_9023,N_9192);
nand U9324 (N_9324,N_9016,N_9071);
nor U9325 (N_9325,N_9078,N_9177);
or U9326 (N_9326,N_9007,N_9035);
or U9327 (N_9327,N_9193,N_9044);
or U9328 (N_9328,N_9044,N_9115);
or U9329 (N_9329,N_9047,N_9045);
nor U9330 (N_9330,N_9149,N_9185);
or U9331 (N_9331,N_9066,N_9191);
nand U9332 (N_9332,N_9038,N_9149);
or U9333 (N_9333,N_9170,N_9061);
and U9334 (N_9334,N_9083,N_9133);
nor U9335 (N_9335,N_9137,N_9010);
and U9336 (N_9336,N_9124,N_9074);
nor U9337 (N_9337,N_9018,N_9102);
or U9338 (N_9338,N_9055,N_9073);
nand U9339 (N_9339,N_9198,N_9025);
nor U9340 (N_9340,N_9149,N_9053);
or U9341 (N_9341,N_9022,N_9014);
and U9342 (N_9342,N_9028,N_9159);
and U9343 (N_9343,N_9198,N_9175);
nand U9344 (N_9344,N_9028,N_9099);
and U9345 (N_9345,N_9070,N_9046);
or U9346 (N_9346,N_9172,N_9031);
xor U9347 (N_9347,N_9156,N_9185);
or U9348 (N_9348,N_9026,N_9048);
or U9349 (N_9349,N_9071,N_9028);
nand U9350 (N_9350,N_9094,N_9053);
nor U9351 (N_9351,N_9066,N_9081);
nor U9352 (N_9352,N_9090,N_9053);
nor U9353 (N_9353,N_9017,N_9176);
nor U9354 (N_9354,N_9168,N_9199);
nor U9355 (N_9355,N_9192,N_9056);
or U9356 (N_9356,N_9025,N_9017);
and U9357 (N_9357,N_9162,N_9130);
and U9358 (N_9358,N_9018,N_9010);
or U9359 (N_9359,N_9055,N_9080);
nor U9360 (N_9360,N_9091,N_9141);
nor U9361 (N_9361,N_9095,N_9172);
and U9362 (N_9362,N_9073,N_9170);
and U9363 (N_9363,N_9185,N_9000);
nand U9364 (N_9364,N_9112,N_9163);
nor U9365 (N_9365,N_9098,N_9023);
and U9366 (N_9366,N_9165,N_9029);
or U9367 (N_9367,N_9082,N_9064);
nor U9368 (N_9368,N_9153,N_9026);
and U9369 (N_9369,N_9075,N_9083);
nor U9370 (N_9370,N_9137,N_9002);
and U9371 (N_9371,N_9115,N_9185);
nand U9372 (N_9372,N_9102,N_9045);
or U9373 (N_9373,N_9098,N_9119);
or U9374 (N_9374,N_9100,N_9165);
or U9375 (N_9375,N_9166,N_9085);
or U9376 (N_9376,N_9164,N_9096);
or U9377 (N_9377,N_9052,N_9193);
nand U9378 (N_9378,N_9046,N_9154);
nor U9379 (N_9379,N_9133,N_9115);
nor U9380 (N_9380,N_9176,N_9056);
xor U9381 (N_9381,N_9038,N_9138);
or U9382 (N_9382,N_9170,N_9006);
nand U9383 (N_9383,N_9172,N_9143);
nand U9384 (N_9384,N_9108,N_9043);
nand U9385 (N_9385,N_9198,N_9052);
or U9386 (N_9386,N_9024,N_9082);
and U9387 (N_9387,N_9148,N_9073);
or U9388 (N_9388,N_9028,N_9108);
xnor U9389 (N_9389,N_9009,N_9001);
or U9390 (N_9390,N_9008,N_9052);
or U9391 (N_9391,N_9100,N_9017);
or U9392 (N_9392,N_9036,N_9073);
and U9393 (N_9393,N_9019,N_9169);
and U9394 (N_9394,N_9009,N_9000);
nor U9395 (N_9395,N_9098,N_9068);
and U9396 (N_9396,N_9171,N_9155);
or U9397 (N_9397,N_9158,N_9062);
nand U9398 (N_9398,N_9078,N_9048);
or U9399 (N_9399,N_9117,N_9197);
nor U9400 (N_9400,N_9284,N_9247);
or U9401 (N_9401,N_9250,N_9218);
nand U9402 (N_9402,N_9384,N_9206);
and U9403 (N_9403,N_9388,N_9300);
nand U9404 (N_9404,N_9338,N_9246);
and U9405 (N_9405,N_9291,N_9251);
or U9406 (N_9406,N_9396,N_9318);
or U9407 (N_9407,N_9343,N_9326);
or U9408 (N_9408,N_9356,N_9216);
and U9409 (N_9409,N_9233,N_9288);
and U9410 (N_9410,N_9319,N_9378);
or U9411 (N_9411,N_9289,N_9221);
or U9412 (N_9412,N_9264,N_9217);
and U9413 (N_9413,N_9276,N_9249);
nand U9414 (N_9414,N_9298,N_9339);
nor U9415 (N_9415,N_9342,N_9364);
and U9416 (N_9416,N_9210,N_9259);
and U9417 (N_9417,N_9395,N_9215);
nand U9418 (N_9418,N_9279,N_9253);
nor U9419 (N_9419,N_9212,N_9260);
nor U9420 (N_9420,N_9351,N_9336);
nor U9421 (N_9421,N_9297,N_9321);
and U9422 (N_9422,N_9286,N_9392);
nand U9423 (N_9423,N_9292,N_9346);
or U9424 (N_9424,N_9312,N_9207);
and U9425 (N_9425,N_9371,N_9219);
nor U9426 (N_9426,N_9245,N_9320);
nor U9427 (N_9427,N_9311,N_9376);
nor U9428 (N_9428,N_9393,N_9274);
nor U9429 (N_9429,N_9267,N_9327);
nor U9430 (N_9430,N_9332,N_9380);
nand U9431 (N_9431,N_9240,N_9359);
or U9432 (N_9432,N_9241,N_9281);
nor U9433 (N_9433,N_9307,N_9345);
and U9434 (N_9434,N_9244,N_9287);
and U9435 (N_9435,N_9381,N_9365);
or U9436 (N_9436,N_9317,N_9283);
nand U9437 (N_9437,N_9255,N_9323);
nor U9438 (N_9438,N_9271,N_9258);
nand U9439 (N_9439,N_9269,N_9261);
xnor U9440 (N_9440,N_9349,N_9397);
or U9441 (N_9441,N_9277,N_9325);
nor U9442 (N_9442,N_9382,N_9357);
or U9443 (N_9443,N_9315,N_9324);
nand U9444 (N_9444,N_9285,N_9290);
nor U9445 (N_9445,N_9330,N_9305);
or U9446 (N_9446,N_9275,N_9329);
nand U9447 (N_9447,N_9322,N_9227);
nor U9448 (N_9448,N_9270,N_9232);
nor U9449 (N_9449,N_9362,N_9243);
or U9450 (N_9450,N_9236,N_9314);
and U9451 (N_9451,N_9370,N_9248);
or U9452 (N_9452,N_9308,N_9398);
nand U9453 (N_9453,N_9262,N_9238);
nand U9454 (N_9454,N_9348,N_9385);
and U9455 (N_9455,N_9368,N_9383);
and U9456 (N_9456,N_9366,N_9387);
or U9457 (N_9457,N_9390,N_9222);
and U9458 (N_9458,N_9201,N_9389);
or U9459 (N_9459,N_9379,N_9220);
nor U9460 (N_9460,N_9200,N_9242);
nor U9461 (N_9461,N_9377,N_9295);
or U9462 (N_9462,N_9344,N_9360);
nor U9463 (N_9463,N_9302,N_9358);
nand U9464 (N_9464,N_9257,N_9235);
nor U9465 (N_9465,N_9266,N_9254);
nor U9466 (N_9466,N_9372,N_9252);
nand U9467 (N_9467,N_9263,N_9205);
and U9468 (N_9468,N_9223,N_9363);
nor U9469 (N_9469,N_9306,N_9231);
and U9470 (N_9470,N_9278,N_9296);
nor U9471 (N_9471,N_9374,N_9333);
or U9472 (N_9472,N_9273,N_9355);
and U9473 (N_9473,N_9391,N_9299);
nand U9474 (N_9474,N_9309,N_9272);
or U9475 (N_9475,N_9214,N_9335);
and U9476 (N_9476,N_9209,N_9226);
and U9477 (N_9477,N_9361,N_9211);
nand U9478 (N_9478,N_9229,N_9367);
or U9479 (N_9479,N_9352,N_9208);
and U9480 (N_9480,N_9224,N_9203);
nor U9481 (N_9481,N_9202,N_9213);
nand U9482 (N_9482,N_9234,N_9204);
nand U9483 (N_9483,N_9313,N_9340);
nor U9484 (N_9484,N_9316,N_9282);
nor U9485 (N_9485,N_9353,N_9350);
nor U9486 (N_9486,N_9303,N_9331);
nand U9487 (N_9487,N_9386,N_9375);
xnor U9488 (N_9488,N_9230,N_9228);
nand U9489 (N_9489,N_9347,N_9337);
and U9490 (N_9490,N_9239,N_9394);
nor U9491 (N_9491,N_9225,N_9369);
nand U9492 (N_9492,N_9294,N_9237);
nand U9493 (N_9493,N_9293,N_9341);
nor U9494 (N_9494,N_9256,N_9354);
xnor U9495 (N_9495,N_9265,N_9334);
and U9496 (N_9496,N_9280,N_9373);
nand U9497 (N_9497,N_9301,N_9304);
nand U9498 (N_9498,N_9399,N_9268);
nand U9499 (N_9499,N_9328,N_9310);
nand U9500 (N_9500,N_9389,N_9300);
nor U9501 (N_9501,N_9378,N_9325);
nor U9502 (N_9502,N_9251,N_9325);
nand U9503 (N_9503,N_9383,N_9234);
or U9504 (N_9504,N_9397,N_9394);
nand U9505 (N_9505,N_9295,N_9381);
nor U9506 (N_9506,N_9366,N_9333);
nor U9507 (N_9507,N_9241,N_9324);
nand U9508 (N_9508,N_9227,N_9253);
and U9509 (N_9509,N_9216,N_9204);
nor U9510 (N_9510,N_9380,N_9251);
or U9511 (N_9511,N_9333,N_9269);
and U9512 (N_9512,N_9319,N_9202);
nand U9513 (N_9513,N_9356,N_9398);
nor U9514 (N_9514,N_9238,N_9320);
or U9515 (N_9515,N_9367,N_9267);
and U9516 (N_9516,N_9226,N_9341);
nor U9517 (N_9517,N_9317,N_9270);
or U9518 (N_9518,N_9397,N_9301);
nand U9519 (N_9519,N_9332,N_9297);
and U9520 (N_9520,N_9263,N_9247);
and U9521 (N_9521,N_9388,N_9297);
or U9522 (N_9522,N_9211,N_9332);
nor U9523 (N_9523,N_9337,N_9395);
nand U9524 (N_9524,N_9327,N_9309);
nand U9525 (N_9525,N_9382,N_9310);
and U9526 (N_9526,N_9207,N_9343);
nand U9527 (N_9527,N_9279,N_9226);
and U9528 (N_9528,N_9392,N_9363);
nand U9529 (N_9529,N_9298,N_9295);
or U9530 (N_9530,N_9222,N_9341);
or U9531 (N_9531,N_9294,N_9260);
nor U9532 (N_9532,N_9380,N_9212);
or U9533 (N_9533,N_9285,N_9359);
nor U9534 (N_9534,N_9205,N_9216);
or U9535 (N_9535,N_9249,N_9394);
nor U9536 (N_9536,N_9254,N_9358);
and U9537 (N_9537,N_9273,N_9382);
nor U9538 (N_9538,N_9256,N_9394);
and U9539 (N_9539,N_9352,N_9360);
or U9540 (N_9540,N_9224,N_9381);
nand U9541 (N_9541,N_9207,N_9250);
or U9542 (N_9542,N_9370,N_9357);
and U9543 (N_9543,N_9310,N_9214);
or U9544 (N_9544,N_9352,N_9229);
or U9545 (N_9545,N_9219,N_9388);
and U9546 (N_9546,N_9289,N_9297);
and U9547 (N_9547,N_9336,N_9392);
nand U9548 (N_9548,N_9253,N_9375);
nor U9549 (N_9549,N_9343,N_9351);
and U9550 (N_9550,N_9225,N_9281);
or U9551 (N_9551,N_9292,N_9289);
or U9552 (N_9552,N_9389,N_9309);
xnor U9553 (N_9553,N_9287,N_9339);
or U9554 (N_9554,N_9363,N_9358);
and U9555 (N_9555,N_9216,N_9229);
nor U9556 (N_9556,N_9282,N_9372);
nand U9557 (N_9557,N_9329,N_9384);
or U9558 (N_9558,N_9349,N_9251);
and U9559 (N_9559,N_9389,N_9369);
and U9560 (N_9560,N_9262,N_9386);
nand U9561 (N_9561,N_9220,N_9336);
or U9562 (N_9562,N_9290,N_9275);
nor U9563 (N_9563,N_9362,N_9334);
or U9564 (N_9564,N_9379,N_9295);
and U9565 (N_9565,N_9254,N_9354);
nor U9566 (N_9566,N_9273,N_9225);
xnor U9567 (N_9567,N_9362,N_9264);
nor U9568 (N_9568,N_9391,N_9310);
nor U9569 (N_9569,N_9333,N_9341);
and U9570 (N_9570,N_9294,N_9385);
nor U9571 (N_9571,N_9395,N_9307);
or U9572 (N_9572,N_9244,N_9237);
and U9573 (N_9573,N_9357,N_9319);
nand U9574 (N_9574,N_9334,N_9226);
nand U9575 (N_9575,N_9340,N_9222);
or U9576 (N_9576,N_9217,N_9297);
and U9577 (N_9577,N_9262,N_9340);
nand U9578 (N_9578,N_9335,N_9291);
nand U9579 (N_9579,N_9221,N_9328);
or U9580 (N_9580,N_9359,N_9260);
or U9581 (N_9581,N_9270,N_9361);
and U9582 (N_9582,N_9291,N_9218);
or U9583 (N_9583,N_9367,N_9215);
or U9584 (N_9584,N_9214,N_9347);
nand U9585 (N_9585,N_9310,N_9290);
nor U9586 (N_9586,N_9262,N_9263);
or U9587 (N_9587,N_9364,N_9265);
and U9588 (N_9588,N_9260,N_9213);
nand U9589 (N_9589,N_9266,N_9267);
nor U9590 (N_9590,N_9382,N_9244);
or U9591 (N_9591,N_9397,N_9318);
nand U9592 (N_9592,N_9283,N_9268);
and U9593 (N_9593,N_9205,N_9388);
and U9594 (N_9594,N_9293,N_9339);
nor U9595 (N_9595,N_9316,N_9395);
nor U9596 (N_9596,N_9271,N_9356);
nor U9597 (N_9597,N_9383,N_9269);
nor U9598 (N_9598,N_9202,N_9360);
or U9599 (N_9599,N_9295,N_9223);
or U9600 (N_9600,N_9591,N_9478);
and U9601 (N_9601,N_9441,N_9592);
nor U9602 (N_9602,N_9451,N_9471);
nor U9603 (N_9603,N_9489,N_9568);
nor U9604 (N_9604,N_9550,N_9516);
and U9605 (N_9605,N_9488,N_9452);
and U9606 (N_9606,N_9599,N_9502);
nor U9607 (N_9607,N_9407,N_9566);
nand U9608 (N_9608,N_9512,N_9561);
and U9609 (N_9609,N_9507,N_9575);
or U9610 (N_9610,N_9560,N_9556);
and U9611 (N_9611,N_9505,N_9521);
nand U9612 (N_9612,N_9477,N_9496);
nor U9613 (N_9613,N_9576,N_9589);
and U9614 (N_9614,N_9424,N_9584);
and U9615 (N_9615,N_9492,N_9569);
or U9616 (N_9616,N_9457,N_9447);
nand U9617 (N_9617,N_9462,N_9433);
or U9618 (N_9618,N_9445,N_9586);
or U9619 (N_9619,N_9444,N_9408);
and U9620 (N_9620,N_9446,N_9526);
and U9621 (N_9621,N_9532,N_9465);
nor U9622 (N_9622,N_9522,N_9443);
nand U9623 (N_9623,N_9406,N_9476);
nor U9624 (N_9624,N_9503,N_9497);
and U9625 (N_9625,N_9494,N_9551);
nor U9626 (N_9626,N_9564,N_9455);
and U9627 (N_9627,N_9475,N_9588);
nand U9628 (N_9628,N_9583,N_9417);
or U9629 (N_9629,N_9423,N_9411);
nand U9630 (N_9630,N_9439,N_9514);
nor U9631 (N_9631,N_9544,N_9429);
and U9632 (N_9632,N_9504,N_9578);
nor U9633 (N_9633,N_9402,N_9437);
nand U9634 (N_9634,N_9416,N_9529);
nand U9635 (N_9635,N_9421,N_9425);
xor U9636 (N_9636,N_9563,N_9539);
xnor U9637 (N_9637,N_9559,N_9519);
and U9638 (N_9638,N_9414,N_9440);
or U9639 (N_9639,N_9453,N_9510);
nor U9640 (N_9640,N_9552,N_9422);
nand U9641 (N_9641,N_9596,N_9579);
nor U9642 (N_9642,N_9483,N_9509);
nand U9643 (N_9643,N_9403,N_9405);
nand U9644 (N_9644,N_9506,N_9543);
nor U9645 (N_9645,N_9523,N_9518);
nor U9646 (N_9646,N_9595,N_9581);
and U9647 (N_9647,N_9580,N_9412);
nor U9648 (N_9648,N_9495,N_9540);
nor U9649 (N_9649,N_9449,N_9585);
or U9650 (N_9650,N_9400,N_9486);
or U9651 (N_9651,N_9463,N_9577);
nor U9652 (N_9652,N_9511,N_9573);
nor U9653 (N_9653,N_9466,N_9474);
or U9654 (N_9654,N_9428,N_9553);
or U9655 (N_9655,N_9554,N_9545);
nand U9656 (N_9656,N_9438,N_9582);
nand U9657 (N_9657,N_9430,N_9415);
nor U9658 (N_9658,N_9537,N_9468);
nor U9659 (N_9659,N_9542,N_9538);
and U9660 (N_9660,N_9448,N_9517);
and U9661 (N_9661,N_9533,N_9469);
nand U9662 (N_9662,N_9470,N_9434);
nor U9663 (N_9663,N_9546,N_9593);
and U9664 (N_9664,N_9572,N_9590);
nor U9665 (N_9665,N_9456,N_9419);
or U9666 (N_9666,N_9513,N_9480);
nand U9667 (N_9667,N_9558,N_9515);
and U9668 (N_9668,N_9565,N_9479);
nand U9669 (N_9669,N_9482,N_9500);
or U9670 (N_9670,N_9459,N_9485);
nand U9671 (N_9671,N_9528,N_9426);
nor U9672 (N_9672,N_9549,N_9534);
and U9673 (N_9673,N_9501,N_9562);
and U9674 (N_9674,N_9490,N_9530);
and U9675 (N_9675,N_9410,N_9547);
or U9676 (N_9676,N_9555,N_9401);
nor U9677 (N_9677,N_9432,N_9570);
and U9678 (N_9678,N_9454,N_9436);
nand U9679 (N_9679,N_9467,N_9409);
or U9680 (N_9680,N_9427,N_9404);
or U9681 (N_9681,N_9535,N_9587);
and U9682 (N_9682,N_9520,N_9548);
and U9683 (N_9683,N_9450,N_9481);
nand U9684 (N_9684,N_9431,N_9524);
or U9685 (N_9685,N_9527,N_9598);
and U9686 (N_9686,N_9472,N_9460);
or U9687 (N_9687,N_9557,N_9435);
or U9688 (N_9688,N_9442,N_9536);
or U9689 (N_9689,N_9574,N_9531);
nand U9690 (N_9690,N_9508,N_9487);
nor U9691 (N_9691,N_9458,N_9484);
nand U9692 (N_9692,N_9461,N_9413);
and U9693 (N_9693,N_9571,N_9498);
nand U9694 (N_9694,N_9541,N_9525);
nor U9695 (N_9695,N_9418,N_9464);
nor U9696 (N_9696,N_9473,N_9594);
nand U9697 (N_9697,N_9567,N_9597);
xnor U9698 (N_9698,N_9491,N_9420);
or U9699 (N_9699,N_9499,N_9493);
or U9700 (N_9700,N_9422,N_9562);
nor U9701 (N_9701,N_9416,N_9481);
and U9702 (N_9702,N_9464,N_9403);
and U9703 (N_9703,N_9462,N_9420);
nor U9704 (N_9704,N_9492,N_9552);
nand U9705 (N_9705,N_9526,N_9567);
and U9706 (N_9706,N_9412,N_9540);
and U9707 (N_9707,N_9508,N_9429);
or U9708 (N_9708,N_9441,N_9454);
nand U9709 (N_9709,N_9550,N_9572);
and U9710 (N_9710,N_9419,N_9541);
nand U9711 (N_9711,N_9473,N_9493);
nand U9712 (N_9712,N_9505,N_9461);
nor U9713 (N_9713,N_9446,N_9535);
nor U9714 (N_9714,N_9439,N_9425);
or U9715 (N_9715,N_9519,N_9579);
nand U9716 (N_9716,N_9551,N_9510);
nand U9717 (N_9717,N_9585,N_9537);
and U9718 (N_9718,N_9422,N_9440);
nand U9719 (N_9719,N_9501,N_9585);
nor U9720 (N_9720,N_9506,N_9552);
or U9721 (N_9721,N_9526,N_9506);
or U9722 (N_9722,N_9469,N_9483);
nor U9723 (N_9723,N_9434,N_9505);
nand U9724 (N_9724,N_9569,N_9528);
or U9725 (N_9725,N_9452,N_9536);
or U9726 (N_9726,N_9476,N_9411);
or U9727 (N_9727,N_9414,N_9462);
and U9728 (N_9728,N_9427,N_9428);
or U9729 (N_9729,N_9492,N_9574);
nand U9730 (N_9730,N_9593,N_9564);
or U9731 (N_9731,N_9464,N_9441);
or U9732 (N_9732,N_9461,N_9490);
and U9733 (N_9733,N_9443,N_9596);
nand U9734 (N_9734,N_9503,N_9448);
and U9735 (N_9735,N_9472,N_9522);
nor U9736 (N_9736,N_9510,N_9509);
nor U9737 (N_9737,N_9504,N_9582);
nor U9738 (N_9738,N_9466,N_9476);
and U9739 (N_9739,N_9426,N_9405);
nor U9740 (N_9740,N_9475,N_9406);
nand U9741 (N_9741,N_9525,N_9570);
nand U9742 (N_9742,N_9513,N_9578);
or U9743 (N_9743,N_9551,N_9541);
or U9744 (N_9744,N_9533,N_9572);
nor U9745 (N_9745,N_9468,N_9406);
nor U9746 (N_9746,N_9578,N_9400);
or U9747 (N_9747,N_9437,N_9576);
nand U9748 (N_9748,N_9552,N_9437);
nor U9749 (N_9749,N_9594,N_9425);
or U9750 (N_9750,N_9442,N_9485);
nand U9751 (N_9751,N_9583,N_9432);
nand U9752 (N_9752,N_9413,N_9491);
nor U9753 (N_9753,N_9466,N_9475);
and U9754 (N_9754,N_9590,N_9599);
nand U9755 (N_9755,N_9526,N_9581);
and U9756 (N_9756,N_9547,N_9509);
nand U9757 (N_9757,N_9422,N_9545);
or U9758 (N_9758,N_9491,N_9571);
nor U9759 (N_9759,N_9485,N_9598);
nor U9760 (N_9760,N_9586,N_9465);
or U9761 (N_9761,N_9494,N_9587);
nor U9762 (N_9762,N_9550,N_9541);
nor U9763 (N_9763,N_9489,N_9495);
nand U9764 (N_9764,N_9481,N_9559);
or U9765 (N_9765,N_9526,N_9427);
or U9766 (N_9766,N_9462,N_9458);
or U9767 (N_9767,N_9466,N_9434);
nand U9768 (N_9768,N_9489,N_9462);
or U9769 (N_9769,N_9483,N_9537);
nor U9770 (N_9770,N_9469,N_9489);
or U9771 (N_9771,N_9487,N_9561);
and U9772 (N_9772,N_9571,N_9434);
nor U9773 (N_9773,N_9580,N_9456);
nand U9774 (N_9774,N_9528,N_9427);
nor U9775 (N_9775,N_9586,N_9492);
or U9776 (N_9776,N_9542,N_9507);
nor U9777 (N_9777,N_9455,N_9413);
nor U9778 (N_9778,N_9435,N_9597);
nor U9779 (N_9779,N_9474,N_9536);
or U9780 (N_9780,N_9599,N_9409);
and U9781 (N_9781,N_9429,N_9570);
or U9782 (N_9782,N_9536,N_9424);
nor U9783 (N_9783,N_9427,N_9598);
and U9784 (N_9784,N_9448,N_9485);
or U9785 (N_9785,N_9515,N_9467);
or U9786 (N_9786,N_9516,N_9424);
and U9787 (N_9787,N_9529,N_9493);
and U9788 (N_9788,N_9515,N_9589);
nand U9789 (N_9789,N_9450,N_9577);
and U9790 (N_9790,N_9475,N_9561);
and U9791 (N_9791,N_9440,N_9559);
nand U9792 (N_9792,N_9569,N_9473);
nand U9793 (N_9793,N_9581,N_9573);
nor U9794 (N_9794,N_9471,N_9587);
or U9795 (N_9795,N_9441,N_9533);
nor U9796 (N_9796,N_9433,N_9538);
nor U9797 (N_9797,N_9409,N_9489);
or U9798 (N_9798,N_9459,N_9400);
and U9799 (N_9799,N_9584,N_9582);
or U9800 (N_9800,N_9626,N_9718);
or U9801 (N_9801,N_9680,N_9684);
nand U9802 (N_9802,N_9747,N_9658);
nand U9803 (N_9803,N_9636,N_9752);
nor U9804 (N_9804,N_9727,N_9635);
and U9805 (N_9805,N_9751,N_9762);
nor U9806 (N_9806,N_9616,N_9639);
nand U9807 (N_9807,N_9646,N_9659);
nand U9808 (N_9808,N_9699,N_9799);
nand U9809 (N_9809,N_9613,N_9783);
or U9810 (N_9810,N_9733,N_9710);
nand U9811 (N_9811,N_9722,N_9771);
nor U9812 (N_9812,N_9707,N_9624);
nor U9813 (N_9813,N_9679,N_9629);
xor U9814 (N_9814,N_9774,N_9760);
nor U9815 (N_9815,N_9661,N_9753);
nor U9816 (N_9816,N_9728,N_9731);
nand U9817 (N_9817,N_9691,N_9706);
and U9818 (N_9818,N_9627,N_9721);
and U9819 (N_9819,N_9677,N_9656);
nor U9820 (N_9820,N_9697,N_9772);
and U9821 (N_9821,N_9605,N_9792);
or U9822 (N_9822,N_9675,N_9609);
or U9823 (N_9823,N_9701,N_9637);
and U9824 (N_9824,N_9734,N_9726);
nor U9825 (N_9825,N_9761,N_9739);
nor U9826 (N_9826,N_9669,N_9730);
and U9827 (N_9827,N_9686,N_9676);
nand U9828 (N_9828,N_9708,N_9600);
nand U9829 (N_9829,N_9786,N_9749);
and U9830 (N_9830,N_9655,N_9615);
xor U9831 (N_9831,N_9693,N_9777);
or U9832 (N_9832,N_9644,N_9740);
or U9833 (N_9833,N_9745,N_9780);
nand U9834 (N_9834,N_9610,N_9689);
or U9835 (N_9835,N_9793,N_9607);
nor U9836 (N_9836,N_9608,N_9744);
xnor U9837 (N_9837,N_9754,N_9711);
nor U9838 (N_9838,N_9647,N_9781);
nand U9839 (N_9839,N_9763,N_9724);
nand U9840 (N_9840,N_9756,N_9723);
nor U9841 (N_9841,N_9787,N_9640);
nand U9842 (N_9842,N_9719,N_9714);
and U9843 (N_9843,N_9736,N_9653);
nor U9844 (N_9844,N_9667,N_9798);
and U9845 (N_9845,N_9601,N_9622);
or U9846 (N_9846,N_9789,N_9611);
nand U9847 (N_9847,N_9758,N_9621);
nand U9848 (N_9848,N_9709,N_9790);
or U9849 (N_9849,N_9769,N_9682);
nor U9850 (N_9850,N_9666,N_9620);
and U9851 (N_9851,N_9654,N_9784);
or U9852 (N_9852,N_9649,N_9770);
and U9853 (N_9853,N_9604,N_9700);
nand U9854 (N_9854,N_9650,N_9750);
or U9855 (N_9855,N_9619,N_9618);
and U9856 (N_9856,N_9795,N_9735);
and U9857 (N_9857,N_9634,N_9757);
nand U9858 (N_9858,N_9705,N_9732);
nand U9859 (N_9859,N_9641,N_9632);
or U9860 (N_9860,N_9746,N_9678);
or U9861 (N_9861,N_9696,N_9743);
nand U9862 (N_9862,N_9741,N_9651);
or U9863 (N_9863,N_9692,N_9778);
nand U9864 (N_9864,N_9704,N_9687);
or U9865 (N_9865,N_9625,N_9665);
nand U9866 (N_9866,N_9788,N_9796);
nor U9867 (N_9867,N_9785,N_9766);
nand U9868 (N_9868,N_9662,N_9695);
and U9869 (N_9869,N_9755,N_9628);
or U9870 (N_9870,N_9794,N_9768);
or U9871 (N_9871,N_9694,N_9648);
nor U9872 (N_9872,N_9603,N_9671);
nor U9873 (N_9873,N_9638,N_9698);
nor U9874 (N_9874,N_9672,N_9738);
and U9875 (N_9875,N_9729,N_9614);
and U9876 (N_9876,N_9779,N_9663);
and U9877 (N_9877,N_9737,N_9657);
or U9878 (N_9878,N_9715,N_9631);
nand U9879 (N_9879,N_9685,N_9602);
or U9880 (N_9880,N_9643,N_9690);
nand U9881 (N_9881,N_9702,N_9617);
or U9882 (N_9882,N_9775,N_9764);
nand U9883 (N_9883,N_9652,N_9645);
or U9884 (N_9884,N_9791,N_9630);
nor U9885 (N_9885,N_9664,N_9606);
or U9886 (N_9886,N_9742,N_9683);
or U9887 (N_9887,N_9681,N_9717);
nand U9888 (N_9888,N_9716,N_9782);
and U9889 (N_9889,N_9767,N_9612);
and U9890 (N_9890,N_9642,N_9668);
and U9891 (N_9891,N_9713,N_9673);
and U9892 (N_9892,N_9773,N_9720);
or U9893 (N_9893,N_9670,N_9633);
xnor U9894 (N_9894,N_9712,N_9748);
nand U9895 (N_9895,N_9688,N_9759);
nor U9896 (N_9896,N_9797,N_9765);
or U9897 (N_9897,N_9703,N_9674);
nor U9898 (N_9898,N_9776,N_9660);
or U9899 (N_9899,N_9725,N_9623);
nor U9900 (N_9900,N_9723,N_9706);
nand U9901 (N_9901,N_9665,N_9747);
nor U9902 (N_9902,N_9797,N_9734);
or U9903 (N_9903,N_9650,N_9742);
nor U9904 (N_9904,N_9744,N_9622);
and U9905 (N_9905,N_9629,N_9783);
nand U9906 (N_9906,N_9670,N_9680);
nand U9907 (N_9907,N_9771,N_9741);
and U9908 (N_9908,N_9614,N_9706);
or U9909 (N_9909,N_9778,N_9723);
or U9910 (N_9910,N_9734,N_9679);
or U9911 (N_9911,N_9617,N_9766);
nand U9912 (N_9912,N_9643,N_9613);
or U9913 (N_9913,N_9662,N_9717);
nor U9914 (N_9914,N_9657,N_9720);
or U9915 (N_9915,N_9644,N_9753);
nand U9916 (N_9916,N_9799,N_9693);
nand U9917 (N_9917,N_9748,N_9661);
or U9918 (N_9918,N_9692,N_9633);
nor U9919 (N_9919,N_9625,N_9645);
or U9920 (N_9920,N_9724,N_9680);
nor U9921 (N_9921,N_9726,N_9769);
and U9922 (N_9922,N_9686,N_9761);
and U9923 (N_9923,N_9664,N_9744);
nor U9924 (N_9924,N_9741,N_9668);
and U9925 (N_9925,N_9738,N_9762);
nand U9926 (N_9926,N_9673,N_9609);
or U9927 (N_9927,N_9614,N_9734);
and U9928 (N_9928,N_9664,N_9725);
nor U9929 (N_9929,N_9764,N_9634);
nand U9930 (N_9930,N_9768,N_9799);
nor U9931 (N_9931,N_9760,N_9747);
and U9932 (N_9932,N_9608,N_9756);
and U9933 (N_9933,N_9728,N_9729);
nor U9934 (N_9934,N_9772,N_9605);
nand U9935 (N_9935,N_9709,N_9739);
nor U9936 (N_9936,N_9664,N_9624);
or U9937 (N_9937,N_9764,N_9708);
and U9938 (N_9938,N_9611,N_9775);
and U9939 (N_9939,N_9705,N_9798);
nor U9940 (N_9940,N_9754,N_9741);
and U9941 (N_9941,N_9676,N_9647);
and U9942 (N_9942,N_9705,N_9685);
and U9943 (N_9943,N_9752,N_9654);
and U9944 (N_9944,N_9798,N_9708);
or U9945 (N_9945,N_9687,N_9722);
nand U9946 (N_9946,N_9703,N_9754);
nor U9947 (N_9947,N_9719,N_9700);
or U9948 (N_9948,N_9616,N_9767);
or U9949 (N_9949,N_9768,N_9683);
or U9950 (N_9950,N_9781,N_9762);
and U9951 (N_9951,N_9627,N_9780);
and U9952 (N_9952,N_9720,N_9618);
or U9953 (N_9953,N_9604,N_9617);
and U9954 (N_9954,N_9674,N_9649);
and U9955 (N_9955,N_9734,N_9654);
or U9956 (N_9956,N_9601,N_9749);
nor U9957 (N_9957,N_9633,N_9744);
or U9958 (N_9958,N_9635,N_9756);
or U9959 (N_9959,N_9725,N_9783);
nor U9960 (N_9960,N_9725,N_9782);
or U9961 (N_9961,N_9779,N_9743);
or U9962 (N_9962,N_9662,N_9750);
nand U9963 (N_9963,N_9694,N_9794);
and U9964 (N_9964,N_9734,N_9652);
nor U9965 (N_9965,N_9734,N_9717);
and U9966 (N_9966,N_9754,N_9782);
or U9967 (N_9967,N_9781,N_9685);
nor U9968 (N_9968,N_9790,N_9756);
and U9969 (N_9969,N_9635,N_9703);
or U9970 (N_9970,N_9739,N_9619);
nand U9971 (N_9971,N_9640,N_9771);
nand U9972 (N_9972,N_9761,N_9647);
nor U9973 (N_9973,N_9690,N_9681);
nand U9974 (N_9974,N_9748,N_9730);
and U9975 (N_9975,N_9619,N_9770);
nand U9976 (N_9976,N_9795,N_9775);
or U9977 (N_9977,N_9662,N_9615);
and U9978 (N_9978,N_9754,N_9660);
nand U9979 (N_9979,N_9744,N_9628);
nand U9980 (N_9980,N_9683,N_9737);
nor U9981 (N_9981,N_9600,N_9651);
nor U9982 (N_9982,N_9675,N_9757);
and U9983 (N_9983,N_9708,N_9635);
and U9984 (N_9984,N_9703,N_9667);
or U9985 (N_9985,N_9786,N_9699);
nand U9986 (N_9986,N_9716,N_9737);
and U9987 (N_9987,N_9783,N_9623);
nor U9988 (N_9988,N_9625,N_9791);
nor U9989 (N_9989,N_9687,N_9767);
nand U9990 (N_9990,N_9667,N_9767);
nor U9991 (N_9991,N_9743,N_9634);
nor U9992 (N_9992,N_9763,N_9697);
or U9993 (N_9993,N_9680,N_9745);
and U9994 (N_9994,N_9699,N_9618);
nor U9995 (N_9995,N_9668,N_9641);
or U9996 (N_9996,N_9731,N_9612);
or U9997 (N_9997,N_9715,N_9716);
or U9998 (N_9998,N_9762,N_9683);
or U9999 (N_9999,N_9710,N_9734);
and UO_0 (O_0,N_9837,N_9938);
nor UO_1 (O_1,N_9974,N_9825);
nand UO_2 (O_2,N_9843,N_9893);
nor UO_3 (O_3,N_9888,N_9852);
nand UO_4 (O_4,N_9981,N_9871);
or UO_5 (O_5,N_9891,N_9889);
or UO_6 (O_6,N_9967,N_9870);
or UO_7 (O_7,N_9965,N_9853);
nor UO_8 (O_8,N_9863,N_9934);
and UO_9 (O_9,N_9840,N_9897);
and UO_10 (O_10,N_9945,N_9961);
or UO_11 (O_11,N_9907,N_9867);
nor UO_12 (O_12,N_9818,N_9994);
and UO_13 (O_13,N_9817,N_9845);
nand UO_14 (O_14,N_9873,N_9808);
nand UO_15 (O_15,N_9856,N_9930);
nor UO_16 (O_16,N_9922,N_9946);
nor UO_17 (O_17,N_9906,N_9892);
nor UO_18 (O_18,N_9958,N_9838);
nor UO_19 (O_19,N_9957,N_9842);
or UO_20 (O_20,N_9857,N_9991);
nand UO_21 (O_21,N_9855,N_9908);
and UO_22 (O_22,N_9882,N_9992);
or UO_23 (O_23,N_9877,N_9803);
or UO_24 (O_24,N_9836,N_9829);
and UO_25 (O_25,N_9848,N_9936);
nor UO_26 (O_26,N_9971,N_9850);
nand UO_27 (O_27,N_9968,N_9869);
or UO_28 (O_28,N_9885,N_9914);
nor UO_29 (O_29,N_9951,N_9821);
nor UO_30 (O_30,N_9831,N_9866);
or UO_31 (O_31,N_9832,N_9802);
or UO_32 (O_32,N_9890,N_9865);
nor UO_33 (O_33,N_9809,N_9966);
or UO_34 (O_34,N_9886,N_9811);
and UO_35 (O_35,N_9833,N_9859);
and UO_36 (O_36,N_9989,N_9985);
and UO_37 (O_37,N_9874,N_9955);
nand UO_38 (O_38,N_9923,N_9804);
nor UO_39 (O_39,N_9827,N_9878);
or UO_40 (O_40,N_9862,N_9800);
nand UO_41 (O_41,N_9988,N_9830);
nand UO_42 (O_42,N_9987,N_9999);
and UO_43 (O_43,N_9844,N_9929);
or UO_44 (O_44,N_9997,N_9998);
nand UO_45 (O_45,N_9933,N_9948);
and UO_46 (O_46,N_9875,N_9953);
and UO_47 (O_47,N_9959,N_9954);
or UO_48 (O_48,N_9903,N_9816);
or UO_49 (O_49,N_9973,N_9916);
or UO_50 (O_50,N_9805,N_9801);
nand UO_51 (O_51,N_9978,N_9847);
nand UO_52 (O_52,N_9883,N_9944);
nand UO_53 (O_53,N_9949,N_9849);
or UO_54 (O_54,N_9943,N_9814);
nand UO_55 (O_55,N_9980,N_9927);
and UO_56 (O_56,N_9928,N_9960);
nand UO_57 (O_57,N_9977,N_9826);
nor UO_58 (O_58,N_9828,N_9900);
and UO_59 (O_59,N_9952,N_9815);
or UO_60 (O_60,N_9919,N_9822);
nor UO_61 (O_61,N_9879,N_9915);
nor UO_62 (O_62,N_9986,N_9824);
or UO_63 (O_63,N_9950,N_9939);
or UO_64 (O_64,N_9932,N_9975);
nor UO_65 (O_65,N_9881,N_9823);
nor UO_66 (O_66,N_9993,N_9872);
nor UO_67 (O_67,N_9920,N_9983);
nand UO_68 (O_68,N_9868,N_9813);
or UO_69 (O_69,N_9931,N_9912);
nor UO_70 (O_70,N_9896,N_9962);
or UO_71 (O_71,N_9851,N_9937);
nand UO_72 (O_72,N_9972,N_9940);
and UO_73 (O_73,N_9901,N_9819);
nor UO_74 (O_74,N_9925,N_9895);
nor UO_75 (O_75,N_9963,N_9941);
nand UO_76 (O_76,N_9947,N_9887);
nor UO_77 (O_77,N_9820,N_9969);
nand UO_78 (O_78,N_9810,N_9905);
or UO_79 (O_79,N_9894,N_9858);
nand UO_80 (O_80,N_9902,N_9964);
nor UO_81 (O_81,N_9904,N_9876);
nor UO_82 (O_82,N_9909,N_9921);
or UO_83 (O_83,N_9880,N_9812);
or UO_84 (O_84,N_9935,N_9924);
nor UO_85 (O_85,N_9898,N_9807);
or UO_86 (O_86,N_9979,N_9861);
nor UO_87 (O_87,N_9976,N_9913);
nor UO_88 (O_88,N_9996,N_9884);
and UO_89 (O_89,N_9864,N_9970);
nand UO_90 (O_90,N_9995,N_9860);
or UO_91 (O_91,N_9911,N_9984);
nand UO_92 (O_92,N_9841,N_9839);
and UO_93 (O_93,N_9942,N_9854);
nor UO_94 (O_94,N_9910,N_9917);
or UO_95 (O_95,N_9982,N_9918);
or UO_96 (O_96,N_9835,N_9990);
nor UO_97 (O_97,N_9834,N_9806);
and UO_98 (O_98,N_9926,N_9956);
nor UO_99 (O_99,N_9899,N_9846);
and UO_100 (O_100,N_9816,N_9997);
or UO_101 (O_101,N_9893,N_9857);
and UO_102 (O_102,N_9997,N_9882);
nand UO_103 (O_103,N_9962,N_9807);
nand UO_104 (O_104,N_9978,N_9880);
and UO_105 (O_105,N_9919,N_9888);
nor UO_106 (O_106,N_9883,N_9933);
nor UO_107 (O_107,N_9932,N_9862);
nor UO_108 (O_108,N_9861,N_9878);
nand UO_109 (O_109,N_9887,N_9831);
and UO_110 (O_110,N_9866,N_9960);
and UO_111 (O_111,N_9873,N_9850);
nand UO_112 (O_112,N_9885,N_9908);
or UO_113 (O_113,N_9809,N_9959);
nand UO_114 (O_114,N_9880,N_9861);
and UO_115 (O_115,N_9831,N_9802);
and UO_116 (O_116,N_9934,N_9837);
or UO_117 (O_117,N_9887,N_9931);
or UO_118 (O_118,N_9948,N_9915);
nand UO_119 (O_119,N_9863,N_9804);
nor UO_120 (O_120,N_9903,N_9880);
nor UO_121 (O_121,N_9902,N_9942);
nor UO_122 (O_122,N_9964,N_9843);
nor UO_123 (O_123,N_9834,N_9940);
or UO_124 (O_124,N_9892,N_9897);
and UO_125 (O_125,N_9827,N_9966);
nand UO_126 (O_126,N_9989,N_9808);
and UO_127 (O_127,N_9972,N_9821);
or UO_128 (O_128,N_9896,N_9977);
nand UO_129 (O_129,N_9968,N_9877);
or UO_130 (O_130,N_9825,N_9897);
and UO_131 (O_131,N_9879,N_9908);
and UO_132 (O_132,N_9857,N_9935);
or UO_133 (O_133,N_9915,N_9914);
or UO_134 (O_134,N_9938,N_9986);
nor UO_135 (O_135,N_9999,N_9904);
and UO_136 (O_136,N_9884,N_9899);
nand UO_137 (O_137,N_9910,N_9808);
nor UO_138 (O_138,N_9979,N_9911);
or UO_139 (O_139,N_9979,N_9918);
and UO_140 (O_140,N_9971,N_9939);
nor UO_141 (O_141,N_9879,N_9992);
or UO_142 (O_142,N_9894,N_9964);
nor UO_143 (O_143,N_9872,N_9804);
or UO_144 (O_144,N_9949,N_9802);
and UO_145 (O_145,N_9874,N_9845);
nand UO_146 (O_146,N_9896,N_9887);
nor UO_147 (O_147,N_9804,N_9888);
and UO_148 (O_148,N_9883,N_9853);
nor UO_149 (O_149,N_9895,N_9911);
nand UO_150 (O_150,N_9904,N_9981);
and UO_151 (O_151,N_9918,N_9944);
nand UO_152 (O_152,N_9941,N_9937);
nor UO_153 (O_153,N_9918,N_9891);
nand UO_154 (O_154,N_9951,N_9940);
and UO_155 (O_155,N_9933,N_9837);
nor UO_156 (O_156,N_9880,N_9901);
or UO_157 (O_157,N_9867,N_9958);
and UO_158 (O_158,N_9912,N_9957);
and UO_159 (O_159,N_9918,N_9991);
nor UO_160 (O_160,N_9846,N_9956);
nand UO_161 (O_161,N_9836,N_9989);
and UO_162 (O_162,N_9871,N_9955);
and UO_163 (O_163,N_9837,N_9820);
nor UO_164 (O_164,N_9972,N_9952);
nand UO_165 (O_165,N_9895,N_9834);
and UO_166 (O_166,N_9821,N_9822);
or UO_167 (O_167,N_9979,N_9949);
nor UO_168 (O_168,N_9878,N_9800);
nor UO_169 (O_169,N_9852,N_9958);
nor UO_170 (O_170,N_9947,N_9991);
and UO_171 (O_171,N_9867,N_9987);
nand UO_172 (O_172,N_9992,N_9959);
or UO_173 (O_173,N_9873,N_9835);
or UO_174 (O_174,N_9856,N_9907);
and UO_175 (O_175,N_9836,N_9801);
and UO_176 (O_176,N_9914,N_9825);
nand UO_177 (O_177,N_9895,N_9972);
nand UO_178 (O_178,N_9943,N_9905);
nor UO_179 (O_179,N_9802,N_9921);
nand UO_180 (O_180,N_9908,N_9930);
and UO_181 (O_181,N_9878,N_9956);
or UO_182 (O_182,N_9889,N_9896);
and UO_183 (O_183,N_9965,N_9959);
nand UO_184 (O_184,N_9802,N_9992);
nor UO_185 (O_185,N_9870,N_9812);
and UO_186 (O_186,N_9889,N_9928);
nor UO_187 (O_187,N_9897,N_9942);
nand UO_188 (O_188,N_9992,N_9814);
nand UO_189 (O_189,N_9869,N_9916);
nand UO_190 (O_190,N_9951,N_9887);
and UO_191 (O_191,N_9933,N_9832);
and UO_192 (O_192,N_9945,N_9851);
and UO_193 (O_193,N_9806,N_9879);
nor UO_194 (O_194,N_9816,N_9978);
and UO_195 (O_195,N_9952,N_9862);
nand UO_196 (O_196,N_9858,N_9926);
or UO_197 (O_197,N_9911,N_9846);
or UO_198 (O_198,N_9851,N_9813);
xor UO_199 (O_199,N_9887,N_9833);
or UO_200 (O_200,N_9832,N_9870);
nand UO_201 (O_201,N_9886,N_9848);
or UO_202 (O_202,N_9862,N_9807);
xnor UO_203 (O_203,N_9869,N_9901);
nand UO_204 (O_204,N_9984,N_9959);
or UO_205 (O_205,N_9998,N_9806);
and UO_206 (O_206,N_9805,N_9961);
nor UO_207 (O_207,N_9869,N_9988);
nor UO_208 (O_208,N_9919,N_9801);
nor UO_209 (O_209,N_9803,N_9989);
nor UO_210 (O_210,N_9862,N_9935);
nor UO_211 (O_211,N_9890,N_9872);
and UO_212 (O_212,N_9972,N_9804);
nand UO_213 (O_213,N_9833,N_9992);
nand UO_214 (O_214,N_9811,N_9957);
nor UO_215 (O_215,N_9859,N_9911);
and UO_216 (O_216,N_9971,N_9977);
nand UO_217 (O_217,N_9807,N_9852);
or UO_218 (O_218,N_9886,N_9971);
nor UO_219 (O_219,N_9827,N_9871);
nor UO_220 (O_220,N_9821,N_9841);
nand UO_221 (O_221,N_9999,N_9959);
nor UO_222 (O_222,N_9889,N_9941);
or UO_223 (O_223,N_9913,N_9800);
nand UO_224 (O_224,N_9812,N_9942);
nor UO_225 (O_225,N_9906,N_9876);
nand UO_226 (O_226,N_9990,N_9894);
nor UO_227 (O_227,N_9807,N_9992);
nand UO_228 (O_228,N_9945,N_9888);
and UO_229 (O_229,N_9857,N_9855);
nor UO_230 (O_230,N_9972,N_9908);
nand UO_231 (O_231,N_9949,N_9804);
or UO_232 (O_232,N_9923,N_9940);
nor UO_233 (O_233,N_9836,N_9943);
and UO_234 (O_234,N_9986,N_9818);
nor UO_235 (O_235,N_9861,N_9951);
or UO_236 (O_236,N_9833,N_9956);
and UO_237 (O_237,N_9803,N_9915);
nand UO_238 (O_238,N_9942,N_9832);
or UO_239 (O_239,N_9866,N_9953);
or UO_240 (O_240,N_9975,N_9866);
nand UO_241 (O_241,N_9816,N_9808);
nand UO_242 (O_242,N_9867,N_9989);
and UO_243 (O_243,N_9826,N_9893);
or UO_244 (O_244,N_9839,N_9973);
or UO_245 (O_245,N_9927,N_9821);
nor UO_246 (O_246,N_9938,N_9849);
nand UO_247 (O_247,N_9999,N_9875);
nor UO_248 (O_248,N_9853,N_9828);
or UO_249 (O_249,N_9844,N_9903);
nand UO_250 (O_250,N_9860,N_9886);
and UO_251 (O_251,N_9826,N_9800);
or UO_252 (O_252,N_9989,N_9941);
nor UO_253 (O_253,N_9975,N_9869);
nand UO_254 (O_254,N_9870,N_9816);
nor UO_255 (O_255,N_9800,N_9837);
and UO_256 (O_256,N_9943,N_9873);
nand UO_257 (O_257,N_9860,N_9878);
nand UO_258 (O_258,N_9937,N_9884);
or UO_259 (O_259,N_9877,N_9810);
and UO_260 (O_260,N_9903,N_9953);
and UO_261 (O_261,N_9914,N_9943);
and UO_262 (O_262,N_9805,N_9874);
and UO_263 (O_263,N_9926,N_9949);
or UO_264 (O_264,N_9939,N_9987);
and UO_265 (O_265,N_9990,N_9888);
nor UO_266 (O_266,N_9845,N_9852);
nor UO_267 (O_267,N_9918,N_9912);
nor UO_268 (O_268,N_9805,N_9881);
or UO_269 (O_269,N_9925,N_9920);
or UO_270 (O_270,N_9882,N_9917);
nand UO_271 (O_271,N_9865,N_9970);
nor UO_272 (O_272,N_9986,N_9893);
and UO_273 (O_273,N_9866,N_9992);
nor UO_274 (O_274,N_9993,N_9843);
and UO_275 (O_275,N_9808,N_9810);
or UO_276 (O_276,N_9971,N_9942);
and UO_277 (O_277,N_9830,N_9832);
or UO_278 (O_278,N_9855,N_9893);
or UO_279 (O_279,N_9904,N_9859);
nor UO_280 (O_280,N_9933,N_9867);
or UO_281 (O_281,N_9839,N_9922);
and UO_282 (O_282,N_9994,N_9970);
nor UO_283 (O_283,N_9809,N_9891);
nand UO_284 (O_284,N_9959,N_9815);
nor UO_285 (O_285,N_9828,N_9892);
nand UO_286 (O_286,N_9852,N_9971);
or UO_287 (O_287,N_9853,N_9815);
nor UO_288 (O_288,N_9929,N_9827);
or UO_289 (O_289,N_9926,N_9831);
nor UO_290 (O_290,N_9824,N_9985);
nor UO_291 (O_291,N_9908,N_9989);
nand UO_292 (O_292,N_9905,N_9914);
nand UO_293 (O_293,N_9804,N_9865);
nor UO_294 (O_294,N_9849,N_9837);
or UO_295 (O_295,N_9865,N_9905);
and UO_296 (O_296,N_9929,N_9860);
and UO_297 (O_297,N_9920,N_9908);
nor UO_298 (O_298,N_9912,N_9894);
nor UO_299 (O_299,N_9989,N_9982);
and UO_300 (O_300,N_9866,N_9835);
or UO_301 (O_301,N_9896,N_9986);
nor UO_302 (O_302,N_9930,N_9887);
and UO_303 (O_303,N_9879,N_9818);
and UO_304 (O_304,N_9988,N_9995);
or UO_305 (O_305,N_9891,N_9817);
or UO_306 (O_306,N_9916,N_9987);
or UO_307 (O_307,N_9864,N_9881);
nor UO_308 (O_308,N_9948,N_9984);
nand UO_309 (O_309,N_9870,N_9840);
or UO_310 (O_310,N_9837,N_9830);
nor UO_311 (O_311,N_9921,N_9919);
or UO_312 (O_312,N_9935,N_9960);
or UO_313 (O_313,N_9917,N_9989);
nor UO_314 (O_314,N_9970,N_9898);
nor UO_315 (O_315,N_9946,N_9844);
nand UO_316 (O_316,N_9897,N_9860);
nand UO_317 (O_317,N_9804,N_9808);
nor UO_318 (O_318,N_9964,N_9853);
or UO_319 (O_319,N_9870,N_9949);
nand UO_320 (O_320,N_9888,N_9898);
and UO_321 (O_321,N_9825,N_9894);
nand UO_322 (O_322,N_9853,N_9836);
xnor UO_323 (O_323,N_9994,N_9894);
nor UO_324 (O_324,N_9826,N_9896);
or UO_325 (O_325,N_9841,N_9880);
or UO_326 (O_326,N_9851,N_9950);
or UO_327 (O_327,N_9923,N_9991);
nand UO_328 (O_328,N_9934,N_9815);
and UO_329 (O_329,N_9921,N_9833);
nand UO_330 (O_330,N_9963,N_9865);
nor UO_331 (O_331,N_9887,N_9867);
nand UO_332 (O_332,N_9837,N_9924);
or UO_333 (O_333,N_9829,N_9831);
or UO_334 (O_334,N_9979,N_9807);
or UO_335 (O_335,N_9946,N_9979);
nor UO_336 (O_336,N_9977,N_9816);
nand UO_337 (O_337,N_9872,N_9821);
and UO_338 (O_338,N_9904,N_9860);
nand UO_339 (O_339,N_9855,N_9926);
nor UO_340 (O_340,N_9860,N_9964);
or UO_341 (O_341,N_9950,N_9982);
nand UO_342 (O_342,N_9872,N_9918);
nor UO_343 (O_343,N_9974,N_9913);
nor UO_344 (O_344,N_9985,N_9971);
and UO_345 (O_345,N_9856,N_9862);
nand UO_346 (O_346,N_9804,N_9977);
nand UO_347 (O_347,N_9943,N_9887);
nand UO_348 (O_348,N_9900,N_9993);
nand UO_349 (O_349,N_9928,N_9872);
or UO_350 (O_350,N_9814,N_9965);
nand UO_351 (O_351,N_9897,N_9889);
and UO_352 (O_352,N_9866,N_9912);
nand UO_353 (O_353,N_9907,N_9902);
or UO_354 (O_354,N_9852,N_9956);
nand UO_355 (O_355,N_9829,N_9875);
nand UO_356 (O_356,N_9966,N_9874);
xnor UO_357 (O_357,N_9903,N_9927);
nand UO_358 (O_358,N_9932,N_9804);
or UO_359 (O_359,N_9944,N_9929);
nor UO_360 (O_360,N_9957,N_9998);
and UO_361 (O_361,N_9899,N_9898);
nand UO_362 (O_362,N_9986,N_9899);
nor UO_363 (O_363,N_9903,N_9979);
and UO_364 (O_364,N_9817,N_9936);
nor UO_365 (O_365,N_9875,N_9913);
nor UO_366 (O_366,N_9932,N_9988);
nor UO_367 (O_367,N_9838,N_9867);
nand UO_368 (O_368,N_9826,N_9942);
nand UO_369 (O_369,N_9891,N_9802);
and UO_370 (O_370,N_9857,N_9847);
nand UO_371 (O_371,N_9885,N_9846);
and UO_372 (O_372,N_9839,N_9947);
and UO_373 (O_373,N_9975,N_9929);
or UO_374 (O_374,N_9852,N_9818);
nand UO_375 (O_375,N_9966,N_9851);
nand UO_376 (O_376,N_9834,N_9801);
and UO_377 (O_377,N_9952,N_9991);
nor UO_378 (O_378,N_9915,N_9811);
nand UO_379 (O_379,N_9967,N_9814);
and UO_380 (O_380,N_9939,N_9815);
nand UO_381 (O_381,N_9814,N_9842);
and UO_382 (O_382,N_9852,N_9800);
nor UO_383 (O_383,N_9966,N_9969);
nor UO_384 (O_384,N_9993,N_9936);
nand UO_385 (O_385,N_9807,N_9993);
nand UO_386 (O_386,N_9943,N_9857);
nand UO_387 (O_387,N_9901,N_9834);
and UO_388 (O_388,N_9867,N_9849);
or UO_389 (O_389,N_9862,N_9852);
or UO_390 (O_390,N_9950,N_9878);
nand UO_391 (O_391,N_9953,N_9951);
nor UO_392 (O_392,N_9831,N_9851);
nor UO_393 (O_393,N_9827,N_9880);
nand UO_394 (O_394,N_9983,N_9978);
nand UO_395 (O_395,N_9879,N_9957);
or UO_396 (O_396,N_9913,N_9813);
nand UO_397 (O_397,N_9858,N_9865);
and UO_398 (O_398,N_9925,N_9849);
nor UO_399 (O_399,N_9996,N_9865);
nor UO_400 (O_400,N_9999,N_9803);
nand UO_401 (O_401,N_9837,N_9815);
xor UO_402 (O_402,N_9933,N_9839);
nand UO_403 (O_403,N_9972,N_9884);
and UO_404 (O_404,N_9928,N_9932);
nor UO_405 (O_405,N_9892,N_9904);
nor UO_406 (O_406,N_9804,N_9907);
nand UO_407 (O_407,N_9872,N_9844);
or UO_408 (O_408,N_9944,N_9880);
nor UO_409 (O_409,N_9952,N_9945);
nor UO_410 (O_410,N_9904,N_9884);
nand UO_411 (O_411,N_9941,N_9904);
nor UO_412 (O_412,N_9904,N_9902);
nor UO_413 (O_413,N_9810,N_9972);
or UO_414 (O_414,N_9827,N_9956);
nand UO_415 (O_415,N_9912,N_9801);
nor UO_416 (O_416,N_9846,N_9927);
or UO_417 (O_417,N_9812,N_9955);
nand UO_418 (O_418,N_9995,N_9863);
or UO_419 (O_419,N_9877,N_9938);
nor UO_420 (O_420,N_9984,N_9815);
nand UO_421 (O_421,N_9936,N_9860);
and UO_422 (O_422,N_9953,N_9800);
nand UO_423 (O_423,N_9879,N_9950);
nor UO_424 (O_424,N_9946,N_9958);
and UO_425 (O_425,N_9964,N_9886);
nand UO_426 (O_426,N_9979,N_9983);
nor UO_427 (O_427,N_9901,N_9804);
nor UO_428 (O_428,N_9868,N_9802);
or UO_429 (O_429,N_9840,N_9948);
and UO_430 (O_430,N_9963,N_9993);
xor UO_431 (O_431,N_9996,N_9965);
nand UO_432 (O_432,N_9941,N_9919);
or UO_433 (O_433,N_9887,N_9928);
nor UO_434 (O_434,N_9976,N_9859);
and UO_435 (O_435,N_9935,N_9814);
and UO_436 (O_436,N_9961,N_9965);
nand UO_437 (O_437,N_9807,N_9986);
or UO_438 (O_438,N_9975,N_9986);
nor UO_439 (O_439,N_9948,N_9874);
and UO_440 (O_440,N_9885,N_9976);
and UO_441 (O_441,N_9876,N_9877);
and UO_442 (O_442,N_9976,N_9947);
or UO_443 (O_443,N_9983,N_9987);
nand UO_444 (O_444,N_9844,N_9830);
or UO_445 (O_445,N_9881,N_9843);
and UO_446 (O_446,N_9934,N_9839);
or UO_447 (O_447,N_9955,N_9932);
nand UO_448 (O_448,N_9895,N_9887);
or UO_449 (O_449,N_9967,N_9977);
nor UO_450 (O_450,N_9830,N_9882);
nor UO_451 (O_451,N_9904,N_9995);
and UO_452 (O_452,N_9957,N_9848);
or UO_453 (O_453,N_9991,N_9888);
or UO_454 (O_454,N_9804,N_9952);
nand UO_455 (O_455,N_9976,N_9806);
nor UO_456 (O_456,N_9824,N_9967);
or UO_457 (O_457,N_9988,N_9821);
and UO_458 (O_458,N_9841,N_9825);
or UO_459 (O_459,N_9979,N_9997);
nand UO_460 (O_460,N_9915,N_9961);
nand UO_461 (O_461,N_9812,N_9948);
nand UO_462 (O_462,N_9896,N_9944);
nor UO_463 (O_463,N_9803,N_9862);
nor UO_464 (O_464,N_9984,N_9854);
or UO_465 (O_465,N_9850,N_9980);
and UO_466 (O_466,N_9812,N_9801);
and UO_467 (O_467,N_9811,N_9890);
nand UO_468 (O_468,N_9931,N_9921);
and UO_469 (O_469,N_9964,N_9896);
nor UO_470 (O_470,N_9851,N_9934);
or UO_471 (O_471,N_9813,N_9945);
nand UO_472 (O_472,N_9965,N_9867);
nand UO_473 (O_473,N_9815,N_9875);
and UO_474 (O_474,N_9885,N_9864);
or UO_475 (O_475,N_9893,N_9874);
and UO_476 (O_476,N_9872,N_9848);
nand UO_477 (O_477,N_9991,N_9864);
nand UO_478 (O_478,N_9801,N_9904);
nand UO_479 (O_479,N_9862,N_9843);
nor UO_480 (O_480,N_9920,N_9880);
or UO_481 (O_481,N_9974,N_9877);
nor UO_482 (O_482,N_9856,N_9806);
or UO_483 (O_483,N_9836,N_9883);
and UO_484 (O_484,N_9886,N_9955);
or UO_485 (O_485,N_9823,N_9923);
nor UO_486 (O_486,N_9859,N_9973);
and UO_487 (O_487,N_9999,N_9947);
or UO_488 (O_488,N_9824,N_9955);
and UO_489 (O_489,N_9966,N_9927);
or UO_490 (O_490,N_9944,N_9876);
and UO_491 (O_491,N_9847,N_9886);
and UO_492 (O_492,N_9988,N_9860);
and UO_493 (O_493,N_9994,N_9870);
nand UO_494 (O_494,N_9988,N_9986);
nor UO_495 (O_495,N_9837,N_9992);
and UO_496 (O_496,N_9970,N_9818);
nor UO_497 (O_497,N_9910,N_9802);
or UO_498 (O_498,N_9872,N_9822);
or UO_499 (O_499,N_9820,N_9979);
or UO_500 (O_500,N_9928,N_9870);
nor UO_501 (O_501,N_9941,N_9979);
nand UO_502 (O_502,N_9895,N_9973);
nand UO_503 (O_503,N_9927,N_9972);
or UO_504 (O_504,N_9924,N_9862);
or UO_505 (O_505,N_9858,N_9956);
nor UO_506 (O_506,N_9835,N_9937);
and UO_507 (O_507,N_9876,N_9963);
nor UO_508 (O_508,N_9839,N_9996);
and UO_509 (O_509,N_9890,N_9917);
and UO_510 (O_510,N_9980,N_9987);
and UO_511 (O_511,N_9820,N_9920);
and UO_512 (O_512,N_9899,N_9836);
nand UO_513 (O_513,N_9943,N_9854);
nor UO_514 (O_514,N_9858,N_9840);
nand UO_515 (O_515,N_9905,N_9800);
nand UO_516 (O_516,N_9874,N_9818);
and UO_517 (O_517,N_9815,N_9969);
and UO_518 (O_518,N_9930,N_9882);
or UO_519 (O_519,N_9825,N_9990);
and UO_520 (O_520,N_9825,N_9840);
nor UO_521 (O_521,N_9853,N_9921);
and UO_522 (O_522,N_9874,N_9814);
nor UO_523 (O_523,N_9811,N_9873);
or UO_524 (O_524,N_9897,N_9816);
and UO_525 (O_525,N_9935,N_9865);
or UO_526 (O_526,N_9845,N_9871);
nor UO_527 (O_527,N_9979,N_9819);
nor UO_528 (O_528,N_9863,N_9909);
nand UO_529 (O_529,N_9818,N_9873);
or UO_530 (O_530,N_9855,N_9897);
and UO_531 (O_531,N_9907,N_9802);
or UO_532 (O_532,N_9971,N_9937);
nor UO_533 (O_533,N_9910,N_9889);
nand UO_534 (O_534,N_9806,N_9958);
or UO_535 (O_535,N_9922,N_9848);
nor UO_536 (O_536,N_9931,N_9967);
nand UO_537 (O_537,N_9822,N_9813);
or UO_538 (O_538,N_9861,N_9851);
or UO_539 (O_539,N_9864,N_9953);
or UO_540 (O_540,N_9954,N_9867);
or UO_541 (O_541,N_9925,N_9873);
xor UO_542 (O_542,N_9889,N_9843);
and UO_543 (O_543,N_9910,N_9977);
and UO_544 (O_544,N_9885,N_9968);
nor UO_545 (O_545,N_9906,N_9802);
or UO_546 (O_546,N_9915,N_9863);
and UO_547 (O_547,N_9814,N_9950);
nand UO_548 (O_548,N_9980,N_9943);
and UO_549 (O_549,N_9886,N_9827);
nand UO_550 (O_550,N_9931,N_9862);
or UO_551 (O_551,N_9971,N_9895);
or UO_552 (O_552,N_9960,N_9851);
nand UO_553 (O_553,N_9828,N_9890);
and UO_554 (O_554,N_9968,N_9814);
nand UO_555 (O_555,N_9979,N_9937);
or UO_556 (O_556,N_9830,N_9868);
and UO_557 (O_557,N_9828,N_9910);
and UO_558 (O_558,N_9842,N_9990);
or UO_559 (O_559,N_9934,N_9885);
or UO_560 (O_560,N_9869,N_9909);
nand UO_561 (O_561,N_9978,N_9962);
or UO_562 (O_562,N_9909,N_9801);
or UO_563 (O_563,N_9993,N_9846);
nor UO_564 (O_564,N_9966,N_9844);
or UO_565 (O_565,N_9876,N_9905);
or UO_566 (O_566,N_9839,N_9939);
nand UO_567 (O_567,N_9991,N_9940);
nand UO_568 (O_568,N_9976,N_9939);
and UO_569 (O_569,N_9974,N_9828);
and UO_570 (O_570,N_9855,N_9875);
or UO_571 (O_571,N_9857,N_9904);
or UO_572 (O_572,N_9925,N_9995);
nand UO_573 (O_573,N_9972,N_9943);
nor UO_574 (O_574,N_9876,N_9860);
and UO_575 (O_575,N_9916,N_9832);
and UO_576 (O_576,N_9966,N_9899);
nor UO_577 (O_577,N_9981,N_9819);
and UO_578 (O_578,N_9956,N_9885);
nand UO_579 (O_579,N_9847,N_9869);
and UO_580 (O_580,N_9935,N_9937);
or UO_581 (O_581,N_9955,N_9860);
and UO_582 (O_582,N_9943,N_9832);
nand UO_583 (O_583,N_9927,N_9823);
or UO_584 (O_584,N_9801,N_9838);
nor UO_585 (O_585,N_9937,N_9826);
and UO_586 (O_586,N_9854,N_9977);
or UO_587 (O_587,N_9848,N_9871);
and UO_588 (O_588,N_9994,N_9859);
or UO_589 (O_589,N_9864,N_9809);
and UO_590 (O_590,N_9804,N_9823);
and UO_591 (O_591,N_9843,N_9863);
nand UO_592 (O_592,N_9870,N_9933);
nor UO_593 (O_593,N_9851,N_9864);
and UO_594 (O_594,N_9928,N_9993);
and UO_595 (O_595,N_9880,N_9854);
nand UO_596 (O_596,N_9978,N_9884);
nand UO_597 (O_597,N_9819,N_9923);
nor UO_598 (O_598,N_9942,N_9833);
and UO_599 (O_599,N_9989,N_9979);
nand UO_600 (O_600,N_9961,N_9955);
or UO_601 (O_601,N_9975,N_9943);
nor UO_602 (O_602,N_9877,N_9996);
or UO_603 (O_603,N_9845,N_9811);
nor UO_604 (O_604,N_9917,N_9993);
nor UO_605 (O_605,N_9939,N_9966);
or UO_606 (O_606,N_9878,N_9830);
nand UO_607 (O_607,N_9892,N_9995);
nor UO_608 (O_608,N_9828,N_9839);
nor UO_609 (O_609,N_9884,N_9922);
nor UO_610 (O_610,N_9924,N_9813);
and UO_611 (O_611,N_9803,N_9871);
nor UO_612 (O_612,N_9885,N_9906);
or UO_613 (O_613,N_9824,N_9880);
and UO_614 (O_614,N_9914,N_9896);
nand UO_615 (O_615,N_9821,N_9939);
and UO_616 (O_616,N_9849,N_9836);
nand UO_617 (O_617,N_9912,N_9895);
nand UO_618 (O_618,N_9926,N_9939);
nand UO_619 (O_619,N_9914,N_9988);
and UO_620 (O_620,N_9965,N_9805);
nand UO_621 (O_621,N_9953,N_9874);
nand UO_622 (O_622,N_9946,N_9871);
or UO_623 (O_623,N_9822,N_9866);
and UO_624 (O_624,N_9830,N_9970);
nand UO_625 (O_625,N_9912,N_9903);
nor UO_626 (O_626,N_9966,N_9848);
nor UO_627 (O_627,N_9915,N_9919);
nor UO_628 (O_628,N_9949,N_9925);
and UO_629 (O_629,N_9801,N_9949);
or UO_630 (O_630,N_9831,N_9956);
nand UO_631 (O_631,N_9966,N_9929);
nand UO_632 (O_632,N_9853,N_9897);
nand UO_633 (O_633,N_9839,N_9884);
nand UO_634 (O_634,N_9811,N_9922);
and UO_635 (O_635,N_9814,N_9838);
nor UO_636 (O_636,N_9928,N_9823);
and UO_637 (O_637,N_9873,N_9858);
nand UO_638 (O_638,N_9847,N_9894);
nand UO_639 (O_639,N_9917,N_9885);
nor UO_640 (O_640,N_9983,N_9810);
and UO_641 (O_641,N_9948,N_9809);
nand UO_642 (O_642,N_9850,N_9899);
and UO_643 (O_643,N_9805,N_9913);
nand UO_644 (O_644,N_9807,N_9846);
nand UO_645 (O_645,N_9913,N_9832);
xnor UO_646 (O_646,N_9975,N_9961);
and UO_647 (O_647,N_9863,N_9969);
and UO_648 (O_648,N_9961,N_9884);
or UO_649 (O_649,N_9810,N_9998);
and UO_650 (O_650,N_9874,N_9882);
nor UO_651 (O_651,N_9821,N_9850);
nand UO_652 (O_652,N_9982,N_9840);
or UO_653 (O_653,N_9993,N_9982);
nand UO_654 (O_654,N_9918,N_9988);
and UO_655 (O_655,N_9928,N_9863);
nand UO_656 (O_656,N_9801,N_9887);
nand UO_657 (O_657,N_9894,N_9903);
nand UO_658 (O_658,N_9845,N_9989);
and UO_659 (O_659,N_9848,N_9986);
nand UO_660 (O_660,N_9970,N_9853);
or UO_661 (O_661,N_9930,N_9920);
nand UO_662 (O_662,N_9893,N_9909);
nand UO_663 (O_663,N_9974,N_9919);
xor UO_664 (O_664,N_9818,N_9884);
nand UO_665 (O_665,N_9999,N_9989);
xor UO_666 (O_666,N_9824,N_9988);
and UO_667 (O_667,N_9808,N_9971);
nor UO_668 (O_668,N_9876,N_9929);
nor UO_669 (O_669,N_9880,N_9863);
nand UO_670 (O_670,N_9995,N_9843);
nor UO_671 (O_671,N_9853,N_9834);
or UO_672 (O_672,N_9922,N_9914);
or UO_673 (O_673,N_9937,N_9965);
or UO_674 (O_674,N_9906,N_9886);
and UO_675 (O_675,N_9810,N_9966);
or UO_676 (O_676,N_9813,N_9847);
nor UO_677 (O_677,N_9807,N_9851);
and UO_678 (O_678,N_9902,N_9833);
or UO_679 (O_679,N_9917,N_9824);
and UO_680 (O_680,N_9850,N_9920);
nand UO_681 (O_681,N_9943,N_9996);
or UO_682 (O_682,N_9988,N_9999);
nor UO_683 (O_683,N_9848,N_9879);
nand UO_684 (O_684,N_9898,N_9917);
nand UO_685 (O_685,N_9909,N_9971);
or UO_686 (O_686,N_9963,N_9858);
and UO_687 (O_687,N_9872,N_9907);
or UO_688 (O_688,N_9943,N_9954);
nor UO_689 (O_689,N_9864,N_9929);
nor UO_690 (O_690,N_9905,N_9959);
or UO_691 (O_691,N_9940,N_9899);
or UO_692 (O_692,N_9933,N_9944);
nand UO_693 (O_693,N_9928,N_9977);
or UO_694 (O_694,N_9999,N_9969);
or UO_695 (O_695,N_9882,N_9923);
or UO_696 (O_696,N_9920,N_9862);
and UO_697 (O_697,N_9940,N_9903);
and UO_698 (O_698,N_9888,N_9843);
nor UO_699 (O_699,N_9842,N_9999);
and UO_700 (O_700,N_9869,N_9965);
nand UO_701 (O_701,N_9806,N_9986);
nand UO_702 (O_702,N_9969,N_9852);
or UO_703 (O_703,N_9853,N_9939);
nor UO_704 (O_704,N_9987,N_9931);
and UO_705 (O_705,N_9930,N_9892);
nor UO_706 (O_706,N_9921,N_9827);
and UO_707 (O_707,N_9911,N_9899);
and UO_708 (O_708,N_9867,N_9848);
and UO_709 (O_709,N_9974,N_9800);
nand UO_710 (O_710,N_9881,N_9951);
or UO_711 (O_711,N_9963,N_9891);
or UO_712 (O_712,N_9899,N_9982);
and UO_713 (O_713,N_9915,N_9921);
nor UO_714 (O_714,N_9911,N_9892);
and UO_715 (O_715,N_9983,N_9881);
or UO_716 (O_716,N_9816,N_9871);
nor UO_717 (O_717,N_9971,N_9941);
nand UO_718 (O_718,N_9884,N_9840);
or UO_719 (O_719,N_9891,N_9985);
and UO_720 (O_720,N_9902,N_9989);
or UO_721 (O_721,N_9930,N_9932);
and UO_722 (O_722,N_9891,N_9862);
and UO_723 (O_723,N_9952,N_9856);
nand UO_724 (O_724,N_9919,N_9972);
nor UO_725 (O_725,N_9869,N_9837);
and UO_726 (O_726,N_9946,N_9898);
nand UO_727 (O_727,N_9803,N_9812);
nand UO_728 (O_728,N_9948,N_9868);
nor UO_729 (O_729,N_9965,N_9854);
or UO_730 (O_730,N_9867,N_9884);
nand UO_731 (O_731,N_9813,N_9997);
or UO_732 (O_732,N_9901,N_9963);
nor UO_733 (O_733,N_9884,N_9852);
nor UO_734 (O_734,N_9944,N_9860);
or UO_735 (O_735,N_9914,N_9931);
nor UO_736 (O_736,N_9820,N_9854);
nor UO_737 (O_737,N_9876,N_9850);
nand UO_738 (O_738,N_9934,N_9918);
nand UO_739 (O_739,N_9819,N_9858);
or UO_740 (O_740,N_9971,N_9876);
and UO_741 (O_741,N_9860,N_9808);
nand UO_742 (O_742,N_9919,N_9932);
nand UO_743 (O_743,N_9937,N_9972);
and UO_744 (O_744,N_9928,N_9983);
nor UO_745 (O_745,N_9943,N_9947);
and UO_746 (O_746,N_9844,N_9867);
nor UO_747 (O_747,N_9847,N_9818);
and UO_748 (O_748,N_9967,N_9846);
nand UO_749 (O_749,N_9893,N_9962);
and UO_750 (O_750,N_9844,N_9904);
nor UO_751 (O_751,N_9980,N_9936);
nand UO_752 (O_752,N_9867,N_9983);
xor UO_753 (O_753,N_9838,N_9954);
nand UO_754 (O_754,N_9975,N_9947);
nor UO_755 (O_755,N_9981,N_9909);
or UO_756 (O_756,N_9837,N_9982);
or UO_757 (O_757,N_9958,N_9998);
nor UO_758 (O_758,N_9844,N_9932);
or UO_759 (O_759,N_9855,N_9953);
and UO_760 (O_760,N_9845,N_9893);
nor UO_761 (O_761,N_9873,N_9935);
nand UO_762 (O_762,N_9939,N_9827);
nor UO_763 (O_763,N_9835,N_9970);
nor UO_764 (O_764,N_9991,N_9819);
nor UO_765 (O_765,N_9951,N_9880);
xnor UO_766 (O_766,N_9939,N_9808);
and UO_767 (O_767,N_9805,N_9891);
xnor UO_768 (O_768,N_9933,N_9811);
nand UO_769 (O_769,N_9802,N_9843);
nor UO_770 (O_770,N_9941,N_9913);
and UO_771 (O_771,N_9924,N_9964);
xnor UO_772 (O_772,N_9960,N_9903);
and UO_773 (O_773,N_9810,N_9890);
or UO_774 (O_774,N_9884,N_9992);
and UO_775 (O_775,N_9812,N_9977);
and UO_776 (O_776,N_9841,N_9956);
and UO_777 (O_777,N_9882,N_9960);
nand UO_778 (O_778,N_9954,N_9802);
nor UO_779 (O_779,N_9928,N_9851);
nor UO_780 (O_780,N_9857,N_9898);
or UO_781 (O_781,N_9957,N_9868);
nor UO_782 (O_782,N_9840,N_9817);
or UO_783 (O_783,N_9915,N_9916);
nand UO_784 (O_784,N_9965,N_9896);
nor UO_785 (O_785,N_9906,N_9914);
nand UO_786 (O_786,N_9850,N_9834);
nand UO_787 (O_787,N_9849,N_9942);
and UO_788 (O_788,N_9945,N_9911);
nand UO_789 (O_789,N_9843,N_9904);
nand UO_790 (O_790,N_9974,N_9898);
or UO_791 (O_791,N_9804,N_9994);
nor UO_792 (O_792,N_9926,N_9958);
or UO_793 (O_793,N_9994,N_9968);
or UO_794 (O_794,N_9827,N_9903);
nor UO_795 (O_795,N_9844,N_9979);
nand UO_796 (O_796,N_9962,N_9857);
and UO_797 (O_797,N_9855,N_9854);
nand UO_798 (O_798,N_9893,N_9965);
or UO_799 (O_799,N_9906,N_9949);
nand UO_800 (O_800,N_9988,N_9974);
and UO_801 (O_801,N_9946,N_9889);
nor UO_802 (O_802,N_9928,N_9883);
nor UO_803 (O_803,N_9947,N_9894);
nand UO_804 (O_804,N_9878,N_9920);
nand UO_805 (O_805,N_9868,N_9866);
nor UO_806 (O_806,N_9836,N_9920);
or UO_807 (O_807,N_9973,N_9821);
and UO_808 (O_808,N_9854,N_9832);
and UO_809 (O_809,N_9850,N_9822);
or UO_810 (O_810,N_9841,N_9947);
and UO_811 (O_811,N_9946,N_9882);
nand UO_812 (O_812,N_9859,N_9933);
nor UO_813 (O_813,N_9994,N_9815);
nor UO_814 (O_814,N_9916,N_9971);
nand UO_815 (O_815,N_9934,N_9900);
nor UO_816 (O_816,N_9810,N_9948);
or UO_817 (O_817,N_9953,N_9823);
nor UO_818 (O_818,N_9975,N_9899);
or UO_819 (O_819,N_9862,N_9828);
nand UO_820 (O_820,N_9809,N_9813);
or UO_821 (O_821,N_9880,N_9971);
nor UO_822 (O_822,N_9809,N_9978);
or UO_823 (O_823,N_9870,N_9905);
nor UO_824 (O_824,N_9983,N_9839);
nor UO_825 (O_825,N_9906,N_9974);
or UO_826 (O_826,N_9873,N_9830);
nand UO_827 (O_827,N_9820,N_9814);
nand UO_828 (O_828,N_9922,N_9925);
and UO_829 (O_829,N_9858,N_9829);
nor UO_830 (O_830,N_9820,N_9952);
and UO_831 (O_831,N_9937,N_9973);
and UO_832 (O_832,N_9863,N_9959);
or UO_833 (O_833,N_9877,N_9862);
or UO_834 (O_834,N_9965,N_9897);
nand UO_835 (O_835,N_9906,N_9956);
nand UO_836 (O_836,N_9913,N_9909);
and UO_837 (O_837,N_9999,N_9923);
and UO_838 (O_838,N_9922,N_9955);
and UO_839 (O_839,N_9914,N_9817);
or UO_840 (O_840,N_9803,N_9980);
or UO_841 (O_841,N_9863,N_9954);
or UO_842 (O_842,N_9865,N_9801);
or UO_843 (O_843,N_9917,N_9940);
nor UO_844 (O_844,N_9885,N_9805);
nor UO_845 (O_845,N_9932,N_9965);
or UO_846 (O_846,N_9932,N_9964);
nor UO_847 (O_847,N_9956,N_9961);
nor UO_848 (O_848,N_9817,N_9800);
and UO_849 (O_849,N_9839,N_9844);
nor UO_850 (O_850,N_9806,N_9801);
or UO_851 (O_851,N_9990,N_9973);
nor UO_852 (O_852,N_9920,N_9807);
nor UO_853 (O_853,N_9929,N_9988);
or UO_854 (O_854,N_9860,N_9962);
nor UO_855 (O_855,N_9902,N_9823);
or UO_856 (O_856,N_9878,N_9912);
nor UO_857 (O_857,N_9834,N_9848);
nand UO_858 (O_858,N_9835,N_9892);
or UO_859 (O_859,N_9911,N_9816);
nand UO_860 (O_860,N_9847,N_9889);
nor UO_861 (O_861,N_9885,N_9875);
xnor UO_862 (O_862,N_9868,N_9880);
nor UO_863 (O_863,N_9885,N_9960);
nor UO_864 (O_864,N_9928,N_9834);
nor UO_865 (O_865,N_9899,N_9984);
nor UO_866 (O_866,N_9980,N_9820);
or UO_867 (O_867,N_9987,N_9902);
nand UO_868 (O_868,N_9964,N_9966);
or UO_869 (O_869,N_9927,N_9877);
or UO_870 (O_870,N_9843,N_9822);
or UO_871 (O_871,N_9959,N_9897);
and UO_872 (O_872,N_9901,N_9805);
and UO_873 (O_873,N_9986,N_9882);
and UO_874 (O_874,N_9993,N_9981);
nand UO_875 (O_875,N_9920,N_9969);
or UO_876 (O_876,N_9899,N_9964);
and UO_877 (O_877,N_9998,N_9884);
or UO_878 (O_878,N_9815,N_9895);
or UO_879 (O_879,N_9804,N_9879);
nor UO_880 (O_880,N_9838,N_9897);
or UO_881 (O_881,N_9907,N_9948);
nor UO_882 (O_882,N_9820,N_9812);
or UO_883 (O_883,N_9818,N_9877);
or UO_884 (O_884,N_9828,N_9858);
and UO_885 (O_885,N_9926,N_9869);
nor UO_886 (O_886,N_9976,N_9952);
nor UO_887 (O_887,N_9829,N_9992);
nand UO_888 (O_888,N_9879,N_9803);
nor UO_889 (O_889,N_9985,N_9977);
nor UO_890 (O_890,N_9834,N_9856);
or UO_891 (O_891,N_9801,N_9952);
and UO_892 (O_892,N_9995,N_9910);
nand UO_893 (O_893,N_9964,N_9889);
nor UO_894 (O_894,N_9893,N_9905);
or UO_895 (O_895,N_9940,N_9876);
or UO_896 (O_896,N_9932,N_9835);
nor UO_897 (O_897,N_9894,N_9887);
or UO_898 (O_898,N_9876,N_9990);
nand UO_899 (O_899,N_9986,N_9907);
nor UO_900 (O_900,N_9939,N_9902);
nand UO_901 (O_901,N_9923,N_9871);
nand UO_902 (O_902,N_9969,N_9990);
xor UO_903 (O_903,N_9917,N_9923);
and UO_904 (O_904,N_9845,N_9904);
nor UO_905 (O_905,N_9936,N_9931);
nand UO_906 (O_906,N_9948,N_9848);
nand UO_907 (O_907,N_9902,N_9997);
nand UO_908 (O_908,N_9946,N_9956);
nand UO_909 (O_909,N_9985,N_9958);
nand UO_910 (O_910,N_9881,N_9865);
nand UO_911 (O_911,N_9827,N_9801);
nor UO_912 (O_912,N_9941,N_9826);
nand UO_913 (O_913,N_9973,N_9823);
or UO_914 (O_914,N_9878,N_9921);
or UO_915 (O_915,N_9957,N_9920);
nand UO_916 (O_916,N_9895,N_9914);
nand UO_917 (O_917,N_9999,N_9950);
nand UO_918 (O_918,N_9825,N_9944);
nor UO_919 (O_919,N_9892,N_9900);
and UO_920 (O_920,N_9999,N_9807);
and UO_921 (O_921,N_9910,N_9902);
nand UO_922 (O_922,N_9875,N_9874);
and UO_923 (O_923,N_9937,N_9913);
or UO_924 (O_924,N_9957,N_9910);
or UO_925 (O_925,N_9927,N_9851);
and UO_926 (O_926,N_9930,N_9980);
or UO_927 (O_927,N_9803,N_9815);
nor UO_928 (O_928,N_9984,N_9875);
and UO_929 (O_929,N_9980,N_9988);
or UO_930 (O_930,N_9807,N_9972);
nand UO_931 (O_931,N_9955,N_9889);
and UO_932 (O_932,N_9954,N_9887);
or UO_933 (O_933,N_9995,N_9965);
nor UO_934 (O_934,N_9989,N_9858);
nor UO_935 (O_935,N_9913,N_9929);
and UO_936 (O_936,N_9992,N_9849);
nand UO_937 (O_937,N_9822,N_9879);
or UO_938 (O_938,N_9828,N_9855);
nand UO_939 (O_939,N_9914,N_9879);
nand UO_940 (O_940,N_9947,N_9832);
nand UO_941 (O_941,N_9947,N_9823);
or UO_942 (O_942,N_9990,N_9968);
nand UO_943 (O_943,N_9832,N_9871);
nor UO_944 (O_944,N_9819,N_9940);
and UO_945 (O_945,N_9871,N_9807);
and UO_946 (O_946,N_9871,N_9918);
or UO_947 (O_947,N_9872,N_9985);
nand UO_948 (O_948,N_9849,N_9900);
nor UO_949 (O_949,N_9826,N_9938);
or UO_950 (O_950,N_9959,N_9926);
or UO_951 (O_951,N_9808,N_9946);
or UO_952 (O_952,N_9923,N_9988);
or UO_953 (O_953,N_9979,N_9894);
and UO_954 (O_954,N_9846,N_9969);
and UO_955 (O_955,N_9871,N_9986);
or UO_956 (O_956,N_9848,N_9817);
and UO_957 (O_957,N_9979,N_9947);
nor UO_958 (O_958,N_9998,N_9987);
and UO_959 (O_959,N_9902,N_9819);
or UO_960 (O_960,N_9801,N_9853);
nor UO_961 (O_961,N_9802,N_9818);
nand UO_962 (O_962,N_9905,N_9929);
nor UO_963 (O_963,N_9885,N_9838);
and UO_964 (O_964,N_9968,N_9807);
or UO_965 (O_965,N_9961,N_9929);
nand UO_966 (O_966,N_9910,N_9960);
or UO_967 (O_967,N_9884,N_9999);
nand UO_968 (O_968,N_9851,N_9946);
or UO_969 (O_969,N_9825,N_9812);
nand UO_970 (O_970,N_9904,N_9806);
or UO_971 (O_971,N_9811,N_9816);
nand UO_972 (O_972,N_9983,N_9925);
nand UO_973 (O_973,N_9902,N_9953);
and UO_974 (O_974,N_9862,N_9965);
or UO_975 (O_975,N_9860,N_9963);
and UO_976 (O_976,N_9838,N_9999);
nand UO_977 (O_977,N_9931,N_9844);
and UO_978 (O_978,N_9912,N_9899);
or UO_979 (O_979,N_9953,N_9968);
nand UO_980 (O_980,N_9938,N_9895);
and UO_981 (O_981,N_9864,N_9985);
or UO_982 (O_982,N_9905,N_9845);
and UO_983 (O_983,N_9989,N_9915);
and UO_984 (O_984,N_9987,N_9972);
nor UO_985 (O_985,N_9933,N_9848);
or UO_986 (O_986,N_9942,N_9924);
nor UO_987 (O_987,N_9838,N_9886);
xor UO_988 (O_988,N_9810,N_9931);
nor UO_989 (O_989,N_9934,N_9814);
nand UO_990 (O_990,N_9895,N_9861);
nand UO_991 (O_991,N_9802,N_9865);
nand UO_992 (O_992,N_9859,N_9834);
nand UO_993 (O_993,N_9913,N_9833);
nand UO_994 (O_994,N_9968,N_9972);
nand UO_995 (O_995,N_9932,N_9876);
nor UO_996 (O_996,N_9873,N_9967);
or UO_997 (O_997,N_9946,N_9822);
nor UO_998 (O_998,N_9907,N_9998);
xnor UO_999 (O_999,N_9842,N_9963);
or UO_1000 (O_1000,N_9892,N_9814);
nor UO_1001 (O_1001,N_9894,N_9962);
nand UO_1002 (O_1002,N_9989,N_9885);
nor UO_1003 (O_1003,N_9955,N_9876);
and UO_1004 (O_1004,N_9887,N_9983);
or UO_1005 (O_1005,N_9865,N_9910);
nor UO_1006 (O_1006,N_9853,N_9847);
nand UO_1007 (O_1007,N_9818,N_9858);
or UO_1008 (O_1008,N_9855,N_9961);
nor UO_1009 (O_1009,N_9894,N_9954);
nor UO_1010 (O_1010,N_9870,N_9966);
nor UO_1011 (O_1011,N_9983,N_9954);
nand UO_1012 (O_1012,N_9952,N_9835);
and UO_1013 (O_1013,N_9845,N_9960);
nor UO_1014 (O_1014,N_9830,N_9807);
nand UO_1015 (O_1015,N_9804,N_9870);
or UO_1016 (O_1016,N_9949,N_9812);
nand UO_1017 (O_1017,N_9879,N_9933);
or UO_1018 (O_1018,N_9910,N_9843);
xnor UO_1019 (O_1019,N_9807,N_9849);
and UO_1020 (O_1020,N_9848,N_9944);
or UO_1021 (O_1021,N_9985,N_9970);
or UO_1022 (O_1022,N_9852,N_9922);
or UO_1023 (O_1023,N_9850,N_9944);
nor UO_1024 (O_1024,N_9840,N_9952);
nand UO_1025 (O_1025,N_9982,N_9828);
nor UO_1026 (O_1026,N_9885,N_9831);
nor UO_1027 (O_1027,N_9946,N_9913);
nand UO_1028 (O_1028,N_9842,N_9994);
nand UO_1029 (O_1029,N_9957,N_9918);
nand UO_1030 (O_1030,N_9821,N_9979);
nand UO_1031 (O_1031,N_9806,N_9893);
or UO_1032 (O_1032,N_9856,N_9888);
nand UO_1033 (O_1033,N_9810,N_9829);
or UO_1034 (O_1034,N_9957,N_9937);
and UO_1035 (O_1035,N_9913,N_9839);
or UO_1036 (O_1036,N_9840,N_9875);
nor UO_1037 (O_1037,N_9854,N_9954);
or UO_1038 (O_1038,N_9808,N_9835);
nand UO_1039 (O_1039,N_9912,N_9800);
and UO_1040 (O_1040,N_9831,N_9990);
and UO_1041 (O_1041,N_9955,N_9803);
and UO_1042 (O_1042,N_9810,N_9937);
nand UO_1043 (O_1043,N_9808,N_9979);
nor UO_1044 (O_1044,N_9873,N_9918);
nand UO_1045 (O_1045,N_9892,N_9885);
and UO_1046 (O_1046,N_9832,N_9902);
and UO_1047 (O_1047,N_9822,N_9951);
or UO_1048 (O_1048,N_9804,N_9848);
and UO_1049 (O_1049,N_9827,N_9908);
nand UO_1050 (O_1050,N_9800,N_9902);
or UO_1051 (O_1051,N_9985,N_9935);
nand UO_1052 (O_1052,N_9957,N_9933);
or UO_1053 (O_1053,N_9926,N_9843);
or UO_1054 (O_1054,N_9940,N_9829);
nand UO_1055 (O_1055,N_9864,N_9913);
nand UO_1056 (O_1056,N_9977,N_9966);
nor UO_1057 (O_1057,N_9987,N_9807);
or UO_1058 (O_1058,N_9880,N_9969);
or UO_1059 (O_1059,N_9935,N_9852);
or UO_1060 (O_1060,N_9912,N_9822);
or UO_1061 (O_1061,N_9922,N_9859);
and UO_1062 (O_1062,N_9952,N_9844);
nor UO_1063 (O_1063,N_9882,N_9906);
nor UO_1064 (O_1064,N_9868,N_9873);
nor UO_1065 (O_1065,N_9894,N_9897);
or UO_1066 (O_1066,N_9884,N_9849);
nor UO_1067 (O_1067,N_9951,N_9839);
nand UO_1068 (O_1068,N_9833,N_9882);
or UO_1069 (O_1069,N_9854,N_9945);
and UO_1070 (O_1070,N_9919,N_9877);
nand UO_1071 (O_1071,N_9804,N_9955);
and UO_1072 (O_1072,N_9954,N_9912);
nor UO_1073 (O_1073,N_9929,N_9889);
and UO_1074 (O_1074,N_9806,N_9857);
nand UO_1075 (O_1075,N_9845,N_9943);
nand UO_1076 (O_1076,N_9850,N_9893);
nand UO_1077 (O_1077,N_9938,N_9841);
nand UO_1078 (O_1078,N_9995,N_9987);
and UO_1079 (O_1079,N_9912,N_9917);
or UO_1080 (O_1080,N_9856,N_9828);
or UO_1081 (O_1081,N_9888,N_9975);
nand UO_1082 (O_1082,N_9925,N_9816);
and UO_1083 (O_1083,N_9879,N_9840);
or UO_1084 (O_1084,N_9967,N_9882);
or UO_1085 (O_1085,N_9909,N_9933);
and UO_1086 (O_1086,N_9979,N_9960);
or UO_1087 (O_1087,N_9987,N_9919);
or UO_1088 (O_1088,N_9934,N_9957);
and UO_1089 (O_1089,N_9882,N_9994);
and UO_1090 (O_1090,N_9912,N_9970);
or UO_1091 (O_1091,N_9875,N_9995);
nor UO_1092 (O_1092,N_9853,N_9854);
nand UO_1093 (O_1093,N_9936,N_9821);
nor UO_1094 (O_1094,N_9869,N_9961);
nor UO_1095 (O_1095,N_9991,N_9810);
nor UO_1096 (O_1096,N_9868,N_9814);
or UO_1097 (O_1097,N_9910,N_9929);
or UO_1098 (O_1098,N_9809,N_9831);
and UO_1099 (O_1099,N_9886,N_9967);
and UO_1100 (O_1100,N_9913,N_9991);
nand UO_1101 (O_1101,N_9950,N_9884);
nand UO_1102 (O_1102,N_9815,N_9841);
nor UO_1103 (O_1103,N_9997,N_9921);
nand UO_1104 (O_1104,N_9891,N_9907);
or UO_1105 (O_1105,N_9808,N_9845);
and UO_1106 (O_1106,N_9818,N_9890);
and UO_1107 (O_1107,N_9987,N_9992);
nor UO_1108 (O_1108,N_9905,N_9896);
nor UO_1109 (O_1109,N_9800,N_9973);
nor UO_1110 (O_1110,N_9851,N_9810);
or UO_1111 (O_1111,N_9997,N_9909);
nand UO_1112 (O_1112,N_9942,N_9905);
nor UO_1113 (O_1113,N_9816,N_9973);
nor UO_1114 (O_1114,N_9911,N_9805);
and UO_1115 (O_1115,N_9927,N_9825);
nor UO_1116 (O_1116,N_9923,N_9806);
nor UO_1117 (O_1117,N_9868,N_9944);
nor UO_1118 (O_1118,N_9895,N_9847);
or UO_1119 (O_1119,N_9959,N_9884);
nand UO_1120 (O_1120,N_9895,N_9954);
nor UO_1121 (O_1121,N_9883,N_9887);
and UO_1122 (O_1122,N_9829,N_9939);
nand UO_1123 (O_1123,N_9835,N_9985);
nor UO_1124 (O_1124,N_9887,N_9814);
nor UO_1125 (O_1125,N_9912,N_9846);
nand UO_1126 (O_1126,N_9921,N_9945);
nand UO_1127 (O_1127,N_9887,N_9997);
or UO_1128 (O_1128,N_9949,N_9860);
nor UO_1129 (O_1129,N_9945,N_9815);
nor UO_1130 (O_1130,N_9827,N_9948);
nand UO_1131 (O_1131,N_9849,N_9918);
nor UO_1132 (O_1132,N_9892,N_9937);
nor UO_1133 (O_1133,N_9852,N_9978);
and UO_1134 (O_1134,N_9984,N_9823);
nand UO_1135 (O_1135,N_9863,N_9941);
or UO_1136 (O_1136,N_9995,N_9977);
or UO_1137 (O_1137,N_9855,N_9951);
and UO_1138 (O_1138,N_9826,N_9843);
and UO_1139 (O_1139,N_9961,N_9983);
and UO_1140 (O_1140,N_9941,N_9800);
nand UO_1141 (O_1141,N_9908,N_9968);
nand UO_1142 (O_1142,N_9894,N_9963);
or UO_1143 (O_1143,N_9960,N_9805);
nor UO_1144 (O_1144,N_9980,N_9894);
and UO_1145 (O_1145,N_9863,N_9858);
and UO_1146 (O_1146,N_9815,N_9977);
nor UO_1147 (O_1147,N_9820,N_9971);
and UO_1148 (O_1148,N_9816,N_9858);
and UO_1149 (O_1149,N_9835,N_9967);
and UO_1150 (O_1150,N_9898,N_9805);
and UO_1151 (O_1151,N_9910,N_9832);
or UO_1152 (O_1152,N_9876,N_9816);
nand UO_1153 (O_1153,N_9813,N_9881);
nand UO_1154 (O_1154,N_9896,N_9865);
nand UO_1155 (O_1155,N_9823,N_9987);
and UO_1156 (O_1156,N_9985,N_9839);
nor UO_1157 (O_1157,N_9938,N_9823);
nor UO_1158 (O_1158,N_9838,N_9984);
or UO_1159 (O_1159,N_9835,N_9801);
or UO_1160 (O_1160,N_9942,N_9980);
nor UO_1161 (O_1161,N_9830,N_9879);
nand UO_1162 (O_1162,N_9998,N_9868);
nor UO_1163 (O_1163,N_9868,N_9829);
nor UO_1164 (O_1164,N_9872,N_9981);
nand UO_1165 (O_1165,N_9928,N_9921);
or UO_1166 (O_1166,N_9992,N_9936);
nand UO_1167 (O_1167,N_9839,N_9930);
or UO_1168 (O_1168,N_9906,N_9841);
and UO_1169 (O_1169,N_9889,N_9953);
xor UO_1170 (O_1170,N_9940,N_9885);
nand UO_1171 (O_1171,N_9997,N_9876);
nand UO_1172 (O_1172,N_9900,N_9846);
or UO_1173 (O_1173,N_9916,N_9887);
or UO_1174 (O_1174,N_9888,N_9832);
nand UO_1175 (O_1175,N_9985,N_9950);
or UO_1176 (O_1176,N_9943,N_9917);
nor UO_1177 (O_1177,N_9847,N_9810);
nor UO_1178 (O_1178,N_9924,N_9890);
nand UO_1179 (O_1179,N_9802,N_9886);
or UO_1180 (O_1180,N_9854,N_9857);
nand UO_1181 (O_1181,N_9837,N_9975);
nor UO_1182 (O_1182,N_9803,N_9971);
nand UO_1183 (O_1183,N_9890,N_9954);
and UO_1184 (O_1184,N_9890,N_9945);
nand UO_1185 (O_1185,N_9839,N_9843);
or UO_1186 (O_1186,N_9951,N_9884);
and UO_1187 (O_1187,N_9894,N_9972);
or UO_1188 (O_1188,N_9883,N_9857);
nand UO_1189 (O_1189,N_9930,N_9914);
nor UO_1190 (O_1190,N_9992,N_9864);
nand UO_1191 (O_1191,N_9926,N_9842);
or UO_1192 (O_1192,N_9958,N_9980);
nand UO_1193 (O_1193,N_9899,N_9857);
or UO_1194 (O_1194,N_9885,N_9977);
or UO_1195 (O_1195,N_9914,N_9870);
or UO_1196 (O_1196,N_9879,N_9868);
and UO_1197 (O_1197,N_9894,N_9958);
or UO_1198 (O_1198,N_9945,N_9885);
nand UO_1199 (O_1199,N_9912,N_9815);
and UO_1200 (O_1200,N_9913,N_9904);
nand UO_1201 (O_1201,N_9810,N_9951);
nand UO_1202 (O_1202,N_9845,N_9832);
nor UO_1203 (O_1203,N_9912,N_9926);
nor UO_1204 (O_1204,N_9942,N_9835);
nand UO_1205 (O_1205,N_9960,N_9888);
and UO_1206 (O_1206,N_9908,N_9984);
or UO_1207 (O_1207,N_9988,N_9928);
nand UO_1208 (O_1208,N_9920,N_9872);
and UO_1209 (O_1209,N_9899,N_9959);
nor UO_1210 (O_1210,N_9958,N_9897);
and UO_1211 (O_1211,N_9983,N_9939);
and UO_1212 (O_1212,N_9929,N_9984);
nand UO_1213 (O_1213,N_9851,N_9801);
nand UO_1214 (O_1214,N_9858,N_9918);
nor UO_1215 (O_1215,N_9904,N_9976);
nand UO_1216 (O_1216,N_9875,N_9811);
nand UO_1217 (O_1217,N_9899,N_9812);
or UO_1218 (O_1218,N_9851,N_9986);
and UO_1219 (O_1219,N_9884,N_9905);
and UO_1220 (O_1220,N_9806,N_9855);
and UO_1221 (O_1221,N_9909,N_9896);
or UO_1222 (O_1222,N_9840,N_9810);
and UO_1223 (O_1223,N_9827,N_9838);
nand UO_1224 (O_1224,N_9977,N_9834);
nor UO_1225 (O_1225,N_9988,N_9856);
nor UO_1226 (O_1226,N_9913,N_9987);
and UO_1227 (O_1227,N_9907,N_9916);
or UO_1228 (O_1228,N_9911,N_9862);
or UO_1229 (O_1229,N_9863,N_9875);
or UO_1230 (O_1230,N_9961,N_9967);
or UO_1231 (O_1231,N_9946,N_9993);
nand UO_1232 (O_1232,N_9914,N_9904);
nand UO_1233 (O_1233,N_9934,N_9894);
and UO_1234 (O_1234,N_9985,N_9973);
or UO_1235 (O_1235,N_9899,N_9852);
and UO_1236 (O_1236,N_9909,N_9876);
or UO_1237 (O_1237,N_9958,N_9993);
or UO_1238 (O_1238,N_9909,N_9947);
and UO_1239 (O_1239,N_9846,N_9894);
nor UO_1240 (O_1240,N_9903,N_9976);
nand UO_1241 (O_1241,N_9951,N_9929);
and UO_1242 (O_1242,N_9937,N_9854);
nor UO_1243 (O_1243,N_9930,N_9803);
or UO_1244 (O_1244,N_9816,N_9853);
or UO_1245 (O_1245,N_9829,N_9965);
and UO_1246 (O_1246,N_9935,N_9941);
or UO_1247 (O_1247,N_9811,N_9964);
nand UO_1248 (O_1248,N_9908,N_9928);
nor UO_1249 (O_1249,N_9841,N_9919);
nand UO_1250 (O_1250,N_9982,N_9933);
or UO_1251 (O_1251,N_9953,N_9913);
nand UO_1252 (O_1252,N_9825,N_9891);
nor UO_1253 (O_1253,N_9882,N_9955);
or UO_1254 (O_1254,N_9994,N_9943);
or UO_1255 (O_1255,N_9802,N_9948);
or UO_1256 (O_1256,N_9864,N_9987);
or UO_1257 (O_1257,N_9912,N_9999);
or UO_1258 (O_1258,N_9850,N_9970);
nand UO_1259 (O_1259,N_9892,N_9997);
nor UO_1260 (O_1260,N_9857,N_9947);
nand UO_1261 (O_1261,N_9941,N_9969);
nand UO_1262 (O_1262,N_9884,N_9906);
nor UO_1263 (O_1263,N_9903,N_9868);
nand UO_1264 (O_1264,N_9976,N_9935);
nand UO_1265 (O_1265,N_9868,N_9807);
and UO_1266 (O_1266,N_9817,N_9847);
nor UO_1267 (O_1267,N_9819,N_9983);
or UO_1268 (O_1268,N_9995,N_9971);
nand UO_1269 (O_1269,N_9873,N_9822);
nor UO_1270 (O_1270,N_9923,N_9908);
or UO_1271 (O_1271,N_9893,N_9899);
nor UO_1272 (O_1272,N_9808,N_9844);
nor UO_1273 (O_1273,N_9828,N_9963);
and UO_1274 (O_1274,N_9939,N_9927);
nor UO_1275 (O_1275,N_9988,N_9984);
and UO_1276 (O_1276,N_9987,N_9874);
or UO_1277 (O_1277,N_9814,N_9995);
and UO_1278 (O_1278,N_9915,N_9938);
nand UO_1279 (O_1279,N_9942,N_9866);
nand UO_1280 (O_1280,N_9931,N_9962);
nand UO_1281 (O_1281,N_9838,N_9915);
nand UO_1282 (O_1282,N_9959,N_9862);
or UO_1283 (O_1283,N_9974,N_9963);
nor UO_1284 (O_1284,N_9845,N_9917);
or UO_1285 (O_1285,N_9928,N_9814);
or UO_1286 (O_1286,N_9863,N_9970);
and UO_1287 (O_1287,N_9951,N_9906);
or UO_1288 (O_1288,N_9975,N_9853);
nor UO_1289 (O_1289,N_9884,N_9930);
xor UO_1290 (O_1290,N_9932,N_9808);
and UO_1291 (O_1291,N_9821,N_9985);
and UO_1292 (O_1292,N_9972,N_9904);
and UO_1293 (O_1293,N_9815,N_9983);
or UO_1294 (O_1294,N_9858,N_9834);
nor UO_1295 (O_1295,N_9860,N_9940);
or UO_1296 (O_1296,N_9887,N_9857);
and UO_1297 (O_1297,N_9968,N_9811);
and UO_1298 (O_1298,N_9824,N_9907);
nand UO_1299 (O_1299,N_9806,N_9823);
nor UO_1300 (O_1300,N_9801,N_9920);
or UO_1301 (O_1301,N_9878,N_9936);
nand UO_1302 (O_1302,N_9837,N_9981);
or UO_1303 (O_1303,N_9952,N_9967);
or UO_1304 (O_1304,N_9965,N_9976);
nor UO_1305 (O_1305,N_9878,N_9993);
nand UO_1306 (O_1306,N_9921,N_9986);
nor UO_1307 (O_1307,N_9800,N_9919);
nand UO_1308 (O_1308,N_9881,N_9816);
and UO_1309 (O_1309,N_9870,N_9820);
and UO_1310 (O_1310,N_9816,N_9960);
or UO_1311 (O_1311,N_9844,N_9967);
nand UO_1312 (O_1312,N_9911,N_9962);
and UO_1313 (O_1313,N_9912,N_9861);
nor UO_1314 (O_1314,N_9939,N_9894);
or UO_1315 (O_1315,N_9848,N_9996);
or UO_1316 (O_1316,N_9949,N_9907);
nand UO_1317 (O_1317,N_9905,N_9947);
nand UO_1318 (O_1318,N_9929,N_9973);
nand UO_1319 (O_1319,N_9990,N_9932);
and UO_1320 (O_1320,N_9851,N_9942);
nor UO_1321 (O_1321,N_9915,N_9894);
nor UO_1322 (O_1322,N_9988,N_9819);
or UO_1323 (O_1323,N_9913,N_9963);
xnor UO_1324 (O_1324,N_9960,N_9930);
nor UO_1325 (O_1325,N_9811,N_9885);
nand UO_1326 (O_1326,N_9853,N_9802);
nand UO_1327 (O_1327,N_9946,N_9980);
nand UO_1328 (O_1328,N_9926,N_9891);
or UO_1329 (O_1329,N_9870,N_9978);
or UO_1330 (O_1330,N_9906,N_9810);
and UO_1331 (O_1331,N_9995,N_9913);
nor UO_1332 (O_1332,N_9874,N_9810);
nand UO_1333 (O_1333,N_9889,N_9816);
and UO_1334 (O_1334,N_9808,N_9964);
and UO_1335 (O_1335,N_9910,N_9875);
nor UO_1336 (O_1336,N_9901,N_9879);
xor UO_1337 (O_1337,N_9880,N_9842);
nand UO_1338 (O_1338,N_9816,N_9865);
and UO_1339 (O_1339,N_9854,N_9823);
nand UO_1340 (O_1340,N_9901,N_9883);
nor UO_1341 (O_1341,N_9971,N_9812);
or UO_1342 (O_1342,N_9924,N_9801);
and UO_1343 (O_1343,N_9847,N_9959);
nand UO_1344 (O_1344,N_9842,N_9811);
or UO_1345 (O_1345,N_9861,N_9850);
nand UO_1346 (O_1346,N_9989,N_9964);
or UO_1347 (O_1347,N_9845,N_9969);
or UO_1348 (O_1348,N_9989,N_9897);
nand UO_1349 (O_1349,N_9884,N_9981);
or UO_1350 (O_1350,N_9849,N_9982);
and UO_1351 (O_1351,N_9984,N_9858);
nor UO_1352 (O_1352,N_9972,N_9931);
and UO_1353 (O_1353,N_9964,N_9929);
and UO_1354 (O_1354,N_9845,N_9887);
or UO_1355 (O_1355,N_9864,N_9821);
or UO_1356 (O_1356,N_9877,N_9892);
nand UO_1357 (O_1357,N_9879,N_9833);
or UO_1358 (O_1358,N_9804,N_9890);
nor UO_1359 (O_1359,N_9999,N_9967);
and UO_1360 (O_1360,N_9948,N_9962);
and UO_1361 (O_1361,N_9855,N_9827);
nand UO_1362 (O_1362,N_9822,N_9950);
or UO_1363 (O_1363,N_9995,N_9818);
nand UO_1364 (O_1364,N_9811,N_9808);
and UO_1365 (O_1365,N_9826,N_9999);
or UO_1366 (O_1366,N_9870,N_9864);
nand UO_1367 (O_1367,N_9899,N_9801);
and UO_1368 (O_1368,N_9960,N_9822);
and UO_1369 (O_1369,N_9824,N_9952);
or UO_1370 (O_1370,N_9955,N_9930);
or UO_1371 (O_1371,N_9939,N_9871);
nor UO_1372 (O_1372,N_9893,N_9971);
nor UO_1373 (O_1373,N_9906,N_9925);
or UO_1374 (O_1374,N_9940,N_9863);
or UO_1375 (O_1375,N_9839,N_9831);
and UO_1376 (O_1376,N_9843,N_9817);
or UO_1377 (O_1377,N_9973,N_9801);
nor UO_1378 (O_1378,N_9813,N_9823);
nand UO_1379 (O_1379,N_9841,N_9920);
nand UO_1380 (O_1380,N_9845,N_9966);
or UO_1381 (O_1381,N_9917,N_9985);
and UO_1382 (O_1382,N_9885,N_9880);
nand UO_1383 (O_1383,N_9843,N_9873);
and UO_1384 (O_1384,N_9960,N_9859);
nor UO_1385 (O_1385,N_9888,N_9915);
nand UO_1386 (O_1386,N_9857,N_9957);
nand UO_1387 (O_1387,N_9891,N_9950);
and UO_1388 (O_1388,N_9814,N_9998);
nand UO_1389 (O_1389,N_9896,N_9901);
nor UO_1390 (O_1390,N_9887,N_9980);
nor UO_1391 (O_1391,N_9929,N_9875);
or UO_1392 (O_1392,N_9938,N_9953);
or UO_1393 (O_1393,N_9840,N_9826);
nand UO_1394 (O_1394,N_9940,N_9945);
or UO_1395 (O_1395,N_9844,N_9889);
or UO_1396 (O_1396,N_9904,N_9912);
or UO_1397 (O_1397,N_9912,N_9860);
and UO_1398 (O_1398,N_9920,N_9864);
and UO_1399 (O_1399,N_9812,N_9912);
and UO_1400 (O_1400,N_9857,N_9819);
or UO_1401 (O_1401,N_9935,N_9953);
nor UO_1402 (O_1402,N_9974,N_9941);
or UO_1403 (O_1403,N_9831,N_9964);
nor UO_1404 (O_1404,N_9875,N_9916);
and UO_1405 (O_1405,N_9977,N_9813);
and UO_1406 (O_1406,N_9805,N_9942);
nand UO_1407 (O_1407,N_9879,N_9829);
nor UO_1408 (O_1408,N_9963,N_9883);
or UO_1409 (O_1409,N_9814,N_9818);
or UO_1410 (O_1410,N_9860,N_9850);
nor UO_1411 (O_1411,N_9865,N_9806);
nor UO_1412 (O_1412,N_9902,N_9936);
nand UO_1413 (O_1413,N_9807,N_9902);
nor UO_1414 (O_1414,N_9847,N_9940);
or UO_1415 (O_1415,N_9866,N_9928);
nand UO_1416 (O_1416,N_9841,N_9873);
nor UO_1417 (O_1417,N_9828,N_9881);
or UO_1418 (O_1418,N_9821,N_9866);
and UO_1419 (O_1419,N_9859,N_9840);
nand UO_1420 (O_1420,N_9803,N_9938);
nand UO_1421 (O_1421,N_9815,N_9975);
nand UO_1422 (O_1422,N_9807,N_9996);
and UO_1423 (O_1423,N_9881,N_9991);
xor UO_1424 (O_1424,N_9980,N_9964);
and UO_1425 (O_1425,N_9975,N_9928);
and UO_1426 (O_1426,N_9835,N_9906);
nor UO_1427 (O_1427,N_9938,N_9997);
nor UO_1428 (O_1428,N_9942,N_9855);
or UO_1429 (O_1429,N_9934,N_9866);
nand UO_1430 (O_1430,N_9985,N_9819);
nor UO_1431 (O_1431,N_9903,N_9914);
nand UO_1432 (O_1432,N_9828,N_9863);
and UO_1433 (O_1433,N_9956,N_9825);
and UO_1434 (O_1434,N_9803,N_9903);
nand UO_1435 (O_1435,N_9948,N_9942);
nand UO_1436 (O_1436,N_9820,N_9981);
and UO_1437 (O_1437,N_9878,N_9811);
nor UO_1438 (O_1438,N_9837,N_9834);
nand UO_1439 (O_1439,N_9801,N_9871);
or UO_1440 (O_1440,N_9895,N_9913);
or UO_1441 (O_1441,N_9859,N_9925);
nand UO_1442 (O_1442,N_9858,N_9852);
and UO_1443 (O_1443,N_9896,N_9908);
nand UO_1444 (O_1444,N_9942,N_9989);
nor UO_1445 (O_1445,N_9925,N_9839);
nand UO_1446 (O_1446,N_9960,N_9917);
xnor UO_1447 (O_1447,N_9845,N_9898);
nor UO_1448 (O_1448,N_9893,N_9996);
xor UO_1449 (O_1449,N_9964,N_9903);
or UO_1450 (O_1450,N_9941,N_9841);
nand UO_1451 (O_1451,N_9811,N_9967);
or UO_1452 (O_1452,N_9934,N_9811);
nand UO_1453 (O_1453,N_9945,N_9893);
nor UO_1454 (O_1454,N_9830,N_9849);
nand UO_1455 (O_1455,N_9968,N_9848);
nand UO_1456 (O_1456,N_9948,N_9804);
nand UO_1457 (O_1457,N_9940,N_9993);
nand UO_1458 (O_1458,N_9928,N_9952);
and UO_1459 (O_1459,N_9870,N_9946);
or UO_1460 (O_1460,N_9803,N_9819);
nand UO_1461 (O_1461,N_9965,N_9848);
and UO_1462 (O_1462,N_9968,N_9882);
and UO_1463 (O_1463,N_9959,N_9873);
and UO_1464 (O_1464,N_9866,N_9955);
nor UO_1465 (O_1465,N_9820,N_9934);
nor UO_1466 (O_1466,N_9958,N_9873);
nand UO_1467 (O_1467,N_9888,N_9992);
or UO_1468 (O_1468,N_9823,N_9840);
nand UO_1469 (O_1469,N_9978,N_9887);
or UO_1470 (O_1470,N_9964,N_9806);
nand UO_1471 (O_1471,N_9859,N_9891);
nor UO_1472 (O_1472,N_9831,N_9905);
nand UO_1473 (O_1473,N_9967,N_9871);
nor UO_1474 (O_1474,N_9811,N_9962);
nand UO_1475 (O_1475,N_9899,N_9828);
nor UO_1476 (O_1476,N_9942,N_9955);
and UO_1477 (O_1477,N_9841,N_9804);
nand UO_1478 (O_1478,N_9812,N_9890);
nor UO_1479 (O_1479,N_9981,N_9986);
or UO_1480 (O_1480,N_9834,N_9988);
and UO_1481 (O_1481,N_9813,N_9991);
and UO_1482 (O_1482,N_9940,N_9879);
nor UO_1483 (O_1483,N_9939,N_9834);
or UO_1484 (O_1484,N_9833,N_9843);
nor UO_1485 (O_1485,N_9833,N_9991);
and UO_1486 (O_1486,N_9982,N_9912);
nor UO_1487 (O_1487,N_9903,N_9834);
and UO_1488 (O_1488,N_9817,N_9900);
or UO_1489 (O_1489,N_9961,N_9872);
and UO_1490 (O_1490,N_9879,N_9889);
nor UO_1491 (O_1491,N_9903,N_9833);
nand UO_1492 (O_1492,N_9864,N_9932);
nand UO_1493 (O_1493,N_9833,N_9961);
nand UO_1494 (O_1494,N_9864,N_9905);
nor UO_1495 (O_1495,N_9816,N_9820);
nand UO_1496 (O_1496,N_9901,N_9990);
and UO_1497 (O_1497,N_9827,N_9950);
nand UO_1498 (O_1498,N_9972,N_9983);
nor UO_1499 (O_1499,N_9828,N_9875);
endmodule