module basic_500_3000_500_60_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_122,In_288);
and U1 (N_1,In_385,In_236);
nor U2 (N_2,In_428,In_191);
or U3 (N_3,In_137,In_93);
nor U4 (N_4,In_318,In_242);
nand U5 (N_5,In_68,In_226);
and U6 (N_6,In_335,In_434);
nor U7 (N_7,In_124,In_5);
nand U8 (N_8,In_159,In_322);
or U9 (N_9,In_212,In_278);
or U10 (N_10,In_310,In_371);
and U11 (N_11,In_350,In_139);
and U12 (N_12,In_197,In_297);
xnor U13 (N_13,In_131,In_491);
nor U14 (N_14,In_337,In_425);
xor U15 (N_15,In_125,In_101);
and U16 (N_16,In_243,In_377);
or U17 (N_17,In_311,In_307);
nor U18 (N_18,In_53,In_18);
nand U19 (N_19,In_327,In_163);
xnor U20 (N_20,In_422,In_312);
nand U21 (N_21,In_479,In_282);
and U22 (N_22,In_25,In_386);
xnor U23 (N_23,In_403,In_215);
or U24 (N_24,In_321,In_23);
nor U25 (N_25,In_272,In_380);
and U26 (N_26,In_416,In_473);
or U27 (N_27,In_61,In_150);
or U28 (N_28,In_280,In_482);
and U29 (N_29,In_201,In_481);
and U30 (N_30,In_22,In_289);
and U31 (N_31,In_302,In_7);
or U32 (N_32,In_248,In_264);
xor U33 (N_33,In_354,In_96);
nand U34 (N_34,In_493,In_56);
nor U35 (N_35,In_194,In_104);
nor U36 (N_36,In_362,In_470);
or U37 (N_37,In_314,In_329);
nand U38 (N_38,In_393,In_384);
or U39 (N_39,In_462,In_443);
or U40 (N_40,In_465,In_82);
or U41 (N_41,In_148,In_246);
and U42 (N_42,In_143,In_235);
nor U43 (N_43,In_169,In_352);
and U44 (N_44,In_144,In_461);
and U45 (N_45,In_63,In_27);
or U46 (N_46,In_132,In_234);
or U47 (N_47,In_138,In_0);
or U48 (N_48,In_256,In_347);
or U49 (N_49,In_88,In_48);
xor U50 (N_50,In_460,In_58);
nand U51 (N_51,In_180,In_437);
and U52 (N_52,N_5,In_486);
or U53 (N_53,N_48,In_432);
nand U54 (N_54,In_214,In_45);
xor U55 (N_55,In_423,In_414);
and U56 (N_56,In_251,In_364);
xnor U57 (N_57,In_490,In_412);
nand U58 (N_58,In_92,In_97);
nand U59 (N_59,In_449,In_303);
and U60 (N_60,In_213,In_219);
nor U61 (N_61,In_119,In_285);
xor U62 (N_62,In_86,In_231);
and U63 (N_63,In_128,In_287);
and U64 (N_64,In_19,In_12);
and U65 (N_65,In_474,N_18);
nand U66 (N_66,In_330,In_55);
nand U67 (N_67,In_346,In_174);
xnor U68 (N_68,In_396,In_165);
nand U69 (N_69,In_66,In_305);
or U70 (N_70,In_472,In_34);
and U71 (N_71,In_149,In_426);
and U72 (N_72,In_75,In_74);
nor U73 (N_73,In_336,In_279);
xnor U74 (N_74,In_40,In_366);
nand U75 (N_75,In_306,In_464);
xnor U76 (N_76,In_77,N_38);
or U77 (N_77,In_485,In_382);
and U78 (N_78,In_253,In_233);
and U79 (N_79,In_395,In_185);
and U80 (N_80,In_487,In_227);
or U81 (N_81,In_152,N_22);
xor U82 (N_82,In_195,In_378);
nand U83 (N_83,N_46,N_10);
nor U84 (N_84,In_49,In_146);
or U85 (N_85,In_161,In_237);
xnor U86 (N_86,In_390,In_444);
nor U87 (N_87,In_351,In_6);
nand U88 (N_88,In_50,In_295);
and U89 (N_89,In_145,In_118);
and U90 (N_90,In_320,In_155);
or U91 (N_91,In_26,In_244);
and U92 (N_92,In_455,In_361);
xor U93 (N_93,In_339,In_269);
nor U94 (N_94,In_98,N_6);
nand U95 (N_95,In_373,In_73);
nand U96 (N_96,N_9,In_223);
nand U97 (N_97,In_52,In_117);
xnor U98 (N_98,In_411,In_308);
xor U99 (N_99,In_170,In_162);
or U100 (N_100,In_331,In_166);
nand U101 (N_101,In_401,In_54);
or U102 (N_102,In_433,In_247);
nand U103 (N_103,In_156,In_9);
nor U104 (N_104,In_484,In_46);
xnor U105 (N_105,N_37,In_181);
nand U106 (N_106,In_47,In_116);
and U107 (N_107,In_172,In_179);
xnor U108 (N_108,In_356,N_81);
xnor U109 (N_109,In_100,In_192);
and U110 (N_110,In_415,In_20);
nor U111 (N_111,In_72,In_198);
and U112 (N_112,In_431,In_355);
or U113 (N_113,N_75,In_276);
nor U114 (N_114,In_277,In_480);
nand U115 (N_115,N_65,In_126);
and U116 (N_116,In_274,In_41);
nor U117 (N_117,In_99,In_467);
nor U118 (N_118,In_57,In_394);
and U119 (N_119,In_316,In_193);
nand U120 (N_120,N_30,N_15);
nor U121 (N_121,In_70,In_267);
and U122 (N_122,In_109,In_370);
or U123 (N_123,N_19,In_21);
nor U124 (N_124,In_463,In_298);
nand U125 (N_125,N_24,In_13);
xor U126 (N_126,In_405,N_74);
xor U127 (N_127,In_142,In_447);
xor U128 (N_128,In_85,In_207);
and U129 (N_129,In_15,In_317);
xor U130 (N_130,In_60,In_292);
nor U131 (N_131,In_59,N_89);
and U132 (N_132,In_451,In_257);
xnor U133 (N_133,In_392,In_333);
xor U134 (N_134,In_134,In_301);
xnor U135 (N_135,In_439,In_176);
nand U136 (N_136,In_35,In_11);
nand U137 (N_137,In_438,In_400);
xnor U138 (N_138,N_60,In_399);
and U139 (N_139,In_435,In_135);
or U140 (N_140,In_200,N_63);
and U141 (N_141,N_55,In_497);
nand U142 (N_142,N_84,In_189);
nor U143 (N_143,N_57,In_183);
nand U144 (N_144,In_39,N_20);
nor U145 (N_145,In_325,In_175);
or U146 (N_146,In_332,N_66);
xor U147 (N_147,In_37,In_471);
nand U148 (N_148,N_90,In_387);
xnor U149 (N_149,In_91,In_222);
nor U150 (N_150,In_216,In_457);
or U151 (N_151,In_51,In_488);
xor U152 (N_152,N_91,In_151);
or U153 (N_153,N_93,In_408);
xnor U154 (N_154,In_168,N_70);
or U155 (N_155,N_25,In_343);
and U156 (N_156,In_30,N_101);
nor U157 (N_157,In_407,In_140);
xor U158 (N_158,In_129,In_36);
xor U159 (N_159,In_105,In_315);
nand U160 (N_160,N_99,In_76);
or U161 (N_161,In_32,In_397);
xnor U162 (N_162,In_188,N_144);
xor U163 (N_163,In_294,N_3);
nor U164 (N_164,In_208,N_149);
xnor U165 (N_165,In_217,In_283);
nand U166 (N_166,N_32,In_342);
and U167 (N_167,N_79,N_117);
and U168 (N_168,In_255,N_56);
xnor U169 (N_169,N_114,N_123);
or U170 (N_170,In_209,N_41);
nor U171 (N_171,N_116,N_95);
or U172 (N_172,In_359,In_483);
nand U173 (N_173,N_129,N_136);
xor U174 (N_174,In_167,In_419);
nor U175 (N_175,In_357,In_81);
nor U176 (N_176,N_141,N_42);
xor U177 (N_177,In_340,In_344);
nand U178 (N_178,In_313,In_65);
and U179 (N_179,N_104,N_85);
xnor U180 (N_180,N_100,In_476);
and U181 (N_181,In_102,In_293);
and U182 (N_182,N_17,In_478);
nand U183 (N_183,In_44,In_121);
or U184 (N_184,In_218,N_105);
xnor U185 (N_185,In_38,In_221);
nor U186 (N_186,N_62,N_14);
nor U187 (N_187,In_263,N_50);
and U188 (N_188,In_89,N_61);
or U189 (N_189,N_7,In_489);
and U190 (N_190,In_14,In_64);
xnor U191 (N_191,In_17,N_121);
or U192 (N_192,N_59,In_78);
nand U193 (N_193,N_71,In_83);
or U194 (N_194,In_187,In_410);
and U195 (N_195,N_94,N_102);
and U196 (N_196,In_113,In_324);
or U197 (N_197,N_27,In_466);
or U198 (N_198,N_120,N_78);
nand U199 (N_199,N_87,In_365);
and U200 (N_200,N_113,In_28);
xor U201 (N_201,In_446,N_162);
or U202 (N_202,N_109,N_128);
xor U203 (N_203,In_328,In_290);
and U204 (N_204,In_186,In_250);
nand U205 (N_205,In_296,N_29);
nand U206 (N_206,In_133,In_304);
nor U207 (N_207,In_204,N_195);
xor U208 (N_208,In_158,In_459);
and U209 (N_209,N_157,N_169);
and U210 (N_210,In_429,In_436);
nor U211 (N_211,N_197,In_271);
nor U212 (N_212,In_427,In_178);
nand U213 (N_213,In_24,In_450);
xor U214 (N_214,In_475,N_161);
nand U215 (N_215,In_220,N_11);
or U216 (N_216,In_87,N_26);
and U217 (N_217,In_260,N_186);
nand U218 (N_218,N_158,N_47);
and U219 (N_219,In_300,In_8);
and U220 (N_220,In_448,In_468);
nand U221 (N_221,N_51,N_134);
xnor U222 (N_222,In_141,In_430);
nor U223 (N_223,In_29,In_309);
xor U224 (N_224,In_173,In_4);
nand U225 (N_225,In_367,In_273);
xor U226 (N_226,In_164,In_130);
and U227 (N_227,In_203,In_210);
nand U228 (N_228,In_275,N_165);
and U229 (N_229,N_33,N_80);
or U230 (N_230,N_198,In_418);
nand U231 (N_231,In_42,In_205);
nor U232 (N_232,In_440,In_245);
xnor U233 (N_233,In_496,In_106);
nor U234 (N_234,N_40,In_238);
xor U235 (N_235,N_166,N_130);
nor U236 (N_236,In_258,In_406);
and U237 (N_237,N_171,N_178);
nand U238 (N_238,In_240,In_177);
nor U239 (N_239,In_196,N_98);
nand U240 (N_240,N_194,In_360);
and U241 (N_241,In_10,In_123);
and U242 (N_242,N_43,N_112);
or U243 (N_243,N_73,In_239);
or U244 (N_244,In_228,In_454);
xnor U245 (N_245,N_172,In_110);
nand U246 (N_246,N_119,In_492);
xor U247 (N_247,In_363,In_265);
or U248 (N_248,N_170,N_111);
nand U249 (N_249,In_358,N_72);
xnor U250 (N_250,N_31,In_127);
xnor U251 (N_251,In_232,N_213);
and U252 (N_252,In_389,N_155);
nor U253 (N_253,N_229,N_4);
nor U254 (N_254,N_34,N_132);
nand U255 (N_255,N_182,In_477);
or U256 (N_256,N_211,N_204);
xnor U257 (N_257,In_3,N_196);
or U258 (N_258,In_388,In_80);
nand U259 (N_259,N_240,In_284);
or U260 (N_260,In_319,In_270);
or U261 (N_261,N_231,N_159);
nand U262 (N_262,N_210,N_68);
and U263 (N_263,In_376,In_421);
nor U264 (N_264,N_249,N_103);
nor U265 (N_265,In_441,N_246);
and U266 (N_266,In_334,N_106);
nand U267 (N_267,In_114,N_150);
nor U268 (N_268,N_64,N_188);
and U269 (N_269,N_245,N_82);
xnor U270 (N_270,N_44,In_160);
or U271 (N_271,In_398,N_176);
and U272 (N_272,N_164,N_115);
nand U273 (N_273,N_203,N_36);
or U274 (N_274,N_206,In_95);
xnor U275 (N_275,N_223,In_90);
and U276 (N_276,In_281,N_233);
nor U277 (N_277,In_94,N_200);
and U278 (N_278,N_28,In_103);
nand U279 (N_279,N_163,In_229);
or U280 (N_280,In_43,N_160);
and U281 (N_281,N_221,In_259);
xnor U282 (N_282,N_69,N_92);
nor U283 (N_283,N_225,In_495);
xnor U284 (N_284,In_452,In_409);
nor U285 (N_285,N_234,In_286);
xnor U286 (N_286,N_222,N_97);
and U287 (N_287,In_442,N_214);
nand U288 (N_288,In_153,In_326);
or U289 (N_289,N_184,N_227);
and U290 (N_290,In_420,N_148);
nand U291 (N_291,N_125,In_62);
and U292 (N_292,N_217,N_0);
nor U293 (N_293,N_215,In_79);
nand U294 (N_294,N_244,In_31);
nor U295 (N_295,N_135,N_191);
or U296 (N_296,N_168,In_16);
and U297 (N_297,In_345,N_218);
nor U298 (N_298,In_249,In_108);
nor U299 (N_299,In_369,N_124);
and U300 (N_300,In_115,N_255);
nand U301 (N_301,N_107,In_154);
and U302 (N_302,N_35,N_235);
nand U303 (N_303,In_348,N_16);
and U304 (N_304,N_201,N_193);
and U305 (N_305,N_295,N_285);
nand U306 (N_306,In_375,N_199);
and U307 (N_307,In_381,N_268);
and U308 (N_308,In_1,N_192);
or U309 (N_309,In_136,N_286);
nor U310 (N_310,N_77,N_239);
nand U311 (N_311,In_349,N_122);
xnor U312 (N_312,N_284,N_52);
nor U313 (N_313,N_243,In_147);
xnor U314 (N_314,N_271,In_469);
nand U315 (N_315,In_69,N_190);
nand U316 (N_316,N_280,N_238);
nor U317 (N_317,N_205,N_277);
nor U318 (N_318,In_67,N_180);
xor U319 (N_319,N_290,In_211);
xor U320 (N_320,In_338,N_147);
nand U321 (N_321,N_185,N_156);
and U322 (N_322,N_67,N_13);
nand U323 (N_323,N_279,N_139);
or U324 (N_324,In_230,N_138);
nand U325 (N_325,N_263,In_268);
or U326 (N_326,N_118,N_49);
nor U327 (N_327,N_23,N_230);
xor U328 (N_328,N_220,N_283);
nor U329 (N_329,N_252,In_372);
xnor U330 (N_330,In_206,N_174);
xor U331 (N_331,N_181,In_224);
or U332 (N_332,In_499,In_171);
xor U333 (N_333,N_2,N_269);
nor U334 (N_334,N_299,N_247);
and U335 (N_335,N_298,N_292);
and U336 (N_336,N_236,N_208);
nand U337 (N_337,N_262,N_207);
and U338 (N_338,N_275,In_299);
or U339 (N_339,N_189,N_266);
nor U340 (N_340,N_140,N_256);
nor U341 (N_341,N_39,In_71);
and U342 (N_342,N_21,In_353);
nor U343 (N_343,N_219,N_212);
and U344 (N_344,N_253,N_254);
and U345 (N_345,N_242,In_199);
and U346 (N_346,N_260,N_251);
or U347 (N_347,N_228,N_96);
nor U348 (N_348,N_241,N_8);
or U349 (N_349,N_282,N_143);
and U350 (N_350,N_310,N_342);
nor U351 (N_351,N_250,N_308);
xnor U352 (N_352,In_417,N_305);
and U353 (N_353,N_300,In_262);
nor U354 (N_354,N_264,In_341);
and U355 (N_355,N_343,N_297);
or U356 (N_356,N_237,N_183);
or U357 (N_357,N_302,In_368);
nor U358 (N_358,In_424,N_314);
nand U359 (N_359,In_458,N_281);
and U360 (N_360,N_331,N_311);
nor U361 (N_361,N_315,In_494);
nand U362 (N_362,N_175,N_303);
nand U363 (N_363,N_1,N_274);
xnor U364 (N_364,N_153,N_167);
and U365 (N_365,In_413,In_241);
nor U366 (N_366,In_84,In_402);
nor U367 (N_367,N_248,In_456);
nand U368 (N_368,In_202,In_383);
xnor U369 (N_369,N_45,N_151);
nand U370 (N_370,N_291,N_289);
xor U371 (N_371,N_326,N_270);
xor U372 (N_372,N_276,N_273);
xnor U373 (N_373,N_110,N_333);
and U374 (N_374,N_341,N_152);
nand U375 (N_375,N_332,N_321);
nand U376 (N_376,In_252,N_317);
or U377 (N_377,N_261,In_266);
and U378 (N_378,N_312,N_216);
xnor U379 (N_379,N_226,N_131);
or U380 (N_380,In_291,N_316);
and U381 (N_381,N_265,N_323);
nor U382 (N_382,N_278,In_182);
nand U383 (N_383,N_179,N_126);
xnor U384 (N_384,In_404,N_294);
nand U385 (N_385,In_323,N_267);
nor U386 (N_386,N_340,N_108);
or U387 (N_387,In_445,N_76);
nor U388 (N_388,N_287,N_337);
or U389 (N_389,In_453,N_133);
nor U390 (N_390,N_301,N_54);
and U391 (N_391,N_320,N_202);
nand U392 (N_392,N_347,N_209);
nor U393 (N_393,In_33,N_349);
and U394 (N_394,N_12,N_187);
xor U395 (N_395,N_127,N_344);
nor U396 (N_396,In_112,In_379);
and U397 (N_397,N_259,N_177);
or U398 (N_398,N_58,In_157);
nor U399 (N_399,N_142,N_83);
nand U400 (N_400,In_374,N_318);
nand U401 (N_401,N_356,In_107);
or U402 (N_402,N_173,N_367);
xnor U403 (N_403,N_379,N_390);
and U404 (N_404,N_145,In_111);
nor U405 (N_405,N_355,N_398);
or U406 (N_406,N_386,In_225);
and U407 (N_407,N_378,N_339);
nor U408 (N_408,N_154,N_368);
xnor U409 (N_409,N_370,N_304);
xor U410 (N_410,N_258,N_327);
xnor U411 (N_411,N_359,N_394);
and U412 (N_412,N_330,N_381);
nor U413 (N_413,N_319,N_335);
nor U414 (N_414,N_353,N_384);
nand U415 (N_415,N_346,N_324);
nor U416 (N_416,N_325,N_88);
or U417 (N_417,N_369,N_391);
and U418 (N_418,In_2,N_348);
xnor U419 (N_419,N_397,N_328);
and U420 (N_420,N_376,N_232);
and U421 (N_421,In_261,N_374);
nand U422 (N_422,N_338,N_86);
nor U423 (N_423,N_357,N_375);
nand U424 (N_424,N_288,N_352);
nor U425 (N_425,N_372,N_345);
nand U426 (N_426,N_362,N_224);
and U427 (N_427,N_387,N_385);
nand U428 (N_428,N_365,N_309);
and U429 (N_429,N_383,N_336);
or U430 (N_430,In_254,N_377);
nor U431 (N_431,N_399,N_334);
nor U432 (N_432,N_366,N_380);
nand U433 (N_433,N_146,N_360);
or U434 (N_434,N_393,N_351);
nand U435 (N_435,N_373,In_391);
nor U436 (N_436,N_361,N_363);
xnor U437 (N_437,In_184,N_257);
and U438 (N_438,N_296,N_389);
or U439 (N_439,N_322,In_190);
and U440 (N_440,N_382,In_120);
and U441 (N_441,N_364,N_388);
nor U442 (N_442,N_395,N_358);
or U443 (N_443,In_498,N_137);
or U444 (N_444,N_306,N_392);
nor U445 (N_445,N_293,N_396);
nor U446 (N_446,N_371,N_307);
or U447 (N_447,N_53,N_313);
or U448 (N_448,N_350,N_354);
and U449 (N_449,N_272,N_329);
and U450 (N_450,N_404,N_408);
nand U451 (N_451,N_445,N_428);
xnor U452 (N_452,N_414,N_407);
and U453 (N_453,N_448,N_412);
or U454 (N_454,N_437,N_434);
and U455 (N_455,N_422,N_432);
and U456 (N_456,N_401,N_443);
or U457 (N_457,N_425,N_430);
or U458 (N_458,N_415,N_423);
nand U459 (N_459,N_417,N_420);
and U460 (N_460,N_416,N_438);
nand U461 (N_461,N_433,N_435);
xor U462 (N_462,N_424,N_421);
nor U463 (N_463,N_413,N_400);
or U464 (N_464,N_429,N_405);
nor U465 (N_465,N_403,N_441);
nor U466 (N_466,N_446,N_419);
nand U467 (N_467,N_427,N_449);
xnor U468 (N_468,N_436,N_431);
nor U469 (N_469,N_411,N_418);
xnor U470 (N_470,N_402,N_439);
nand U471 (N_471,N_409,N_447);
xor U472 (N_472,N_426,N_406);
or U473 (N_473,N_410,N_440);
and U474 (N_474,N_444,N_442);
nand U475 (N_475,N_448,N_430);
nand U476 (N_476,N_439,N_438);
and U477 (N_477,N_402,N_407);
nand U478 (N_478,N_427,N_448);
and U479 (N_479,N_400,N_410);
xnor U480 (N_480,N_425,N_411);
nor U481 (N_481,N_404,N_416);
xor U482 (N_482,N_425,N_449);
nand U483 (N_483,N_430,N_415);
or U484 (N_484,N_439,N_431);
nor U485 (N_485,N_449,N_409);
xor U486 (N_486,N_444,N_447);
or U487 (N_487,N_424,N_437);
xor U488 (N_488,N_417,N_440);
nor U489 (N_489,N_426,N_444);
nand U490 (N_490,N_435,N_434);
xor U491 (N_491,N_417,N_423);
and U492 (N_492,N_410,N_406);
nand U493 (N_493,N_445,N_404);
nor U494 (N_494,N_407,N_410);
nand U495 (N_495,N_428,N_431);
nor U496 (N_496,N_423,N_405);
nand U497 (N_497,N_413,N_404);
nand U498 (N_498,N_436,N_434);
and U499 (N_499,N_432,N_415);
and U500 (N_500,N_453,N_457);
and U501 (N_501,N_468,N_465);
and U502 (N_502,N_452,N_497);
nor U503 (N_503,N_461,N_463);
xor U504 (N_504,N_450,N_474);
nor U505 (N_505,N_464,N_455);
and U506 (N_506,N_456,N_470);
nand U507 (N_507,N_477,N_476);
xor U508 (N_508,N_482,N_486);
or U509 (N_509,N_495,N_496);
xor U510 (N_510,N_485,N_481);
xnor U511 (N_511,N_488,N_472);
and U512 (N_512,N_479,N_462);
nand U513 (N_513,N_491,N_494);
nor U514 (N_514,N_490,N_467);
nand U515 (N_515,N_454,N_493);
nand U516 (N_516,N_487,N_460);
nor U517 (N_517,N_499,N_466);
or U518 (N_518,N_459,N_498);
and U519 (N_519,N_458,N_480);
or U520 (N_520,N_478,N_471);
nor U521 (N_521,N_483,N_473);
and U522 (N_522,N_451,N_475);
or U523 (N_523,N_492,N_469);
nand U524 (N_524,N_484,N_489);
nand U525 (N_525,N_489,N_461);
nor U526 (N_526,N_464,N_458);
or U527 (N_527,N_468,N_466);
xnor U528 (N_528,N_485,N_493);
nor U529 (N_529,N_482,N_483);
nand U530 (N_530,N_486,N_494);
nor U531 (N_531,N_467,N_480);
or U532 (N_532,N_493,N_457);
nor U533 (N_533,N_461,N_497);
nor U534 (N_534,N_493,N_489);
nand U535 (N_535,N_457,N_498);
and U536 (N_536,N_454,N_495);
nor U537 (N_537,N_466,N_484);
xor U538 (N_538,N_460,N_481);
nand U539 (N_539,N_453,N_495);
or U540 (N_540,N_479,N_478);
nor U541 (N_541,N_450,N_455);
nor U542 (N_542,N_490,N_479);
or U543 (N_543,N_469,N_494);
or U544 (N_544,N_499,N_483);
or U545 (N_545,N_459,N_491);
xor U546 (N_546,N_487,N_470);
nand U547 (N_547,N_457,N_475);
nand U548 (N_548,N_470,N_473);
and U549 (N_549,N_463,N_454);
nor U550 (N_550,N_543,N_520);
nor U551 (N_551,N_525,N_545);
nor U552 (N_552,N_506,N_541);
and U553 (N_553,N_527,N_528);
nor U554 (N_554,N_549,N_501);
and U555 (N_555,N_512,N_505);
xnor U556 (N_556,N_503,N_536);
and U557 (N_557,N_529,N_518);
nand U558 (N_558,N_532,N_531);
xnor U559 (N_559,N_538,N_509);
xor U560 (N_560,N_504,N_515);
and U561 (N_561,N_502,N_510);
xor U562 (N_562,N_513,N_522);
or U563 (N_563,N_524,N_547);
or U564 (N_564,N_540,N_526);
xnor U565 (N_565,N_516,N_530);
and U566 (N_566,N_534,N_517);
nand U567 (N_567,N_544,N_546);
and U568 (N_568,N_523,N_539);
and U569 (N_569,N_535,N_514);
or U570 (N_570,N_507,N_519);
nor U571 (N_571,N_511,N_521);
and U572 (N_572,N_542,N_500);
or U573 (N_573,N_533,N_508);
or U574 (N_574,N_537,N_548);
nand U575 (N_575,N_521,N_502);
nor U576 (N_576,N_540,N_533);
nor U577 (N_577,N_510,N_532);
xnor U578 (N_578,N_529,N_532);
and U579 (N_579,N_536,N_506);
xnor U580 (N_580,N_525,N_538);
or U581 (N_581,N_501,N_544);
or U582 (N_582,N_514,N_545);
xnor U583 (N_583,N_510,N_519);
and U584 (N_584,N_529,N_546);
xor U585 (N_585,N_546,N_514);
or U586 (N_586,N_530,N_535);
nor U587 (N_587,N_506,N_546);
xor U588 (N_588,N_534,N_545);
or U589 (N_589,N_512,N_532);
or U590 (N_590,N_542,N_503);
nor U591 (N_591,N_527,N_514);
or U592 (N_592,N_518,N_528);
nand U593 (N_593,N_538,N_532);
or U594 (N_594,N_541,N_539);
nand U595 (N_595,N_502,N_515);
or U596 (N_596,N_506,N_517);
xor U597 (N_597,N_515,N_505);
nand U598 (N_598,N_539,N_527);
and U599 (N_599,N_513,N_504);
xor U600 (N_600,N_581,N_565);
or U601 (N_601,N_570,N_590);
xnor U602 (N_602,N_580,N_583);
nor U603 (N_603,N_571,N_592);
nor U604 (N_604,N_550,N_586);
nor U605 (N_605,N_562,N_556);
and U606 (N_606,N_558,N_579);
and U607 (N_607,N_551,N_597);
and U608 (N_608,N_598,N_594);
nor U609 (N_609,N_566,N_588);
nor U610 (N_610,N_599,N_582);
nand U611 (N_611,N_572,N_554);
xnor U612 (N_612,N_564,N_561);
or U613 (N_613,N_559,N_596);
and U614 (N_614,N_568,N_593);
and U615 (N_615,N_552,N_560);
and U616 (N_616,N_589,N_591);
nand U617 (N_617,N_574,N_573);
and U618 (N_618,N_585,N_578);
nor U619 (N_619,N_584,N_553);
nor U620 (N_620,N_587,N_563);
or U621 (N_621,N_595,N_569);
xor U622 (N_622,N_557,N_567);
or U623 (N_623,N_555,N_575);
nor U624 (N_624,N_576,N_577);
and U625 (N_625,N_570,N_583);
nand U626 (N_626,N_559,N_586);
and U627 (N_627,N_566,N_581);
nor U628 (N_628,N_554,N_570);
or U629 (N_629,N_588,N_568);
or U630 (N_630,N_587,N_584);
nand U631 (N_631,N_573,N_569);
xnor U632 (N_632,N_592,N_564);
or U633 (N_633,N_590,N_583);
nand U634 (N_634,N_581,N_560);
or U635 (N_635,N_598,N_585);
nor U636 (N_636,N_575,N_581);
or U637 (N_637,N_592,N_583);
xnor U638 (N_638,N_574,N_557);
nor U639 (N_639,N_568,N_597);
nand U640 (N_640,N_586,N_551);
or U641 (N_641,N_599,N_554);
nand U642 (N_642,N_578,N_552);
and U643 (N_643,N_597,N_554);
xnor U644 (N_644,N_561,N_581);
nand U645 (N_645,N_559,N_598);
nor U646 (N_646,N_554,N_552);
nor U647 (N_647,N_588,N_575);
nand U648 (N_648,N_553,N_569);
or U649 (N_649,N_564,N_551);
nor U650 (N_650,N_630,N_610);
nand U651 (N_651,N_603,N_606);
nor U652 (N_652,N_628,N_644);
nor U653 (N_653,N_636,N_624);
and U654 (N_654,N_605,N_635);
or U655 (N_655,N_612,N_604);
and U656 (N_656,N_623,N_629);
xor U657 (N_657,N_615,N_613);
xor U658 (N_658,N_614,N_648);
and U659 (N_659,N_625,N_622);
and U660 (N_660,N_640,N_616);
or U661 (N_661,N_618,N_619);
or U662 (N_662,N_642,N_641);
nor U663 (N_663,N_643,N_607);
xnor U664 (N_664,N_617,N_600);
and U665 (N_665,N_638,N_647);
and U666 (N_666,N_649,N_626);
or U667 (N_667,N_632,N_645);
or U668 (N_668,N_611,N_601);
and U669 (N_669,N_633,N_646);
and U670 (N_670,N_637,N_608);
xor U671 (N_671,N_621,N_639);
or U672 (N_672,N_627,N_620);
nor U673 (N_673,N_631,N_634);
nor U674 (N_674,N_609,N_602);
or U675 (N_675,N_646,N_609);
or U676 (N_676,N_600,N_604);
xnor U677 (N_677,N_602,N_610);
nand U678 (N_678,N_615,N_622);
nor U679 (N_679,N_621,N_604);
and U680 (N_680,N_602,N_627);
xor U681 (N_681,N_602,N_626);
nor U682 (N_682,N_636,N_648);
xor U683 (N_683,N_630,N_617);
or U684 (N_684,N_604,N_623);
xnor U685 (N_685,N_602,N_613);
and U686 (N_686,N_641,N_644);
and U687 (N_687,N_620,N_625);
nand U688 (N_688,N_626,N_622);
xor U689 (N_689,N_604,N_628);
or U690 (N_690,N_636,N_632);
nand U691 (N_691,N_646,N_620);
nand U692 (N_692,N_634,N_644);
xor U693 (N_693,N_643,N_603);
nand U694 (N_694,N_612,N_623);
nor U695 (N_695,N_632,N_644);
and U696 (N_696,N_610,N_636);
or U697 (N_697,N_643,N_629);
nand U698 (N_698,N_641,N_634);
and U699 (N_699,N_646,N_639);
or U700 (N_700,N_659,N_673);
nor U701 (N_701,N_665,N_699);
nor U702 (N_702,N_670,N_688);
and U703 (N_703,N_655,N_679);
xor U704 (N_704,N_663,N_667);
nor U705 (N_705,N_692,N_677);
nand U706 (N_706,N_687,N_674);
or U707 (N_707,N_661,N_664);
nor U708 (N_708,N_668,N_666);
xnor U709 (N_709,N_678,N_682);
or U710 (N_710,N_696,N_651);
nand U711 (N_711,N_685,N_691);
nor U712 (N_712,N_693,N_654);
nand U713 (N_713,N_681,N_683);
nor U714 (N_714,N_669,N_680);
xnor U715 (N_715,N_697,N_675);
nand U716 (N_716,N_672,N_653);
or U717 (N_717,N_694,N_695);
and U718 (N_718,N_660,N_690);
nand U719 (N_719,N_662,N_686);
nand U720 (N_720,N_656,N_698);
nor U721 (N_721,N_684,N_658);
or U722 (N_722,N_671,N_689);
and U723 (N_723,N_676,N_650);
nand U724 (N_724,N_652,N_657);
xor U725 (N_725,N_693,N_659);
nor U726 (N_726,N_675,N_678);
nor U727 (N_727,N_689,N_696);
nand U728 (N_728,N_655,N_678);
nor U729 (N_729,N_688,N_691);
nor U730 (N_730,N_657,N_669);
or U731 (N_731,N_654,N_664);
nor U732 (N_732,N_690,N_657);
or U733 (N_733,N_695,N_677);
xor U734 (N_734,N_657,N_673);
and U735 (N_735,N_698,N_695);
xor U736 (N_736,N_696,N_655);
nand U737 (N_737,N_692,N_655);
xnor U738 (N_738,N_675,N_662);
nand U739 (N_739,N_696,N_662);
and U740 (N_740,N_697,N_658);
and U741 (N_741,N_666,N_697);
nor U742 (N_742,N_667,N_680);
nor U743 (N_743,N_699,N_664);
or U744 (N_744,N_676,N_653);
and U745 (N_745,N_655,N_680);
nand U746 (N_746,N_670,N_677);
and U747 (N_747,N_684,N_665);
and U748 (N_748,N_690,N_675);
nor U749 (N_749,N_693,N_670);
nor U750 (N_750,N_713,N_719);
nor U751 (N_751,N_747,N_743);
and U752 (N_752,N_727,N_720);
xor U753 (N_753,N_728,N_741);
nor U754 (N_754,N_738,N_730);
xnor U755 (N_755,N_722,N_717);
xor U756 (N_756,N_707,N_724);
xor U757 (N_757,N_711,N_704);
or U758 (N_758,N_737,N_731);
nand U759 (N_759,N_745,N_716);
or U760 (N_760,N_749,N_729);
and U761 (N_761,N_746,N_709);
nand U762 (N_762,N_714,N_739);
xnor U763 (N_763,N_703,N_712);
or U764 (N_764,N_726,N_706);
nor U765 (N_765,N_721,N_733);
or U766 (N_766,N_705,N_708);
and U767 (N_767,N_736,N_735);
or U768 (N_768,N_701,N_718);
nor U769 (N_769,N_732,N_742);
and U770 (N_770,N_700,N_748);
xor U771 (N_771,N_702,N_725);
xnor U772 (N_772,N_740,N_723);
nand U773 (N_773,N_710,N_734);
or U774 (N_774,N_715,N_744);
xor U775 (N_775,N_702,N_734);
and U776 (N_776,N_744,N_704);
nand U777 (N_777,N_725,N_734);
nand U778 (N_778,N_717,N_725);
nor U779 (N_779,N_739,N_700);
nand U780 (N_780,N_707,N_723);
and U781 (N_781,N_714,N_733);
xnor U782 (N_782,N_700,N_720);
xor U783 (N_783,N_729,N_705);
or U784 (N_784,N_747,N_734);
nand U785 (N_785,N_705,N_736);
xnor U786 (N_786,N_703,N_740);
xor U787 (N_787,N_749,N_732);
nor U788 (N_788,N_728,N_722);
nor U789 (N_789,N_735,N_709);
nand U790 (N_790,N_724,N_701);
or U791 (N_791,N_719,N_720);
and U792 (N_792,N_720,N_733);
or U793 (N_793,N_710,N_715);
and U794 (N_794,N_730,N_722);
nand U795 (N_795,N_702,N_700);
nor U796 (N_796,N_730,N_709);
nor U797 (N_797,N_724,N_711);
and U798 (N_798,N_717,N_719);
and U799 (N_799,N_735,N_745);
or U800 (N_800,N_757,N_760);
or U801 (N_801,N_783,N_764);
nor U802 (N_802,N_796,N_768);
xnor U803 (N_803,N_755,N_779);
or U804 (N_804,N_766,N_777);
xnor U805 (N_805,N_776,N_756);
nand U806 (N_806,N_792,N_769);
nor U807 (N_807,N_758,N_774);
and U808 (N_808,N_763,N_788);
and U809 (N_809,N_773,N_750);
and U810 (N_810,N_790,N_759);
or U811 (N_811,N_771,N_781);
or U812 (N_812,N_765,N_794);
and U813 (N_813,N_798,N_770);
or U814 (N_814,N_754,N_753);
and U815 (N_815,N_752,N_795);
and U816 (N_816,N_784,N_762);
or U817 (N_817,N_775,N_786);
xor U818 (N_818,N_793,N_761);
nor U819 (N_819,N_797,N_799);
xnor U820 (N_820,N_789,N_778);
nand U821 (N_821,N_767,N_787);
xnor U822 (N_822,N_791,N_772);
xnor U823 (N_823,N_785,N_751);
xnor U824 (N_824,N_780,N_782);
or U825 (N_825,N_782,N_752);
or U826 (N_826,N_758,N_762);
nor U827 (N_827,N_787,N_792);
nor U828 (N_828,N_783,N_756);
and U829 (N_829,N_796,N_795);
nand U830 (N_830,N_752,N_763);
xnor U831 (N_831,N_781,N_757);
nand U832 (N_832,N_794,N_760);
or U833 (N_833,N_792,N_755);
xor U834 (N_834,N_798,N_778);
nand U835 (N_835,N_791,N_768);
and U836 (N_836,N_777,N_783);
xnor U837 (N_837,N_766,N_779);
nor U838 (N_838,N_785,N_784);
and U839 (N_839,N_772,N_752);
and U840 (N_840,N_787,N_764);
nand U841 (N_841,N_757,N_759);
nor U842 (N_842,N_784,N_754);
or U843 (N_843,N_795,N_788);
xnor U844 (N_844,N_782,N_751);
nor U845 (N_845,N_756,N_752);
or U846 (N_846,N_785,N_765);
xor U847 (N_847,N_759,N_755);
or U848 (N_848,N_764,N_755);
or U849 (N_849,N_757,N_779);
or U850 (N_850,N_830,N_811);
xor U851 (N_851,N_845,N_833);
or U852 (N_852,N_832,N_822);
nor U853 (N_853,N_817,N_841);
nor U854 (N_854,N_805,N_818);
nor U855 (N_855,N_842,N_825);
and U856 (N_856,N_844,N_824);
nand U857 (N_857,N_821,N_848);
xor U858 (N_858,N_810,N_829);
or U859 (N_859,N_802,N_801);
and U860 (N_860,N_831,N_808);
and U861 (N_861,N_807,N_827);
and U862 (N_862,N_839,N_834);
and U863 (N_863,N_849,N_838);
xnor U864 (N_864,N_814,N_815);
xor U865 (N_865,N_800,N_846);
xnor U866 (N_866,N_847,N_809);
nor U867 (N_867,N_820,N_819);
nand U868 (N_868,N_840,N_804);
xnor U869 (N_869,N_826,N_836);
nor U870 (N_870,N_843,N_828);
and U871 (N_871,N_816,N_837);
nand U872 (N_872,N_813,N_806);
nor U873 (N_873,N_835,N_803);
xor U874 (N_874,N_823,N_812);
or U875 (N_875,N_829,N_828);
xnor U876 (N_876,N_803,N_817);
and U877 (N_877,N_845,N_814);
xnor U878 (N_878,N_831,N_814);
or U879 (N_879,N_846,N_811);
and U880 (N_880,N_844,N_845);
or U881 (N_881,N_848,N_814);
nor U882 (N_882,N_847,N_828);
xnor U883 (N_883,N_835,N_802);
nand U884 (N_884,N_802,N_814);
xor U885 (N_885,N_806,N_807);
nand U886 (N_886,N_815,N_837);
or U887 (N_887,N_832,N_849);
nor U888 (N_888,N_819,N_808);
nor U889 (N_889,N_817,N_839);
xor U890 (N_890,N_847,N_831);
nand U891 (N_891,N_822,N_817);
nor U892 (N_892,N_821,N_849);
and U893 (N_893,N_801,N_845);
xor U894 (N_894,N_813,N_802);
nand U895 (N_895,N_846,N_807);
and U896 (N_896,N_817,N_835);
xnor U897 (N_897,N_843,N_849);
or U898 (N_898,N_843,N_836);
and U899 (N_899,N_840,N_848);
or U900 (N_900,N_886,N_851);
xor U901 (N_901,N_880,N_858);
nand U902 (N_902,N_875,N_888);
nand U903 (N_903,N_856,N_871);
xnor U904 (N_904,N_899,N_877);
and U905 (N_905,N_868,N_898);
xnor U906 (N_906,N_864,N_876);
and U907 (N_907,N_892,N_857);
nand U908 (N_908,N_885,N_863);
or U909 (N_909,N_861,N_866);
xnor U910 (N_910,N_894,N_870);
nor U911 (N_911,N_874,N_862);
xnor U912 (N_912,N_860,N_882);
nor U913 (N_913,N_869,N_893);
or U914 (N_914,N_891,N_879);
nor U915 (N_915,N_896,N_883);
and U916 (N_916,N_897,N_853);
nand U917 (N_917,N_854,N_881);
nand U918 (N_918,N_878,N_852);
nor U919 (N_919,N_895,N_887);
nand U920 (N_920,N_872,N_889);
or U921 (N_921,N_855,N_850);
or U922 (N_922,N_859,N_890);
nor U923 (N_923,N_873,N_867);
or U924 (N_924,N_884,N_865);
and U925 (N_925,N_862,N_881);
xor U926 (N_926,N_894,N_869);
nand U927 (N_927,N_882,N_878);
nor U928 (N_928,N_888,N_872);
xnor U929 (N_929,N_875,N_867);
xor U930 (N_930,N_852,N_873);
nor U931 (N_931,N_853,N_892);
nor U932 (N_932,N_884,N_895);
xnor U933 (N_933,N_890,N_868);
or U934 (N_934,N_851,N_866);
nand U935 (N_935,N_865,N_860);
xnor U936 (N_936,N_879,N_886);
nor U937 (N_937,N_865,N_855);
nand U938 (N_938,N_888,N_891);
and U939 (N_939,N_878,N_895);
nor U940 (N_940,N_863,N_896);
xor U941 (N_941,N_887,N_873);
nor U942 (N_942,N_898,N_865);
or U943 (N_943,N_881,N_894);
nor U944 (N_944,N_893,N_888);
nor U945 (N_945,N_866,N_852);
xnor U946 (N_946,N_878,N_854);
nor U947 (N_947,N_886,N_874);
nand U948 (N_948,N_897,N_855);
nor U949 (N_949,N_874,N_869);
nand U950 (N_950,N_941,N_902);
xnor U951 (N_951,N_924,N_939);
nand U952 (N_952,N_912,N_945);
xor U953 (N_953,N_926,N_921);
and U954 (N_954,N_942,N_907);
or U955 (N_955,N_937,N_943);
xor U956 (N_956,N_905,N_922);
nand U957 (N_957,N_919,N_925);
or U958 (N_958,N_906,N_944);
nor U959 (N_959,N_932,N_928);
or U960 (N_960,N_913,N_915);
nand U961 (N_961,N_935,N_938);
xor U962 (N_962,N_916,N_949);
nand U963 (N_963,N_920,N_910);
or U964 (N_964,N_908,N_934);
xnor U965 (N_965,N_947,N_917);
nand U966 (N_966,N_909,N_933);
and U967 (N_967,N_946,N_948);
or U968 (N_968,N_936,N_900);
xor U969 (N_969,N_923,N_927);
or U970 (N_970,N_930,N_901);
nand U971 (N_971,N_931,N_914);
and U972 (N_972,N_911,N_929);
nand U973 (N_973,N_918,N_940);
nand U974 (N_974,N_904,N_903);
and U975 (N_975,N_912,N_930);
nor U976 (N_976,N_947,N_948);
nor U977 (N_977,N_909,N_915);
or U978 (N_978,N_933,N_946);
nand U979 (N_979,N_918,N_907);
xnor U980 (N_980,N_948,N_903);
or U981 (N_981,N_925,N_909);
nand U982 (N_982,N_928,N_926);
nand U983 (N_983,N_940,N_949);
nor U984 (N_984,N_904,N_913);
xnor U985 (N_985,N_917,N_906);
and U986 (N_986,N_945,N_935);
xnor U987 (N_987,N_937,N_905);
nor U988 (N_988,N_941,N_924);
nand U989 (N_989,N_938,N_911);
or U990 (N_990,N_947,N_924);
nor U991 (N_991,N_933,N_913);
xnor U992 (N_992,N_929,N_901);
xor U993 (N_993,N_903,N_902);
and U994 (N_994,N_946,N_905);
and U995 (N_995,N_923,N_926);
or U996 (N_996,N_935,N_918);
and U997 (N_997,N_938,N_943);
or U998 (N_998,N_903,N_946);
nand U999 (N_999,N_926,N_905);
or U1000 (N_1000,N_969,N_972);
xor U1001 (N_1001,N_971,N_954);
or U1002 (N_1002,N_968,N_970);
or U1003 (N_1003,N_991,N_987);
nand U1004 (N_1004,N_985,N_992);
and U1005 (N_1005,N_960,N_961);
and U1006 (N_1006,N_963,N_973);
and U1007 (N_1007,N_958,N_993);
nor U1008 (N_1008,N_959,N_967);
nand U1009 (N_1009,N_986,N_950);
nand U1010 (N_1010,N_984,N_998);
or U1011 (N_1011,N_962,N_955);
or U1012 (N_1012,N_957,N_964);
nand U1013 (N_1013,N_980,N_981);
xnor U1014 (N_1014,N_953,N_977);
nand U1015 (N_1015,N_965,N_989);
nor U1016 (N_1016,N_951,N_956);
nand U1017 (N_1017,N_983,N_994);
or U1018 (N_1018,N_990,N_966);
or U1019 (N_1019,N_975,N_952);
or U1020 (N_1020,N_995,N_988);
nor U1021 (N_1021,N_976,N_978);
nand U1022 (N_1022,N_997,N_996);
nor U1023 (N_1023,N_974,N_982);
or U1024 (N_1024,N_979,N_999);
nor U1025 (N_1025,N_990,N_983);
and U1026 (N_1026,N_984,N_960);
nor U1027 (N_1027,N_987,N_961);
nand U1028 (N_1028,N_969,N_998);
nor U1029 (N_1029,N_988,N_994);
nor U1030 (N_1030,N_962,N_970);
nor U1031 (N_1031,N_990,N_956);
nor U1032 (N_1032,N_953,N_987);
or U1033 (N_1033,N_988,N_973);
nand U1034 (N_1034,N_980,N_954);
nor U1035 (N_1035,N_958,N_985);
xnor U1036 (N_1036,N_968,N_962);
or U1037 (N_1037,N_987,N_977);
or U1038 (N_1038,N_959,N_955);
nand U1039 (N_1039,N_995,N_951);
nor U1040 (N_1040,N_996,N_986);
xor U1041 (N_1041,N_950,N_999);
nand U1042 (N_1042,N_952,N_960);
and U1043 (N_1043,N_993,N_969);
nand U1044 (N_1044,N_986,N_976);
or U1045 (N_1045,N_978,N_955);
nand U1046 (N_1046,N_971,N_962);
nand U1047 (N_1047,N_999,N_987);
nor U1048 (N_1048,N_965,N_952);
xnor U1049 (N_1049,N_959,N_991);
or U1050 (N_1050,N_1047,N_1043);
and U1051 (N_1051,N_1015,N_1008);
xor U1052 (N_1052,N_1005,N_1009);
or U1053 (N_1053,N_1034,N_1003);
nand U1054 (N_1054,N_1032,N_1004);
xnor U1055 (N_1055,N_1049,N_1018);
or U1056 (N_1056,N_1022,N_1010);
nor U1057 (N_1057,N_1035,N_1038);
nand U1058 (N_1058,N_1025,N_1014);
and U1059 (N_1059,N_1021,N_1020);
nor U1060 (N_1060,N_1002,N_1006);
or U1061 (N_1061,N_1016,N_1024);
nand U1062 (N_1062,N_1033,N_1030);
nand U1063 (N_1063,N_1044,N_1040);
nand U1064 (N_1064,N_1001,N_1013);
xor U1065 (N_1065,N_1048,N_1031);
nand U1066 (N_1066,N_1023,N_1037);
nand U1067 (N_1067,N_1000,N_1045);
nand U1068 (N_1068,N_1036,N_1019);
nand U1069 (N_1069,N_1028,N_1042);
nor U1070 (N_1070,N_1041,N_1039);
nand U1071 (N_1071,N_1011,N_1026);
nand U1072 (N_1072,N_1029,N_1017);
xor U1073 (N_1073,N_1012,N_1027);
xnor U1074 (N_1074,N_1046,N_1007);
or U1075 (N_1075,N_1002,N_1007);
xor U1076 (N_1076,N_1004,N_1023);
nor U1077 (N_1077,N_1013,N_1046);
and U1078 (N_1078,N_1026,N_1046);
xor U1079 (N_1079,N_1041,N_1026);
nor U1080 (N_1080,N_1031,N_1009);
nand U1081 (N_1081,N_1048,N_1043);
nand U1082 (N_1082,N_1040,N_1049);
nand U1083 (N_1083,N_1046,N_1047);
xnor U1084 (N_1084,N_1001,N_1017);
and U1085 (N_1085,N_1037,N_1015);
and U1086 (N_1086,N_1017,N_1031);
xor U1087 (N_1087,N_1028,N_1031);
and U1088 (N_1088,N_1022,N_1040);
and U1089 (N_1089,N_1022,N_1035);
and U1090 (N_1090,N_1028,N_1019);
xnor U1091 (N_1091,N_1015,N_1023);
or U1092 (N_1092,N_1031,N_1035);
nand U1093 (N_1093,N_1031,N_1032);
or U1094 (N_1094,N_1001,N_1029);
xnor U1095 (N_1095,N_1008,N_1048);
and U1096 (N_1096,N_1011,N_1033);
xor U1097 (N_1097,N_1032,N_1021);
and U1098 (N_1098,N_1008,N_1016);
nand U1099 (N_1099,N_1005,N_1032);
xor U1100 (N_1100,N_1056,N_1094);
xnor U1101 (N_1101,N_1055,N_1091);
or U1102 (N_1102,N_1069,N_1063);
and U1103 (N_1103,N_1084,N_1076);
or U1104 (N_1104,N_1082,N_1093);
or U1105 (N_1105,N_1064,N_1090);
and U1106 (N_1106,N_1073,N_1068);
and U1107 (N_1107,N_1099,N_1061);
and U1108 (N_1108,N_1053,N_1054);
xor U1109 (N_1109,N_1086,N_1065);
and U1110 (N_1110,N_1085,N_1052);
and U1111 (N_1111,N_1050,N_1095);
or U1112 (N_1112,N_1097,N_1060);
or U1113 (N_1113,N_1074,N_1098);
or U1114 (N_1114,N_1066,N_1058);
nand U1115 (N_1115,N_1051,N_1080);
xnor U1116 (N_1116,N_1071,N_1059);
xnor U1117 (N_1117,N_1096,N_1067);
nor U1118 (N_1118,N_1092,N_1075);
nand U1119 (N_1119,N_1070,N_1089);
and U1120 (N_1120,N_1083,N_1079);
or U1121 (N_1121,N_1088,N_1087);
and U1122 (N_1122,N_1072,N_1078);
nand U1123 (N_1123,N_1057,N_1081);
and U1124 (N_1124,N_1062,N_1077);
xor U1125 (N_1125,N_1076,N_1095);
or U1126 (N_1126,N_1075,N_1068);
and U1127 (N_1127,N_1088,N_1068);
or U1128 (N_1128,N_1098,N_1094);
or U1129 (N_1129,N_1052,N_1078);
or U1130 (N_1130,N_1061,N_1068);
and U1131 (N_1131,N_1094,N_1072);
nor U1132 (N_1132,N_1065,N_1097);
nand U1133 (N_1133,N_1085,N_1065);
and U1134 (N_1134,N_1050,N_1098);
nand U1135 (N_1135,N_1054,N_1062);
or U1136 (N_1136,N_1065,N_1083);
and U1137 (N_1137,N_1094,N_1077);
and U1138 (N_1138,N_1062,N_1081);
xnor U1139 (N_1139,N_1067,N_1086);
and U1140 (N_1140,N_1069,N_1061);
nand U1141 (N_1141,N_1070,N_1080);
and U1142 (N_1142,N_1068,N_1080);
nand U1143 (N_1143,N_1090,N_1099);
nor U1144 (N_1144,N_1097,N_1059);
or U1145 (N_1145,N_1085,N_1078);
nor U1146 (N_1146,N_1077,N_1089);
nor U1147 (N_1147,N_1054,N_1076);
or U1148 (N_1148,N_1086,N_1052);
xor U1149 (N_1149,N_1057,N_1070);
and U1150 (N_1150,N_1116,N_1111);
and U1151 (N_1151,N_1100,N_1135);
and U1152 (N_1152,N_1121,N_1144);
or U1153 (N_1153,N_1102,N_1136);
or U1154 (N_1154,N_1137,N_1118);
nor U1155 (N_1155,N_1104,N_1103);
or U1156 (N_1156,N_1131,N_1128);
xnor U1157 (N_1157,N_1114,N_1145);
nor U1158 (N_1158,N_1147,N_1129);
nand U1159 (N_1159,N_1124,N_1133);
or U1160 (N_1160,N_1148,N_1141);
or U1161 (N_1161,N_1106,N_1132);
xnor U1162 (N_1162,N_1110,N_1125);
and U1163 (N_1163,N_1122,N_1146);
and U1164 (N_1164,N_1139,N_1101);
nand U1165 (N_1165,N_1138,N_1126);
and U1166 (N_1166,N_1105,N_1107);
and U1167 (N_1167,N_1134,N_1113);
or U1168 (N_1168,N_1140,N_1117);
or U1169 (N_1169,N_1130,N_1127);
or U1170 (N_1170,N_1149,N_1109);
xor U1171 (N_1171,N_1143,N_1142);
nor U1172 (N_1172,N_1112,N_1123);
nor U1173 (N_1173,N_1119,N_1108);
nand U1174 (N_1174,N_1115,N_1120);
or U1175 (N_1175,N_1144,N_1136);
xor U1176 (N_1176,N_1103,N_1143);
nand U1177 (N_1177,N_1134,N_1131);
and U1178 (N_1178,N_1148,N_1142);
nand U1179 (N_1179,N_1148,N_1127);
nor U1180 (N_1180,N_1129,N_1108);
nor U1181 (N_1181,N_1146,N_1133);
and U1182 (N_1182,N_1130,N_1111);
or U1183 (N_1183,N_1141,N_1132);
xnor U1184 (N_1184,N_1110,N_1120);
or U1185 (N_1185,N_1136,N_1139);
xor U1186 (N_1186,N_1145,N_1131);
nor U1187 (N_1187,N_1112,N_1104);
and U1188 (N_1188,N_1121,N_1101);
nand U1189 (N_1189,N_1102,N_1144);
nor U1190 (N_1190,N_1124,N_1131);
or U1191 (N_1191,N_1141,N_1117);
nand U1192 (N_1192,N_1119,N_1104);
xor U1193 (N_1193,N_1107,N_1114);
nor U1194 (N_1194,N_1140,N_1125);
or U1195 (N_1195,N_1128,N_1142);
or U1196 (N_1196,N_1146,N_1116);
nand U1197 (N_1197,N_1145,N_1100);
and U1198 (N_1198,N_1139,N_1118);
and U1199 (N_1199,N_1114,N_1113);
nor U1200 (N_1200,N_1190,N_1152);
and U1201 (N_1201,N_1180,N_1172);
nand U1202 (N_1202,N_1183,N_1186);
xor U1203 (N_1203,N_1160,N_1157);
or U1204 (N_1204,N_1167,N_1164);
xor U1205 (N_1205,N_1168,N_1182);
nand U1206 (N_1206,N_1185,N_1177);
xor U1207 (N_1207,N_1198,N_1194);
nand U1208 (N_1208,N_1179,N_1192);
xor U1209 (N_1209,N_1189,N_1188);
nand U1210 (N_1210,N_1162,N_1169);
nor U1211 (N_1211,N_1184,N_1156);
or U1212 (N_1212,N_1163,N_1154);
nor U1213 (N_1213,N_1153,N_1170);
and U1214 (N_1214,N_1176,N_1197);
and U1215 (N_1215,N_1199,N_1196);
nand U1216 (N_1216,N_1158,N_1166);
and U1217 (N_1217,N_1175,N_1173);
nand U1218 (N_1218,N_1181,N_1171);
or U1219 (N_1219,N_1165,N_1187);
xor U1220 (N_1220,N_1174,N_1161);
and U1221 (N_1221,N_1155,N_1191);
or U1222 (N_1222,N_1195,N_1193);
xor U1223 (N_1223,N_1151,N_1159);
nand U1224 (N_1224,N_1178,N_1150);
nand U1225 (N_1225,N_1181,N_1162);
or U1226 (N_1226,N_1151,N_1176);
xor U1227 (N_1227,N_1175,N_1176);
nor U1228 (N_1228,N_1176,N_1162);
and U1229 (N_1229,N_1160,N_1191);
nand U1230 (N_1230,N_1185,N_1182);
nor U1231 (N_1231,N_1150,N_1165);
or U1232 (N_1232,N_1183,N_1189);
xor U1233 (N_1233,N_1179,N_1172);
nor U1234 (N_1234,N_1167,N_1183);
or U1235 (N_1235,N_1162,N_1175);
xnor U1236 (N_1236,N_1160,N_1159);
and U1237 (N_1237,N_1156,N_1190);
nor U1238 (N_1238,N_1198,N_1181);
nand U1239 (N_1239,N_1183,N_1174);
or U1240 (N_1240,N_1179,N_1166);
or U1241 (N_1241,N_1173,N_1160);
nor U1242 (N_1242,N_1157,N_1154);
nor U1243 (N_1243,N_1187,N_1151);
and U1244 (N_1244,N_1163,N_1194);
or U1245 (N_1245,N_1179,N_1156);
and U1246 (N_1246,N_1178,N_1173);
nor U1247 (N_1247,N_1197,N_1151);
nor U1248 (N_1248,N_1163,N_1195);
xnor U1249 (N_1249,N_1182,N_1169);
and U1250 (N_1250,N_1212,N_1246);
nand U1251 (N_1251,N_1210,N_1248);
nor U1252 (N_1252,N_1244,N_1215);
xor U1253 (N_1253,N_1202,N_1208);
and U1254 (N_1254,N_1203,N_1245);
nand U1255 (N_1255,N_1249,N_1219);
xor U1256 (N_1256,N_1240,N_1220);
xnor U1257 (N_1257,N_1207,N_1235);
and U1258 (N_1258,N_1221,N_1247);
and U1259 (N_1259,N_1238,N_1216);
and U1260 (N_1260,N_1223,N_1224);
nand U1261 (N_1261,N_1236,N_1242);
and U1262 (N_1262,N_1201,N_1218);
and U1263 (N_1263,N_1205,N_1241);
and U1264 (N_1264,N_1226,N_1232);
and U1265 (N_1265,N_1211,N_1214);
xor U1266 (N_1266,N_1234,N_1243);
and U1267 (N_1267,N_1228,N_1206);
or U1268 (N_1268,N_1225,N_1209);
nor U1269 (N_1269,N_1230,N_1213);
and U1270 (N_1270,N_1233,N_1239);
xnor U1271 (N_1271,N_1222,N_1229);
and U1272 (N_1272,N_1204,N_1227);
or U1273 (N_1273,N_1217,N_1231);
nor U1274 (N_1274,N_1237,N_1200);
nand U1275 (N_1275,N_1232,N_1228);
and U1276 (N_1276,N_1223,N_1206);
and U1277 (N_1277,N_1235,N_1236);
or U1278 (N_1278,N_1231,N_1243);
xnor U1279 (N_1279,N_1223,N_1233);
nor U1280 (N_1280,N_1218,N_1211);
nand U1281 (N_1281,N_1205,N_1240);
nor U1282 (N_1282,N_1220,N_1211);
xnor U1283 (N_1283,N_1223,N_1212);
or U1284 (N_1284,N_1246,N_1222);
or U1285 (N_1285,N_1224,N_1235);
or U1286 (N_1286,N_1248,N_1205);
nand U1287 (N_1287,N_1234,N_1230);
nand U1288 (N_1288,N_1229,N_1217);
and U1289 (N_1289,N_1221,N_1235);
or U1290 (N_1290,N_1224,N_1231);
or U1291 (N_1291,N_1229,N_1213);
xnor U1292 (N_1292,N_1244,N_1223);
and U1293 (N_1293,N_1200,N_1210);
or U1294 (N_1294,N_1229,N_1232);
or U1295 (N_1295,N_1228,N_1212);
or U1296 (N_1296,N_1216,N_1240);
nor U1297 (N_1297,N_1200,N_1245);
and U1298 (N_1298,N_1200,N_1244);
or U1299 (N_1299,N_1248,N_1225);
and U1300 (N_1300,N_1252,N_1253);
xnor U1301 (N_1301,N_1290,N_1285);
nand U1302 (N_1302,N_1251,N_1266);
or U1303 (N_1303,N_1299,N_1264);
or U1304 (N_1304,N_1294,N_1261);
or U1305 (N_1305,N_1279,N_1258);
and U1306 (N_1306,N_1259,N_1272);
or U1307 (N_1307,N_1282,N_1283);
nand U1308 (N_1308,N_1254,N_1274);
nor U1309 (N_1309,N_1260,N_1277);
or U1310 (N_1310,N_1269,N_1271);
nand U1311 (N_1311,N_1298,N_1287);
xnor U1312 (N_1312,N_1257,N_1292);
xor U1313 (N_1313,N_1275,N_1256);
nor U1314 (N_1314,N_1278,N_1288);
and U1315 (N_1315,N_1268,N_1284);
nand U1316 (N_1316,N_1297,N_1295);
and U1317 (N_1317,N_1280,N_1293);
nor U1318 (N_1318,N_1296,N_1267);
nor U1319 (N_1319,N_1281,N_1270);
xor U1320 (N_1320,N_1291,N_1289);
nor U1321 (N_1321,N_1263,N_1262);
nand U1322 (N_1322,N_1276,N_1255);
and U1323 (N_1323,N_1250,N_1265);
or U1324 (N_1324,N_1273,N_1286);
xor U1325 (N_1325,N_1299,N_1273);
and U1326 (N_1326,N_1292,N_1297);
nor U1327 (N_1327,N_1251,N_1283);
and U1328 (N_1328,N_1255,N_1261);
nand U1329 (N_1329,N_1270,N_1289);
nand U1330 (N_1330,N_1277,N_1256);
and U1331 (N_1331,N_1287,N_1275);
nor U1332 (N_1332,N_1275,N_1295);
nor U1333 (N_1333,N_1269,N_1274);
and U1334 (N_1334,N_1266,N_1280);
and U1335 (N_1335,N_1289,N_1256);
or U1336 (N_1336,N_1263,N_1289);
and U1337 (N_1337,N_1272,N_1297);
and U1338 (N_1338,N_1274,N_1286);
nand U1339 (N_1339,N_1281,N_1264);
nor U1340 (N_1340,N_1262,N_1292);
nand U1341 (N_1341,N_1290,N_1284);
nand U1342 (N_1342,N_1268,N_1287);
nand U1343 (N_1343,N_1264,N_1292);
xnor U1344 (N_1344,N_1284,N_1299);
or U1345 (N_1345,N_1266,N_1253);
nand U1346 (N_1346,N_1297,N_1267);
and U1347 (N_1347,N_1250,N_1281);
xor U1348 (N_1348,N_1265,N_1264);
or U1349 (N_1349,N_1266,N_1296);
or U1350 (N_1350,N_1347,N_1310);
and U1351 (N_1351,N_1309,N_1340);
and U1352 (N_1352,N_1341,N_1345);
xor U1353 (N_1353,N_1331,N_1332);
xor U1354 (N_1354,N_1311,N_1321);
xor U1355 (N_1355,N_1328,N_1317);
xnor U1356 (N_1356,N_1304,N_1303);
nor U1357 (N_1357,N_1320,N_1324);
and U1358 (N_1358,N_1307,N_1344);
nor U1359 (N_1359,N_1330,N_1326);
or U1360 (N_1360,N_1336,N_1313);
and U1361 (N_1361,N_1318,N_1315);
nand U1362 (N_1362,N_1337,N_1348);
nand U1363 (N_1363,N_1339,N_1302);
or U1364 (N_1364,N_1308,N_1334);
and U1365 (N_1365,N_1322,N_1316);
nand U1366 (N_1366,N_1314,N_1349);
nor U1367 (N_1367,N_1342,N_1325);
nand U1368 (N_1368,N_1333,N_1319);
xnor U1369 (N_1369,N_1300,N_1305);
or U1370 (N_1370,N_1312,N_1306);
nand U1371 (N_1371,N_1301,N_1343);
nor U1372 (N_1372,N_1327,N_1335);
and U1373 (N_1373,N_1346,N_1338);
or U1374 (N_1374,N_1323,N_1329);
or U1375 (N_1375,N_1324,N_1301);
and U1376 (N_1376,N_1344,N_1312);
nand U1377 (N_1377,N_1320,N_1336);
nand U1378 (N_1378,N_1314,N_1300);
nor U1379 (N_1379,N_1337,N_1305);
and U1380 (N_1380,N_1308,N_1346);
nor U1381 (N_1381,N_1314,N_1309);
xor U1382 (N_1382,N_1307,N_1349);
and U1383 (N_1383,N_1330,N_1340);
and U1384 (N_1384,N_1331,N_1321);
nor U1385 (N_1385,N_1335,N_1337);
or U1386 (N_1386,N_1332,N_1312);
xor U1387 (N_1387,N_1349,N_1334);
and U1388 (N_1388,N_1331,N_1316);
and U1389 (N_1389,N_1303,N_1328);
nand U1390 (N_1390,N_1335,N_1349);
and U1391 (N_1391,N_1339,N_1324);
nand U1392 (N_1392,N_1306,N_1314);
xnor U1393 (N_1393,N_1345,N_1324);
nor U1394 (N_1394,N_1323,N_1302);
xnor U1395 (N_1395,N_1333,N_1310);
and U1396 (N_1396,N_1324,N_1314);
or U1397 (N_1397,N_1320,N_1307);
xnor U1398 (N_1398,N_1311,N_1345);
nor U1399 (N_1399,N_1314,N_1315);
xor U1400 (N_1400,N_1384,N_1357);
xor U1401 (N_1401,N_1388,N_1360);
and U1402 (N_1402,N_1370,N_1364);
nor U1403 (N_1403,N_1359,N_1391);
nor U1404 (N_1404,N_1378,N_1381);
nor U1405 (N_1405,N_1363,N_1393);
nand U1406 (N_1406,N_1383,N_1395);
and U1407 (N_1407,N_1353,N_1394);
and U1408 (N_1408,N_1355,N_1366);
and U1409 (N_1409,N_1387,N_1371);
and U1410 (N_1410,N_1386,N_1397);
or U1411 (N_1411,N_1367,N_1382);
nor U1412 (N_1412,N_1389,N_1390);
and U1413 (N_1413,N_1385,N_1369);
and U1414 (N_1414,N_1373,N_1365);
nor U1415 (N_1415,N_1361,N_1376);
nor U1416 (N_1416,N_1396,N_1399);
nor U1417 (N_1417,N_1354,N_1358);
nand U1418 (N_1418,N_1350,N_1380);
nor U1419 (N_1419,N_1392,N_1374);
nand U1420 (N_1420,N_1352,N_1398);
or U1421 (N_1421,N_1362,N_1375);
or U1422 (N_1422,N_1351,N_1368);
or U1423 (N_1423,N_1356,N_1377);
or U1424 (N_1424,N_1379,N_1372);
xnor U1425 (N_1425,N_1388,N_1352);
nor U1426 (N_1426,N_1384,N_1378);
xnor U1427 (N_1427,N_1352,N_1353);
nor U1428 (N_1428,N_1384,N_1362);
and U1429 (N_1429,N_1365,N_1374);
and U1430 (N_1430,N_1366,N_1386);
or U1431 (N_1431,N_1391,N_1382);
and U1432 (N_1432,N_1353,N_1354);
xor U1433 (N_1433,N_1359,N_1367);
and U1434 (N_1434,N_1378,N_1369);
nand U1435 (N_1435,N_1388,N_1390);
xnor U1436 (N_1436,N_1387,N_1356);
and U1437 (N_1437,N_1389,N_1374);
nand U1438 (N_1438,N_1375,N_1376);
xnor U1439 (N_1439,N_1371,N_1390);
and U1440 (N_1440,N_1351,N_1396);
nand U1441 (N_1441,N_1391,N_1395);
or U1442 (N_1442,N_1385,N_1357);
and U1443 (N_1443,N_1354,N_1382);
nand U1444 (N_1444,N_1381,N_1387);
xor U1445 (N_1445,N_1382,N_1394);
and U1446 (N_1446,N_1375,N_1387);
nand U1447 (N_1447,N_1350,N_1363);
nand U1448 (N_1448,N_1390,N_1367);
nand U1449 (N_1449,N_1390,N_1372);
and U1450 (N_1450,N_1417,N_1428);
xor U1451 (N_1451,N_1419,N_1447);
xnor U1452 (N_1452,N_1415,N_1409);
or U1453 (N_1453,N_1410,N_1401);
xor U1454 (N_1454,N_1406,N_1438);
nor U1455 (N_1455,N_1425,N_1432);
nor U1456 (N_1456,N_1402,N_1449);
and U1457 (N_1457,N_1400,N_1411);
and U1458 (N_1458,N_1443,N_1403);
nand U1459 (N_1459,N_1416,N_1448);
xor U1460 (N_1460,N_1433,N_1408);
nor U1461 (N_1461,N_1434,N_1444);
or U1462 (N_1462,N_1441,N_1407);
or U1463 (N_1463,N_1446,N_1412);
or U1464 (N_1464,N_1423,N_1435);
nand U1465 (N_1465,N_1426,N_1413);
nand U1466 (N_1466,N_1424,N_1405);
nand U1467 (N_1467,N_1431,N_1440);
nand U1468 (N_1468,N_1445,N_1414);
nand U1469 (N_1469,N_1421,N_1418);
nand U1470 (N_1470,N_1427,N_1436);
or U1471 (N_1471,N_1420,N_1429);
nand U1472 (N_1472,N_1422,N_1439);
and U1473 (N_1473,N_1442,N_1404);
nand U1474 (N_1474,N_1430,N_1437);
nor U1475 (N_1475,N_1430,N_1402);
and U1476 (N_1476,N_1429,N_1445);
nor U1477 (N_1477,N_1441,N_1418);
nand U1478 (N_1478,N_1406,N_1407);
nor U1479 (N_1479,N_1443,N_1417);
nand U1480 (N_1480,N_1406,N_1447);
nand U1481 (N_1481,N_1434,N_1440);
xnor U1482 (N_1482,N_1443,N_1430);
or U1483 (N_1483,N_1400,N_1408);
xnor U1484 (N_1484,N_1409,N_1403);
nor U1485 (N_1485,N_1426,N_1427);
nand U1486 (N_1486,N_1405,N_1430);
xnor U1487 (N_1487,N_1422,N_1448);
nor U1488 (N_1488,N_1413,N_1442);
xor U1489 (N_1489,N_1434,N_1445);
and U1490 (N_1490,N_1434,N_1442);
or U1491 (N_1491,N_1400,N_1403);
nor U1492 (N_1492,N_1424,N_1442);
xnor U1493 (N_1493,N_1402,N_1400);
nor U1494 (N_1494,N_1420,N_1414);
or U1495 (N_1495,N_1422,N_1406);
xor U1496 (N_1496,N_1447,N_1432);
and U1497 (N_1497,N_1431,N_1402);
xnor U1498 (N_1498,N_1430,N_1410);
and U1499 (N_1499,N_1415,N_1418);
or U1500 (N_1500,N_1486,N_1498);
nand U1501 (N_1501,N_1459,N_1463);
and U1502 (N_1502,N_1497,N_1469);
and U1503 (N_1503,N_1475,N_1468);
or U1504 (N_1504,N_1461,N_1460);
xor U1505 (N_1505,N_1458,N_1491);
or U1506 (N_1506,N_1485,N_1487);
xnor U1507 (N_1507,N_1499,N_1454);
nand U1508 (N_1508,N_1465,N_1457);
nor U1509 (N_1509,N_1466,N_1493);
xor U1510 (N_1510,N_1451,N_1484);
xor U1511 (N_1511,N_1450,N_1489);
nor U1512 (N_1512,N_1477,N_1464);
nor U1513 (N_1513,N_1453,N_1479);
nor U1514 (N_1514,N_1456,N_1472);
nor U1515 (N_1515,N_1476,N_1480);
or U1516 (N_1516,N_1482,N_1494);
xnor U1517 (N_1517,N_1462,N_1495);
nor U1518 (N_1518,N_1452,N_1490);
and U1519 (N_1519,N_1455,N_1473);
and U1520 (N_1520,N_1496,N_1488);
nand U1521 (N_1521,N_1492,N_1478);
nand U1522 (N_1522,N_1483,N_1467);
and U1523 (N_1523,N_1481,N_1474);
nor U1524 (N_1524,N_1470,N_1471);
and U1525 (N_1525,N_1491,N_1455);
nor U1526 (N_1526,N_1495,N_1464);
and U1527 (N_1527,N_1495,N_1472);
and U1528 (N_1528,N_1466,N_1498);
nand U1529 (N_1529,N_1455,N_1499);
xor U1530 (N_1530,N_1498,N_1454);
and U1531 (N_1531,N_1450,N_1462);
or U1532 (N_1532,N_1492,N_1472);
or U1533 (N_1533,N_1480,N_1461);
or U1534 (N_1534,N_1465,N_1485);
nand U1535 (N_1535,N_1456,N_1497);
and U1536 (N_1536,N_1454,N_1467);
nand U1537 (N_1537,N_1497,N_1457);
nor U1538 (N_1538,N_1469,N_1452);
xnor U1539 (N_1539,N_1487,N_1458);
or U1540 (N_1540,N_1493,N_1478);
nor U1541 (N_1541,N_1494,N_1450);
nor U1542 (N_1542,N_1485,N_1472);
xor U1543 (N_1543,N_1473,N_1485);
nand U1544 (N_1544,N_1466,N_1472);
or U1545 (N_1545,N_1485,N_1470);
xor U1546 (N_1546,N_1466,N_1495);
and U1547 (N_1547,N_1474,N_1465);
nor U1548 (N_1548,N_1478,N_1469);
nor U1549 (N_1549,N_1491,N_1492);
nand U1550 (N_1550,N_1541,N_1549);
or U1551 (N_1551,N_1522,N_1543);
nor U1552 (N_1552,N_1529,N_1506);
xnor U1553 (N_1553,N_1502,N_1537);
nor U1554 (N_1554,N_1544,N_1518);
or U1555 (N_1555,N_1525,N_1509);
nand U1556 (N_1556,N_1533,N_1528);
and U1557 (N_1557,N_1536,N_1534);
nor U1558 (N_1558,N_1515,N_1527);
nor U1559 (N_1559,N_1507,N_1514);
nand U1560 (N_1560,N_1530,N_1532);
or U1561 (N_1561,N_1519,N_1531);
nor U1562 (N_1562,N_1501,N_1535);
nand U1563 (N_1563,N_1523,N_1500);
nor U1564 (N_1564,N_1542,N_1513);
nand U1565 (N_1565,N_1503,N_1511);
xor U1566 (N_1566,N_1521,N_1520);
and U1567 (N_1567,N_1504,N_1505);
nand U1568 (N_1568,N_1516,N_1546);
nor U1569 (N_1569,N_1538,N_1512);
or U1570 (N_1570,N_1526,N_1540);
xnor U1571 (N_1571,N_1548,N_1508);
xnor U1572 (N_1572,N_1517,N_1539);
nand U1573 (N_1573,N_1547,N_1545);
nand U1574 (N_1574,N_1524,N_1510);
nand U1575 (N_1575,N_1532,N_1535);
nor U1576 (N_1576,N_1510,N_1545);
nand U1577 (N_1577,N_1508,N_1505);
xnor U1578 (N_1578,N_1538,N_1533);
nand U1579 (N_1579,N_1508,N_1529);
nor U1580 (N_1580,N_1503,N_1521);
xnor U1581 (N_1581,N_1547,N_1529);
and U1582 (N_1582,N_1530,N_1539);
and U1583 (N_1583,N_1522,N_1544);
nand U1584 (N_1584,N_1505,N_1523);
xnor U1585 (N_1585,N_1521,N_1516);
xnor U1586 (N_1586,N_1527,N_1530);
nor U1587 (N_1587,N_1532,N_1539);
nand U1588 (N_1588,N_1531,N_1547);
and U1589 (N_1589,N_1538,N_1536);
and U1590 (N_1590,N_1520,N_1507);
nor U1591 (N_1591,N_1510,N_1544);
or U1592 (N_1592,N_1547,N_1532);
or U1593 (N_1593,N_1519,N_1532);
nand U1594 (N_1594,N_1516,N_1535);
nand U1595 (N_1595,N_1508,N_1546);
and U1596 (N_1596,N_1501,N_1549);
nor U1597 (N_1597,N_1505,N_1544);
nor U1598 (N_1598,N_1538,N_1526);
xnor U1599 (N_1599,N_1505,N_1548);
nand U1600 (N_1600,N_1570,N_1577);
nand U1601 (N_1601,N_1589,N_1593);
nor U1602 (N_1602,N_1573,N_1588);
or U1603 (N_1603,N_1590,N_1563);
xor U1604 (N_1604,N_1591,N_1585);
or U1605 (N_1605,N_1596,N_1581);
nor U1606 (N_1606,N_1560,N_1599);
or U1607 (N_1607,N_1583,N_1565);
or U1608 (N_1608,N_1566,N_1587);
nand U1609 (N_1609,N_1575,N_1559);
xor U1610 (N_1610,N_1562,N_1578);
nand U1611 (N_1611,N_1550,N_1582);
nor U1612 (N_1612,N_1584,N_1592);
xnor U1613 (N_1613,N_1598,N_1576);
and U1614 (N_1614,N_1557,N_1595);
and U1615 (N_1615,N_1551,N_1567);
or U1616 (N_1616,N_1555,N_1597);
and U1617 (N_1617,N_1572,N_1554);
nor U1618 (N_1618,N_1561,N_1586);
and U1619 (N_1619,N_1571,N_1556);
nand U1620 (N_1620,N_1594,N_1580);
or U1621 (N_1621,N_1579,N_1569);
nand U1622 (N_1622,N_1553,N_1558);
nor U1623 (N_1623,N_1568,N_1552);
and U1624 (N_1624,N_1574,N_1564);
or U1625 (N_1625,N_1555,N_1562);
or U1626 (N_1626,N_1560,N_1580);
nor U1627 (N_1627,N_1593,N_1551);
xnor U1628 (N_1628,N_1552,N_1579);
nand U1629 (N_1629,N_1566,N_1554);
xor U1630 (N_1630,N_1587,N_1580);
xor U1631 (N_1631,N_1569,N_1582);
or U1632 (N_1632,N_1565,N_1557);
nor U1633 (N_1633,N_1565,N_1589);
xnor U1634 (N_1634,N_1558,N_1562);
or U1635 (N_1635,N_1580,N_1596);
and U1636 (N_1636,N_1559,N_1555);
or U1637 (N_1637,N_1569,N_1599);
and U1638 (N_1638,N_1555,N_1550);
and U1639 (N_1639,N_1583,N_1581);
nor U1640 (N_1640,N_1569,N_1561);
or U1641 (N_1641,N_1572,N_1553);
nand U1642 (N_1642,N_1565,N_1578);
or U1643 (N_1643,N_1591,N_1574);
xor U1644 (N_1644,N_1558,N_1552);
nand U1645 (N_1645,N_1566,N_1590);
and U1646 (N_1646,N_1578,N_1567);
nor U1647 (N_1647,N_1583,N_1597);
nor U1648 (N_1648,N_1592,N_1598);
nand U1649 (N_1649,N_1550,N_1583);
nor U1650 (N_1650,N_1628,N_1612);
xor U1651 (N_1651,N_1622,N_1646);
xor U1652 (N_1652,N_1643,N_1639);
xor U1653 (N_1653,N_1604,N_1621);
and U1654 (N_1654,N_1617,N_1644);
and U1655 (N_1655,N_1602,N_1611);
or U1656 (N_1656,N_1629,N_1605);
nand U1657 (N_1657,N_1614,N_1606);
nand U1658 (N_1658,N_1635,N_1645);
xor U1659 (N_1659,N_1633,N_1631);
and U1660 (N_1660,N_1648,N_1609);
nor U1661 (N_1661,N_1608,N_1625);
and U1662 (N_1662,N_1624,N_1623);
or U1663 (N_1663,N_1601,N_1636);
nor U1664 (N_1664,N_1618,N_1620);
and U1665 (N_1665,N_1610,N_1619);
xor U1666 (N_1666,N_1637,N_1616);
and U1667 (N_1667,N_1603,N_1626);
nand U1668 (N_1668,N_1600,N_1641);
nor U1669 (N_1669,N_1630,N_1615);
nor U1670 (N_1670,N_1649,N_1642);
or U1671 (N_1671,N_1632,N_1627);
and U1672 (N_1672,N_1640,N_1607);
nor U1673 (N_1673,N_1634,N_1638);
and U1674 (N_1674,N_1613,N_1647);
and U1675 (N_1675,N_1627,N_1639);
nor U1676 (N_1676,N_1631,N_1619);
and U1677 (N_1677,N_1642,N_1621);
nand U1678 (N_1678,N_1640,N_1645);
xnor U1679 (N_1679,N_1629,N_1613);
nor U1680 (N_1680,N_1623,N_1636);
xnor U1681 (N_1681,N_1609,N_1614);
xnor U1682 (N_1682,N_1606,N_1620);
nor U1683 (N_1683,N_1645,N_1611);
nand U1684 (N_1684,N_1613,N_1631);
or U1685 (N_1685,N_1638,N_1626);
xnor U1686 (N_1686,N_1625,N_1614);
nand U1687 (N_1687,N_1610,N_1637);
nand U1688 (N_1688,N_1630,N_1635);
nand U1689 (N_1689,N_1602,N_1644);
and U1690 (N_1690,N_1618,N_1615);
xor U1691 (N_1691,N_1615,N_1627);
and U1692 (N_1692,N_1613,N_1600);
nor U1693 (N_1693,N_1625,N_1646);
nand U1694 (N_1694,N_1600,N_1648);
xor U1695 (N_1695,N_1629,N_1630);
nor U1696 (N_1696,N_1604,N_1624);
and U1697 (N_1697,N_1640,N_1603);
nor U1698 (N_1698,N_1600,N_1628);
nand U1699 (N_1699,N_1613,N_1636);
and U1700 (N_1700,N_1696,N_1678);
and U1701 (N_1701,N_1680,N_1684);
or U1702 (N_1702,N_1659,N_1681);
and U1703 (N_1703,N_1652,N_1691);
or U1704 (N_1704,N_1686,N_1650);
nand U1705 (N_1705,N_1677,N_1683);
nor U1706 (N_1706,N_1661,N_1672);
or U1707 (N_1707,N_1662,N_1697);
xnor U1708 (N_1708,N_1653,N_1667);
nand U1709 (N_1709,N_1685,N_1695);
nor U1710 (N_1710,N_1676,N_1668);
or U1711 (N_1711,N_1689,N_1654);
or U1712 (N_1712,N_1690,N_1660);
nand U1713 (N_1713,N_1692,N_1655);
and U1714 (N_1714,N_1664,N_1674);
or U1715 (N_1715,N_1666,N_1693);
nor U1716 (N_1716,N_1656,N_1657);
or U1717 (N_1717,N_1698,N_1671);
nand U1718 (N_1718,N_1663,N_1665);
and U1719 (N_1719,N_1682,N_1679);
xor U1720 (N_1720,N_1687,N_1651);
and U1721 (N_1721,N_1669,N_1699);
nor U1722 (N_1722,N_1688,N_1673);
nor U1723 (N_1723,N_1694,N_1675);
or U1724 (N_1724,N_1658,N_1670);
xnor U1725 (N_1725,N_1698,N_1670);
and U1726 (N_1726,N_1660,N_1693);
and U1727 (N_1727,N_1697,N_1659);
xor U1728 (N_1728,N_1661,N_1676);
nor U1729 (N_1729,N_1661,N_1651);
nor U1730 (N_1730,N_1653,N_1665);
xor U1731 (N_1731,N_1697,N_1652);
nand U1732 (N_1732,N_1692,N_1650);
and U1733 (N_1733,N_1667,N_1692);
xor U1734 (N_1734,N_1662,N_1676);
xor U1735 (N_1735,N_1662,N_1671);
and U1736 (N_1736,N_1684,N_1658);
nor U1737 (N_1737,N_1660,N_1687);
nor U1738 (N_1738,N_1666,N_1652);
or U1739 (N_1739,N_1693,N_1668);
xnor U1740 (N_1740,N_1684,N_1678);
and U1741 (N_1741,N_1665,N_1671);
nand U1742 (N_1742,N_1659,N_1654);
nand U1743 (N_1743,N_1678,N_1665);
or U1744 (N_1744,N_1688,N_1694);
nor U1745 (N_1745,N_1654,N_1650);
nand U1746 (N_1746,N_1688,N_1672);
and U1747 (N_1747,N_1671,N_1678);
and U1748 (N_1748,N_1673,N_1657);
or U1749 (N_1749,N_1680,N_1666);
xnor U1750 (N_1750,N_1731,N_1727);
and U1751 (N_1751,N_1701,N_1743);
and U1752 (N_1752,N_1710,N_1749);
xor U1753 (N_1753,N_1737,N_1711);
xnor U1754 (N_1754,N_1746,N_1724);
nor U1755 (N_1755,N_1704,N_1712);
nand U1756 (N_1756,N_1707,N_1719);
and U1757 (N_1757,N_1729,N_1705);
xor U1758 (N_1758,N_1702,N_1735);
nand U1759 (N_1759,N_1740,N_1715);
nand U1760 (N_1760,N_1747,N_1721);
nor U1761 (N_1761,N_1722,N_1726);
nor U1762 (N_1762,N_1734,N_1745);
nand U1763 (N_1763,N_1744,N_1725);
or U1764 (N_1764,N_1748,N_1741);
or U1765 (N_1765,N_1739,N_1703);
or U1766 (N_1766,N_1706,N_1732);
or U1767 (N_1767,N_1742,N_1717);
xnor U1768 (N_1768,N_1700,N_1730);
xnor U1769 (N_1769,N_1723,N_1716);
nand U1770 (N_1770,N_1708,N_1736);
nor U1771 (N_1771,N_1733,N_1714);
xor U1772 (N_1772,N_1738,N_1728);
nor U1773 (N_1773,N_1720,N_1718);
xor U1774 (N_1774,N_1713,N_1709);
nand U1775 (N_1775,N_1737,N_1713);
nor U1776 (N_1776,N_1714,N_1708);
or U1777 (N_1777,N_1730,N_1737);
xor U1778 (N_1778,N_1713,N_1717);
and U1779 (N_1779,N_1724,N_1739);
xor U1780 (N_1780,N_1703,N_1708);
nand U1781 (N_1781,N_1744,N_1724);
nand U1782 (N_1782,N_1719,N_1731);
nand U1783 (N_1783,N_1733,N_1739);
or U1784 (N_1784,N_1702,N_1717);
nand U1785 (N_1785,N_1724,N_1735);
nor U1786 (N_1786,N_1712,N_1727);
or U1787 (N_1787,N_1742,N_1701);
nor U1788 (N_1788,N_1742,N_1721);
or U1789 (N_1789,N_1739,N_1746);
or U1790 (N_1790,N_1701,N_1738);
and U1791 (N_1791,N_1700,N_1738);
xor U1792 (N_1792,N_1737,N_1742);
or U1793 (N_1793,N_1733,N_1720);
and U1794 (N_1794,N_1730,N_1707);
xor U1795 (N_1795,N_1714,N_1726);
xnor U1796 (N_1796,N_1728,N_1737);
and U1797 (N_1797,N_1708,N_1728);
nand U1798 (N_1798,N_1721,N_1741);
nor U1799 (N_1799,N_1703,N_1706);
and U1800 (N_1800,N_1781,N_1754);
nand U1801 (N_1801,N_1773,N_1795);
xor U1802 (N_1802,N_1779,N_1752);
or U1803 (N_1803,N_1772,N_1796);
nand U1804 (N_1804,N_1797,N_1788);
nand U1805 (N_1805,N_1783,N_1793);
nor U1806 (N_1806,N_1776,N_1789);
xnor U1807 (N_1807,N_1761,N_1755);
nor U1808 (N_1808,N_1798,N_1785);
nand U1809 (N_1809,N_1767,N_1784);
nor U1810 (N_1810,N_1780,N_1762);
and U1811 (N_1811,N_1790,N_1777);
nand U1812 (N_1812,N_1769,N_1763);
xor U1813 (N_1813,N_1765,N_1794);
and U1814 (N_1814,N_1753,N_1750);
or U1815 (N_1815,N_1787,N_1764);
nor U1816 (N_1816,N_1775,N_1766);
nor U1817 (N_1817,N_1759,N_1768);
and U1818 (N_1818,N_1757,N_1782);
or U1819 (N_1819,N_1786,N_1791);
and U1820 (N_1820,N_1771,N_1770);
nor U1821 (N_1821,N_1778,N_1751);
and U1822 (N_1822,N_1756,N_1774);
and U1823 (N_1823,N_1758,N_1792);
and U1824 (N_1824,N_1760,N_1799);
nor U1825 (N_1825,N_1793,N_1796);
nand U1826 (N_1826,N_1773,N_1796);
nand U1827 (N_1827,N_1761,N_1773);
xor U1828 (N_1828,N_1755,N_1781);
nand U1829 (N_1829,N_1795,N_1754);
or U1830 (N_1830,N_1757,N_1766);
nor U1831 (N_1831,N_1763,N_1787);
nor U1832 (N_1832,N_1758,N_1775);
xor U1833 (N_1833,N_1779,N_1767);
xnor U1834 (N_1834,N_1780,N_1769);
or U1835 (N_1835,N_1778,N_1756);
xnor U1836 (N_1836,N_1756,N_1797);
xor U1837 (N_1837,N_1781,N_1770);
nor U1838 (N_1838,N_1770,N_1777);
nand U1839 (N_1839,N_1757,N_1797);
and U1840 (N_1840,N_1781,N_1787);
nor U1841 (N_1841,N_1761,N_1785);
nand U1842 (N_1842,N_1784,N_1770);
or U1843 (N_1843,N_1769,N_1784);
nand U1844 (N_1844,N_1780,N_1783);
xnor U1845 (N_1845,N_1777,N_1793);
xor U1846 (N_1846,N_1789,N_1768);
or U1847 (N_1847,N_1782,N_1775);
nand U1848 (N_1848,N_1799,N_1761);
nor U1849 (N_1849,N_1789,N_1769);
nor U1850 (N_1850,N_1802,N_1848);
nand U1851 (N_1851,N_1847,N_1812);
and U1852 (N_1852,N_1803,N_1825);
nand U1853 (N_1853,N_1819,N_1845);
xor U1854 (N_1854,N_1815,N_1830);
xnor U1855 (N_1855,N_1844,N_1811);
and U1856 (N_1856,N_1846,N_1809);
nor U1857 (N_1857,N_1836,N_1837);
and U1858 (N_1858,N_1835,N_1838);
and U1859 (N_1859,N_1814,N_1818);
or U1860 (N_1860,N_1821,N_1807);
nor U1861 (N_1861,N_1826,N_1831);
and U1862 (N_1862,N_1834,N_1816);
nor U1863 (N_1863,N_1843,N_1840);
nor U1864 (N_1864,N_1833,N_1829);
xor U1865 (N_1865,N_1813,N_1824);
and U1866 (N_1866,N_1817,N_1801);
or U1867 (N_1867,N_1806,N_1805);
nand U1868 (N_1868,N_1820,N_1849);
nor U1869 (N_1869,N_1828,N_1810);
nand U1870 (N_1870,N_1832,N_1842);
and U1871 (N_1871,N_1827,N_1822);
or U1872 (N_1872,N_1800,N_1841);
nor U1873 (N_1873,N_1823,N_1808);
nand U1874 (N_1874,N_1804,N_1839);
or U1875 (N_1875,N_1831,N_1800);
xor U1876 (N_1876,N_1819,N_1802);
and U1877 (N_1877,N_1808,N_1820);
nor U1878 (N_1878,N_1835,N_1822);
nand U1879 (N_1879,N_1844,N_1807);
nor U1880 (N_1880,N_1806,N_1848);
xor U1881 (N_1881,N_1802,N_1800);
and U1882 (N_1882,N_1821,N_1846);
xor U1883 (N_1883,N_1842,N_1841);
or U1884 (N_1884,N_1823,N_1807);
nor U1885 (N_1885,N_1833,N_1806);
nor U1886 (N_1886,N_1846,N_1812);
and U1887 (N_1887,N_1837,N_1823);
and U1888 (N_1888,N_1831,N_1835);
xor U1889 (N_1889,N_1840,N_1822);
and U1890 (N_1890,N_1846,N_1830);
nand U1891 (N_1891,N_1817,N_1825);
nand U1892 (N_1892,N_1838,N_1828);
nand U1893 (N_1893,N_1803,N_1839);
nor U1894 (N_1894,N_1843,N_1832);
nor U1895 (N_1895,N_1824,N_1826);
xor U1896 (N_1896,N_1802,N_1836);
xnor U1897 (N_1897,N_1821,N_1818);
xor U1898 (N_1898,N_1815,N_1820);
nor U1899 (N_1899,N_1847,N_1817);
nand U1900 (N_1900,N_1860,N_1882);
nor U1901 (N_1901,N_1868,N_1855);
nor U1902 (N_1902,N_1870,N_1875);
nand U1903 (N_1903,N_1898,N_1872);
and U1904 (N_1904,N_1881,N_1857);
or U1905 (N_1905,N_1874,N_1864);
and U1906 (N_1906,N_1891,N_1889);
or U1907 (N_1907,N_1893,N_1880);
nor U1908 (N_1908,N_1885,N_1863);
nor U1909 (N_1909,N_1869,N_1852);
xor U1910 (N_1910,N_1887,N_1856);
xnor U1911 (N_1911,N_1861,N_1883);
and U1912 (N_1912,N_1850,N_1899);
and U1913 (N_1913,N_1853,N_1866);
nand U1914 (N_1914,N_1854,N_1896);
xor U1915 (N_1915,N_1858,N_1873);
or U1916 (N_1916,N_1892,N_1884);
xnor U1917 (N_1917,N_1877,N_1876);
xor U1918 (N_1918,N_1865,N_1888);
and U1919 (N_1919,N_1878,N_1859);
or U1920 (N_1920,N_1894,N_1879);
nand U1921 (N_1921,N_1871,N_1862);
nor U1922 (N_1922,N_1895,N_1867);
and U1923 (N_1923,N_1851,N_1886);
nand U1924 (N_1924,N_1897,N_1890);
nand U1925 (N_1925,N_1870,N_1891);
or U1926 (N_1926,N_1889,N_1870);
xnor U1927 (N_1927,N_1887,N_1855);
nor U1928 (N_1928,N_1883,N_1879);
nor U1929 (N_1929,N_1870,N_1881);
or U1930 (N_1930,N_1896,N_1851);
or U1931 (N_1931,N_1862,N_1852);
nor U1932 (N_1932,N_1862,N_1865);
and U1933 (N_1933,N_1858,N_1851);
and U1934 (N_1934,N_1877,N_1866);
and U1935 (N_1935,N_1885,N_1890);
nor U1936 (N_1936,N_1878,N_1851);
xor U1937 (N_1937,N_1879,N_1898);
nand U1938 (N_1938,N_1896,N_1883);
and U1939 (N_1939,N_1860,N_1855);
and U1940 (N_1940,N_1888,N_1882);
or U1941 (N_1941,N_1870,N_1896);
nor U1942 (N_1942,N_1899,N_1865);
nand U1943 (N_1943,N_1879,N_1872);
nand U1944 (N_1944,N_1866,N_1899);
or U1945 (N_1945,N_1868,N_1890);
xnor U1946 (N_1946,N_1889,N_1868);
and U1947 (N_1947,N_1888,N_1871);
nor U1948 (N_1948,N_1883,N_1863);
and U1949 (N_1949,N_1857,N_1886);
and U1950 (N_1950,N_1937,N_1938);
nor U1951 (N_1951,N_1907,N_1909);
nor U1952 (N_1952,N_1942,N_1949);
and U1953 (N_1953,N_1900,N_1916);
xor U1954 (N_1954,N_1933,N_1929);
nand U1955 (N_1955,N_1936,N_1918);
xnor U1956 (N_1956,N_1901,N_1940);
xnor U1957 (N_1957,N_1910,N_1915);
xor U1958 (N_1958,N_1917,N_1931);
nor U1959 (N_1959,N_1920,N_1911);
xor U1960 (N_1960,N_1939,N_1922);
nor U1961 (N_1961,N_1927,N_1923);
nand U1962 (N_1962,N_1903,N_1944);
xor U1963 (N_1963,N_1902,N_1921);
nand U1964 (N_1964,N_1924,N_1919);
and U1965 (N_1965,N_1946,N_1914);
nand U1966 (N_1966,N_1947,N_1913);
nor U1967 (N_1967,N_1943,N_1935);
or U1968 (N_1968,N_1930,N_1905);
xnor U1969 (N_1969,N_1932,N_1925);
nor U1970 (N_1970,N_1928,N_1906);
xor U1971 (N_1971,N_1908,N_1912);
xnor U1972 (N_1972,N_1945,N_1904);
nand U1973 (N_1973,N_1934,N_1941);
nand U1974 (N_1974,N_1948,N_1926);
and U1975 (N_1975,N_1929,N_1909);
nand U1976 (N_1976,N_1943,N_1913);
or U1977 (N_1977,N_1910,N_1933);
nor U1978 (N_1978,N_1943,N_1907);
xnor U1979 (N_1979,N_1917,N_1921);
nor U1980 (N_1980,N_1907,N_1923);
nand U1981 (N_1981,N_1928,N_1924);
and U1982 (N_1982,N_1940,N_1905);
and U1983 (N_1983,N_1908,N_1926);
nor U1984 (N_1984,N_1916,N_1918);
or U1985 (N_1985,N_1906,N_1914);
and U1986 (N_1986,N_1911,N_1924);
nor U1987 (N_1987,N_1949,N_1935);
xnor U1988 (N_1988,N_1901,N_1900);
xor U1989 (N_1989,N_1920,N_1924);
and U1990 (N_1990,N_1949,N_1928);
and U1991 (N_1991,N_1901,N_1921);
nor U1992 (N_1992,N_1926,N_1911);
or U1993 (N_1993,N_1904,N_1920);
and U1994 (N_1994,N_1918,N_1945);
xnor U1995 (N_1995,N_1928,N_1945);
or U1996 (N_1996,N_1949,N_1904);
or U1997 (N_1997,N_1902,N_1943);
and U1998 (N_1998,N_1926,N_1941);
nor U1999 (N_1999,N_1948,N_1904);
or U2000 (N_2000,N_1983,N_1995);
nor U2001 (N_2001,N_1994,N_1953);
or U2002 (N_2002,N_1971,N_1950);
nand U2003 (N_2003,N_1962,N_1960);
xor U2004 (N_2004,N_1968,N_1980);
nand U2005 (N_2005,N_1986,N_1973);
or U2006 (N_2006,N_1982,N_1959);
xnor U2007 (N_2007,N_1963,N_1990);
and U2008 (N_2008,N_1972,N_1979);
xnor U2009 (N_2009,N_1951,N_1952);
xor U2010 (N_2010,N_1985,N_1998);
or U2011 (N_2011,N_1978,N_1974);
or U2012 (N_2012,N_1955,N_1989);
nor U2013 (N_2013,N_1988,N_1964);
or U2014 (N_2014,N_1987,N_1969);
xor U2015 (N_2015,N_1970,N_1993);
nand U2016 (N_2016,N_1965,N_1957);
nand U2017 (N_2017,N_1996,N_1966);
nor U2018 (N_2018,N_1977,N_1992);
or U2019 (N_2019,N_1997,N_1967);
xor U2020 (N_2020,N_1975,N_1999);
nor U2021 (N_2021,N_1958,N_1984);
and U2022 (N_2022,N_1961,N_1991);
or U2023 (N_2023,N_1976,N_1981);
or U2024 (N_2024,N_1956,N_1954);
nand U2025 (N_2025,N_1995,N_1988);
and U2026 (N_2026,N_1961,N_1970);
xor U2027 (N_2027,N_1962,N_1982);
nand U2028 (N_2028,N_1972,N_1997);
xor U2029 (N_2029,N_1988,N_1982);
nand U2030 (N_2030,N_1991,N_1985);
and U2031 (N_2031,N_1970,N_1977);
and U2032 (N_2032,N_1970,N_1956);
nand U2033 (N_2033,N_1968,N_1988);
and U2034 (N_2034,N_1997,N_1988);
or U2035 (N_2035,N_1977,N_1971);
or U2036 (N_2036,N_1993,N_1989);
xor U2037 (N_2037,N_1969,N_1968);
or U2038 (N_2038,N_1990,N_1967);
and U2039 (N_2039,N_1980,N_1969);
and U2040 (N_2040,N_1992,N_1961);
xor U2041 (N_2041,N_1966,N_1989);
xnor U2042 (N_2042,N_1982,N_1996);
or U2043 (N_2043,N_1982,N_1998);
and U2044 (N_2044,N_1977,N_1982);
or U2045 (N_2045,N_1978,N_1981);
nor U2046 (N_2046,N_1958,N_1964);
nor U2047 (N_2047,N_1985,N_1951);
and U2048 (N_2048,N_1989,N_1975);
nand U2049 (N_2049,N_1961,N_1975);
nor U2050 (N_2050,N_2046,N_2017);
nor U2051 (N_2051,N_2005,N_2028);
nor U2052 (N_2052,N_2006,N_2007);
and U2053 (N_2053,N_2030,N_2019);
nor U2054 (N_2054,N_2043,N_2048);
or U2055 (N_2055,N_2039,N_2036);
and U2056 (N_2056,N_2021,N_2022);
xnor U2057 (N_2057,N_2037,N_2008);
nor U2058 (N_2058,N_2000,N_2047);
or U2059 (N_2059,N_2027,N_2034);
and U2060 (N_2060,N_2044,N_2020);
or U2061 (N_2061,N_2029,N_2023);
xnor U2062 (N_2062,N_2031,N_2016);
or U2063 (N_2063,N_2038,N_2015);
and U2064 (N_2064,N_2014,N_2024);
nor U2065 (N_2065,N_2041,N_2003);
and U2066 (N_2066,N_2045,N_2025);
xnor U2067 (N_2067,N_2032,N_2009);
nand U2068 (N_2068,N_2018,N_2049);
nand U2069 (N_2069,N_2040,N_2010);
nand U2070 (N_2070,N_2013,N_2012);
and U2071 (N_2071,N_2026,N_2002);
or U2072 (N_2072,N_2011,N_2042);
and U2073 (N_2073,N_2033,N_2004);
or U2074 (N_2074,N_2035,N_2001);
or U2075 (N_2075,N_2003,N_2040);
or U2076 (N_2076,N_2005,N_2037);
and U2077 (N_2077,N_2007,N_2031);
xnor U2078 (N_2078,N_2028,N_2018);
nand U2079 (N_2079,N_2014,N_2004);
nand U2080 (N_2080,N_2030,N_2008);
and U2081 (N_2081,N_2014,N_2031);
nor U2082 (N_2082,N_2032,N_2039);
xor U2083 (N_2083,N_2022,N_2025);
nor U2084 (N_2084,N_2036,N_2046);
nand U2085 (N_2085,N_2031,N_2026);
and U2086 (N_2086,N_2004,N_2035);
or U2087 (N_2087,N_2009,N_2002);
or U2088 (N_2088,N_2016,N_2044);
and U2089 (N_2089,N_2008,N_2025);
nand U2090 (N_2090,N_2040,N_2021);
xor U2091 (N_2091,N_2034,N_2040);
or U2092 (N_2092,N_2020,N_2034);
or U2093 (N_2093,N_2025,N_2019);
nand U2094 (N_2094,N_2034,N_2013);
nor U2095 (N_2095,N_2004,N_2037);
xnor U2096 (N_2096,N_2022,N_2020);
and U2097 (N_2097,N_2004,N_2018);
and U2098 (N_2098,N_2000,N_2021);
nor U2099 (N_2099,N_2026,N_2007);
nand U2100 (N_2100,N_2070,N_2060);
xnor U2101 (N_2101,N_2085,N_2093);
or U2102 (N_2102,N_2065,N_2069);
nand U2103 (N_2103,N_2088,N_2059);
nand U2104 (N_2104,N_2052,N_2066);
and U2105 (N_2105,N_2097,N_2051);
or U2106 (N_2106,N_2099,N_2078);
or U2107 (N_2107,N_2076,N_2086);
xnor U2108 (N_2108,N_2072,N_2084);
nor U2109 (N_2109,N_2071,N_2055);
nand U2110 (N_2110,N_2080,N_2098);
or U2111 (N_2111,N_2091,N_2082);
and U2112 (N_2112,N_2087,N_2062);
nor U2113 (N_2113,N_2057,N_2079);
or U2114 (N_2114,N_2050,N_2095);
nor U2115 (N_2115,N_2056,N_2083);
nand U2116 (N_2116,N_2090,N_2089);
xor U2117 (N_2117,N_2077,N_2094);
nand U2118 (N_2118,N_2067,N_2075);
nor U2119 (N_2119,N_2058,N_2053);
nand U2120 (N_2120,N_2073,N_2081);
xnor U2121 (N_2121,N_2064,N_2092);
nand U2122 (N_2122,N_2054,N_2096);
and U2123 (N_2123,N_2061,N_2074);
or U2124 (N_2124,N_2063,N_2068);
or U2125 (N_2125,N_2077,N_2082);
nand U2126 (N_2126,N_2053,N_2097);
and U2127 (N_2127,N_2092,N_2089);
nand U2128 (N_2128,N_2095,N_2082);
nor U2129 (N_2129,N_2092,N_2065);
or U2130 (N_2130,N_2066,N_2054);
nand U2131 (N_2131,N_2086,N_2056);
nand U2132 (N_2132,N_2063,N_2094);
nor U2133 (N_2133,N_2051,N_2085);
xnor U2134 (N_2134,N_2087,N_2085);
nor U2135 (N_2135,N_2090,N_2069);
and U2136 (N_2136,N_2079,N_2073);
or U2137 (N_2137,N_2056,N_2087);
xor U2138 (N_2138,N_2060,N_2059);
and U2139 (N_2139,N_2096,N_2066);
and U2140 (N_2140,N_2089,N_2063);
and U2141 (N_2141,N_2052,N_2074);
and U2142 (N_2142,N_2090,N_2085);
and U2143 (N_2143,N_2089,N_2083);
nand U2144 (N_2144,N_2077,N_2060);
and U2145 (N_2145,N_2066,N_2059);
nand U2146 (N_2146,N_2096,N_2082);
nor U2147 (N_2147,N_2067,N_2099);
or U2148 (N_2148,N_2090,N_2094);
nor U2149 (N_2149,N_2077,N_2084);
or U2150 (N_2150,N_2148,N_2143);
or U2151 (N_2151,N_2128,N_2142);
nor U2152 (N_2152,N_2133,N_2116);
or U2153 (N_2153,N_2114,N_2130);
or U2154 (N_2154,N_2101,N_2119);
nor U2155 (N_2155,N_2108,N_2132);
xor U2156 (N_2156,N_2127,N_2104);
nand U2157 (N_2157,N_2144,N_2139);
xnor U2158 (N_2158,N_2124,N_2120);
nand U2159 (N_2159,N_2134,N_2110);
xnor U2160 (N_2160,N_2105,N_2121);
and U2161 (N_2161,N_2125,N_2111);
and U2162 (N_2162,N_2103,N_2149);
xnor U2163 (N_2163,N_2109,N_2126);
xor U2164 (N_2164,N_2122,N_2100);
and U2165 (N_2165,N_2141,N_2115);
nor U2166 (N_2166,N_2107,N_2145);
nor U2167 (N_2167,N_2112,N_2131);
nand U2168 (N_2168,N_2147,N_2136);
xnor U2169 (N_2169,N_2129,N_2118);
nand U2170 (N_2170,N_2137,N_2106);
xnor U2171 (N_2171,N_2123,N_2113);
nor U2172 (N_2172,N_2102,N_2146);
xnor U2173 (N_2173,N_2138,N_2117);
xor U2174 (N_2174,N_2135,N_2140);
nand U2175 (N_2175,N_2139,N_2133);
xnor U2176 (N_2176,N_2140,N_2108);
nand U2177 (N_2177,N_2110,N_2125);
or U2178 (N_2178,N_2149,N_2126);
xnor U2179 (N_2179,N_2116,N_2104);
nand U2180 (N_2180,N_2128,N_2109);
nand U2181 (N_2181,N_2147,N_2118);
nor U2182 (N_2182,N_2129,N_2145);
nand U2183 (N_2183,N_2109,N_2103);
and U2184 (N_2184,N_2145,N_2110);
xnor U2185 (N_2185,N_2106,N_2141);
and U2186 (N_2186,N_2140,N_2145);
or U2187 (N_2187,N_2117,N_2107);
or U2188 (N_2188,N_2134,N_2112);
nor U2189 (N_2189,N_2104,N_2113);
nor U2190 (N_2190,N_2147,N_2131);
xor U2191 (N_2191,N_2103,N_2145);
nand U2192 (N_2192,N_2137,N_2134);
nor U2193 (N_2193,N_2119,N_2114);
and U2194 (N_2194,N_2119,N_2148);
and U2195 (N_2195,N_2125,N_2142);
nand U2196 (N_2196,N_2138,N_2113);
nand U2197 (N_2197,N_2125,N_2118);
nor U2198 (N_2198,N_2101,N_2122);
or U2199 (N_2199,N_2139,N_2127);
and U2200 (N_2200,N_2164,N_2150);
xnor U2201 (N_2201,N_2156,N_2166);
nand U2202 (N_2202,N_2183,N_2165);
nor U2203 (N_2203,N_2161,N_2154);
or U2204 (N_2204,N_2163,N_2174);
xnor U2205 (N_2205,N_2179,N_2186);
xor U2206 (N_2206,N_2170,N_2178);
nor U2207 (N_2207,N_2182,N_2160);
or U2208 (N_2208,N_2195,N_2152);
nor U2209 (N_2209,N_2162,N_2190);
and U2210 (N_2210,N_2159,N_2151);
xor U2211 (N_2211,N_2175,N_2197);
nand U2212 (N_2212,N_2196,N_2167);
nor U2213 (N_2213,N_2184,N_2193);
or U2214 (N_2214,N_2158,N_2192);
and U2215 (N_2215,N_2189,N_2157);
and U2216 (N_2216,N_2187,N_2199);
nor U2217 (N_2217,N_2194,N_2185);
nor U2218 (N_2218,N_2198,N_2172);
and U2219 (N_2219,N_2191,N_2177);
and U2220 (N_2220,N_2188,N_2171);
and U2221 (N_2221,N_2168,N_2173);
nand U2222 (N_2222,N_2169,N_2176);
nand U2223 (N_2223,N_2181,N_2155);
xor U2224 (N_2224,N_2180,N_2153);
xor U2225 (N_2225,N_2185,N_2157);
and U2226 (N_2226,N_2193,N_2186);
and U2227 (N_2227,N_2191,N_2167);
and U2228 (N_2228,N_2158,N_2178);
xor U2229 (N_2229,N_2166,N_2178);
xnor U2230 (N_2230,N_2175,N_2156);
and U2231 (N_2231,N_2172,N_2161);
nand U2232 (N_2232,N_2176,N_2192);
nor U2233 (N_2233,N_2180,N_2176);
xnor U2234 (N_2234,N_2185,N_2189);
nand U2235 (N_2235,N_2167,N_2157);
or U2236 (N_2236,N_2175,N_2168);
or U2237 (N_2237,N_2191,N_2183);
and U2238 (N_2238,N_2155,N_2176);
xnor U2239 (N_2239,N_2166,N_2155);
nor U2240 (N_2240,N_2175,N_2190);
or U2241 (N_2241,N_2193,N_2160);
nand U2242 (N_2242,N_2181,N_2191);
or U2243 (N_2243,N_2194,N_2177);
and U2244 (N_2244,N_2155,N_2189);
and U2245 (N_2245,N_2156,N_2196);
nand U2246 (N_2246,N_2185,N_2154);
and U2247 (N_2247,N_2160,N_2166);
xor U2248 (N_2248,N_2189,N_2152);
nand U2249 (N_2249,N_2194,N_2173);
or U2250 (N_2250,N_2214,N_2224);
nor U2251 (N_2251,N_2228,N_2201);
and U2252 (N_2252,N_2238,N_2249);
or U2253 (N_2253,N_2204,N_2213);
nor U2254 (N_2254,N_2229,N_2232);
xnor U2255 (N_2255,N_2217,N_2209);
and U2256 (N_2256,N_2241,N_2244);
nand U2257 (N_2257,N_2211,N_2235);
nor U2258 (N_2258,N_2220,N_2223);
xor U2259 (N_2259,N_2243,N_2215);
and U2260 (N_2260,N_2221,N_2242);
nand U2261 (N_2261,N_2231,N_2212);
nor U2262 (N_2262,N_2225,N_2240);
nor U2263 (N_2263,N_2230,N_2216);
or U2264 (N_2264,N_2208,N_2233);
or U2265 (N_2265,N_2227,N_2202);
and U2266 (N_2266,N_2200,N_2210);
nor U2267 (N_2267,N_2248,N_2234);
nand U2268 (N_2268,N_2218,N_2222);
and U2269 (N_2269,N_2219,N_2247);
or U2270 (N_2270,N_2237,N_2246);
xnor U2271 (N_2271,N_2203,N_2205);
or U2272 (N_2272,N_2226,N_2206);
nand U2273 (N_2273,N_2207,N_2245);
nand U2274 (N_2274,N_2236,N_2239);
nand U2275 (N_2275,N_2207,N_2219);
nor U2276 (N_2276,N_2230,N_2211);
xor U2277 (N_2277,N_2222,N_2215);
nand U2278 (N_2278,N_2244,N_2223);
xor U2279 (N_2279,N_2234,N_2228);
nand U2280 (N_2280,N_2241,N_2238);
xnor U2281 (N_2281,N_2219,N_2242);
nor U2282 (N_2282,N_2247,N_2202);
or U2283 (N_2283,N_2224,N_2230);
xor U2284 (N_2284,N_2231,N_2208);
nand U2285 (N_2285,N_2218,N_2204);
xnor U2286 (N_2286,N_2209,N_2227);
xor U2287 (N_2287,N_2221,N_2227);
nor U2288 (N_2288,N_2240,N_2227);
and U2289 (N_2289,N_2243,N_2235);
xnor U2290 (N_2290,N_2216,N_2214);
nor U2291 (N_2291,N_2206,N_2207);
xor U2292 (N_2292,N_2231,N_2221);
xnor U2293 (N_2293,N_2248,N_2215);
and U2294 (N_2294,N_2234,N_2227);
xnor U2295 (N_2295,N_2202,N_2237);
xnor U2296 (N_2296,N_2243,N_2227);
nand U2297 (N_2297,N_2234,N_2246);
nand U2298 (N_2298,N_2247,N_2242);
xor U2299 (N_2299,N_2213,N_2216);
nand U2300 (N_2300,N_2285,N_2274);
and U2301 (N_2301,N_2288,N_2277);
xnor U2302 (N_2302,N_2276,N_2287);
nand U2303 (N_2303,N_2271,N_2273);
nor U2304 (N_2304,N_2257,N_2295);
nand U2305 (N_2305,N_2250,N_2296);
xnor U2306 (N_2306,N_2272,N_2262);
and U2307 (N_2307,N_2289,N_2292);
and U2308 (N_2308,N_2297,N_2251);
xnor U2309 (N_2309,N_2290,N_2256);
nor U2310 (N_2310,N_2252,N_2260);
nand U2311 (N_2311,N_2284,N_2255);
xnor U2312 (N_2312,N_2279,N_2294);
and U2313 (N_2313,N_2298,N_2278);
nand U2314 (N_2314,N_2291,N_2299);
nand U2315 (N_2315,N_2282,N_2264);
nand U2316 (N_2316,N_2265,N_2266);
xor U2317 (N_2317,N_2261,N_2268);
or U2318 (N_2318,N_2280,N_2281);
nor U2319 (N_2319,N_2259,N_2253);
nor U2320 (N_2320,N_2293,N_2254);
xnor U2321 (N_2321,N_2267,N_2275);
nand U2322 (N_2322,N_2286,N_2283);
xor U2323 (N_2323,N_2263,N_2270);
xnor U2324 (N_2324,N_2258,N_2269);
or U2325 (N_2325,N_2299,N_2269);
nand U2326 (N_2326,N_2279,N_2259);
and U2327 (N_2327,N_2264,N_2267);
nand U2328 (N_2328,N_2274,N_2287);
or U2329 (N_2329,N_2293,N_2269);
nor U2330 (N_2330,N_2294,N_2258);
and U2331 (N_2331,N_2277,N_2287);
nand U2332 (N_2332,N_2270,N_2287);
xor U2333 (N_2333,N_2252,N_2294);
nand U2334 (N_2334,N_2280,N_2283);
xnor U2335 (N_2335,N_2262,N_2288);
or U2336 (N_2336,N_2268,N_2255);
xor U2337 (N_2337,N_2299,N_2283);
nor U2338 (N_2338,N_2298,N_2251);
xor U2339 (N_2339,N_2250,N_2265);
nor U2340 (N_2340,N_2286,N_2280);
nand U2341 (N_2341,N_2297,N_2262);
xnor U2342 (N_2342,N_2286,N_2279);
xnor U2343 (N_2343,N_2250,N_2299);
nand U2344 (N_2344,N_2255,N_2262);
and U2345 (N_2345,N_2275,N_2283);
xnor U2346 (N_2346,N_2259,N_2262);
xnor U2347 (N_2347,N_2270,N_2294);
xor U2348 (N_2348,N_2253,N_2267);
or U2349 (N_2349,N_2275,N_2287);
nand U2350 (N_2350,N_2330,N_2310);
and U2351 (N_2351,N_2338,N_2305);
nor U2352 (N_2352,N_2332,N_2304);
nand U2353 (N_2353,N_2336,N_2312);
nand U2354 (N_2354,N_2328,N_2323);
or U2355 (N_2355,N_2315,N_2318);
xor U2356 (N_2356,N_2339,N_2344);
nand U2357 (N_2357,N_2329,N_2324);
nor U2358 (N_2358,N_2349,N_2314);
xor U2359 (N_2359,N_2317,N_2337);
and U2360 (N_2360,N_2331,N_2308);
nand U2361 (N_2361,N_2301,N_2333);
nor U2362 (N_2362,N_2313,N_2326);
nor U2363 (N_2363,N_2345,N_2322);
or U2364 (N_2364,N_2335,N_2307);
or U2365 (N_2365,N_2300,N_2302);
xor U2366 (N_2366,N_2341,N_2325);
xnor U2367 (N_2367,N_2320,N_2306);
xnor U2368 (N_2368,N_2311,N_2316);
or U2369 (N_2369,N_2348,N_2343);
xor U2370 (N_2370,N_2321,N_2319);
or U2371 (N_2371,N_2327,N_2347);
nor U2372 (N_2372,N_2309,N_2342);
or U2373 (N_2373,N_2334,N_2340);
or U2374 (N_2374,N_2303,N_2346);
nand U2375 (N_2375,N_2324,N_2305);
nand U2376 (N_2376,N_2306,N_2329);
nand U2377 (N_2377,N_2341,N_2339);
nand U2378 (N_2378,N_2346,N_2325);
or U2379 (N_2379,N_2303,N_2344);
or U2380 (N_2380,N_2324,N_2328);
xor U2381 (N_2381,N_2320,N_2301);
nor U2382 (N_2382,N_2326,N_2310);
xnor U2383 (N_2383,N_2345,N_2349);
and U2384 (N_2384,N_2303,N_2332);
and U2385 (N_2385,N_2330,N_2341);
nand U2386 (N_2386,N_2318,N_2341);
xor U2387 (N_2387,N_2339,N_2334);
xnor U2388 (N_2388,N_2346,N_2328);
nor U2389 (N_2389,N_2309,N_2330);
nor U2390 (N_2390,N_2346,N_2318);
nand U2391 (N_2391,N_2324,N_2321);
nor U2392 (N_2392,N_2316,N_2330);
xnor U2393 (N_2393,N_2330,N_2304);
nor U2394 (N_2394,N_2349,N_2324);
nand U2395 (N_2395,N_2345,N_2307);
nand U2396 (N_2396,N_2309,N_2340);
nand U2397 (N_2397,N_2347,N_2301);
and U2398 (N_2398,N_2310,N_2343);
and U2399 (N_2399,N_2305,N_2306);
or U2400 (N_2400,N_2361,N_2351);
nor U2401 (N_2401,N_2394,N_2354);
nor U2402 (N_2402,N_2362,N_2367);
or U2403 (N_2403,N_2377,N_2396);
and U2404 (N_2404,N_2358,N_2357);
nand U2405 (N_2405,N_2382,N_2365);
or U2406 (N_2406,N_2387,N_2381);
or U2407 (N_2407,N_2393,N_2360);
xnor U2408 (N_2408,N_2388,N_2373);
xor U2409 (N_2409,N_2371,N_2390);
or U2410 (N_2410,N_2375,N_2398);
xnor U2411 (N_2411,N_2395,N_2376);
and U2412 (N_2412,N_2386,N_2366);
or U2413 (N_2413,N_2378,N_2359);
and U2414 (N_2414,N_2391,N_2392);
or U2415 (N_2415,N_2353,N_2380);
and U2416 (N_2416,N_2397,N_2364);
nor U2417 (N_2417,N_2350,N_2379);
nand U2418 (N_2418,N_2372,N_2356);
or U2419 (N_2419,N_2369,N_2385);
nand U2420 (N_2420,N_2384,N_2383);
nand U2421 (N_2421,N_2352,N_2399);
xnor U2422 (N_2422,N_2368,N_2374);
nand U2423 (N_2423,N_2363,N_2355);
or U2424 (N_2424,N_2370,N_2389);
and U2425 (N_2425,N_2396,N_2398);
nand U2426 (N_2426,N_2387,N_2379);
nor U2427 (N_2427,N_2369,N_2375);
nor U2428 (N_2428,N_2368,N_2379);
nor U2429 (N_2429,N_2390,N_2373);
or U2430 (N_2430,N_2380,N_2354);
nor U2431 (N_2431,N_2377,N_2356);
xnor U2432 (N_2432,N_2377,N_2395);
xor U2433 (N_2433,N_2380,N_2367);
or U2434 (N_2434,N_2386,N_2361);
nor U2435 (N_2435,N_2368,N_2367);
nand U2436 (N_2436,N_2389,N_2359);
or U2437 (N_2437,N_2387,N_2364);
nor U2438 (N_2438,N_2361,N_2360);
and U2439 (N_2439,N_2396,N_2378);
or U2440 (N_2440,N_2395,N_2386);
or U2441 (N_2441,N_2389,N_2367);
or U2442 (N_2442,N_2399,N_2388);
or U2443 (N_2443,N_2370,N_2379);
nand U2444 (N_2444,N_2386,N_2397);
or U2445 (N_2445,N_2359,N_2373);
or U2446 (N_2446,N_2396,N_2397);
nor U2447 (N_2447,N_2392,N_2380);
and U2448 (N_2448,N_2363,N_2375);
xnor U2449 (N_2449,N_2355,N_2370);
nor U2450 (N_2450,N_2436,N_2416);
and U2451 (N_2451,N_2446,N_2412);
and U2452 (N_2452,N_2415,N_2422);
xnor U2453 (N_2453,N_2437,N_2411);
nand U2454 (N_2454,N_2431,N_2403);
xnor U2455 (N_2455,N_2413,N_2410);
xor U2456 (N_2456,N_2426,N_2448);
nor U2457 (N_2457,N_2438,N_2409);
xor U2458 (N_2458,N_2420,N_2414);
or U2459 (N_2459,N_2435,N_2424);
xor U2460 (N_2460,N_2443,N_2427);
and U2461 (N_2461,N_2406,N_2421);
or U2462 (N_2462,N_2405,N_2407);
nand U2463 (N_2463,N_2428,N_2401);
or U2464 (N_2464,N_2434,N_2444);
or U2465 (N_2465,N_2449,N_2418);
or U2466 (N_2466,N_2423,N_2408);
or U2467 (N_2467,N_2417,N_2447);
and U2468 (N_2468,N_2445,N_2430);
xnor U2469 (N_2469,N_2432,N_2400);
nor U2470 (N_2470,N_2419,N_2439);
nor U2471 (N_2471,N_2429,N_2441);
xnor U2472 (N_2472,N_2402,N_2404);
nor U2473 (N_2473,N_2433,N_2442);
and U2474 (N_2474,N_2425,N_2440);
nand U2475 (N_2475,N_2436,N_2408);
xnor U2476 (N_2476,N_2444,N_2433);
nand U2477 (N_2477,N_2440,N_2424);
or U2478 (N_2478,N_2448,N_2432);
nand U2479 (N_2479,N_2421,N_2400);
nand U2480 (N_2480,N_2410,N_2406);
xor U2481 (N_2481,N_2427,N_2422);
nor U2482 (N_2482,N_2440,N_2444);
nand U2483 (N_2483,N_2433,N_2421);
xnor U2484 (N_2484,N_2429,N_2444);
and U2485 (N_2485,N_2414,N_2421);
or U2486 (N_2486,N_2402,N_2442);
xnor U2487 (N_2487,N_2441,N_2438);
nand U2488 (N_2488,N_2418,N_2435);
nor U2489 (N_2489,N_2409,N_2416);
xnor U2490 (N_2490,N_2443,N_2440);
xor U2491 (N_2491,N_2406,N_2438);
nor U2492 (N_2492,N_2426,N_2414);
nand U2493 (N_2493,N_2430,N_2437);
nand U2494 (N_2494,N_2404,N_2415);
or U2495 (N_2495,N_2402,N_2400);
or U2496 (N_2496,N_2439,N_2440);
or U2497 (N_2497,N_2435,N_2406);
or U2498 (N_2498,N_2408,N_2407);
xor U2499 (N_2499,N_2445,N_2416);
xor U2500 (N_2500,N_2497,N_2469);
xnor U2501 (N_2501,N_2482,N_2489);
nand U2502 (N_2502,N_2483,N_2492);
xor U2503 (N_2503,N_2466,N_2450);
xnor U2504 (N_2504,N_2473,N_2464);
nor U2505 (N_2505,N_2487,N_2475);
nand U2506 (N_2506,N_2472,N_2476);
nand U2507 (N_2507,N_2486,N_2499);
and U2508 (N_2508,N_2491,N_2452);
and U2509 (N_2509,N_2481,N_2456);
xor U2510 (N_2510,N_2453,N_2495);
and U2511 (N_2511,N_2474,N_2477);
nor U2512 (N_2512,N_2463,N_2455);
nor U2513 (N_2513,N_2478,N_2493);
nor U2514 (N_2514,N_2494,N_2451);
and U2515 (N_2515,N_2488,N_2458);
nor U2516 (N_2516,N_2459,N_2498);
or U2517 (N_2517,N_2465,N_2485);
xnor U2518 (N_2518,N_2490,N_2468);
or U2519 (N_2519,N_2471,N_2467);
or U2520 (N_2520,N_2462,N_2480);
and U2521 (N_2521,N_2479,N_2457);
xnor U2522 (N_2522,N_2470,N_2484);
and U2523 (N_2523,N_2460,N_2454);
and U2524 (N_2524,N_2496,N_2461);
nand U2525 (N_2525,N_2499,N_2469);
nor U2526 (N_2526,N_2499,N_2479);
or U2527 (N_2527,N_2490,N_2458);
and U2528 (N_2528,N_2477,N_2479);
and U2529 (N_2529,N_2487,N_2495);
and U2530 (N_2530,N_2492,N_2474);
and U2531 (N_2531,N_2462,N_2496);
xor U2532 (N_2532,N_2495,N_2481);
nand U2533 (N_2533,N_2480,N_2488);
and U2534 (N_2534,N_2499,N_2460);
and U2535 (N_2535,N_2480,N_2457);
nand U2536 (N_2536,N_2498,N_2455);
or U2537 (N_2537,N_2489,N_2467);
nor U2538 (N_2538,N_2472,N_2450);
and U2539 (N_2539,N_2493,N_2469);
nand U2540 (N_2540,N_2488,N_2482);
xnor U2541 (N_2541,N_2493,N_2486);
nand U2542 (N_2542,N_2457,N_2488);
nand U2543 (N_2543,N_2459,N_2473);
nand U2544 (N_2544,N_2452,N_2472);
or U2545 (N_2545,N_2497,N_2481);
nor U2546 (N_2546,N_2469,N_2464);
xor U2547 (N_2547,N_2464,N_2458);
nand U2548 (N_2548,N_2490,N_2485);
xnor U2549 (N_2549,N_2452,N_2479);
and U2550 (N_2550,N_2507,N_2540);
and U2551 (N_2551,N_2515,N_2545);
nor U2552 (N_2552,N_2509,N_2529);
and U2553 (N_2553,N_2544,N_2519);
xor U2554 (N_2554,N_2524,N_2542);
nand U2555 (N_2555,N_2503,N_2504);
xor U2556 (N_2556,N_2537,N_2508);
or U2557 (N_2557,N_2500,N_2527);
and U2558 (N_2558,N_2547,N_2511);
nor U2559 (N_2559,N_2536,N_2546);
or U2560 (N_2560,N_2530,N_2506);
nand U2561 (N_2561,N_2505,N_2518);
nand U2562 (N_2562,N_2521,N_2531);
xnor U2563 (N_2563,N_2514,N_2516);
xnor U2564 (N_2564,N_2532,N_2538);
nand U2565 (N_2565,N_2510,N_2543);
xnor U2566 (N_2566,N_2522,N_2501);
or U2567 (N_2567,N_2523,N_2520);
nand U2568 (N_2568,N_2502,N_2533);
xor U2569 (N_2569,N_2549,N_2528);
nand U2570 (N_2570,N_2534,N_2525);
xnor U2571 (N_2571,N_2517,N_2548);
nand U2572 (N_2572,N_2526,N_2541);
and U2573 (N_2573,N_2535,N_2513);
nor U2574 (N_2574,N_2539,N_2512);
nor U2575 (N_2575,N_2523,N_2519);
and U2576 (N_2576,N_2544,N_2502);
xor U2577 (N_2577,N_2503,N_2533);
nand U2578 (N_2578,N_2518,N_2526);
or U2579 (N_2579,N_2544,N_2503);
and U2580 (N_2580,N_2532,N_2506);
xnor U2581 (N_2581,N_2515,N_2505);
nor U2582 (N_2582,N_2518,N_2537);
and U2583 (N_2583,N_2539,N_2507);
nor U2584 (N_2584,N_2529,N_2504);
or U2585 (N_2585,N_2514,N_2507);
nand U2586 (N_2586,N_2539,N_2528);
nand U2587 (N_2587,N_2530,N_2501);
xnor U2588 (N_2588,N_2528,N_2529);
or U2589 (N_2589,N_2522,N_2527);
nand U2590 (N_2590,N_2510,N_2537);
nand U2591 (N_2591,N_2516,N_2529);
nand U2592 (N_2592,N_2500,N_2533);
or U2593 (N_2593,N_2549,N_2508);
nand U2594 (N_2594,N_2513,N_2522);
or U2595 (N_2595,N_2543,N_2545);
nor U2596 (N_2596,N_2512,N_2546);
nor U2597 (N_2597,N_2527,N_2545);
nand U2598 (N_2598,N_2549,N_2520);
and U2599 (N_2599,N_2515,N_2540);
or U2600 (N_2600,N_2571,N_2590);
and U2601 (N_2601,N_2596,N_2570);
nor U2602 (N_2602,N_2552,N_2586);
and U2603 (N_2603,N_2577,N_2576);
or U2604 (N_2604,N_2563,N_2566);
and U2605 (N_2605,N_2568,N_2579);
nand U2606 (N_2606,N_2580,N_2591);
and U2607 (N_2607,N_2578,N_2555);
xnor U2608 (N_2608,N_2550,N_2594);
and U2609 (N_2609,N_2588,N_2593);
xor U2610 (N_2610,N_2574,N_2598);
xnor U2611 (N_2611,N_2584,N_2573);
nand U2612 (N_2612,N_2560,N_2583);
xnor U2613 (N_2613,N_2561,N_2582);
and U2614 (N_2614,N_2572,N_2558);
nor U2615 (N_2615,N_2587,N_2559);
nor U2616 (N_2616,N_2581,N_2589);
or U2617 (N_2617,N_2597,N_2595);
or U2618 (N_2618,N_2569,N_2564);
and U2619 (N_2619,N_2556,N_2557);
or U2620 (N_2620,N_2554,N_2592);
xor U2621 (N_2621,N_2551,N_2565);
and U2622 (N_2622,N_2599,N_2553);
nand U2623 (N_2623,N_2585,N_2567);
or U2624 (N_2624,N_2575,N_2562);
nor U2625 (N_2625,N_2599,N_2570);
or U2626 (N_2626,N_2593,N_2562);
nor U2627 (N_2627,N_2574,N_2578);
and U2628 (N_2628,N_2554,N_2556);
nor U2629 (N_2629,N_2562,N_2586);
nand U2630 (N_2630,N_2554,N_2595);
xor U2631 (N_2631,N_2554,N_2564);
nor U2632 (N_2632,N_2558,N_2551);
nand U2633 (N_2633,N_2599,N_2561);
nand U2634 (N_2634,N_2552,N_2581);
xor U2635 (N_2635,N_2558,N_2555);
xor U2636 (N_2636,N_2588,N_2582);
xnor U2637 (N_2637,N_2558,N_2563);
or U2638 (N_2638,N_2578,N_2586);
xnor U2639 (N_2639,N_2587,N_2597);
and U2640 (N_2640,N_2561,N_2596);
xnor U2641 (N_2641,N_2564,N_2558);
or U2642 (N_2642,N_2573,N_2572);
nor U2643 (N_2643,N_2583,N_2593);
nor U2644 (N_2644,N_2551,N_2587);
and U2645 (N_2645,N_2595,N_2590);
xnor U2646 (N_2646,N_2560,N_2572);
and U2647 (N_2647,N_2556,N_2586);
or U2648 (N_2648,N_2553,N_2597);
xor U2649 (N_2649,N_2565,N_2552);
nor U2650 (N_2650,N_2641,N_2628);
and U2651 (N_2651,N_2636,N_2633);
and U2652 (N_2652,N_2621,N_2623);
and U2653 (N_2653,N_2645,N_2606);
nor U2654 (N_2654,N_2613,N_2646);
xnor U2655 (N_2655,N_2637,N_2630);
and U2656 (N_2656,N_2639,N_2635);
and U2657 (N_2657,N_2649,N_2625);
and U2658 (N_2658,N_2608,N_2647);
and U2659 (N_2659,N_2642,N_2607);
xnor U2660 (N_2660,N_2627,N_2610);
or U2661 (N_2661,N_2620,N_2609);
nor U2662 (N_2662,N_2632,N_2604);
nor U2663 (N_2663,N_2634,N_2648);
and U2664 (N_2664,N_2612,N_2619);
or U2665 (N_2665,N_2643,N_2616);
or U2666 (N_2666,N_2631,N_2603);
nor U2667 (N_2667,N_2601,N_2611);
nand U2668 (N_2668,N_2622,N_2615);
nor U2669 (N_2669,N_2638,N_2644);
or U2670 (N_2670,N_2614,N_2618);
nand U2671 (N_2671,N_2640,N_2602);
nand U2672 (N_2672,N_2605,N_2617);
xor U2673 (N_2673,N_2626,N_2624);
nand U2674 (N_2674,N_2629,N_2600);
and U2675 (N_2675,N_2605,N_2615);
and U2676 (N_2676,N_2618,N_2629);
and U2677 (N_2677,N_2637,N_2612);
or U2678 (N_2678,N_2626,N_2611);
or U2679 (N_2679,N_2603,N_2609);
nand U2680 (N_2680,N_2648,N_2625);
and U2681 (N_2681,N_2638,N_2620);
xor U2682 (N_2682,N_2645,N_2634);
or U2683 (N_2683,N_2625,N_2618);
xnor U2684 (N_2684,N_2610,N_2600);
or U2685 (N_2685,N_2605,N_2640);
nor U2686 (N_2686,N_2629,N_2604);
nand U2687 (N_2687,N_2644,N_2613);
nand U2688 (N_2688,N_2606,N_2625);
xnor U2689 (N_2689,N_2603,N_2604);
or U2690 (N_2690,N_2622,N_2636);
or U2691 (N_2691,N_2601,N_2647);
and U2692 (N_2692,N_2613,N_2630);
nand U2693 (N_2693,N_2602,N_2636);
nand U2694 (N_2694,N_2602,N_2609);
or U2695 (N_2695,N_2622,N_2614);
xnor U2696 (N_2696,N_2622,N_2612);
nor U2697 (N_2697,N_2619,N_2630);
or U2698 (N_2698,N_2616,N_2621);
xor U2699 (N_2699,N_2628,N_2635);
nand U2700 (N_2700,N_2699,N_2654);
nor U2701 (N_2701,N_2695,N_2679);
nor U2702 (N_2702,N_2668,N_2698);
nand U2703 (N_2703,N_2669,N_2681);
xnor U2704 (N_2704,N_2650,N_2653);
xor U2705 (N_2705,N_2666,N_2680);
nand U2706 (N_2706,N_2688,N_2662);
nand U2707 (N_2707,N_2683,N_2651);
xor U2708 (N_2708,N_2661,N_2674);
or U2709 (N_2709,N_2665,N_2686);
nor U2710 (N_2710,N_2691,N_2658);
xnor U2711 (N_2711,N_2676,N_2675);
xnor U2712 (N_2712,N_2655,N_2657);
nand U2713 (N_2713,N_2659,N_2682);
and U2714 (N_2714,N_2678,N_2670);
and U2715 (N_2715,N_2696,N_2656);
or U2716 (N_2716,N_2672,N_2663);
and U2717 (N_2717,N_2671,N_2667);
or U2718 (N_2718,N_2694,N_2685);
or U2719 (N_2719,N_2690,N_2660);
nand U2720 (N_2720,N_2697,N_2693);
nor U2721 (N_2721,N_2689,N_2652);
or U2722 (N_2722,N_2687,N_2673);
nand U2723 (N_2723,N_2692,N_2664);
nand U2724 (N_2724,N_2684,N_2677);
nor U2725 (N_2725,N_2697,N_2692);
nor U2726 (N_2726,N_2662,N_2699);
or U2727 (N_2727,N_2666,N_2699);
or U2728 (N_2728,N_2650,N_2696);
nand U2729 (N_2729,N_2686,N_2661);
or U2730 (N_2730,N_2671,N_2690);
and U2731 (N_2731,N_2692,N_2654);
xnor U2732 (N_2732,N_2650,N_2687);
and U2733 (N_2733,N_2696,N_2652);
nand U2734 (N_2734,N_2676,N_2661);
or U2735 (N_2735,N_2678,N_2685);
xor U2736 (N_2736,N_2682,N_2695);
xor U2737 (N_2737,N_2659,N_2664);
nand U2738 (N_2738,N_2671,N_2672);
nor U2739 (N_2739,N_2671,N_2669);
nand U2740 (N_2740,N_2682,N_2685);
and U2741 (N_2741,N_2693,N_2656);
nor U2742 (N_2742,N_2670,N_2666);
and U2743 (N_2743,N_2692,N_2669);
nand U2744 (N_2744,N_2657,N_2650);
and U2745 (N_2745,N_2691,N_2652);
nand U2746 (N_2746,N_2698,N_2684);
nand U2747 (N_2747,N_2669,N_2673);
and U2748 (N_2748,N_2670,N_2688);
or U2749 (N_2749,N_2671,N_2660);
or U2750 (N_2750,N_2716,N_2704);
nor U2751 (N_2751,N_2740,N_2722);
and U2752 (N_2752,N_2744,N_2738);
or U2753 (N_2753,N_2727,N_2742);
and U2754 (N_2754,N_2732,N_2737);
nand U2755 (N_2755,N_2724,N_2701);
or U2756 (N_2756,N_2748,N_2710);
nand U2757 (N_2757,N_2707,N_2718);
and U2758 (N_2758,N_2726,N_2734);
or U2759 (N_2759,N_2746,N_2720);
nor U2760 (N_2760,N_2741,N_2743);
nand U2761 (N_2761,N_2747,N_2711);
xor U2762 (N_2762,N_2702,N_2729);
nor U2763 (N_2763,N_2749,N_2739);
and U2764 (N_2764,N_2712,N_2725);
and U2765 (N_2765,N_2700,N_2730);
and U2766 (N_2766,N_2735,N_2745);
nand U2767 (N_2767,N_2719,N_2723);
nor U2768 (N_2768,N_2715,N_2703);
nor U2769 (N_2769,N_2713,N_2714);
or U2770 (N_2770,N_2706,N_2733);
xnor U2771 (N_2771,N_2736,N_2731);
nand U2772 (N_2772,N_2717,N_2708);
xor U2773 (N_2773,N_2709,N_2705);
nand U2774 (N_2774,N_2721,N_2728);
nor U2775 (N_2775,N_2736,N_2748);
and U2776 (N_2776,N_2730,N_2706);
and U2777 (N_2777,N_2701,N_2715);
xor U2778 (N_2778,N_2704,N_2746);
or U2779 (N_2779,N_2743,N_2703);
xor U2780 (N_2780,N_2722,N_2716);
nand U2781 (N_2781,N_2746,N_2743);
xor U2782 (N_2782,N_2738,N_2703);
nor U2783 (N_2783,N_2715,N_2716);
nor U2784 (N_2784,N_2710,N_2732);
nand U2785 (N_2785,N_2700,N_2748);
xnor U2786 (N_2786,N_2746,N_2738);
nor U2787 (N_2787,N_2722,N_2728);
and U2788 (N_2788,N_2719,N_2746);
or U2789 (N_2789,N_2713,N_2729);
and U2790 (N_2790,N_2741,N_2704);
xor U2791 (N_2791,N_2747,N_2748);
nor U2792 (N_2792,N_2741,N_2733);
nor U2793 (N_2793,N_2737,N_2713);
nand U2794 (N_2794,N_2740,N_2706);
nor U2795 (N_2795,N_2710,N_2709);
xor U2796 (N_2796,N_2720,N_2742);
nor U2797 (N_2797,N_2713,N_2702);
nor U2798 (N_2798,N_2700,N_2714);
and U2799 (N_2799,N_2734,N_2718);
and U2800 (N_2800,N_2795,N_2774);
or U2801 (N_2801,N_2776,N_2755);
nor U2802 (N_2802,N_2750,N_2783);
xnor U2803 (N_2803,N_2767,N_2751);
nor U2804 (N_2804,N_2799,N_2797);
nor U2805 (N_2805,N_2756,N_2773);
xor U2806 (N_2806,N_2772,N_2786);
and U2807 (N_2807,N_2775,N_2794);
and U2808 (N_2808,N_2754,N_2759);
or U2809 (N_2809,N_2769,N_2761);
xnor U2810 (N_2810,N_2790,N_2762);
or U2811 (N_2811,N_2766,N_2793);
and U2812 (N_2812,N_2753,N_2789);
and U2813 (N_2813,N_2757,N_2791);
or U2814 (N_2814,N_2787,N_2780);
nor U2815 (N_2815,N_2798,N_2788);
nand U2816 (N_2816,N_2781,N_2752);
xor U2817 (N_2817,N_2768,N_2770);
nand U2818 (N_2818,N_2765,N_2785);
nor U2819 (N_2819,N_2792,N_2784);
nor U2820 (N_2820,N_2782,N_2771);
and U2821 (N_2821,N_2779,N_2778);
xnor U2822 (N_2822,N_2777,N_2758);
nor U2823 (N_2823,N_2764,N_2796);
xnor U2824 (N_2824,N_2763,N_2760);
or U2825 (N_2825,N_2783,N_2758);
nand U2826 (N_2826,N_2758,N_2798);
nand U2827 (N_2827,N_2776,N_2785);
nand U2828 (N_2828,N_2775,N_2781);
nor U2829 (N_2829,N_2789,N_2776);
nor U2830 (N_2830,N_2754,N_2787);
or U2831 (N_2831,N_2776,N_2760);
nor U2832 (N_2832,N_2750,N_2753);
and U2833 (N_2833,N_2751,N_2795);
xnor U2834 (N_2834,N_2793,N_2765);
nand U2835 (N_2835,N_2761,N_2759);
and U2836 (N_2836,N_2794,N_2751);
or U2837 (N_2837,N_2791,N_2759);
or U2838 (N_2838,N_2756,N_2776);
nor U2839 (N_2839,N_2763,N_2765);
nand U2840 (N_2840,N_2755,N_2774);
nand U2841 (N_2841,N_2783,N_2797);
and U2842 (N_2842,N_2794,N_2755);
and U2843 (N_2843,N_2788,N_2757);
nand U2844 (N_2844,N_2786,N_2795);
or U2845 (N_2845,N_2794,N_2760);
xnor U2846 (N_2846,N_2757,N_2771);
and U2847 (N_2847,N_2775,N_2756);
or U2848 (N_2848,N_2792,N_2780);
or U2849 (N_2849,N_2793,N_2751);
or U2850 (N_2850,N_2811,N_2812);
nor U2851 (N_2851,N_2800,N_2822);
and U2852 (N_2852,N_2842,N_2818);
or U2853 (N_2853,N_2847,N_2843);
nand U2854 (N_2854,N_2807,N_2830);
nor U2855 (N_2855,N_2838,N_2840);
xor U2856 (N_2856,N_2844,N_2810);
or U2857 (N_2857,N_2814,N_2832);
xor U2858 (N_2858,N_2846,N_2815);
xor U2859 (N_2859,N_2841,N_2821);
nand U2860 (N_2860,N_2803,N_2817);
and U2861 (N_2861,N_2845,N_2805);
nand U2862 (N_2862,N_2813,N_2802);
nor U2863 (N_2863,N_2831,N_2823);
or U2864 (N_2864,N_2816,N_2806);
or U2865 (N_2865,N_2837,N_2828);
nor U2866 (N_2866,N_2839,N_2819);
or U2867 (N_2867,N_2835,N_2826);
nand U2868 (N_2868,N_2825,N_2833);
and U2869 (N_2869,N_2801,N_2829);
nand U2870 (N_2870,N_2848,N_2827);
nor U2871 (N_2871,N_2820,N_2849);
nor U2872 (N_2872,N_2809,N_2836);
and U2873 (N_2873,N_2804,N_2834);
nor U2874 (N_2874,N_2808,N_2824);
nor U2875 (N_2875,N_2807,N_2823);
or U2876 (N_2876,N_2825,N_2803);
and U2877 (N_2877,N_2828,N_2843);
xnor U2878 (N_2878,N_2847,N_2820);
nor U2879 (N_2879,N_2840,N_2832);
nor U2880 (N_2880,N_2841,N_2840);
and U2881 (N_2881,N_2842,N_2833);
or U2882 (N_2882,N_2834,N_2813);
xor U2883 (N_2883,N_2837,N_2814);
or U2884 (N_2884,N_2800,N_2813);
or U2885 (N_2885,N_2838,N_2836);
or U2886 (N_2886,N_2844,N_2814);
nand U2887 (N_2887,N_2832,N_2836);
and U2888 (N_2888,N_2816,N_2821);
nand U2889 (N_2889,N_2806,N_2840);
xnor U2890 (N_2890,N_2807,N_2843);
nor U2891 (N_2891,N_2837,N_2826);
nor U2892 (N_2892,N_2839,N_2827);
xor U2893 (N_2893,N_2830,N_2825);
nand U2894 (N_2894,N_2844,N_2803);
nor U2895 (N_2895,N_2802,N_2834);
nor U2896 (N_2896,N_2801,N_2828);
or U2897 (N_2897,N_2825,N_2843);
xor U2898 (N_2898,N_2806,N_2813);
nand U2899 (N_2899,N_2827,N_2828);
nand U2900 (N_2900,N_2857,N_2882);
xnor U2901 (N_2901,N_2869,N_2887);
and U2902 (N_2902,N_2886,N_2863);
nor U2903 (N_2903,N_2893,N_2865);
and U2904 (N_2904,N_2895,N_2890);
nand U2905 (N_2905,N_2866,N_2870);
nand U2906 (N_2906,N_2860,N_2876);
nor U2907 (N_2907,N_2854,N_2855);
nand U2908 (N_2908,N_2871,N_2872);
xnor U2909 (N_2909,N_2889,N_2851);
nand U2910 (N_2910,N_2852,N_2879);
or U2911 (N_2911,N_2867,N_2877);
nand U2912 (N_2912,N_2875,N_2874);
or U2913 (N_2913,N_2896,N_2878);
nor U2914 (N_2914,N_2880,N_2850);
or U2915 (N_2915,N_2864,N_2858);
or U2916 (N_2916,N_2873,N_2856);
nand U2917 (N_2917,N_2899,N_2861);
nor U2918 (N_2918,N_2881,N_2898);
or U2919 (N_2919,N_2894,N_2888);
or U2920 (N_2920,N_2885,N_2862);
xor U2921 (N_2921,N_2859,N_2884);
nor U2922 (N_2922,N_2868,N_2883);
and U2923 (N_2923,N_2891,N_2853);
or U2924 (N_2924,N_2897,N_2892);
and U2925 (N_2925,N_2880,N_2890);
nand U2926 (N_2926,N_2873,N_2876);
and U2927 (N_2927,N_2860,N_2896);
or U2928 (N_2928,N_2866,N_2859);
nor U2929 (N_2929,N_2859,N_2857);
nand U2930 (N_2930,N_2876,N_2871);
or U2931 (N_2931,N_2852,N_2891);
or U2932 (N_2932,N_2855,N_2865);
nor U2933 (N_2933,N_2880,N_2879);
xnor U2934 (N_2934,N_2897,N_2856);
nand U2935 (N_2935,N_2865,N_2875);
or U2936 (N_2936,N_2864,N_2884);
and U2937 (N_2937,N_2873,N_2884);
and U2938 (N_2938,N_2871,N_2877);
xor U2939 (N_2939,N_2877,N_2882);
and U2940 (N_2940,N_2875,N_2892);
nor U2941 (N_2941,N_2855,N_2857);
or U2942 (N_2942,N_2892,N_2866);
xor U2943 (N_2943,N_2892,N_2865);
nor U2944 (N_2944,N_2851,N_2888);
xnor U2945 (N_2945,N_2858,N_2857);
nor U2946 (N_2946,N_2868,N_2891);
nor U2947 (N_2947,N_2870,N_2891);
and U2948 (N_2948,N_2886,N_2870);
nand U2949 (N_2949,N_2876,N_2898);
nor U2950 (N_2950,N_2946,N_2935);
or U2951 (N_2951,N_2932,N_2916);
nand U2952 (N_2952,N_2933,N_2943);
nor U2953 (N_2953,N_2942,N_2901);
nand U2954 (N_2954,N_2902,N_2947);
nor U2955 (N_2955,N_2941,N_2924);
xnor U2956 (N_2956,N_2904,N_2938);
or U2957 (N_2957,N_2925,N_2900);
nor U2958 (N_2958,N_2931,N_2903);
xnor U2959 (N_2959,N_2945,N_2936);
nand U2960 (N_2960,N_2928,N_2912);
nand U2961 (N_2961,N_2930,N_2927);
nand U2962 (N_2962,N_2937,N_2940);
nand U2963 (N_2963,N_2923,N_2939);
nand U2964 (N_2964,N_2908,N_2913);
or U2965 (N_2965,N_2917,N_2929);
nor U2966 (N_2966,N_2918,N_2906);
and U2967 (N_2967,N_2921,N_2907);
or U2968 (N_2968,N_2944,N_2914);
nor U2969 (N_2969,N_2905,N_2949);
and U2970 (N_2970,N_2926,N_2911);
nor U2971 (N_2971,N_2948,N_2934);
nand U2972 (N_2972,N_2922,N_2909);
and U2973 (N_2973,N_2910,N_2915);
or U2974 (N_2974,N_2920,N_2919);
or U2975 (N_2975,N_2933,N_2911);
and U2976 (N_2976,N_2915,N_2949);
nor U2977 (N_2977,N_2911,N_2946);
xnor U2978 (N_2978,N_2944,N_2913);
and U2979 (N_2979,N_2920,N_2944);
and U2980 (N_2980,N_2915,N_2938);
nor U2981 (N_2981,N_2922,N_2906);
and U2982 (N_2982,N_2923,N_2947);
and U2983 (N_2983,N_2916,N_2927);
xor U2984 (N_2984,N_2935,N_2911);
xnor U2985 (N_2985,N_2942,N_2909);
xnor U2986 (N_2986,N_2930,N_2944);
and U2987 (N_2987,N_2947,N_2942);
nand U2988 (N_2988,N_2940,N_2905);
nor U2989 (N_2989,N_2907,N_2927);
nand U2990 (N_2990,N_2941,N_2936);
or U2991 (N_2991,N_2915,N_2908);
xor U2992 (N_2992,N_2918,N_2943);
or U2993 (N_2993,N_2921,N_2948);
or U2994 (N_2994,N_2946,N_2944);
xor U2995 (N_2995,N_2905,N_2931);
nor U2996 (N_2996,N_2942,N_2920);
nand U2997 (N_2997,N_2909,N_2949);
and U2998 (N_2998,N_2921,N_2915);
xor U2999 (N_2999,N_2912,N_2919);
nor UO_0 (O_0,N_2959,N_2957);
nand UO_1 (O_1,N_2956,N_2992);
nand UO_2 (O_2,N_2972,N_2998);
xnor UO_3 (O_3,N_2961,N_2988);
nor UO_4 (O_4,N_2967,N_2958);
xor UO_5 (O_5,N_2995,N_2966);
and UO_6 (O_6,N_2974,N_2965);
xor UO_7 (O_7,N_2994,N_2971);
nand UO_8 (O_8,N_2984,N_2968);
nor UO_9 (O_9,N_2953,N_2973);
nand UO_10 (O_10,N_2986,N_2969);
or UO_11 (O_11,N_2987,N_2962);
nor UO_12 (O_12,N_2982,N_2996);
nor UO_13 (O_13,N_2970,N_2964);
or UO_14 (O_14,N_2954,N_2981);
and UO_15 (O_15,N_2980,N_2952);
nor UO_16 (O_16,N_2960,N_2993);
xnor UO_17 (O_17,N_2976,N_2963);
and UO_18 (O_18,N_2991,N_2978);
xor UO_19 (O_19,N_2977,N_2989);
or UO_20 (O_20,N_2983,N_2997);
xnor UO_21 (O_21,N_2999,N_2979);
or UO_22 (O_22,N_2951,N_2990);
or UO_23 (O_23,N_2955,N_2950);
or UO_24 (O_24,N_2975,N_2985);
nor UO_25 (O_25,N_2958,N_2964);
nand UO_26 (O_26,N_2980,N_2962);
nand UO_27 (O_27,N_2980,N_2982);
nand UO_28 (O_28,N_2954,N_2965);
nor UO_29 (O_29,N_2963,N_2996);
nor UO_30 (O_30,N_2971,N_2966);
nand UO_31 (O_31,N_2986,N_2961);
nand UO_32 (O_32,N_2979,N_2961);
or UO_33 (O_33,N_2993,N_2957);
nor UO_34 (O_34,N_2993,N_2989);
nor UO_35 (O_35,N_2991,N_2977);
xor UO_36 (O_36,N_2963,N_2990);
and UO_37 (O_37,N_2964,N_2950);
nand UO_38 (O_38,N_2952,N_2999);
nor UO_39 (O_39,N_2979,N_2969);
and UO_40 (O_40,N_2992,N_2964);
nand UO_41 (O_41,N_2967,N_2972);
xor UO_42 (O_42,N_2983,N_2969);
nand UO_43 (O_43,N_2974,N_2961);
nand UO_44 (O_44,N_2998,N_2986);
and UO_45 (O_45,N_2995,N_2955);
nand UO_46 (O_46,N_2970,N_2965);
and UO_47 (O_47,N_2959,N_2963);
nand UO_48 (O_48,N_2958,N_2986);
and UO_49 (O_49,N_2983,N_2967);
or UO_50 (O_50,N_2978,N_2981);
or UO_51 (O_51,N_2979,N_2967);
xor UO_52 (O_52,N_2982,N_2993);
nor UO_53 (O_53,N_2994,N_2968);
and UO_54 (O_54,N_2965,N_2968);
and UO_55 (O_55,N_2963,N_2951);
nor UO_56 (O_56,N_2984,N_2987);
xnor UO_57 (O_57,N_2956,N_2984);
nor UO_58 (O_58,N_2989,N_2973);
and UO_59 (O_59,N_2968,N_2998);
xor UO_60 (O_60,N_2993,N_2974);
nand UO_61 (O_61,N_2996,N_2991);
xnor UO_62 (O_62,N_2965,N_2960);
or UO_63 (O_63,N_2985,N_2981);
nand UO_64 (O_64,N_2992,N_2986);
xnor UO_65 (O_65,N_2973,N_2969);
xnor UO_66 (O_66,N_2980,N_2976);
nand UO_67 (O_67,N_2977,N_2997);
and UO_68 (O_68,N_2953,N_2994);
nor UO_69 (O_69,N_2967,N_2951);
nor UO_70 (O_70,N_2956,N_2995);
and UO_71 (O_71,N_2990,N_2958);
xor UO_72 (O_72,N_2964,N_2983);
and UO_73 (O_73,N_2958,N_2973);
nor UO_74 (O_74,N_2992,N_2981);
nor UO_75 (O_75,N_2961,N_2983);
nand UO_76 (O_76,N_2951,N_2977);
nand UO_77 (O_77,N_2997,N_2964);
nand UO_78 (O_78,N_2957,N_2955);
xnor UO_79 (O_79,N_2973,N_2975);
or UO_80 (O_80,N_2986,N_2954);
nor UO_81 (O_81,N_2993,N_2996);
nor UO_82 (O_82,N_2991,N_2997);
and UO_83 (O_83,N_2963,N_2978);
nand UO_84 (O_84,N_2978,N_2979);
or UO_85 (O_85,N_2995,N_2980);
or UO_86 (O_86,N_2972,N_2969);
and UO_87 (O_87,N_2950,N_2966);
xor UO_88 (O_88,N_2987,N_2966);
or UO_89 (O_89,N_2970,N_2998);
and UO_90 (O_90,N_2955,N_2974);
and UO_91 (O_91,N_2990,N_2954);
xor UO_92 (O_92,N_2977,N_2976);
xor UO_93 (O_93,N_2971,N_2951);
and UO_94 (O_94,N_2974,N_2975);
xnor UO_95 (O_95,N_2982,N_2963);
nor UO_96 (O_96,N_2954,N_2974);
and UO_97 (O_97,N_2966,N_2972);
and UO_98 (O_98,N_2962,N_2971);
nand UO_99 (O_99,N_2973,N_2992);
nand UO_100 (O_100,N_2958,N_2956);
nand UO_101 (O_101,N_2999,N_2954);
and UO_102 (O_102,N_2964,N_2975);
nor UO_103 (O_103,N_2984,N_2963);
or UO_104 (O_104,N_2950,N_2962);
nor UO_105 (O_105,N_2974,N_2967);
nor UO_106 (O_106,N_2985,N_2953);
nand UO_107 (O_107,N_2977,N_2958);
xor UO_108 (O_108,N_2984,N_2996);
xnor UO_109 (O_109,N_2958,N_2961);
or UO_110 (O_110,N_2952,N_2960);
nand UO_111 (O_111,N_2954,N_2991);
nand UO_112 (O_112,N_2975,N_2952);
or UO_113 (O_113,N_2954,N_2980);
or UO_114 (O_114,N_2987,N_2973);
nor UO_115 (O_115,N_2971,N_2957);
or UO_116 (O_116,N_2964,N_2976);
nand UO_117 (O_117,N_2962,N_2982);
or UO_118 (O_118,N_2987,N_2981);
nor UO_119 (O_119,N_2996,N_2968);
xnor UO_120 (O_120,N_2950,N_2968);
and UO_121 (O_121,N_2960,N_2973);
and UO_122 (O_122,N_2995,N_2968);
nand UO_123 (O_123,N_2964,N_2980);
xor UO_124 (O_124,N_2995,N_2964);
xor UO_125 (O_125,N_2959,N_2955);
xor UO_126 (O_126,N_2975,N_2972);
and UO_127 (O_127,N_2962,N_2975);
or UO_128 (O_128,N_2990,N_2972);
or UO_129 (O_129,N_2954,N_2970);
nand UO_130 (O_130,N_2962,N_2994);
xor UO_131 (O_131,N_2990,N_2952);
xnor UO_132 (O_132,N_2969,N_2993);
and UO_133 (O_133,N_2955,N_2986);
xnor UO_134 (O_134,N_2967,N_2976);
and UO_135 (O_135,N_2976,N_2997);
nand UO_136 (O_136,N_2981,N_2996);
or UO_137 (O_137,N_2975,N_2958);
or UO_138 (O_138,N_2969,N_2958);
and UO_139 (O_139,N_2978,N_2967);
nor UO_140 (O_140,N_2984,N_2998);
nor UO_141 (O_141,N_2958,N_2974);
xnor UO_142 (O_142,N_2960,N_2994);
nor UO_143 (O_143,N_2982,N_2973);
nor UO_144 (O_144,N_2998,N_2973);
or UO_145 (O_145,N_2953,N_2972);
and UO_146 (O_146,N_2954,N_2993);
and UO_147 (O_147,N_2963,N_2981);
nor UO_148 (O_148,N_2994,N_2967);
xnor UO_149 (O_149,N_2979,N_2994);
nand UO_150 (O_150,N_2965,N_2999);
nor UO_151 (O_151,N_2967,N_2988);
nand UO_152 (O_152,N_2969,N_2996);
nand UO_153 (O_153,N_2957,N_2950);
or UO_154 (O_154,N_2991,N_2963);
nand UO_155 (O_155,N_2996,N_2973);
nand UO_156 (O_156,N_2967,N_2963);
or UO_157 (O_157,N_2987,N_2964);
and UO_158 (O_158,N_2961,N_2999);
and UO_159 (O_159,N_2988,N_2989);
nand UO_160 (O_160,N_2960,N_2972);
nand UO_161 (O_161,N_2999,N_2978);
nor UO_162 (O_162,N_2966,N_2955);
or UO_163 (O_163,N_2998,N_2963);
xnor UO_164 (O_164,N_2979,N_2993);
or UO_165 (O_165,N_2959,N_2983);
nand UO_166 (O_166,N_2952,N_2964);
nor UO_167 (O_167,N_2971,N_2981);
xnor UO_168 (O_168,N_2991,N_2988);
nor UO_169 (O_169,N_2999,N_2970);
nand UO_170 (O_170,N_2978,N_2952);
and UO_171 (O_171,N_2950,N_2983);
nand UO_172 (O_172,N_2995,N_2950);
nand UO_173 (O_173,N_2999,N_2973);
xnor UO_174 (O_174,N_2968,N_2986);
nor UO_175 (O_175,N_2965,N_2987);
or UO_176 (O_176,N_2968,N_2956);
or UO_177 (O_177,N_2960,N_2962);
and UO_178 (O_178,N_2999,N_2994);
nand UO_179 (O_179,N_2969,N_2999);
nand UO_180 (O_180,N_2987,N_2988);
nor UO_181 (O_181,N_2958,N_2984);
nor UO_182 (O_182,N_2989,N_2958);
or UO_183 (O_183,N_2964,N_2996);
xor UO_184 (O_184,N_2954,N_2988);
and UO_185 (O_185,N_2970,N_2971);
nand UO_186 (O_186,N_2979,N_2990);
and UO_187 (O_187,N_2963,N_2987);
or UO_188 (O_188,N_2966,N_2964);
and UO_189 (O_189,N_2969,N_2968);
nor UO_190 (O_190,N_2959,N_2961);
or UO_191 (O_191,N_2986,N_2994);
nand UO_192 (O_192,N_2952,N_2971);
nand UO_193 (O_193,N_2961,N_2963);
nor UO_194 (O_194,N_2967,N_2954);
xor UO_195 (O_195,N_2971,N_2987);
nand UO_196 (O_196,N_2977,N_2953);
or UO_197 (O_197,N_2981,N_2961);
nor UO_198 (O_198,N_2973,N_2962);
nor UO_199 (O_199,N_2971,N_2973);
or UO_200 (O_200,N_2959,N_2950);
or UO_201 (O_201,N_2971,N_2950);
and UO_202 (O_202,N_2965,N_2993);
and UO_203 (O_203,N_2960,N_2997);
xor UO_204 (O_204,N_2999,N_2993);
xor UO_205 (O_205,N_2980,N_2965);
nor UO_206 (O_206,N_2950,N_2989);
nand UO_207 (O_207,N_2972,N_2984);
nand UO_208 (O_208,N_2995,N_2978);
or UO_209 (O_209,N_2979,N_2982);
and UO_210 (O_210,N_2996,N_2974);
nand UO_211 (O_211,N_2953,N_2961);
nand UO_212 (O_212,N_2972,N_2962);
nand UO_213 (O_213,N_2986,N_2956);
and UO_214 (O_214,N_2990,N_2982);
or UO_215 (O_215,N_2976,N_2970);
and UO_216 (O_216,N_2963,N_2956);
and UO_217 (O_217,N_2990,N_2984);
nand UO_218 (O_218,N_2988,N_2986);
and UO_219 (O_219,N_2970,N_2978);
xnor UO_220 (O_220,N_2982,N_2987);
or UO_221 (O_221,N_2989,N_2996);
and UO_222 (O_222,N_2967,N_2952);
or UO_223 (O_223,N_2968,N_2980);
nand UO_224 (O_224,N_2987,N_2989);
nor UO_225 (O_225,N_2970,N_2960);
nand UO_226 (O_226,N_2986,N_2976);
nor UO_227 (O_227,N_2978,N_2986);
xor UO_228 (O_228,N_2995,N_2970);
nand UO_229 (O_229,N_2954,N_2984);
and UO_230 (O_230,N_2985,N_2982);
or UO_231 (O_231,N_2992,N_2957);
nand UO_232 (O_232,N_2950,N_2998);
nand UO_233 (O_233,N_2982,N_2989);
or UO_234 (O_234,N_2955,N_2989);
and UO_235 (O_235,N_2953,N_2988);
nand UO_236 (O_236,N_2978,N_2959);
xor UO_237 (O_237,N_2958,N_2982);
xor UO_238 (O_238,N_2975,N_2960);
and UO_239 (O_239,N_2959,N_2956);
xor UO_240 (O_240,N_2981,N_2965);
and UO_241 (O_241,N_2998,N_2989);
and UO_242 (O_242,N_2983,N_2979);
nand UO_243 (O_243,N_2992,N_2950);
nand UO_244 (O_244,N_2978,N_2977);
nor UO_245 (O_245,N_2992,N_2993);
or UO_246 (O_246,N_2991,N_2971);
nand UO_247 (O_247,N_2969,N_2970);
and UO_248 (O_248,N_2983,N_2957);
or UO_249 (O_249,N_2963,N_2964);
or UO_250 (O_250,N_2995,N_2976);
and UO_251 (O_251,N_2969,N_2997);
and UO_252 (O_252,N_2963,N_2994);
or UO_253 (O_253,N_2952,N_2953);
nand UO_254 (O_254,N_2988,N_2979);
nor UO_255 (O_255,N_2960,N_2999);
nor UO_256 (O_256,N_2981,N_2967);
or UO_257 (O_257,N_2978,N_2961);
xor UO_258 (O_258,N_2992,N_2955);
or UO_259 (O_259,N_2977,N_2964);
nor UO_260 (O_260,N_2989,N_2953);
or UO_261 (O_261,N_2969,N_2977);
or UO_262 (O_262,N_2957,N_2990);
or UO_263 (O_263,N_2969,N_2998);
nor UO_264 (O_264,N_2950,N_2973);
xor UO_265 (O_265,N_2997,N_2966);
nor UO_266 (O_266,N_2987,N_2990);
nor UO_267 (O_267,N_2993,N_2997);
or UO_268 (O_268,N_2962,N_2954);
nor UO_269 (O_269,N_2967,N_2955);
xor UO_270 (O_270,N_2975,N_2970);
and UO_271 (O_271,N_2951,N_2992);
or UO_272 (O_272,N_2961,N_2989);
nand UO_273 (O_273,N_2971,N_2989);
xor UO_274 (O_274,N_2957,N_2958);
nor UO_275 (O_275,N_2974,N_2966);
nand UO_276 (O_276,N_2990,N_2976);
nor UO_277 (O_277,N_2968,N_2967);
and UO_278 (O_278,N_2974,N_2959);
xnor UO_279 (O_279,N_2957,N_2984);
and UO_280 (O_280,N_2951,N_2998);
xor UO_281 (O_281,N_2974,N_2950);
and UO_282 (O_282,N_2978,N_2951);
nand UO_283 (O_283,N_2962,N_2998);
xnor UO_284 (O_284,N_2970,N_2961);
nand UO_285 (O_285,N_2963,N_2952);
or UO_286 (O_286,N_2955,N_2964);
and UO_287 (O_287,N_2992,N_2959);
and UO_288 (O_288,N_2996,N_2955);
nand UO_289 (O_289,N_2983,N_2987);
nor UO_290 (O_290,N_2991,N_2962);
or UO_291 (O_291,N_2958,N_2955);
and UO_292 (O_292,N_2997,N_2988);
nor UO_293 (O_293,N_2969,N_2952);
nor UO_294 (O_294,N_2983,N_2999);
xnor UO_295 (O_295,N_2953,N_2969);
xnor UO_296 (O_296,N_2951,N_2964);
nor UO_297 (O_297,N_2958,N_2963);
and UO_298 (O_298,N_2999,N_2951);
and UO_299 (O_299,N_2962,N_2977);
xnor UO_300 (O_300,N_2966,N_2994);
and UO_301 (O_301,N_2966,N_2985);
xnor UO_302 (O_302,N_2982,N_2976);
nand UO_303 (O_303,N_2978,N_2988);
xor UO_304 (O_304,N_2985,N_2987);
xor UO_305 (O_305,N_2953,N_2993);
xor UO_306 (O_306,N_2988,N_2998);
nand UO_307 (O_307,N_2975,N_2991);
nand UO_308 (O_308,N_2976,N_2960);
nor UO_309 (O_309,N_2993,N_2967);
nand UO_310 (O_310,N_2976,N_2956);
xnor UO_311 (O_311,N_2952,N_2974);
and UO_312 (O_312,N_2990,N_2973);
and UO_313 (O_313,N_2997,N_2980);
xnor UO_314 (O_314,N_2995,N_2992);
or UO_315 (O_315,N_2994,N_2965);
or UO_316 (O_316,N_2970,N_2968);
nor UO_317 (O_317,N_2968,N_2989);
or UO_318 (O_318,N_2975,N_2968);
xnor UO_319 (O_319,N_2961,N_2965);
nand UO_320 (O_320,N_2999,N_2988);
and UO_321 (O_321,N_2978,N_2968);
or UO_322 (O_322,N_2954,N_2982);
nand UO_323 (O_323,N_2953,N_2955);
nand UO_324 (O_324,N_2957,N_2994);
nor UO_325 (O_325,N_2970,N_2983);
and UO_326 (O_326,N_2985,N_2995);
nand UO_327 (O_327,N_2960,N_2977);
nor UO_328 (O_328,N_2989,N_2986);
nor UO_329 (O_329,N_2987,N_2991);
nand UO_330 (O_330,N_2981,N_2957);
nor UO_331 (O_331,N_2992,N_2954);
nand UO_332 (O_332,N_2959,N_2975);
nand UO_333 (O_333,N_2980,N_2957);
nand UO_334 (O_334,N_2987,N_2958);
or UO_335 (O_335,N_2972,N_2958);
and UO_336 (O_336,N_2996,N_2965);
nand UO_337 (O_337,N_2994,N_2983);
and UO_338 (O_338,N_2974,N_2985);
or UO_339 (O_339,N_2973,N_2968);
nor UO_340 (O_340,N_2951,N_2979);
nand UO_341 (O_341,N_2998,N_2983);
nand UO_342 (O_342,N_2966,N_2961);
and UO_343 (O_343,N_2976,N_2955);
and UO_344 (O_344,N_2963,N_2997);
nor UO_345 (O_345,N_2985,N_2968);
or UO_346 (O_346,N_2968,N_2981);
nor UO_347 (O_347,N_2975,N_2995);
or UO_348 (O_348,N_2987,N_2968);
nor UO_349 (O_349,N_2968,N_2971);
nor UO_350 (O_350,N_2974,N_2984);
xnor UO_351 (O_351,N_2953,N_2998);
or UO_352 (O_352,N_2979,N_2972);
and UO_353 (O_353,N_2967,N_2964);
and UO_354 (O_354,N_2975,N_2997);
nor UO_355 (O_355,N_2990,N_2999);
xor UO_356 (O_356,N_2963,N_2974);
nor UO_357 (O_357,N_2982,N_2969);
and UO_358 (O_358,N_2955,N_2979);
nand UO_359 (O_359,N_2976,N_2962);
and UO_360 (O_360,N_2995,N_2991);
and UO_361 (O_361,N_2983,N_2955);
and UO_362 (O_362,N_2988,N_2958);
nand UO_363 (O_363,N_2997,N_2951);
or UO_364 (O_364,N_2971,N_2997);
and UO_365 (O_365,N_2971,N_2980);
and UO_366 (O_366,N_2966,N_2967);
xor UO_367 (O_367,N_2970,N_2974);
and UO_368 (O_368,N_2975,N_2993);
and UO_369 (O_369,N_2984,N_2952);
xnor UO_370 (O_370,N_2969,N_2989);
xnor UO_371 (O_371,N_2980,N_2978);
and UO_372 (O_372,N_2996,N_2998);
xnor UO_373 (O_373,N_2984,N_2995);
nand UO_374 (O_374,N_2953,N_2950);
xor UO_375 (O_375,N_2957,N_2985);
nor UO_376 (O_376,N_2992,N_2998);
or UO_377 (O_377,N_2954,N_2973);
nand UO_378 (O_378,N_2988,N_2996);
xnor UO_379 (O_379,N_2975,N_2977);
and UO_380 (O_380,N_2957,N_2974);
nor UO_381 (O_381,N_2976,N_2953);
nor UO_382 (O_382,N_2995,N_2962);
or UO_383 (O_383,N_2969,N_2992);
or UO_384 (O_384,N_2960,N_2984);
or UO_385 (O_385,N_2986,N_2999);
xnor UO_386 (O_386,N_2966,N_2981);
and UO_387 (O_387,N_2971,N_2961);
and UO_388 (O_388,N_2989,N_2985);
nor UO_389 (O_389,N_2956,N_2966);
nand UO_390 (O_390,N_2951,N_2959);
nor UO_391 (O_391,N_2967,N_2997);
nand UO_392 (O_392,N_2977,N_2950);
and UO_393 (O_393,N_2966,N_2998);
or UO_394 (O_394,N_2962,N_2997);
xnor UO_395 (O_395,N_2998,N_2965);
nor UO_396 (O_396,N_2959,N_2965);
and UO_397 (O_397,N_2962,N_2970);
xnor UO_398 (O_398,N_2997,N_2999);
or UO_399 (O_399,N_2973,N_2993);
nor UO_400 (O_400,N_2979,N_2997);
xnor UO_401 (O_401,N_2998,N_2975);
and UO_402 (O_402,N_2985,N_2962);
nor UO_403 (O_403,N_2996,N_2999);
or UO_404 (O_404,N_2972,N_2961);
and UO_405 (O_405,N_2998,N_2981);
nand UO_406 (O_406,N_2957,N_2966);
nand UO_407 (O_407,N_2999,N_2974);
nor UO_408 (O_408,N_2993,N_2984);
nor UO_409 (O_409,N_2986,N_2983);
nor UO_410 (O_410,N_2988,N_2959);
or UO_411 (O_411,N_2992,N_2979);
and UO_412 (O_412,N_2954,N_2976);
xor UO_413 (O_413,N_2976,N_2966);
or UO_414 (O_414,N_2999,N_2964);
xor UO_415 (O_415,N_2965,N_2956);
and UO_416 (O_416,N_2975,N_2965);
or UO_417 (O_417,N_2980,N_2977);
or UO_418 (O_418,N_2983,N_2971);
nand UO_419 (O_419,N_2957,N_2976);
xnor UO_420 (O_420,N_2981,N_2974);
nor UO_421 (O_421,N_2965,N_2976);
nand UO_422 (O_422,N_2951,N_2995);
or UO_423 (O_423,N_2956,N_2972);
or UO_424 (O_424,N_2985,N_2988);
nand UO_425 (O_425,N_2995,N_2993);
xor UO_426 (O_426,N_2987,N_2976);
or UO_427 (O_427,N_2987,N_2957);
and UO_428 (O_428,N_2972,N_2968);
and UO_429 (O_429,N_2977,N_2984);
or UO_430 (O_430,N_2991,N_2964);
nor UO_431 (O_431,N_2994,N_2985);
nand UO_432 (O_432,N_2951,N_2972);
xnor UO_433 (O_433,N_2966,N_2993);
nor UO_434 (O_434,N_2963,N_2992);
or UO_435 (O_435,N_2960,N_2958);
and UO_436 (O_436,N_2961,N_2996);
xnor UO_437 (O_437,N_2959,N_2976);
nor UO_438 (O_438,N_2961,N_2968);
nor UO_439 (O_439,N_2997,N_2972);
nand UO_440 (O_440,N_2988,N_2982);
nand UO_441 (O_441,N_2999,N_2998);
or UO_442 (O_442,N_2987,N_2952);
and UO_443 (O_443,N_2996,N_2986);
nand UO_444 (O_444,N_2982,N_2971);
and UO_445 (O_445,N_2959,N_2964);
or UO_446 (O_446,N_2963,N_2986);
and UO_447 (O_447,N_2991,N_2956);
nor UO_448 (O_448,N_2972,N_2963);
nor UO_449 (O_449,N_2971,N_2988);
xnor UO_450 (O_450,N_2961,N_2997);
or UO_451 (O_451,N_2969,N_2991);
nand UO_452 (O_452,N_2964,N_2984);
or UO_453 (O_453,N_2975,N_2978);
nand UO_454 (O_454,N_2982,N_2978);
nor UO_455 (O_455,N_2980,N_2974);
nor UO_456 (O_456,N_2994,N_2980);
and UO_457 (O_457,N_2998,N_2991);
nand UO_458 (O_458,N_2990,N_2974);
nand UO_459 (O_459,N_2995,N_2959);
or UO_460 (O_460,N_2990,N_2956);
or UO_461 (O_461,N_2999,N_2980);
or UO_462 (O_462,N_2953,N_2999);
xor UO_463 (O_463,N_2986,N_2953);
nand UO_464 (O_464,N_2968,N_2951);
xnor UO_465 (O_465,N_2979,N_2973);
nand UO_466 (O_466,N_2952,N_2955);
or UO_467 (O_467,N_2965,N_2990);
nand UO_468 (O_468,N_2958,N_2995);
and UO_469 (O_469,N_2959,N_2981);
nor UO_470 (O_470,N_2970,N_2987);
nand UO_471 (O_471,N_2960,N_2987);
and UO_472 (O_472,N_2979,N_2957);
or UO_473 (O_473,N_2998,N_2958);
xnor UO_474 (O_474,N_2995,N_2996);
nand UO_475 (O_475,N_2990,N_2988);
nand UO_476 (O_476,N_2954,N_2989);
nor UO_477 (O_477,N_2952,N_2958);
nand UO_478 (O_478,N_2958,N_2965);
and UO_479 (O_479,N_2984,N_2967);
nand UO_480 (O_480,N_2983,N_2988);
nor UO_481 (O_481,N_2991,N_2972);
nand UO_482 (O_482,N_2954,N_2969);
nor UO_483 (O_483,N_2972,N_2955);
and UO_484 (O_484,N_2983,N_2960);
xor UO_485 (O_485,N_2979,N_2975);
or UO_486 (O_486,N_2997,N_2950);
and UO_487 (O_487,N_2954,N_2951);
or UO_488 (O_488,N_2965,N_2988);
or UO_489 (O_489,N_2960,N_2996);
or UO_490 (O_490,N_2981,N_2969);
or UO_491 (O_491,N_2983,N_2965);
nand UO_492 (O_492,N_2989,N_2963);
or UO_493 (O_493,N_2952,N_2998);
and UO_494 (O_494,N_2986,N_2967);
nor UO_495 (O_495,N_2992,N_2977);
or UO_496 (O_496,N_2989,N_2951);
or UO_497 (O_497,N_2952,N_2956);
xnor UO_498 (O_498,N_2995,N_2979);
nor UO_499 (O_499,N_2986,N_2977);
endmodule