module basic_3000_30000_3500_6_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1736,In_2397);
or U1 (N_1,In_2612,In_57);
xnor U2 (N_2,In_318,In_1776);
nor U3 (N_3,In_2507,In_2090);
and U4 (N_4,In_433,In_2384);
or U5 (N_5,In_2263,In_820);
xor U6 (N_6,In_2874,In_2050);
and U7 (N_7,In_1810,In_677);
and U8 (N_8,In_1099,In_1060);
nor U9 (N_9,In_2550,In_2887);
and U10 (N_10,In_1301,In_2149);
xnor U11 (N_11,In_1862,In_354);
nor U12 (N_12,In_587,In_1198);
xnor U13 (N_13,In_2759,In_878);
and U14 (N_14,In_2431,In_2578);
and U15 (N_15,In_394,In_1430);
xor U16 (N_16,In_213,In_2861);
and U17 (N_17,In_1069,In_1408);
and U18 (N_18,In_1400,In_1108);
nand U19 (N_19,In_2940,In_1895);
xnor U20 (N_20,In_1019,In_1002);
or U21 (N_21,In_1160,In_1864);
nand U22 (N_22,In_1992,In_325);
and U23 (N_23,In_1815,In_1879);
nand U24 (N_24,In_2753,In_1372);
nor U25 (N_25,In_74,In_558);
nor U26 (N_26,In_173,In_1312);
or U27 (N_27,In_1467,In_602);
or U28 (N_28,In_2453,In_1351);
and U29 (N_29,In_2497,In_1650);
nor U30 (N_30,In_1619,In_2871);
or U31 (N_31,In_2772,In_1696);
nor U32 (N_32,In_2699,In_2601);
xnor U33 (N_33,In_2985,In_2841);
nand U34 (N_34,In_431,In_1273);
or U35 (N_35,In_653,In_2478);
nor U36 (N_36,In_2820,In_902);
or U37 (N_37,In_2588,In_687);
and U38 (N_38,In_5,In_942);
or U39 (N_39,In_1582,In_829);
nor U40 (N_40,In_2230,In_307);
xor U41 (N_41,In_969,In_1017);
and U42 (N_42,In_1603,In_2857);
and U43 (N_43,In_299,In_1536);
or U44 (N_44,In_957,In_2071);
nand U45 (N_45,In_2986,In_1165);
nor U46 (N_46,In_999,In_1898);
nor U47 (N_47,In_35,In_1846);
nand U48 (N_48,In_2977,In_2675);
xor U49 (N_49,In_808,In_718);
or U50 (N_50,In_1770,In_792);
and U51 (N_51,In_1739,In_1018);
or U52 (N_52,In_2734,In_2850);
nor U53 (N_53,In_2953,In_1322);
xor U54 (N_54,In_1252,In_2942);
and U55 (N_55,In_1791,In_126);
nand U56 (N_56,In_1595,In_76);
nor U57 (N_57,In_21,In_2632);
xnor U58 (N_58,In_2115,In_2282);
nand U59 (N_59,In_2698,In_1462);
and U60 (N_60,In_1821,In_1882);
nor U61 (N_61,In_1440,In_1071);
nand U62 (N_62,In_2472,In_1174);
or U63 (N_63,In_108,In_2756);
xor U64 (N_64,In_2014,In_1422);
nor U65 (N_65,In_2564,In_392);
nand U66 (N_66,In_2034,In_1403);
or U67 (N_67,In_1214,In_236);
and U68 (N_68,In_1386,In_965);
nor U69 (N_69,In_331,In_713);
nor U70 (N_70,In_1905,In_549);
or U71 (N_71,In_1253,In_1208);
and U72 (N_72,In_2521,In_1145);
nor U73 (N_73,In_921,In_405);
and U74 (N_74,In_1124,In_1218);
nand U75 (N_75,In_545,In_1872);
xor U76 (N_76,In_658,In_632);
xor U77 (N_77,In_1844,In_1067);
and U78 (N_78,In_2931,In_2897);
xnor U79 (N_79,In_2875,In_2943);
nor U80 (N_80,In_692,In_890);
or U81 (N_81,In_1284,In_1868);
nor U82 (N_82,In_1854,In_20);
or U83 (N_83,In_2215,In_2720);
or U84 (N_84,In_1550,In_2484);
or U85 (N_85,In_2278,In_815);
and U86 (N_86,In_2370,In_1149);
nand U87 (N_87,In_1795,In_1187);
or U88 (N_88,In_2829,In_642);
or U89 (N_89,In_2555,In_2424);
and U90 (N_90,In_1327,In_2800);
or U91 (N_91,In_427,In_852);
or U92 (N_92,In_2962,In_2690);
or U93 (N_93,In_168,In_1936);
or U94 (N_94,In_860,In_409);
nand U95 (N_95,In_2427,In_2520);
xor U96 (N_96,In_104,In_1420);
or U97 (N_97,In_577,In_998);
nand U98 (N_98,In_2996,In_744);
nor U99 (N_99,In_2523,In_2443);
and U100 (N_100,In_943,In_8);
nor U101 (N_101,In_458,In_248);
and U102 (N_102,In_2544,In_2651);
or U103 (N_103,In_488,In_1942);
and U104 (N_104,In_862,In_2480);
nor U105 (N_105,In_2456,In_1633);
nand U106 (N_106,In_1326,In_2912);
nor U107 (N_107,In_1200,In_2190);
nor U108 (N_108,In_2933,In_2979);
nand U109 (N_109,In_570,In_2538);
nand U110 (N_110,In_241,In_1238);
or U111 (N_111,In_1998,In_1323);
and U112 (N_112,In_2131,In_529);
nor U113 (N_113,In_1672,In_2814);
nand U114 (N_114,In_1801,In_1355);
and U115 (N_115,In_2316,In_1688);
and U116 (N_116,In_1941,In_1438);
nand U117 (N_117,In_2364,In_956);
nor U118 (N_118,In_2870,In_1144);
nand U119 (N_119,In_784,In_2628);
xor U120 (N_120,In_2046,In_94);
nand U121 (N_121,In_941,In_1677);
nor U122 (N_122,In_2091,In_668);
or U123 (N_123,In_1909,In_2893);
nor U124 (N_124,In_1051,In_1883);
nand U125 (N_125,In_2633,In_2345);
or U126 (N_126,In_2062,In_2303);
nand U127 (N_127,In_2540,In_2929);
or U128 (N_128,In_2923,In_2958);
xnor U129 (N_129,In_865,In_1915);
nor U130 (N_130,In_1107,In_531);
and U131 (N_131,In_1041,In_1388);
xor U132 (N_132,In_2832,In_13);
nor U133 (N_133,In_2179,In_2495);
xnor U134 (N_134,In_1518,In_2666);
and U135 (N_135,In_2355,In_1399);
and U136 (N_136,In_1084,In_2739);
and U137 (N_137,In_398,In_1102);
or U138 (N_138,In_2679,In_169);
nor U139 (N_139,In_2853,In_1893);
and U140 (N_140,In_1162,In_1761);
or U141 (N_141,In_1395,In_159);
or U142 (N_142,In_970,In_2199);
nor U143 (N_143,In_2765,In_982);
nor U144 (N_144,In_2662,In_1207);
nand U145 (N_145,In_1638,In_216);
or U146 (N_146,In_2840,In_1706);
nand U147 (N_147,In_238,In_134);
xnor U148 (N_148,In_475,In_930);
or U149 (N_149,In_2566,In_1690);
nand U150 (N_150,In_918,In_1337);
and U151 (N_151,In_2955,In_167);
nand U152 (N_152,In_1063,In_682);
and U153 (N_153,In_434,In_419);
nand U154 (N_154,In_1606,In_2936);
nor U155 (N_155,In_34,In_2452);
xnor U156 (N_156,In_2415,In_147);
nand U157 (N_157,In_2950,In_1257);
nor U158 (N_158,In_2064,In_699);
and U159 (N_159,In_287,In_1250);
or U160 (N_160,In_1014,In_1753);
nor U161 (N_161,In_283,In_2890);
and U162 (N_162,In_2191,In_2783);
nor U163 (N_163,In_840,In_186);
or U164 (N_164,In_1956,In_1092);
and U165 (N_165,In_1705,In_2919);
nand U166 (N_166,In_2811,In_2037);
nor U167 (N_167,In_53,In_912);
nand U168 (N_168,In_1151,In_1015);
xor U169 (N_169,In_2554,In_684);
or U170 (N_170,In_882,In_2323);
nand U171 (N_171,In_2403,In_2806);
or U172 (N_172,In_2856,In_2560);
nor U173 (N_173,In_1762,In_2058);
nand U174 (N_174,In_2937,In_1365);
nand U175 (N_175,In_708,In_1542);
nand U176 (N_176,In_1793,In_1343);
nor U177 (N_177,In_2008,In_2998);
nand U178 (N_178,In_1576,In_980);
or U179 (N_179,In_1535,In_317);
nand U180 (N_180,In_559,In_2838);
nor U181 (N_181,In_156,In_377);
or U182 (N_182,In_91,In_2208);
or U183 (N_183,In_2188,In_1485);
or U184 (N_184,In_2997,In_2755);
and U185 (N_185,In_2300,In_1533);
or U186 (N_186,In_1889,In_2313);
nor U187 (N_187,In_2846,In_137);
nand U188 (N_188,In_774,In_2619);
or U189 (N_189,In_1404,In_1782);
and U190 (N_190,In_1141,In_2500);
xor U191 (N_191,In_1938,In_474);
nor U192 (N_192,In_2294,In_2731);
nand U193 (N_193,In_2154,In_675);
and U194 (N_194,In_2982,In_1627);
and U195 (N_195,In_1010,In_1419);
nor U196 (N_196,In_1554,In_1734);
nor U197 (N_197,In_525,In_2580);
nor U198 (N_198,In_2388,In_1264);
or U199 (N_199,In_1733,In_1928);
xor U200 (N_200,In_2989,In_2895);
and U201 (N_201,In_1531,In_2182);
nor U202 (N_202,In_1949,In_796);
nor U203 (N_203,In_1483,In_1106);
nor U204 (N_204,In_2180,In_810);
nor U205 (N_205,In_1959,In_1196);
nand U206 (N_206,In_858,In_818);
and U207 (N_207,In_2005,In_2048);
nand U208 (N_208,In_927,In_1901);
and U209 (N_209,In_1841,In_2166);
and U210 (N_210,In_452,In_1973);
nand U211 (N_211,In_1480,In_499);
nor U212 (N_212,In_2854,In_760);
nand U213 (N_213,In_2760,In_483);
and U214 (N_214,In_2470,In_1368);
and U215 (N_215,In_2541,In_2237);
nor U216 (N_216,In_428,In_981);
or U217 (N_217,In_844,In_1549);
xnor U218 (N_218,In_1985,In_715);
nor U219 (N_219,In_297,In_2726);
nand U220 (N_220,In_1293,In_2645);
or U221 (N_221,In_2219,In_800);
or U222 (N_222,In_622,In_1006);
nor U223 (N_223,In_1479,In_268);
or U224 (N_224,In_496,In_1498);
nand U225 (N_225,In_994,In_223);
and U226 (N_226,In_1565,In_1148);
or U227 (N_227,In_2105,In_1152);
nand U228 (N_228,In_1963,In_1974);
or U229 (N_229,In_280,In_2128);
xor U230 (N_230,In_386,In_2851);
xor U231 (N_231,In_2983,In_451);
or U232 (N_232,In_649,In_757);
or U233 (N_233,In_1506,In_543);
nand U234 (N_234,In_1217,In_2471);
and U235 (N_235,In_2297,In_2098);
nand U236 (N_236,In_1222,In_1103);
and U237 (N_237,In_568,In_2900);
nor U238 (N_238,In_1742,In_2409);
nand U239 (N_239,In_688,In_1823);
nor U240 (N_240,In_769,In_583);
nand U241 (N_241,In_1131,In_1530);
or U242 (N_242,In_669,In_254);
or U243 (N_243,In_2824,In_2410);
and U244 (N_244,In_144,In_1086);
or U245 (N_245,In_2202,In_1173);
xor U246 (N_246,In_2697,In_1887);
or U247 (N_247,In_1227,In_64);
or U248 (N_248,In_37,In_278);
or U249 (N_249,In_1505,In_81);
nand U250 (N_250,In_158,In_2175);
or U251 (N_251,In_889,In_131);
nor U252 (N_252,In_2905,In_2086);
nor U253 (N_253,In_1089,In_2606);
or U254 (N_254,In_526,In_1435);
and U255 (N_255,In_676,In_512);
nand U256 (N_256,In_1512,In_1026);
or U257 (N_257,In_1698,In_2053);
nor U258 (N_258,In_696,In_887);
and U259 (N_259,In_1358,In_2852);
xor U260 (N_260,In_1401,In_50);
nand U261 (N_261,In_539,In_2421);
nor U262 (N_262,In_24,In_2626);
nor U263 (N_263,In_1588,In_1328);
or U264 (N_264,In_2296,In_1951);
and U265 (N_265,In_1033,In_2575);
xnor U266 (N_266,In_1517,In_2459);
nand U267 (N_267,In_542,In_1119);
nor U268 (N_268,In_2904,In_804);
and U269 (N_269,In_2302,In_1824);
and U270 (N_270,In_1153,In_2586);
nor U271 (N_271,In_770,In_891);
nand U272 (N_272,In_2163,In_1784);
nand U273 (N_273,In_876,In_1261);
or U274 (N_274,In_1248,In_193);
nand U275 (N_275,In_901,In_2797);
nor U276 (N_276,In_544,In_783);
nor U277 (N_277,In_2019,In_1797);
xor U278 (N_278,In_230,In_1085);
nand U279 (N_279,In_2280,In_445);
or U280 (N_280,In_1157,In_1656);
nand U281 (N_281,In_975,In_2348);
nand U282 (N_282,In_2206,In_1039);
and U283 (N_283,In_2903,In_420);
or U284 (N_284,In_799,In_555);
nor U285 (N_285,In_679,In_2009);
nor U286 (N_286,In_2172,In_2552);
xnor U287 (N_287,In_329,In_252);
and U288 (N_288,In_634,In_421);
nor U289 (N_289,In_2308,In_220);
and U290 (N_290,In_2864,In_1452);
nand U291 (N_291,In_1635,In_1658);
and U292 (N_292,In_339,In_17);
and U293 (N_293,In_2151,In_2437);
or U294 (N_294,In_58,In_1476);
nand U295 (N_295,In_811,In_877);
nor U296 (N_296,In_1743,In_2684);
and U297 (N_297,In_839,In_565);
xnor U298 (N_298,In_2822,In_447);
nand U299 (N_299,In_2957,In_664);
or U300 (N_300,In_1912,In_1256);
and U301 (N_301,In_2381,In_2129);
and U302 (N_302,In_2200,In_2284);
nand U303 (N_303,In_1968,In_249);
or U304 (N_304,In_2174,In_2203);
or U305 (N_305,In_183,In_1121);
nor U306 (N_306,In_841,In_1990);
nor U307 (N_307,In_2250,In_182);
nor U308 (N_308,In_2291,In_1335);
and U309 (N_309,In_2984,In_415);
nand U310 (N_310,In_1083,In_923);
or U311 (N_311,In_2255,In_2789);
and U312 (N_312,In_1670,In_291);
nand U313 (N_313,In_490,In_2321);
nor U314 (N_314,In_295,In_2494);
and U315 (N_315,In_2006,In_552);
nor U316 (N_316,In_1800,In_603);
and U317 (N_317,In_2272,In_574);
nand U318 (N_318,In_240,In_2959);
nor U319 (N_319,In_1109,In_1578);
nor U320 (N_320,In_1504,In_2269);
xnor U321 (N_321,In_244,In_2499);
or U322 (N_322,In_2573,In_2044);
or U323 (N_323,In_2295,In_2026);
or U324 (N_324,In_2326,In_1822);
nor U325 (N_325,In_166,In_2788);
and U326 (N_326,In_2392,In_2139);
nor U327 (N_327,In_1710,In_2609);
nand U328 (N_328,In_979,In_260);
nor U329 (N_329,In_1272,In_370);
nor U330 (N_330,In_524,In_264);
nand U331 (N_331,In_2109,In_1147);
nor U332 (N_332,In_305,In_1640);
or U333 (N_333,In_1631,In_2032);
xnor U334 (N_334,In_650,In_1870);
and U335 (N_335,In_2031,In_1225);
and U336 (N_336,In_1826,In_1867);
xor U337 (N_337,In_1373,In_1035);
xnor U338 (N_338,In_1502,In_1387);
or U339 (N_339,In_2072,In_919);
or U340 (N_340,In_680,In_1376);
nor U341 (N_341,In_2167,In_467);
xor U342 (N_342,In_1210,In_1838);
nor U343 (N_343,In_2477,In_2995);
or U344 (N_344,In_1247,In_1697);
and U345 (N_345,In_1538,In_594);
nor U346 (N_346,In_362,In_605);
xor U347 (N_347,In_2655,In_1843);
xnor U348 (N_348,In_1481,In_2455);
and U349 (N_349,In_2359,In_689);
xnor U350 (N_350,In_983,In_628);
nand U351 (N_351,In_564,In_1712);
and U352 (N_352,In_1484,In_2542);
or U353 (N_353,In_7,In_497);
or U354 (N_354,In_1624,In_2569);
nor U355 (N_355,In_107,In_2591);
nor U356 (N_356,In_259,In_2077);
nor U357 (N_357,In_1031,In_2357);
and U358 (N_358,In_2892,In_1296);
nor U359 (N_359,In_1120,In_1667);
and U360 (N_360,In_617,In_546);
or U361 (N_361,In_2374,In_2750);
nor U362 (N_362,In_590,In_1394);
and U363 (N_363,In_794,In_1643);
xor U364 (N_364,In_2450,In_1655);
and U365 (N_365,In_184,In_734);
xor U366 (N_366,In_2956,In_2971);
and U367 (N_367,In_621,In_212);
nand U368 (N_368,In_446,In_1647);
or U369 (N_369,In_2967,In_2217);
xnor U370 (N_370,In_2705,In_2717);
or U371 (N_371,In_338,In_1907);
and U372 (N_372,In_1313,In_1622);
or U373 (N_373,In_1439,In_206);
nor U374 (N_374,In_185,In_365);
nand U375 (N_375,In_2240,In_1216);
nor U376 (N_376,In_1433,In_2599);
or U377 (N_377,In_111,In_2727);
nand U378 (N_378,In_340,In_1837);
and U379 (N_379,In_2428,In_1470);
or U380 (N_380,In_397,In_203);
xor U381 (N_381,In_506,In_199);
xor U382 (N_382,In_1477,In_2022);
or U383 (N_383,In_1073,In_2987);
or U384 (N_384,In_830,In_2980);
and U385 (N_385,In_60,In_384);
nand U386 (N_386,In_1799,In_1679);
nand U387 (N_387,In_1379,In_2362);
nor U388 (N_388,In_875,In_407);
nor U389 (N_389,In_2685,In_1919);
nor U390 (N_390,In_2778,In_1308);
and U391 (N_391,In_481,In_541);
nor U392 (N_392,In_1999,In_2379);
and U393 (N_393,In_1828,In_1297);
nor U394 (N_394,In_2401,In_2615);
nand U395 (N_395,In_472,In_1819);
xor U396 (N_396,In_790,In_2387);
nor U397 (N_397,In_2425,In_1371);
and U398 (N_398,In_1787,In_155);
nor U399 (N_399,In_2299,In_1771);
and U400 (N_400,In_566,In_2741);
xnor U401 (N_401,In_2068,In_2040);
nand U402 (N_402,In_2325,In_1964);
nor U403 (N_403,In_1555,In_1118);
and U404 (N_404,In_1052,In_2310);
and U405 (N_405,In_2382,In_833);
and U406 (N_406,In_1113,In_2350);
and U407 (N_407,In_1792,In_1378);
nand U408 (N_408,In_356,In_578);
and U409 (N_409,In_1055,In_764);
or U410 (N_410,In_1314,In_2503);
and U411 (N_411,In_2636,In_1453);
and U412 (N_412,In_195,In_2650);
nor U413 (N_413,In_1298,In_707);
and U414 (N_414,In_1860,In_2176);
nor U415 (N_415,In_1050,In_2003);
nor U416 (N_416,In_1544,In_581);
or U417 (N_417,In_614,In_105);
and U418 (N_418,In_2536,In_2334);
and U419 (N_419,In_864,In_100);
or U420 (N_420,In_2873,In_801);
or U421 (N_421,In_1344,In_1429);
or U422 (N_422,In_2426,In_1240);
and U423 (N_423,In_371,In_328);
nor U424 (N_424,In_1030,In_275);
nand U425 (N_425,In_1906,In_2027);
or U426 (N_426,In_2074,In_1366);
and U427 (N_427,In_827,In_176);
nand U428 (N_428,In_1436,In_672);
xnor U429 (N_429,In_261,In_2143);
and U430 (N_430,In_2061,In_502);
nand U431 (N_431,In_1560,In_188);
nand U432 (N_432,In_1281,In_266);
xnor U433 (N_433,In_2423,In_1417);
and U434 (N_434,In_2918,In_2277);
and U435 (N_435,In_779,In_842);
and U436 (N_436,In_379,In_1577);
xnor U437 (N_437,In_2848,In_1503);
or U438 (N_438,In_2352,In_432);
nor U439 (N_439,In_1763,In_2162);
nor U440 (N_440,In_1236,In_847);
or U441 (N_441,In_1921,In_2458);
and U442 (N_442,In_1354,In_146);
nand U443 (N_443,In_1032,In_1023);
nor U444 (N_444,In_2947,In_1421);
and U445 (N_445,In_286,In_1123);
and U446 (N_446,In_947,In_1457);
and U447 (N_447,In_2101,In_1431);
or U448 (N_448,In_2669,In_995);
or U449 (N_449,In_217,In_99);
xor U450 (N_450,In_916,In_493);
or U451 (N_451,In_722,In_2290);
nor U452 (N_452,In_413,In_855);
and U453 (N_453,In_1356,In_1649);
xor U454 (N_454,In_2531,In_357);
and U455 (N_455,In_1888,In_540);
nand U456 (N_456,In_1700,In_1036);
and U457 (N_457,In_532,In_1197);
or U458 (N_458,In_1288,In_1972);
nand U459 (N_459,In_1853,In_87);
and U460 (N_460,In_2584,In_2589);
and U461 (N_461,In_1415,In_2059);
nor U462 (N_462,In_1223,In_2331);
nor U463 (N_463,In_996,In_1294);
or U464 (N_464,In_2914,In_2867);
xnor U465 (N_465,In_1184,In_2968);
and U466 (N_466,In_953,In_1442);
nand U467 (N_467,In_2429,In_767);
and U468 (N_468,In_1011,In_778);
nand U469 (N_469,In_1780,In_2468);
or U470 (N_470,In_2417,In_1866);
or U471 (N_471,In_298,In_2405);
nand U472 (N_472,In_1045,In_2570);
nor U473 (N_473,In_1129,In_1665);
nand U474 (N_474,In_1451,In_514);
nor U475 (N_475,In_1923,In_775);
nor U476 (N_476,In_2492,In_2389);
nand U477 (N_477,In_71,In_1246);
nor U478 (N_478,In_1007,In_2860);
xor U479 (N_479,In_4,In_709);
or U480 (N_480,In_314,In_300);
or U481 (N_481,In_443,In_2884);
and U482 (N_482,In_1520,In_1789);
nand U483 (N_483,In_869,In_161);
nor U484 (N_484,In_1454,In_97);
nor U485 (N_485,In_2205,In_2548);
xor U486 (N_486,In_1960,In_360);
and U487 (N_487,In_2878,In_977);
nor U488 (N_488,In_2365,In_1345);
nor U489 (N_489,In_984,In_548);
or U490 (N_490,In_1571,In_2135);
nor U491 (N_491,In_469,In_2600);
nand U492 (N_492,In_1384,In_1268);
nand U493 (N_493,In_1262,In_2235);
xor U494 (N_494,In_2782,In_2532);
nor U495 (N_495,In_348,In_1925);
xnor U496 (N_496,In_189,In_2204);
or U497 (N_497,In_1874,In_630);
nor U498 (N_498,In_2689,In_1913);
or U499 (N_499,In_332,In_1612);
nand U500 (N_500,In_1459,In_19);
nand U501 (N_501,In_886,In_935);
nand U502 (N_502,In_1899,In_2309);
nor U503 (N_503,In_1329,In_1332);
and U504 (N_504,In_1114,In_118);
nor U505 (N_505,In_2928,In_2275);
nor U506 (N_506,In_2946,In_655);
and U507 (N_507,In_638,In_1474);
or U508 (N_508,In_1607,In_2603);
nand U509 (N_509,In_950,In_1316);
nor U510 (N_510,In_2652,In_2681);
nor U511 (N_511,In_2226,In_1475);
nor U512 (N_512,In_1585,In_550);
and U513 (N_513,In_922,In_1170);
nor U514 (N_514,In_939,In_898);
nor U515 (N_515,In_1087,In_1970);
or U516 (N_516,In_1962,In_1871);
nand U517 (N_517,In_515,In_2665);
nor U518 (N_518,In_289,In_2328);
and U519 (N_519,In_2862,In_1955);
xnor U520 (N_520,In_385,In_142);
nor U521 (N_521,In_1034,In_2836);
nor U522 (N_522,In_1139,In_2396);
and U523 (N_523,In_1855,In_1251);
or U524 (N_524,In_245,In_2639);
nor U525 (N_525,In_2178,In_756);
nor U526 (N_526,In_1231,In_482);
or U527 (N_527,In_1463,In_501);
nor U528 (N_528,In_1993,In_538);
nand U529 (N_529,In_1500,In_1717);
nand U530 (N_530,In_366,In_1441);
and U531 (N_531,In_785,In_2610);
and U532 (N_532,In_1958,In_1781);
xor U533 (N_533,In_429,In_1933);
nand U534 (N_534,In_410,In_1673);
or U535 (N_535,In_1727,In_14);
nor U536 (N_536,In_2837,In_2385);
nand U537 (N_537,In_2253,In_2076);
nand U538 (N_538,In_42,In_2108);
or U539 (N_539,In_359,In_2899);
xor U540 (N_540,In_861,In_2324);
and U541 (N_541,In_72,In_417);
or U542 (N_542,In_1110,In_519);
or U543 (N_543,In_2342,In_798);
and U544 (N_544,In_1054,In_1563);
nor U545 (N_545,In_674,In_1760);
nor U546 (N_546,In_511,In_2736);
or U547 (N_547,In_55,In_293);
and U548 (N_548,In_1597,In_1428);
or U549 (N_549,In_851,In_1154);
or U550 (N_550,In_2742,In_2616);
or U551 (N_551,In_2049,In_1211);
nand U552 (N_552,In_1835,In_643);
xnor U553 (N_553,In_2268,In_2932);
or U554 (N_554,In_1004,In_2333);
and U555 (N_555,In_2539,In_1192);
xnor U556 (N_556,In_381,In_1965);
or U557 (N_557,In_573,In_313);
nand U558 (N_558,In_86,In_1230);
or U559 (N_559,In_1830,In_393);
and U560 (N_560,In_224,In_1586);
or U561 (N_561,In_1637,In_372);
and U562 (N_562,In_2758,In_2795);
nand U563 (N_563,In_1920,In_2948);
and U564 (N_564,In_1553,In_2769);
and U565 (N_565,In_2896,In_485);
nand U566 (N_566,In_267,In_598);
nor U567 (N_567,In_2430,In_1728);
nor U568 (N_568,In_619,In_1685);
xnor U569 (N_569,In_2451,In_2465);
or U570 (N_570,In_1886,In_2723);
nor U571 (N_571,In_934,In_1725);
nor U572 (N_572,In_1674,In_2413);
nor U573 (N_573,In_888,In_763);
or U574 (N_574,In_1957,In_2888);
or U575 (N_575,In_2843,In_685);
or U576 (N_576,In_1813,In_2454);
or U577 (N_577,In_929,In_2084);
and U578 (N_578,In_113,In_2360);
nor U579 (N_579,In_940,In_1981);
nand U580 (N_580,In_2537,In_2894);
or U581 (N_581,In_196,In_966);
xnor U582 (N_582,In_334,In_303);
or U583 (N_583,In_1300,In_2881);
nand U584 (N_584,In_2404,In_1097);
nand U585 (N_585,In_2319,In_2124);
nor U586 (N_586,In_2969,In_1596);
nor U587 (N_587,In_1449,In_2827);
nor U588 (N_588,In_1601,In_2483);
nor U589 (N_589,In_491,In_1363);
and U590 (N_590,In_2673,In_751);
nor U591 (N_591,In_1183,In_1306);
xnor U592 (N_592,In_2587,In_2201);
nor U593 (N_593,In_2161,In_116);
nor U594 (N_594,In_787,In_933);
and U595 (N_595,In_1012,In_1486);
and U596 (N_596,In_486,In_2785);
nand U597 (N_597,In_2559,In_1303);
or U598 (N_598,In_470,In_1896);
or U599 (N_599,In_1802,In_2629);
nand U600 (N_600,In_1024,In_227);
nand U601 (N_601,In_1935,In_1767);
nand U602 (N_602,In_620,In_2613);
nor U603 (N_603,In_1393,In_232);
or U604 (N_604,In_285,In_2744);
nand U605 (N_605,In_2522,In_2412);
nor U606 (N_606,In_2358,In_712);
xor U607 (N_607,In_1775,In_1759);
and U608 (N_608,In_345,In_1833);
nor U609 (N_609,In_2549,In_522);
and U610 (N_610,In_2393,In_745);
or U611 (N_611,In_2624,In_2236);
and U612 (N_612,In_480,In_636);
or U613 (N_613,In_102,In_1243);
and U614 (N_614,In_920,In_1164);
and U615 (N_615,In_2620,In_1046);
xnor U616 (N_616,In_312,In_2444);
and U617 (N_617,In_2186,In_1156);
nand U618 (N_618,In_2315,In_1668);
nor U619 (N_619,In_276,In_1515);
nor U620 (N_620,In_2485,In_1382);
or U621 (N_621,In_557,In_579);
nor U622 (N_622,In_2512,In_1095);
nor U623 (N_623,In_1747,In_711);
nand U624 (N_624,In_2653,In_1195);
nor U625 (N_625,In_938,In_1013);
and U626 (N_626,In_51,In_2146);
and U627 (N_627,In_468,In_2446);
nand U628 (N_628,In_462,In_1494);
or U629 (N_629,In_1692,In_351);
nand U630 (N_630,In_1460,In_2891);
nand U631 (N_631,In_1028,In_1450);
or U632 (N_632,In_907,In_1749);
or U633 (N_633,In_2356,In_2732);
nor U634 (N_634,In_2514,In_2519);
and U635 (N_635,In_1204,In_835);
and U636 (N_636,In_990,In_1471);
nor U637 (N_637,In_2677,In_946);
and U638 (N_638,In_2057,In_138);
or U639 (N_639,In_63,In_1158);
and U640 (N_640,In_444,In_1142);
or U641 (N_641,In_2593,In_1620);
nor U642 (N_642,In_2719,In_904);
nor U643 (N_643,In_2322,In_2292);
xor U644 (N_644,In_198,In_2780);
or U645 (N_645,In_2821,In_1037);
or U646 (N_646,In_2102,In_611);
nand U647 (N_647,In_755,In_1730);
nand U648 (N_648,In_1632,In_2212);
and U649 (N_649,In_2792,In_629);
nor U650 (N_650,In_575,In_1407);
nor U651 (N_651,In_1592,In_1064);
nor U652 (N_652,In_361,In_1790);
nand U653 (N_653,In_521,In_219);
nand U654 (N_654,In_2643,In_955);
nand U655 (N_655,In_1876,In_40);
or U656 (N_656,In_2754,In_2378);
or U657 (N_657,In_2097,In_2801);
or U658 (N_658,In_1971,In_1334);
and U659 (N_659,In_1409,In_145);
or U660 (N_660,In_507,In_1657);
nand U661 (N_661,In_2728,In_1581);
xnor U662 (N_662,In_26,In_2013);
xnor U663 (N_663,In_1932,In_1931);
nor U664 (N_664,In_460,In_2749);
nor U665 (N_665,In_1719,In_1750);
nor U666 (N_666,In_1798,In_2347);
nor U667 (N_667,In_773,In_2729);
nand U668 (N_668,In_225,In_1397);
or U669 (N_669,In_554,In_383);
nor U670 (N_670,In_461,In_2960);
nand U671 (N_671,In_1413,In_2210);
and U672 (N_672,In_737,In_2901);
and U673 (N_673,In_2524,In_2416);
and U674 (N_674,In_1339,In_659);
xor U675 (N_675,In_121,In_1310);
and U676 (N_676,In_2158,In_2515);
and U677 (N_677,In_937,In_1807);
or U678 (N_678,In_2341,In_2036);
nand U679 (N_679,In_344,In_1336);
xor U680 (N_680,In_2751,In_2419);
nor U681 (N_681,In_2533,In_404);
and U682 (N_682,In_2000,In_2411);
nor U683 (N_683,In_974,In_2383);
xnor U684 (N_684,In_2833,In_1547);
nor U685 (N_685,In_2380,In_2460);
nand U686 (N_686,In_2819,In_797);
and U687 (N_687,In_1722,In_2964);
nand U688 (N_688,In_1735,In_2259);
nor U689 (N_689,In_2695,In_1662);
and U690 (N_690,In_1856,In_2194);
and U691 (N_691,In_1519,In_399);
nand U692 (N_692,In_1861,In_2733);
or U693 (N_693,In_2305,In_2908);
nand U694 (N_694,In_1651,In_1385);
or U695 (N_695,In_2781,In_691);
or U696 (N_696,In_828,In_2551);
or U697 (N_697,In_819,In_831);
nand U698 (N_698,In_534,In_2474);
or U699 (N_699,In_1777,In_1130);
and U700 (N_700,In_2713,In_604);
or U701 (N_701,In_1369,In_1377);
xnor U702 (N_702,In_2002,In_457);
xor U703 (N_703,In_976,In_2709);
nand U704 (N_704,In_1309,In_2095);
or U705 (N_705,In_2055,In_177);
nand U706 (N_706,In_723,In_1292);
nand U707 (N_707,In_2975,In_323);
nand U708 (N_708,In_54,In_250);
or U709 (N_709,In_455,In_15);
nand U710 (N_710,In_1492,In_1564);
xor U711 (N_711,In_1402,In_353);
or U712 (N_712,In_233,In_1765);
nor U713 (N_713,In_239,In_1299);
nand U714 (N_714,In_637,In_2508);
and U715 (N_715,In_782,In_845);
or U716 (N_716,In_1628,In_120);
or U717 (N_717,In_1444,In_657);
nand U718 (N_718,In_1521,In_2670);
nand U719 (N_719,In_2630,In_805);
or U720 (N_720,In_881,In_125);
nand U721 (N_721,In_1020,In_2688);
or U722 (N_722,In_2637,In_187);
and U723 (N_723,In_1331,In_1930);
or U724 (N_724,In_989,In_47);
and U725 (N_725,In_1078,In_1137);
and U726 (N_726,In_695,In_2525);
or U727 (N_727,In_1022,In_2646);
nand U728 (N_728,In_1858,In_67);
nand U729 (N_729,In_1661,In_1274);
or U730 (N_730,In_41,In_2298);
nor U731 (N_731,In_704,In_2281);
or U732 (N_732,In_2001,In_1695);
nand U733 (N_733,In_477,In_324);
nand U734 (N_734,In_716,In_1491);
or U735 (N_735,In_2052,In_505);
or U736 (N_736,In_106,In_2776);
nor U737 (N_737,In_714,In_569);
and U738 (N_738,In_2794,In_2288);
xnor U739 (N_739,In_1832,In_2096);
or U740 (N_740,In_1572,In_1877);
nor U741 (N_741,In_2433,In_1621);
and U742 (N_742,In_1809,In_2747);
and U743 (N_743,In_739,In_2092);
or U744 (N_744,In_130,In_2830);
and U745 (N_745,In_1820,In_180);
nor U746 (N_746,In_1249,In_2361);
and U747 (N_747,In_2661,In_471);
or U748 (N_748,In_635,In_1788);
or U749 (N_749,In_2735,In_1279);
and U750 (N_750,In_45,In_1191);
nand U751 (N_751,In_2173,In_226);
or U752 (N_752,In_1583,In_913);
nand U753 (N_753,In_1283,In_616);
nor U754 (N_754,In_1370,In_2245);
xor U755 (N_755,In_2842,In_337);
and U756 (N_756,In_2118,In_2018);
nor U757 (N_757,In_2337,In_1104);
nor U758 (N_758,In_1570,In_2876);
xor U759 (N_759,In_162,In_758);
or U760 (N_760,In_1271,In_2951);
and U761 (N_761,In_171,In_2283);
nand U762 (N_762,In_1478,In_412);
or U763 (N_763,In_536,In_440);
nor U764 (N_764,In_84,In_2825);
or U765 (N_765,In_1466,In_148);
or U766 (N_766,In_2099,In_153);
nand U767 (N_767,In_846,In_2889);
nor U768 (N_768,In_2696,In_968);
or U769 (N_769,In_464,In_1594);
nor U770 (N_770,In_724,In_665);
nor U771 (N_771,In_1244,In_1125);
nand U772 (N_772,In_2224,In_1254);
nor U773 (N_773,In_197,In_1465);
nand U774 (N_774,In_2439,In_2622);
xnor U775 (N_775,In_1188,In_2016);
xor U776 (N_776,In_892,In_1526);
nor U777 (N_777,In_2574,In_1025);
nor U778 (N_778,In_932,In_2658);
nand U779 (N_779,In_671,In_1937);
nand U780 (N_780,In_2702,In_1469);
nor U781 (N_781,In_2193,In_834);
and U782 (N_782,In_258,In_742);
nand U783 (N_783,In_2715,In_1827);
or U784 (N_784,In_2011,In_1495);
nand U785 (N_785,In_9,In_1146);
or U786 (N_786,In_2518,In_1199);
nand U787 (N_787,In_1663,In_2568);
or U788 (N_788,In_23,In_1890);
xnor U789 (N_789,In_202,In_868);
xnor U790 (N_790,In_2121,In_2476);
xor U791 (N_791,In_1239,In_2138);
nor U792 (N_792,In_1115,In_2087);
nor U793 (N_793,In_1265,In_12);
and U794 (N_794,In_101,In_1686);
nor U795 (N_795,In_2577,In_2516);
nor U796 (N_796,In_2376,In_2056);
nand U797 (N_797,In_2966,In_2686);
and U798 (N_798,In_1528,In_1350);
nor U799 (N_799,In_1950,In_194);
nand U800 (N_800,In_27,In_2314);
nand U801 (N_801,In_2528,In_1282);
nor U802 (N_802,In_759,In_1065);
or U803 (N_803,In_270,In_1245);
nor U804 (N_804,In_164,In_1903);
nor U805 (N_805,In_478,In_2039);
nor U806 (N_806,In_400,In_1609);
nand U807 (N_807,In_2683,In_2625);
or U808 (N_808,In_2974,In_364);
or U809 (N_809,In_1111,In_1194);
xnor U810 (N_810,In_79,In_1464);
nor U811 (N_811,In_1587,In_1732);
nand U812 (N_812,In_1708,In_1785);
nand U813 (N_813,In_1851,In_2771);
xor U814 (N_814,In_1716,In_1221);
or U815 (N_815,In_2813,In_1829);
nand U816 (N_816,In_2676,In_1885);
and U817 (N_817,In_16,In_2231);
nand U818 (N_818,In_2481,In_1599);
and U819 (N_819,In_1729,In_609);
nor U820 (N_820,In_597,In_408);
xor U821 (N_821,In_1320,In_866);
nor U822 (N_822,In_2442,In_1341);
xnor U823 (N_823,In_596,In_1140);
nor U824 (N_824,In_175,In_1617);
nor U825 (N_825,In_2192,In_1333);
or U826 (N_826,In_1163,In_1133);
and U827 (N_827,In_988,In_157);
nor U828 (N_828,In_824,In_2145);
nor U829 (N_829,In_1641,In_1574);
nand U830 (N_830,In_1307,In_1911);
or U831 (N_831,In_2116,In_466);
or U832 (N_832,In_1718,In_644);
and U833 (N_833,In_311,In_1808);
and U834 (N_834,In_1389,In_1944);
nor U835 (N_835,In_853,In_1380);
and U836 (N_836,In_909,In_22);
nand U837 (N_837,In_1414,In_1233);
nor U838 (N_838,In_2844,In_961);
nor U839 (N_839,In_2103,In_750);
and U840 (N_840,In_1580,In_172);
or U841 (N_841,In_903,In_2351);
and U842 (N_842,In_1954,In_456);
nand U843 (N_843,In_1509,In_2693);
nand U844 (N_844,In_1212,In_265);
nand U845 (N_845,In_1066,In_80);
nor U846 (N_846,In_1437,In_368);
nand U847 (N_847,In_911,In_863);
or U848 (N_848,In_1740,In_917);
and U849 (N_849,In_1280,In_2510);
nor U850 (N_850,In_46,In_2007);
xnor U851 (N_851,In_1796,In_1410);
or U852 (N_852,In_2222,In_972);
and U853 (N_853,In_2120,In_1489);
nand U854 (N_854,In_1112,In_533);
or U855 (N_855,In_388,In_1258);
nand U856 (N_856,In_2491,In_702);
nand U857 (N_857,In_2527,In_2799);
nor U858 (N_858,In_2635,In_1902);
and U859 (N_859,In_473,In_1875);
nor U860 (N_860,In_2089,In_836);
nor U861 (N_861,In_2790,In_2526);
and U862 (N_862,In_986,In_281);
nor U863 (N_863,In_1751,In_562);
and U864 (N_864,In_1226,In_690);
nor U865 (N_865,In_1664,In_1132);
nand U866 (N_866,In_646,In_2535);
and U867 (N_867,In_2227,In_648);
xor U868 (N_868,In_1737,In_1934);
nand U869 (N_869,In_1573,In_1644);
nor U870 (N_870,In_44,In_1724);
nand U871 (N_871,In_640,In_2701);
nor U872 (N_872,In_817,In_1390);
nor U873 (N_873,In_2114,In_62);
nor U874 (N_874,In_1473,In_2196);
or U875 (N_875,In_1948,In_1398);
nor U876 (N_876,In_296,In_1219);
nand U877 (N_877,In_2663,In_2398);
or U878 (N_878,In_1458,In_1042);
nor U879 (N_879,In_1713,In_2373);
and U880 (N_880,In_1897,In_498);
xor U881 (N_881,In_508,In_2927);
nor U882 (N_882,In_1731,In_1150);
and U883 (N_883,In_205,In_2228);
xnor U884 (N_884,In_985,In_900);
nand U885 (N_885,In_2858,In_1468);
nor U886 (N_886,In_2490,In_2798);
nand U887 (N_887,In_2440,In_2372);
or U888 (N_888,In_424,In_310);
nor U889 (N_889,In_18,In_228);
nor U890 (N_890,In_1305,In_872);
xnor U891 (N_891,In_2093,In_1616);
nor U892 (N_892,In_2336,In_181);
and U893 (N_893,In_1694,In_1134);
nand U894 (N_894,In_1922,In_623);
or U895 (N_895,In_1324,In_2170);
nand U896 (N_896,In_2126,In_1325);
nand U897 (N_897,In_1352,In_28);
nand U898 (N_898,In_1057,In_129);
or U899 (N_899,In_1953,In_1318);
nand U900 (N_900,In_1579,In_1383);
and U901 (N_901,In_567,In_2125);
or U902 (N_902,In_78,In_510);
and U903 (N_903,In_141,In_2804);
and U904 (N_904,In_2276,In_1881);
or U905 (N_905,In_178,In_135);
and U906 (N_906,In_2447,In_595);
and U907 (N_907,In_765,In_2576);
or U908 (N_908,In_576,In_1768);
or U909 (N_909,In_32,In_2238);
nor U910 (N_910,In_92,In_1381);
or U911 (N_911,In_1070,In_2479);
nor U912 (N_912,In_1290,In_1374);
xnor U913 (N_913,In_367,In_1260);
nand U914 (N_914,In_825,In_2543);
nor U915 (N_915,In_2209,In_601);
nand U916 (N_916,In_1786,In_2165);
nor U917 (N_917,In_382,In_896);
nor U918 (N_918,In_479,In_651);
nand U919 (N_919,In_214,In_2945);
or U920 (N_920,In_49,In_2618);
nor U921 (N_921,In_719,In_2993);
or U922 (N_922,In_2069,In_1349);
nor U923 (N_923,In_1741,In_1255);
and U924 (N_924,In_237,In_290);
nor U925 (N_925,In_123,In_850);
nor U926 (N_926,In_1185,In_1081);
and U927 (N_927,In_1952,In_2505);
nor U928 (N_928,In_1049,In_654);
or U929 (N_929,In_2488,In_2082);
nor U930 (N_930,In_1047,In_438);
or U931 (N_931,In_1997,In_1671);
xor U932 (N_932,In_2081,In_414);
or U933 (N_933,In_2565,In_1003);
nand U934 (N_934,In_703,In_1061);
nand U935 (N_935,In_2023,In_2320);
or U936 (N_936,In_2710,In_2706);
nor U937 (N_937,In_1101,In_1745);
nand U938 (N_938,In_342,In_2594);
nand U939 (N_939,In_1600,In_2886);
nor U940 (N_940,In_517,In_1080);
nand U941 (N_941,In_2775,In_1016);
or U942 (N_942,In_2761,In_2976);
and U943 (N_943,In_1840,In_2088);
nand U944 (N_944,In_2249,In_520);
or U945 (N_945,In_1654,In_1406);
or U946 (N_946,In_2434,In_2796);
nor U947 (N_947,In_547,In_2762);
and U948 (N_948,In_2708,In_1682);
or U949 (N_949,In_150,In_746);
xnor U950 (N_950,In_1589,In_591);
xor U951 (N_951,In_2786,In_673);
nor U952 (N_952,In_2664,In_1908);
nand U953 (N_953,In_1987,In_89);
xor U954 (N_954,In_2262,In_1105);
nand U955 (N_955,In_93,In_2464);
nand U956 (N_956,In_683,In_2287);
nor U957 (N_957,In_2304,In_1100);
nand U958 (N_958,In_284,In_2920);
or U959 (N_959,In_553,In_2763);
or U960 (N_960,In_2286,In_743);
xor U961 (N_961,In_2930,In_1278);
or U962 (N_962,In_1646,In_2572);
or U963 (N_963,In_803,In_1986);
nor U964 (N_964,In_2181,In_2486);
or U965 (N_965,In_2988,In_2913);
and U966 (N_966,In_1626,In_1455);
or U967 (N_967,In_561,In_109);
nor U968 (N_968,In_2344,In_11);
nand U969 (N_969,In_77,In_885);
and U970 (N_970,In_3,In_2021);
nand U971 (N_971,In_2952,In_251);
or U972 (N_972,In_2847,In_2375);
nand U973 (N_973,In_2067,In_2660);
or U974 (N_974,In_68,In_2656);
and U975 (N_975,In_971,In_2711);
and U976 (N_976,In_2273,In_897);
and U977 (N_977,In_416,In_1311);
nor U978 (N_978,In_2441,In_2941);
or U979 (N_979,In_1947,In_2868);
and U980 (N_980,In_65,In_2547);
or U981 (N_981,In_2511,In_48);
nand U982 (N_982,In_2106,In_771);
nor U983 (N_983,In_1516,In_1088);
nand U984 (N_984,In_333,In_1831);
nor U985 (N_985,In_964,In_1426);
nor U986 (N_986,In_2766,In_165);
nor U987 (N_987,In_2634,In_1559);
nor U988 (N_988,In_380,In_2764);
and U989 (N_989,In_6,In_1077);
nor U990 (N_990,In_321,In_1127);
and U991 (N_991,In_870,In_2211);
and U992 (N_992,In_1270,In_2132);
or U993 (N_993,In_2631,In_1259);
or U994 (N_994,In_459,In_2017);
and U995 (N_995,In_854,In_1979);
nor U996 (N_996,In_88,In_1575);
and U997 (N_997,In_1914,In_2123);
or U998 (N_998,In_2065,In_2915);
nor U999 (N_999,In_967,In_112);
nor U1000 (N_1000,In_2534,In_1424);
or U1001 (N_1001,In_122,In_667);
and U1002 (N_1002,In_2232,In_2390);
or U1003 (N_1003,In_2595,In_1090);
nor U1004 (N_1004,In_425,In_2244);
and U1005 (N_1005,In_626,In_1203);
nand U1006 (N_1006,In_2935,In_1878);
nor U1007 (N_1007,In_500,In_1234);
xor U1008 (N_1008,In_29,In_492);
and U1009 (N_1009,In_396,In_1929);
nor U1010 (N_1010,In_2621,In_2902);
nand U1011 (N_1011,In_2107,In_647);
and U1012 (N_1012,In_1276,In_221);
nor U1013 (N_1013,In_822,In_2718);
xnor U1014 (N_1014,In_1044,In_728);
nand U1015 (N_1015,In_2054,In_586);
or U1016 (N_1016,In_426,In_1598);
nand U1017 (N_1017,In_2289,In_1396);
or U1018 (N_1018,In_1367,In_1346);
nor U1019 (N_1019,In_256,In_2911);
and U1020 (N_1020,In_2330,In_2859);
xnor U1021 (N_1021,In_2436,In_2150);
or U1022 (N_1022,In_2556,In_762);
and U1023 (N_1023,In_253,In_2184);
or U1024 (N_1024,In_2317,In_373);
nand U1025 (N_1025,In_2839,In_954);
or U1026 (N_1026,In_1079,In_2394);
nand U1027 (N_1027,In_1834,In_2834);
nor U1028 (N_1028,In_1675,In_316);
or U1029 (N_1029,In_1038,In_2869);
nand U1030 (N_1030,In_717,In_387);
xor U1031 (N_1031,In_2614,In_1317);
or U1032 (N_1032,In_1072,In_463);
and U1033 (N_1033,In_2703,In_958);
xor U1034 (N_1034,In_663,In_2448);
or U1035 (N_1035,In_2159,In_139);
xor U1036 (N_1036,In_369,In_1448);
or U1037 (N_1037,In_761,In_1507);
nor U1038 (N_1038,In_2746,In_1839);
nor U1039 (N_1039,In_727,In_2546);
nor U1040 (N_1040,In_793,In_2712);
xnor U1041 (N_1041,In_2704,In_2369);
or U1042 (N_1042,In_209,In_1416);
nand U1043 (N_1043,In_1360,In_257);
nand U1044 (N_1044,In_401,In_1359);
nand U1045 (N_1045,In_418,In_1074);
nand U1046 (N_1046,In_788,In_2866);
nor U1047 (N_1047,In_1446,In_56);
and U1048 (N_1048,In_2218,In_210);
and U1049 (N_1049,In_1982,In_1676);
nand U1050 (N_1050,In_661,In_218);
nand U1051 (N_1051,In_2994,In_612);
nand U1052 (N_1052,In_997,In_1269);
nand U1053 (N_1053,In_1869,In_422);
nand U1054 (N_1054,In_355,In_1857);
and U1055 (N_1055,In_1094,In_528);
and U1056 (N_1056,In_1847,In_211);
xnor U1057 (N_1057,In_2924,In_694);
and U1058 (N_1058,In_2327,In_2882);
and U1059 (N_1059,In_1224,In_2414);
nand U1060 (N_1060,In_959,In_1143);
and U1061 (N_1061,In_0,In_1704);
nor U1062 (N_1062,In_2605,In_2725);
nor U1063 (N_1063,In_1746,In_1171);
and U1064 (N_1064,In_874,In_1842);
nor U1065 (N_1065,In_2144,In_70);
nor U1066 (N_1066,In_600,In_732);
or U1067 (N_1067,In_1523,In_2692);
and U1068 (N_1068,In_375,In_883);
and U1069 (N_1069,In_2029,In_154);
or U1070 (N_1070,In_949,In_476);
or U1071 (N_1071,In_1900,In_2078);
nand U1072 (N_1072,In_741,In_1652);
nor U1073 (N_1073,In_867,In_2674);
and U1074 (N_1074,In_309,In_36);
and U1075 (N_1075,In_449,In_606);
nand U1076 (N_1076,In_766,In_1975);
and U1077 (N_1077,In_1639,In_2787);
nor U1078 (N_1078,In_736,In_2815);
nor U1079 (N_1079,In_1098,In_2641);
nand U1080 (N_1080,In_2501,In_1319);
and U1081 (N_1081,In_945,In_618);
or U1082 (N_1082,In_2517,In_2258);
and U1083 (N_1083,In_119,In_2737);
and U1084 (N_1084,In_733,In_1939);
nand U1085 (N_1085,In_2879,In_2133);
and U1086 (N_1086,In_1642,In_772);
and U1087 (N_1087,In_1434,In_1213);
xnor U1088 (N_1088,In_132,In_1522);
and U1089 (N_1089,In_2590,In_777);
xor U1090 (N_1090,In_411,In_962);
and U1091 (N_1091,In_143,In_235);
and U1092 (N_1092,In_2293,In_905);
xnor U1093 (N_1093,In_1539,In_589);
nor U1094 (N_1094,In_1513,In_1361);
or U1095 (N_1095,In_2949,In_1940);
nand U1096 (N_1096,In_2583,In_1779);
xor U1097 (N_1097,In_1005,In_2285);
and U1098 (N_1098,In_117,In_2070);
nand U1099 (N_1099,In_2368,In_963);
nand U1100 (N_1100,In_2774,In_1117);
xor U1101 (N_1101,In_2432,In_1610);
or U1102 (N_1102,In_1205,In_503);
or U1103 (N_1103,In_1427,In_1991);
nor U1104 (N_1104,In_1556,In_2608);
nand U1105 (N_1105,In_2349,In_2970);
or U1106 (N_1106,In_1175,In_246);
nor U1107 (N_1107,In_776,In_1180);
and U1108 (N_1108,In_2020,In_516);
nor U1109 (N_1109,In_435,In_625);
nor U1110 (N_1110,In_2248,In_2865);
or U1111 (N_1111,In_1043,In_2234);
nor U1112 (N_1112,In_2335,In_1669);
nand U1113 (N_1113,In_518,In_2079);
xnor U1114 (N_1114,In_2722,In_2466);
or U1115 (N_1115,In_1501,In_390);
and U1116 (N_1116,In_391,In_149);
nor U1117 (N_1117,In_1873,In_330);
and U1118 (N_1118,In_1241,In_2243);
and U1119 (N_1119,In_1720,In_2083);
or U1120 (N_1120,In_2147,In_2934);
or U1121 (N_1121,In_2247,In_350);
nand U1122 (N_1122,In_729,In_2164);
xor U1123 (N_1123,In_2812,In_319);
nand U1124 (N_1124,In_39,In_2831);
nand U1125 (N_1125,In_2877,In_786);
nand U1126 (N_1126,In_814,In_2467);
nand U1127 (N_1127,In_1764,In_2743);
nand U1128 (N_1128,In_2033,In_2402);
nor U1129 (N_1129,In_2802,In_2047);
xor U1130 (N_1130,In_871,In_1209);
or U1131 (N_1131,In_2475,In_1508);
nand U1132 (N_1132,In_812,In_1988);
nand U1133 (N_1133,In_1511,In_2779);
nand U1134 (N_1134,In_124,In_1613);
and U1135 (N_1135,In_1524,In_1966);
and U1136 (N_1136,In_2907,In_1136);
or U1137 (N_1137,In_952,In_363);
nor U1138 (N_1138,In_2898,In_639);
or U1139 (N_1139,In_2038,In_2922);
or U1140 (N_1140,In_1490,In_288);
or U1141 (N_1141,In_1493,In_1405);
or U1142 (N_1142,In_2716,In_1179);
and U1143 (N_1143,In_242,In_163);
and U1144 (N_1144,In_2168,In_2241);
nor U1145 (N_1145,In_2012,In_1541);
nor U1146 (N_1146,In_700,In_1977);
nor U1147 (N_1147,In_1275,In_2773);
nand U1148 (N_1148,In_1548,In_1910);
or U1149 (N_1149,In_1849,In_795);
nand U1150 (N_1150,In_1773,In_951);
or U1151 (N_1151,In_2978,In_2141);
nand U1152 (N_1152,In_1995,In_2965);
nand U1153 (N_1153,In_936,In_1347);
and U1154 (N_1154,In_2435,In_1412);
or U1155 (N_1155,In_731,In_698);
nor U1156 (N_1156,In_1978,In_1138);
nor U1157 (N_1157,In_453,In_1418);
or U1158 (N_1158,In_376,In_1228);
or U1159 (N_1159,In_928,In_1748);
nor U1160 (N_1160,In_1126,In_2504);
xnor U1161 (N_1161,In_1315,In_484);
or U1162 (N_1162,In_1945,In_823);
nor U1163 (N_1163,In_2585,In_152);
nand U1164 (N_1164,In_133,In_2596);
nor U1165 (N_1165,In_2130,In_1558);
and U1166 (N_1166,In_781,In_2938);
or U1167 (N_1167,In_2377,In_1357);
nand U1168 (N_1168,In_2909,In_2917);
nand U1169 (N_1169,In_910,In_1128);
nor U1170 (N_1170,In_2925,In_1021);
nor U1171 (N_1171,In_2592,In_1590);
or U1172 (N_1172,In_2582,In_1068);
nand U1173 (N_1173,In_1806,In_1561);
nor U1174 (N_1174,In_1056,In_2627);
xor U1175 (N_1175,In_1689,In_1814);
xnor U1176 (N_1176,In_1756,In_1983);
xor U1177 (N_1177,In_1009,In_753);
or U1178 (N_1178,In_1811,In_523);
nand U1179 (N_1179,In_2961,In_454);
and U1180 (N_1180,In_2563,In_273);
nand U1181 (N_1181,In_880,In_2513);
xnor U1182 (N_1182,In_115,In_1604);
nor U1183 (N_1183,In_128,In_489);
and U1184 (N_1184,In_1186,In_2939);
nor U1185 (N_1185,In_2571,In_2803);
nor U1186 (N_1186,In_494,In_1302);
nor U1187 (N_1187,In_656,In_2338);
nand U1188 (N_1188,In_2346,In_1917);
and U1189 (N_1189,In_1392,In_1291);
or U1190 (N_1190,In_666,In_277);
xor U1191 (N_1191,In_2418,In_791);
or U1192 (N_1192,In_1757,In_1946);
nor U1193 (N_1193,In_2042,In_1391);
and U1194 (N_1194,In_906,In_1884);
and U1195 (N_1195,In_1267,In_592);
nand U1196 (N_1196,In_1769,In_2332);
nor U1197 (N_1197,In_838,In_2808);
and U1198 (N_1198,In_90,In_1008);
or U1199 (N_1199,In_2122,In_1075);
nor U1200 (N_1200,In_2252,In_2678);
nand U1201 (N_1201,In_341,In_1984);
and U1202 (N_1202,In_1593,In_1629);
and U1203 (N_1203,In_2445,In_1058);
nand U1204 (N_1204,In_2991,In_2597);
nor U1205 (N_1205,In_1053,In_2691);
or U1206 (N_1206,In_2926,In_2312);
and U1207 (N_1207,In_1891,In_1660);
nand U1208 (N_1208,In_747,In_1726);
or U1209 (N_1209,In_987,In_1499);
xor U1210 (N_1210,In_1805,In_1172);
nand U1211 (N_1211,In_1634,In_1062);
or U1212 (N_1212,In_2791,In_2260);
nor U1213 (N_1213,In_423,In_495);
xnor U1214 (N_1214,In_2954,In_1169);
nand U1215 (N_1215,In_884,In_2301);
nand U1216 (N_1216,In_914,In_2910);
nand U1217 (N_1217,In_2111,In_2714);
nor U1218 (N_1218,In_1989,In_1608);
and U1219 (N_1219,In_1048,In_2999);
or U1220 (N_1220,In_179,In_563);
nand U1221 (N_1221,In_2489,In_336);
or U1222 (N_1222,In_915,In_1687);
nor U1223 (N_1223,In_1514,In_2113);
nand U1224 (N_1224,In_1752,In_1648);
and U1225 (N_1225,In_2035,In_2270);
or U1226 (N_1226,In_1321,In_437);
xor U1227 (N_1227,In_1623,In_2136);
and U1228 (N_1228,In_641,In_992);
nand U1229 (N_1229,In_1529,In_2251);
nand U1230 (N_1230,In_2818,In_1691);
and U1231 (N_1231,In_2724,In_2740);
nor U1232 (N_1232,In_821,In_2306);
or U1233 (N_1233,In_2721,In_1166);
nor U1234 (N_1234,In_1852,In_2225);
and U1235 (N_1235,In_2119,In_527);
xnor U1236 (N_1236,In_2100,In_1924);
and U1237 (N_1237,In_705,In_513);
nor U1238 (N_1238,In_2137,In_2195);
nor U1239 (N_1239,In_2187,In_43);
nand U1240 (N_1240,In_2264,In_813);
nor U1241 (N_1241,In_610,In_1916);
or U1242 (N_1242,In_271,In_114);
or U1243 (N_1243,In_2399,In_2343);
nand U1244 (N_1244,In_1482,In_110);
nand U1245 (N_1245,In_2558,In_2767);
nor U1246 (N_1246,In_2469,In_1263);
nor U1247 (N_1247,In_2828,In_2809);
or U1248 (N_1248,In_2642,In_1190);
or U1249 (N_1249,In_2921,In_1348);
nor U1250 (N_1250,In_326,In_2473);
or U1251 (N_1251,In_2363,In_2793);
xor U1252 (N_1252,In_1182,In_1848);
and U1253 (N_1253,In_2502,In_993);
or U1254 (N_1254,In_584,In_1527);
nor U1255 (N_1255,In_1772,In_2784);
nor U1256 (N_1256,In_160,In_448);
nor U1257 (N_1257,In_2682,In_2816);
xnor U1258 (N_1258,In_98,In_895);
or U1259 (N_1259,In_1803,In_1202);
and U1260 (N_1260,In_1546,In_1625);
nor U1261 (N_1261,In_926,In_2422);
and U1262 (N_1262,In_2506,In_1342);
nor U1263 (N_1263,In_243,In_1681);
nand U1264 (N_1264,In_2367,In_389);
xor U1265 (N_1265,In_1456,In_627);
nand U1266 (N_1266,In_192,In_1159);
and U1267 (N_1267,In_2707,In_190);
or U1268 (N_1268,In_1364,In_1178);
and U1269 (N_1269,In_2607,In_2579);
nor U1270 (N_1270,In_1155,In_1567);
nor U1271 (N_1271,In_2183,In_1976);
or U1272 (N_1272,In_2274,In_1967);
xor U1273 (N_1273,In_662,In_802);
nor U1274 (N_1274,In_2529,In_1699);
and U1275 (N_1275,In_2142,In_504);
nor U1276 (N_1276,In_349,In_306);
or U1277 (N_1277,In_1569,In_2197);
and U1278 (N_1278,In_2153,In_2213);
nand U1279 (N_1279,In_2449,In_2687);
nand U1280 (N_1280,In_931,In_2777);
nor U1281 (N_1281,In_1996,In_615);
xor U1282 (N_1282,In_2817,In_1189);
and U1283 (N_1283,In_1059,In_2160);
nor U1284 (N_1284,In_1865,In_2045);
xnor U1285 (N_1285,In_304,In_2863);
nor U1286 (N_1286,In_2318,In_1534);
nor U1287 (N_1287,In_1702,In_551);
nand U1288 (N_1288,In_25,In_1201);
and U1289 (N_1289,In_30,In_10);
nand U1290 (N_1290,In_2198,In_678);
nor U1291 (N_1291,In_2257,In_1425);
nor U1292 (N_1292,In_1181,In_2672);
nand U1293 (N_1293,In_1229,In_136);
nor U1294 (N_1294,In_1266,In_2051);
or U1295 (N_1295,In_530,In_1362);
nor U1296 (N_1296,In_2094,In_127);
nor U1297 (N_1297,In_1353,In_52);
nand U1298 (N_1298,In_1825,In_509);
nand U1299 (N_1299,In_1605,In_82);
or U1300 (N_1300,In_2043,In_103);
or U1301 (N_1301,In_2845,In_2671);
and U1302 (N_1302,In_1289,In_1602);
nand U1303 (N_1303,In_1817,In_1591);
and U1304 (N_1304,In_374,In_908);
nand U1305 (N_1305,In_1711,In_1091);
nor U1306 (N_1306,In_607,In_1754);
nor U1307 (N_1307,In_151,In_1566);
and U1308 (N_1308,In_2617,In_2700);
and U1309 (N_1309,In_1135,In_1076);
nand U1310 (N_1310,In_2567,In_754);
nand U1311 (N_1311,In_2972,In_1);
nand U1312 (N_1312,In_2254,In_1678);
and U1313 (N_1313,In_1863,In_1859);
nor U1314 (N_1314,In_2177,In_2463);
and U1315 (N_1315,In_2371,In_1659);
nor U1316 (N_1316,In_725,In_2849);
and U1317 (N_1317,In_2647,In_1680);
and U1318 (N_1318,In_2134,In_608);
and U1319 (N_1319,In_670,In_1001);
or U1320 (N_1320,In_925,In_1168);
and U1321 (N_1321,In_2493,In_1447);
nor U1322 (N_1322,In_2112,In_1715);
or U1323 (N_1323,In_582,In_343);
or U1324 (N_1324,In_1904,In_738);
or U1325 (N_1325,In_2265,In_1411);
nand U1326 (N_1326,In_315,In_2855);
nor U1327 (N_1327,In_1755,In_2770);
or U1328 (N_1328,In_2752,In_686);
and U1329 (N_1329,In_2611,In_347);
nand U1330 (N_1330,In_208,In_832);
and U1331 (N_1331,In_255,In_1040);
or U1332 (N_1332,In_1707,In_1738);
xnor U1333 (N_1333,In_2654,In_1794);
xnor U1334 (N_1334,In_207,In_2073);
and U1335 (N_1335,In_73,In_2659);
xnor U1336 (N_1336,In_735,In_2562);
nand U1337 (N_1337,In_1029,In_2025);
xor U1338 (N_1338,In_2015,In_2992);
and U1339 (N_1339,In_1703,In_2553);
nor U1340 (N_1340,In_1287,In_262);
and U1341 (N_1341,In_2117,In_857);
nor U1342 (N_1342,In_2156,In_789);
nand U1343 (N_1343,In_301,In_2835);
nand U1344 (N_1344,In_1943,In_200);
xor U1345 (N_1345,In_660,In_856);
nor U1346 (N_1346,In_487,In_2638);
and U1347 (N_1347,In_633,In_2498);
or U1348 (N_1348,In_1532,In_1892);
nor U1349 (N_1349,In_1497,In_730);
and U1350 (N_1350,In_1562,In_229);
or U1351 (N_1351,In_2906,In_1774);
and U1352 (N_1352,In_571,In_1918);
nor U1353 (N_1353,In_2386,In_894);
nand U1354 (N_1354,In_2233,In_1545);
or U1355 (N_1355,In_2805,In_2267);
nand U1356 (N_1356,In_69,In_1375);
or U1357 (N_1357,In_1330,In_96);
or U1358 (N_1358,In_2157,In_1443);
nor U1359 (N_1359,In_2545,In_1472);
nand U1360 (N_1360,In_710,In_191);
or U1361 (N_1361,In_1167,In_2823);
nor U1362 (N_1362,In_2339,In_2140);
nand U1363 (N_1363,In_1096,In_2242);
nand U1364 (N_1364,In_2944,In_2207);
and U1365 (N_1365,In_1778,In_1812);
nor U1366 (N_1366,In_924,In_1206);
nor U1367 (N_1367,In_585,In_2973);
nor U1368 (N_1368,In_2990,In_2004);
nor U1369 (N_1369,In_2256,In_991);
and U1370 (N_1370,In_556,In_2085);
nor U1371 (N_1371,In_2216,In_1557);
nor U1372 (N_1372,In_302,In_1684);
and U1373 (N_1373,In_572,In_1543);
and U1374 (N_1374,In_2623,In_1235);
nand U1375 (N_1375,In_204,In_599);
nor U1376 (N_1376,In_294,In_2757);
and U1377 (N_1377,In_560,In_222);
nor U1378 (N_1378,In_681,In_1969);
nand U1379 (N_1379,In_269,In_837);
nand U1380 (N_1380,In_2075,In_2155);
or U1381 (N_1381,In_2169,In_580);
and U1382 (N_1382,In_1237,In_1525);
nand U1383 (N_1383,In_465,In_1744);
and U1384 (N_1384,In_2266,In_2807);
xor U1385 (N_1385,In_879,In_1653);
nor U1386 (N_1386,In_2340,In_2189);
or U1387 (N_1387,In_263,In_809);
and U1388 (N_1388,In_215,In_1568);
and U1389 (N_1389,In_1980,In_2060);
and U1390 (N_1390,In_893,In_2271);
nand U1391 (N_1391,In_1804,In_1636);
or U1392 (N_1392,In_170,In_1666);
nor U1393 (N_1393,In_613,In_1487);
nand U1394 (N_1394,In_2730,In_320);
or U1395 (N_1395,In_2239,In_1766);
xnor U1396 (N_1396,In_2229,In_1161);
and U1397 (N_1397,In_1723,In_1423);
nand U1398 (N_1398,In_231,In_948);
nor U1399 (N_1399,In_2826,In_2311);
nand U1400 (N_1400,In_66,In_1611);
nor U1401 (N_1401,In_2810,In_1215);
nand U1402 (N_1402,In_2407,In_2104);
nor U1403 (N_1403,In_2010,In_1432);
and U1404 (N_1404,In_247,In_849);
nand U1405 (N_1405,In_201,In_2604);
nand U1406 (N_1406,In_720,In_2220);
and U1407 (N_1407,In_2581,In_1714);
nand U1408 (N_1408,In_1880,In_140);
and U1409 (N_1409,In_2649,In_1927);
or U1410 (N_1410,In_31,In_403);
or U1411 (N_1411,In_1295,In_1618);
nand U1412 (N_1412,In_631,In_2391);
nor U1413 (N_1413,In_899,In_2127);
and U1414 (N_1414,In_1721,In_2680);
xnor U1415 (N_1415,In_282,In_1836);
nand U1416 (N_1416,In_1818,In_274);
nor U1417 (N_1417,In_1552,In_1277);
nand U1418 (N_1418,In_2885,In_1926);
and U1419 (N_1419,In_308,In_1304);
and U1420 (N_1420,In_2171,In_2110);
or U1421 (N_1421,In_83,In_2400);
nor U1422 (N_1422,In_2768,In_442);
nor U1423 (N_1423,In_740,In_2024);
nand U1424 (N_1424,In_2530,In_2745);
and U1425 (N_1425,In_33,In_2030);
xor U1426 (N_1426,In_1683,In_873);
or U1427 (N_1427,In_2066,In_2872);
nor U1428 (N_1428,In_2657,In_1894);
or U1429 (N_1429,In_1816,In_652);
and U1430 (N_1430,In_2667,In_1000);
nor U1431 (N_1431,In_859,In_973);
nand U1432 (N_1432,In_1551,In_234);
nor U1433 (N_1433,In_816,In_2221);
nor U1434 (N_1434,In_2557,In_1220);
and U1435 (N_1435,In_2406,In_721);
xnor U1436 (N_1436,In_2438,In_2963);
xor U1437 (N_1437,In_1783,In_2353);
nor U1438 (N_1438,In_978,In_843);
nor U1439 (N_1439,In_2261,In_1630);
or U1440 (N_1440,In_61,In_1845);
nor U1441 (N_1441,In_535,In_1709);
and U1442 (N_1442,In_807,In_1116);
xnor U1443 (N_1443,In_1510,In_768);
and U1444 (N_1444,In_436,In_2408);
nand U1445 (N_1445,In_2668,In_2);
or U1446 (N_1446,In_439,In_1082);
nor U1447 (N_1447,In_2329,In_1177);
nand U1448 (N_1448,In_2420,In_749);
nand U1449 (N_1449,In_406,In_2487);
nor U1450 (N_1450,In_430,In_1338);
nor U1451 (N_1451,In_358,In_2063);
nand U1452 (N_1452,In_2366,In_1994);
or U1453 (N_1453,In_2509,In_2883);
nand U1454 (N_1454,In_693,In_2246);
or U1455 (N_1455,In_848,In_1027);
nor U1456 (N_1456,In_697,In_1445);
nand U1457 (N_1457,In_537,In_395);
and U1458 (N_1458,In_748,In_1122);
xnor U1459 (N_1459,In_174,In_1176);
and U1460 (N_1460,In_1496,In_2496);
nand U1461 (N_1461,In_2748,In_2738);
xor U1462 (N_1462,In_327,In_1340);
and U1463 (N_1463,In_2461,In_2482);
xor U1464 (N_1464,In_322,In_292);
or U1465 (N_1465,In_1537,In_1285);
nand U1466 (N_1466,In_2981,In_726);
nor U1467 (N_1467,In_59,In_1461);
and U1468 (N_1468,In_85,In_1961);
nand U1469 (N_1469,In_645,In_1614);
xnor U1470 (N_1470,In_624,In_1232);
xor U1471 (N_1471,In_588,In_2880);
xor U1472 (N_1472,In_38,In_2185);
xor U1473 (N_1473,In_1286,In_1488);
nor U1474 (N_1474,In_95,In_1758);
nand U1475 (N_1475,In_2028,In_1693);
or U1476 (N_1476,In_2395,In_2648);
nand U1477 (N_1477,In_75,In_346);
and U1478 (N_1478,In_2148,In_1584);
nor U1479 (N_1479,In_378,In_272);
or U1480 (N_1480,In_2307,In_2561);
nand U1481 (N_1481,In_2223,In_335);
xor U1482 (N_1482,In_593,In_2080);
nor U1483 (N_1483,In_2640,In_1701);
and U1484 (N_1484,In_2462,In_1850);
or U1485 (N_1485,In_2694,In_1645);
nor U1486 (N_1486,In_2457,In_701);
nor U1487 (N_1487,In_2598,In_780);
nand U1488 (N_1488,In_706,In_352);
or U1489 (N_1489,In_2214,In_752);
and U1490 (N_1490,In_2916,In_2279);
nand U1491 (N_1491,In_2602,In_960);
nor U1492 (N_1492,In_1615,In_806);
and U1493 (N_1493,In_2152,In_944);
and U1494 (N_1494,In_1540,In_2041);
nor U1495 (N_1495,In_402,In_826);
and U1496 (N_1496,In_279,In_2354);
nor U1497 (N_1497,In_1242,In_2644);
and U1498 (N_1498,In_441,In_1193);
or U1499 (N_1499,In_1093,In_450);
nor U1500 (N_1500,In_1072,In_1179);
nand U1501 (N_1501,In_2276,In_2191);
nand U1502 (N_1502,In_2606,In_2851);
or U1503 (N_1503,In_2897,In_1285);
nand U1504 (N_1504,In_1098,In_525);
nand U1505 (N_1505,In_137,In_1893);
nor U1506 (N_1506,In_1198,In_1053);
or U1507 (N_1507,In_173,In_2321);
nor U1508 (N_1508,In_694,In_2446);
nor U1509 (N_1509,In_630,In_832);
and U1510 (N_1510,In_1904,In_1277);
and U1511 (N_1511,In_2073,In_2611);
xnor U1512 (N_1512,In_1705,In_1013);
or U1513 (N_1513,In_254,In_2229);
or U1514 (N_1514,In_1454,In_2542);
or U1515 (N_1515,In_535,In_2188);
nor U1516 (N_1516,In_2221,In_1077);
and U1517 (N_1517,In_1044,In_656);
nor U1518 (N_1518,In_776,In_2431);
and U1519 (N_1519,In_1046,In_2465);
or U1520 (N_1520,In_1478,In_1848);
nand U1521 (N_1521,In_1760,In_2768);
nand U1522 (N_1522,In_2736,In_787);
and U1523 (N_1523,In_2508,In_1663);
or U1524 (N_1524,In_261,In_2940);
nor U1525 (N_1525,In_987,In_673);
and U1526 (N_1526,In_102,In_1959);
nor U1527 (N_1527,In_2828,In_1897);
nor U1528 (N_1528,In_105,In_1437);
or U1529 (N_1529,In_2521,In_744);
or U1530 (N_1530,In_65,In_44);
or U1531 (N_1531,In_2772,In_2403);
nor U1532 (N_1532,In_800,In_600);
nand U1533 (N_1533,In_1085,In_2037);
and U1534 (N_1534,In_2135,In_1143);
nand U1535 (N_1535,In_2114,In_84);
and U1536 (N_1536,In_25,In_2070);
or U1537 (N_1537,In_988,In_1780);
and U1538 (N_1538,In_341,In_888);
nand U1539 (N_1539,In_1751,In_52);
or U1540 (N_1540,In_922,In_1965);
xnor U1541 (N_1541,In_639,In_999);
nor U1542 (N_1542,In_683,In_197);
nor U1543 (N_1543,In_2704,In_2219);
nand U1544 (N_1544,In_622,In_134);
or U1545 (N_1545,In_526,In_1204);
and U1546 (N_1546,In_1083,In_1884);
nand U1547 (N_1547,In_2828,In_2097);
nand U1548 (N_1548,In_1403,In_1372);
xnor U1549 (N_1549,In_2297,In_1958);
nor U1550 (N_1550,In_745,In_940);
and U1551 (N_1551,In_2304,In_1557);
xnor U1552 (N_1552,In_1728,In_1159);
xor U1553 (N_1553,In_1229,In_1754);
nand U1554 (N_1554,In_2425,In_979);
or U1555 (N_1555,In_120,In_1931);
nor U1556 (N_1556,In_1365,In_1165);
nand U1557 (N_1557,In_45,In_1192);
nor U1558 (N_1558,In_2382,In_2439);
xnor U1559 (N_1559,In_1325,In_822);
nand U1560 (N_1560,In_2134,In_1220);
nand U1561 (N_1561,In_1351,In_2277);
nand U1562 (N_1562,In_1793,In_1456);
or U1563 (N_1563,In_2770,In_887);
and U1564 (N_1564,In_1968,In_727);
and U1565 (N_1565,In_885,In_194);
xnor U1566 (N_1566,In_1139,In_1064);
nor U1567 (N_1567,In_596,In_1617);
or U1568 (N_1568,In_2386,In_2959);
and U1569 (N_1569,In_676,In_1934);
nor U1570 (N_1570,In_128,In_2304);
or U1571 (N_1571,In_7,In_2480);
nor U1572 (N_1572,In_1785,In_1003);
nor U1573 (N_1573,In_1381,In_538);
and U1574 (N_1574,In_384,In_1257);
and U1575 (N_1575,In_870,In_2912);
or U1576 (N_1576,In_2434,In_909);
nor U1577 (N_1577,In_423,In_598);
and U1578 (N_1578,In_1568,In_13);
xnor U1579 (N_1579,In_1794,In_2910);
or U1580 (N_1580,In_1128,In_1161);
or U1581 (N_1581,In_2716,In_2593);
and U1582 (N_1582,In_2201,In_1251);
and U1583 (N_1583,In_2028,In_2877);
or U1584 (N_1584,In_2356,In_1672);
and U1585 (N_1585,In_2018,In_2468);
nor U1586 (N_1586,In_2772,In_2505);
and U1587 (N_1587,In_1121,In_1669);
or U1588 (N_1588,In_1913,In_25);
and U1589 (N_1589,In_1510,In_182);
nor U1590 (N_1590,In_2810,In_2314);
or U1591 (N_1591,In_2053,In_2507);
or U1592 (N_1592,In_2179,In_608);
nand U1593 (N_1593,In_570,In_2922);
nand U1594 (N_1594,In_2657,In_1988);
or U1595 (N_1595,In_255,In_1622);
and U1596 (N_1596,In_281,In_2598);
and U1597 (N_1597,In_665,In_598);
or U1598 (N_1598,In_549,In_693);
nand U1599 (N_1599,In_2006,In_438);
nand U1600 (N_1600,In_2420,In_2648);
and U1601 (N_1601,In_1586,In_1258);
or U1602 (N_1602,In_1220,In_550);
or U1603 (N_1603,In_1570,In_777);
nor U1604 (N_1604,In_1474,In_2999);
nand U1605 (N_1605,In_871,In_2203);
xor U1606 (N_1606,In_2558,In_208);
and U1607 (N_1607,In_2689,In_2919);
nand U1608 (N_1608,In_291,In_2420);
or U1609 (N_1609,In_904,In_400);
or U1610 (N_1610,In_464,In_2933);
nand U1611 (N_1611,In_1305,In_1817);
nand U1612 (N_1612,In_1973,In_2712);
and U1613 (N_1613,In_2495,In_2140);
nor U1614 (N_1614,In_2048,In_1704);
nor U1615 (N_1615,In_1791,In_542);
nor U1616 (N_1616,In_204,In_1820);
xor U1617 (N_1617,In_671,In_855);
nand U1618 (N_1618,In_1736,In_2845);
or U1619 (N_1619,In_150,In_19);
nand U1620 (N_1620,In_1259,In_69);
or U1621 (N_1621,In_539,In_1818);
or U1622 (N_1622,In_2265,In_2173);
nor U1623 (N_1623,In_1224,In_1594);
nand U1624 (N_1624,In_340,In_189);
nor U1625 (N_1625,In_1292,In_1974);
and U1626 (N_1626,In_1896,In_2952);
or U1627 (N_1627,In_2074,In_1592);
nand U1628 (N_1628,In_1287,In_2520);
and U1629 (N_1629,In_69,In_356);
and U1630 (N_1630,In_1376,In_1392);
and U1631 (N_1631,In_1062,In_1851);
nand U1632 (N_1632,In_2648,In_1126);
and U1633 (N_1633,In_1545,In_1603);
and U1634 (N_1634,In_142,In_1501);
nand U1635 (N_1635,In_730,In_2480);
nor U1636 (N_1636,In_1129,In_2662);
nor U1637 (N_1637,In_2382,In_593);
nand U1638 (N_1638,In_217,In_2636);
nand U1639 (N_1639,In_1838,In_2857);
or U1640 (N_1640,In_43,In_81);
nor U1641 (N_1641,In_335,In_1308);
nand U1642 (N_1642,In_1533,In_2096);
nor U1643 (N_1643,In_567,In_287);
nand U1644 (N_1644,In_2619,In_1900);
xor U1645 (N_1645,In_2179,In_1372);
nor U1646 (N_1646,In_743,In_2833);
nor U1647 (N_1647,In_2891,In_1052);
or U1648 (N_1648,In_2246,In_814);
or U1649 (N_1649,In_2043,In_706);
or U1650 (N_1650,In_2263,In_2868);
or U1651 (N_1651,In_286,In_1047);
nor U1652 (N_1652,In_2544,In_2028);
or U1653 (N_1653,In_974,In_1249);
and U1654 (N_1654,In_763,In_764);
and U1655 (N_1655,In_417,In_475);
and U1656 (N_1656,In_2563,In_670);
and U1657 (N_1657,In_2787,In_2895);
nand U1658 (N_1658,In_1209,In_2998);
and U1659 (N_1659,In_1522,In_1418);
nand U1660 (N_1660,In_1918,In_947);
nor U1661 (N_1661,In_805,In_978);
nand U1662 (N_1662,In_1740,In_2006);
or U1663 (N_1663,In_2476,In_1956);
xnor U1664 (N_1664,In_742,In_1180);
nand U1665 (N_1665,In_2232,In_2362);
and U1666 (N_1666,In_2569,In_39);
nand U1667 (N_1667,In_1816,In_1331);
nand U1668 (N_1668,In_1525,In_2820);
or U1669 (N_1669,In_2433,In_704);
or U1670 (N_1670,In_2017,In_1229);
or U1671 (N_1671,In_1118,In_627);
and U1672 (N_1672,In_1584,In_1662);
nand U1673 (N_1673,In_2648,In_225);
nor U1674 (N_1674,In_1527,In_1055);
nor U1675 (N_1675,In_1656,In_976);
nor U1676 (N_1676,In_662,In_48);
xor U1677 (N_1677,In_2087,In_1946);
and U1678 (N_1678,In_963,In_2077);
nor U1679 (N_1679,In_1448,In_22);
nor U1680 (N_1680,In_2372,In_1758);
nor U1681 (N_1681,In_645,In_2338);
or U1682 (N_1682,In_1086,In_1561);
and U1683 (N_1683,In_1037,In_570);
nand U1684 (N_1684,In_1131,In_1828);
or U1685 (N_1685,In_1222,In_2798);
nand U1686 (N_1686,In_1475,In_364);
nand U1687 (N_1687,In_1168,In_2690);
nor U1688 (N_1688,In_1751,In_2449);
nand U1689 (N_1689,In_125,In_493);
xor U1690 (N_1690,In_1214,In_1623);
nand U1691 (N_1691,In_636,In_704);
or U1692 (N_1692,In_42,In_1609);
nand U1693 (N_1693,In_2067,In_2530);
or U1694 (N_1694,In_2983,In_2685);
or U1695 (N_1695,In_2133,In_486);
nand U1696 (N_1696,In_883,In_1570);
and U1697 (N_1697,In_460,In_1563);
and U1698 (N_1698,In_2120,In_1852);
nand U1699 (N_1699,In_2373,In_96);
nand U1700 (N_1700,In_1244,In_2241);
xor U1701 (N_1701,In_2121,In_265);
or U1702 (N_1702,In_1663,In_766);
xnor U1703 (N_1703,In_2515,In_2965);
and U1704 (N_1704,In_902,In_2965);
or U1705 (N_1705,In_489,In_2447);
nor U1706 (N_1706,In_2829,In_686);
and U1707 (N_1707,In_1315,In_127);
and U1708 (N_1708,In_187,In_2738);
nand U1709 (N_1709,In_2255,In_1004);
or U1710 (N_1710,In_1510,In_1951);
or U1711 (N_1711,In_1143,In_2091);
and U1712 (N_1712,In_400,In_1165);
nand U1713 (N_1713,In_1021,In_159);
or U1714 (N_1714,In_402,In_6);
nand U1715 (N_1715,In_2071,In_1872);
nor U1716 (N_1716,In_2986,In_2230);
nor U1717 (N_1717,In_2828,In_1155);
or U1718 (N_1718,In_2759,In_2559);
nor U1719 (N_1719,In_565,In_1534);
nand U1720 (N_1720,In_1044,In_2512);
nor U1721 (N_1721,In_1830,In_458);
nand U1722 (N_1722,In_37,In_966);
xor U1723 (N_1723,In_2298,In_911);
nand U1724 (N_1724,In_1021,In_2905);
or U1725 (N_1725,In_1655,In_599);
nor U1726 (N_1726,In_2203,In_310);
nand U1727 (N_1727,In_899,In_52);
and U1728 (N_1728,In_1761,In_1173);
and U1729 (N_1729,In_1721,In_2253);
nand U1730 (N_1730,In_283,In_1172);
and U1731 (N_1731,In_172,In_133);
xor U1732 (N_1732,In_137,In_2057);
nor U1733 (N_1733,In_88,In_2983);
and U1734 (N_1734,In_2415,In_1020);
xnor U1735 (N_1735,In_2631,In_2496);
nand U1736 (N_1736,In_168,In_592);
nor U1737 (N_1737,In_1744,In_2343);
nand U1738 (N_1738,In_1439,In_23);
nand U1739 (N_1739,In_1831,In_2828);
nor U1740 (N_1740,In_277,In_1059);
nand U1741 (N_1741,In_1926,In_175);
and U1742 (N_1742,In_1921,In_2001);
or U1743 (N_1743,In_34,In_2089);
xor U1744 (N_1744,In_2339,In_802);
or U1745 (N_1745,In_1154,In_1933);
nor U1746 (N_1746,In_726,In_297);
and U1747 (N_1747,In_1158,In_380);
or U1748 (N_1748,In_988,In_443);
nor U1749 (N_1749,In_625,In_2433);
nand U1750 (N_1750,In_1313,In_1903);
and U1751 (N_1751,In_42,In_2554);
or U1752 (N_1752,In_1008,In_2660);
nand U1753 (N_1753,In_2199,In_1078);
and U1754 (N_1754,In_2169,In_1356);
or U1755 (N_1755,In_1893,In_1703);
or U1756 (N_1756,In_248,In_1078);
and U1757 (N_1757,In_2624,In_1709);
nor U1758 (N_1758,In_565,In_1821);
nor U1759 (N_1759,In_1924,In_5);
or U1760 (N_1760,In_1847,In_1032);
and U1761 (N_1761,In_519,In_467);
or U1762 (N_1762,In_2589,In_1918);
nor U1763 (N_1763,In_1301,In_38);
xnor U1764 (N_1764,In_2472,In_1448);
nand U1765 (N_1765,In_2221,In_368);
or U1766 (N_1766,In_1676,In_1972);
nand U1767 (N_1767,In_1133,In_1537);
xnor U1768 (N_1768,In_2656,In_2267);
and U1769 (N_1769,In_1078,In_18);
or U1770 (N_1770,In_1237,In_1829);
nand U1771 (N_1771,In_2288,In_2565);
nor U1772 (N_1772,In_1575,In_1858);
nand U1773 (N_1773,In_1798,In_1874);
nand U1774 (N_1774,In_581,In_481);
nor U1775 (N_1775,In_2396,In_1234);
and U1776 (N_1776,In_2608,In_1119);
xor U1777 (N_1777,In_2443,In_1898);
or U1778 (N_1778,In_247,In_2644);
and U1779 (N_1779,In_118,In_61);
nor U1780 (N_1780,In_742,In_352);
nand U1781 (N_1781,In_8,In_1480);
xor U1782 (N_1782,In_2919,In_2765);
or U1783 (N_1783,In_2494,In_1405);
or U1784 (N_1784,In_141,In_2035);
or U1785 (N_1785,In_1278,In_1145);
and U1786 (N_1786,In_1734,In_2762);
nand U1787 (N_1787,In_1830,In_740);
nor U1788 (N_1788,In_1696,In_2848);
nand U1789 (N_1789,In_1524,In_173);
and U1790 (N_1790,In_287,In_2097);
xnor U1791 (N_1791,In_1967,In_2196);
xor U1792 (N_1792,In_1190,In_1868);
nand U1793 (N_1793,In_2304,In_2785);
nor U1794 (N_1794,In_2197,In_2611);
nor U1795 (N_1795,In_1311,In_1921);
nor U1796 (N_1796,In_1257,In_2357);
nor U1797 (N_1797,In_1308,In_1507);
nor U1798 (N_1798,In_2453,In_547);
or U1799 (N_1799,In_193,In_2032);
nand U1800 (N_1800,In_2856,In_5);
nor U1801 (N_1801,In_1664,In_1808);
or U1802 (N_1802,In_1084,In_2423);
nor U1803 (N_1803,In_1887,In_483);
nor U1804 (N_1804,In_2804,In_2450);
xnor U1805 (N_1805,In_831,In_1232);
nor U1806 (N_1806,In_951,In_2774);
nor U1807 (N_1807,In_1518,In_636);
or U1808 (N_1808,In_349,In_2536);
nand U1809 (N_1809,In_2690,In_1103);
nand U1810 (N_1810,In_973,In_1373);
and U1811 (N_1811,In_2227,In_2151);
nand U1812 (N_1812,In_2604,In_1037);
nor U1813 (N_1813,In_2498,In_2234);
or U1814 (N_1814,In_1167,In_155);
or U1815 (N_1815,In_686,In_1601);
nand U1816 (N_1816,In_1407,In_2285);
and U1817 (N_1817,In_1940,In_2237);
or U1818 (N_1818,In_899,In_1033);
or U1819 (N_1819,In_554,In_964);
nand U1820 (N_1820,In_1028,In_2576);
nor U1821 (N_1821,In_1517,In_1475);
and U1822 (N_1822,In_2113,In_1516);
nand U1823 (N_1823,In_273,In_618);
nor U1824 (N_1824,In_241,In_248);
xnor U1825 (N_1825,In_460,In_2249);
nand U1826 (N_1826,In_1748,In_191);
or U1827 (N_1827,In_660,In_1645);
xor U1828 (N_1828,In_432,In_2080);
xnor U1829 (N_1829,In_807,In_255);
nand U1830 (N_1830,In_1581,In_2475);
or U1831 (N_1831,In_2179,In_2806);
nor U1832 (N_1832,In_2585,In_1639);
xor U1833 (N_1833,In_260,In_1357);
nand U1834 (N_1834,In_2350,In_2450);
nor U1835 (N_1835,In_61,In_260);
and U1836 (N_1836,In_2092,In_2907);
nand U1837 (N_1837,In_2335,In_423);
xnor U1838 (N_1838,In_1119,In_965);
xnor U1839 (N_1839,In_2492,In_1140);
or U1840 (N_1840,In_1276,In_2764);
or U1841 (N_1841,In_627,In_1612);
nand U1842 (N_1842,In_1890,In_2322);
and U1843 (N_1843,In_680,In_1636);
and U1844 (N_1844,In_2693,In_2497);
nand U1845 (N_1845,In_418,In_2170);
xor U1846 (N_1846,In_2342,In_1663);
nand U1847 (N_1847,In_2732,In_2943);
nor U1848 (N_1848,In_1964,In_2543);
nor U1849 (N_1849,In_684,In_1406);
or U1850 (N_1850,In_816,In_1556);
nand U1851 (N_1851,In_2726,In_1630);
nand U1852 (N_1852,In_2288,In_2762);
nand U1853 (N_1853,In_764,In_2814);
and U1854 (N_1854,In_692,In_210);
or U1855 (N_1855,In_1114,In_1552);
nor U1856 (N_1856,In_2581,In_1115);
and U1857 (N_1857,In_2909,In_1235);
and U1858 (N_1858,In_325,In_2898);
and U1859 (N_1859,In_2926,In_2536);
xnor U1860 (N_1860,In_109,In_2324);
xor U1861 (N_1861,In_1535,In_957);
xor U1862 (N_1862,In_2720,In_1118);
xnor U1863 (N_1863,In_2630,In_1479);
or U1864 (N_1864,In_1734,In_1231);
nor U1865 (N_1865,In_1864,In_1539);
xor U1866 (N_1866,In_283,In_43);
or U1867 (N_1867,In_1423,In_1357);
and U1868 (N_1868,In_692,In_1331);
or U1869 (N_1869,In_837,In_658);
nor U1870 (N_1870,In_1009,In_1060);
and U1871 (N_1871,In_1318,In_1025);
xnor U1872 (N_1872,In_787,In_1324);
nand U1873 (N_1873,In_2451,In_1474);
nor U1874 (N_1874,In_1797,In_2507);
xor U1875 (N_1875,In_2705,In_348);
nand U1876 (N_1876,In_2562,In_2315);
or U1877 (N_1877,In_2205,In_493);
nand U1878 (N_1878,In_1737,In_1910);
and U1879 (N_1879,In_2355,In_1159);
nand U1880 (N_1880,In_26,In_537);
and U1881 (N_1881,In_215,In_838);
nor U1882 (N_1882,In_1383,In_2312);
nor U1883 (N_1883,In_186,In_2878);
nand U1884 (N_1884,In_1795,In_996);
nand U1885 (N_1885,In_2597,In_2057);
nand U1886 (N_1886,In_644,In_2192);
or U1887 (N_1887,In_1011,In_2401);
and U1888 (N_1888,In_1530,In_2295);
or U1889 (N_1889,In_2155,In_1823);
nor U1890 (N_1890,In_460,In_1300);
and U1891 (N_1891,In_930,In_1205);
and U1892 (N_1892,In_356,In_1367);
nand U1893 (N_1893,In_2871,In_738);
xnor U1894 (N_1894,In_1446,In_1433);
xnor U1895 (N_1895,In_1376,In_153);
and U1896 (N_1896,In_1712,In_99);
or U1897 (N_1897,In_1043,In_59);
nand U1898 (N_1898,In_2422,In_1027);
nand U1899 (N_1899,In_2747,In_2416);
nor U1900 (N_1900,In_413,In_175);
nand U1901 (N_1901,In_899,In_950);
xnor U1902 (N_1902,In_1559,In_74);
or U1903 (N_1903,In_1346,In_5);
nand U1904 (N_1904,In_2674,In_981);
and U1905 (N_1905,In_1754,In_298);
nand U1906 (N_1906,In_1354,In_2964);
or U1907 (N_1907,In_923,In_2222);
xor U1908 (N_1908,In_2262,In_2719);
nand U1909 (N_1909,In_2484,In_894);
and U1910 (N_1910,In_627,In_1035);
nand U1911 (N_1911,In_1188,In_571);
or U1912 (N_1912,In_2037,In_831);
nor U1913 (N_1913,In_203,In_706);
nand U1914 (N_1914,In_858,In_72);
nand U1915 (N_1915,In_2401,In_9);
or U1916 (N_1916,In_1631,In_2788);
nor U1917 (N_1917,In_40,In_571);
nand U1918 (N_1918,In_1119,In_1000);
xnor U1919 (N_1919,In_1922,In_2194);
nor U1920 (N_1920,In_970,In_1860);
or U1921 (N_1921,In_2511,In_2459);
xor U1922 (N_1922,In_2108,In_461);
or U1923 (N_1923,In_203,In_1665);
and U1924 (N_1924,In_503,In_1917);
or U1925 (N_1925,In_782,In_2769);
nor U1926 (N_1926,In_1178,In_2348);
and U1927 (N_1927,In_36,In_2421);
and U1928 (N_1928,In_762,In_1040);
xor U1929 (N_1929,In_1370,In_1037);
or U1930 (N_1930,In_14,In_948);
or U1931 (N_1931,In_2039,In_91);
nand U1932 (N_1932,In_1122,In_417);
nand U1933 (N_1933,In_2679,In_2078);
nor U1934 (N_1934,In_1433,In_200);
and U1935 (N_1935,In_1187,In_1755);
and U1936 (N_1936,In_784,In_1603);
and U1937 (N_1937,In_1532,In_2142);
nand U1938 (N_1938,In_1219,In_1623);
or U1939 (N_1939,In_2265,In_1820);
or U1940 (N_1940,In_2331,In_2001);
nand U1941 (N_1941,In_2663,In_549);
nor U1942 (N_1942,In_1632,In_523);
nor U1943 (N_1943,In_1420,In_2896);
nand U1944 (N_1944,In_322,In_1836);
or U1945 (N_1945,In_822,In_96);
nand U1946 (N_1946,In_2063,In_748);
or U1947 (N_1947,In_2878,In_1385);
xor U1948 (N_1948,In_478,In_2279);
or U1949 (N_1949,In_224,In_2839);
nand U1950 (N_1950,In_1734,In_2747);
nor U1951 (N_1951,In_515,In_66);
and U1952 (N_1952,In_1619,In_21);
nand U1953 (N_1953,In_2941,In_1079);
xnor U1954 (N_1954,In_1153,In_2584);
or U1955 (N_1955,In_2581,In_2153);
and U1956 (N_1956,In_445,In_1636);
and U1957 (N_1957,In_2010,In_1183);
nor U1958 (N_1958,In_2992,In_1366);
or U1959 (N_1959,In_1634,In_183);
or U1960 (N_1960,In_2959,In_2215);
nor U1961 (N_1961,In_740,In_1577);
nand U1962 (N_1962,In_1706,In_1496);
and U1963 (N_1963,In_2816,In_1190);
nand U1964 (N_1964,In_2683,In_2736);
nand U1965 (N_1965,In_1652,In_256);
and U1966 (N_1966,In_1671,In_1464);
nor U1967 (N_1967,In_226,In_124);
or U1968 (N_1968,In_2952,In_1994);
nand U1969 (N_1969,In_2021,In_108);
nand U1970 (N_1970,In_1843,In_1515);
nand U1971 (N_1971,In_1442,In_2544);
nand U1972 (N_1972,In_1041,In_2986);
nor U1973 (N_1973,In_1779,In_1061);
or U1974 (N_1974,In_1253,In_2214);
and U1975 (N_1975,In_77,In_2204);
or U1976 (N_1976,In_2606,In_167);
nand U1977 (N_1977,In_2686,In_2502);
or U1978 (N_1978,In_364,In_83);
nand U1979 (N_1979,In_1243,In_189);
nand U1980 (N_1980,In_671,In_737);
nand U1981 (N_1981,In_955,In_1648);
or U1982 (N_1982,In_1012,In_775);
nand U1983 (N_1983,In_2296,In_1454);
nand U1984 (N_1984,In_688,In_737);
nand U1985 (N_1985,In_486,In_1991);
or U1986 (N_1986,In_646,In_692);
and U1987 (N_1987,In_1793,In_56);
or U1988 (N_1988,In_1092,In_686);
nand U1989 (N_1989,In_842,In_2511);
and U1990 (N_1990,In_700,In_88);
xnor U1991 (N_1991,In_1204,In_768);
and U1992 (N_1992,In_92,In_1656);
nand U1993 (N_1993,In_1863,In_990);
and U1994 (N_1994,In_58,In_1891);
nor U1995 (N_1995,In_1521,In_141);
and U1996 (N_1996,In_2349,In_1423);
or U1997 (N_1997,In_895,In_1971);
and U1998 (N_1998,In_2041,In_2580);
and U1999 (N_1999,In_1494,In_2900);
or U2000 (N_2000,In_1711,In_2459);
xor U2001 (N_2001,In_2140,In_2680);
or U2002 (N_2002,In_1764,In_2175);
nor U2003 (N_2003,In_1397,In_1271);
nand U2004 (N_2004,In_1888,In_146);
and U2005 (N_2005,In_234,In_1495);
and U2006 (N_2006,In_2303,In_664);
nor U2007 (N_2007,In_1071,In_1027);
xor U2008 (N_2008,In_28,In_2149);
or U2009 (N_2009,In_2914,In_1120);
or U2010 (N_2010,In_817,In_414);
nor U2011 (N_2011,In_2183,In_681);
or U2012 (N_2012,In_709,In_843);
nand U2013 (N_2013,In_2246,In_713);
or U2014 (N_2014,In_192,In_1481);
xor U2015 (N_2015,In_312,In_2480);
or U2016 (N_2016,In_2463,In_2027);
and U2017 (N_2017,In_229,In_2537);
xor U2018 (N_2018,In_2203,In_2528);
xnor U2019 (N_2019,In_433,In_2193);
nor U2020 (N_2020,In_308,In_2890);
and U2021 (N_2021,In_450,In_2908);
and U2022 (N_2022,In_32,In_1187);
nor U2023 (N_2023,In_661,In_1796);
or U2024 (N_2024,In_242,In_1403);
or U2025 (N_2025,In_2589,In_195);
nand U2026 (N_2026,In_2615,In_2273);
xor U2027 (N_2027,In_2825,In_494);
nand U2028 (N_2028,In_2196,In_1736);
nand U2029 (N_2029,In_2811,In_872);
or U2030 (N_2030,In_971,In_2294);
and U2031 (N_2031,In_1493,In_112);
nor U2032 (N_2032,In_1043,In_2968);
or U2033 (N_2033,In_22,In_1843);
nor U2034 (N_2034,In_2564,In_1714);
xnor U2035 (N_2035,In_15,In_2824);
nand U2036 (N_2036,In_1095,In_376);
nand U2037 (N_2037,In_1099,In_2934);
xor U2038 (N_2038,In_1535,In_51);
and U2039 (N_2039,In_1820,In_2227);
xor U2040 (N_2040,In_2316,In_733);
nand U2041 (N_2041,In_2666,In_2342);
nand U2042 (N_2042,In_661,In_2199);
xnor U2043 (N_2043,In_216,In_2686);
or U2044 (N_2044,In_1795,In_2152);
and U2045 (N_2045,In_25,In_1054);
nor U2046 (N_2046,In_2806,In_1263);
xnor U2047 (N_2047,In_2881,In_2330);
or U2048 (N_2048,In_589,In_2133);
nor U2049 (N_2049,In_2268,In_2488);
or U2050 (N_2050,In_2828,In_1824);
or U2051 (N_2051,In_17,In_2822);
and U2052 (N_2052,In_1044,In_1306);
or U2053 (N_2053,In_2886,In_2214);
nor U2054 (N_2054,In_2476,In_1668);
or U2055 (N_2055,In_2960,In_2306);
nor U2056 (N_2056,In_1861,In_1815);
or U2057 (N_2057,In_1037,In_1832);
nand U2058 (N_2058,In_2526,In_1540);
or U2059 (N_2059,In_1604,In_200);
nand U2060 (N_2060,In_1634,In_302);
nor U2061 (N_2061,In_1675,In_933);
nor U2062 (N_2062,In_2399,In_1647);
nand U2063 (N_2063,In_206,In_1731);
nand U2064 (N_2064,In_2957,In_2530);
nand U2065 (N_2065,In_1119,In_95);
or U2066 (N_2066,In_486,In_823);
or U2067 (N_2067,In_1702,In_1200);
or U2068 (N_2068,In_2759,In_925);
nor U2069 (N_2069,In_1317,In_1767);
nand U2070 (N_2070,In_1918,In_2576);
nor U2071 (N_2071,In_1936,In_2795);
nor U2072 (N_2072,In_2134,In_2445);
and U2073 (N_2073,In_2042,In_2310);
xnor U2074 (N_2074,In_409,In_1208);
and U2075 (N_2075,In_2997,In_2498);
or U2076 (N_2076,In_2450,In_22);
and U2077 (N_2077,In_2161,In_2053);
or U2078 (N_2078,In_986,In_1711);
and U2079 (N_2079,In_2573,In_163);
nand U2080 (N_2080,In_789,In_732);
nor U2081 (N_2081,In_1945,In_135);
or U2082 (N_2082,In_2291,In_2058);
or U2083 (N_2083,In_314,In_821);
and U2084 (N_2084,In_715,In_1109);
and U2085 (N_2085,In_891,In_1894);
or U2086 (N_2086,In_992,In_777);
xor U2087 (N_2087,In_2374,In_2289);
and U2088 (N_2088,In_1727,In_1477);
nor U2089 (N_2089,In_1032,In_1678);
and U2090 (N_2090,In_43,In_568);
or U2091 (N_2091,In_1595,In_887);
nor U2092 (N_2092,In_2585,In_1633);
nand U2093 (N_2093,In_147,In_18);
nor U2094 (N_2094,In_2577,In_2432);
or U2095 (N_2095,In_162,In_1008);
and U2096 (N_2096,In_2180,In_1297);
xor U2097 (N_2097,In_384,In_913);
and U2098 (N_2098,In_1566,In_2559);
and U2099 (N_2099,In_2862,In_553);
or U2100 (N_2100,In_900,In_1958);
or U2101 (N_2101,In_334,In_747);
xor U2102 (N_2102,In_1085,In_1585);
and U2103 (N_2103,In_330,In_2061);
and U2104 (N_2104,In_1898,In_1146);
nand U2105 (N_2105,In_2336,In_2770);
and U2106 (N_2106,In_2167,In_623);
nor U2107 (N_2107,In_696,In_1260);
or U2108 (N_2108,In_2024,In_1785);
nor U2109 (N_2109,In_116,In_2205);
or U2110 (N_2110,In_2150,In_1748);
and U2111 (N_2111,In_190,In_94);
or U2112 (N_2112,In_2462,In_363);
nor U2113 (N_2113,In_165,In_2282);
or U2114 (N_2114,In_2260,In_1156);
nor U2115 (N_2115,In_2789,In_2573);
nor U2116 (N_2116,In_2747,In_2195);
and U2117 (N_2117,In_1242,In_384);
nand U2118 (N_2118,In_1144,In_2048);
nand U2119 (N_2119,In_2209,In_2639);
or U2120 (N_2120,In_2387,In_710);
or U2121 (N_2121,In_1089,In_2102);
or U2122 (N_2122,In_1645,In_1520);
xnor U2123 (N_2123,In_436,In_809);
nor U2124 (N_2124,In_474,In_2234);
nand U2125 (N_2125,In_2032,In_345);
nor U2126 (N_2126,In_334,In_2477);
nand U2127 (N_2127,In_1675,In_453);
nor U2128 (N_2128,In_2202,In_2792);
nand U2129 (N_2129,In_746,In_1700);
and U2130 (N_2130,In_236,In_2760);
and U2131 (N_2131,In_2826,In_763);
and U2132 (N_2132,In_419,In_2456);
nor U2133 (N_2133,In_2836,In_1233);
and U2134 (N_2134,In_2349,In_1358);
nor U2135 (N_2135,In_1555,In_1360);
nand U2136 (N_2136,In_2207,In_2747);
or U2137 (N_2137,In_2086,In_2308);
or U2138 (N_2138,In_479,In_2957);
nor U2139 (N_2139,In_398,In_1738);
xor U2140 (N_2140,In_1252,In_2435);
and U2141 (N_2141,In_902,In_1260);
nor U2142 (N_2142,In_935,In_247);
nor U2143 (N_2143,In_881,In_2806);
or U2144 (N_2144,In_1985,In_1242);
xor U2145 (N_2145,In_2260,In_2565);
xnor U2146 (N_2146,In_2604,In_2935);
nor U2147 (N_2147,In_2253,In_318);
xnor U2148 (N_2148,In_2927,In_1041);
nor U2149 (N_2149,In_2994,In_1656);
nor U2150 (N_2150,In_1653,In_1948);
and U2151 (N_2151,In_2744,In_511);
and U2152 (N_2152,In_489,In_573);
nor U2153 (N_2153,In_139,In_2161);
nand U2154 (N_2154,In_710,In_351);
nor U2155 (N_2155,In_2189,In_2072);
xnor U2156 (N_2156,In_781,In_38);
and U2157 (N_2157,In_616,In_858);
nand U2158 (N_2158,In_1499,In_2448);
nand U2159 (N_2159,In_354,In_1212);
and U2160 (N_2160,In_2154,In_2820);
and U2161 (N_2161,In_2218,In_2959);
and U2162 (N_2162,In_558,In_1393);
or U2163 (N_2163,In_399,In_174);
nand U2164 (N_2164,In_970,In_242);
and U2165 (N_2165,In_1252,In_910);
and U2166 (N_2166,In_1730,In_965);
and U2167 (N_2167,In_633,In_318);
or U2168 (N_2168,In_1317,In_1724);
or U2169 (N_2169,In_2465,In_797);
xor U2170 (N_2170,In_2629,In_829);
xnor U2171 (N_2171,In_2247,In_2454);
and U2172 (N_2172,In_1615,In_80);
and U2173 (N_2173,In_666,In_2906);
nor U2174 (N_2174,In_2057,In_370);
xor U2175 (N_2175,In_2377,In_1258);
and U2176 (N_2176,In_2827,In_2417);
and U2177 (N_2177,In_1688,In_2663);
nor U2178 (N_2178,In_1493,In_1163);
xnor U2179 (N_2179,In_2562,In_2706);
xor U2180 (N_2180,In_1464,In_1430);
nand U2181 (N_2181,In_1581,In_2918);
or U2182 (N_2182,In_1850,In_502);
or U2183 (N_2183,In_1050,In_2367);
nand U2184 (N_2184,In_2864,In_217);
and U2185 (N_2185,In_2725,In_152);
nand U2186 (N_2186,In_2338,In_1384);
xor U2187 (N_2187,In_2388,In_1267);
and U2188 (N_2188,In_2331,In_1291);
xor U2189 (N_2189,In_1151,In_1785);
nand U2190 (N_2190,In_1218,In_2814);
and U2191 (N_2191,In_394,In_1625);
and U2192 (N_2192,In_2459,In_829);
and U2193 (N_2193,In_2987,In_2636);
nor U2194 (N_2194,In_2284,In_2054);
nor U2195 (N_2195,In_1751,In_829);
nand U2196 (N_2196,In_2082,In_1745);
and U2197 (N_2197,In_2690,In_1073);
xor U2198 (N_2198,In_1168,In_1169);
nand U2199 (N_2199,In_2806,In_599);
nor U2200 (N_2200,In_1722,In_1864);
nor U2201 (N_2201,In_453,In_37);
and U2202 (N_2202,In_1040,In_418);
or U2203 (N_2203,In_949,In_1);
nor U2204 (N_2204,In_315,In_1550);
nand U2205 (N_2205,In_2167,In_266);
nand U2206 (N_2206,In_2354,In_2291);
and U2207 (N_2207,In_1560,In_2223);
nor U2208 (N_2208,In_1823,In_2499);
nor U2209 (N_2209,In_708,In_1285);
nand U2210 (N_2210,In_1998,In_176);
nand U2211 (N_2211,In_2638,In_1631);
nor U2212 (N_2212,In_1927,In_2838);
and U2213 (N_2213,In_548,In_1808);
nor U2214 (N_2214,In_2693,In_484);
nand U2215 (N_2215,In_1601,In_2525);
nand U2216 (N_2216,In_190,In_865);
or U2217 (N_2217,In_2610,In_1786);
nand U2218 (N_2218,In_241,In_105);
or U2219 (N_2219,In_787,In_1265);
nor U2220 (N_2220,In_209,In_1864);
or U2221 (N_2221,In_1437,In_2681);
nor U2222 (N_2222,In_2238,In_2539);
nor U2223 (N_2223,In_192,In_1150);
or U2224 (N_2224,In_2876,In_2313);
nand U2225 (N_2225,In_855,In_1959);
or U2226 (N_2226,In_2002,In_2544);
or U2227 (N_2227,In_1498,In_2774);
nand U2228 (N_2228,In_2972,In_877);
or U2229 (N_2229,In_2368,In_1511);
and U2230 (N_2230,In_2694,In_2477);
and U2231 (N_2231,In_2764,In_2829);
and U2232 (N_2232,In_1573,In_312);
nor U2233 (N_2233,In_1148,In_2748);
nand U2234 (N_2234,In_1679,In_1433);
and U2235 (N_2235,In_2015,In_277);
nand U2236 (N_2236,In_2787,In_2667);
and U2237 (N_2237,In_1255,In_676);
nand U2238 (N_2238,In_69,In_2850);
nand U2239 (N_2239,In_2522,In_770);
or U2240 (N_2240,In_468,In_1173);
nand U2241 (N_2241,In_1567,In_1892);
nand U2242 (N_2242,In_950,In_685);
nor U2243 (N_2243,In_2342,In_2366);
nand U2244 (N_2244,In_269,In_1061);
or U2245 (N_2245,In_2598,In_452);
and U2246 (N_2246,In_155,In_2321);
nand U2247 (N_2247,In_1252,In_230);
and U2248 (N_2248,In_596,In_94);
nand U2249 (N_2249,In_1007,In_438);
nor U2250 (N_2250,In_1038,In_1438);
xor U2251 (N_2251,In_1600,In_852);
nand U2252 (N_2252,In_763,In_2032);
nor U2253 (N_2253,In_100,In_2843);
or U2254 (N_2254,In_445,In_2785);
nand U2255 (N_2255,In_2696,In_2564);
or U2256 (N_2256,In_2275,In_2948);
and U2257 (N_2257,In_2892,In_2688);
and U2258 (N_2258,In_1130,In_2697);
nor U2259 (N_2259,In_2096,In_2010);
xor U2260 (N_2260,In_1840,In_1823);
and U2261 (N_2261,In_106,In_1448);
nor U2262 (N_2262,In_2150,In_1813);
or U2263 (N_2263,In_2141,In_1104);
and U2264 (N_2264,In_187,In_226);
nand U2265 (N_2265,In_1195,In_961);
nand U2266 (N_2266,In_1796,In_1181);
nor U2267 (N_2267,In_900,In_101);
nand U2268 (N_2268,In_417,In_957);
and U2269 (N_2269,In_518,In_303);
xor U2270 (N_2270,In_2251,In_101);
and U2271 (N_2271,In_512,In_233);
and U2272 (N_2272,In_2395,In_2932);
nor U2273 (N_2273,In_486,In_1548);
xnor U2274 (N_2274,In_565,In_2910);
and U2275 (N_2275,In_1127,In_1307);
nand U2276 (N_2276,In_552,In_2283);
nor U2277 (N_2277,In_1941,In_2872);
and U2278 (N_2278,In_1698,In_1971);
or U2279 (N_2279,In_2993,In_2330);
nor U2280 (N_2280,In_543,In_601);
or U2281 (N_2281,In_2279,In_461);
and U2282 (N_2282,In_2104,In_2436);
or U2283 (N_2283,In_2571,In_2579);
xor U2284 (N_2284,In_2852,In_1405);
nand U2285 (N_2285,In_2837,In_528);
or U2286 (N_2286,In_2452,In_1737);
nand U2287 (N_2287,In_357,In_461);
nor U2288 (N_2288,In_1473,In_318);
nand U2289 (N_2289,In_1545,In_59);
nand U2290 (N_2290,In_381,In_2194);
nor U2291 (N_2291,In_2431,In_925);
nand U2292 (N_2292,In_2729,In_2458);
or U2293 (N_2293,In_1096,In_986);
xnor U2294 (N_2294,In_2396,In_740);
nor U2295 (N_2295,In_2967,In_846);
xor U2296 (N_2296,In_278,In_472);
xnor U2297 (N_2297,In_2034,In_2448);
or U2298 (N_2298,In_84,In_268);
nor U2299 (N_2299,In_2213,In_1884);
and U2300 (N_2300,In_2387,In_2838);
nand U2301 (N_2301,In_912,In_570);
nand U2302 (N_2302,In_319,In_1215);
nand U2303 (N_2303,In_2702,In_783);
or U2304 (N_2304,In_542,In_562);
nand U2305 (N_2305,In_401,In_65);
or U2306 (N_2306,In_2656,In_2686);
nand U2307 (N_2307,In_1254,In_804);
xnor U2308 (N_2308,In_1099,In_768);
nand U2309 (N_2309,In_1700,In_2088);
and U2310 (N_2310,In_1769,In_587);
xnor U2311 (N_2311,In_2602,In_2683);
nor U2312 (N_2312,In_826,In_838);
nor U2313 (N_2313,In_569,In_2879);
or U2314 (N_2314,In_981,In_717);
nand U2315 (N_2315,In_147,In_461);
nor U2316 (N_2316,In_1618,In_1585);
nand U2317 (N_2317,In_247,In_1532);
and U2318 (N_2318,In_2452,In_496);
nand U2319 (N_2319,In_1372,In_1056);
nor U2320 (N_2320,In_2218,In_2128);
nor U2321 (N_2321,In_784,In_680);
and U2322 (N_2322,In_126,In_2930);
nand U2323 (N_2323,In_2897,In_2900);
or U2324 (N_2324,In_122,In_2951);
nor U2325 (N_2325,In_647,In_213);
or U2326 (N_2326,In_1982,In_611);
nand U2327 (N_2327,In_1874,In_2832);
nand U2328 (N_2328,In_1389,In_107);
nor U2329 (N_2329,In_378,In_152);
nor U2330 (N_2330,In_1501,In_1208);
nor U2331 (N_2331,In_2946,In_1084);
and U2332 (N_2332,In_1213,In_2312);
nor U2333 (N_2333,In_2104,In_1435);
nand U2334 (N_2334,In_2736,In_1480);
and U2335 (N_2335,In_1601,In_2657);
or U2336 (N_2336,In_1222,In_1240);
and U2337 (N_2337,In_86,In_793);
nor U2338 (N_2338,In_357,In_2480);
and U2339 (N_2339,In_2523,In_2227);
or U2340 (N_2340,In_352,In_211);
nand U2341 (N_2341,In_2124,In_1407);
xor U2342 (N_2342,In_1353,In_2624);
nand U2343 (N_2343,In_1740,In_1552);
nand U2344 (N_2344,In_905,In_1112);
or U2345 (N_2345,In_2715,In_1210);
xor U2346 (N_2346,In_1257,In_2943);
and U2347 (N_2347,In_1671,In_841);
or U2348 (N_2348,In_1658,In_1433);
nand U2349 (N_2349,In_213,In_2313);
nor U2350 (N_2350,In_2059,In_392);
and U2351 (N_2351,In_1242,In_1596);
nor U2352 (N_2352,In_1332,In_237);
nand U2353 (N_2353,In_2130,In_1937);
and U2354 (N_2354,In_1710,In_1354);
nor U2355 (N_2355,In_2658,In_768);
or U2356 (N_2356,In_1857,In_1385);
or U2357 (N_2357,In_359,In_763);
and U2358 (N_2358,In_565,In_1973);
nor U2359 (N_2359,In_1293,In_1521);
or U2360 (N_2360,In_1590,In_556);
or U2361 (N_2361,In_1071,In_1808);
nand U2362 (N_2362,In_1475,In_1618);
nand U2363 (N_2363,In_1939,In_2388);
nand U2364 (N_2364,In_2819,In_2161);
nand U2365 (N_2365,In_1564,In_2593);
nor U2366 (N_2366,In_362,In_2383);
nor U2367 (N_2367,In_105,In_1464);
xnor U2368 (N_2368,In_2939,In_411);
nand U2369 (N_2369,In_2992,In_1662);
or U2370 (N_2370,In_2578,In_1095);
or U2371 (N_2371,In_2920,In_2081);
nand U2372 (N_2372,In_519,In_2765);
nor U2373 (N_2373,In_2996,In_2653);
xnor U2374 (N_2374,In_2027,In_1204);
nor U2375 (N_2375,In_1632,In_2532);
and U2376 (N_2376,In_1929,In_2932);
nor U2377 (N_2377,In_131,In_2976);
and U2378 (N_2378,In_731,In_1595);
and U2379 (N_2379,In_210,In_1744);
nand U2380 (N_2380,In_377,In_2433);
nor U2381 (N_2381,In_1930,In_1859);
or U2382 (N_2382,In_341,In_1543);
nand U2383 (N_2383,In_1921,In_649);
nor U2384 (N_2384,In_1031,In_1781);
or U2385 (N_2385,In_2680,In_2085);
or U2386 (N_2386,In_1452,In_2590);
nor U2387 (N_2387,In_1016,In_1611);
or U2388 (N_2388,In_2388,In_1189);
nor U2389 (N_2389,In_1844,In_1100);
nand U2390 (N_2390,In_726,In_308);
or U2391 (N_2391,In_2035,In_2618);
or U2392 (N_2392,In_1150,In_1754);
nand U2393 (N_2393,In_1623,In_258);
nand U2394 (N_2394,In_807,In_474);
or U2395 (N_2395,In_1507,In_949);
nand U2396 (N_2396,In_2501,In_2441);
and U2397 (N_2397,In_1831,In_128);
and U2398 (N_2398,In_100,In_1209);
nand U2399 (N_2399,In_2098,In_893);
and U2400 (N_2400,In_450,In_1068);
xor U2401 (N_2401,In_2398,In_493);
or U2402 (N_2402,In_2055,In_2428);
nand U2403 (N_2403,In_2539,In_1298);
xnor U2404 (N_2404,In_773,In_1638);
and U2405 (N_2405,In_128,In_1823);
and U2406 (N_2406,In_1378,In_1058);
or U2407 (N_2407,In_1742,In_2356);
or U2408 (N_2408,In_2394,In_130);
and U2409 (N_2409,In_1039,In_1982);
or U2410 (N_2410,In_886,In_1409);
nand U2411 (N_2411,In_2791,In_878);
or U2412 (N_2412,In_1275,In_2469);
or U2413 (N_2413,In_2242,In_2647);
and U2414 (N_2414,In_1385,In_2329);
or U2415 (N_2415,In_2605,In_813);
xor U2416 (N_2416,In_1798,In_1796);
xor U2417 (N_2417,In_999,In_1093);
or U2418 (N_2418,In_139,In_2916);
or U2419 (N_2419,In_2062,In_1423);
and U2420 (N_2420,In_287,In_2754);
or U2421 (N_2421,In_1216,In_1936);
nor U2422 (N_2422,In_1086,In_2638);
nand U2423 (N_2423,In_1374,In_1792);
and U2424 (N_2424,In_1633,In_234);
xnor U2425 (N_2425,In_1613,In_914);
or U2426 (N_2426,In_2548,In_28);
and U2427 (N_2427,In_2054,In_1097);
and U2428 (N_2428,In_2579,In_279);
and U2429 (N_2429,In_669,In_2590);
or U2430 (N_2430,In_310,In_1671);
nor U2431 (N_2431,In_114,In_1971);
nor U2432 (N_2432,In_2908,In_1121);
nand U2433 (N_2433,In_2391,In_655);
and U2434 (N_2434,In_354,In_2632);
or U2435 (N_2435,In_2372,In_566);
and U2436 (N_2436,In_2217,In_1492);
nor U2437 (N_2437,In_2629,In_1276);
nand U2438 (N_2438,In_1568,In_1024);
or U2439 (N_2439,In_2057,In_925);
and U2440 (N_2440,In_1505,In_507);
xnor U2441 (N_2441,In_1509,In_1921);
nand U2442 (N_2442,In_2701,In_1765);
nand U2443 (N_2443,In_1144,In_1685);
and U2444 (N_2444,In_742,In_2281);
and U2445 (N_2445,In_375,In_2847);
nor U2446 (N_2446,In_2023,In_2336);
nand U2447 (N_2447,In_702,In_2706);
nand U2448 (N_2448,In_2577,In_2258);
or U2449 (N_2449,In_2422,In_2084);
and U2450 (N_2450,In_1168,In_1202);
or U2451 (N_2451,In_1641,In_2937);
nor U2452 (N_2452,In_2360,In_1950);
nor U2453 (N_2453,In_930,In_1395);
or U2454 (N_2454,In_687,In_2368);
or U2455 (N_2455,In_612,In_856);
and U2456 (N_2456,In_2000,In_2361);
or U2457 (N_2457,In_1025,In_2101);
and U2458 (N_2458,In_29,In_21);
nand U2459 (N_2459,In_958,In_1191);
nand U2460 (N_2460,In_2682,In_1799);
nand U2461 (N_2461,In_1889,In_2707);
nor U2462 (N_2462,In_2336,In_2923);
nor U2463 (N_2463,In_518,In_1046);
xnor U2464 (N_2464,In_2124,In_2686);
or U2465 (N_2465,In_1077,In_1349);
nand U2466 (N_2466,In_672,In_1986);
xnor U2467 (N_2467,In_954,In_2271);
nand U2468 (N_2468,In_818,In_1292);
nand U2469 (N_2469,In_260,In_1004);
and U2470 (N_2470,In_468,In_1369);
and U2471 (N_2471,In_706,In_2909);
nor U2472 (N_2472,In_491,In_2653);
and U2473 (N_2473,In_2283,In_1280);
and U2474 (N_2474,In_2760,In_1955);
or U2475 (N_2475,In_1996,In_1684);
and U2476 (N_2476,In_1909,In_690);
xnor U2477 (N_2477,In_2995,In_1546);
or U2478 (N_2478,In_373,In_336);
nand U2479 (N_2479,In_445,In_1618);
xnor U2480 (N_2480,In_2568,In_164);
nand U2481 (N_2481,In_2266,In_33);
or U2482 (N_2482,In_1615,In_2819);
nand U2483 (N_2483,In_814,In_367);
or U2484 (N_2484,In_788,In_1601);
nand U2485 (N_2485,In_1140,In_1442);
nand U2486 (N_2486,In_1736,In_768);
nand U2487 (N_2487,In_2177,In_1249);
xnor U2488 (N_2488,In_986,In_427);
nand U2489 (N_2489,In_156,In_1530);
nand U2490 (N_2490,In_2663,In_130);
or U2491 (N_2491,In_1324,In_1103);
or U2492 (N_2492,In_2378,In_1670);
nand U2493 (N_2493,In_1099,In_960);
or U2494 (N_2494,In_2717,In_2293);
nand U2495 (N_2495,In_1997,In_1761);
nand U2496 (N_2496,In_2023,In_736);
nor U2497 (N_2497,In_288,In_2987);
nand U2498 (N_2498,In_397,In_33);
or U2499 (N_2499,In_2021,In_1026);
xnor U2500 (N_2500,In_2811,In_88);
nand U2501 (N_2501,In_1612,In_874);
nor U2502 (N_2502,In_1875,In_2096);
nand U2503 (N_2503,In_2567,In_59);
xnor U2504 (N_2504,In_1324,In_366);
nor U2505 (N_2505,In_56,In_1532);
or U2506 (N_2506,In_2809,In_1163);
nor U2507 (N_2507,In_763,In_2020);
nand U2508 (N_2508,In_652,In_369);
nor U2509 (N_2509,In_1834,In_926);
xor U2510 (N_2510,In_2646,In_1249);
and U2511 (N_2511,In_849,In_1228);
or U2512 (N_2512,In_2117,In_2020);
or U2513 (N_2513,In_2796,In_2243);
nand U2514 (N_2514,In_120,In_794);
or U2515 (N_2515,In_1846,In_2281);
and U2516 (N_2516,In_371,In_1720);
and U2517 (N_2517,In_2145,In_1932);
nand U2518 (N_2518,In_2252,In_2296);
or U2519 (N_2519,In_1768,In_500);
xnor U2520 (N_2520,In_2938,In_2885);
or U2521 (N_2521,In_720,In_1889);
or U2522 (N_2522,In_2110,In_1583);
or U2523 (N_2523,In_2362,In_1174);
nand U2524 (N_2524,In_1424,In_1737);
nor U2525 (N_2525,In_1599,In_729);
and U2526 (N_2526,In_1118,In_633);
nand U2527 (N_2527,In_2763,In_241);
and U2528 (N_2528,In_1101,In_351);
and U2529 (N_2529,In_721,In_2123);
or U2530 (N_2530,In_747,In_1111);
nand U2531 (N_2531,In_504,In_1104);
and U2532 (N_2532,In_866,In_1857);
and U2533 (N_2533,In_145,In_2353);
nor U2534 (N_2534,In_1409,In_2263);
nand U2535 (N_2535,In_924,In_2275);
nor U2536 (N_2536,In_2495,In_333);
nor U2537 (N_2537,In_1790,In_1634);
nor U2538 (N_2538,In_2503,In_1231);
nor U2539 (N_2539,In_456,In_1234);
xnor U2540 (N_2540,In_2389,In_1819);
and U2541 (N_2541,In_2289,In_1617);
nor U2542 (N_2542,In_808,In_50);
and U2543 (N_2543,In_2943,In_2865);
or U2544 (N_2544,In_2962,In_393);
nand U2545 (N_2545,In_869,In_1800);
and U2546 (N_2546,In_1871,In_2848);
nand U2547 (N_2547,In_2741,In_1516);
nor U2548 (N_2548,In_2807,In_2069);
nand U2549 (N_2549,In_2385,In_849);
nand U2550 (N_2550,In_2373,In_493);
or U2551 (N_2551,In_1916,In_2541);
or U2552 (N_2552,In_817,In_943);
nand U2553 (N_2553,In_532,In_1233);
xnor U2554 (N_2554,In_2151,In_2633);
or U2555 (N_2555,In_1121,In_499);
or U2556 (N_2556,In_1969,In_1225);
nor U2557 (N_2557,In_2644,In_2833);
xor U2558 (N_2558,In_371,In_1884);
and U2559 (N_2559,In_2657,In_310);
or U2560 (N_2560,In_1190,In_1004);
or U2561 (N_2561,In_19,In_594);
xnor U2562 (N_2562,In_2714,In_1454);
xnor U2563 (N_2563,In_2072,In_2675);
and U2564 (N_2564,In_519,In_389);
and U2565 (N_2565,In_1343,In_2602);
nand U2566 (N_2566,In_2998,In_2540);
and U2567 (N_2567,In_2786,In_2904);
and U2568 (N_2568,In_1838,In_1554);
nor U2569 (N_2569,In_105,In_1358);
nor U2570 (N_2570,In_1148,In_2802);
or U2571 (N_2571,In_708,In_2759);
nand U2572 (N_2572,In_2766,In_1788);
or U2573 (N_2573,In_455,In_2768);
or U2574 (N_2574,In_1483,In_1408);
nor U2575 (N_2575,In_1938,In_2344);
or U2576 (N_2576,In_1599,In_1630);
and U2577 (N_2577,In_2351,In_119);
and U2578 (N_2578,In_2483,In_698);
xnor U2579 (N_2579,In_298,In_1894);
or U2580 (N_2580,In_1789,In_2077);
nand U2581 (N_2581,In_303,In_2777);
xor U2582 (N_2582,In_1141,In_209);
nand U2583 (N_2583,In_1007,In_2806);
nand U2584 (N_2584,In_804,In_1489);
nor U2585 (N_2585,In_1250,In_890);
nand U2586 (N_2586,In_1458,In_2065);
or U2587 (N_2587,In_2541,In_367);
nor U2588 (N_2588,In_1723,In_2899);
or U2589 (N_2589,In_2420,In_2365);
nor U2590 (N_2590,In_2754,In_2557);
nand U2591 (N_2591,In_1674,In_1889);
or U2592 (N_2592,In_1941,In_1394);
nor U2593 (N_2593,In_1422,In_217);
nand U2594 (N_2594,In_1709,In_1966);
nor U2595 (N_2595,In_272,In_1657);
or U2596 (N_2596,In_2861,In_2377);
nor U2597 (N_2597,In_2338,In_1746);
nor U2598 (N_2598,In_1131,In_1543);
or U2599 (N_2599,In_81,In_2143);
nand U2600 (N_2600,In_2379,In_2848);
or U2601 (N_2601,In_1506,In_1604);
nor U2602 (N_2602,In_2276,In_1338);
nor U2603 (N_2603,In_2411,In_2772);
nor U2604 (N_2604,In_2163,In_2300);
and U2605 (N_2605,In_1575,In_2642);
nand U2606 (N_2606,In_1718,In_67);
nand U2607 (N_2607,In_2358,In_1814);
nand U2608 (N_2608,In_2762,In_2165);
nand U2609 (N_2609,In_2319,In_2800);
nand U2610 (N_2610,In_2672,In_2476);
nand U2611 (N_2611,In_1793,In_2714);
nor U2612 (N_2612,In_890,In_1102);
xor U2613 (N_2613,In_1101,In_2798);
or U2614 (N_2614,In_546,In_88);
nand U2615 (N_2615,In_864,In_2898);
nand U2616 (N_2616,In_405,In_2462);
nor U2617 (N_2617,In_1070,In_2786);
or U2618 (N_2618,In_399,In_1302);
or U2619 (N_2619,In_2294,In_913);
nand U2620 (N_2620,In_1445,In_230);
and U2621 (N_2621,In_1922,In_2218);
or U2622 (N_2622,In_1994,In_2285);
nand U2623 (N_2623,In_1134,In_276);
and U2624 (N_2624,In_258,In_1229);
or U2625 (N_2625,In_2395,In_2215);
nor U2626 (N_2626,In_1432,In_2051);
nand U2627 (N_2627,In_474,In_526);
nor U2628 (N_2628,In_2051,In_121);
nand U2629 (N_2629,In_308,In_1386);
or U2630 (N_2630,In_2100,In_2326);
nand U2631 (N_2631,In_936,In_2316);
nor U2632 (N_2632,In_2662,In_1727);
and U2633 (N_2633,In_2130,In_2580);
nand U2634 (N_2634,In_1123,In_902);
or U2635 (N_2635,In_380,In_2907);
nand U2636 (N_2636,In_1257,In_2600);
nand U2637 (N_2637,In_36,In_2984);
or U2638 (N_2638,In_575,In_1788);
nor U2639 (N_2639,In_1581,In_1256);
and U2640 (N_2640,In_1728,In_2340);
nand U2641 (N_2641,In_2122,In_1833);
nor U2642 (N_2642,In_882,In_532);
and U2643 (N_2643,In_1646,In_722);
xnor U2644 (N_2644,In_596,In_2464);
and U2645 (N_2645,In_1520,In_463);
or U2646 (N_2646,In_1276,In_1123);
or U2647 (N_2647,In_1733,In_34);
nand U2648 (N_2648,In_1047,In_177);
or U2649 (N_2649,In_279,In_565);
nand U2650 (N_2650,In_740,In_1898);
and U2651 (N_2651,In_1332,In_80);
nand U2652 (N_2652,In_1432,In_1499);
and U2653 (N_2653,In_724,In_631);
nand U2654 (N_2654,In_2488,In_613);
nand U2655 (N_2655,In_1156,In_2205);
and U2656 (N_2656,In_1532,In_2073);
nor U2657 (N_2657,In_621,In_2761);
nor U2658 (N_2658,In_1648,In_645);
or U2659 (N_2659,In_2585,In_1694);
or U2660 (N_2660,In_899,In_2577);
nand U2661 (N_2661,In_2307,In_2711);
or U2662 (N_2662,In_899,In_715);
nor U2663 (N_2663,In_1685,In_1858);
nand U2664 (N_2664,In_2030,In_1816);
or U2665 (N_2665,In_2110,In_1880);
or U2666 (N_2666,In_1931,In_252);
nor U2667 (N_2667,In_1478,In_1209);
and U2668 (N_2668,In_2474,In_1751);
and U2669 (N_2669,In_147,In_435);
xor U2670 (N_2670,In_953,In_2111);
xor U2671 (N_2671,In_1093,In_361);
nand U2672 (N_2672,In_1290,In_2995);
and U2673 (N_2673,In_2719,In_378);
and U2674 (N_2674,In_525,In_2589);
and U2675 (N_2675,In_465,In_1185);
or U2676 (N_2676,In_2073,In_2630);
nand U2677 (N_2677,In_2098,In_224);
xor U2678 (N_2678,In_1025,In_984);
or U2679 (N_2679,In_1638,In_2713);
nor U2680 (N_2680,In_2192,In_630);
or U2681 (N_2681,In_1851,In_1373);
nor U2682 (N_2682,In_2503,In_307);
nor U2683 (N_2683,In_2575,In_1636);
or U2684 (N_2684,In_1816,In_317);
or U2685 (N_2685,In_745,In_807);
or U2686 (N_2686,In_1403,In_1487);
nand U2687 (N_2687,In_1728,In_2126);
xor U2688 (N_2688,In_1448,In_873);
nand U2689 (N_2689,In_2864,In_176);
nor U2690 (N_2690,In_1371,In_758);
or U2691 (N_2691,In_1417,In_206);
and U2692 (N_2692,In_915,In_2128);
nand U2693 (N_2693,In_2275,In_406);
nand U2694 (N_2694,In_1692,In_182);
nand U2695 (N_2695,In_638,In_659);
nand U2696 (N_2696,In_1706,In_1548);
and U2697 (N_2697,In_92,In_1348);
and U2698 (N_2698,In_2706,In_295);
or U2699 (N_2699,In_1178,In_453);
nand U2700 (N_2700,In_797,In_2333);
and U2701 (N_2701,In_1586,In_1005);
xor U2702 (N_2702,In_1551,In_2924);
nor U2703 (N_2703,In_1000,In_822);
nor U2704 (N_2704,In_1946,In_2883);
and U2705 (N_2705,In_1176,In_1223);
or U2706 (N_2706,In_13,In_2317);
nor U2707 (N_2707,In_2361,In_2305);
nor U2708 (N_2708,In_946,In_80);
nor U2709 (N_2709,In_1975,In_289);
nor U2710 (N_2710,In_2341,In_284);
nor U2711 (N_2711,In_2382,In_2434);
or U2712 (N_2712,In_1115,In_537);
or U2713 (N_2713,In_2265,In_1266);
nor U2714 (N_2714,In_1862,In_1621);
nand U2715 (N_2715,In_2728,In_2525);
and U2716 (N_2716,In_4,In_1030);
xor U2717 (N_2717,In_1570,In_102);
nor U2718 (N_2718,In_2629,In_2126);
or U2719 (N_2719,In_1358,In_542);
and U2720 (N_2720,In_2258,In_2882);
or U2721 (N_2721,In_94,In_24);
nor U2722 (N_2722,In_194,In_720);
nor U2723 (N_2723,In_2600,In_1726);
and U2724 (N_2724,In_1878,In_707);
nand U2725 (N_2725,In_2725,In_1646);
or U2726 (N_2726,In_1452,In_796);
nand U2727 (N_2727,In_1634,In_1961);
nor U2728 (N_2728,In_2771,In_68);
nand U2729 (N_2729,In_2977,In_1078);
or U2730 (N_2730,In_2113,In_2460);
and U2731 (N_2731,In_1662,In_1095);
and U2732 (N_2732,In_1284,In_349);
nor U2733 (N_2733,In_2981,In_2316);
and U2734 (N_2734,In_1782,In_1818);
or U2735 (N_2735,In_386,In_1832);
nand U2736 (N_2736,In_2604,In_2616);
and U2737 (N_2737,In_303,In_1046);
xnor U2738 (N_2738,In_703,In_1524);
nor U2739 (N_2739,In_456,In_1743);
nand U2740 (N_2740,In_2763,In_180);
nor U2741 (N_2741,In_1571,In_660);
and U2742 (N_2742,In_1333,In_1795);
nand U2743 (N_2743,In_241,In_393);
or U2744 (N_2744,In_973,In_1045);
nor U2745 (N_2745,In_1026,In_763);
nand U2746 (N_2746,In_879,In_2902);
nor U2747 (N_2747,In_2265,In_91);
xnor U2748 (N_2748,In_310,In_2347);
or U2749 (N_2749,In_289,In_1916);
nand U2750 (N_2750,In_2657,In_76);
nand U2751 (N_2751,In_1029,In_1007);
nor U2752 (N_2752,In_2546,In_1897);
nor U2753 (N_2753,In_529,In_1435);
nor U2754 (N_2754,In_1787,In_2976);
and U2755 (N_2755,In_726,In_518);
and U2756 (N_2756,In_1898,In_1379);
nor U2757 (N_2757,In_2237,In_2059);
xnor U2758 (N_2758,In_2079,In_2975);
xnor U2759 (N_2759,In_539,In_2693);
nand U2760 (N_2760,In_626,In_1144);
nand U2761 (N_2761,In_2506,In_753);
or U2762 (N_2762,In_2727,In_1847);
nand U2763 (N_2763,In_92,In_111);
or U2764 (N_2764,In_2639,In_2789);
nor U2765 (N_2765,In_2657,In_1174);
xor U2766 (N_2766,In_429,In_1055);
and U2767 (N_2767,In_1852,In_403);
and U2768 (N_2768,In_2990,In_1366);
and U2769 (N_2769,In_1047,In_2230);
nand U2770 (N_2770,In_1000,In_2484);
nand U2771 (N_2771,In_1685,In_2800);
nor U2772 (N_2772,In_802,In_721);
nor U2773 (N_2773,In_243,In_177);
and U2774 (N_2774,In_1814,In_2661);
or U2775 (N_2775,In_660,In_1270);
and U2776 (N_2776,In_1709,In_1556);
nor U2777 (N_2777,In_678,In_103);
and U2778 (N_2778,In_1350,In_125);
nor U2779 (N_2779,In_2968,In_535);
nor U2780 (N_2780,In_2385,In_1722);
nand U2781 (N_2781,In_1121,In_1040);
and U2782 (N_2782,In_2894,In_1372);
or U2783 (N_2783,In_1683,In_1956);
nor U2784 (N_2784,In_2380,In_994);
or U2785 (N_2785,In_47,In_216);
and U2786 (N_2786,In_1091,In_1099);
nor U2787 (N_2787,In_1500,In_447);
nor U2788 (N_2788,In_2588,In_2849);
nor U2789 (N_2789,In_1352,In_607);
or U2790 (N_2790,In_1375,In_1853);
nand U2791 (N_2791,In_2786,In_2052);
nand U2792 (N_2792,In_1169,In_737);
xor U2793 (N_2793,In_1809,In_2776);
nand U2794 (N_2794,In_83,In_1046);
or U2795 (N_2795,In_1412,In_2878);
nor U2796 (N_2796,In_2710,In_612);
nor U2797 (N_2797,In_547,In_400);
nor U2798 (N_2798,In_1435,In_2050);
and U2799 (N_2799,In_1552,In_661);
nand U2800 (N_2800,In_2995,In_121);
or U2801 (N_2801,In_2985,In_270);
nand U2802 (N_2802,In_1367,In_2278);
and U2803 (N_2803,In_1958,In_420);
and U2804 (N_2804,In_618,In_2926);
nand U2805 (N_2805,In_1956,In_1240);
nand U2806 (N_2806,In_2526,In_108);
nand U2807 (N_2807,In_1048,In_1525);
or U2808 (N_2808,In_1289,In_2824);
nor U2809 (N_2809,In_274,In_47);
xor U2810 (N_2810,In_57,In_975);
nor U2811 (N_2811,In_231,In_1458);
and U2812 (N_2812,In_1469,In_2019);
and U2813 (N_2813,In_2268,In_308);
nor U2814 (N_2814,In_2419,In_1667);
and U2815 (N_2815,In_1522,In_1651);
nand U2816 (N_2816,In_454,In_2997);
nand U2817 (N_2817,In_2905,In_2407);
nand U2818 (N_2818,In_2839,In_1403);
or U2819 (N_2819,In_2959,In_1317);
nor U2820 (N_2820,In_1363,In_898);
nand U2821 (N_2821,In_793,In_2869);
xnor U2822 (N_2822,In_2621,In_1181);
or U2823 (N_2823,In_763,In_1680);
or U2824 (N_2824,In_1817,In_1216);
and U2825 (N_2825,In_2166,In_2983);
or U2826 (N_2826,In_1485,In_2521);
nand U2827 (N_2827,In_416,In_1367);
nor U2828 (N_2828,In_116,In_346);
or U2829 (N_2829,In_414,In_2506);
and U2830 (N_2830,In_2625,In_321);
nand U2831 (N_2831,In_2710,In_666);
nand U2832 (N_2832,In_1499,In_1357);
or U2833 (N_2833,In_2184,In_2366);
nor U2834 (N_2834,In_1610,In_1027);
and U2835 (N_2835,In_2720,In_1514);
nand U2836 (N_2836,In_1124,In_740);
and U2837 (N_2837,In_1670,In_2893);
nor U2838 (N_2838,In_109,In_847);
nand U2839 (N_2839,In_22,In_2288);
nand U2840 (N_2840,In_2358,In_1685);
xor U2841 (N_2841,In_2004,In_1921);
nor U2842 (N_2842,In_446,In_2225);
or U2843 (N_2843,In_1827,In_1816);
or U2844 (N_2844,In_2480,In_1284);
nor U2845 (N_2845,In_2401,In_1661);
or U2846 (N_2846,In_2749,In_1326);
nor U2847 (N_2847,In_1080,In_1773);
nand U2848 (N_2848,In_1878,In_2187);
nand U2849 (N_2849,In_2760,In_1753);
nand U2850 (N_2850,In_2031,In_641);
or U2851 (N_2851,In_466,In_1020);
or U2852 (N_2852,In_1860,In_2387);
or U2853 (N_2853,In_668,In_7);
or U2854 (N_2854,In_1496,In_984);
or U2855 (N_2855,In_201,In_1580);
nor U2856 (N_2856,In_1878,In_1222);
and U2857 (N_2857,In_1518,In_549);
or U2858 (N_2858,In_1562,In_826);
or U2859 (N_2859,In_1057,In_2892);
or U2860 (N_2860,In_2905,In_1712);
xor U2861 (N_2861,In_1681,In_2318);
nand U2862 (N_2862,In_1936,In_2130);
xnor U2863 (N_2863,In_1549,In_34);
nor U2864 (N_2864,In_787,In_2768);
nand U2865 (N_2865,In_2290,In_2241);
or U2866 (N_2866,In_1122,In_1060);
nor U2867 (N_2867,In_497,In_618);
and U2868 (N_2868,In_1409,In_1677);
nor U2869 (N_2869,In_1705,In_916);
nand U2870 (N_2870,In_448,In_2821);
nand U2871 (N_2871,In_2427,In_1010);
nor U2872 (N_2872,In_2713,In_2042);
nand U2873 (N_2873,In_828,In_2340);
or U2874 (N_2874,In_582,In_2425);
and U2875 (N_2875,In_2661,In_2643);
and U2876 (N_2876,In_1121,In_1290);
and U2877 (N_2877,In_1644,In_2274);
and U2878 (N_2878,In_115,In_2320);
nand U2879 (N_2879,In_1616,In_1225);
or U2880 (N_2880,In_840,In_813);
or U2881 (N_2881,In_1023,In_1404);
and U2882 (N_2882,In_573,In_1645);
nor U2883 (N_2883,In_359,In_2988);
nor U2884 (N_2884,In_1228,In_2264);
xnor U2885 (N_2885,In_461,In_711);
or U2886 (N_2886,In_1968,In_1842);
or U2887 (N_2887,In_496,In_2855);
xor U2888 (N_2888,In_1583,In_2957);
nor U2889 (N_2889,In_259,In_315);
nand U2890 (N_2890,In_404,In_154);
nor U2891 (N_2891,In_624,In_2864);
xnor U2892 (N_2892,In_1676,In_86);
nand U2893 (N_2893,In_2630,In_636);
or U2894 (N_2894,In_1809,In_2047);
and U2895 (N_2895,In_2158,In_784);
or U2896 (N_2896,In_1857,In_2742);
or U2897 (N_2897,In_2195,In_1492);
or U2898 (N_2898,In_1481,In_844);
or U2899 (N_2899,In_978,In_907);
and U2900 (N_2900,In_747,In_2141);
nor U2901 (N_2901,In_1250,In_769);
and U2902 (N_2902,In_1429,In_2963);
and U2903 (N_2903,In_928,In_2064);
nand U2904 (N_2904,In_1713,In_886);
or U2905 (N_2905,In_2288,In_2920);
nand U2906 (N_2906,In_1041,In_1720);
xnor U2907 (N_2907,In_197,In_401);
nand U2908 (N_2908,In_1168,In_2819);
nand U2909 (N_2909,In_1942,In_1041);
nor U2910 (N_2910,In_1442,In_1898);
nand U2911 (N_2911,In_1983,In_152);
nor U2912 (N_2912,In_2642,In_2953);
nor U2913 (N_2913,In_815,In_1538);
or U2914 (N_2914,In_2923,In_2481);
nand U2915 (N_2915,In_2551,In_1241);
nand U2916 (N_2916,In_675,In_2436);
nor U2917 (N_2917,In_379,In_2811);
or U2918 (N_2918,In_288,In_933);
and U2919 (N_2919,In_1124,In_1507);
and U2920 (N_2920,In_1759,In_2679);
nor U2921 (N_2921,In_2607,In_994);
xor U2922 (N_2922,In_904,In_581);
nor U2923 (N_2923,In_1971,In_1798);
nor U2924 (N_2924,In_299,In_1211);
nand U2925 (N_2925,In_2231,In_600);
nor U2926 (N_2926,In_302,In_1022);
or U2927 (N_2927,In_1814,In_939);
nor U2928 (N_2928,In_371,In_1029);
nand U2929 (N_2929,In_428,In_2326);
nor U2930 (N_2930,In_2999,In_2766);
nand U2931 (N_2931,In_1176,In_260);
and U2932 (N_2932,In_843,In_2079);
or U2933 (N_2933,In_883,In_1224);
nor U2934 (N_2934,In_1470,In_2535);
nor U2935 (N_2935,In_2158,In_977);
and U2936 (N_2936,In_2720,In_1526);
or U2937 (N_2937,In_2477,In_1867);
nand U2938 (N_2938,In_1435,In_994);
nand U2939 (N_2939,In_524,In_230);
and U2940 (N_2940,In_9,In_957);
or U2941 (N_2941,In_2761,In_430);
and U2942 (N_2942,In_1993,In_741);
and U2943 (N_2943,In_170,In_2293);
and U2944 (N_2944,In_1001,In_1116);
or U2945 (N_2945,In_473,In_511);
or U2946 (N_2946,In_806,In_2673);
nor U2947 (N_2947,In_739,In_1759);
and U2948 (N_2948,In_1228,In_1617);
nor U2949 (N_2949,In_1957,In_2262);
and U2950 (N_2950,In_431,In_2012);
or U2951 (N_2951,In_1008,In_2814);
nand U2952 (N_2952,In_1355,In_462);
xor U2953 (N_2953,In_2099,In_2536);
nand U2954 (N_2954,In_1604,In_619);
xnor U2955 (N_2955,In_1457,In_1918);
and U2956 (N_2956,In_847,In_681);
nand U2957 (N_2957,In_2521,In_532);
nand U2958 (N_2958,In_73,In_213);
nor U2959 (N_2959,In_2055,In_2871);
nor U2960 (N_2960,In_1074,In_1724);
or U2961 (N_2961,In_2369,In_1136);
xor U2962 (N_2962,In_1070,In_194);
nor U2963 (N_2963,In_699,In_365);
nor U2964 (N_2964,In_376,In_282);
or U2965 (N_2965,In_624,In_2519);
nor U2966 (N_2966,In_1163,In_2117);
nor U2967 (N_2967,In_931,In_1112);
or U2968 (N_2968,In_781,In_1212);
xor U2969 (N_2969,In_2257,In_882);
nand U2970 (N_2970,In_2475,In_861);
nand U2971 (N_2971,In_2197,In_2134);
nor U2972 (N_2972,In_2132,In_574);
xnor U2973 (N_2973,In_2780,In_483);
nand U2974 (N_2974,In_2134,In_2786);
and U2975 (N_2975,In_655,In_615);
and U2976 (N_2976,In_2827,In_2159);
or U2977 (N_2977,In_595,In_203);
nor U2978 (N_2978,In_168,In_1094);
nand U2979 (N_2979,In_1702,In_813);
nor U2980 (N_2980,In_151,In_539);
nand U2981 (N_2981,In_753,In_1209);
xor U2982 (N_2982,In_1987,In_466);
and U2983 (N_2983,In_181,In_2038);
and U2984 (N_2984,In_2113,In_1032);
nor U2985 (N_2985,In_1001,In_2094);
or U2986 (N_2986,In_117,In_2853);
and U2987 (N_2987,In_2392,In_2562);
nor U2988 (N_2988,In_2771,In_1393);
or U2989 (N_2989,In_2181,In_224);
nand U2990 (N_2990,In_2249,In_2714);
nand U2991 (N_2991,In_1939,In_932);
nor U2992 (N_2992,In_706,In_2000);
nand U2993 (N_2993,In_208,In_745);
and U2994 (N_2994,In_344,In_2520);
and U2995 (N_2995,In_2537,In_651);
nand U2996 (N_2996,In_153,In_2981);
or U2997 (N_2997,In_82,In_1729);
and U2998 (N_2998,In_153,In_2811);
nor U2999 (N_2999,In_771,In_143);
and U3000 (N_3000,In_1459,In_1808);
nor U3001 (N_3001,In_2588,In_1205);
or U3002 (N_3002,In_2712,In_1369);
and U3003 (N_3003,In_1077,In_2170);
nand U3004 (N_3004,In_2034,In_2025);
nor U3005 (N_3005,In_1691,In_74);
nor U3006 (N_3006,In_1844,In_1040);
or U3007 (N_3007,In_1239,In_2407);
nor U3008 (N_3008,In_2765,In_2726);
nand U3009 (N_3009,In_2180,In_2590);
nand U3010 (N_3010,In_2201,In_938);
nor U3011 (N_3011,In_2454,In_1664);
nor U3012 (N_3012,In_984,In_191);
nor U3013 (N_3013,In_2726,In_1557);
xnor U3014 (N_3014,In_2981,In_2441);
nor U3015 (N_3015,In_876,In_1360);
and U3016 (N_3016,In_2196,In_1040);
or U3017 (N_3017,In_1071,In_2510);
or U3018 (N_3018,In_1433,In_847);
or U3019 (N_3019,In_1036,In_159);
and U3020 (N_3020,In_762,In_516);
and U3021 (N_3021,In_2824,In_1297);
nand U3022 (N_3022,In_52,In_404);
nand U3023 (N_3023,In_2822,In_1982);
and U3024 (N_3024,In_2555,In_2309);
or U3025 (N_3025,In_2051,In_2075);
nor U3026 (N_3026,In_2694,In_178);
nand U3027 (N_3027,In_2251,In_500);
nand U3028 (N_3028,In_2525,In_562);
nand U3029 (N_3029,In_2105,In_1051);
or U3030 (N_3030,In_2007,In_1774);
and U3031 (N_3031,In_2311,In_1928);
nor U3032 (N_3032,In_465,In_1503);
and U3033 (N_3033,In_1812,In_929);
or U3034 (N_3034,In_1992,In_2382);
and U3035 (N_3035,In_1725,In_1271);
nand U3036 (N_3036,In_2566,In_1635);
or U3037 (N_3037,In_10,In_1653);
or U3038 (N_3038,In_2807,In_2525);
or U3039 (N_3039,In_1859,In_1701);
or U3040 (N_3040,In_2735,In_1962);
nand U3041 (N_3041,In_1189,In_29);
xor U3042 (N_3042,In_2464,In_2544);
xnor U3043 (N_3043,In_195,In_1029);
nand U3044 (N_3044,In_363,In_499);
nand U3045 (N_3045,In_78,In_343);
nor U3046 (N_3046,In_1330,In_2914);
and U3047 (N_3047,In_389,In_1107);
xor U3048 (N_3048,In_1492,In_1917);
nand U3049 (N_3049,In_2971,In_1172);
nand U3050 (N_3050,In_2832,In_2633);
and U3051 (N_3051,In_848,In_1898);
nor U3052 (N_3052,In_322,In_2375);
nor U3053 (N_3053,In_2601,In_2384);
and U3054 (N_3054,In_193,In_569);
xnor U3055 (N_3055,In_2583,In_1826);
or U3056 (N_3056,In_1740,In_2797);
or U3057 (N_3057,In_1572,In_2658);
or U3058 (N_3058,In_799,In_1532);
nand U3059 (N_3059,In_2246,In_836);
nor U3060 (N_3060,In_1318,In_2002);
and U3061 (N_3061,In_1667,In_880);
and U3062 (N_3062,In_1761,In_1176);
and U3063 (N_3063,In_1598,In_147);
nand U3064 (N_3064,In_1981,In_2801);
and U3065 (N_3065,In_2969,In_107);
nand U3066 (N_3066,In_2859,In_1894);
and U3067 (N_3067,In_1677,In_2439);
nor U3068 (N_3068,In_1105,In_2097);
nor U3069 (N_3069,In_387,In_920);
nor U3070 (N_3070,In_1414,In_2008);
nor U3071 (N_3071,In_1853,In_1992);
nor U3072 (N_3072,In_158,In_978);
nand U3073 (N_3073,In_2093,In_252);
or U3074 (N_3074,In_627,In_765);
and U3075 (N_3075,In_2348,In_184);
or U3076 (N_3076,In_329,In_2946);
xor U3077 (N_3077,In_1163,In_888);
and U3078 (N_3078,In_9,In_2115);
and U3079 (N_3079,In_1479,In_973);
and U3080 (N_3080,In_1995,In_2087);
nor U3081 (N_3081,In_1532,In_640);
nand U3082 (N_3082,In_2972,In_325);
nand U3083 (N_3083,In_2019,In_2060);
nand U3084 (N_3084,In_1665,In_2090);
nor U3085 (N_3085,In_2657,In_1844);
and U3086 (N_3086,In_2610,In_1583);
nor U3087 (N_3087,In_1413,In_411);
nand U3088 (N_3088,In_220,In_2788);
and U3089 (N_3089,In_1759,In_1605);
nand U3090 (N_3090,In_2673,In_1464);
and U3091 (N_3091,In_747,In_2618);
and U3092 (N_3092,In_1794,In_510);
nand U3093 (N_3093,In_2247,In_2620);
nor U3094 (N_3094,In_298,In_285);
nand U3095 (N_3095,In_895,In_741);
nand U3096 (N_3096,In_186,In_2860);
nor U3097 (N_3097,In_1964,In_1905);
xor U3098 (N_3098,In_2481,In_978);
and U3099 (N_3099,In_1447,In_2689);
and U3100 (N_3100,In_2798,In_1631);
or U3101 (N_3101,In_4,In_249);
and U3102 (N_3102,In_1971,In_1796);
and U3103 (N_3103,In_2145,In_2765);
or U3104 (N_3104,In_2191,In_1915);
nand U3105 (N_3105,In_903,In_1942);
or U3106 (N_3106,In_2800,In_712);
xnor U3107 (N_3107,In_1099,In_114);
nand U3108 (N_3108,In_1547,In_392);
and U3109 (N_3109,In_2796,In_1160);
nor U3110 (N_3110,In_1384,In_2218);
nand U3111 (N_3111,In_1059,In_2275);
nand U3112 (N_3112,In_2692,In_2959);
nand U3113 (N_3113,In_1986,In_338);
and U3114 (N_3114,In_2738,In_2233);
and U3115 (N_3115,In_48,In_2186);
nor U3116 (N_3116,In_1475,In_1408);
and U3117 (N_3117,In_2183,In_1647);
nor U3118 (N_3118,In_2759,In_127);
nor U3119 (N_3119,In_2521,In_1611);
nor U3120 (N_3120,In_1617,In_201);
nand U3121 (N_3121,In_797,In_1732);
nor U3122 (N_3122,In_166,In_491);
nand U3123 (N_3123,In_1945,In_990);
nand U3124 (N_3124,In_704,In_2636);
and U3125 (N_3125,In_759,In_2649);
nor U3126 (N_3126,In_509,In_1804);
nor U3127 (N_3127,In_1399,In_2347);
nand U3128 (N_3128,In_768,In_1737);
nand U3129 (N_3129,In_2127,In_2476);
and U3130 (N_3130,In_1233,In_1520);
nor U3131 (N_3131,In_2550,In_1346);
nand U3132 (N_3132,In_721,In_1006);
or U3133 (N_3133,In_2370,In_2495);
or U3134 (N_3134,In_379,In_1873);
xnor U3135 (N_3135,In_2465,In_1407);
or U3136 (N_3136,In_505,In_2636);
nor U3137 (N_3137,In_363,In_1882);
or U3138 (N_3138,In_2987,In_1887);
nand U3139 (N_3139,In_1858,In_1850);
nor U3140 (N_3140,In_2691,In_1723);
nor U3141 (N_3141,In_1521,In_2896);
xnor U3142 (N_3142,In_310,In_276);
xor U3143 (N_3143,In_1701,In_2723);
nand U3144 (N_3144,In_1843,In_413);
nor U3145 (N_3145,In_2281,In_2559);
nor U3146 (N_3146,In_612,In_364);
and U3147 (N_3147,In_1943,In_882);
or U3148 (N_3148,In_2154,In_142);
or U3149 (N_3149,In_2623,In_89);
nor U3150 (N_3150,In_2762,In_657);
and U3151 (N_3151,In_929,In_1773);
and U3152 (N_3152,In_778,In_661);
or U3153 (N_3153,In_2626,In_2855);
nor U3154 (N_3154,In_704,In_161);
nand U3155 (N_3155,In_2965,In_2329);
and U3156 (N_3156,In_1484,In_2917);
nand U3157 (N_3157,In_2737,In_2322);
and U3158 (N_3158,In_2587,In_2929);
nor U3159 (N_3159,In_2603,In_2261);
nor U3160 (N_3160,In_1560,In_2828);
nor U3161 (N_3161,In_2215,In_1466);
or U3162 (N_3162,In_628,In_2424);
and U3163 (N_3163,In_20,In_2990);
and U3164 (N_3164,In_944,In_178);
nor U3165 (N_3165,In_2633,In_1078);
nor U3166 (N_3166,In_2643,In_1119);
and U3167 (N_3167,In_1775,In_1163);
xnor U3168 (N_3168,In_1067,In_1);
nand U3169 (N_3169,In_2314,In_1858);
xor U3170 (N_3170,In_1748,In_1979);
nand U3171 (N_3171,In_2683,In_273);
nor U3172 (N_3172,In_2693,In_898);
nor U3173 (N_3173,In_2488,In_2786);
or U3174 (N_3174,In_882,In_655);
nand U3175 (N_3175,In_1140,In_428);
nor U3176 (N_3176,In_1802,In_241);
nor U3177 (N_3177,In_2220,In_1836);
or U3178 (N_3178,In_1789,In_721);
nand U3179 (N_3179,In_1478,In_534);
and U3180 (N_3180,In_891,In_1296);
or U3181 (N_3181,In_288,In_1733);
nand U3182 (N_3182,In_1048,In_2567);
xor U3183 (N_3183,In_280,In_862);
or U3184 (N_3184,In_1271,In_2697);
nor U3185 (N_3185,In_1260,In_2282);
and U3186 (N_3186,In_1385,In_2243);
and U3187 (N_3187,In_898,In_2137);
xor U3188 (N_3188,In_2400,In_2722);
or U3189 (N_3189,In_2941,In_2628);
or U3190 (N_3190,In_1458,In_724);
nand U3191 (N_3191,In_2974,In_2165);
or U3192 (N_3192,In_2263,In_2642);
or U3193 (N_3193,In_2731,In_302);
or U3194 (N_3194,In_1783,In_1097);
and U3195 (N_3195,In_1530,In_804);
xnor U3196 (N_3196,In_1563,In_1864);
and U3197 (N_3197,In_275,In_1759);
and U3198 (N_3198,In_323,In_368);
xor U3199 (N_3199,In_2433,In_2854);
nor U3200 (N_3200,In_1053,In_298);
or U3201 (N_3201,In_1715,In_2910);
or U3202 (N_3202,In_2497,In_933);
nor U3203 (N_3203,In_1044,In_2847);
and U3204 (N_3204,In_1942,In_2472);
nand U3205 (N_3205,In_415,In_726);
or U3206 (N_3206,In_572,In_1304);
or U3207 (N_3207,In_549,In_17);
nand U3208 (N_3208,In_1290,In_271);
nand U3209 (N_3209,In_1152,In_2480);
nor U3210 (N_3210,In_2994,In_2944);
nand U3211 (N_3211,In_1873,In_1906);
and U3212 (N_3212,In_2731,In_2329);
nor U3213 (N_3213,In_793,In_632);
and U3214 (N_3214,In_719,In_513);
nand U3215 (N_3215,In_1349,In_236);
nor U3216 (N_3216,In_2433,In_893);
or U3217 (N_3217,In_1899,In_2048);
nand U3218 (N_3218,In_2690,In_425);
and U3219 (N_3219,In_2911,In_1995);
nand U3220 (N_3220,In_1511,In_2123);
nor U3221 (N_3221,In_2932,In_1498);
and U3222 (N_3222,In_2057,In_2704);
nor U3223 (N_3223,In_1512,In_2458);
xor U3224 (N_3224,In_1673,In_2607);
nor U3225 (N_3225,In_887,In_673);
xor U3226 (N_3226,In_2366,In_2009);
nor U3227 (N_3227,In_2628,In_2874);
nand U3228 (N_3228,In_1169,In_619);
xor U3229 (N_3229,In_1903,In_2136);
nor U3230 (N_3230,In_1054,In_2536);
or U3231 (N_3231,In_2715,In_2761);
xor U3232 (N_3232,In_1572,In_2311);
nor U3233 (N_3233,In_2542,In_637);
or U3234 (N_3234,In_1399,In_2775);
nor U3235 (N_3235,In_474,In_2422);
and U3236 (N_3236,In_1450,In_1673);
nand U3237 (N_3237,In_615,In_100);
nor U3238 (N_3238,In_2100,In_725);
nand U3239 (N_3239,In_2520,In_1181);
nor U3240 (N_3240,In_2546,In_2136);
xnor U3241 (N_3241,In_1028,In_2292);
nor U3242 (N_3242,In_2785,In_1080);
nor U3243 (N_3243,In_1844,In_2670);
nor U3244 (N_3244,In_1296,In_1954);
or U3245 (N_3245,In_2116,In_353);
and U3246 (N_3246,In_2088,In_2559);
or U3247 (N_3247,In_562,In_592);
and U3248 (N_3248,In_2819,In_1428);
or U3249 (N_3249,In_537,In_1740);
xor U3250 (N_3250,In_1402,In_1139);
nor U3251 (N_3251,In_2600,In_739);
nor U3252 (N_3252,In_1775,In_1922);
xor U3253 (N_3253,In_1345,In_298);
and U3254 (N_3254,In_1846,In_2843);
nand U3255 (N_3255,In_524,In_2874);
nand U3256 (N_3256,In_887,In_2898);
nand U3257 (N_3257,In_838,In_558);
nor U3258 (N_3258,In_1021,In_745);
and U3259 (N_3259,In_1590,In_2770);
and U3260 (N_3260,In_33,In_1188);
and U3261 (N_3261,In_2865,In_279);
and U3262 (N_3262,In_2139,In_1226);
nor U3263 (N_3263,In_859,In_1123);
xnor U3264 (N_3264,In_382,In_2827);
nor U3265 (N_3265,In_2030,In_279);
and U3266 (N_3266,In_2785,In_2637);
or U3267 (N_3267,In_2986,In_1175);
or U3268 (N_3268,In_803,In_1932);
xor U3269 (N_3269,In_2832,In_476);
nor U3270 (N_3270,In_183,In_780);
nor U3271 (N_3271,In_1881,In_2866);
or U3272 (N_3272,In_2410,In_1811);
nand U3273 (N_3273,In_2390,In_265);
and U3274 (N_3274,In_25,In_2607);
or U3275 (N_3275,In_1447,In_1228);
nand U3276 (N_3276,In_1649,In_820);
nand U3277 (N_3277,In_744,In_264);
nand U3278 (N_3278,In_1091,In_2755);
or U3279 (N_3279,In_1229,In_639);
and U3280 (N_3280,In_392,In_789);
or U3281 (N_3281,In_67,In_1455);
nand U3282 (N_3282,In_1387,In_883);
nand U3283 (N_3283,In_2443,In_2209);
and U3284 (N_3284,In_2942,In_1981);
or U3285 (N_3285,In_109,In_230);
and U3286 (N_3286,In_1706,In_2583);
or U3287 (N_3287,In_1346,In_1787);
or U3288 (N_3288,In_1592,In_1241);
nor U3289 (N_3289,In_294,In_1944);
and U3290 (N_3290,In_969,In_2722);
nand U3291 (N_3291,In_2248,In_2345);
nor U3292 (N_3292,In_1908,In_360);
nor U3293 (N_3293,In_2516,In_63);
nor U3294 (N_3294,In_2202,In_1300);
xor U3295 (N_3295,In_1739,In_2730);
xnor U3296 (N_3296,In_25,In_852);
or U3297 (N_3297,In_616,In_2755);
and U3298 (N_3298,In_2517,In_2125);
nand U3299 (N_3299,In_1449,In_909);
nand U3300 (N_3300,In_1869,In_2654);
nor U3301 (N_3301,In_913,In_2490);
or U3302 (N_3302,In_1582,In_572);
nor U3303 (N_3303,In_2492,In_764);
and U3304 (N_3304,In_2898,In_2211);
and U3305 (N_3305,In_1203,In_1524);
nor U3306 (N_3306,In_1296,In_2490);
nor U3307 (N_3307,In_1332,In_543);
or U3308 (N_3308,In_1895,In_2951);
nor U3309 (N_3309,In_844,In_2183);
nand U3310 (N_3310,In_1896,In_2851);
nor U3311 (N_3311,In_2298,In_1885);
and U3312 (N_3312,In_2542,In_828);
or U3313 (N_3313,In_2378,In_2038);
or U3314 (N_3314,In_1773,In_82);
and U3315 (N_3315,In_2211,In_501);
or U3316 (N_3316,In_2707,In_2282);
nor U3317 (N_3317,In_2454,In_2227);
or U3318 (N_3318,In_1165,In_1526);
and U3319 (N_3319,In_643,In_1035);
nand U3320 (N_3320,In_2765,In_2969);
and U3321 (N_3321,In_992,In_978);
and U3322 (N_3322,In_1117,In_1495);
xor U3323 (N_3323,In_318,In_707);
xnor U3324 (N_3324,In_1001,In_2619);
or U3325 (N_3325,In_1164,In_1811);
nand U3326 (N_3326,In_1790,In_2901);
nand U3327 (N_3327,In_2635,In_380);
and U3328 (N_3328,In_879,In_2762);
nand U3329 (N_3329,In_2771,In_1158);
and U3330 (N_3330,In_1745,In_2609);
or U3331 (N_3331,In_2903,In_2077);
xor U3332 (N_3332,In_179,In_1979);
nor U3333 (N_3333,In_2068,In_464);
nor U3334 (N_3334,In_2905,In_1855);
or U3335 (N_3335,In_1707,In_2302);
xor U3336 (N_3336,In_2896,In_25);
nand U3337 (N_3337,In_1088,In_379);
or U3338 (N_3338,In_314,In_2705);
xnor U3339 (N_3339,In_2149,In_937);
or U3340 (N_3340,In_1072,In_2170);
or U3341 (N_3341,In_67,In_557);
nand U3342 (N_3342,In_2448,In_1188);
nor U3343 (N_3343,In_755,In_641);
nand U3344 (N_3344,In_355,In_2518);
xnor U3345 (N_3345,In_2954,In_1614);
xnor U3346 (N_3346,In_2995,In_903);
nor U3347 (N_3347,In_1108,In_2951);
nor U3348 (N_3348,In_494,In_857);
or U3349 (N_3349,In_2330,In_1096);
and U3350 (N_3350,In_1862,In_47);
nor U3351 (N_3351,In_798,In_2358);
or U3352 (N_3352,In_912,In_1227);
nor U3353 (N_3353,In_271,In_1407);
nor U3354 (N_3354,In_2883,In_2059);
nand U3355 (N_3355,In_1407,In_2692);
xor U3356 (N_3356,In_1201,In_293);
nand U3357 (N_3357,In_2672,In_795);
nand U3358 (N_3358,In_2665,In_366);
or U3359 (N_3359,In_113,In_199);
xor U3360 (N_3360,In_2658,In_2538);
nor U3361 (N_3361,In_754,In_1027);
and U3362 (N_3362,In_864,In_560);
xor U3363 (N_3363,In_1779,In_439);
nand U3364 (N_3364,In_290,In_2687);
nand U3365 (N_3365,In_2340,In_1640);
or U3366 (N_3366,In_1057,In_142);
nand U3367 (N_3367,In_159,In_2675);
nor U3368 (N_3368,In_77,In_2531);
xor U3369 (N_3369,In_682,In_1074);
nor U3370 (N_3370,In_2481,In_1591);
or U3371 (N_3371,In_1817,In_2612);
xnor U3372 (N_3372,In_897,In_2117);
nor U3373 (N_3373,In_1200,In_2374);
nand U3374 (N_3374,In_1922,In_2702);
nand U3375 (N_3375,In_359,In_2553);
xor U3376 (N_3376,In_2153,In_2432);
or U3377 (N_3377,In_273,In_2609);
nand U3378 (N_3378,In_1303,In_2430);
and U3379 (N_3379,In_2624,In_2097);
nor U3380 (N_3380,In_868,In_1497);
nand U3381 (N_3381,In_898,In_735);
or U3382 (N_3382,In_1470,In_527);
and U3383 (N_3383,In_1260,In_2835);
and U3384 (N_3384,In_1456,In_1296);
and U3385 (N_3385,In_891,In_640);
and U3386 (N_3386,In_248,In_1919);
nor U3387 (N_3387,In_67,In_2594);
xnor U3388 (N_3388,In_1183,In_2228);
nand U3389 (N_3389,In_2473,In_877);
or U3390 (N_3390,In_343,In_378);
nor U3391 (N_3391,In_1801,In_2269);
or U3392 (N_3392,In_767,In_53);
and U3393 (N_3393,In_2536,In_2864);
or U3394 (N_3394,In_2253,In_1745);
nand U3395 (N_3395,In_267,In_31);
nor U3396 (N_3396,In_98,In_849);
xnor U3397 (N_3397,In_2206,In_1191);
xor U3398 (N_3398,In_1930,In_1108);
and U3399 (N_3399,In_135,In_724);
nor U3400 (N_3400,In_443,In_2179);
or U3401 (N_3401,In_2999,In_1040);
nor U3402 (N_3402,In_1593,In_1895);
or U3403 (N_3403,In_2729,In_751);
and U3404 (N_3404,In_1331,In_904);
nand U3405 (N_3405,In_2587,In_670);
nand U3406 (N_3406,In_2418,In_2411);
nand U3407 (N_3407,In_1390,In_118);
and U3408 (N_3408,In_1382,In_2580);
xnor U3409 (N_3409,In_1412,In_2357);
nand U3410 (N_3410,In_1448,In_1461);
nor U3411 (N_3411,In_2391,In_2884);
or U3412 (N_3412,In_2603,In_1150);
and U3413 (N_3413,In_1780,In_2170);
or U3414 (N_3414,In_1095,In_1260);
xor U3415 (N_3415,In_1810,In_1209);
xor U3416 (N_3416,In_1873,In_1780);
or U3417 (N_3417,In_913,In_943);
and U3418 (N_3418,In_2107,In_1035);
and U3419 (N_3419,In_316,In_417);
nand U3420 (N_3420,In_2012,In_1648);
and U3421 (N_3421,In_2408,In_114);
nor U3422 (N_3422,In_719,In_1229);
nand U3423 (N_3423,In_1518,In_2640);
nor U3424 (N_3424,In_342,In_2726);
nand U3425 (N_3425,In_844,In_974);
or U3426 (N_3426,In_941,In_1669);
nand U3427 (N_3427,In_1224,In_2595);
nand U3428 (N_3428,In_1807,In_1649);
nor U3429 (N_3429,In_1499,In_1193);
nor U3430 (N_3430,In_1121,In_572);
nand U3431 (N_3431,In_2027,In_530);
and U3432 (N_3432,In_925,In_2056);
nand U3433 (N_3433,In_2086,In_757);
or U3434 (N_3434,In_2512,In_12);
xor U3435 (N_3435,In_2704,In_2839);
xor U3436 (N_3436,In_1140,In_2182);
and U3437 (N_3437,In_497,In_1224);
xnor U3438 (N_3438,In_2098,In_389);
and U3439 (N_3439,In_806,In_2474);
nand U3440 (N_3440,In_836,In_2705);
xnor U3441 (N_3441,In_2446,In_2421);
nor U3442 (N_3442,In_501,In_1444);
nor U3443 (N_3443,In_840,In_640);
or U3444 (N_3444,In_890,In_2000);
nor U3445 (N_3445,In_2919,In_1613);
nand U3446 (N_3446,In_1396,In_157);
nor U3447 (N_3447,In_1699,In_2651);
nand U3448 (N_3448,In_2123,In_95);
or U3449 (N_3449,In_1973,In_2949);
nor U3450 (N_3450,In_1663,In_2255);
and U3451 (N_3451,In_602,In_1134);
and U3452 (N_3452,In_2161,In_941);
xor U3453 (N_3453,In_1017,In_2371);
and U3454 (N_3454,In_1233,In_1462);
nor U3455 (N_3455,In_2974,In_359);
or U3456 (N_3456,In_383,In_1802);
and U3457 (N_3457,In_139,In_662);
and U3458 (N_3458,In_1508,In_2902);
or U3459 (N_3459,In_1100,In_1433);
and U3460 (N_3460,In_2377,In_112);
or U3461 (N_3461,In_41,In_2430);
nand U3462 (N_3462,In_556,In_546);
nand U3463 (N_3463,In_602,In_1117);
nand U3464 (N_3464,In_717,In_1935);
and U3465 (N_3465,In_2249,In_1838);
or U3466 (N_3466,In_2288,In_526);
or U3467 (N_3467,In_171,In_914);
or U3468 (N_3468,In_2765,In_2159);
and U3469 (N_3469,In_2600,In_703);
or U3470 (N_3470,In_438,In_630);
xnor U3471 (N_3471,In_2503,In_1328);
nor U3472 (N_3472,In_1423,In_302);
xor U3473 (N_3473,In_505,In_161);
nand U3474 (N_3474,In_903,In_769);
and U3475 (N_3475,In_485,In_2336);
nor U3476 (N_3476,In_2422,In_2634);
or U3477 (N_3477,In_147,In_679);
nor U3478 (N_3478,In_1164,In_11);
or U3479 (N_3479,In_845,In_2832);
nor U3480 (N_3480,In_1279,In_2229);
nor U3481 (N_3481,In_1178,In_2213);
or U3482 (N_3482,In_402,In_2772);
xnor U3483 (N_3483,In_1217,In_65);
nor U3484 (N_3484,In_2104,In_2412);
xnor U3485 (N_3485,In_2303,In_1151);
and U3486 (N_3486,In_2169,In_1141);
nand U3487 (N_3487,In_972,In_1333);
nor U3488 (N_3488,In_562,In_1911);
or U3489 (N_3489,In_1924,In_1020);
nor U3490 (N_3490,In_2374,In_481);
xnor U3491 (N_3491,In_1314,In_494);
nor U3492 (N_3492,In_2711,In_1577);
and U3493 (N_3493,In_2490,In_390);
nor U3494 (N_3494,In_218,In_2160);
nand U3495 (N_3495,In_438,In_1453);
nand U3496 (N_3496,In_230,In_1263);
nand U3497 (N_3497,In_969,In_1342);
nor U3498 (N_3498,In_2750,In_1251);
and U3499 (N_3499,In_1422,In_2376);
or U3500 (N_3500,In_2079,In_552);
and U3501 (N_3501,In_1426,In_1270);
or U3502 (N_3502,In_2061,In_712);
or U3503 (N_3503,In_224,In_1140);
and U3504 (N_3504,In_2166,In_2283);
xnor U3505 (N_3505,In_1117,In_2663);
or U3506 (N_3506,In_2513,In_1928);
xnor U3507 (N_3507,In_1869,In_844);
and U3508 (N_3508,In_593,In_2091);
nor U3509 (N_3509,In_1404,In_882);
and U3510 (N_3510,In_1897,In_289);
and U3511 (N_3511,In_949,In_2354);
nor U3512 (N_3512,In_2532,In_1413);
nand U3513 (N_3513,In_2700,In_31);
nor U3514 (N_3514,In_2855,In_2495);
nor U3515 (N_3515,In_2855,In_2980);
nand U3516 (N_3516,In_165,In_2359);
nand U3517 (N_3517,In_2037,In_1661);
nor U3518 (N_3518,In_1607,In_255);
nand U3519 (N_3519,In_2679,In_551);
and U3520 (N_3520,In_1139,In_2724);
and U3521 (N_3521,In_695,In_1431);
nand U3522 (N_3522,In_120,In_842);
and U3523 (N_3523,In_1554,In_41);
and U3524 (N_3524,In_2143,In_307);
nand U3525 (N_3525,In_1694,In_2426);
and U3526 (N_3526,In_2012,In_292);
and U3527 (N_3527,In_2561,In_505);
nor U3528 (N_3528,In_2596,In_2223);
nand U3529 (N_3529,In_1640,In_902);
or U3530 (N_3530,In_51,In_2193);
or U3531 (N_3531,In_2156,In_599);
or U3532 (N_3532,In_1773,In_947);
nor U3533 (N_3533,In_2407,In_1639);
or U3534 (N_3534,In_2521,In_1338);
nor U3535 (N_3535,In_2881,In_2333);
or U3536 (N_3536,In_514,In_2641);
or U3537 (N_3537,In_2679,In_1806);
and U3538 (N_3538,In_2533,In_1579);
and U3539 (N_3539,In_207,In_1268);
nor U3540 (N_3540,In_2918,In_799);
or U3541 (N_3541,In_1963,In_82);
xor U3542 (N_3542,In_1873,In_827);
nand U3543 (N_3543,In_2589,In_188);
or U3544 (N_3544,In_427,In_402);
nor U3545 (N_3545,In_82,In_601);
nand U3546 (N_3546,In_2619,In_2080);
nand U3547 (N_3547,In_1949,In_2732);
and U3548 (N_3548,In_1420,In_724);
and U3549 (N_3549,In_486,In_2373);
nor U3550 (N_3550,In_2644,In_2641);
or U3551 (N_3551,In_572,In_575);
nor U3552 (N_3552,In_14,In_1687);
nand U3553 (N_3553,In_2911,In_901);
nor U3554 (N_3554,In_1834,In_2797);
and U3555 (N_3555,In_779,In_2725);
nand U3556 (N_3556,In_123,In_1962);
nand U3557 (N_3557,In_1077,In_2888);
and U3558 (N_3558,In_293,In_748);
and U3559 (N_3559,In_2196,In_764);
and U3560 (N_3560,In_718,In_2966);
or U3561 (N_3561,In_552,In_2349);
xor U3562 (N_3562,In_1306,In_2845);
or U3563 (N_3563,In_1188,In_2869);
nand U3564 (N_3564,In_2010,In_458);
and U3565 (N_3565,In_2940,In_515);
nor U3566 (N_3566,In_1850,In_2763);
nand U3567 (N_3567,In_2460,In_2635);
nand U3568 (N_3568,In_836,In_2464);
nand U3569 (N_3569,In_2719,In_1401);
or U3570 (N_3570,In_176,In_434);
nand U3571 (N_3571,In_1801,In_1279);
xor U3572 (N_3572,In_2552,In_24);
or U3573 (N_3573,In_216,In_2850);
nand U3574 (N_3574,In_2632,In_545);
nor U3575 (N_3575,In_1580,In_560);
nor U3576 (N_3576,In_867,In_764);
and U3577 (N_3577,In_1559,In_1068);
nor U3578 (N_3578,In_1533,In_579);
or U3579 (N_3579,In_881,In_333);
nor U3580 (N_3580,In_1073,In_654);
and U3581 (N_3581,In_1625,In_1611);
nor U3582 (N_3582,In_2489,In_2777);
and U3583 (N_3583,In_1190,In_1102);
or U3584 (N_3584,In_1122,In_2505);
nor U3585 (N_3585,In_2082,In_842);
and U3586 (N_3586,In_256,In_2114);
and U3587 (N_3587,In_1954,In_1243);
or U3588 (N_3588,In_2414,In_453);
or U3589 (N_3589,In_812,In_2593);
nand U3590 (N_3590,In_729,In_2712);
and U3591 (N_3591,In_1167,In_115);
nor U3592 (N_3592,In_2618,In_631);
nor U3593 (N_3593,In_917,In_2120);
nand U3594 (N_3594,In_1615,In_2297);
nand U3595 (N_3595,In_2022,In_2563);
nand U3596 (N_3596,In_2959,In_2301);
and U3597 (N_3597,In_1883,In_652);
nor U3598 (N_3598,In_483,In_2783);
nor U3599 (N_3599,In_2708,In_494);
nand U3600 (N_3600,In_2222,In_2622);
and U3601 (N_3601,In_2772,In_995);
nor U3602 (N_3602,In_163,In_883);
or U3603 (N_3603,In_95,In_1181);
nor U3604 (N_3604,In_467,In_1538);
and U3605 (N_3605,In_2342,In_1871);
xnor U3606 (N_3606,In_1330,In_1031);
nor U3607 (N_3607,In_1243,In_943);
and U3608 (N_3608,In_495,In_2364);
nor U3609 (N_3609,In_1678,In_151);
and U3610 (N_3610,In_2420,In_2073);
xnor U3611 (N_3611,In_2776,In_1480);
nand U3612 (N_3612,In_1103,In_776);
or U3613 (N_3613,In_1295,In_266);
xnor U3614 (N_3614,In_1520,In_2551);
or U3615 (N_3615,In_1825,In_201);
nor U3616 (N_3616,In_1338,In_1424);
and U3617 (N_3617,In_1046,In_1297);
xor U3618 (N_3618,In_1533,In_1877);
or U3619 (N_3619,In_1707,In_2288);
nor U3620 (N_3620,In_672,In_1288);
nor U3621 (N_3621,In_320,In_1378);
nand U3622 (N_3622,In_797,In_2870);
nor U3623 (N_3623,In_2875,In_2871);
or U3624 (N_3624,In_224,In_1835);
nand U3625 (N_3625,In_294,In_1000);
nand U3626 (N_3626,In_2164,In_2838);
xor U3627 (N_3627,In_2002,In_1209);
nor U3628 (N_3628,In_125,In_2839);
and U3629 (N_3629,In_2023,In_1749);
nor U3630 (N_3630,In_1566,In_2832);
or U3631 (N_3631,In_1442,In_1181);
xnor U3632 (N_3632,In_717,In_595);
and U3633 (N_3633,In_2941,In_2557);
xor U3634 (N_3634,In_220,In_733);
nor U3635 (N_3635,In_1203,In_1452);
nor U3636 (N_3636,In_2047,In_1692);
xor U3637 (N_3637,In_176,In_2528);
nor U3638 (N_3638,In_2025,In_2782);
or U3639 (N_3639,In_883,In_1146);
and U3640 (N_3640,In_1207,In_2238);
and U3641 (N_3641,In_181,In_2378);
nand U3642 (N_3642,In_1860,In_2687);
or U3643 (N_3643,In_1143,In_598);
nand U3644 (N_3644,In_2859,In_2695);
nand U3645 (N_3645,In_898,In_45);
nand U3646 (N_3646,In_1841,In_2623);
nor U3647 (N_3647,In_889,In_2772);
nor U3648 (N_3648,In_168,In_2073);
and U3649 (N_3649,In_2371,In_1084);
nand U3650 (N_3650,In_236,In_2083);
and U3651 (N_3651,In_96,In_459);
nand U3652 (N_3652,In_2587,In_1995);
nor U3653 (N_3653,In_944,In_2833);
xor U3654 (N_3654,In_2950,In_2981);
xor U3655 (N_3655,In_771,In_2295);
nand U3656 (N_3656,In_1769,In_47);
and U3657 (N_3657,In_2171,In_2671);
nand U3658 (N_3658,In_1626,In_503);
nor U3659 (N_3659,In_1432,In_826);
nor U3660 (N_3660,In_690,In_762);
nand U3661 (N_3661,In_2712,In_957);
nand U3662 (N_3662,In_2068,In_475);
and U3663 (N_3663,In_1835,In_2379);
or U3664 (N_3664,In_1489,In_453);
and U3665 (N_3665,In_153,In_2200);
and U3666 (N_3666,In_2448,In_1409);
nand U3667 (N_3667,In_61,In_1153);
or U3668 (N_3668,In_342,In_266);
nand U3669 (N_3669,In_1873,In_2340);
xnor U3670 (N_3670,In_2713,In_2903);
or U3671 (N_3671,In_2879,In_6);
nor U3672 (N_3672,In_298,In_481);
or U3673 (N_3673,In_1052,In_2612);
nor U3674 (N_3674,In_167,In_2813);
nor U3675 (N_3675,In_2677,In_1294);
and U3676 (N_3676,In_2852,In_2246);
or U3677 (N_3677,In_2013,In_2624);
or U3678 (N_3678,In_2373,In_438);
nor U3679 (N_3679,In_899,In_1476);
nand U3680 (N_3680,In_2578,In_2084);
nand U3681 (N_3681,In_481,In_889);
nor U3682 (N_3682,In_1018,In_957);
or U3683 (N_3683,In_293,In_604);
and U3684 (N_3684,In_194,In_1790);
or U3685 (N_3685,In_781,In_1937);
nor U3686 (N_3686,In_274,In_1883);
xnor U3687 (N_3687,In_300,In_1539);
and U3688 (N_3688,In_1346,In_977);
nor U3689 (N_3689,In_1322,In_1273);
and U3690 (N_3690,In_2838,In_1467);
or U3691 (N_3691,In_1202,In_1520);
and U3692 (N_3692,In_1356,In_1550);
and U3693 (N_3693,In_339,In_2606);
xnor U3694 (N_3694,In_2663,In_582);
nor U3695 (N_3695,In_2826,In_1102);
nor U3696 (N_3696,In_2511,In_2576);
nand U3697 (N_3697,In_97,In_2323);
nand U3698 (N_3698,In_353,In_2014);
nand U3699 (N_3699,In_2591,In_47);
and U3700 (N_3700,In_1255,In_326);
and U3701 (N_3701,In_2380,In_2562);
nand U3702 (N_3702,In_2311,In_2300);
nor U3703 (N_3703,In_2777,In_2591);
nor U3704 (N_3704,In_1895,In_2707);
or U3705 (N_3705,In_402,In_1827);
nor U3706 (N_3706,In_418,In_2787);
nor U3707 (N_3707,In_507,In_1427);
and U3708 (N_3708,In_1678,In_1517);
nand U3709 (N_3709,In_2627,In_2999);
or U3710 (N_3710,In_557,In_1138);
or U3711 (N_3711,In_523,In_2109);
and U3712 (N_3712,In_1336,In_2042);
xnor U3713 (N_3713,In_1589,In_825);
and U3714 (N_3714,In_895,In_2150);
nand U3715 (N_3715,In_2888,In_389);
nand U3716 (N_3716,In_1350,In_1056);
nand U3717 (N_3717,In_1215,In_230);
nand U3718 (N_3718,In_1240,In_186);
nor U3719 (N_3719,In_2094,In_325);
and U3720 (N_3720,In_653,In_274);
and U3721 (N_3721,In_1762,In_2397);
nand U3722 (N_3722,In_667,In_1036);
nor U3723 (N_3723,In_2313,In_2411);
nand U3724 (N_3724,In_2946,In_838);
nand U3725 (N_3725,In_2046,In_1437);
nor U3726 (N_3726,In_2520,In_2820);
nand U3727 (N_3727,In_296,In_1039);
xnor U3728 (N_3728,In_2403,In_1218);
xor U3729 (N_3729,In_1705,In_1413);
nand U3730 (N_3730,In_2051,In_1819);
nor U3731 (N_3731,In_635,In_333);
nor U3732 (N_3732,In_1109,In_2658);
nand U3733 (N_3733,In_140,In_787);
xnor U3734 (N_3734,In_1168,In_1929);
nand U3735 (N_3735,In_724,In_2494);
and U3736 (N_3736,In_1385,In_2141);
xor U3737 (N_3737,In_2921,In_244);
or U3738 (N_3738,In_1205,In_2985);
and U3739 (N_3739,In_959,In_2212);
xnor U3740 (N_3740,In_1316,In_513);
nand U3741 (N_3741,In_2215,In_1906);
nor U3742 (N_3742,In_1968,In_2214);
and U3743 (N_3743,In_187,In_1556);
nand U3744 (N_3744,In_2322,In_1035);
and U3745 (N_3745,In_2832,In_931);
nor U3746 (N_3746,In_2103,In_254);
nand U3747 (N_3747,In_142,In_2872);
and U3748 (N_3748,In_1544,In_2166);
or U3749 (N_3749,In_1093,In_2211);
nand U3750 (N_3750,In_825,In_2832);
and U3751 (N_3751,In_1621,In_59);
xor U3752 (N_3752,In_1295,In_360);
nor U3753 (N_3753,In_569,In_2946);
xnor U3754 (N_3754,In_1271,In_1574);
nand U3755 (N_3755,In_1862,In_2182);
and U3756 (N_3756,In_207,In_381);
or U3757 (N_3757,In_2324,In_2149);
nor U3758 (N_3758,In_2276,In_881);
or U3759 (N_3759,In_1134,In_876);
xor U3760 (N_3760,In_1285,In_2228);
nor U3761 (N_3761,In_760,In_2267);
and U3762 (N_3762,In_1563,In_354);
or U3763 (N_3763,In_204,In_261);
or U3764 (N_3764,In_2554,In_868);
and U3765 (N_3765,In_2905,In_1865);
xnor U3766 (N_3766,In_606,In_1045);
and U3767 (N_3767,In_192,In_902);
nor U3768 (N_3768,In_967,In_2322);
and U3769 (N_3769,In_2159,In_1451);
nor U3770 (N_3770,In_1264,In_1103);
nor U3771 (N_3771,In_1855,In_1820);
or U3772 (N_3772,In_1751,In_698);
or U3773 (N_3773,In_1825,In_2491);
nand U3774 (N_3774,In_114,In_2483);
or U3775 (N_3775,In_2261,In_1579);
or U3776 (N_3776,In_1259,In_2808);
xor U3777 (N_3777,In_1851,In_277);
xnor U3778 (N_3778,In_2779,In_1670);
nand U3779 (N_3779,In_2305,In_1927);
nor U3780 (N_3780,In_985,In_309);
xor U3781 (N_3781,In_2432,In_2024);
nor U3782 (N_3782,In_1990,In_1248);
or U3783 (N_3783,In_244,In_974);
and U3784 (N_3784,In_413,In_2036);
nor U3785 (N_3785,In_1570,In_2275);
and U3786 (N_3786,In_480,In_2535);
or U3787 (N_3787,In_851,In_956);
and U3788 (N_3788,In_1515,In_1985);
or U3789 (N_3789,In_451,In_311);
or U3790 (N_3790,In_2025,In_996);
or U3791 (N_3791,In_2385,In_1551);
or U3792 (N_3792,In_1661,In_377);
or U3793 (N_3793,In_776,In_1797);
nor U3794 (N_3794,In_2833,In_1870);
nand U3795 (N_3795,In_2548,In_2690);
and U3796 (N_3796,In_1616,In_2235);
or U3797 (N_3797,In_356,In_588);
nand U3798 (N_3798,In_2161,In_2224);
nand U3799 (N_3799,In_1541,In_1518);
nand U3800 (N_3800,In_164,In_1795);
nand U3801 (N_3801,In_1216,In_1108);
or U3802 (N_3802,In_2291,In_1727);
and U3803 (N_3803,In_782,In_1731);
or U3804 (N_3804,In_2359,In_1768);
or U3805 (N_3805,In_1587,In_2605);
or U3806 (N_3806,In_2353,In_2849);
nand U3807 (N_3807,In_949,In_705);
or U3808 (N_3808,In_1754,In_1460);
or U3809 (N_3809,In_198,In_847);
and U3810 (N_3810,In_2338,In_240);
xnor U3811 (N_3811,In_1944,In_2473);
nor U3812 (N_3812,In_92,In_1808);
nand U3813 (N_3813,In_2532,In_338);
or U3814 (N_3814,In_2545,In_1462);
nand U3815 (N_3815,In_1530,In_223);
nor U3816 (N_3816,In_2619,In_1326);
or U3817 (N_3817,In_177,In_551);
and U3818 (N_3818,In_2688,In_2642);
xnor U3819 (N_3819,In_1590,In_2142);
and U3820 (N_3820,In_168,In_2561);
or U3821 (N_3821,In_2213,In_1390);
and U3822 (N_3822,In_105,In_2488);
or U3823 (N_3823,In_1511,In_1591);
and U3824 (N_3824,In_2677,In_1648);
and U3825 (N_3825,In_2553,In_1180);
or U3826 (N_3826,In_1885,In_89);
nand U3827 (N_3827,In_2586,In_111);
and U3828 (N_3828,In_1493,In_795);
and U3829 (N_3829,In_2899,In_184);
or U3830 (N_3830,In_1601,In_1529);
and U3831 (N_3831,In_2037,In_2804);
and U3832 (N_3832,In_654,In_1418);
nor U3833 (N_3833,In_1176,In_352);
nand U3834 (N_3834,In_698,In_199);
nand U3835 (N_3835,In_438,In_856);
and U3836 (N_3836,In_1714,In_1117);
nand U3837 (N_3837,In_1721,In_365);
or U3838 (N_3838,In_82,In_2449);
nand U3839 (N_3839,In_1608,In_482);
nor U3840 (N_3840,In_1905,In_1163);
nand U3841 (N_3841,In_434,In_1632);
and U3842 (N_3842,In_425,In_2026);
nand U3843 (N_3843,In_312,In_2683);
nor U3844 (N_3844,In_1042,In_1543);
nand U3845 (N_3845,In_2846,In_1909);
xnor U3846 (N_3846,In_2164,In_557);
xor U3847 (N_3847,In_2433,In_131);
nor U3848 (N_3848,In_709,In_205);
nand U3849 (N_3849,In_511,In_1612);
or U3850 (N_3850,In_2207,In_726);
and U3851 (N_3851,In_13,In_1778);
nand U3852 (N_3852,In_1686,In_1330);
and U3853 (N_3853,In_117,In_2097);
nor U3854 (N_3854,In_1175,In_1126);
and U3855 (N_3855,In_1050,In_273);
and U3856 (N_3856,In_986,In_1858);
and U3857 (N_3857,In_1019,In_929);
and U3858 (N_3858,In_1647,In_2558);
and U3859 (N_3859,In_2643,In_20);
and U3860 (N_3860,In_236,In_2545);
nor U3861 (N_3861,In_1894,In_2000);
nor U3862 (N_3862,In_1437,In_1191);
nor U3863 (N_3863,In_2981,In_242);
nor U3864 (N_3864,In_467,In_2187);
nand U3865 (N_3865,In_1540,In_1622);
or U3866 (N_3866,In_586,In_2185);
nor U3867 (N_3867,In_495,In_1205);
or U3868 (N_3868,In_889,In_19);
xnor U3869 (N_3869,In_13,In_1924);
nor U3870 (N_3870,In_1642,In_2223);
nor U3871 (N_3871,In_2263,In_2447);
xnor U3872 (N_3872,In_2261,In_1846);
or U3873 (N_3873,In_1219,In_1080);
nor U3874 (N_3874,In_2917,In_2113);
or U3875 (N_3875,In_2523,In_1979);
nor U3876 (N_3876,In_1670,In_2533);
nand U3877 (N_3877,In_1203,In_640);
nand U3878 (N_3878,In_2066,In_132);
or U3879 (N_3879,In_631,In_2451);
or U3880 (N_3880,In_2505,In_684);
nor U3881 (N_3881,In_2889,In_1432);
and U3882 (N_3882,In_2957,In_899);
nor U3883 (N_3883,In_574,In_2453);
and U3884 (N_3884,In_2981,In_1435);
nand U3885 (N_3885,In_505,In_1767);
and U3886 (N_3886,In_378,In_1654);
nor U3887 (N_3887,In_1085,In_1755);
or U3888 (N_3888,In_1165,In_2457);
nand U3889 (N_3889,In_1030,In_794);
nand U3890 (N_3890,In_2410,In_2548);
or U3891 (N_3891,In_2844,In_75);
nor U3892 (N_3892,In_997,In_2548);
nand U3893 (N_3893,In_1637,In_1189);
or U3894 (N_3894,In_1751,In_2722);
or U3895 (N_3895,In_2420,In_2999);
and U3896 (N_3896,In_2029,In_186);
nor U3897 (N_3897,In_371,In_1467);
or U3898 (N_3898,In_893,In_1329);
or U3899 (N_3899,In_2295,In_694);
nor U3900 (N_3900,In_515,In_361);
and U3901 (N_3901,In_107,In_2221);
or U3902 (N_3902,In_2636,In_1427);
xnor U3903 (N_3903,In_2754,In_2829);
nor U3904 (N_3904,In_2446,In_1397);
or U3905 (N_3905,In_1087,In_1453);
or U3906 (N_3906,In_866,In_2247);
nand U3907 (N_3907,In_844,In_2349);
or U3908 (N_3908,In_2213,In_893);
and U3909 (N_3909,In_2638,In_1157);
nor U3910 (N_3910,In_702,In_1633);
and U3911 (N_3911,In_2193,In_516);
or U3912 (N_3912,In_2830,In_2664);
nor U3913 (N_3913,In_1286,In_448);
nand U3914 (N_3914,In_1220,In_103);
and U3915 (N_3915,In_1137,In_1712);
or U3916 (N_3916,In_2191,In_514);
and U3917 (N_3917,In_1728,In_2191);
nor U3918 (N_3918,In_878,In_1474);
or U3919 (N_3919,In_1046,In_695);
xnor U3920 (N_3920,In_2492,In_646);
nand U3921 (N_3921,In_1963,In_1739);
xnor U3922 (N_3922,In_904,In_1461);
and U3923 (N_3923,In_2142,In_1520);
nand U3924 (N_3924,In_2311,In_1216);
xor U3925 (N_3925,In_298,In_1031);
nand U3926 (N_3926,In_636,In_1617);
nor U3927 (N_3927,In_2133,In_2938);
xnor U3928 (N_3928,In_2560,In_2542);
nor U3929 (N_3929,In_2233,In_2687);
nand U3930 (N_3930,In_1664,In_62);
xnor U3931 (N_3931,In_2356,In_481);
or U3932 (N_3932,In_1600,In_2826);
or U3933 (N_3933,In_1328,In_690);
nor U3934 (N_3934,In_2539,In_12);
nor U3935 (N_3935,In_2723,In_1190);
nand U3936 (N_3936,In_2716,In_1591);
nand U3937 (N_3937,In_2920,In_89);
and U3938 (N_3938,In_2003,In_2444);
nand U3939 (N_3939,In_1773,In_1103);
and U3940 (N_3940,In_2518,In_1201);
or U3941 (N_3941,In_1328,In_402);
and U3942 (N_3942,In_2186,In_2236);
and U3943 (N_3943,In_1854,In_661);
or U3944 (N_3944,In_2020,In_1999);
or U3945 (N_3945,In_436,In_1979);
and U3946 (N_3946,In_939,In_2468);
nor U3947 (N_3947,In_2355,In_526);
nand U3948 (N_3948,In_1325,In_128);
nand U3949 (N_3949,In_1559,In_248);
and U3950 (N_3950,In_2433,In_1428);
nor U3951 (N_3951,In_2668,In_538);
nor U3952 (N_3952,In_1818,In_2302);
or U3953 (N_3953,In_666,In_1761);
nand U3954 (N_3954,In_744,In_1577);
nor U3955 (N_3955,In_852,In_2363);
and U3956 (N_3956,In_808,In_1551);
and U3957 (N_3957,In_1482,In_2220);
and U3958 (N_3958,In_1640,In_1366);
and U3959 (N_3959,In_1177,In_2523);
nand U3960 (N_3960,In_239,In_732);
xnor U3961 (N_3961,In_1509,In_82);
nand U3962 (N_3962,In_2725,In_2190);
and U3963 (N_3963,In_2928,In_2901);
and U3964 (N_3964,In_194,In_1850);
xnor U3965 (N_3965,In_627,In_1014);
nand U3966 (N_3966,In_988,In_1878);
xnor U3967 (N_3967,In_1376,In_134);
and U3968 (N_3968,In_298,In_1080);
or U3969 (N_3969,In_2282,In_1614);
nand U3970 (N_3970,In_2695,In_1497);
or U3971 (N_3971,In_63,In_1546);
nor U3972 (N_3972,In_76,In_1497);
or U3973 (N_3973,In_1094,In_1328);
xnor U3974 (N_3974,In_2422,In_2843);
or U3975 (N_3975,In_2441,In_2479);
nand U3976 (N_3976,In_1510,In_912);
nand U3977 (N_3977,In_239,In_776);
nand U3978 (N_3978,In_438,In_2269);
or U3979 (N_3979,In_2650,In_2510);
and U3980 (N_3980,In_288,In_508);
or U3981 (N_3981,In_677,In_688);
nand U3982 (N_3982,In_1212,In_2224);
and U3983 (N_3983,In_2216,In_774);
xor U3984 (N_3984,In_1613,In_354);
nand U3985 (N_3985,In_705,In_1083);
and U3986 (N_3986,In_375,In_2116);
and U3987 (N_3987,In_937,In_220);
nor U3988 (N_3988,In_2083,In_1930);
or U3989 (N_3989,In_2212,In_1420);
xnor U3990 (N_3990,In_2206,In_1924);
or U3991 (N_3991,In_1138,In_1069);
and U3992 (N_3992,In_1830,In_1193);
or U3993 (N_3993,In_424,In_103);
xnor U3994 (N_3994,In_1069,In_329);
nor U3995 (N_3995,In_2652,In_281);
and U3996 (N_3996,In_2158,In_196);
nor U3997 (N_3997,In_2534,In_2512);
and U3998 (N_3998,In_2016,In_2105);
nand U3999 (N_3999,In_1705,In_409);
and U4000 (N_4000,In_2867,In_2063);
and U4001 (N_4001,In_2650,In_1489);
and U4002 (N_4002,In_2499,In_622);
xnor U4003 (N_4003,In_13,In_2297);
nand U4004 (N_4004,In_1058,In_421);
nor U4005 (N_4005,In_1153,In_1571);
nor U4006 (N_4006,In_106,In_588);
or U4007 (N_4007,In_542,In_1523);
or U4008 (N_4008,In_847,In_2363);
nor U4009 (N_4009,In_2326,In_627);
nand U4010 (N_4010,In_938,In_1265);
nand U4011 (N_4011,In_525,In_231);
nor U4012 (N_4012,In_2761,In_527);
nor U4013 (N_4013,In_2488,In_546);
and U4014 (N_4014,In_2228,In_1579);
and U4015 (N_4015,In_374,In_838);
and U4016 (N_4016,In_2319,In_2404);
and U4017 (N_4017,In_786,In_354);
nand U4018 (N_4018,In_2272,In_385);
nor U4019 (N_4019,In_1542,In_1109);
or U4020 (N_4020,In_1879,In_409);
nor U4021 (N_4021,In_1915,In_2367);
and U4022 (N_4022,In_1303,In_397);
and U4023 (N_4023,In_654,In_2911);
and U4024 (N_4024,In_1250,In_721);
nor U4025 (N_4025,In_1450,In_1011);
nor U4026 (N_4026,In_853,In_54);
or U4027 (N_4027,In_539,In_1512);
nor U4028 (N_4028,In_1474,In_1877);
and U4029 (N_4029,In_2363,In_1160);
nand U4030 (N_4030,In_2091,In_1355);
and U4031 (N_4031,In_1810,In_2359);
or U4032 (N_4032,In_1925,In_1744);
or U4033 (N_4033,In_452,In_1516);
or U4034 (N_4034,In_547,In_1607);
nor U4035 (N_4035,In_739,In_479);
nor U4036 (N_4036,In_2994,In_1762);
nand U4037 (N_4037,In_2451,In_2537);
and U4038 (N_4038,In_2778,In_2679);
nor U4039 (N_4039,In_1637,In_645);
nand U4040 (N_4040,In_2433,In_1604);
or U4041 (N_4041,In_886,In_632);
nor U4042 (N_4042,In_309,In_1439);
or U4043 (N_4043,In_890,In_2120);
xnor U4044 (N_4044,In_581,In_375);
nor U4045 (N_4045,In_1618,In_544);
nand U4046 (N_4046,In_98,In_2253);
or U4047 (N_4047,In_223,In_1620);
nor U4048 (N_4048,In_2470,In_1413);
nand U4049 (N_4049,In_210,In_1315);
and U4050 (N_4050,In_1377,In_1892);
and U4051 (N_4051,In_1971,In_701);
nor U4052 (N_4052,In_2072,In_1058);
xor U4053 (N_4053,In_1149,In_1363);
xor U4054 (N_4054,In_676,In_1485);
or U4055 (N_4055,In_2861,In_2944);
and U4056 (N_4056,In_617,In_769);
nand U4057 (N_4057,In_1141,In_1437);
or U4058 (N_4058,In_544,In_739);
and U4059 (N_4059,In_919,In_333);
nand U4060 (N_4060,In_1507,In_2527);
nor U4061 (N_4061,In_1121,In_2271);
and U4062 (N_4062,In_227,In_2415);
xnor U4063 (N_4063,In_2343,In_2690);
or U4064 (N_4064,In_1455,In_2765);
xnor U4065 (N_4065,In_13,In_2411);
nand U4066 (N_4066,In_2614,In_1128);
and U4067 (N_4067,In_2822,In_2544);
or U4068 (N_4068,In_111,In_381);
nand U4069 (N_4069,In_1338,In_455);
nand U4070 (N_4070,In_974,In_1974);
nor U4071 (N_4071,In_1962,In_14);
and U4072 (N_4072,In_932,In_1122);
nand U4073 (N_4073,In_408,In_2460);
nor U4074 (N_4074,In_278,In_1145);
or U4075 (N_4075,In_1700,In_852);
or U4076 (N_4076,In_501,In_2196);
nand U4077 (N_4077,In_549,In_1293);
xnor U4078 (N_4078,In_2318,In_1225);
nand U4079 (N_4079,In_1705,In_25);
nand U4080 (N_4080,In_1634,In_2596);
and U4081 (N_4081,In_1880,In_144);
and U4082 (N_4082,In_2334,In_2721);
and U4083 (N_4083,In_1765,In_2436);
nand U4084 (N_4084,In_1453,In_1194);
nor U4085 (N_4085,In_657,In_2394);
nor U4086 (N_4086,In_2700,In_194);
nor U4087 (N_4087,In_841,In_781);
nor U4088 (N_4088,In_1646,In_833);
and U4089 (N_4089,In_482,In_404);
and U4090 (N_4090,In_2405,In_2582);
nand U4091 (N_4091,In_50,In_459);
and U4092 (N_4092,In_2357,In_2941);
xnor U4093 (N_4093,In_1473,In_1456);
and U4094 (N_4094,In_2283,In_2031);
and U4095 (N_4095,In_1088,In_450);
nor U4096 (N_4096,In_1914,In_1356);
or U4097 (N_4097,In_1947,In_1958);
nor U4098 (N_4098,In_2110,In_1238);
and U4099 (N_4099,In_2835,In_2684);
xor U4100 (N_4100,In_367,In_2835);
nand U4101 (N_4101,In_2925,In_1449);
or U4102 (N_4102,In_2742,In_2719);
nor U4103 (N_4103,In_706,In_532);
nand U4104 (N_4104,In_2792,In_950);
nand U4105 (N_4105,In_1270,In_2524);
xor U4106 (N_4106,In_2041,In_1045);
or U4107 (N_4107,In_1245,In_174);
nand U4108 (N_4108,In_249,In_2016);
nor U4109 (N_4109,In_2053,In_182);
or U4110 (N_4110,In_2618,In_1695);
and U4111 (N_4111,In_1783,In_1722);
nand U4112 (N_4112,In_2175,In_1739);
nand U4113 (N_4113,In_1844,In_2503);
nor U4114 (N_4114,In_325,In_1394);
nor U4115 (N_4115,In_1485,In_2276);
or U4116 (N_4116,In_2251,In_2056);
nor U4117 (N_4117,In_399,In_2422);
nand U4118 (N_4118,In_1327,In_1934);
nor U4119 (N_4119,In_2158,In_2323);
nor U4120 (N_4120,In_2875,In_544);
xor U4121 (N_4121,In_27,In_2466);
and U4122 (N_4122,In_2671,In_2497);
or U4123 (N_4123,In_105,In_1101);
xor U4124 (N_4124,In_56,In_1139);
and U4125 (N_4125,In_1192,In_476);
and U4126 (N_4126,In_1584,In_331);
or U4127 (N_4127,In_849,In_929);
and U4128 (N_4128,In_2340,In_2633);
nand U4129 (N_4129,In_2002,In_2183);
or U4130 (N_4130,In_2746,In_1410);
and U4131 (N_4131,In_587,In_2706);
xnor U4132 (N_4132,In_1722,In_1320);
nand U4133 (N_4133,In_1861,In_632);
or U4134 (N_4134,In_2524,In_128);
nand U4135 (N_4135,In_2658,In_2515);
and U4136 (N_4136,In_2457,In_1254);
and U4137 (N_4137,In_87,In_1423);
and U4138 (N_4138,In_483,In_2314);
or U4139 (N_4139,In_1171,In_1262);
nor U4140 (N_4140,In_2868,In_2020);
and U4141 (N_4141,In_693,In_2675);
xnor U4142 (N_4142,In_871,In_2862);
xnor U4143 (N_4143,In_1889,In_1883);
and U4144 (N_4144,In_379,In_2565);
or U4145 (N_4145,In_1479,In_2114);
xnor U4146 (N_4146,In_2638,In_1998);
nor U4147 (N_4147,In_420,In_1913);
nor U4148 (N_4148,In_859,In_2137);
xor U4149 (N_4149,In_1810,In_1159);
nand U4150 (N_4150,In_1431,In_2165);
and U4151 (N_4151,In_1499,In_2538);
nor U4152 (N_4152,In_2282,In_1548);
nand U4153 (N_4153,In_550,In_1175);
and U4154 (N_4154,In_2206,In_2707);
nand U4155 (N_4155,In_2344,In_886);
nor U4156 (N_4156,In_417,In_971);
or U4157 (N_4157,In_2071,In_2294);
nand U4158 (N_4158,In_999,In_2814);
or U4159 (N_4159,In_2055,In_1806);
nand U4160 (N_4160,In_776,In_176);
nor U4161 (N_4161,In_1201,In_1387);
nand U4162 (N_4162,In_511,In_1406);
nand U4163 (N_4163,In_921,In_912);
or U4164 (N_4164,In_342,In_1258);
nor U4165 (N_4165,In_500,In_1275);
and U4166 (N_4166,In_881,In_2985);
nand U4167 (N_4167,In_1378,In_2645);
and U4168 (N_4168,In_104,In_657);
nand U4169 (N_4169,In_2784,In_2895);
or U4170 (N_4170,In_1379,In_1357);
nor U4171 (N_4171,In_2335,In_2212);
nor U4172 (N_4172,In_190,In_1322);
nor U4173 (N_4173,In_2943,In_949);
nand U4174 (N_4174,In_2841,In_1481);
xor U4175 (N_4175,In_843,In_1088);
nor U4176 (N_4176,In_738,In_2047);
and U4177 (N_4177,In_2414,In_436);
nor U4178 (N_4178,In_787,In_1397);
and U4179 (N_4179,In_768,In_1789);
nor U4180 (N_4180,In_2177,In_2712);
or U4181 (N_4181,In_2887,In_1660);
nand U4182 (N_4182,In_202,In_1332);
nor U4183 (N_4183,In_1420,In_585);
nand U4184 (N_4184,In_1936,In_1200);
and U4185 (N_4185,In_624,In_674);
and U4186 (N_4186,In_2022,In_2259);
nor U4187 (N_4187,In_1868,In_860);
and U4188 (N_4188,In_2476,In_959);
or U4189 (N_4189,In_293,In_1246);
or U4190 (N_4190,In_900,In_1333);
or U4191 (N_4191,In_883,In_62);
or U4192 (N_4192,In_1069,In_1638);
xnor U4193 (N_4193,In_1884,In_2636);
nor U4194 (N_4194,In_208,In_1212);
or U4195 (N_4195,In_527,In_966);
and U4196 (N_4196,In_1885,In_1526);
xor U4197 (N_4197,In_1358,In_1480);
nor U4198 (N_4198,In_0,In_2612);
and U4199 (N_4199,In_1887,In_120);
nand U4200 (N_4200,In_2789,In_880);
or U4201 (N_4201,In_2721,In_2799);
nand U4202 (N_4202,In_2122,In_333);
and U4203 (N_4203,In_2955,In_2316);
and U4204 (N_4204,In_1335,In_2236);
nor U4205 (N_4205,In_875,In_732);
and U4206 (N_4206,In_2820,In_1714);
or U4207 (N_4207,In_1300,In_2102);
nand U4208 (N_4208,In_942,In_2049);
nand U4209 (N_4209,In_1640,In_2516);
xnor U4210 (N_4210,In_95,In_2060);
xnor U4211 (N_4211,In_2724,In_1461);
nor U4212 (N_4212,In_1064,In_2866);
xnor U4213 (N_4213,In_1195,In_1797);
nand U4214 (N_4214,In_622,In_1886);
nor U4215 (N_4215,In_837,In_1951);
nor U4216 (N_4216,In_1776,In_359);
nor U4217 (N_4217,In_1528,In_2540);
nor U4218 (N_4218,In_2779,In_1931);
nor U4219 (N_4219,In_2810,In_1400);
and U4220 (N_4220,In_2547,In_2647);
nand U4221 (N_4221,In_1328,In_1901);
nor U4222 (N_4222,In_1978,In_1787);
xor U4223 (N_4223,In_2583,In_2373);
or U4224 (N_4224,In_2020,In_1176);
and U4225 (N_4225,In_221,In_1773);
xor U4226 (N_4226,In_1262,In_1983);
nand U4227 (N_4227,In_1777,In_2866);
nor U4228 (N_4228,In_584,In_118);
and U4229 (N_4229,In_223,In_1624);
and U4230 (N_4230,In_2086,In_1968);
nor U4231 (N_4231,In_136,In_328);
nand U4232 (N_4232,In_2141,In_2174);
or U4233 (N_4233,In_650,In_696);
nand U4234 (N_4234,In_129,In_2763);
nand U4235 (N_4235,In_794,In_1438);
or U4236 (N_4236,In_190,In_245);
nand U4237 (N_4237,In_849,In_173);
and U4238 (N_4238,In_2067,In_46);
nor U4239 (N_4239,In_2341,In_1482);
nor U4240 (N_4240,In_2417,In_837);
or U4241 (N_4241,In_2141,In_2211);
or U4242 (N_4242,In_2929,In_2882);
or U4243 (N_4243,In_1093,In_2356);
and U4244 (N_4244,In_2254,In_2219);
nor U4245 (N_4245,In_217,In_634);
or U4246 (N_4246,In_664,In_2575);
xnor U4247 (N_4247,In_2700,In_1558);
xor U4248 (N_4248,In_949,In_1683);
nor U4249 (N_4249,In_2712,In_348);
nand U4250 (N_4250,In_2328,In_1111);
nor U4251 (N_4251,In_1789,In_358);
or U4252 (N_4252,In_2212,In_893);
or U4253 (N_4253,In_10,In_1170);
nand U4254 (N_4254,In_1854,In_1563);
and U4255 (N_4255,In_1503,In_940);
nor U4256 (N_4256,In_621,In_995);
or U4257 (N_4257,In_281,In_2585);
nand U4258 (N_4258,In_1914,In_1930);
or U4259 (N_4259,In_1384,In_109);
nand U4260 (N_4260,In_206,In_2301);
and U4261 (N_4261,In_1784,In_1946);
or U4262 (N_4262,In_778,In_645);
nand U4263 (N_4263,In_1005,In_1799);
or U4264 (N_4264,In_1581,In_2178);
nor U4265 (N_4265,In_956,In_1712);
nor U4266 (N_4266,In_282,In_2887);
nor U4267 (N_4267,In_739,In_1618);
nand U4268 (N_4268,In_1178,In_859);
and U4269 (N_4269,In_976,In_1965);
xor U4270 (N_4270,In_1812,In_71);
and U4271 (N_4271,In_929,In_2174);
nor U4272 (N_4272,In_368,In_2176);
nor U4273 (N_4273,In_1562,In_17);
or U4274 (N_4274,In_2846,In_1508);
or U4275 (N_4275,In_2070,In_2054);
nor U4276 (N_4276,In_1605,In_2956);
nand U4277 (N_4277,In_420,In_1158);
and U4278 (N_4278,In_447,In_1010);
nor U4279 (N_4279,In_781,In_304);
or U4280 (N_4280,In_2648,In_64);
nand U4281 (N_4281,In_316,In_2246);
nor U4282 (N_4282,In_1474,In_2996);
and U4283 (N_4283,In_260,In_2754);
and U4284 (N_4284,In_519,In_1373);
or U4285 (N_4285,In_1108,In_1638);
nand U4286 (N_4286,In_1755,In_1);
and U4287 (N_4287,In_518,In_2451);
nand U4288 (N_4288,In_477,In_493);
and U4289 (N_4289,In_452,In_346);
nor U4290 (N_4290,In_1803,In_565);
nand U4291 (N_4291,In_2414,In_2388);
nor U4292 (N_4292,In_971,In_1793);
xor U4293 (N_4293,In_2257,In_2820);
nand U4294 (N_4294,In_80,In_1715);
nand U4295 (N_4295,In_1146,In_539);
and U4296 (N_4296,In_2891,In_1488);
nand U4297 (N_4297,In_3,In_497);
nand U4298 (N_4298,In_2292,In_2064);
and U4299 (N_4299,In_2348,In_594);
and U4300 (N_4300,In_1176,In_685);
and U4301 (N_4301,In_619,In_2960);
or U4302 (N_4302,In_2720,In_1204);
nor U4303 (N_4303,In_1465,In_1684);
nand U4304 (N_4304,In_923,In_426);
nor U4305 (N_4305,In_403,In_1819);
or U4306 (N_4306,In_2446,In_707);
nand U4307 (N_4307,In_1579,In_2514);
xor U4308 (N_4308,In_1860,In_1053);
and U4309 (N_4309,In_2804,In_658);
and U4310 (N_4310,In_2722,In_2255);
or U4311 (N_4311,In_644,In_2543);
or U4312 (N_4312,In_2010,In_1533);
nor U4313 (N_4313,In_529,In_214);
nor U4314 (N_4314,In_754,In_1978);
or U4315 (N_4315,In_2917,In_16);
or U4316 (N_4316,In_972,In_311);
or U4317 (N_4317,In_826,In_2507);
nor U4318 (N_4318,In_2768,In_2856);
or U4319 (N_4319,In_2593,In_1136);
and U4320 (N_4320,In_1401,In_458);
nand U4321 (N_4321,In_1932,In_2046);
or U4322 (N_4322,In_102,In_1651);
or U4323 (N_4323,In_2152,In_461);
nor U4324 (N_4324,In_147,In_1565);
and U4325 (N_4325,In_1508,In_2187);
nor U4326 (N_4326,In_2916,In_2769);
or U4327 (N_4327,In_1167,In_2524);
nand U4328 (N_4328,In_2340,In_880);
nor U4329 (N_4329,In_1334,In_369);
nor U4330 (N_4330,In_2983,In_2817);
or U4331 (N_4331,In_1053,In_969);
nor U4332 (N_4332,In_2625,In_1270);
nand U4333 (N_4333,In_457,In_2490);
xnor U4334 (N_4334,In_1731,In_396);
and U4335 (N_4335,In_2645,In_2271);
nor U4336 (N_4336,In_832,In_1269);
or U4337 (N_4337,In_633,In_1888);
or U4338 (N_4338,In_244,In_563);
and U4339 (N_4339,In_2091,In_2223);
nor U4340 (N_4340,In_446,In_2367);
nor U4341 (N_4341,In_1713,In_779);
or U4342 (N_4342,In_2918,In_217);
nand U4343 (N_4343,In_816,In_2062);
or U4344 (N_4344,In_1884,In_556);
nand U4345 (N_4345,In_939,In_1570);
and U4346 (N_4346,In_2269,In_761);
or U4347 (N_4347,In_22,In_330);
or U4348 (N_4348,In_1392,In_281);
xor U4349 (N_4349,In_2732,In_2447);
nor U4350 (N_4350,In_2357,In_825);
or U4351 (N_4351,In_940,In_297);
nand U4352 (N_4352,In_2668,In_571);
or U4353 (N_4353,In_1007,In_328);
and U4354 (N_4354,In_2926,In_2756);
nand U4355 (N_4355,In_1178,In_2542);
nor U4356 (N_4356,In_2068,In_2178);
nand U4357 (N_4357,In_1302,In_1974);
or U4358 (N_4358,In_1996,In_2323);
nor U4359 (N_4359,In_1864,In_1196);
nand U4360 (N_4360,In_1681,In_2328);
nor U4361 (N_4361,In_987,In_1689);
nor U4362 (N_4362,In_386,In_2912);
xnor U4363 (N_4363,In_2528,In_1604);
nand U4364 (N_4364,In_1537,In_440);
nor U4365 (N_4365,In_1873,In_2328);
and U4366 (N_4366,In_441,In_2236);
or U4367 (N_4367,In_554,In_444);
nand U4368 (N_4368,In_951,In_2915);
or U4369 (N_4369,In_1866,In_1389);
nand U4370 (N_4370,In_1750,In_1811);
and U4371 (N_4371,In_113,In_402);
and U4372 (N_4372,In_1913,In_2546);
and U4373 (N_4373,In_1635,In_135);
or U4374 (N_4374,In_1102,In_2179);
or U4375 (N_4375,In_1369,In_2466);
and U4376 (N_4376,In_333,In_2993);
nand U4377 (N_4377,In_1072,In_338);
nor U4378 (N_4378,In_2150,In_314);
and U4379 (N_4379,In_2205,In_1546);
and U4380 (N_4380,In_2713,In_2128);
and U4381 (N_4381,In_1864,In_2287);
or U4382 (N_4382,In_2877,In_287);
nor U4383 (N_4383,In_876,In_36);
or U4384 (N_4384,In_2925,In_2725);
nor U4385 (N_4385,In_9,In_1944);
nor U4386 (N_4386,In_2597,In_39);
nor U4387 (N_4387,In_431,In_2297);
nand U4388 (N_4388,In_954,In_2457);
or U4389 (N_4389,In_2192,In_286);
nor U4390 (N_4390,In_264,In_1685);
xnor U4391 (N_4391,In_510,In_59);
and U4392 (N_4392,In_1172,In_2690);
and U4393 (N_4393,In_1531,In_245);
and U4394 (N_4394,In_266,In_2911);
nand U4395 (N_4395,In_144,In_1517);
nor U4396 (N_4396,In_1783,In_2375);
and U4397 (N_4397,In_2539,In_311);
and U4398 (N_4398,In_988,In_2257);
xor U4399 (N_4399,In_266,In_1068);
nand U4400 (N_4400,In_1629,In_585);
nor U4401 (N_4401,In_1074,In_2837);
nand U4402 (N_4402,In_590,In_133);
or U4403 (N_4403,In_1539,In_2061);
and U4404 (N_4404,In_2513,In_896);
and U4405 (N_4405,In_680,In_1380);
xnor U4406 (N_4406,In_1581,In_448);
nand U4407 (N_4407,In_2968,In_2928);
or U4408 (N_4408,In_1571,In_1626);
or U4409 (N_4409,In_2892,In_957);
nand U4410 (N_4410,In_924,In_2817);
nor U4411 (N_4411,In_2829,In_753);
and U4412 (N_4412,In_2496,In_2788);
nor U4413 (N_4413,In_1664,In_314);
or U4414 (N_4414,In_566,In_1759);
or U4415 (N_4415,In_1373,In_716);
nand U4416 (N_4416,In_1963,In_1777);
xnor U4417 (N_4417,In_1254,In_451);
nand U4418 (N_4418,In_1771,In_679);
nand U4419 (N_4419,In_1321,In_342);
nand U4420 (N_4420,In_2378,In_2531);
nand U4421 (N_4421,In_1517,In_2933);
and U4422 (N_4422,In_109,In_735);
nand U4423 (N_4423,In_2704,In_2209);
and U4424 (N_4424,In_2111,In_993);
or U4425 (N_4425,In_1102,In_115);
nor U4426 (N_4426,In_2278,In_1051);
and U4427 (N_4427,In_78,In_176);
or U4428 (N_4428,In_2247,In_2175);
nor U4429 (N_4429,In_1668,In_2218);
or U4430 (N_4430,In_2298,In_202);
and U4431 (N_4431,In_2107,In_2908);
or U4432 (N_4432,In_724,In_1041);
or U4433 (N_4433,In_2649,In_99);
xnor U4434 (N_4434,In_2827,In_1753);
nand U4435 (N_4435,In_2942,In_739);
and U4436 (N_4436,In_2851,In_1488);
nand U4437 (N_4437,In_1904,In_2518);
or U4438 (N_4438,In_1415,In_2171);
nand U4439 (N_4439,In_1479,In_2417);
nor U4440 (N_4440,In_2274,In_1070);
nand U4441 (N_4441,In_2953,In_2166);
or U4442 (N_4442,In_782,In_2709);
xnor U4443 (N_4443,In_115,In_2242);
nand U4444 (N_4444,In_2766,In_2584);
nor U4445 (N_4445,In_168,In_2407);
or U4446 (N_4446,In_1158,In_165);
and U4447 (N_4447,In_1036,In_717);
or U4448 (N_4448,In_105,In_370);
and U4449 (N_4449,In_1191,In_322);
and U4450 (N_4450,In_1285,In_1443);
and U4451 (N_4451,In_2630,In_2237);
or U4452 (N_4452,In_2971,In_1165);
nor U4453 (N_4453,In_1504,In_1246);
nand U4454 (N_4454,In_1262,In_1945);
xnor U4455 (N_4455,In_55,In_187);
nand U4456 (N_4456,In_981,In_2684);
or U4457 (N_4457,In_801,In_1874);
nand U4458 (N_4458,In_962,In_349);
and U4459 (N_4459,In_2947,In_192);
xnor U4460 (N_4460,In_2499,In_1209);
or U4461 (N_4461,In_384,In_1613);
or U4462 (N_4462,In_298,In_1538);
nand U4463 (N_4463,In_1939,In_331);
nand U4464 (N_4464,In_651,In_363);
nand U4465 (N_4465,In_960,In_125);
or U4466 (N_4466,In_2208,In_2886);
and U4467 (N_4467,In_835,In_2965);
or U4468 (N_4468,In_1493,In_2477);
nor U4469 (N_4469,In_743,In_1387);
and U4470 (N_4470,In_2344,In_1401);
nor U4471 (N_4471,In_1509,In_2887);
or U4472 (N_4472,In_2577,In_2658);
or U4473 (N_4473,In_2087,In_939);
and U4474 (N_4474,In_1686,In_1941);
nor U4475 (N_4475,In_1837,In_1397);
and U4476 (N_4476,In_445,In_1622);
or U4477 (N_4477,In_1210,In_2039);
nand U4478 (N_4478,In_708,In_2381);
xor U4479 (N_4479,In_747,In_2777);
nor U4480 (N_4480,In_2802,In_2054);
nand U4481 (N_4481,In_601,In_1149);
nand U4482 (N_4482,In_983,In_2921);
and U4483 (N_4483,In_1173,In_2981);
and U4484 (N_4484,In_2576,In_624);
nor U4485 (N_4485,In_1791,In_932);
and U4486 (N_4486,In_1235,In_1145);
or U4487 (N_4487,In_634,In_272);
nor U4488 (N_4488,In_2462,In_139);
or U4489 (N_4489,In_763,In_1329);
nand U4490 (N_4490,In_1606,In_714);
nand U4491 (N_4491,In_264,In_1050);
and U4492 (N_4492,In_2429,In_2701);
or U4493 (N_4493,In_979,In_2334);
and U4494 (N_4494,In_396,In_1173);
or U4495 (N_4495,In_1318,In_0);
and U4496 (N_4496,In_577,In_1336);
nor U4497 (N_4497,In_906,In_1263);
nand U4498 (N_4498,In_2155,In_1994);
or U4499 (N_4499,In_2317,In_1962);
and U4500 (N_4500,In_731,In_1478);
nand U4501 (N_4501,In_2230,In_1166);
and U4502 (N_4502,In_2109,In_1445);
and U4503 (N_4503,In_789,In_931);
xor U4504 (N_4504,In_1460,In_1070);
and U4505 (N_4505,In_2197,In_1409);
or U4506 (N_4506,In_762,In_2639);
xor U4507 (N_4507,In_2666,In_19);
nand U4508 (N_4508,In_2013,In_1711);
or U4509 (N_4509,In_2542,In_2387);
and U4510 (N_4510,In_491,In_113);
nand U4511 (N_4511,In_2896,In_2002);
nor U4512 (N_4512,In_140,In_1135);
nor U4513 (N_4513,In_622,In_2829);
nor U4514 (N_4514,In_463,In_2161);
nand U4515 (N_4515,In_1017,In_1957);
and U4516 (N_4516,In_1345,In_238);
and U4517 (N_4517,In_250,In_701);
and U4518 (N_4518,In_2179,In_609);
nand U4519 (N_4519,In_1631,In_1125);
and U4520 (N_4520,In_1,In_475);
or U4521 (N_4521,In_1928,In_785);
nand U4522 (N_4522,In_2618,In_1018);
nor U4523 (N_4523,In_555,In_763);
nor U4524 (N_4524,In_2099,In_2379);
xnor U4525 (N_4525,In_2695,In_959);
and U4526 (N_4526,In_2940,In_199);
nor U4527 (N_4527,In_395,In_221);
and U4528 (N_4528,In_1297,In_2235);
and U4529 (N_4529,In_2555,In_1918);
xnor U4530 (N_4530,In_2064,In_2897);
nor U4531 (N_4531,In_1223,In_1726);
nand U4532 (N_4532,In_585,In_1840);
or U4533 (N_4533,In_370,In_2267);
nand U4534 (N_4534,In_149,In_1794);
and U4535 (N_4535,In_2959,In_1909);
and U4536 (N_4536,In_1972,In_1476);
nor U4537 (N_4537,In_2253,In_2603);
xor U4538 (N_4538,In_160,In_1605);
and U4539 (N_4539,In_401,In_1062);
or U4540 (N_4540,In_1207,In_21);
and U4541 (N_4541,In_1409,In_356);
or U4542 (N_4542,In_1361,In_163);
nand U4543 (N_4543,In_1718,In_312);
nand U4544 (N_4544,In_654,In_1812);
xnor U4545 (N_4545,In_2187,In_1131);
or U4546 (N_4546,In_1891,In_2557);
or U4547 (N_4547,In_2626,In_1469);
nand U4548 (N_4548,In_2435,In_2378);
and U4549 (N_4549,In_1893,In_91);
or U4550 (N_4550,In_2461,In_329);
or U4551 (N_4551,In_1175,In_2957);
or U4552 (N_4552,In_300,In_2195);
nand U4553 (N_4553,In_2026,In_373);
or U4554 (N_4554,In_1291,In_2686);
or U4555 (N_4555,In_2262,In_1162);
nand U4556 (N_4556,In_2742,In_2975);
and U4557 (N_4557,In_2000,In_2596);
and U4558 (N_4558,In_2643,In_2215);
and U4559 (N_4559,In_2512,In_1472);
and U4560 (N_4560,In_428,In_811);
nand U4561 (N_4561,In_1536,In_2426);
and U4562 (N_4562,In_2798,In_288);
xnor U4563 (N_4563,In_863,In_43);
and U4564 (N_4564,In_1141,In_2634);
and U4565 (N_4565,In_1859,In_2483);
or U4566 (N_4566,In_2548,In_860);
or U4567 (N_4567,In_2263,In_2178);
xor U4568 (N_4568,In_2456,In_403);
or U4569 (N_4569,In_1065,In_739);
nor U4570 (N_4570,In_1922,In_2898);
or U4571 (N_4571,In_2278,In_623);
nor U4572 (N_4572,In_2228,In_2161);
nor U4573 (N_4573,In_1809,In_1272);
and U4574 (N_4574,In_533,In_48);
nand U4575 (N_4575,In_2860,In_2574);
or U4576 (N_4576,In_145,In_2647);
nand U4577 (N_4577,In_2764,In_2214);
nor U4578 (N_4578,In_16,In_2890);
nor U4579 (N_4579,In_1431,In_1522);
or U4580 (N_4580,In_2120,In_57);
or U4581 (N_4581,In_1929,In_2301);
or U4582 (N_4582,In_2941,In_2174);
nor U4583 (N_4583,In_827,In_2598);
or U4584 (N_4584,In_2787,In_791);
or U4585 (N_4585,In_2063,In_1313);
nor U4586 (N_4586,In_1400,In_2988);
or U4587 (N_4587,In_2208,In_2738);
nor U4588 (N_4588,In_667,In_833);
nand U4589 (N_4589,In_2310,In_2000);
and U4590 (N_4590,In_2124,In_2938);
or U4591 (N_4591,In_488,In_1869);
nand U4592 (N_4592,In_1335,In_20);
nand U4593 (N_4593,In_1768,In_51);
nand U4594 (N_4594,In_1058,In_285);
nand U4595 (N_4595,In_966,In_585);
or U4596 (N_4596,In_459,In_2844);
and U4597 (N_4597,In_2058,In_154);
and U4598 (N_4598,In_1103,In_259);
nor U4599 (N_4599,In_1073,In_1076);
and U4600 (N_4600,In_109,In_206);
nand U4601 (N_4601,In_813,In_515);
and U4602 (N_4602,In_2728,In_2582);
and U4603 (N_4603,In_1273,In_581);
nand U4604 (N_4604,In_2121,In_345);
and U4605 (N_4605,In_1571,In_1072);
xnor U4606 (N_4606,In_842,In_1469);
and U4607 (N_4607,In_237,In_772);
and U4608 (N_4608,In_825,In_296);
and U4609 (N_4609,In_921,In_2064);
and U4610 (N_4610,In_969,In_2493);
and U4611 (N_4611,In_353,In_1332);
or U4612 (N_4612,In_1095,In_918);
and U4613 (N_4613,In_555,In_684);
nor U4614 (N_4614,In_545,In_1027);
nor U4615 (N_4615,In_2144,In_1717);
or U4616 (N_4616,In_309,In_663);
or U4617 (N_4617,In_1711,In_1701);
or U4618 (N_4618,In_15,In_1894);
xnor U4619 (N_4619,In_1520,In_626);
or U4620 (N_4620,In_995,In_71);
nand U4621 (N_4621,In_546,In_2472);
nand U4622 (N_4622,In_642,In_1623);
and U4623 (N_4623,In_898,In_1493);
xnor U4624 (N_4624,In_1720,In_660);
nor U4625 (N_4625,In_2768,In_1549);
nand U4626 (N_4626,In_1340,In_1427);
nand U4627 (N_4627,In_871,In_1078);
or U4628 (N_4628,In_2859,In_795);
or U4629 (N_4629,In_2313,In_2567);
xnor U4630 (N_4630,In_887,In_2901);
or U4631 (N_4631,In_2282,In_1495);
or U4632 (N_4632,In_1296,In_295);
nor U4633 (N_4633,In_1224,In_1190);
nor U4634 (N_4634,In_548,In_114);
and U4635 (N_4635,In_2844,In_2159);
nand U4636 (N_4636,In_2017,In_1742);
or U4637 (N_4637,In_2017,In_1769);
nor U4638 (N_4638,In_1529,In_1288);
nor U4639 (N_4639,In_937,In_214);
or U4640 (N_4640,In_453,In_768);
nand U4641 (N_4641,In_1097,In_1722);
nand U4642 (N_4642,In_2398,In_2068);
and U4643 (N_4643,In_1257,In_783);
nor U4644 (N_4644,In_1483,In_1705);
or U4645 (N_4645,In_1146,In_2849);
and U4646 (N_4646,In_245,In_686);
nor U4647 (N_4647,In_982,In_1497);
or U4648 (N_4648,In_2692,In_567);
nand U4649 (N_4649,In_906,In_2924);
or U4650 (N_4650,In_887,In_715);
or U4651 (N_4651,In_2578,In_2229);
and U4652 (N_4652,In_899,In_1093);
or U4653 (N_4653,In_467,In_1081);
xor U4654 (N_4654,In_227,In_2824);
nor U4655 (N_4655,In_790,In_1586);
nand U4656 (N_4656,In_2839,In_89);
and U4657 (N_4657,In_862,In_202);
nor U4658 (N_4658,In_1312,In_1988);
nor U4659 (N_4659,In_2400,In_2283);
xor U4660 (N_4660,In_1572,In_1933);
and U4661 (N_4661,In_175,In_921);
and U4662 (N_4662,In_2549,In_2245);
xor U4663 (N_4663,In_1372,In_2126);
and U4664 (N_4664,In_2182,In_1332);
nand U4665 (N_4665,In_2709,In_2532);
and U4666 (N_4666,In_2602,In_736);
nor U4667 (N_4667,In_1087,In_556);
nor U4668 (N_4668,In_485,In_362);
nor U4669 (N_4669,In_303,In_2468);
and U4670 (N_4670,In_313,In_1007);
nand U4671 (N_4671,In_548,In_814);
nand U4672 (N_4672,In_2693,In_2374);
xnor U4673 (N_4673,In_1494,In_757);
nand U4674 (N_4674,In_1581,In_854);
and U4675 (N_4675,In_2500,In_2779);
nand U4676 (N_4676,In_1387,In_2219);
or U4677 (N_4677,In_817,In_1311);
xor U4678 (N_4678,In_396,In_860);
nand U4679 (N_4679,In_93,In_1013);
and U4680 (N_4680,In_461,In_873);
nand U4681 (N_4681,In_1302,In_1097);
xor U4682 (N_4682,In_2925,In_2372);
and U4683 (N_4683,In_1547,In_1865);
nand U4684 (N_4684,In_1703,In_1241);
or U4685 (N_4685,In_1627,In_1843);
and U4686 (N_4686,In_2104,In_1627);
nor U4687 (N_4687,In_1644,In_551);
xor U4688 (N_4688,In_770,In_2465);
nor U4689 (N_4689,In_1606,In_1912);
or U4690 (N_4690,In_523,In_1287);
or U4691 (N_4691,In_365,In_332);
or U4692 (N_4692,In_592,In_2990);
or U4693 (N_4693,In_475,In_2108);
nor U4694 (N_4694,In_2665,In_417);
nand U4695 (N_4695,In_2258,In_1060);
nand U4696 (N_4696,In_2849,In_804);
nor U4697 (N_4697,In_1786,In_1243);
nand U4698 (N_4698,In_1031,In_349);
or U4699 (N_4699,In_2483,In_2095);
xor U4700 (N_4700,In_2645,In_162);
nor U4701 (N_4701,In_1713,In_2834);
and U4702 (N_4702,In_1186,In_2498);
and U4703 (N_4703,In_1641,In_2729);
or U4704 (N_4704,In_2659,In_941);
or U4705 (N_4705,In_1272,In_367);
nand U4706 (N_4706,In_156,In_46);
or U4707 (N_4707,In_852,In_1744);
and U4708 (N_4708,In_848,In_99);
xnor U4709 (N_4709,In_969,In_95);
and U4710 (N_4710,In_414,In_2525);
or U4711 (N_4711,In_1872,In_1587);
or U4712 (N_4712,In_1606,In_1412);
nand U4713 (N_4713,In_284,In_2785);
and U4714 (N_4714,In_2660,In_411);
nor U4715 (N_4715,In_2918,In_2949);
xor U4716 (N_4716,In_69,In_954);
nand U4717 (N_4717,In_1109,In_1475);
xnor U4718 (N_4718,In_2215,In_1538);
and U4719 (N_4719,In_1121,In_1536);
nand U4720 (N_4720,In_80,In_2837);
and U4721 (N_4721,In_926,In_35);
nand U4722 (N_4722,In_334,In_458);
nor U4723 (N_4723,In_1898,In_284);
nand U4724 (N_4724,In_2571,In_777);
nand U4725 (N_4725,In_896,In_1292);
or U4726 (N_4726,In_1357,In_2638);
or U4727 (N_4727,In_1586,In_1562);
or U4728 (N_4728,In_1114,In_717);
nor U4729 (N_4729,In_2516,In_2085);
nor U4730 (N_4730,In_261,In_2615);
and U4731 (N_4731,In_2124,In_662);
and U4732 (N_4732,In_894,In_1251);
or U4733 (N_4733,In_1556,In_1972);
or U4734 (N_4734,In_1424,In_1711);
nor U4735 (N_4735,In_182,In_126);
or U4736 (N_4736,In_1307,In_1094);
and U4737 (N_4737,In_2407,In_1440);
nand U4738 (N_4738,In_491,In_454);
nor U4739 (N_4739,In_130,In_2169);
xor U4740 (N_4740,In_2679,In_326);
and U4741 (N_4741,In_1659,In_1137);
and U4742 (N_4742,In_1777,In_1796);
nor U4743 (N_4743,In_525,In_2109);
and U4744 (N_4744,In_177,In_1327);
nor U4745 (N_4745,In_923,In_757);
and U4746 (N_4746,In_517,In_2698);
nand U4747 (N_4747,In_718,In_956);
nand U4748 (N_4748,In_2535,In_1114);
nand U4749 (N_4749,In_1382,In_246);
nand U4750 (N_4750,In_1404,In_1717);
nand U4751 (N_4751,In_1013,In_1847);
or U4752 (N_4752,In_2285,In_2936);
xnor U4753 (N_4753,In_1955,In_1008);
and U4754 (N_4754,In_2701,In_989);
nor U4755 (N_4755,In_2292,In_2079);
xor U4756 (N_4756,In_103,In_143);
nor U4757 (N_4757,In_2936,In_1718);
and U4758 (N_4758,In_550,In_944);
and U4759 (N_4759,In_2791,In_1573);
and U4760 (N_4760,In_2051,In_1676);
and U4761 (N_4761,In_1356,In_840);
or U4762 (N_4762,In_1973,In_110);
or U4763 (N_4763,In_1941,In_268);
nand U4764 (N_4764,In_389,In_1256);
xnor U4765 (N_4765,In_2913,In_353);
nand U4766 (N_4766,In_1978,In_1559);
nand U4767 (N_4767,In_48,In_2682);
nor U4768 (N_4768,In_1434,In_1951);
nor U4769 (N_4769,In_757,In_526);
or U4770 (N_4770,In_520,In_409);
or U4771 (N_4771,In_1262,In_2792);
nand U4772 (N_4772,In_459,In_2868);
xor U4773 (N_4773,In_1096,In_1145);
nand U4774 (N_4774,In_956,In_874);
or U4775 (N_4775,In_478,In_1443);
xor U4776 (N_4776,In_788,In_2520);
nor U4777 (N_4777,In_2605,In_2680);
and U4778 (N_4778,In_1776,In_852);
xnor U4779 (N_4779,In_345,In_2453);
or U4780 (N_4780,In_1576,In_1159);
nor U4781 (N_4781,In_184,In_2696);
or U4782 (N_4782,In_418,In_265);
nor U4783 (N_4783,In_915,In_1987);
or U4784 (N_4784,In_2276,In_1807);
and U4785 (N_4785,In_2066,In_1313);
nand U4786 (N_4786,In_630,In_2093);
or U4787 (N_4787,In_1436,In_1069);
and U4788 (N_4788,In_2043,In_2815);
nand U4789 (N_4789,In_1968,In_2446);
or U4790 (N_4790,In_2671,In_741);
nand U4791 (N_4791,In_359,In_2378);
nand U4792 (N_4792,In_685,In_973);
and U4793 (N_4793,In_396,In_2011);
xor U4794 (N_4794,In_273,In_817);
or U4795 (N_4795,In_1844,In_747);
nor U4796 (N_4796,In_2321,In_2270);
nand U4797 (N_4797,In_2931,In_1867);
or U4798 (N_4798,In_466,In_2136);
nor U4799 (N_4799,In_1507,In_765);
or U4800 (N_4800,In_1239,In_1167);
or U4801 (N_4801,In_1702,In_151);
or U4802 (N_4802,In_1009,In_78);
or U4803 (N_4803,In_2180,In_1057);
or U4804 (N_4804,In_2617,In_2131);
xnor U4805 (N_4805,In_1301,In_2998);
nor U4806 (N_4806,In_1536,In_1560);
or U4807 (N_4807,In_1323,In_2688);
and U4808 (N_4808,In_1404,In_1828);
nand U4809 (N_4809,In_2149,In_1289);
or U4810 (N_4810,In_2765,In_2404);
nand U4811 (N_4811,In_305,In_103);
or U4812 (N_4812,In_1023,In_2135);
and U4813 (N_4813,In_143,In_2981);
nor U4814 (N_4814,In_2342,In_965);
nand U4815 (N_4815,In_1668,In_746);
nor U4816 (N_4816,In_2717,In_1933);
nor U4817 (N_4817,In_2764,In_788);
or U4818 (N_4818,In_2151,In_1808);
xor U4819 (N_4819,In_2677,In_1897);
and U4820 (N_4820,In_2026,In_2182);
and U4821 (N_4821,In_1611,In_304);
nand U4822 (N_4822,In_259,In_862);
nor U4823 (N_4823,In_1756,In_733);
and U4824 (N_4824,In_2130,In_23);
or U4825 (N_4825,In_328,In_1933);
nor U4826 (N_4826,In_1083,In_2542);
nor U4827 (N_4827,In_2377,In_1134);
or U4828 (N_4828,In_2213,In_2232);
nor U4829 (N_4829,In_564,In_1675);
nand U4830 (N_4830,In_1487,In_1129);
nand U4831 (N_4831,In_745,In_1824);
nor U4832 (N_4832,In_2150,In_204);
nand U4833 (N_4833,In_1957,In_1812);
or U4834 (N_4834,In_481,In_1740);
and U4835 (N_4835,In_1402,In_2);
and U4836 (N_4836,In_92,In_2629);
nand U4837 (N_4837,In_2292,In_2988);
or U4838 (N_4838,In_259,In_1613);
or U4839 (N_4839,In_2768,In_1094);
xor U4840 (N_4840,In_1692,In_118);
or U4841 (N_4841,In_2320,In_532);
and U4842 (N_4842,In_2662,In_2508);
nand U4843 (N_4843,In_2697,In_2480);
or U4844 (N_4844,In_2656,In_1185);
nor U4845 (N_4845,In_1541,In_1350);
nand U4846 (N_4846,In_922,In_489);
nor U4847 (N_4847,In_2621,In_1600);
nand U4848 (N_4848,In_1596,In_2706);
nand U4849 (N_4849,In_2866,In_1586);
and U4850 (N_4850,In_1749,In_2799);
nor U4851 (N_4851,In_793,In_1626);
nor U4852 (N_4852,In_1091,In_2704);
nor U4853 (N_4853,In_1559,In_1211);
nor U4854 (N_4854,In_2175,In_1527);
and U4855 (N_4855,In_20,In_1987);
and U4856 (N_4856,In_2927,In_2988);
and U4857 (N_4857,In_2937,In_1141);
nor U4858 (N_4858,In_2779,In_554);
and U4859 (N_4859,In_1492,In_2550);
and U4860 (N_4860,In_282,In_1584);
nand U4861 (N_4861,In_1787,In_1328);
nand U4862 (N_4862,In_2198,In_152);
nor U4863 (N_4863,In_2577,In_946);
or U4864 (N_4864,In_2429,In_976);
nand U4865 (N_4865,In_1705,In_451);
or U4866 (N_4866,In_889,In_1601);
nor U4867 (N_4867,In_767,In_2345);
and U4868 (N_4868,In_894,In_2655);
nand U4869 (N_4869,In_2608,In_161);
or U4870 (N_4870,In_1514,In_1100);
nand U4871 (N_4871,In_2659,In_2864);
or U4872 (N_4872,In_2324,In_1431);
nand U4873 (N_4873,In_1994,In_420);
or U4874 (N_4874,In_270,In_1087);
nor U4875 (N_4875,In_2634,In_2306);
and U4876 (N_4876,In_199,In_586);
and U4877 (N_4877,In_207,In_202);
nand U4878 (N_4878,In_182,In_448);
and U4879 (N_4879,In_2057,In_1070);
nand U4880 (N_4880,In_1432,In_1908);
xnor U4881 (N_4881,In_1334,In_1868);
xor U4882 (N_4882,In_1361,In_2466);
nand U4883 (N_4883,In_1743,In_238);
nand U4884 (N_4884,In_2741,In_1895);
xnor U4885 (N_4885,In_1605,In_739);
or U4886 (N_4886,In_1858,In_1360);
nand U4887 (N_4887,In_1592,In_1457);
or U4888 (N_4888,In_1975,In_2332);
or U4889 (N_4889,In_2431,In_1319);
or U4890 (N_4890,In_1152,In_1424);
xnor U4891 (N_4891,In_1641,In_102);
and U4892 (N_4892,In_113,In_1821);
and U4893 (N_4893,In_149,In_1317);
nand U4894 (N_4894,In_1515,In_1136);
or U4895 (N_4895,In_2612,In_977);
and U4896 (N_4896,In_1129,In_697);
and U4897 (N_4897,In_697,In_2988);
and U4898 (N_4898,In_540,In_1001);
xnor U4899 (N_4899,In_1215,In_90);
or U4900 (N_4900,In_2002,In_2821);
or U4901 (N_4901,In_257,In_1630);
and U4902 (N_4902,In_2707,In_1225);
nand U4903 (N_4903,In_981,In_2186);
and U4904 (N_4904,In_1270,In_357);
nand U4905 (N_4905,In_321,In_1597);
and U4906 (N_4906,In_2775,In_53);
or U4907 (N_4907,In_1424,In_1213);
xnor U4908 (N_4908,In_2041,In_932);
nor U4909 (N_4909,In_2394,In_2114);
nand U4910 (N_4910,In_2567,In_1274);
nand U4911 (N_4911,In_2981,In_1899);
or U4912 (N_4912,In_433,In_2225);
or U4913 (N_4913,In_2463,In_68);
and U4914 (N_4914,In_63,In_2233);
and U4915 (N_4915,In_340,In_1610);
or U4916 (N_4916,In_2371,In_2427);
nor U4917 (N_4917,In_2936,In_2870);
nand U4918 (N_4918,In_2284,In_2836);
and U4919 (N_4919,In_248,In_2895);
or U4920 (N_4920,In_784,In_2288);
nand U4921 (N_4921,In_421,In_1001);
nor U4922 (N_4922,In_2890,In_1908);
nor U4923 (N_4923,In_2798,In_2665);
and U4924 (N_4924,In_2606,In_875);
nor U4925 (N_4925,In_1178,In_378);
nor U4926 (N_4926,In_506,In_2018);
nand U4927 (N_4927,In_2098,In_2298);
nor U4928 (N_4928,In_2604,In_1219);
xor U4929 (N_4929,In_2290,In_1724);
nor U4930 (N_4930,In_117,In_2333);
or U4931 (N_4931,In_225,In_1579);
nor U4932 (N_4932,In_180,In_1206);
xnor U4933 (N_4933,In_1917,In_294);
nor U4934 (N_4934,In_1326,In_804);
nand U4935 (N_4935,In_1129,In_649);
or U4936 (N_4936,In_477,In_2848);
nand U4937 (N_4937,In_1901,In_273);
and U4938 (N_4938,In_1345,In_2349);
or U4939 (N_4939,In_1233,In_1171);
xor U4940 (N_4940,In_1814,In_1692);
xor U4941 (N_4941,In_2974,In_2758);
nor U4942 (N_4942,In_1314,In_1320);
nand U4943 (N_4943,In_299,In_405);
nor U4944 (N_4944,In_1182,In_991);
and U4945 (N_4945,In_1097,In_2429);
nand U4946 (N_4946,In_1087,In_2095);
nor U4947 (N_4947,In_124,In_1752);
and U4948 (N_4948,In_1325,In_1152);
nand U4949 (N_4949,In_907,In_456);
xnor U4950 (N_4950,In_169,In_176);
and U4951 (N_4951,In_2898,In_520);
or U4952 (N_4952,In_1061,In_162);
nand U4953 (N_4953,In_1623,In_1385);
or U4954 (N_4954,In_1624,In_1572);
nand U4955 (N_4955,In_1771,In_474);
nand U4956 (N_4956,In_1407,In_2960);
nor U4957 (N_4957,In_2365,In_1960);
nor U4958 (N_4958,In_51,In_2);
nor U4959 (N_4959,In_33,In_2613);
nand U4960 (N_4960,In_275,In_163);
or U4961 (N_4961,In_1899,In_2535);
and U4962 (N_4962,In_1124,In_1111);
and U4963 (N_4963,In_697,In_1788);
and U4964 (N_4964,In_2400,In_1505);
and U4965 (N_4965,In_2727,In_2112);
and U4966 (N_4966,In_2066,In_234);
xnor U4967 (N_4967,In_1752,In_1169);
and U4968 (N_4968,In_1280,In_1639);
or U4969 (N_4969,In_65,In_489);
or U4970 (N_4970,In_2009,In_2550);
nor U4971 (N_4971,In_349,In_2508);
nor U4972 (N_4972,In_928,In_342);
and U4973 (N_4973,In_2035,In_2802);
nor U4974 (N_4974,In_2850,In_612);
or U4975 (N_4975,In_9,In_1199);
nor U4976 (N_4976,In_2357,In_1315);
nor U4977 (N_4977,In_2620,In_317);
nand U4978 (N_4978,In_2588,In_1615);
or U4979 (N_4979,In_593,In_2532);
and U4980 (N_4980,In_1347,In_559);
and U4981 (N_4981,In_1451,In_2982);
nor U4982 (N_4982,In_1749,In_87);
nor U4983 (N_4983,In_2272,In_1613);
nand U4984 (N_4984,In_1595,In_1123);
and U4985 (N_4985,In_2166,In_1184);
or U4986 (N_4986,In_2776,In_248);
and U4987 (N_4987,In_838,In_943);
or U4988 (N_4988,In_2073,In_1145);
nand U4989 (N_4989,In_2207,In_1565);
or U4990 (N_4990,In_854,In_420);
or U4991 (N_4991,In_2141,In_2269);
nor U4992 (N_4992,In_189,In_1584);
or U4993 (N_4993,In_1614,In_2792);
and U4994 (N_4994,In_10,In_1596);
nand U4995 (N_4995,In_221,In_577);
xor U4996 (N_4996,In_2736,In_834);
and U4997 (N_4997,In_766,In_1779);
nand U4998 (N_4998,In_340,In_299);
nor U4999 (N_4999,In_934,In_2525);
nand U5000 (N_5000,N_2033,N_968);
xnor U5001 (N_5001,N_3213,N_394);
nor U5002 (N_5002,N_2859,N_3816);
or U5003 (N_5003,N_3784,N_4408);
xor U5004 (N_5004,N_3436,N_1731);
nand U5005 (N_5005,N_2023,N_361);
nor U5006 (N_5006,N_3651,N_1497);
or U5007 (N_5007,N_3366,N_1231);
nand U5008 (N_5008,N_2899,N_3129);
xor U5009 (N_5009,N_3778,N_1927);
nand U5010 (N_5010,N_2190,N_4047);
nand U5011 (N_5011,N_3602,N_325);
or U5012 (N_5012,N_2642,N_3068);
and U5013 (N_5013,N_3496,N_4777);
or U5014 (N_5014,N_4182,N_2312);
nor U5015 (N_5015,N_2466,N_4950);
nor U5016 (N_5016,N_1397,N_935);
and U5017 (N_5017,N_3363,N_2932);
and U5018 (N_5018,N_1585,N_644);
and U5019 (N_5019,N_4011,N_2933);
nand U5020 (N_5020,N_2557,N_1429);
or U5021 (N_5021,N_3373,N_2350);
and U5022 (N_5022,N_4079,N_2357);
or U5023 (N_5023,N_91,N_1437);
and U5024 (N_5024,N_1123,N_667);
or U5025 (N_5025,N_4945,N_2527);
nor U5026 (N_5026,N_2979,N_943);
nand U5027 (N_5027,N_2674,N_4872);
or U5028 (N_5028,N_987,N_2739);
nand U5029 (N_5029,N_4202,N_1803);
and U5030 (N_5030,N_4068,N_972);
and U5031 (N_5031,N_1897,N_932);
nand U5032 (N_5032,N_2040,N_1906);
nor U5033 (N_5033,N_1118,N_1716);
nor U5034 (N_5034,N_1145,N_3697);
nor U5035 (N_5035,N_3769,N_3395);
nor U5036 (N_5036,N_3327,N_4978);
and U5037 (N_5037,N_2305,N_3276);
and U5038 (N_5038,N_1626,N_1923);
or U5039 (N_5039,N_3793,N_4262);
nor U5040 (N_5040,N_822,N_1156);
or U5041 (N_5041,N_3702,N_4063);
and U5042 (N_5042,N_475,N_1637);
xor U5043 (N_5043,N_1841,N_3114);
or U5044 (N_5044,N_2605,N_365);
or U5045 (N_5045,N_3192,N_211);
nor U5046 (N_5046,N_537,N_3779);
xor U5047 (N_5047,N_3111,N_4897);
and U5048 (N_5048,N_4748,N_3918);
nor U5049 (N_5049,N_1606,N_800);
and U5050 (N_5050,N_3689,N_582);
nand U5051 (N_5051,N_4100,N_185);
and U5052 (N_5052,N_3903,N_4775);
nand U5053 (N_5053,N_4380,N_2953);
xnor U5054 (N_5054,N_4649,N_1845);
nand U5055 (N_5055,N_508,N_3818);
xnor U5056 (N_5056,N_4814,N_230);
or U5057 (N_5057,N_2798,N_696);
nand U5058 (N_5058,N_3226,N_848);
nor U5059 (N_5059,N_2637,N_2839);
or U5060 (N_5060,N_2247,N_4264);
nor U5061 (N_5061,N_4903,N_2036);
and U5062 (N_5062,N_3522,N_1763);
nand U5063 (N_5063,N_445,N_846);
or U5064 (N_5064,N_3355,N_4732);
or U5065 (N_5065,N_3569,N_1571);
nor U5066 (N_5066,N_3584,N_853);
nor U5067 (N_5067,N_3583,N_2081);
or U5068 (N_5068,N_3016,N_1873);
xor U5069 (N_5069,N_4270,N_3259);
nor U5070 (N_5070,N_766,N_1);
or U5071 (N_5071,N_633,N_3251);
or U5072 (N_5072,N_1456,N_1146);
and U5073 (N_5073,N_864,N_425);
or U5074 (N_5074,N_1255,N_1227);
nand U5075 (N_5075,N_1382,N_3150);
or U5076 (N_5076,N_2266,N_3973);
or U5077 (N_5077,N_99,N_3336);
and U5078 (N_5078,N_958,N_4967);
and U5079 (N_5079,N_659,N_3834);
nor U5080 (N_5080,N_3293,N_4888);
and U5081 (N_5081,N_676,N_3037);
nor U5082 (N_5082,N_2311,N_4679);
or U5083 (N_5083,N_1620,N_4933);
or U5084 (N_5084,N_1291,N_4420);
and U5085 (N_5085,N_2892,N_3298);
or U5086 (N_5086,N_3369,N_262);
nand U5087 (N_5087,N_44,N_1813);
nand U5088 (N_5088,N_3578,N_1475);
nor U5089 (N_5089,N_336,N_1423);
nand U5090 (N_5090,N_1868,N_926);
xnor U5091 (N_5091,N_2157,N_4625);
nor U5092 (N_5092,N_1838,N_2070);
nand U5093 (N_5093,N_287,N_4163);
nor U5094 (N_5094,N_2594,N_3688);
and U5095 (N_5095,N_173,N_4103);
xnor U5096 (N_5096,N_1165,N_248);
and U5097 (N_5097,N_1371,N_123);
nor U5098 (N_5098,N_3085,N_4158);
and U5099 (N_5099,N_3675,N_4746);
and U5100 (N_5100,N_2884,N_3864);
or U5101 (N_5101,N_493,N_594);
and U5102 (N_5102,N_803,N_1024);
or U5103 (N_5103,N_3380,N_4818);
or U5104 (N_5104,N_993,N_4980);
nand U5105 (N_5105,N_3310,N_3938);
nor U5106 (N_5106,N_3167,N_4648);
nor U5107 (N_5107,N_4533,N_218);
or U5108 (N_5108,N_1132,N_1455);
and U5109 (N_5109,N_2998,N_1934);
nor U5110 (N_5110,N_4144,N_2046);
nand U5111 (N_5111,N_2608,N_3690);
and U5112 (N_5112,N_4567,N_4469);
nand U5113 (N_5113,N_2283,N_2349);
nand U5114 (N_5114,N_4651,N_4132);
and U5115 (N_5115,N_1966,N_3617);
nand U5116 (N_5116,N_1912,N_1018);
xnor U5117 (N_5117,N_2090,N_3108);
nor U5118 (N_5118,N_3283,N_4785);
nand U5119 (N_5119,N_1721,N_1680);
and U5120 (N_5120,N_4200,N_3655);
nor U5121 (N_5121,N_3539,N_3370);
nor U5122 (N_5122,N_3252,N_1312);
and U5123 (N_5123,N_4225,N_3997);
nor U5124 (N_5124,N_4689,N_3764);
nor U5125 (N_5125,N_4383,N_2614);
nor U5126 (N_5126,N_1183,N_4143);
or U5127 (N_5127,N_1301,N_4924);
and U5128 (N_5128,N_4621,N_1764);
and U5129 (N_5129,N_884,N_4823);
nor U5130 (N_5130,N_4570,N_3971);
nor U5131 (N_5131,N_2927,N_1267);
xnor U5132 (N_5132,N_2352,N_1494);
or U5133 (N_5133,N_2624,N_2420);
xor U5134 (N_5134,N_1222,N_1150);
or U5135 (N_5135,N_4882,N_2497);
or U5136 (N_5136,N_754,N_3763);
and U5137 (N_5137,N_776,N_3233);
or U5138 (N_5138,N_4471,N_78);
and U5139 (N_5139,N_811,N_3475);
and U5140 (N_5140,N_1970,N_3679);
xor U5141 (N_5141,N_1619,N_1493);
xor U5142 (N_5142,N_16,N_3450);
nand U5143 (N_5143,N_42,N_1916);
nor U5144 (N_5144,N_3739,N_912);
or U5145 (N_5145,N_2567,N_4551);
xor U5146 (N_5146,N_3603,N_1653);
or U5147 (N_5147,N_3711,N_4083);
xnor U5148 (N_5148,N_1939,N_4759);
and U5149 (N_5149,N_1263,N_3976);
nand U5150 (N_5150,N_2801,N_774);
nand U5151 (N_5151,N_921,N_453);
nand U5152 (N_5152,N_1561,N_2316);
nand U5153 (N_5153,N_670,N_4682);
nor U5154 (N_5154,N_1209,N_4582);
nor U5155 (N_5155,N_4437,N_975);
nand U5156 (N_5156,N_3714,N_1305);
nand U5157 (N_5157,N_37,N_3017);
nand U5158 (N_5158,N_818,N_4261);
nand U5159 (N_5159,N_2340,N_4465);
nand U5160 (N_5160,N_4634,N_1818);
and U5161 (N_5161,N_748,N_1586);
or U5162 (N_5162,N_4805,N_4877);
xor U5163 (N_5163,N_2203,N_282);
nand U5164 (N_5164,N_2843,N_3926);
or U5165 (N_5165,N_1082,N_4711);
nand U5166 (N_5166,N_4628,N_519);
xor U5167 (N_5167,N_4138,N_4377);
xnor U5168 (N_5168,N_624,N_2758);
and U5169 (N_5169,N_3383,N_4535);
nand U5170 (N_5170,N_2573,N_4052);
and U5171 (N_5171,N_4658,N_1746);
nor U5172 (N_5172,N_4911,N_1609);
nor U5173 (N_5173,N_3038,N_4055);
nor U5174 (N_5174,N_1472,N_4678);
nand U5175 (N_5175,N_4384,N_291);
or U5176 (N_5176,N_59,N_4479);
xor U5177 (N_5177,N_1468,N_2235);
or U5178 (N_5178,N_2286,N_3178);
and U5179 (N_5179,N_63,N_1749);
or U5180 (N_5180,N_1590,N_2812);
or U5181 (N_5181,N_3703,N_2776);
and U5182 (N_5182,N_551,N_2525);
or U5183 (N_5183,N_3908,N_552);
and U5184 (N_5184,N_2067,N_1499);
or U5185 (N_5185,N_3507,N_573);
and U5186 (N_5186,N_2610,N_572);
nor U5187 (N_5187,N_665,N_1323);
nor U5188 (N_5188,N_1216,N_3521);
nand U5189 (N_5189,N_2285,N_4970);
and U5190 (N_5190,N_2313,N_2178);
and U5191 (N_5191,N_3883,N_2727);
nand U5192 (N_5192,N_1117,N_1965);
nor U5193 (N_5193,N_3007,N_3154);
nand U5194 (N_5194,N_1668,N_75);
nand U5195 (N_5195,N_3061,N_167);
nand U5196 (N_5196,N_3439,N_4485);
nor U5197 (N_5197,N_4425,N_3237);
nor U5198 (N_5198,N_4695,N_4547);
xnor U5199 (N_5199,N_4604,N_1706);
nand U5200 (N_5200,N_2034,N_4273);
nand U5201 (N_5201,N_4293,N_1135);
or U5202 (N_5202,N_2869,N_4107);
or U5203 (N_5203,N_4253,N_2849);
nand U5204 (N_5204,N_3901,N_227);
nor U5205 (N_5205,N_3429,N_47);
nand U5206 (N_5206,N_4507,N_2086);
or U5207 (N_5207,N_386,N_619);
nand U5208 (N_5208,N_370,N_1019);
and U5209 (N_5209,N_1023,N_3664);
nand U5210 (N_5210,N_208,N_547);
xnor U5211 (N_5211,N_2214,N_3282);
nand U5212 (N_5212,N_2707,N_3188);
nand U5213 (N_5213,N_1346,N_1751);
and U5214 (N_5214,N_1377,N_3073);
or U5215 (N_5215,N_1967,N_2022);
or U5216 (N_5216,N_4358,N_2621);
and U5217 (N_5217,N_1277,N_2684);
nand U5218 (N_5218,N_829,N_1618);
nor U5219 (N_5219,N_201,N_2465);
and U5220 (N_5220,N_1390,N_3033);
nand U5221 (N_5221,N_2765,N_1553);
nand U5222 (N_5222,N_3771,N_4162);
and U5223 (N_5223,N_4925,N_1199);
nor U5224 (N_5224,N_4976,N_423);
or U5225 (N_5225,N_511,N_1781);
nor U5226 (N_5226,N_3914,N_2031);
nand U5227 (N_5227,N_1385,N_653);
nor U5228 (N_5228,N_3090,N_436);
nand U5229 (N_5229,N_4954,N_807);
and U5230 (N_5230,N_1115,N_2631);
nor U5231 (N_5231,N_3579,N_1104);
or U5232 (N_5232,N_4378,N_3054);
nor U5233 (N_5233,N_334,N_990);
or U5234 (N_5234,N_2717,N_2576);
or U5235 (N_5235,N_3257,N_1252);
or U5236 (N_5236,N_1896,N_528);
nor U5237 (N_5237,N_1401,N_3483);
or U5238 (N_5238,N_3790,N_723);
xnor U5239 (N_5239,N_1948,N_2781);
nand U5240 (N_5240,N_1414,N_859);
nand U5241 (N_5241,N_4815,N_2623);
xor U5242 (N_5242,N_4643,N_1032);
nor U5243 (N_5243,N_3216,N_3208);
nand U5244 (N_5244,N_4607,N_204);
nand U5245 (N_5245,N_4444,N_3828);
and U5246 (N_5246,N_2719,N_1476);
and U5247 (N_5247,N_1839,N_4140);
or U5248 (N_5248,N_3833,N_84);
nand U5249 (N_5249,N_3631,N_137);
xnor U5250 (N_5250,N_2289,N_843);
or U5251 (N_5251,N_3665,N_1396);
nand U5252 (N_5252,N_2653,N_2800);
xor U5253 (N_5253,N_2873,N_1114);
nor U5254 (N_5254,N_728,N_410);
nand U5255 (N_5255,N_3887,N_4630);
and U5256 (N_5256,N_2991,N_247);
or U5257 (N_5257,N_3094,N_3406);
and U5258 (N_5258,N_2968,N_589);
or U5259 (N_5259,N_816,N_601);
and U5260 (N_5260,N_925,N_1030);
xor U5261 (N_5261,N_4065,N_4269);
or U5262 (N_5262,N_4589,N_4185);
and U5263 (N_5263,N_3528,N_839);
or U5264 (N_5264,N_1353,N_160);
or U5265 (N_5265,N_4537,N_1313);
nor U5266 (N_5266,N_320,N_3983);
nand U5267 (N_5267,N_3142,N_4310);
xnor U5268 (N_5268,N_3855,N_1715);
and U5269 (N_5269,N_109,N_153);
nor U5270 (N_5270,N_641,N_4769);
or U5271 (N_5271,N_3845,N_179);
and U5272 (N_5272,N_1003,N_3131);
nand U5273 (N_5273,N_1614,N_409);
nor U5274 (N_5274,N_2087,N_1142);
and U5275 (N_5275,N_2137,N_513);
or U5276 (N_5276,N_3411,N_304);
nor U5277 (N_5277,N_885,N_3510);
nor U5278 (N_5278,N_3506,N_408);
or U5279 (N_5279,N_2520,N_1355);
and U5280 (N_5280,N_1737,N_3840);
nor U5281 (N_5281,N_2750,N_4306);
xor U5282 (N_5282,N_4744,N_1098);
nand U5283 (N_5283,N_3235,N_2460);
xnor U5284 (N_5284,N_317,N_3091);
or U5285 (N_5285,N_4865,N_4700);
nand U5286 (N_5286,N_3354,N_4540);
nor U5287 (N_5287,N_1727,N_4553);
nor U5288 (N_5288,N_4228,N_2192);
and U5289 (N_5289,N_4265,N_2029);
or U5290 (N_5290,N_1513,N_627);
or U5291 (N_5291,N_597,N_4749);
or U5292 (N_5292,N_4025,N_801);
nand U5293 (N_5293,N_1000,N_95);
nor U5294 (N_5294,N_1331,N_554);
or U5295 (N_5295,N_3721,N_4821);
nor U5296 (N_5296,N_3117,N_2381);
or U5297 (N_5297,N_3805,N_707);
or U5298 (N_5298,N_3403,N_1230);
nand U5299 (N_5299,N_4274,N_3180);
nor U5300 (N_5300,N_4160,N_2200);
and U5301 (N_5301,N_1449,N_3468);
nor U5302 (N_5302,N_4327,N_2508);
or U5303 (N_5303,N_634,N_1459);
nor U5304 (N_5304,N_2229,N_4910);
nor U5305 (N_5305,N_1771,N_4247);
and U5306 (N_5306,N_3338,N_3624);
or U5307 (N_5307,N_420,N_2320);
nand U5308 (N_5308,N_3044,N_79);
nor U5309 (N_5309,N_4472,N_13);
or U5310 (N_5310,N_1411,N_1596);
nand U5311 (N_5311,N_3254,N_4586);
nor U5312 (N_5312,N_253,N_3944);
nor U5313 (N_5313,N_2282,N_3802);
xnor U5314 (N_5314,N_2771,N_4217);
nand U5315 (N_5315,N_3952,N_3303);
nor U5316 (N_5316,N_622,N_404);
nor U5317 (N_5317,N_2387,N_2894);
nor U5318 (N_5318,N_4867,N_649);
and U5319 (N_5319,N_1028,N_4027);
nor U5320 (N_5320,N_4892,N_3486);
nand U5321 (N_5321,N_3656,N_2291);
or U5322 (N_5322,N_4928,N_4347);
or U5323 (N_5323,N_1792,N_1406);
or U5324 (N_5324,N_2575,N_3968);
or U5325 (N_5325,N_1926,N_1239);
nand U5326 (N_5326,N_3018,N_3286);
xor U5327 (N_5327,N_2685,N_2026);
or U5328 (N_5328,N_3045,N_2754);
nand U5329 (N_5329,N_4098,N_719);
nor U5330 (N_5330,N_2397,N_559);
and U5331 (N_5331,N_1833,N_12);
nand U5332 (N_5332,N_2210,N_4677);
or U5333 (N_5333,N_359,N_4135);
or U5334 (N_5334,N_372,N_1014);
nor U5335 (N_5335,N_4277,N_3994);
and U5336 (N_5336,N_446,N_1631);
nand U5337 (N_5337,N_283,N_2622);
nor U5338 (N_5338,N_4955,N_2233);
or U5339 (N_5339,N_3342,N_2515);
nor U5340 (N_5340,N_11,N_1478);
or U5341 (N_5341,N_2396,N_4803);
nor U5342 (N_5342,N_1648,N_3939);
or U5343 (N_5343,N_2524,N_4434);
or U5344 (N_5344,N_2261,N_3497);
and U5345 (N_5345,N_4451,N_646);
and U5346 (N_5346,N_4354,N_712);
and U5347 (N_5347,N_4716,N_371);
or U5348 (N_5348,N_996,N_2384);
nand U5349 (N_5349,N_3667,N_1365);
or U5350 (N_5350,N_233,N_3893);
xor U5351 (N_5351,N_440,N_4004);
and U5352 (N_5352,N_1726,N_1791);
and U5353 (N_5353,N_2786,N_1369);
or U5354 (N_5354,N_3807,N_507);
or U5355 (N_5355,N_3272,N_1127);
nor U5356 (N_5356,N_4934,N_3869);
nor U5357 (N_5357,N_2636,N_2926);
or U5358 (N_5358,N_1198,N_1848);
and U5359 (N_5359,N_2250,N_550);
nor U5360 (N_5360,N_3135,N_900);
nand U5361 (N_5361,N_998,N_772);
nor U5362 (N_5362,N_2655,N_1482);
or U5363 (N_5363,N_1684,N_690);
nor U5364 (N_5364,N_396,N_1774);
or U5365 (N_5365,N_3055,N_963);
or U5366 (N_5366,N_3894,N_3511);
xnor U5367 (N_5367,N_4614,N_4433);
xor U5368 (N_5368,N_1678,N_3242);
nor U5369 (N_5369,N_4216,N_32);
and U5370 (N_5370,N_2904,N_868);
and U5371 (N_5371,N_4526,N_2102);
nor U5372 (N_5372,N_3284,N_200);
nand U5373 (N_5373,N_309,N_1563);
nor U5374 (N_5374,N_1254,N_3132);
or U5375 (N_5375,N_3144,N_3653);
and U5376 (N_5376,N_4020,N_4263);
and U5377 (N_5377,N_21,N_2517);
nand U5378 (N_5378,N_4164,N_2072);
xnor U5379 (N_5379,N_180,N_4176);
nor U5380 (N_5380,N_3074,N_2428);
nand U5381 (N_5381,N_3531,N_4379);
and U5382 (N_5382,N_347,N_2035);
nand U5383 (N_5383,N_294,N_4542);
nand U5384 (N_5384,N_2394,N_2767);
or U5385 (N_5385,N_2133,N_845);
or U5386 (N_5386,N_1775,N_4345);
and U5387 (N_5387,N_1006,N_3947);
nor U5388 (N_5388,N_451,N_1416);
nor U5389 (N_5389,N_2480,N_3059);
or U5390 (N_5390,N_2867,N_1153);
and U5391 (N_5391,N_4985,N_2516);
nor U5392 (N_5392,N_3707,N_3123);
or U5393 (N_5393,N_4671,N_380);
nor U5394 (N_5394,N_1919,N_3351);
or U5395 (N_5395,N_2723,N_3409);
or U5396 (N_5396,N_1575,N_3534);
nor U5397 (N_5397,N_3937,N_4667);
nand U5398 (N_5398,N_1220,N_2984);
nand U5399 (N_5399,N_4598,N_1201);
or U5400 (N_5400,N_1880,N_362);
nor U5401 (N_5401,N_3480,N_4305);
nor U5402 (N_5402,N_2531,N_1802);
xor U5403 (N_5403,N_2977,N_389);
nand U5404 (N_5404,N_4364,N_3970);
nor U5405 (N_5405,N_473,N_852);
nand U5406 (N_5406,N_4308,N_4923);
nor U5407 (N_5407,N_1736,N_3072);
nand U5408 (N_5408,N_3517,N_3043);
nor U5409 (N_5409,N_3568,N_2364);
and U5410 (N_5410,N_102,N_1889);
xnor U5411 (N_5411,N_490,N_2549);
nor U5412 (N_5412,N_50,N_2736);
nand U5413 (N_5413,N_1084,N_2947);
and U5414 (N_5414,N_1533,N_1203);
and U5415 (N_5415,N_2073,N_2014);
nand U5416 (N_5416,N_1712,N_1167);
nor U5417 (N_5417,N_2789,N_3164);
nand U5418 (N_5418,N_2016,N_1643);
and U5419 (N_5419,N_1959,N_4617);
nor U5420 (N_5420,N_2220,N_4307);
and U5421 (N_5421,N_4854,N_4901);
xor U5422 (N_5422,N_4483,N_1647);
xnor U5423 (N_5423,N_4812,N_2589);
nor U5424 (N_5424,N_2960,N_1767);
and U5425 (N_5425,N_3102,N_31);
and U5426 (N_5426,N_447,N_2355);
nor U5427 (N_5427,N_730,N_3999);
or U5428 (N_5428,N_3389,N_3122);
or U5429 (N_5429,N_4067,N_3339);
nand U5430 (N_5430,N_4381,N_971);
nand U5431 (N_5431,N_2345,N_2940);
and U5432 (N_5432,N_1722,N_1567);
xor U5433 (N_5433,N_1995,N_2779);
or U5434 (N_5434,N_1915,N_1122);
nand U5435 (N_5435,N_3485,N_112);
nand U5436 (N_5436,N_849,N_40);
nor U5437 (N_5437,N_4258,N_566);
nand U5438 (N_5438,N_4106,N_2080);
or U5439 (N_5439,N_4195,N_955);
nand U5440 (N_5440,N_4544,N_3230);
and U5441 (N_5441,N_1956,N_2710);
and U5442 (N_5442,N_1753,N_545);
nor U5443 (N_5443,N_1809,N_3481);
or U5444 (N_5444,N_1213,N_1107);
nor U5445 (N_5445,N_3444,N_243);
and U5446 (N_5446,N_4757,N_4870);
nor U5447 (N_5447,N_3321,N_534);
nand U5448 (N_5448,N_1730,N_4424);
and U5449 (N_5449,N_3227,N_4858);
xor U5450 (N_5450,N_4478,N_738);
nand U5451 (N_5451,N_4342,N_1496);
and U5452 (N_5452,N_4272,N_2239);
nand U5453 (N_5453,N_3787,N_3799);
or U5454 (N_5454,N_2060,N_2265);
xor U5455 (N_5455,N_139,N_4828);
nand U5456 (N_5456,N_4992,N_888);
nor U5457 (N_5457,N_4656,N_82);
nand U5458 (N_5458,N_3052,N_4611);
xor U5459 (N_5459,N_1744,N_2756);
or U5460 (N_5460,N_382,N_3716);
and U5461 (N_5461,N_1253,N_349);
or U5462 (N_5462,N_2415,N_1450);
nor U5463 (N_5463,N_4319,N_2696);
or U5464 (N_5464,N_2954,N_3039);
nor U5465 (N_5465,N_2537,N_1679);
and U5466 (N_5466,N_3533,N_3095);
nand U5467 (N_5467,N_1874,N_4240);
xnor U5468 (N_5468,N_563,N_2809);
nand U5469 (N_5469,N_2906,N_4007);
nand U5470 (N_5470,N_4766,N_3979);
xnor U5471 (N_5471,N_2053,N_2383);
nand U5472 (N_5472,N_1384,N_1392);
nor U5473 (N_5473,N_2783,N_191);
or U5474 (N_5474,N_1428,N_1527);
nand U5475 (N_5475,N_3385,N_4987);
or U5476 (N_5476,N_1034,N_3446);
nor U5477 (N_5477,N_556,N_4654);
nor U5478 (N_5478,N_4413,N_1560);
or U5479 (N_5479,N_1974,N_1177);
nor U5480 (N_5480,N_4491,N_3184);
and U5481 (N_5481,N_3698,N_3873);
or U5482 (N_5482,N_1458,N_1228);
nor U5483 (N_5483,N_4593,N_890);
and U5484 (N_5484,N_695,N_2901);
or U5485 (N_5485,N_3299,N_2187);
nand U5486 (N_5486,N_2482,N_4005);
nor U5487 (N_5487,N_3660,N_4154);
and U5488 (N_5488,N_1599,N_4565);
nand U5489 (N_5489,N_4122,N_1992);
nand U5490 (N_5490,N_3929,N_441);
nand U5491 (N_5491,N_722,N_1403);
or U5492 (N_5492,N_2025,N_4276);
or U5493 (N_5493,N_4811,N_163);
nand U5494 (N_5494,N_2663,N_3889);
xor U5495 (N_5495,N_4119,N_2772);
nor U5496 (N_5496,N_3582,N_1010);
or U5497 (N_5497,N_443,N_2408);
or U5498 (N_5498,N_737,N_412);
and U5499 (N_5499,N_1794,N_3713);
and U5500 (N_5500,N_2540,N_1502);
or U5501 (N_5501,N_1436,N_2139);
xor U5502 (N_5502,N_506,N_444);
and U5503 (N_5503,N_2962,N_3843);
or U5504 (N_5504,N_4998,N_1281);
nor U5505 (N_5505,N_510,N_989);
and U5506 (N_5506,N_2834,N_562);
nand U5507 (N_5507,N_2686,N_4833);
xor U5508 (N_5508,N_4800,N_976);
or U5509 (N_5509,N_35,N_1284);
and U5510 (N_5510,N_4816,N_2218);
and U5511 (N_5511,N_1233,N_841);
nand U5512 (N_5512,N_1507,N_4602);
and U5513 (N_5513,N_4819,N_4780);
nand U5514 (N_5514,N_2082,N_3307);
nor U5515 (N_5515,N_3562,N_194);
and U5516 (N_5516,N_2820,N_2918);
nor U5517 (N_5517,N_2356,N_3348);
or U5518 (N_5518,N_3625,N_1988);
xnor U5519 (N_5519,N_535,N_3695);
xor U5520 (N_5520,N_33,N_3718);
or U5521 (N_5521,N_3767,N_2755);
xor U5522 (N_5522,N_855,N_3505);
or U5523 (N_5523,N_4281,N_3410);
and U5524 (N_5524,N_1264,N_742);
or U5525 (N_5525,N_4531,N_3113);
and U5526 (N_5526,N_4443,N_2230);
and U5527 (N_5527,N_413,N_2437);
or U5528 (N_5528,N_2738,N_2188);
and U5529 (N_5529,N_1826,N_1480);
and U5530 (N_5530,N_4524,N_4450);
nor U5531 (N_5531,N_3783,N_810);
and U5532 (N_5532,N_1309,N_1785);
nor U5533 (N_5533,N_1665,N_3008);
xnor U5534 (N_5534,N_2981,N_2470);
nand U5535 (N_5535,N_3431,N_4093);
nand U5536 (N_5536,N_245,N_143);
nand U5537 (N_5537,N_3954,N_709);
and U5538 (N_5538,N_3905,N_4387);
or U5539 (N_5539,N_502,N_2169);
nor U5540 (N_5540,N_1061,N_1197);
nand U5541 (N_5541,N_1602,N_3036);
and U5542 (N_5542,N_3417,N_2116);
or U5543 (N_5543,N_3300,N_904);
nand U5544 (N_5544,N_3975,N_1116);
nand U5545 (N_5545,N_4584,N_1588);
or U5546 (N_5546,N_2092,N_3100);
nand U5547 (N_5547,N_3646,N_1705);
and U5548 (N_5548,N_3331,N_428);
nand U5549 (N_5549,N_2691,N_949);
and U5550 (N_5550,N_1587,N_1989);
or U5551 (N_5551,N_2418,N_3217);
nor U5552 (N_5552,N_711,N_1574);
nor U5553 (N_5553,N_2601,N_2909);
nand U5554 (N_5554,N_38,N_3109);
nand U5555 (N_5555,N_3426,N_3515);
and U5556 (N_5556,N_3542,N_3232);
and U5557 (N_5557,N_4840,N_4906);
nand U5558 (N_5558,N_4049,N_1299);
or U5559 (N_5559,N_4346,N_2294);
or U5560 (N_5560,N_1795,N_3610);
and U5561 (N_5561,N_1936,N_3756);
or U5562 (N_5562,N_3384,N_778);
xor U5563 (N_5563,N_526,N_769);
nand U5564 (N_5564,N_3564,N_3669);
xor U5565 (N_5565,N_2654,N_2949);
or U5566 (N_5566,N_1985,N_3757);
nand U5567 (N_5567,N_292,N_3988);
nand U5568 (N_5568,N_3501,N_666);
xnor U5569 (N_5569,N_2193,N_3347);
nand U5570 (N_5570,N_246,N_2056);
nand U5571 (N_5571,N_2659,N_4422);
or U5572 (N_5572,N_4129,N_1538);
nor U5573 (N_5573,N_2296,N_1304);
and U5574 (N_5574,N_2359,N_3773);
or U5575 (N_5575,N_3852,N_1711);
xnor U5576 (N_5576,N_2385,N_4784);
and U5577 (N_5577,N_4574,N_1981);
nor U5578 (N_5578,N_802,N_3158);
and U5579 (N_5579,N_339,N_3482);
nor U5580 (N_5580,N_4040,N_3320);
and U5581 (N_5581,N_4454,N_3723);
and U5582 (N_5582,N_255,N_3459);
or U5583 (N_5583,N_3719,N_4141);
nand U5584 (N_5584,N_3677,N_3075);
and U5585 (N_5585,N_1242,N_107);
nor U5586 (N_5586,N_4931,N_62);
nor U5587 (N_5587,N_4014,N_3762);
xnor U5588 (N_5588,N_731,N_4991);
nand U5589 (N_5589,N_2241,N_1387);
xor U5590 (N_5590,N_569,N_4760);
xor U5591 (N_5591,N_2613,N_4986);
or U5592 (N_5592,N_2993,N_1607);
and U5593 (N_5593,N_1805,N_4073);
and U5594 (N_5594,N_643,N_4529);
xor U5595 (N_5595,N_2201,N_4605);
nor U5596 (N_5596,N_1520,N_3642);
and U5597 (N_5597,N_1036,N_2403);
and U5598 (N_5598,N_4230,N_2761);
nand U5599 (N_5599,N_1526,N_3553);
or U5600 (N_5600,N_564,N_4686);
and U5601 (N_5601,N_4576,N_1302);
xnor U5602 (N_5602,N_182,N_3014);
nand U5603 (N_5603,N_3357,N_3911);
or U5604 (N_5604,N_4546,N_4555);
and U5605 (N_5605,N_953,N_4359);
or U5606 (N_5606,N_2380,N_4208);
nor U5607 (N_5607,N_3931,N_3815);
nand U5608 (N_5608,N_1770,N_3492);
xnor U5609 (N_5609,N_3626,N_697);
xor U5610 (N_5610,N_817,N_1272);
or U5611 (N_5611,N_4650,N_2429);
xor U5612 (N_5612,N_735,N_2249);
or U5613 (N_5613,N_692,N_4112);
or U5614 (N_5614,N_1734,N_3589);
nand U5615 (N_5615,N_276,N_1976);
nor U5616 (N_5616,N_4841,N_664);
xnor U5617 (N_5617,N_293,N_2599);
or U5618 (N_5618,N_1860,N_4254);
and U5619 (N_5619,N_4837,N_1293);
and U5620 (N_5620,N_4974,N_1415);
or U5621 (N_5621,N_4826,N_4461);
or U5622 (N_5622,N_3138,N_1993);
nor U5623 (N_5623,N_2254,N_4070);
or U5624 (N_5624,N_1953,N_3266);
nor U5625 (N_5625,N_2150,N_725);
nand U5626 (N_5626,N_2919,N_2143);
and U5627 (N_5627,N_1669,N_3831);
or U5628 (N_5628,N_4613,N_3738);
nand U5629 (N_5629,N_2720,N_836);
or U5630 (N_5630,N_2713,N_4039);
nand U5631 (N_5631,N_3765,N_3604);
nor U5632 (N_5632,N_1854,N_3524);
nor U5633 (N_5633,N_93,N_1613);
nand U5634 (N_5634,N_252,N_3886);
or U5635 (N_5635,N_4782,N_4001);
or U5636 (N_5636,N_1893,N_1720);
and U5637 (N_5637,N_934,N_375);
or U5638 (N_5638,N_4740,N_3523);
nor U5639 (N_5639,N_2476,N_2002);
nand U5640 (N_5640,N_2475,N_54);
xor U5641 (N_5641,N_4879,N_2122);
or U5642 (N_5642,N_470,N_2128);
nor U5643 (N_5643,N_3715,N_4398);
nor U5644 (N_5644,N_4117,N_4999);
nor U5645 (N_5645,N_4224,N_2329);
nor U5646 (N_5646,N_630,N_710);
xnor U5647 (N_5647,N_1361,N_1210);
nor U5648 (N_5648,N_2591,N_2021);
nor U5649 (N_5649,N_405,N_2632);
and U5650 (N_5650,N_3277,N_488);
nand U5651 (N_5651,N_174,N_587);
nand U5652 (N_5652,N_4245,N_1550);
or U5653 (N_5653,N_4029,N_277);
xor U5654 (N_5654,N_1528,N_1110);
or U5655 (N_5655,N_2522,N_4249);
or U5656 (N_5656,N_4623,N_2743);
nand U5657 (N_5657,N_663,N_4883);
and U5658 (N_5658,N_2708,N_1963);
xnor U5659 (N_5659,N_2413,N_3456);
nand U5660 (N_5660,N_1928,N_2732);
nor U5661 (N_5661,N_4693,N_1251);
or U5662 (N_5662,N_1687,N_838);
xnor U5663 (N_5663,N_96,N_256);
nor U5664 (N_5664,N_4366,N_4763);
and U5665 (N_5665,N_2896,N_1627);
and U5666 (N_5666,N_2641,N_3494);
nand U5667 (N_5667,N_636,N_1022);
or U5668 (N_5668,N_2764,N_2536);
or U5669 (N_5669,N_1077,N_285);
nand U5670 (N_5670,N_2135,N_4764);
and U5671 (N_5671,N_1799,N_3161);
nor U5672 (N_5672,N_1784,N_4951);
nand U5673 (N_5673,N_3658,N_2735);
or U5674 (N_5674,N_2609,N_4661);
nor U5675 (N_5675,N_3169,N_580);
nand U5676 (N_5676,N_3004,N_1195);
and U5677 (N_5677,N_1957,N_2174);
nor U5678 (N_5678,N_683,N_2395);
nand U5679 (N_5679,N_2593,N_4511);
nand U5680 (N_5680,N_1578,N_1225);
nand U5681 (N_5681,N_570,N_1383);
nor U5682 (N_5682,N_2489,N_3030);
nand U5683 (N_5683,N_4187,N_4058);
nor U5684 (N_5684,N_1950,N_966);
nor U5685 (N_5685,N_2745,N_2793);
and U5686 (N_5686,N_4324,N_1202);
or U5687 (N_5687,N_4969,N_319);
nor U5688 (N_5688,N_1329,N_1120);
nand U5689 (N_5689,N_2242,N_2173);
and U5690 (N_5690,N_4313,N_721);
and U5691 (N_5691,N_1692,N_4971);
nand U5692 (N_5692,N_4875,N_3071);
or U5693 (N_5693,N_4958,N_2512);
and U5694 (N_5694,N_4074,N_1470);
and U5695 (N_5695,N_223,N_895);
nand U5696 (N_5696,N_4300,N_145);
xor U5697 (N_5697,N_3408,N_4099);
and U5698 (N_5698,N_605,N_169);
and U5699 (N_5699,N_4552,N_4385);
nand U5700 (N_5700,N_2948,N_199);
and U5701 (N_5701,N_3935,N_2191);
or U5702 (N_5702,N_2414,N_4590);
or U5703 (N_5703,N_4588,N_381);
xnor U5704 (N_5704,N_4720,N_3223);
or U5705 (N_5705,N_3498,N_2132);
and U5706 (N_5706,N_1288,N_4431);
and U5707 (N_5707,N_1871,N_752);
nor U5708 (N_5708,N_4309,N_3200);
nor U5709 (N_5709,N_98,N_3897);
nor U5710 (N_5710,N_3632,N_2872);
nand U5711 (N_5711,N_165,N_2392);
nor U5712 (N_5712,N_2238,N_3441);
or U5713 (N_5713,N_3925,N_3195);
or U5714 (N_5714,N_269,N_1568);
nor U5715 (N_5715,N_4199,N_3414);
nand U5716 (N_5716,N_3166,N_1243);
nor U5717 (N_5717,N_1196,N_3238);
and U5718 (N_5718,N_3029,N_3681);
nor U5719 (N_5719,N_2880,N_2432);
nand U5720 (N_5720,N_3218,N_296);
nor U5721 (N_5721,N_2318,N_3933);
or U5722 (N_5722,N_4799,N_4108);
nor U5723 (N_5723,N_172,N_4449);
and U5724 (N_5724,N_2071,N_3982);
nor U5725 (N_5725,N_863,N_4370);
nand U5726 (N_5726,N_4735,N_4635);
or U5727 (N_5727,N_3424,N_1856);
nand U5728 (N_5728,N_1261,N_3934);
nand U5729 (N_5729,N_1424,N_369);
or U5730 (N_5730,N_1859,N_1836);
and U5731 (N_5731,N_2222,N_3652);
nor U5732 (N_5732,N_4874,N_2630);
nor U5733 (N_5733,N_739,N_3440);
and U5734 (N_5734,N_450,N_3416);
and U5735 (N_5735,N_2509,N_2042);
or U5736 (N_5736,N_2204,N_4575);
and U5737 (N_5737,N_3659,N_261);
or U5738 (N_5738,N_3089,N_4862);
nor U5739 (N_5739,N_3580,N_1136);
xor U5740 (N_5740,N_2952,N_4124);
nor U5741 (N_5741,N_1846,N_1628);
or U5742 (N_5742,N_3177,N_4706);
nand U5743 (N_5743,N_3532,N_2439);
nor U5744 (N_5744,N_3326,N_1469);
nand U5745 (N_5745,N_1521,N_1181);
nor U5746 (N_5746,N_936,N_532);
and U5747 (N_5747,N_3813,N_4034);
or U5748 (N_5748,N_585,N_1258);
and U5749 (N_5749,N_640,N_1902);
nand U5750 (N_5750,N_295,N_4930);
and U5751 (N_5751,N_4560,N_4340);
and U5752 (N_5752,N_819,N_1464);
and U5753 (N_5753,N_950,N_2149);
xor U5754 (N_5754,N_3907,N_3879);
nor U5755 (N_5755,N_3335,N_1109);
or U5756 (N_5756,N_2821,N_3844);
and U5757 (N_5757,N_1872,N_4845);
or U5758 (N_5758,N_4,N_2513);
and U5759 (N_5759,N_3847,N_3777);
nand U5760 (N_5760,N_1310,N_2093);
and U5761 (N_5761,N_4417,N_637);
and U5762 (N_5762,N_306,N_3317);
nand U5763 (N_5763,N_4639,N_2393);
or U5764 (N_5764,N_4490,N_1891);
nand U5765 (N_5765,N_3780,N_4412);
and U5766 (N_5766,N_3860,N_1582);
nor U5767 (N_5767,N_3400,N_214);
and U5768 (N_5768,N_2196,N_3112);
nor U5769 (N_5769,N_784,N_3174);
xor U5770 (N_5770,N_3912,N_3140);
nand U5771 (N_5771,N_629,N_1463);
nor U5772 (N_5772,N_3885,N_947);
nor U5773 (N_5773,N_2183,N_4804);
or U5774 (N_5774,N_2103,N_4715);
nor U5775 (N_5775,N_700,N_4665);
nor U5776 (N_5776,N_2519,N_1584);
or U5777 (N_5777,N_4932,N_1645);
nand U5778 (N_5778,N_3876,N_4778);
nor U5779 (N_5779,N_4212,N_259);
nor U5780 (N_5780,N_2768,N_3923);
xor U5781 (N_5781,N_4670,N_4032);
and U5782 (N_5782,N_1960,N_1247);
nand U5783 (N_5783,N_1997,N_4131);
or U5784 (N_5784,N_2592,N_750);
nand U5785 (N_5785,N_2965,N_350);
nand U5786 (N_5786,N_2787,N_3854);
or U5787 (N_5787,N_694,N_2309);
or U5788 (N_5788,N_1847,N_195);
nor U5789 (N_5789,N_4400,N_4282);
and U5790 (N_5790,N_2077,N_2644);
nand U5791 (N_5791,N_3995,N_4054);
nand U5792 (N_5792,N_1442,N_1983);
nor U5793 (N_5793,N_1176,N_4077);
nor U5794 (N_5794,N_3228,N_751);
or U5795 (N_5795,N_2374,N_3047);
nor U5796 (N_5796,N_4183,N_1204);
xor U5797 (N_5797,N_274,N_3449);
nand U5798 (N_5798,N_3211,N_4729);
or U5799 (N_5799,N_281,N_1131);
nand U5800 (N_5800,N_4239,N_2860);
or U5801 (N_5801,N_787,N_3856);
and U5802 (N_5802,N_931,N_4959);
xnor U5803 (N_5803,N_2182,N_1646);
or U5804 (N_5804,N_964,N_2897);
and U5805 (N_5805,N_4994,N_3323);
or U5806 (N_5806,N_2134,N_2687);
or U5807 (N_5807,N_2121,N_3119);
and U5808 (N_5808,N_2404,N_525);
xor U5809 (N_5809,N_366,N_1040);
and U5810 (N_5810,N_1009,N_1445);
xor U5811 (N_5811,N_2185,N_4975);
xnor U5812 (N_5812,N_820,N_4241);
and U5813 (N_5813,N_608,N_4081);
and U5814 (N_5814,N_4852,N_2411);
and U5815 (N_5815,N_4513,N_4087);
or U5816 (N_5816,N_2759,N_515);
nor U5817 (N_5817,N_837,N_4942);
nor U5818 (N_5818,N_2670,N_4330);
nand U5819 (N_5819,N_3990,N_4355);
or U5820 (N_5820,N_4538,N_1725);
nand U5821 (N_5821,N_3924,N_3495);
nand U5822 (N_5822,N_260,N_1076);
nor U5823 (N_5823,N_3280,N_1595);
or U5824 (N_5824,N_301,N_3623);
xor U5825 (N_5825,N_4045,N_1697);
and U5826 (N_5826,N_672,N_2101);
or U5827 (N_5827,N_3792,N_1327);
nand U5828 (N_5828,N_4922,N_2700);
nor U5829 (N_5829,N_2579,N_106);
nor U5830 (N_5830,N_2096,N_755);
and U5831 (N_5831,N_2123,N_1017);
xor U5832 (N_5832,N_2590,N_1259);
nor U5833 (N_5833,N_3010,N_1755);
nor U5834 (N_5834,N_2423,N_74);
and U5835 (N_5835,N_271,N_3493);
nor U5836 (N_5836,N_1279,N_484);
or U5837 (N_5837,N_2234,N_3191);
and U5838 (N_5838,N_4295,N_1529);
or U5839 (N_5839,N_1961,N_4714);
and U5840 (N_5840,N_1714,N_1326);
or U5841 (N_5841,N_3747,N_684);
nand U5842 (N_5842,N_2620,N_4303);
nand U5843 (N_5843,N_4076,N_631);
xnor U5844 (N_5844,N_2063,N_1400);
nand U5845 (N_5845,N_249,N_3557);
nand U5846 (N_5846,N_3839,N_1699);
nand U5847 (N_5847,N_4773,N_1565);
nand U5848 (N_5848,N_956,N_560);
or U5849 (N_5849,N_565,N_4724);
nor U5850 (N_5850,N_1776,N_1140);
nand U5851 (N_5851,N_2791,N_1556);
or U5852 (N_5852,N_2541,N_1696);
xor U5853 (N_5853,N_4397,N_503);
or U5854 (N_5854,N_4292,N_3577);
and U5855 (N_5855,N_2503,N_1147);
nand U5856 (N_5856,N_3267,N_1151);
and U5857 (N_5857,N_567,N_4904);
and U5858 (N_5858,N_1282,N_1765);
nor U5859 (N_5859,N_4936,N_2505);
xnor U5860 (N_5860,N_393,N_2994);
and U5861 (N_5861,N_3638,N_1941);
nor U5862 (N_5862,N_1824,N_10);
and U5863 (N_5863,N_941,N_3592);
or U5864 (N_5864,N_2769,N_4562);
or U5865 (N_5865,N_2752,N_3084);
and U5866 (N_5866,N_648,N_18);
nor U5867 (N_5867,N_1832,N_2162);
or U5868 (N_5868,N_2278,N_3199);
or U5869 (N_5869,N_1256,N_414);
nand U5870 (N_5870,N_813,N_4898);
and U5871 (N_5871,N_924,N_1949);
nand U5872 (N_5872,N_1484,N_3183);
or U5873 (N_5873,N_681,N_3306);
nand U5874 (N_5874,N_4033,N_889);
nor U5875 (N_5875,N_4294,N_471);
or U5876 (N_5876,N_4624,N_2438);
and U5877 (N_5877,N_1067,N_477);
or U5878 (N_5878,N_3910,N_862);
nand U5879 (N_5879,N_894,N_3198);
nand U5880 (N_5880,N_2595,N_729);
xnor U5881 (N_5881,N_3086,N_3356);
or U5882 (N_5882,N_1515,N_4563);
nor U5883 (N_5883,N_327,N_312);
nand U5884 (N_5884,N_674,N_2510);
nor U5885 (N_5885,N_1636,N_4000);
and U5886 (N_5886,N_263,N_3455);
nor U5887 (N_5887,N_2929,N_3786);
xor U5888 (N_5888,N_2574,N_66);
nand U5889 (N_5889,N_3105,N_4973);
nand U5890 (N_5890,N_87,N_4988);
or U5891 (N_5891,N_4909,N_202);
nand U5892 (N_5892,N_1430,N_1439);
nand U5893 (N_5893,N_4596,N_4056);
nor U5894 (N_5894,N_4520,N_1801);
and U5895 (N_5895,N_4113,N_4415);
nor U5896 (N_5896,N_4503,N_3098);
nand U5897 (N_5897,N_356,N_4701);
nand U5898 (N_5898,N_2486,N_1850);
or U5899 (N_5899,N_4522,N_449);
and U5900 (N_5900,N_2815,N_2863);
nand U5901 (N_5901,N_459,N_4145);
and U5902 (N_5902,N_3358,N_2270);
nand U5903 (N_5903,N_575,N_2773);
or U5904 (N_5904,N_3575,N_1486);
nor U5905 (N_5905,N_1322,N_4406);
or U5906 (N_5906,N_3241,N_3985);
or U5907 (N_5907,N_4301,N_4977);
and U5908 (N_5908,N_4776,N_833);
nor U5909 (N_5909,N_2030,N_875);
or U5910 (N_5910,N_3717,N_4008);
nand U5911 (N_5911,N_1652,N_685);
or U5912 (N_5912,N_4151,N_3551);
nand U5913 (N_5913,N_2672,N_760);
nor U5914 (N_5914,N_3536,N_2225);
and U5915 (N_5915,N_3627,N_2237);
and U5916 (N_5916,N_919,N_3572);
xor U5917 (N_5917,N_3377,N_3643);
nor U5918 (N_5918,N_4085,N_929);
or U5919 (N_5919,N_3221,N_3759);
nand U5920 (N_5920,N_364,N_679);
or U5921 (N_5921,N_4642,N_2705);
nand U5922 (N_5922,N_72,N_4500);
or U5923 (N_5923,N_224,N_2890);
and U5924 (N_5924,N_2496,N_2003);
or U5925 (N_5925,N_3003,N_4527);
nor U5926 (N_5926,N_1958,N_1192);
and U5927 (N_5927,N_1883,N_3127);
nor U5928 (N_5928,N_3115,N_3556);
or U5929 (N_5929,N_4842,N_1987);
nand U5930 (N_5930,N_2050,N_2967);
nand U5931 (N_5931,N_3404,N_4376);
nand U5932 (N_5932,N_4506,N_1048);
nand U5933 (N_5933,N_4652,N_3798);
xnor U5934 (N_5934,N_3157,N_2124);
nor U5935 (N_5935,N_24,N_25);
or U5936 (N_5936,N_2477,N_1244);
xor U5937 (N_5937,N_1101,N_3050);
nor U5938 (N_5938,N_2879,N_395);
and U5939 (N_5939,N_4918,N_3028);
and U5940 (N_5940,N_2699,N_1540);
or U5941 (N_5941,N_147,N_3246);
or U5942 (N_5942,N_3210,N_2259);
and U5943 (N_5943,N_3205,N_4734);
or U5944 (N_5944,N_2701,N_1295);
and U5945 (N_5945,N_43,N_2275);
nand U5946 (N_5946,N_610,N_3106);
and U5947 (N_5947,N_632,N_485);
and U5948 (N_5948,N_720,N_49);
or U5949 (N_5949,N_1581,N_3308);
and U5950 (N_5950,N_3187,N_2348);
or U5951 (N_5951,N_2430,N_4246);
nor U5952 (N_5952,N_3120,N_4111);
nor U5953 (N_5953,N_1212,N_2246);
xor U5954 (N_5954,N_4488,N_4259);
nand U5955 (N_5955,N_2792,N_2577);
nor U5956 (N_5956,N_3618,N_1103);
or U5957 (N_5957,N_1375,N_2539);
or U5958 (N_5958,N_181,N_4459);
or U5959 (N_5959,N_4556,N_3212);
and U5960 (N_5960,N_4620,N_4421);
or U5961 (N_5961,N_125,N_2570);
or U5962 (N_5962,N_4846,N_1547);
and U5963 (N_5963,N_2645,N_2095);
or U5964 (N_5964,N_2521,N_480);
and U5965 (N_5965,N_4288,N_1747);
and U5966 (N_5966,N_3474,N_3647);
and U5967 (N_5967,N_981,N_1265);
or U5968 (N_5968,N_1191,N_1016);
nand U5969 (N_5969,N_2597,N_1661);
and U5970 (N_5970,N_1063,N_1681);
and U5971 (N_5971,N_132,N_1739);
or U5972 (N_5972,N_1126,N_2100);
nor U5973 (N_5973,N_4418,N_4357);
and U5974 (N_5974,N_1420,N_785);
or U5975 (N_5975,N_3909,N_4688);
nand U5976 (N_5976,N_1788,N_3422);
and U5977 (N_5977,N_4136,N_2054);
nor U5978 (N_5978,N_1688,N_650);
nor U5979 (N_5979,N_844,N_2995);
nor U5980 (N_5980,N_2228,N_3362);
or U5981 (N_5981,N_1058,N_2741);
nand U5982 (N_5982,N_343,N_3744);
or U5983 (N_5983,N_4363,N_1787);
nand U5984 (N_5984,N_2862,N_3065);
or U5985 (N_5985,N_600,N_4935);
xor U5986 (N_5986,N_4227,N_3797);
nor U5987 (N_5987,N_4403,N_2431);
nor U5988 (N_5988,N_1338,N_4880);
nand U5989 (N_5989,N_2427,N_284);
and U5990 (N_5990,N_4458,N_4419);
or U5991 (N_5991,N_108,N_487);
nor U5992 (N_5992,N_1557,N_1662);
nor U5993 (N_5993,N_1004,N_2562);
and U5994 (N_5994,N_122,N_1178);
nor U5995 (N_5995,N_3253,N_1986);
nor U5996 (N_5996,N_4889,N_3836);
and U5997 (N_5997,N_4125,N_4687);
and U5998 (N_5998,N_4753,N_2112);
nand U5999 (N_5999,N_3710,N_1080);
or U6000 (N_6000,N_2322,N_4184);
and U6001 (N_6001,N_3388,N_4473);
nand U6002 (N_6002,N_498,N_4896);
nand U6003 (N_6003,N_687,N_3992);
nor U6004 (N_6004,N_3741,N_1097);
or U6005 (N_6005,N_1359,N_492);
nand U6006 (N_6006,N_1921,N_995);
or U6007 (N_6007,N_439,N_168);
or U6008 (N_6008,N_430,N_2886);
xnor U6009 (N_6009,N_2709,N_1591);
or U6010 (N_6010,N_1830,N_2526);
nand U6011 (N_6011,N_1685,N_2245);
nand U6012 (N_6012,N_918,N_4475);
nor U6013 (N_6013,N_3445,N_2647);
xnor U6014 (N_6014,N_3561,N_2665);
or U6015 (N_6015,N_81,N_1994);
xor U6016 (N_6016,N_2934,N_2883);
nor U6017 (N_6017,N_3692,N_1095);
and U6018 (N_6018,N_4887,N_3770);
nand U6019 (N_6019,N_2680,N_2308);
nand U6020 (N_6020,N_4102,N_3247);
nor U6021 (N_6021,N_1870,N_1710);
or U6022 (N_6022,N_1853,N_29);
xor U6023 (N_6023,N_452,N_3471);
and U6024 (N_6024,N_2478,N_4830);
and U6025 (N_6025,N_4298,N_354);
nand U6026 (N_6026,N_1852,N_3243);
nor U6027 (N_6027,N_2001,N_3570);
nor U6028 (N_6028,N_3273,N_3152);
and U6029 (N_6029,N_4869,N_3460);
nor U6030 (N_6030,N_3936,N_991);
nor U6031 (N_6031,N_2479,N_2874);
nor U6032 (N_6032,N_3165,N_1980);
or U6033 (N_6033,N_1234,N_724);
nand U6034 (N_6034,N_3311,N_2231);
xnor U6035 (N_6035,N_1157,N_4336);
and U6036 (N_6036,N_1039,N_726);
and U6037 (N_6037,N_1641,N_2032);
or U6038 (N_6038,N_982,N_3674);
and U6039 (N_6039,N_1898,N_1633);
and U6040 (N_6040,N_1704,N_3605);
nand U6041 (N_6041,N_1215,N_3508);
and U6042 (N_6042,N_4266,N_3957);
nor U6043 (N_6043,N_3136,N_4314);
nor U6044 (N_6044,N_1056,N_4619);
and U6045 (N_6045,N_1709,N_1005);
and U6046 (N_6046,N_1807,N_3462);
nor U6047 (N_6047,N_3466,N_2194);
and U6048 (N_6048,N_1479,N_1427);
and U6049 (N_6049,N_4360,N_4927);
or U6050 (N_6050,N_1489,N_2850);
nand U6051 (N_6051,N_4884,N_2219);
and U6052 (N_6052,N_4989,N_4929);
nand U6053 (N_6053,N_3451,N_2810);
and U6054 (N_6054,N_1290,N_588);
or U6055 (N_6055,N_3088,N_1903);
or U6056 (N_6056,N_4456,N_2928);
nor U6057 (N_6057,N_1786,N_1828);
nand U6058 (N_6058,N_3015,N_1292);
or U6059 (N_6059,N_910,N_1121);
nor U6060 (N_6060,N_4036,N_76);
nor U6061 (N_6061,N_3963,N_1938);
and U6062 (N_6062,N_4941,N_2091);
xnor U6063 (N_6063,N_4375,N_4468);
nor U6064 (N_6064,N_2400,N_3841);
nand U6065 (N_6065,N_3835,N_2272);
nand U6066 (N_6066,N_345,N_1844);
and U6067 (N_6067,N_2504,N_2078);
or U6068 (N_6068,N_887,N_2681);
xnor U6069 (N_6069,N_3270,N_4843);
nor U6070 (N_6070,N_215,N_583);
or U6071 (N_6071,N_2494,N_2583);
or U6072 (N_6072,N_1465,N_759);
nand U6073 (N_6073,N_387,N_1477);
and U6074 (N_6074,N_3964,N_203);
nand U6075 (N_6075,N_3941,N_2618);
nor U6076 (N_6076,N_2288,N_363);
nand U6077 (N_6077,N_539,N_3437);
nor U6078 (N_6078,N_662,N_3868);
xor U6079 (N_6079,N_3182,N_2059);
nand U6080 (N_6080,N_3746,N_4868);
nor U6081 (N_6081,N_3316,N_797);
or U6082 (N_6082,N_1074,N_4244);
nor U6083 (N_6083,N_36,N_4578);
nor U6084 (N_6084,N_4190,N_4159);
nand U6085 (N_6085,N_39,N_1866);
and U6086 (N_6086,N_2164,N_2138);
and U6087 (N_6087,N_970,N_3734);
or U6088 (N_6088,N_2668,N_3057);
nand U6089 (N_6089,N_2307,N_308);
nand U6090 (N_6090,N_658,N_216);
or U6091 (N_6091,N_1724,N_746);
or U6092 (N_6092,N_1911,N_1454);
or U6093 (N_6093,N_3682,N_2664);
or U6094 (N_6094,N_2131,N_4737);
nand U6095 (N_6095,N_466,N_4616);
and U6096 (N_6096,N_2744,N_878);
nand U6097 (N_6097,N_68,N_3529);
nor U6098 (N_6098,N_4718,N_433);
nor U6099 (N_6099,N_2256,N_61);
and U6100 (N_6100,N_4139,N_4236);
nor U6101 (N_6101,N_4146,N_2017);
nand U6102 (N_6102,N_2184,N_2419);
xor U6103 (N_6103,N_2445,N_541);
and U6104 (N_6104,N_2453,N_821);
or U6105 (N_6105,N_3423,N_2662);
and U6106 (N_6106,N_4368,N_783);
or U6107 (N_6107,N_1342,N_3292);
nor U6108 (N_6108,N_1796,N_2818);
or U6109 (N_6109,N_1395,N_2544);
or U6110 (N_6110,N_2398,N_3173);
or U6111 (N_6111,N_3945,N_3881);
nand U6112 (N_6112,N_4672,N_307);
or U6113 (N_6113,N_3181,N_4082);
xnor U6114 (N_6114,N_3093,N_3960);
xnor U6115 (N_6115,N_911,N_3133);
and U6116 (N_6116,N_3644,N_4150);
and U6117 (N_6117,N_2925,N_747);
and U6118 (N_6118,N_4549,N_1597);
xor U6119 (N_6119,N_4114,N_4016);
or U6120 (N_6120,N_3791,N_1399);
xor U6121 (N_6121,N_2145,N_4675);
and U6122 (N_6122,N_2692,N_4427);
and U6123 (N_6123,N_149,N_2747);
or U6124 (N_6124,N_3882,N_3151);
nor U6125 (N_6125,N_3633,N_1656);
or U6126 (N_6126,N_3491,N_2416);
nor U6127 (N_6127,N_1448,N_3981);
or U6128 (N_6128,N_2617,N_1180);
nor U6129 (N_6129,N_969,N_3962);
or U6130 (N_6130,N_1554,N_20);
or U6131 (N_6131,N_3884,N_3176);
nor U6132 (N_6132,N_4983,N_4523);
xor U6133 (N_6133,N_4411,N_555);
and U6134 (N_6134,N_2331,N_3022);
nand U6135 (N_6135,N_4464,N_2425);
and U6136 (N_6136,N_3250,N_753);
and U6137 (N_6137,N_2177,N_1990);
or U6138 (N_6138,N_2760,N_3895);
nor U6139 (N_6139,N_1184,N_4723);
nand U6140 (N_6140,N_2584,N_3160);
nor U6141 (N_6141,N_142,N_463);
nand U6142 (N_6142,N_2114,N_1823);
or U6143 (N_6143,N_2604,N_4134);
nand U6144 (N_6144,N_3754,N_222);
and U6145 (N_6145,N_2209,N_1374);
and U6146 (N_6146,N_812,N_2675);
or U6147 (N_6147,N_3124,N_892);
nand U6148 (N_6148,N_4629,N_1328);
nand U6149 (N_6149,N_1815,N_1524);
and U6150 (N_6150,N_2853,N_3663);
nor U6151 (N_6151,N_1119,N_329);
and U6152 (N_6152,N_1163,N_1885);
nand U6153 (N_6153,N_3694,N_2224);
nor U6154 (N_6154,N_915,N_1402);
nor U6155 (N_6155,N_3699,N_1611);
nor U6156 (N_6156,N_4168,N_4219);
nor U6157 (N_6157,N_4329,N_2153);
xor U6158 (N_6158,N_903,N_0);
nand U6159 (N_6159,N_2794,N_4291);
nor U6160 (N_6160,N_4754,N_1408);
xnor U6161 (N_6161,N_3600,N_1071);
and U6162 (N_6162,N_2725,N_479);
nor U6163 (N_6163,N_1572,N_2297);
and U6164 (N_6164,N_4953,N_2891);
and U6165 (N_6165,N_4155,N_2941);
nor U6166 (N_6166,N_3785,N_2612);
or U6167 (N_6167,N_4343,N_4772);
or U6168 (N_6168,N_4915,N_4946);
and U6169 (N_6169,N_4248,N_1360);
nor U6170 (N_6170,N_3046,N_1011);
or U6171 (N_6171,N_961,N_3141);
or U6172 (N_6172,N_1954,N_2436);
or U6173 (N_6173,N_4493,N_4765);
nor U6174 (N_6174,N_154,N_2461);
nor U6175 (N_6175,N_913,N_478);
xor U6176 (N_6176,N_4166,N_4997);
and U6177 (N_6177,N_2198,N_3240);
nor U6178 (N_6178,N_2472,N_2619);
nand U6179 (N_6179,N_4891,N_4118);
nand U6180 (N_6180,N_948,N_1708);
and U6181 (N_6181,N_3204,N_4762);
or U6182 (N_6182,N_221,N_4964);
nor U6183 (N_6183,N_2762,N_4926);
nand U6184 (N_6184,N_2363,N_3467);
nand U6185 (N_6185,N_1982,N_2066);
xor U6186 (N_6186,N_3064,N_3987);
nand U6187 (N_6187,N_2277,N_1168);
and U6188 (N_6188,N_1689,N_2111);
nor U6189 (N_6189,N_1105,N_1702);
and U6190 (N_6190,N_4585,N_2068);
nand U6191 (N_6191,N_86,N_4043);
and U6192 (N_6192,N_3330,N_1742);
or U6193 (N_6193,N_1551,N_2803);
and U6194 (N_6194,N_2542,N_1878);
and U6195 (N_6195,N_300,N_1908);
nand U6196 (N_6196,N_757,N_512);
nand U6197 (N_6197,N_3956,N_3576);
and U6198 (N_6198,N_2588,N_1466);
or U6199 (N_6199,N_2332,N_2969);
or U6200 (N_6200,N_3268,N_4152);
and U6201 (N_6201,N_2559,N_4743);
nor U6202 (N_6202,N_1440,N_2734);
nand U6203 (N_6203,N_2774,N_73);
and U6204 (N_6204,N_3432,N_1616);
xor U6205 (N_6205,N_4940,N_2866);
or U6206 (N_6206,N_4137,N_777);
nand U6207 (N_6207,N_2455,N_628);
or U6208 (N_6208,N_1296,N_4631);
and U6209 (N_6209,N_1683,N_3333);
or U6210 (N_6210,N_2351,N_3391);
and U6211 (N_6211,N_3853,N_1171);
nor U6212 (N_6212,N_2817,N_4399);
nand U6213 (N_6213,N_4388,N_708);
or U6214 (N_6214,N_162,N_2253);
nor U6215 (N_6215,N_4995,N_3657);
nor U6216 (N_6216,N_1417,N_2903);
nor U6217 (N_6217,N_3991,N_4013);
and U6218 (N_6218,N_2409,N_796);
xor U6219 (N_6219,N_2391,N_861);
nor U6220 (N_6220,N_930,N_4878);
nand U6221 (N_6221,N_429,N_2712);
xnor U6222 (N_6222,N_118,N_761);
nor U6223 (N_6223,N_3670,N_4484);
nor U6224 (N_6224,N_4536,N_3825);
and U6225 (N_6225,N_907,N_1137);
or U6226 (N_6226,N_4919,N_713);
nor U6227 (N_6227,N_4813,N_3552);
xor U6228 (N_6228,N_791,N_2069);
nor U6229 (N_6229,N_3190,N_1573);
nor U6230 (N_6230,N_198,N_2971);
or U6231 (N_6231,N_2916,N_2353);
nand U6232 (N_6232,N_942,N_335);
and U6233 (N_6233,N_1350,N_1733);
or U6234 (N_6234,N_402,N_1431);
or U6235 (N_6235,N_2199,N_1214);
nand U6236 (N_6236,N_2043,N_2378);
nor U6237 (N_6237,N_3766,N_2302);
or U6238 (N_6238,N_1851,N_4002);
or U6239 (N_6239,N_4153,N_497);
and U6240 (N_6240,N_873,N_1977);
and U6241 (N_6241,N_1541,N_4435);
and U6242 (N_6242,N_717,N_348);
and U6243 (N_6243,N_1160,N_2673);
nor U6244 (N_6244,N_3559,N_1677);
or U6245 (N_6245,N_652,N_1522);
nand U6246 (N_6246,N_3635,N_4514);
and U6247 (N_6247,N_2325,N_1211);
or U6248 (N_6248,N_3147,N_2808);
nor U6249 (N_6249,N_3526,N_2568);
nor U6250 (N_6250,N_432,N_4369);
nor U6251 (N_6251,N_1506,N_2825);
or U6252 (N_6252,N_4982,N_2751);
and U6253 (N_6253,N_2500,N_4501);
nand U6254 (N_6254,N_3731,N_3587);
or U6255 (N_6255,N_353,N_1410);
nor U6256 (N_6256,N_2334,N_3827);
nor U6257 (N_6257,N_954,N_1659);
and U6258 (N_6258,N_4010,N_1073);
or U6259 (N_6259,N_673,N_2799);
or U6260 (N_6260,N_1558,N_909);
xor U6261 (N_6261,N_4351,N_4993);
nand U6262 (N_6262,N_280,N_792);
or U6263 (N_6263,N_851,N_92);
nand U6264 (N_6264,N_2939,N_264);
nor U6265 (N_6265,N_1044,N_4831);
and U6266 (N_6266,N_2611,N_3365);
and U6267 (N_6267,N_4747,N_4952);
nand U6268 (N_6268,N_3622,N_4751);
xor U6269 (N_6269,N_1372,N_138);
xor U6270 (N_6270,N_3156,N_158);
xnor U6271 (N_6271,N_4853,N_2388);
nand U6272 (N_6272,N_3056,N_3812);
or U6273 (N_6273,N_3069,N_3011);
and U6274 (N_6274,N_2660,N_2598);
nor U6275 (N_6275,N_4834,N_1615);
nor U6276 (N_6276,N_3980,N_3571);
and U6277 (N_6277,N_4393,N_2816);
nor U6278 (N_6278,N_457,N_1102);
nand U6279 (N_6279,N_192,N_332);
or U6280 (N_6280,N_2703,N_2840);
xor U6281 (N_6281,N_1294,N_1670);
nand U6282 (N_6282,N_2006,N_3146);
nor U6283 (N_6283,N_3312,N_3943);
nand U6284 (N_6284,N_2766,N_4069);
nand U6285 (N_6285,N_4404,N_2045);
and U6286 (N_6286,N_4807,N_645);
nor U6287 (N_6287,N_1033,N_879);
nand U6288 (N_6288,N_1495,N_1154);
nand U6289 (N_6289,N_2236,N_830);
or U6290 (N_6290,N_3851,N_3566);
nand U6291 (N_6291,N_1492,N_4873);
xor U6292 (N_6292,N_1434,N_3520);
and U6293 (N_6293,N_962,N_461);
and U6294 (N_6294,N_1625,N_1043);
nand U6295 (N_6295,N_251,N_419);
nor U6296 (N_6296,N_3096,N_85);
or U6297 (N_6297,N_299,N_4201);
and U6298 (N_6298,N_1318,N_4615);
nor U6299 (N_6299,N_2697,N_524);
nor U6300 (N_6300,N_1393,N_804);
and U6301 (N_6301,N_1315,N_2822);
or U6302 (N_6302,N_1800,N_3231);
xor U6303 (N_6303,N_4028,N_2858);
nor U6304 (N_6304,N_2020,N_1366);
or U6305 (N_6305,N_1713,N_2155);
nor U6306 (N_6306,N_3899,N_422);
nand U6307 (N_6307,N_4205,N_767);
and U6308 (N_6308,N_1345,N_310);
nor U6309 (N_6309,N_1542,N_939);
nor U6310 (N_6310,N_2118,N_3544);
or U6311 (N_6311,N_3104,N_2973);
and U6312 (N_6312,N_1031,N_2706);
or U6313 (N_6313,N_431,N_4229);
or U6314 (N_6314,N_3405,N_1773);
nand U6315 (N_6315,N_1857,N_3880);
or U6316 (N_6316,N_1843,N_3435);
xnor U6317 (N_6317,N_4771,N_3081);
xnor U6318 (N_6318,N_847,N_2);
or U6319 (N_6319,N_226,N_270);
nor U6320 (N_6320,N_3027,N_1025);
nor U6321 (N_6321,N_1593,N_808);
or U6322 (N_6322,N_741,N_1280);
xnor U6323 (N_6323,N_2946,N_2473);
nor U6324 (N_6324,N_3020,N_1447);
nand U6325 (N_6325,N_3499,N_2956);
or U6326 (N_6326,N_2151,N_254);
nor U6327 (N_6327,N_3809,N_2269);
and U6328 (N_6328,N_2823,N_945);
and U6329 (N_6329,N_1979,N_2154);
and U6330 (N_6330,N_4965,N_58);
nor U6331 (N_6331,N_1576,N_1594);
and U6332 (N_6332,N_2401,N_3185);
nand U6333 (N_6333,N_166,N_4495);
or U6334 (N_6334,N_3371,N_3287);
and U6335 (N_6335,N_1274,N_3998);
or U6336 (N_6336,N_4062,N_1610);
and U6337 (N_6337,N_568,N_4902);
xor U6338 (N_6338,N_7,N_2454);
nor U6339 (N_6339,N_1855,N_4832);
or U6340 (N_6340,N_4126,N_1188);
nor U6341 (N_6341,N_626,N_2893);
nand U6342 (N_6342,N_4730,N_793);
or U6343 (N_6343,N_474,N_4750);
and U6344 (N_6344,N_4827,N_1909);
xnor U6345 (N_6345,N_2377,N_2587);
or U6346 (N_6346,N_983,N_2533);
nand U6347 (N_6347,N_2126,N_4696);
xor U6348 (N_6348,N_1512,N_4321);
and U6349 (N_6349,N_1134,N_3846);
and U6350 (N_6350,N_1549,N_2770);
nor U6351 (N_6351,N_2910,N_3168);
nand U6352 (N_6352,N_4323,N_4966);
and U6353 (N_6353,N_763,N_4610);
nand U6354 (N_6354,N_870,N_1943);
and U6355 (N_6355,N_2310,N_3878);
or U6356 (N_6356,N_3438,N_213);
nor U6357 (N_6357,N_3428,N_1229);
nor U6358 (N_6358,N_2217,N_4448);
and U6359 (N_6359,N_1605,N_2804);
and U6360 (N_6360,N_330,N_3360);
or U6361 (N_6361,N_2572,N_1363);
nand U6362 (N_6362,N_4169,N_4571);
nor U6363 (N_6363,N_3541,N_538);
nand U6364 (N_6364,N_418,N_240);
nand U6365 (N_6365,N_2013,N_244);
or U6366 (N_6366,N_3469,N_3420);
or U6367 (N_6367,N_1837,N_3302);
and U6368 (N_6368,N_654,N_1888);
and U6369 (N_6369,N_1933,N_4943);
nand U6370 (N_6370,N_780,N_1059);
nor U6371 (N_6371,N_3671,N_2502);
nor U6372 (N_6372,N_1223,N_236);
nor U6373 (N_6373,N_2514,N_4188);
or U6374 (N_6374,N_986,N_3281);
nor U6375 (N_6375,N_398,N_2451);
and U6376 (N_6376,N_1138,N_1270);
nor U6377 (N_6377,N_3305,N_1901);
and U6378 (N_6378,N_3025,N_3051);
or U6379 (N_6379,N_2499,N_3224);
or U6380 (N_6380,N_2807,N_2417);
nor U6381 (N_6381,N_999,N_3637);
and U6382 (N_6382,N_2457,N_1703);
nor U6383 (N_6383,N_4839,N_3826);
nor U6384 (N_6384,N_1682,N_2715);
nand U6385 (N_6385,N_4609,N_2306);
or U6386 (N_6386,N_4439,N_1308);
nor U6387 (N_6387,N_4165,N_3916);
nand U6388 (N_6388,N_2596,N_2298);
nand U6389 (N_6389,N_3222,N_2152);
nand U6390 (N_6390,N_768,N_3817);
nor U6391 (N_6391,N_3913,N_1300);
and U6392 (N_6392,N_3634,N_2722);
nand U6393 (N_6393,N_2226,N_2008);
or U6394 (N_6394,N_4233,N_4820);
nor U6395 (N_6395,N_2327,N_3830);
nor U6396 (N_6396,N_4920,N_1161);
and U6397 (N_6397,N_4968,N_1812);
or U6398 (N_6398,N_3751,N_4719);
and U6399 (N_6399,N_4463,N_902);
nor U6400 (N_6400,N_2581,N_3863);
or U6401 (N_6401,N_311,N_3130);
and U6402 (N_6402,N_1864,N_795);
nor U6403 (N_6403,N_1086,N_9);
and U6404 (N_6404,N_2161,N_2689);
xor U6405 (N_6405,N_4430,N_2186);
or U6406 (N_6406,N_2290,N_427);
nand U6407 (N_6407,N_4597,N_1672);
and U6408 (N_6408,N_3955,N_4710);
and U6409 (N_6409,N_2711,N_1971);
and U6410 (N_6410,N_2690,N_3344);
xnor U6411 (N_6411,N_734,N_3742);
or U6412 (N_6412,N_2299,N_620);
nand U6413 (N_6413,N_1752,N_618);
nand U6414 (N_6414,N_2777,N_209);
and U6415 (N_6415,N_3687,N_4350);
nor U6416 (N_6416,N_1819,N_3361);
nand U6417 (N_6417,N_4685,N_57);
and U6418 (N_6418,N_1760,N_379);
nor U6419 (N_6419,N_4697,N_188);
or U6420 (N_6420,N_905,N_3484);
nand U6421 (N_6421,N_4172,N_881);
nand U6422 (N_6422,N_2264,N_3078);
or U6423 (N_6423,N_3229,N_2104);
nor U6424 (N_6424,N_592,N_756);
nor U6425 (N_6425,N_3461,N_4600);
and U6426 (N_6426,N_4090,N_2197);
xnor U6427 (N_6427,N_4890,N_2980);
nand U6428 (N_6428,N_190,N_34);
nor U6429 (N_6429,N_4618,N_4673);
nor U6430 (N_6430,N_3752,N_2136);
and U6431 (N_6431,N_1343,N_2015);
or U6432 (N_6432,N_2937,N_3932);
nor U6433 (N_6433,N_3949,N_4792);
nor U6434 (N_6434,N_2992,N_4637);
or U6435 (N_6435,N_815,N_476);
and U6436 (N_6436,N_1099,N_2323);
nor U6437 (N_6437,N_1673,N_2885);
or U6438 (N_6438,N_1432,N_2915);
or U6439 (N_6439,N_3367,N_1762);
nand U6440 (N_6440,N_495,N_2582);
nand U6441 (N_6441,N_1412,N_1289);
nor U6442 (N_6442,N_4089,N_1869);
or U6443 (N_6443,N_2920,N_3795);
xnor U6444 (N_6444,N_228,N_121);
and U6445 (N_6445,N_1185,N_1905);
or U6446 (N_6446,N_155,N_2372);
nor U6447 (N_6447,N_920,N_1822);
nor U6448 (N_6448,N_2651,N_2109);
nor U6449 (N_6449,N_2898,N_4061);
and U6450 (N_6450,N_4390,N_2065);
and U6451 (N_6451,N_1877,N_4316);
nor U6452 (N_6452,N_2532,N_2125);
and U6453 (N_6453,N_4372,N_2938);
nor U6454 (N_6454,N_2650,N_857);
nor U6455 (N_6455,N_4096,N_3628);
nand U6456 (N_6456,N_491,N_3236);
nor U6457 (N_6457,N_788,N_1068);
nand U6458 (N_6458,N_1769,N_1108);
or U6459 (N_6459,N_4367,N_2847);
and U6460 (N_6460,N_3001,N_1206);
nand U6461 (N_6461,N_4335,N_1340);
xor U6462 (N_6462,N_4626,N_486);
and U6463 (N_6463,N_170,N_4532);
and U6464 (N_6464,N_1013,N_3352);
or U6465 (N_6465,N_1504,N_1078);
and U6466 (N_6466,N_53,N_2857);
and U6467 (N_6467,N_606,N_3434);
nand U6468 (N_6468,N_4497,N_2358);
nand U6469 (N_6469,N_2211,N_4662);
or U6470 (N_6470,N_2301,N_3465);
and U6471 (N_6471,N_1750,N_1370);
nor U6472 (N_6472,N_3875,N_1996);
or U6473 (N_6473,N_267,N_2704);
nor U6474 (N_6474,N_3567,N_1045);
nand U6475 (N_6475,N_4698,N_4371);
nand U6476 (N_6476,N_3808,N_3381);
and U6477 (N_6477,N_3630,N_3972);
or U6478 (N_6478,N_2788,N_2227);
nor U6479 (N_6479,N_2935,N_4286);
nand U6480 (N_6480,N_2740,N_4234);
nand U6481 (N_6481,N_4810,N_3189);
nand U6482 (N_6482,N_4059,N_2518);
nor U6483 (N_6483,N_2495,N_2369);
nor U6484 (N_6484,N_549,N_3782);
xnor U6485 (N_6485,N_4825,N_3279);
nor U6486 (N_6486,N_2176,N_3761);
xnor U6487 (N_6487,N_591,N_4211);
nand U6488 (N_6488,N_4194,N_1317);
xnor U6489 (N_6489,N_3986,N_435);
nand U6490 (N_6490,N_3996,N_974);
nor U6491 (N_6491,N_4913,N_867);
or U6492 (N_6492,N_577,N_1728);
xnor U6493 (N_6493,N_4048,N_2627);
or U6494 (N_6494,N_2441,N_3928);
nand U6495 (N_6495,N_603,N_2990);
or U6496 (N_6496,N_1634,N_4856);
or U6497 (N_6497,N_2997,N_2076);
nand U6498 (N_6498,N_4285,N_727);
nand U6499 (N_6499,N_426,N_2749);
and U6500 (N_6500,N_4525,N_4736);
and U6501 (N_6501,N_860,N_3488);
nand U6502 (N_6502,N_3977,N_3002);
nand U6503 (N_6503,N_1904,N_4235);
and U6504 (N_6504,N_3382,N_4037);
or U6505 (N_6505,N_1332,N_1269);
and U6506 (N_6506,N_2671,N_3209);
or U6507 (N_6507,N_4322,N_2276);
or U6508 (N_6508,N_2098,N_273);
nor U6509 (N_6509,N_3349,N_3418);
nor U6510 (N_6510,N_1453,N_1089);
and U6511 (N_6511,N_1398,N_3203);
and U6512 (N_6512,N_3728,N_3865);
nor U6513 (N_6513,N_416,N_2469);
and U6514 (N_6514,N_3867,N_2447);
or U6515 (N_6515,N_2538,N_3386);
xor U6516 (N_6516,N_781,N_882);
nor U6517 (N_6517,N_3678,N_3504);
and U6518 (N_6518,N_4409,N_3442);
or U6519 (N_6519,N_2931,N_4177);
nand U6520 (N_6520,N_2870,N_2113);
and U6521 (N_6521,N_2911,N_1907);
nand U6522 (N_6522,N_467,N_3641);
xor U6523 (N_6523,N_3413,N_3070);
nand U6524 (N_6524,N_3538,N_458);
nor U6525 (N_6525,N_2730,N_4179);
and U6526 (N_6526,N_4612,N_3107);
nand U6527 (N_6527,N_1303,N_23);
nand U6528 (N_6528,N_2957,N_1564);
xor U6529 (N_6529,N_2037,N_184);
and U6530 (N_6530,N_660,N_4554);
and U6531 (N_6531,N_3588,N_689);
nor U6532 (N_6532,N_1623,N_2841);
or U6533 (N_6533,N_3376,N_2586);
xnor U6534 (N_6534,N_1096,N_164);
nor U6535 (N_6535,N_688,N_4791);
and U6536 (N_6536,N_235,N_4580);
and U6537 (N_6537,N_392,N_2639);
and U6538 (N_6538,N_3832,N_2202);
and U6539 (N_6539,N_4770,N_1535);
xnor U6540 (N_6540,N_1337,N_1218);
or U6541 (N_6541,N_762,N_3629);
and U6542 (N_6542,N_579,N_898);
nand U6543 (N_6543,N_1287,N_1187);
nor U6544 (N_6544,N_1598,N_2678);
nand U6545 (N_6545,N_2287,N_4296);
and U6546 (N_6546,N_1505,N_927);
xnor U6547 (N_6547,N_1182,N_4847);
or U6548 (N_6548,N_4220,N_4756);
nand U6549 (N_6549,N_2263,N_1079);
nor U6550 (N_6550,N_2657,N_1951);
and U6551 (N_6551,N_232,N_2633);
nand U6552 (N_6552,N_1498,N_4599);
nor U6553 (N_6553,N_323,N_2170);
or U6554 (N_6554,N_3,N_826);
or U6555 (N_6555,N_4664,N_3329);
nor U6556 (N_6556,N_357,N_2775);
and U6557 (N_6557,N_704,N_732);
nor U6558 (N_6558,N_383,N_4638);
nor U6559 (N_6559,N_468,N_2189);
nor U6560 (N_6560,N_2362,N_4457);
nor U6561 (N_6561,N_3558,N_3732);
xnor U6562 (N_6562,N_3745,N_3041);
or U6563 (N_6563,N_4690,N_3781);
nor U6564 (N_6564,N_3824,N_2347);
and U6565 (N_6565,N_4466,N_2802);
and U6566 (N_6566,N_186,N_4683);
nor U6567 (N_6567,N_4545,N_3811);
nor U6568 (N_6568,N_46,N_2467);
or U6569 (N_6569,N_4312,N_3518);
nand U6570 (N_6570,N_988,N_1654);
or U6571 (N_6571,N_4110,N_3803);
and U6572 (N_6572,N_4474,N_4401);
nor U6573 (N_6573,N_2985,N_1409);
nor U6574 (N_6574,N_1148,N_4426);
or U6575 (N_6575,N_2561,N_4018);
or U6576 (N_6576,N_4481,N_595);
nand U6577 (N_6577,N_1362,N_4251);
or U6578 (N_6578,N_4518,N_576);
nor U6579 (N_6579,N_1825,N_992);
nand U6580 (N_6580,N_4808,N_1491);
nor U6581 (N_6581,N_1875,N_3397);
or U6582 (N_6582,N_2742,N_3593);
nor U6583 (N_6583,N_2785,N_4204);
nor U6584 (N_6584,N_2344,N_4797);
nor U6585 (N_6585,N_229,N_4521);
nand U6586 (N_6586,N_2120,N_3919);
nor U6587 (N_6587,N_655,N_30);
nor U6588 (N_6588,N_1516,N_401);
xnor U6589 (N_6589,N_1054,N_4512);
or U6590 (N_6590,N_2868,N_342);
or U6591 (N_6591,N_3993,N_2160);
nand U6592 (N_6592,N_1169,N_1579);
or U6593 (N_6593,N_2778,N_4822);
and U6594 (N_6594,N_2379,N_4072);
or U6595 (N_6595,N_4260,N_2468);
xnor U6596 (N_6596,N_4577,N_4558);
nor U6597 (N_6597,N_4899,N_2171);
nor U6598 (N_6598,N_88,N_6);
and U6599 (N_6599,N_3989,N_2481);
nor U6600 (N_6600,N_3463,N_3296);
nor U6601 (N_6601,N_4550,N_2097);
nand U6602 (N_6602,N_4218,N_4257);
or U6603 (N_6603,N_3519,N_3820);
and U6604 (N_6604,N_1297,N_4866);
or U6605 (N_6605,N_4802,N_3082);
and U6606 (N_6606,N_3297,N_2966);
and U6607 (N_6607,N_3477,N_4787);
and U6608 (N_6608,N_3776,N_854);
nand U6609 (N_6609,N_4467,N_2606);
or U6610 (N_6610,N_2335,N_1421);
nand U6611 (N_6611,N_744,N_3394);
and U6612 (N_6612,N_4708,N_3207);
nor U6613 (N_6613,N_1376,N_1748);
nand U6614 (N_6614,N_4829,N_2450);
or U6615 (N_6615,N_789,N_3640);
nor U6616 (N_6616,N_2566,N_231);
or U6617 (N_6617,N_4705,N_1248);
nor U6618 (N_6618,N_351,N_1644);
and U6619 (N_6619,N_1457,N_2452);
and U6620 (N_6620,N_3648,N_3148);
nor U6621 (N_6621,N_2107,N_212);
nor U6622 (N_6622,N_2790,N_2337);
and U6623 (N_6623,N_1278,N_765);
xor U6624 (N_6624,N_1536,N_2175);
nand U6625 (N_6625,N_2748,N_3374);
nand U6626 (N_6626,N_4581,N_2248);
nand U6627 (N_6627,N_3704,N_609);
nand U6628 (N_6628,N_2038,N_3244);
or U6629 (N_6629,N_2851,N_4774);
xnor U6630 (N_6630,N_4207,N_3774);
nor U6631 (N_6631,N_3379,N_2051);
nor U6632 (N_6632,N_1621,N_2964);
xnor U6633 (N_6633,N_4519,N_3012);
nand U6634 (N_6634,N_2262,N_4731);
or U6635 (N_6635,N_4907,N_3649);
or U6636 (N_6636,N_827,N_3547);
and U6637 (N_6637,N_3345,N_4026);
nand U6638 (N_6638,N_3560,N_1671);
and U6639 (N_6639,N_3619,N_2733);
xor U6640 (N_6640,N_1306,N_4157);
or U6641 (N_6641,N_1125,N_2172);
and U6642 (N_6642,N_4492,N_2341);
xor U6643 (N_6643,N_2324,N_3261);
and U6644 (N_6644,N_1351,N_4908);
or U6645 (N_6645,N_1500,N_2004);
or U6646 (N_6646,N_115,N_1519);
or U6647 (N_6647,N_4684,N_3586);
or U6648 (N_6648,N_1336,N_4455);
or U6649 (N_6649,N_2523,N_3325);
and U6650 (N_6650,N_3639,N_2728);
nor U6651 (N_6651,N_3304,N_2127);
nand U6652 (N_6652,N_2718,N_2005);
or U6653 (N_6653,N_2702,N_1691);
or U6654 (N_6654,N_4121,N_3725);
nor U6655 (N_6655,N_2007,N_3804);
or U6656 (N_6656,N_1945,N_4275);
and U6657 (N_6657,N_1501,N_809);
and U6658 (N_6658,N_1978,N_3613);
xnor U6659 (N_6659,N_686,N_4916);
and U6660 (N_6660,N_2796,N_1642);
and U6661 (N_6661,N_4962,N_1205);
nand U6662 (N_6662,N_4091,N_3128);
and U6663 (N_6663,N_4859,N_2424);
or U6664 (N_6664,N_4886,N_718);
and U6665 (N_6665,N_4395,N_3396);
and U6666 (N_6666,N_4702,N_302);
nor U6667 (N_6667,N_883,N_3904);
nand U6668 (N_6668,N_2922,N_4362);
xor U6669 (N_6669,N_4541,N_2163);
nor U6670 (N_6670,N_1570,N_2084);
nand U6671 (N_6671,N_2406,N_3693);
and U6672 (N_6672,N_2563,N_1064);
xnor U6673 (N_6673,N_4669,N_3125);
nor U6674 (N_6674,N_3000,N_4783);
or U6675 (N_6675,N_3581,N_2833);
xnor U6676 (N_6676,N_4088,N_3953);
and U6677 (N_6677,N_1055,N_3162);
and U6678 (N_6678,N_1900,N_136);
or U6679 (N_6679,N_897,N_764);
and U6680 (N_6680,N_272,N_4836);
or U6681 (N_6681,N_4167,N_1729);
xor U6682 (N_6682,N_1651,N_3143);
or U6683 (N_6683,N_3454,N_940);
and U6684 (N_6684,N_1441,N_8);
nor U6685 (N_6685,N_3350,N_2629);
nand U6686 (N_6686,N_1509,N_814);
nor U6687 (N_6687,N_1947,N_874);
xor U6688 (N_6688,N_1999,N_1266);
or U6689 (N_6689,N_3859,N_2462);
or U6690 (N_6690,N_4086,N_651);
and U6691 (N_6691,N_4636,N_3478);
and U6692 (N_6692,N_3470,N_4704);
or U6693 (N_6693,N_1532,N_3196);
nand U6694 (N_6694,N_1368,N_1940);
xor U6695 (N_6695,N_2554,N_3917);
and U6696 (N_6696,N_2999,N_2142);
or U6697 (N_6697,N_908,N_1918);
or U6698 (N_6698,N_278,N_3902);
and U6699 (N_6699,N_1379,N_3891);
nand U6700 (N_6700,N_2534,N_3509);
or U6701 (N_6701,N_574,N_250);
nand U6702 (N_6702,N_3573,N_1422);
or U6703 (N_6703,N_4402,N_2011);
or U6704 (N_6704,N_3958,N_1461);
nor U6705 (N_6705,N_4728,N_2682);
nand U6706 (N_6706,N_656,N_1124);
nor U6707 (N_6707,N_872,N_1639);
nor U6708 (N_6708,N_4981,N_1600);
and U6709 (N_6709,N_1922,N_3906);
nand U6710 (N_6710,N_2165,N_355);
nor U6711 (N_6711,N_2529,N_944);
and U6712 (N_6712,N_3705,N_286);
nand U6713 (N_6713,N_1113,N_1130);
or U6714 (N_6714,N_1389,N_4779);
nor U6715 (N_6715,N_1539,N_4566);
nor U6716 (N_6716,N_3319,N_994);
nand U6717 (N_6717,N_1955,N_1307);
nor U6718 (N_6718,N_2943,N_28);
nor U6719 (N_6719,N_979,N_2180);
and U6720 (N_6720,N_2252,N_2996);
xor U6721 (N_6721,N_786,N_2564);
nor U6722 (N_6722,N_120,N_2147);
nor U6723 (N_6723,N_51,N_2950);
nand U6724 (N_6724,N_4215,N_2724);
nand U6725 (N_6725,N_3616,N_951);
and U6726 (N_6726,N_1738,N_1325);
nand U6727 (N_6727,N_1240,N_1462);
xor U6728 (N_6728,N_1200,N_3315);
and U6729 (N_6729,N_2753,N_3464);
nand U6730 (N_6730,N_4972,N_1021);
nand U6731 (N_6731,N_2490,N_2864);
nor U6732 (N_6732,N_2861,N_316);
nor U6733 (N_6733,N_2882,N_716);
nor U6734 (N_6734,N_3749,N_368);
and U6735 (N_6735,N_127,N_3278);
or U6736 (N_6736,N_442,N_1394);
xnor U6737 (N_6737,N_2458,N_2829);
and U6738 (N_6738,N_322,N_388);
nand U6739 (N_6739,N_1657,N_2780);
and U6740 (N_6740,N_3392,N_4084);
or U6741 (N_6741,N_3543,N_3206);
or U6742 (N_6742,N_1046,N_4893);
or U6743 (N_6743,N_1155,N_4105);
xnor U6744 (N_6744,N_303,N_144);
or U6745 (N_6745,N_2975,N_1969);
nand U6746 (N_6746,N_1735,N_4739);
or U6747 (N_6747,N_403,N_3814);
nand U6748 (N_6748,N_504,N_2698);
nand U6749 (N_6749,N_1861,N_2640);
nand U6750 (N_6750,N_151,N_1487);
nand U6751 (N_6751,N_275,N_4738);
and U6752 (N_6752,N_1311,N_4587);
nand U6753 (N_6753,N_1655,N_4594);
and U6754 (N_6754,N_1964,N_3197);
nand U6755 (N_6755,N_1164,N_3712);
and U6756 (N_6756,N_2679,N_1426);
nor U6757 (N_6757,N_4394,N_2336);
xor U6758 (N_6758,N_2900,N_1276);
nor U6759 (N_6759,N_1698,N_1518);
nor U6760 (N_6760,N_3821,N_1863);
or U6761 (N_6761,N_126,N_3262);
or U6762 (N_6762,N_3341,N_237);
nor U6763 (N_6763,N_3314,N_4325);
and U6764 (N_6764,N_3399,N_3220);
or U6765 (N_6765,N_3896,N_3023);
or U6766 (N_6766,N_923,N_1060);
and U6767 (N_6767,N_2955,N_1562);
and U6768 (N_6768,N_2558,N_1624);
nor U6769 (N_6769,N_1275,N_1083);
nor U6770 (N_6770,N_2047,N_1062);
nor U6771 (N_6771,N_578,N_2580);
or U6772 (N_6772,N_3819,N_790);
or U6773 (N_6773,N_2914,N_4482);
xnor U6774 (N_6774,N_1298,N_678);
nand U6775 (N_6775,N_2694,N_2361);
nand U6776 (N_6776,N_3285,N_374);
or U6777 (N_6777,N_80,N_159);
nor U6778 (N_6778,N_397,N_257);
or U6779 (N_6779,N_1418,N_101);
nand U6780 (N_6780,N_1766,N_1693);
or U6781 (N_6781,N_1260,N_4583);
or U6782 (N_6782,N_3060,N_1189);
or U6783 (N_6783,N_1268,N_4256);
nand U6784 (N_6784,N_1072,N_3654);
nand U6785 (N_6785,N_3948,N_1754);
and U6786 (N_6786,N_613,N_4876);
nand U6787 (N_6787,N_1143,N_3419);
and U6788 (N_6788,N_1879,N_2487);
or U6789 (N_6789,N_2039,N_1910);
xnor U6790 (N_6790,N_3684,N_288);
or U6791 (N_6791,N_835,N_454);
nand U6792 (N_6792,N_698,N_2159);
nand U6793 (N_6793,N_3301,N_48);
nand U6794 (N_6794,N_3516,N_4741);
and U6795 (N_6795,N_530,N_4237);
or U6796 (N_6796,N_1638,N_1075);
and U6797 (N_6797,N_3134,N_3574);
or U6798 (N_6798,N_318,N_4591);
nor U6799 (N_6799,N_3034,N_2195);
nor U6800 (N_6800,N_4850,N_798);
nand U6801 (N_6801,N_2019,N_4477);
or U6802 (N_6802,N_625,N_3857);
nor U6803 (N_6803,N_1451,N_4441);
and U6804 (N_6804,N_4365,N_1316);
nor U6805 (N_6805,N_134,N_4289);
nor U6806 (N_6806,N_3775,N_2616);
nand U6807 (N_6807,N_3092,N_1091);
or U6808 (N_6808,N_3636,N_4644);
and U6809 (N_6809,N_1530,N_4641);
nand U6810 (N_6810,N_2338,N_2784);
or U6811 (N_6811,N_1820,N_2552);
nor U6812 (N_6812,N_4023,N_869);
and U6813 (N_6813,N_2878,N_1603);
or U6814 (N_6814,N_2105,N_472);
nor U6815 (N_6815,N_3295,N_460);
or U6816 (N_6816,N_4956,N_22);
and U6817 (N_6817,N_2945,N_1798);
or U6818 (N_6818,N_148,N_279);
nor U6819 (N_6819,N_3263,N_196);
nand U6820 (N_6820,N_4046,N_4148);
nand U6821 (N_6821,N_2405,N_206);
nand U6822 (N_6822,N_4861,N_771);
nor U6823 (N_6823,N_2284,N_4894);
nand U6824 (N_6824,N_4331,N_4857);
nand U6825 (N_6825,N_2148,N_1756);
nand U6826 (N_6826,N_2986,N_1347);
or U6827 (N_6827,N_3239,N_1676);
xor U6828 (N_6828,N_4078,N_4252);
xnor U6829 (N_6829,N_2961,N_1285);
nand U6830 (N_6830,N_2553,N_4130);
nor U6831 (N_6831,N_980,N_1224);
or U6832 (N_6832,N_1112,N_1435);
and U6833 (N_6833,N_2895,N_4905);
nand U6834 (N_6834,N_2638,N_2600);
or U6835 (N_6835,N_1834,N_3810);
nand U6836 (N_6836,N_1723,N_3264);
nand U6837 (N_6837,N_4214,N_4733);
xor U6838 (N_6838,N_1835,N_1425);
nand U6839 (N_6839,N_3448,N_3537);
and U6840 (N_6840,N_2012,N_3110);
nor U6841 (N_6841,N_1467,N_4382);
nand U6842 (N_6842,N_1566,N_501);
xor U6843 (N_6843,N_1768,N_2511);
and U6844 (N_6844,N_3040,N_1629);
or U6845 (N_6845,N_1460,N_3024);
nand U6846 (N_6846,N_1589,N_2666);
and U6847 (N_6847,N_2446,N_19);
and U6848 (N_6848,N_2471,N_1849);
nor U6849 (N_6849,N_3256,N_2887);
and U6850 (N_6850,N_3685,N_4320);
and U6851 (N_6851,N_2842,N_133);
and U6852 (N_6852,N_360,N_1789);
nand U6853 (N_6853,N_3500,N_824);
or U6854 (N_6854,N_77,N_1894);
nand U6855 (N_6855,N_2550,N_2978);
and U6856 (N_6856,N_1660,N_3447);
xnor U6857 (N_6857,N_4721,N_4031);
nor U6858 (N_6858,N_2339,N_3691);
or U6859 (N_6859,N_2936,N_4189);
and U6860 (N_6860,N_2281,N_1758);
nor U6861 (N_6861,N_4374,N_1814);
xnor U6862 (N_6862,N_3421,N_2551);
nor U6863 (N_6863,N_3842,N_3837);
nor U6864 (N_6864,N_3324,N_2483);
nand U6865 (N_6865,N_4573,N_1051);
nand U6866 (N_6866,N_3565,N_1330);
nor U6867 (N_6867,N_2099,N_15);
xor U6868 (N_6868,N_2243,N_3877);
and U6869 (N_6869,N_2158,N_4123);
or U6870 (N_6870,N_465,N_4447);
nor U6871 (N_6871,N_1876,N_669);
nor U6872 (N_6872,N_156,N_2625);
nor U6873 (N_6873,N_3343,N_2491);
xnor U6874 (N_6874,N_4075,N_52);
nor U6875 (N_6875,N_3974,N_4489);
and U6876 (N_6876,N_3736,N_4095);
nor U6877 (N_6877,N_593,N_4937);
or U6878 (N_6878,N_2746,N_2846);
nand U6879 (N_6879,N_2106,N_3201);
nor U6880 (N_6880,N_4504,N_1892);
and U6881 (N_6881,N_4173,N_3245);
or U6882 (N_6882,N_344,N_4660);
and U6883 (N_6883,N_3922,N_3472);
and U6884 (N_6884,N_456,N_187);
and U6885 (N_6885,N_3019,N_3042);
nor U6886 (N_6886,N_1037,N_4844);
and U6887 (N_6887,N_2865,N_680);
nor U6888 (N_6888,N_635,N_104);
or U6889 (N_6889,N_241,N_4094);
and U6890 (N_6890,N_1029,N_1488);
xor U6891 (N_6891,N_4712,N_3248);
nor U6892 (N_6892,N_2402,N_1667);
or U6893 (N_6893,N_2304,N_3476);
xnor U6894 (N_6894,N_4092,N_2208);
nand U6895 (N_6895,N_2333,N_4632);
nand U6896 (N_6896,N_557,N_3116);
nor U6897 (N_6897,N_1592,N_4674);
nor U6898 (N_6898,N_2813,N_3801);
nand U6899 (N_6899,N_2763,N_3530);
nand U6900 (N_6900,N_3364,N_3053);
nor U6901 (N_6901,N_3103,N_4963);
and U6902 (N_6902,N_100,N_3607);
and U6903 (N_6903,N_2407,N_2052);
or U6904 (N_6904,N_2412,N_4539);
nand U6905 (N_6905,N_1273,N_775);
nor U6906 (N_6906,N_850,N_4603);
nor U6907 (N_6907,N_2089,N_2634);
and U6908 (N_6908,N_3730,N_1577);
xor U6909 (N_6909,N_2917,N_1219);
or U6910 (N_6910,N_3457,N_4752);
xor U6911 (N_6911,N_171,N_481);
or U6912 (N_6912,N_1931,N_4543);
and U6913 (N_6913,N_1069,N_4041);
nand U6914 (N_6914,N_338,N_832);
nor U6915 (N_6915,N_2319,N_522);
nor U6916 (N_6916,N_4104,N_4442);
nor U6917 (N_6917,N_1162,N_1930);
or U6918 (N_6918,N_4713,N_1088);
and U6919 (N_6919,N_1700,N_1481);
nand U6920 (N_6920,N_611,N_518);
or U6921 (N_6921,N_604,N_2731);
or U6922 (N_6922,N_3540,N_242);
or U6923 (N_6923,N_4280,N_4009);
and U6924 (N_6924,N_3265,N_1694);
nor U6925 (N_6925,N_3596,N_1221);
nand U6926 (N_6926,N_4120,N_1246);
nor U6927 (N_6927,N_3621,N_2181);
nor U6928 (N_6928,N_2688,N_140);
or U6929 (N_6929,N_4655,N_2376);
nand U6930 (N_6930,N_1831,N_4436);
and U6931 (N_6931,N_114,N_110);
nand U6932 (N_6932,N_1348,N_1027);
and U6933 (N_6933,N_4405,N_733);
or U6934 (N_6934,N_1172,N_3966);
nand U6935 (N_6935,N_4429,N_219);
nor U6936 (N_6936,N_3430,N_27);
nand U6937 (N_6937,N_1793,N_4210);
and U6938 (N_6938,N_2560,N_4283);
or U6939 (N_6939,N_1925,N_1404);
nand U6940 (N_6940,N_2354,N_4339);
or U6941 (N_6941,N_2166,N_2546);
nand U6942 (N_6942,N_2267,N_558);
or U6943 (N_6943,N_2565,N_1913);
xor U6944 (N_6944,N_691,N_3453);
nor U6945 (N_6945,N_2141,N_4133);
nor U6946 (N_6946,N_1630,N_4559);
nor U6947 (N_6947,N_745,N_297);
nor U6948 (N_6948,N_4222,N_4175);
nand U6949 (N_6949,N_3097,N_1050);
nand U6950 (N_6950,N_3608,N_4128);
nor U6951 (N_6951,N_671,N_3077);
nand U6952 (N_6952,N_415,N_4438);
xor U6953 (N_6953,N_438,N_4509);
nand U6954 (N_6954,N_152,N_3258);
nand U6955 (N_6955,N_1914,N_2848);
nor U6956 (N_6956,N_3275,N_3202);
nand U6957 (N_6957,N_3866,N_2852);
nand U6958 (N_6958,N_2326,N_1650);
nor U6959 (N_6959,N_3031,N_1810);
nand U6960 (N_6960,N_3170,N_2485);
nand U6961 (N_6961,N_1531,N_2545);
or U6962 (N_6962,N_1840,N_1190);
nand U6963 (N_6963,N_3951,N_1741);
nor U6964 (N_6964,N_3768,N_1333);
xnor U6965 (N_6965,N_2824,N_1675);
nand U6966 (N_6966,N_26,N_4564);
xor U6967 (N_6967,N_4640,N_4180);
and U6968 (N_6968,N_2615,N_2140);
and U6969 (N_6969,N_2370,N_462);
nand U6970 (N_6970,N_3696,N_4453);
nand U6971 (N_6971,N_1158,N_2342);
and U6972 (N_6972,N_90,N_740);
nand U6973 (N_6973,N_3171,N_157);
or U6974 (N_6974,N_1144,N_1580);
nor U6975 (N_6975,N_3194,N_2110);
nor U6976 (N_6976,N_4606,N_4793);
xnor U6977 (N_6977,N_3291,N_3921);
and U6978 (N_6978,N_4801,N_4707);
or U6979 (N_6979,N_1537,N_3706);
nor U6980 (N_6980,N_4947,N_2028);
and U6981 (N_6981,N_1890,N_97);
or U6982 (N_6982,N_1490,N_3862);
and U6983 (N_6983,N_4353,N_4064);
and U6984 (N_6984,N_1517,N_3013);
and U6985 (N_6985,N_4290,N_1962);
nor U6986 (N_6986,N_499,N_2876);
and U6987 (N_6987,N_3415,N_4315);
and U6988 (N_6988,N_4486,N_3965);
and U6989 (N_6989,N_193,N_3961);
nor U6990 (N_6990,N_1170,N_1617);
and U6991 (N_6991,N_1236,N_805);
xnor U6992 (N_6992,N_3049,N_3585);
nor U6993 (N_6993,N_1895,N_1047);
nor U6994 (N_6994,N_3726,N_1319);
nor U6995 (N_6995,N_4203,N_614);
and U6996 (N_6996,N_928,N_1139);
and U6997 (N_6997,N_3359,N_1106);
nand U6998 (N_6998,N_4761,N_543);
nor U6999 (N_6999,N_4921,N_4250);
and U7000 (N_7000,N_411,N_314);
nor U7001 (N_7001,N_1937,N_1984);
nor U7002 (N_7002,N_2055,N_4328);
and U7003 (N_7003,N_2365,N_1232);
xnor U7004 (N_7004,N_1929,N_952);
and U7005 (N_7005,N_4758,N_4692);
nor U7006 (N_7006,N_2049,N_189);
xor U7007 (N_7007,N_2501,N_135);
and U7008 (N_7008,N_4515,N_4646);
nand U7009 (N_7009,N_4979,N_3848);
or U7010 (N_7010,N_4024,N_4569);
and U7011 (N_7011,N_584,N_298);
nor U7012 (N_7012,N_1407,N_3260);
and U7013 (N_7013,N_384,N_315);
and U7014 (N_7014,N_2543,N_1858);
or U7015 (N_7015,N_3549,N_1087);
and U7016 (N_7016,N_500,N_2677);
xnor U7017 (N_7017,N_4115,N_1053);
or U7018 (N_7018,N_1842,N_4279);
or U7019 (N_7019,N_1779,N_3172);
nand U7020 (N_7020,N_1093,N_2167);
xnor U7021 (N_7021,N_1972,N_840);
and U7022 (N_7022,N_424,N_647);
and U7023 (N_7023,N_865,N_1341);
or U7024 (N_7024,N_469,N_1356);
or U7025 (N_7025,N_639,N_1241);
or U7026 (N_7026,N_2212,N_3729);
nor U7027 (N_7027,N_1674,N_1035);
or U7028 (N_7028,N_4193,N_69);
nor U7029 (N_7029,N_346,N_2902);
nor U7030 (N_7030,N_2827,N_2716);
nor U7031 (N_7031,N_677,N_238);
and U7032 (N_7032,N_2737,N_331);
nand U7033 (N_7033,N_3796,N_917);
nor U7034 (N_7034,N_1514,N_1334);
xor U7035 (N_7035,N_1052,N_494);
nor U7036 (N_7036,N_3662,N_2556);
nand U7037 (N_7037,N_4221,N_984);
nand U7038 (N_7038,N_1257,N_886);
or U7039 (N_7039,N_1065,N_258);
and U7040 (N_7040,N_1701,N_2875);
or U7041 (N_7041,N_4939,N_3393);
or U7042 (N_7042,N_3611,N_2389);
or U7043 (N_7043,N_4197,N_3890);
or U7044 (N_7044,N_1601,N_4181);
or U7045 (N_7045,N_3676,N_4196);
nand U7046 (N_7046,N_4627,N_1707);
nor U7047 (N_7047,N_1583,N_1344);
or U7048 (N_7048,N_1391,N_377);
or U7049 (N_7049,N_2027,N_234);
nor U7050 (N_7050,N_2838,N_1175);
nor U7051 (N_7051,N_3513,N_2293);
nor U7052 (N_7052,N_3433,N_3288);
nor U7053 (N_7053,N_2464,N_448);
or U7054 (N_7054,N_2368,N_183);
and U7055 (N_7055,N_3724,N_1364);
nor U7056 (N_7056,N_116,N_965);
nor U7057 (N_7057,N_4885,N_3076);
nand U7058 (N_7058,N_4304,N_1935);
or U7059 (N_7059,N_4788,N_675);
nand U7060 (N_7060,N_1804,N_1503);
or U7061 (N_7061,N_130,N_3378);
or U7062 (N_7062,N_1485,N_937);
nand U7063 (N_7063,N_4948,N_3555);
and U7064 (N_7064,N_378,N_2492);
nor U7065 (N_7065,N_1001,N_290);
and U7066 (N_7066,N_4510,N_3035);
and U7067 (N_7067,N_3823,N_4352);
nor U7068 (N_7068,N_3554,N_615);
or U7069 (N_7069,N_2987,N_2315);
nand U7070 (N_7070,N_1283,N_3163);
or U7071 (N_7071,N_505,N_2855);
or U7072 (N_7072,N_985,N_5);
nand U7073 (N_7073,N_1483,N_2944);
nand U7074 (N_7074,N_1608,N_2205);
nand U7075 (N_7075,N_417,N_407);
and U7076 (N_7076,N_1649,N_14);
nor U7077 (N_7077,N_4755,N_758);
nand U7078 (N_7078,N_2877,N_1008);
and U7079 (N_7079,N_561,N_2280);
and U7080 (N_7080,N_4789,N_4242);
nor U7081 (N_7081,N_1141,N_2321);
xor U7082 (N_7082,N_977,N_4191);
nand U7083 (N_7083,N_4432,N_3615);
and U7084 (N_7084,N_2044,N_3153);
and U7085 (N_7085,N_434,N_3121);
nand U7086 (N_7086,N_2854,N_4622);
nor U7087 (N_7087,N_2244,N_701);
xor U7088 (N_7088,N_3645,N_4035);
nand U7089 (N_7089,N_3722,N_3967);
or U7090 (N_7090,N_3179,N_3006);
and U7091 (N_7091,N_4668,N_1546);
nor U7092 (N_7092,N_1085,N_4015);
nand U7093 (N_7093,N_2410,N_1100);
xnor U7094 (N_7094,N_4338,N_4428);
nand U7095 (N_7095,N_141,N_358);
nor U7096 (N_7096,N_3969,N_1405);
or U7097 (N_7097,N_553,N_4318);
or U7098 (N_7098,N_4691,N_2223);
and U7099 (N_7099,N_150,N_967);
or U7100 (N_7100,N_2079,N_3407);
and U7101 (N_7101,N_702,N_599);
or U7102 (N_7102,N_328,N_4302);
and U7103 (N_7103,N_1510,N_2130);
nor U7104 (N_7104,N_1783,N_642);
nand U7105 (N_7105,N_2923,N_4561);
nor U7106 (N_7106,N_71,N_1658);
nand U7107 (N_7107,N_3599,N_3800);
xnor U7108 (N_7108,N_1386,N_3332);
nand U7109 (N_7109,N_4012,N_4389);
and U7110 (N_7110,N_617,N_2913);
nand U7111 (N_7111,N_2064,N_4149);
nand U7112 (N_7112,N_2057,N_1740);
nor U7113 (N_7113,N_3048,N_1217);
nand U7114 (N_7114,N_3672,N_4271);
xnor U7115 (N_7115,N_2498,N_2271);
nor U7116 (N_7116,N_455,N_2117);
nor U7117 (N_7117,N_705,N_1041);
nand U7118 (N_7118,N_2168,N_4223);
or U7119 (N_7119,N_1718,N_2179);
or U7120 (N_7120,N_205,N_1174);
nor U7121 (N_7121,N_3087,N_806);
and U7122 (N_7122,N_337,N_4476);
and U7123 (N_7123,N_2805,N_4961);
or U7124 (N_7124,N_4297,N_2216);
nand U7125 (N_7125,N_321,N_2555);
and U7126 (N_7126,N_1761,N_3099);
or U7127 (N_7127,N_3874,N_2366);
nand U7128 (N_7128,N_3900,N_2129);
nor U7129 (N_7129,N_540,N_527);
nand U7130 (N_7130,N_1772,N_714);
or U7131 (N_7131,N_4871,N_1829);
nand U7132 (N_7132,N_638,N_2474);
or U7133 (N_7133,N_2646,N_2578);
or U7134 (N_7134,N_2603,N_2835);
nor U7135 (N_7135,N_3145,N_1932);
nand U7136 (N_7136,N_4156,N_1640);
nor U7137 (N_7137,N_2845,N_3269);
or U7138 (N_7138,N_3322,N_483);
nand U7139 (N_7139,N_3959,N_1354);
or U7140 (N_7140,N_4881,N_2488);
nand U7141 (N_7141,N_4017,N_3489);
and U7142 (N_7142,N_4790,N_3390);
and U7143 (N_7143,N_1433,N_2232);
or U7144 (N_7144,N_1886,N_1865);
and U7145 (N_7145,N_3353,N_4243);
and U7146 (N_7146,N_2856,N_177);
nand U7147 (N_7147,N_4502,N_2959);
and U7148 (N_7148,N_2888,N_4487);
nor U7149 (N_7149,N_3737,N_4392);
nor U7150 (N_7150,N_4653,N_3502);
nor U7151 (N_7151,N_2652,N_1186);
and U7152 (N_7152,N_4178,N_1717);
and U7153 (N_7153,N_1817,N_1881);
nand U7154 (N_7154,N_2635,N_4703);
or U7155 (N_7155,N_3598,N_2206);
nor U7156 (N_7156,N_4053,N_2661);
xnor U7157 (N_7157,N_3666,N_373);
nor U7158 (N_7158,N_1816,N_2221);
and U7159 (N_7159,N_3673,N_773);
or U7160 (N_7160,N_3512,N_111);
and U7161 (N_7161,N_1070,N_1245);
xnor U7162 (N_7162,N_2300,N_326);
nand U7163 (N_7163,N_2274,N_4633);
or U7164 (N_7164,N_225,N_3009);
nor U7165 (N_7165,N_4895,N_4348);
nand U7166 (N_7166,N_2912,N_324);
nand U7167 (N_7167,N_1827,N_4042);
nand U7168 (N_7168,N_2571,N_2832);
and U7169 (N_7169,N_571,N_3701);
nand U7170 (N_7170,N_2434,N_3021);
or U7171 (N_7171,N_896,N_83);
or U7172 (N_7172,N_4864,N_2382);
nor U7173 (N_7173,N_607,N_2399);
or U7174 (N_7174,N_1152,N_4745);
or U7175 (N_7175,N_1444,N_4022);
and U7176 (N_7176,N_4044,N_2976);
xor U7177 (N_7177,N_3789,N_4647);
nor U7178 (N_7178,N_3850,N_482);
nand U7179 (N_7179,N_3425,N_1543);
xnor U7180 (N_7180,N_715,N_1159);
or U7181 (N_7181,N_3337,N_2983);
and U7182 (N_7182,N_3822,N_400);
nand U7183 (N_7183,N_4860,N_1020);
and U7184 (N_7184,N_3984,N_2440);
or U7185 (N_7185,N_4786,N_4681);
nor U7186 (N_7186,N_3838,N_946);
or U7187 (N_7187,N_3888,N_2085);
and U7188 (N_7188,N_4462,N_489);
nand U7189 (N_7189,N_3829,N_1473);
or U7190 (N_7190,N_3700,N_3597);
or U7191 (N_7191,N_2830,N_3137);
xnor U7192 (N_7192,N_3872,N_4781);
and U7193 (N_7193,N_2908,N_4333);
or U7194 (N_7194,N_3609,N_4317);
or U7195 (N_7195,N_586,N_4341);
nor U7196 (N_7196,N_4109,N_1686);
and U7197 (N_7197,N_2213,N_4666);
nand U7198 (N_7198,N_1380,N_782);
or U7199 (N_7199,N_2240,N_1612);
nand U7200 (N_7200,N_794,N_4494);
and U7201 (N_7201,N_4480,N_4326);
nor U7202 (N_7202,N_4798,N_2088);
nor U7203 (N_7203,N_4676,N_4116);
nand U7204 (N_7204,N_3149,N_421);
and U7205 (N_7205,N_2119,N_1128);
xor U7206 (N_7206,N_1090,N_3387);
nor U7207 (N_7207,N_4592,N_4021);
or U7208 (N_7208,N_706,N_4579);
nand U7209 (N_7209,N_1226,N_3372);
and U7210 (N_7210,N_1508,N_3289);
xor U7211 (N_7211,N_3915,N_4914);
nand U7212 (N_7212,N_4446,N_341);
or U7213 (N_7213,N_1695,N_4373);
and U7214 (N_7214,N_1249,N_1471);
xor U7215 (N_7215,N_1778,N_2989);
nor U7216 (N_7216,N_899,N_3978);
nand U7217 (N_7217,N_4337,N_2988);
nor U7218 (N_7218,N_4344,N_2658);
or U7219 (N_7219,N_2144,N_4595);
nor U7220 (N_7220,N_1373,N_4407);
and U7221 (N_7221,N_2058,N_2303);
nand U7222 (N_7222,N_1632,N_891);
nand U7223 (N_7223,N_4809,N_2314);
and U7224 (N_7224,N_1821,N_2602);
and U7225 (N_7225,N_2797,N_3215);
or U7226 (N_7226,N_3079,N_2585);
nand U7227 (N_7227,N_3398,N_520);
or U7228 (N_7228,N_2905,N_4019);
and U7229 (N_7229,N_4709,N_4284);
or U7230 (N_7230,N_657,N_3668);
xnor U7231 (N_7231,N_4516,N_4795);
nor U7232 (N_7232,N_64,N_3427);
or U7233 (N_7233,N_3452,N_2094);
nor U7234 (N_7234,N_1321,N_2982);
nor U7235 (N_7235,N_3155,N_2871);
or U7236 (N_7236,N_4938,N_2714);
or U7237 (N_7237,N_4835,N_1811);
nor U7238 (N_7238,N_1973,N_3101);
nand U7239 (N_7239,N_2048,N_1166);
nor U7240 (N_7240,N_1719,N_4949);
or U7241 (N_7241,N_2974,N_3772);
nand U7242 (N_7242,N_957,N_4396);
or U7243 (N_7243,N_3733,N_340);
nor U7244 (N_7244,N_1777,N_113);
or U7245 (N_7245,N_3758,N_2444);
and U7246 (N_7246,N_41,N_2828);
and U7247 (N_7247,N_2814,N_4912);
nand U7248 (N_7248,N_4722,N_67);
nand U7249 (N_7249,N_390,N_4699);
and U7250 (N_7250,N_1179,N_3683);
nand U7251 (N_7251,N_3920,N_2628);
nand U7252 (N_7252,N_4445,N_699);
or U7253 (N_7253,N_4528,N_2018);
nor U7254 (N_7254,N_4198,N_1446);
or U7255 (N_7255,N_3080,N_3274);
nor U7256 (N_7256,N_4848,N_4003);
or U7257 (N_7257,N_529,N_2656);
nor U7258 (N_7258,N_623,N_3563);
or U7259 (N_7259,N_1968,N_3083);
or U7260 (N_7260,N_536,N_3606);
nor U7261 (N_7261,N_2831,N_2449);
nand U7262 (N_7262,N_1015,N_3545);
nand U7263 (N_7263,N_1525,N_3340);
nor U7264 (N_7264,N_305,N_56);
xnor U7265 (N_7265,N_3898,N_3126);
and U7266 (N_7266,N_1548,N_3294);
nand U7267 (N_7267,N_4984,N_922);
nor U7268 (N_7268,N_399,N_523);
or U7269 (N_7269,N_2683,N_598);
and U7270 (N_7270,N_3686,N_2881);
nand U7271 (N_7271,N_4996,N_3594);
and U7272 (N_7272,N_2317,N_3271);
or U7273 (N_7273,N_3067,N_2330);
xor U7274 (N_7274,N_4900,N_105);
nor U7275 (N_7275,N_4213,N_2062);
nand U7276 (N_7276,N_4209,N_119);
or U7277 (N_7277,N_1092,N_4663);
and U7278 (N_7278,N_4824,N_3309);
or U7279 (N_7279,N_4960,N_2951);
or U7280 (N_7280,N_2422,N_3186);
and U7281 (N_7281,N_178,N_4287);
nand U7282 (N_7282,N_3479,N_4608);
nand U7283 (N_7283,N_1555,N_3794);
and U7284 (N_7284,N_3806,N_2535);
xnor U7285 (N_7285,N_1194,N_1635);
or U7286 (N_7286,N_978,N_2547);
nor U7287 (N_7287,N_2146,N_2421);
or U7288 (N_7288,N_933,N_1862);
xnor U7289 (N_7289,N_1419,N_1208);
or U7290 (N_7290,N_3458,N_352);
or U7291 (N_7291,N_1664,N_1438);
nor U7292 (N_7292,N_2958,N_3328);
nor U7293 (N_7293,N_779,N_3473);
nor U7294 (N_7294,N_1381,N_2292);
or U7295 (N_7295,N_743,N_2607);
or U7296 (N_7296,N_17,N_4080);
nor U7297 (N_7297,N_3753,N_2924);
nor U7298 (N_7298,N_4990,N_161);
nor U7299 (N_7299,N_1690,N_146);
and U7300 (N_7300,N_4557,N_514);
nand U7301 (N_7301,N_1388,N_3503);
nand U7302 (N_7302,N_3159,N_3546);
nor U7303 (N_7303,N_1920,N_4944);
nand U7304 (N_7304,N_3870,N_2083);
and U7305 (N_7305,N_3946,N_4097);
nor U7306 (N_7306,N_1286,N_1066);
nand U7307 (N_7307,N_959,N_367);
and U7308 (N_7308,N_406,N_1899);
nor U7309 (N_7309,N_3930,N_4851);
nor U7310 (N_7310,N_496,N_2260);
xnor U7311 (N_7311,N_2371,N_4855);
or U7312 (N_7312,N_3595,N_4817);
nand U7313 (N_7313,N_3032,N_3760);
xor U7314 (N_7314,N_2484,N_517);
and U7315 (N_7315,N_1808,N_901);
nor U7316 (N_7316,N_1358,N_542);
nand U7317 (N_7317,N_1952,N_2108);
nor U7318 (N_7318,N_3727,N_313);
xnor U7319 (N_7319,N_4174,N_1666);
nor U7320 (N_7320,N_239,N_1133);
or U7321 (N_7321,N_1569,N_4499);
nor U7322 (N_7322,N_1743,N_1474);
nand U7323 (N_7323,N_4460,N_4060);
nand U7324 (N_7324,N_176,N_880);
and U7325 (N_7325,N_914,N_1339);
xnor U7326 (N_7326,N_2273,N_4726);
nor U7327 (N_7327,N_1207,N_3062);
nand U7328 (N_7328,N_3788,N_546);
or U7329 (N_7329,N_3720,N_1324);
and U7330 (N_7330,N_464,N_3234);
nor U7331 (N_7331,N_682,N_1867);
or U7332 (N_7332,N_4768,N_2726);
or U7333 (N_7333,N_3849,N_3620);
xor U7334 (N_7334,N_2942,N_4332);
nor U7335 (N_7335,N_4838,N_4232);
nand U7336 (N_7336,N_1534,N_2041);
nand U7337 (N_7337,N_4030,N_2463);
nand U7338 (N_7338,N_4957,N_2970);
and U7339 (N_7339,N_4057,N_581);
nor U7340 (N_7340,N_197,N_4391);
or U7341 (N_7341,N_4051,N_2972);
nand U7342 (N_7342,N_531,N_2279);
or U7343 (N_7343,N_4505,N_1942);
and U7344 (N_7344,N_1352,N_2930);
xnor U7345 (N_7345,N_3735,N_2548);
and U7346 (N_7346,N_3661,N_2695);
and U7347 (N_7347,N_1917,N_544);
and U7348 (N_7348,N_266,N_45);
nor U7349 (N_7349,N_3005,N_509);
nor U7350 (N_7350,N_4410,N_1663);
xnor U7351 (N_7351,N_2907,N_2569);
nor U7352 (N_7352,N_2921,N_131);
and U7353 (N_7353,N_2373,N_3601);
nand U7354 (N_7354,N_3871,N_3412);
and U7355 (N_7355,N_4694,N_1378);
nand U7356 (N_7356,N_4038,N_265);
xnor U7357 (N_7357,N_1094,N_3219);
and U7358 (N_7358,N_1745,N_2819);
or U7359 (N_7359,N_3950,N_3225);
or U7360 (N_7360,N_4572,N_612);
and U7361 (N_7361,N_4727,N_2343);
nor U7362 (N_7362,N_1038,N_4680);
or U7363 (N_7363,N_3740,N_1780);
xor U7364 (N_7364,N_217,N_3858);
and U7365 (N_7365,N_3548,N_2251);
xnor U7366 (N_7366,N_736,N_997);
nor U7367 (N_7367,N_2442,N_1002);
and U7368 (N_7368,N_3334,N_2346);
or U7369 (N_7369,N_1081,N_2433);
nor U7370 (N_7370,N_548,N_2530);
nor U7371 (N_7371,N_856,N_2795);
and U7372 (N_7372,N_4452,N_4530);
or U7373 (N_7373,N_1357,N_1552);
and U7374 (N_7374,N_4440,N_4186);
nand U7375 (N_7375,N_3193,N_4917);
nor U7376 (N_7376,N_916,N_1235);
nor U7377 (N_7377,N_616,N_2676);
xor U7378 (N_7378,N_2024,N_2667);
xor U7379 (N_7379,N_1511,N_1887);
or U7380 (N_7380,N_1042,N_668);
nand U7381 (N_7381,N_3748,N_3535);
nand U7382 (N_7382,N_2328,N_1604);
nor U7383 (N_7383,N_4568,N_89);
nand U7384 (N_7384,N_1757,N_3525);
and U7385 (N_7385,N_2837,N_621);
and U7386 (N_7386,N_1946,N_4659);
nand U7387 (N_7387,N_893,N_3443);
nand U7388 (N_7388,N_2426,N_2268);
nor U7389 (N_7389,N_1782,N_2010);
and U7390 (N_7390,N_4311,N_2493);
nor U7391 (N_7391,N_1237,N_2000);
and U7392 (N_7392,N_4725,N_3743);
and U7393 (N_7393,N_1443,N_4334);
nor U7394 (N_7394,N_703,N_4806);
nor U7395 (N_7395,N_4349,N_55);
xor U7396 (N_7396,N_3612,N_4796);
and U7397 (N_7397,N_2669,N_1975);
or U7398 (N_7398,N_834,N_2507);
or U7399 (N_7399,N_4238,N_1998);
nand U7400 (N_7400,N_4496,N_4255);
and U7401 (N_7401,N_2215,N_1544);
nor U7402 (N_7402,N_103,N_2729);
and U7403 (N_7403,N_3402,N_1149);
and U7404 (N_7404,N_4161,N_749);
and U7405 (N_7405,N_4127,N_1545);
nor U7406 (N_7406,N_2889,N_960);
or U7407 (N_7407,N_60,N_828);
nand U7408 (N_7408,N_3590,N_333);
and U7409 (N_7409,N_3487,N_70);
nor U7410 (N_7410,N_4006,N_4226);
and U7411 (N_7411,N_4416,N_4231);
nor U7412 (N_7412,N_124,N_4050);
or U7413 (N_7413,N_1759,N_1173);
and U7414 (N_7414,N_3249,N_2626);
nor U7415 (N_7415,N_693,N_3861);
nor U7416 (N_7416,N_2528,N_1884);
and U7417 (N_7417,N_2648,N_4147);
nand U7418 (N_7418,N_4717,N_4863);
nor U7419 (N_7419,N_4171,N_3680);
and U7420 (N_7420,N_4414,N_65);
or U7421 (N_7421,N_4268,N_385);
and U7422 (N_7422,N_4170,N_1238);
nand U7423 (N_7423,N_4192,N_825);
or U7424 (N_7424,N_94,N_3755);
and U7425 (N_7425,N_3066,N_3255);
or U7426 (N_7426,N_3709,N_3527);
and U7427 (N_7427,N_3614,N_3550);
nor U7428 (N_7428,N_376,N_1924);
or U7429 (N_7429,N_2115,N_1271);
or U7430 (N_7430,N_2074,N_4142);
xor U7431 (N_7431,N_1413,N_1012);
nor U7432 (N_7432,N_3058,N_770);
nand U7433 (N_7433,N_4601,N_1057);
and U7434 (N_7434,N_4767,N_2806);
nor U7435 (N_7435,N_516,N_1523);
nand U7436 (N_7436,N_4361,N_3368);
and U7437 (N_7437,N_799,N_2257);
nor U7438 (N_7438,N_3708,N_3175);
xnor U7439 (N_7439,N_1129,N_4742);
nor U7440 (N_7440,N_4534,N_220);
and U7441 (N_7441,N_1049,N_3290);
and U7442 (N_7442,N_2156,N_823);
nor U7443 (N_7443,N_4299,N_1335);
xnor U7444 (N_7444,N_2375,N_3514);
and U7445 (N_7445,N_876,N_2435);
or U7446 (N_7446,N_1349,N_3490);
nand U7447 (N_7447,N_4657,N_2390);
or U7448 (N_7448,N_877,N_1882);
and U7449 (N_7449,N_2295,N_4645);
or U7450 (N_7450,N_4206,N_4278);
nand U7451 (N_7451,N_2811,N_1314);
xor U7452 (N_7452,N_4071,N_4498);
nand U7453 (N_7453,N_2782,N_3927);
nor U7454 (N_7454,N_4267,N_3892);
xnor U7455 (N_7455,N_2255,N_3375);
nand U7456 (N_7456,N_4423,N_2360);
nand U7457 (N_7457,N_2258,N_973);
nor U7458 (N_7458,N_2643,N_1367);
xnor U7459 (N_7459,N_391,N_3063);
or U7460 (N_7460,N_866,N_602);
or U7461 (N_7461,N_2009,N_590);
nand U7462 (N_7462,N_2721,N_4066);
nand U7463 (N_7463,N_521,N_210);
nand U7464 (N_7464,N_1944,N_1111);
xor U7465 (N_7465,N_207,N_1452);
and U7466 (N_7466,N_3026,N_3591);
nor U7467 (N_7467,N_906,N_3214);
nand U7468 (N_7468,N_2386,N_3346);
nor U7469 (N_7469,N_871,N_2448);
nor U7470 (N_7470,N_175,N_4470);
or U7471 (N_7471,N_128,N_289);
and U7472 (N_7472,N_842,N_2844);
nand U7473 (N_7473,N_1559,N_858);
xor U7474 (N_7474,N_3942,N_4101);
nand U7475 (N_7475,N_437,N_2693);
and U7476 (N_7476,N_2836,N_1262);
and U7477 (N_7477,N_2075,N_1320);
or U7478 (N_7478,N_596,N_3118);
and U7479 (N_7479,N_3940,N_2757);
nor U7480 (N_7480,N_2061,N_1732);
and U7481 (N_7481,N_2649,N_4356);
and U7482 (N_7482,N_4548,N_2207);
nand U7483 (N_7483,N_3650,N_1026);
and U7484 (N_7484,N_117,N_1622);
or U7485 (N_7485,N_2506,N_4517);
nor U7486 (N_7486,N_2367,N_1250);
nor U7487 (N_7487,N_4794,N_3318);
or U7488 (N_7488,N_2443,N_831);
and U7489 (N_7489,N_4508,N_3401);
or U7490 (N_7490,N_2963,N_1193);
or U7491 (N_7491,N_1797,N_938);
or U7492 (N_7492,N_4386,N_2826);
or U7493 (N_7493,N_3139,N_3750);
nor U7494 (N_7494,N_129,N_268);
nand U7495 (N_7495,N_1991,N_4849);
nand U7496 (N_7496,N_1806,N_2459);
or U7497 (N_7497,N_533,N_1790);
nor U7498 (N_7498,N_3313,N_1007);
or U7499 (N_7499,N_2456,N_661);
xor U7500 (N_7500,N_3292,N_4540);
nor U7501 (N_7501,N_4902,N_4031);
and U7502 (N_7502,N_2963,N_877);
and U7503 (N_7503,N_622,N_4230);
and U7504 (N_7504,N_168,N_4011);
and U7505 (N_7505,N_3385,N_2723);
nand U7506 (N_7506,N_748,N_277);
nand U7507 (N_7507,N_1894,N_1370);
nor U7508 (N_7508,N_3410,N_4222);
or U7509 (N_7509,N_1764,N_2933);
xnor U7510 (N_7510,N_902,N_1891);
nand U7511 (N_7511,N_1253,N_61);
nand U7512 (N_7512,N_1161,N_3676);
nor U7513 (N_7513,N_3242,N_1936);
nand U7514 (N_7514,N_1355,N_2720);
xnor U7515 (N_7515,N_3834,N_4434);
and U7516 (N_7516,N_2539,N_4401);
nor U7517 (N_7517,N_3542,N_4398);
and U7518 (N_7518,N_4095,N_2423);
or U7519 (N_7519,N_622,N_3781);
or U7520 (N_7520,N_3484,N_685);
xnor U7521 (N_7521,N_2525,N_2298);
nor U7522 (N_7522,N_1454,N_2788);
nand U7523 (N_7523,N_290,N_2766);
nand U7524 (N_7524,N_2855,N_749);
nand U7525 (N_7525,N_1475,N_1836);
and U7526 (N_7526,N_3354,N_4576);
xnor U7527 (N_7527,N_3541,N_2772);
xor U7528 (N_7528,N_4983,N_615);
and U7529 (N_7529,N_3862,N_1032);
or U7530 (N_7530,N_3897,N_731);
xnor U7531 (N_7531,N_4392,N_2594);
nand U7532 (N_7532,N_235,N_4559);
nor U7533 (N_7533,N_614,N_4861);
xnor U7534 (N_7534,N_4563,N_2764);
xor U7535 (N_7535,N_3657,N_1963);
and U7536 (N_7536,N_1802,N_2968);
and U7537 (N_7537,N_3269,N_3977);
xor U7538 (N_7538,N_1593,N_2324);
or U7539 (N_7539,N_1322,N_4489);
xor U7540 (N_7540,N_4869,N_856);
nand U7541 (N_7541,N_4394,N_777);
nand U7542 (N_7542,N_2891,N_317);
nand U7543 (N_7543,N_3748,N_2468);
or U7544 (N_7544,N_3112,N_2931);
nor U7545 (N_7545,N_529,N_1153);
xor U7546 (N_7546,N_2866,N_2096);
nor U7547 (N_7547,N_2612,N_414);
or U7548 (N_7548,N_3804,N_259);
nand U7549 (N_7549,N_2448,N_311);
nor U7550 (N_7550,N_1150,N_4629);
nor U7551 (N_7551,N_1023,N_3579);
or U7552 (N_7552,N_2344,N_3852);
xor U7553 (N_7553,N_4565,N_1059);
nand U7554 (N_7554,N_2875,N_1415);
and U7555 (N_7555,N_2476,N_2108);
nand U7556 (N_7556,N_238,N_4552);
and U7557 (N_7557,N_3385,N_2483);
and U7558 (N_7558,N_1551,N_4208);
nor U7559 (N_7559,N_1350,N_4681);
or U7560 (N_7560,N_4338,N_3782);
xnor U7561 (N_7561,N_3304,N_379);
and U7562 (N_7562,N_2091,N_2121);
or U7563 (N_7563,N_2405,N_2883);
xor U7564 (N_7564,N_1541,N_9);
and U7565 (N_7565,N_558,N_2375);
nand U7566 (N_7566,N_65,N_214);
and U7567 (N_7567,N_4315,N_751);
nor U7568 (N_7568,N_771,N_2726);
or U7569 (N_7569,N_4648,N_39);
nand U7570 (N_7570,N_4347,N_1700);
or U7571 (N_7571,N_2451,N_3465);
nor U7572 (N_7572,N_4603,N_563);
nor U7573 (N_7573,N_4054,N_828);
xnor U7574 (N_7574,N_2358,N_1300);
nor U7575 (N_7575,N_1472,N_834);
nor U7576 (N_7576,N_1140,N_1162);
or U7577 (N_7577,N_3484,N_1418);
nor U7578 (N_7578,N_1029,N_4835);
nand U7579 (N_7579,N_610,N_2964);
nand U7580 (N_7580,N_1219,N_4482);
and U7581 (N_7581,N_1283,N_3298);
nor U7582 (N_7582,N_3646,N_4972);
xor U7583 (N_7583,N_3188,N_1328);
nand U7584 (N_7584,N_4914,N_4120);
and U7585 (N_7585,N_2718,N_4941);
or U7586 (N_7586,N_3442,N_2364);
and U7587 (N_7587,N_157,N_2152);
nor U7588 (N_7588,N_2470,N_1872);
xnor U7589 (N_7589,N_3576,N_1187);
nand U7590 (N_7590,N_4916,N_3874);
nor U7591 (N_7591,N_1797,N_3055);
or U7592 (N_7592,N_3820,N_414);
nand U7593 (N_7593,N_2397,N_2879);
nor U7594 (N_7594,N_3646,N_1368);
nor U7595 (N_7595,N_2134,N_4468);
nand U7596 (N_7596,N_3334,N_733);
nor U7597 (N_7597,N_1838,N_1132);
or U7598 (N_7598,N_3845,N_707);
nand U7599 (N_7599,N_1462,N_3033);
nand U7600 (N_7600,N_2073,N_846);
nand U7601 (N_7601,N_1915,N_4980);
nor U7602 (N_7602,N_1416,N_944);
and U7603 (N_7603,N_34,N_2635);
xnor U7604 (N_7604,N_86,N_2057);
or U7605 (N_7605,N_3889,N_2464);
nand U7606 (N_7606,N_181,N_2396);
nor U7607 (N_7607,N_541,N_3530);
or U7608 (N_7608,N_2549,N_321);
and U7609 (N_7609,N_4463,N_1666);
xor U7610 (N_7610,N_4908,N_2545);
and U7611 (N_7611,N_1341,N_2450);
nand U7612 (N_7612,N_2467,N_318);
xor U7613 (N_7613,N_857,N_1083);
and U7614 (N_7614,N_4890,N_116);
or U7615 (N_7615,N_4572,N_4701);
xnor U7616 (N_7616,N_806,N_2279);
nand U7617 (N_7617,N_3274,N_849);
and U7618 (N_7618,N_379,N_2520);
and U7619 (N_7619,N_2136,N_2838);
or U7620 (N_7620,N_867,N_862);
or U7621 (N_7621,N_3144,N_577);
and U7622 (N_7622,N_4391,N_2435);
nor U7623 (N_7623,N_1011,N_3783);
and U7624 (N_7624,N_3397,N_1816);
or U7625 (N_7625,N_3633,N_4625);
and U7626 (N_7626,N_2088,N_378);
or U7627 (N_7627,N_59,N_1914);
nand U7628 (N_7628,N_1046,N_4909);
nand U7629 (N_7629,N_3011,N_1648);
and U7630 (N_7630,N_4373,N_1328);
and U7631 (N_7631,N_1603,N_587);
and U7632 (N_7632,N_591,N_318);
and U7633 (N_7633,N_1119,N_281);
and U7634 (N_7634,N_3724,N_2497);
and U7635 (N_7635,N_608,N_4048);
xnor U7636 (N_7636,N_4933,N_3235);
nor U7637 (N_7637,N_3915,N_1994);
and U7638 (N_7638,N_764,N_4155);
nor U7639 (N_7639,N_2765,N_1175);
xnor U7640 (N_7640,N_3424,N_3894);
or U7641 (N_7641,N_709,N_4555);
xor U7642 (N_7642,N_724,N_4581);
nor U7643 (N_7643,N_1969,N_3503);
or U7644 (N_7644,N_4779,N_3671);
nor U7645 (N_7645,N_4944,N_2899);
nand U7646 (N_7646,N_4577,N_1177);
nand U7647 (N_7647,N_3940,N_1923);
nand U7648 (N_7648,N_578,N_1852);
and U7649 (N_7649,N_4356,N_597);
and U7650 (N_7650,N_1960,N_1136);
xnor U7651 (N_7651,N_2298,N_443);
nand U7652 (N_7652,N_366,N_958);
xor U7653 (N_7653,N_4519,N_1487);
and U7654 (N_7654,N_2428,N_3688);
and U7655 (N_7655,N_3270,N_1850);
nor U7656 (N_7656,N_3501,N_641);
nor U7657 (N_7657,N_1634,N_394);
nand U7658 (N_7658,N_4572,N_543);
nand U7659 (N_7659,N_2067,N_3252);
or U7660 (N_7660,N_4694,N_2157);
nand U7661 (N_7661,N_2756,N_2297);
nand U7662 (N_7662,N_1925,N_1506);
or U7663 (N_7663,N_2230,N_4479);
nor U7664 (N_7664,N_3729,N_3803);
nor U7665 (N_7665,N_1402,N_4074);
nand U7666 (N_7666,N_4056,N_3549);
and U7667 (N_7667,N_1401,N_3669);
and U7668 (N_7668,N_247,N_684);
nand U7669 (N_7669,N_4690,N_4093);
nor U7670 (N_7670,N_367,N_2772);
or U7671 (N_7671,N_964,N_4691);
or U7672 (N_7672,N_406,N_2687);
xnor U7673 (N_7673,N_463,N_3385);
and U7674 (N_7674,N_1015,N_3003);
and U7675 (N_7675,N_559,N_2158);
nand U7676 (N_7676,N_327,N_2334);
and U7677 (N_7677,N_1558,N_1749);
nand U7678 (N_7678,N_547,N_2023);
or U7679 (N_7679,N_4190,N_237);
or U7680 (N_7680,N_3776,N_3712);
nand U7681 (N_7681,N_1582,N_3741);
nand U7682 (N_7682,N_2721,N_3427);
xor U7683 (N_7683,N_3652,N_1023);
or U7684 (N_7684,N_247,N_4567);
or U7685 (N_7685,N_3460,N_697);
nand U7686 (N_7686,N_4429,N_1047);
xnor U7687 (N_7687,N_812,N_1936);
or U7688 (N_7688,N_2202,N_2429);
or U7689 (N_7689,N_4111,N_1970);
nor U7690 (N_7690,N_320,N_367);
and U7691 (N_7691,N_3784,N_2845);
and U7692 (N_7692,N_3306,N_1305);
nor U7693 (N_7693,N_1736,N_750);
and U7694 (N_7694,N_4391,N_3004);
or U7695 (N_7695,N_3362,N_2205);
nor U7696 (N_7696,N_3748,N_4967);
or U7697 (N_7697,N_2084,N_2957);
or U7698 (N_7698,N_1922,N_887);
nor U7699 (N_7699,N_2425,N_2841);
nor U7700 (N_7700,N_2787,N_4608);
nand U7701 (N_7701,N_3042,N_3556);
xnor U7702 (N_7702,N_832,N_3906);
and U7703 (N_7703,N_4806,N_1693);
or U7704 (N_7704,N_1203,N_3679);
nor U7705 (N_7705,N_1462,N_347);
and U7706 (N_7706,N_1842,N_3768);
and U7707 (N_7707,N_4985,N_3183);
or U7708 (N_7708,N_3427,N_3113);
nand U7709 (N_7709,N_1142,N_1677);
or U7710 (N_7710,N_3825,N_2500);
nor U7711 (N_7711,N_1800,N_854);
or U7712 (N_7712,N_2398,N_1505);
or U7713 (N_7713,N_3938,N_2961);
nor U7714 (N_7714,N_4125,N_2351);
nor U7715 (N_7715,N_3973,N_2236);
xnor U7716 (N_7716,N_133,N_2148);
or U7717 (N_7717,N_2819,N_4630);
nor U7718 (N_7718,N_1633,N_4306);
xnor U7719 (N_7719,N_2672,N_4677);
nand U7720 (N_7720,N_4688,N_3393);
nand U7721 (N_7721,N_3833,N_3837);
or U7722 (N_7722,N_301,N_1434);
nor U7723 (N_7723,N_2373,N_2872);
nand U7724 (N_7724,N_3920,N_2586);
nor U7725 (N_7725,N_3961,N_1017);
or U7726 (N_7726,N_4390,N_3192);
or U7727 (N_7727,N_4406,N_1159);
nor U7728 (N_7728,N_3177,N_4606);
nand U7729 (N_7729,N_1965,N_307);
and U7730 (N_7730,N_4296,N_869);
and U7731 (N_7731,N_1900,N_1823);
nor U7732 (N_7732,N_3344,N_4597);
nand U7733 (N_7733,N_2038,N_660);
or U7734 (N_7734,N_58,N_2546);
or U7735 (N_7735,N_2378,N_2331);
nor U7736 (N_7736,N_199,N_1061);
nand U7737 (N_7737,N_2282,N_1641);
and U7738 (N_7738,N_3510,N_4979);
or U7739 (N_7739,N_237,N_1980);
or U7740 (N_7740,N_2379,N_2718);
nand U7741 (N_7741,N_4184,N_1050);
nand U7742 (N_7742,N_3769,N_2471);
nor U7743 (N_7743,N_3371,N_1072);
nor U7744 (N_7744,N_2798,N_3468);
and U7745 (N_7745,N_619,N_3958);
and U7746 (N_7746,N_4670,N_3142);
or U7747 (N_7747,N_687,N_1291);
nand U7748 (N_7748,N_1290,N_4207);
xnor U7749 (N_7749,N_2847,N_372);
or U7750 (N_7750,N_2296,N_4166);
nand U7751 (N_7751,N_36,N_3327);
or U7752 (N_7752,N_2866,N_3433);
or U7753 (N_7753,N_4777,N_2743);
nor U7754 (N_7754,N_722,N_1729);
nand U7755 (N_7755,N_155,N_1579);
or U7756 (N_7756,N_1886,N_4580);
and U7757 (N_7757,N_4421,N_108);
nor U7758 (N_7758,N_4667,N_1885);
or U7759 (N_7759,N_3058,N_4980);
nor U7760 (N_7760,N_237,N_4155);
or U7761 (N_7761,N_1258,N_3749);
and U7762 (N_7762,N_2215,N_405);
or U7763 (N_7763,N_3868,N_426);
or U7764 (N_7764,N_896,N_506);
nor U7765 (N_7765,N_1278,N_2449);
nor U7766 (N_7766,N_322,N_1611);
and U7767 (N_7767,N_1298,N_4471);
nor U7768 (N_7768,N_3976,N_2983);
and U7769 (N_7769,N_2606,N_508);
xnor U7770 (N_7770,N_213,N_1416);
nand U7771 (N_7771,N_4434,N_1571);
nor U7772 (N_7772,N_1120,N_117);
and U7773 (N_7773,N_4414,N_4953);
nand U7774 (N_7774,N_3921,N_1737);
nor U7775 (N_7775,N_1412,N_3201);
xor U7776 (N_7776,N_703,N_666);
nor U7777 (N_7777,N_4879,N_4388);
and U7778 (N_7778,N_2170,N_2516);
and U7779 (N_7779,N_510,N_2509);
and U7780 (N_7780,N_3130,N_436);
nand U7781 (N_7781,N_313,N_621);
nor U7782 (N_7782,N_853,N_2101);
and U7783 (N_7783,N_3212,N_4801);
nor U7784 (N_7784,N_3565,N_2170);
and U7785 (N_7785,N_3120,N_487);
nand U7786 (N_7786,N_2836,N_2141);
xor U7787 (N_7787,N_942,N_814);
and U7788 (N_7788,N_3314,N_1184);
nand U7789 (N_7789,N_4077,N_91);
or U7790 (N_7790,N_3611,N_4454);
and U7791 (N_7791,N_379,N_4096);
nor U7792 (N_7792,N_4737,N_331);
nor U7793 (N_7793,N_365,N_3736);
nand U7794 (N_7794,N_707,N_4381);
or U7795 (N_7795,N_4450,N_2689);
or U7796 (N_7796,N_3794,N_719);
nand U7797 (N_7797,N_2924,N_3429);
nor U7798 (N_7798,N_4299,N_2703);
and U7799 (N_7799,N_4491,N_4975);
nor U7800 (N_7800,N_2319,N_4739);
and U7801 (N_7801,N_1911,N_1979);
and U7802 (N_7802,N_1441,N_2463);
nand U7803 (N_7803,N_2652,N_177);
and U7804 (N_7804,N_1095,N_2851);
nand U7805 (N_7805,N_4355,N_2564);
nand U7806 (N_7806,N_2306,N_552);
nor U7807 (N_7807,N_4464,N_3179);
or U7808 (N_7808,N_2081,N_3408);
and U7809 (N_7809,N_1464,N_2917);
xor U7810 (N_7810,N_944,N_4272);
nand U7811 (N_7811,N_3326,N_3556);
nor U7812 (N_7812,N_4342,N_3175);
xnor U7813 (N_7813,N_2097,N_462);
or U7814 (N_7814,N_4636,N_2824);
and U7815 (N_7815,N_4038,N_2751);
xnor U7816 (N_7816,N_3209,N_446);
nor U7817 (N_7817,N_2495,N_4925);
or U7818 (N_7818,N_1988,N_2506);
nand U7819 (N_7819,N_3547,N_82);
or U7820 (N_7820,N_1101,N_3249);
nand U7821 (N_7821,N_822,N_3997);
and U7822 (N_7822,N_3741,N_1470);
and U7823 (N_7823,N_430,N_4284);
nor U7824 (N_7824,N_4409,N_4433);
and U7825 (N_7825,N_4746,N_4029);
nand U7826 (N_7826,N_630,N_4452);
nor U7827 (N_7827,N_3195,N_3596);
xnor U7828 (N_7828,N_881,N_4330);
and U7829 (N_7829,N_4594,N_197);
xor U7830 (N_7830,N_4060,N_914);
nor U7831 (N_7831,N_4891,N_1724);
nand U7832 (N_7832,N_2792,N_1035);
xor U7833 (N_7833,N_3562,N_1750);
and U7834 (N_7834,N_2783,N_952);
nand U7835 (N_7835,N_745,N_4657);
or U7836 (N_7836,N_1637,N_305);
or U7837 (N_7837,N_415,N_532);
and U7838 (N_7838,N_2434,N_2775);
xor U7839 (N_7839,N_1087,N_1416);
nor U7840 (N_7840,N_1734,N_1625);
nand U7841 (N_7841,N_7,N_779);
nor U7842 (N_7842,N_722,N_3967);
nand U7843 (N_7843,N_1439,N_398);
nand U7844 (N_7844,N_3892,N_2608);
and U7845 (N_7845,N_491,N_849);
and U7846 (N_7846,N_1826,N_1341);
and U7847 (N_7847,N_304,N_4102);
nand U7848 (N_7848,N_534,N_1970);
and U7849 (N_7849,N_2528,N_2519);
or U7850 (N_7850,N_1171,N_4298);
nor U7851 (N_7851,N_2703,N_886);
nand U7852 (N_7852,N_1635,N_3274);
nor U7853 (N_7853,N_4171,N_4414);
and U7854 (N_7854,N_3917,N_3763);
nor U7855 (N_7855,N_3747,N_3959);
or U7856 (N_7856,N_3726,N_4977);
xnor U7857 (N_7857,N_4103,N_1627);
nor U7858 (N_7858,N_4470,N_4690);
or U7859 (N_7859,N_845,N_3439);
and U7860 (N_7860,N_4124,N_4399);
or U7861 (N_7861,N_2770,N_2701);
or U7862 (N_7862,N_2318,N_4762);
and U7863 (N_7863,N_1287,N_497);
and U7864 (N_7864,N_3051,N_430);
nor U7865 (N_7865,N_1349,N_1850);
and U7866 (N_7866,N_3987,N_1722);
or U7867 (N_7867,N_1048,N_4407);
nand U7868 (N_7868,N_2375,N_3611);
nor U7869 (N_7869,N_2440,N_4646);
nand U7870 (N_7870,N_1397,N_766);
or U7871 (N_7871,N_3995,N_3203);
nor U7872 (N_7872,N_1828,N_2688);
nor U7873 (N_7873,N_1305,N_3307);
or U7874 (N_7874,N_98,N_2262);
nand U7875 (N_7875,N_69,N_2538);
and U7876 (N_7876,N_3393,N_3008);
or U7877 (N_7877,N_393,N_2906);
nor U7878 (N_7878,N_1160,N_2538);
nor U7879 (N_7879,N_2123,N_2006);
or U7880 (N_7880,N_3905,N_1173);
and U7881 (N_7881,N_1376,N_1289);
or U7882 (N_7882,N_2105,N_4790);
nand U7883 (N_7883,N_4891,N_3495);
and U7884 (N_7884,N_4203,N_832);
nand U7885 (N_7885,N_3218,N_1882);
nor U7886 (N_7886,N_2497,N_3317);
and U7887 (N_7887,N_3847,N_3722);
nor U7888 (N_7888,N_1283,N_4917);
nor U7889 (N_7889,N_1205,N_2343);
nor U7890 (N_7890,N_1923,N_4830);
and U7891 (N_7891,N_3548,N_3748);
nor U7892 (N_7892,N_1906,N_1331);
and U7893 (N_7893,N_3233,N_1379);
or U7894 (N_7894,N_1395,N_4833);
xnor U7895 (N_7895,N_2679,N_1568);
nor U7896 (N_7896,N_3691,N_2279);
or U7897 (N_7897,N_871,N_2945);
nor U7898 (N_7898,N_4045,N_2159);
or U7899 (N_7899,N_4493,N_4107);
and U7900 (N_7900,N_1390,N_4412);
and U7901 (N_7901,N_4890,N_2163);
xor U7902 (N_7902,N_987,N_4254);
or U7903 (N_7903,N_3248,N_4692);
xnor U7904 (N_7904,N_2267,N_420);
nor U7905 (N_7905,N_3349,N_1751);
and U7906 (N_7906,N_4844,N_137);
nand U7907 (N_7907,N_2678,N_2566);
and U7908 (N_7908,N_2162,N_4358);
xor U7909 (N_7909,N_463,N_2047);
xor U7910 (N_7910,N_1764,N_1064);
or U7911 (N_7911,N_4709,N_319);
or U7912 (N_7912,N_3939,N_1762);
and U7913 (N_7913,N_29,N_2211);
nand U7914 (N_7914,N_1237,N_3093);
nand U7915 (N_7915,N_4011,N_1951);
nor U7916 (N_7916,N_2820,N_730);
nor U7917 (N_7917,N_3377,N_4921);
and U7918 (N_7918,N_4637,N_2425);
nor U7919 (N_7919,N_2848,N_2646);
and U7920 (N_7920,N_4560,N_352);
xor U7921 (N_7921,N_994,N_3795);
nand U7922 (N_7922,N_1700,N_1892);
or U7923 (N_7923,N_294,N_1276);
or U7924 (N_7924,N_4398,N_3135);
or U7925 (N_7925,N_3375,N_4971);
xor U7926 (N_7926,N_70,N_807);
nor U7927 (N_7927,N_3761,N_3567);
or U7928 (N_7928,N_1653,N_4196);
nor U7929 (N_7929,N_4313,N_3234);
nor U7930 (N_7930,N_2438,N_4404);
nor U7931 (N_7931,N_4956,N_3889);
or U7932 (N_7932,N_1250,N_2087);
nor U7933 (N_7933,N_3795,N_3831);
and U7934 (N_7934,N_2830,N_1802);
or U7935 (N_7935,N_237,N_4228);
and U7936 (N_7936,N_949,N_4322);
or U7937 (N_7937,N_4068,N_2292);
nand U7938 (N_7938,N_418,N_4184);
or U7939 (N_7939,N_1688,N_1452);
nand U7940 (N_7940,N_2234,N_1797);
nand U7941 (N_7941,N_1347,N_1956);
nand U7942 (N_7942,N_1478,N_2887);
or U7943 (N_7943,N_1402,N_1718);
or U7944 (N_7944,N_4317,N_2439);
or U7945 (N_7945,N_687,N_2197);
xnor U7946 (N_7946,N_4939,N_4144);
nor U7947 (N_7947,N_3947,N_167);
nor U7948 (N_7948,N_2483,N_1529);
nor U7949 (N_7949,N_2313,N_304);
nand U7950 (N_7950,N_2844,N_1010);
nand U7951 (N_7951,N_2539,N_3976);
nor U7952 (N_7952,N_2394,N_1730);
nand U7953 (N_7953,N_3397,N_2499);
xnor U7954 (N_7954,N_4756,N_4962);
and U7955 (N_7955,N_4006,N_890);
nor U7956 (N_7956,N_3621,N_1691);
and U7957 (N_7957,N_4061,N_2865);
nand U7958 (N_7958,N_266,N_4869);
nand U7959 (N_7959,N_1769,N_2693);
nor U7960 (N_7960,N_2446,N_4424);
xor U7961 (N_7961,N_4141,N_3152);
nand U7962 (N_7962,N_1,N_4134);
or U7963 (N_7963,N_12,N_3484);
nor U7964 (N_7964,N_2155,N_3092);
and U7965 (N_7965,N_3620,N_3712);
nor U7966 (N_7966,N_3521,N_4008);
nand U7967 (N_7967,N_3516,N_1411);
nand U7968 (N_7968,N_4197,N_350);
and U7969 (N_7969,N_3800,N_3931);
or U7970 (N_7970,N_2086,N_4882);
nor U7971 (N_7971,N_4683,N_2407);
nand U7972 (N_7972,N_1403,N_70);
or U7973 (N_7973,N_2707,N_2480);
or U7974 (N_7974,N_2026,N_301);
nand U7975 (N_7975,N_2816,N_4352);
nand U7976 (N_7976,N_2673,N_3533);
nand U7977 (N_7977,N_1892,N_1293);
and U7978 (N_7978,N_4411,N_4747);
and U7979 (N_7979,N_614,N_3281);
or U7980 (N_7980,N_138,N_204);
or U7981 (N_7981,N_3295,N_743);
nor U7982 (N_7982,N_816,N_1465);
nor U7983 (N_7983,N_1074,N_3708);
or U7984 (N_7984,N_156,N_3313);
nand U7985 (N_7985,N_731,N_3447);
nand U7986 (N_7986,N_3258,N_62);
or U7987 (N_7987,N_4285,N_2478);
nand U7988 (N_7988,N_902,N_1638);
and U7989 (N_7989,N_256,N_3158);
or U7990 (N_7990,N_3186,N_3809);
and U7991 (N_7991,N_276,N_1673);
xnor U7992 (N_7992,N_3971,N_78);
nor U7993 (N_7993,N_2454,N_3665);
or U7994 (N_7994,N_4846,N_3570);
nor U7995 (N_7995,N_1179,N_874);
or U7996 (N_7996,N_1443,N_2956);
xor U7997 (N_7997,N_4051,N_1424);
xor U7998 (N_7998,N_2564,N_4747);
xor U7999 (N_7999,N_2813,N_225);
nor U8000 (N_8000,N_4004,N_653);
nor U8001 (N_8001,N_3854,N_4736);
or U8002 (N_8002,N_3219,N_1217);
nor U8003 (N_8003,N_1206,N_4684);
and U8004 (N_8004,N_1904,N_1535);
nor U8005 (N_8005,N_833,N_4245);
nor U8006 (N_8006,N_1466,N_2165);
or U8007 (N_8007,N_3629,N_4927);
nand U8008 (N_8008,N_2324,N_1508);
nor U8009 (N_8009,N_4134,N_4250);
or U8010 (N_8010,N_2770,N_579);
nor U8011 (N_8011,N_3852,N_2832);
and U8012 (N_8012,N_3114,N_3313);
and U8013 (N_8013,N_1472,N_1412);
nand U8014 (N_8014,N_1478,N_4175);
nor U8015 (N_8015,N_571,N_3378);
xnor U8016 (N_8016,N_3425,N_2501);
nor U8017 (N_8017,N_1018,N_2938);
nand U8018 (N_8018,N_357,N_3284);
nand U8019 (N_8019,N_1304,N_4167);
and U8020 (N_8020,N_2775,N_4031);
or U8021 (N_8021,N_1774,N_4490);
and U8022 (N_8022,N_3146,N_290);
xor U8023 (N_8023,N_1242,N_280);
or U8024 (N_8024,N_124,N_4884);
nor U8025 (N_8025,N_998,N_2243);
nand U8026 (N_8026,N_4246,N_4187);
and U8027 (N_8027,N_4719,N_3139);
nor U8028 (N_8028,N_2055,N_1591);
nand U8029 (N_8029,N_4738,N_1634);
nand U8030 (N_8030,N_3543,N_1603);
or U8031 (N_8031,N_2446,N_166);
or U8032 (N_8032,N_2709,N_759);
and U8033 (N_8033,N_2747,N_1954);
nor U8034 (N_8034,N_1059,N_26);
nand U8035 (N_8035,N_4086,N_4186);
nand U8036 (N_8036,N_4759,N_4803);
nand U8037 (N_8037,N_4473,N_2888);
nand U8038 (N_8038,N_1812,N_1540);
nand U8039 (N_8039,N_185,N_2593);
xor U8040 (N_8040,N_2168,N_3526);
and U8041 (N_8041,N_3848,N_1924);
xnor U8042 (N_8042,N_4444,N_3506);
or U8043 (N_8043,N_3905,N_4782);
nor U8044 (N_8044,N_3778,N_2508);
nand U8045 (N_8045,N_4511,N_52);
and U8046 (N_8046,N_2917,N_1135);
nand U8047 (N_8047,N_212,N_1541);
nor U8048 (N_8048,N_4445,N_1257);
or U8049 (N_8049,N_1843,N_2010);
nor U8050 (N_8050,N_480,N_1497);
xor U8051 (N_8051,N_3653,N_3520);
or U8052 (N_8052,N_4371,N_1392);
or U8053 (N_8053,N_304,N_4707);
and U8054 (N_8054,N_3039,N_1666);
nand U8055 (N_8055,N_1761,N_1674);
or U8056 (N_8056,N_1348,N_2616);
or U8057 (N_8057,N_741,N_1062);
xor U8058 (N_8058,N_3189,N_1601);
and U8059 (N_8059,N_3697,N_4998);
or U8060 (N_8060,N_1193,N_3492);
nand U8061 (N_8061,N_4640,N_628);
and U8062 (N_8062,N_2011,N_3370);
or U8063 (N_8063,N_745,N_3131);
xnor U8064 (N_8064,N_1419,N_2722);
nand U8065 (N_8065,N_1549,N_3748);
nand U8066 (N_8066,N_1511,N_3174);
nor U8067 (N_8067,N_3678,N_1007);
nor U8068 (N_8068,N_3802,N_4521);
nand U8069 (N_8069,N_2162,N_4972);
xor U8070 (N_8070,N_824,N_960);
nor U8071 (N_8071,N_1307,N_3008);
or U8072 (N_8072,N_3713,N_381);
or U8073 (N_8073,N_3481,N_3127);
and U8074 (N_8074,N_457,N_851);
nand U8075 (N_8075,N_877,N_1372);
nand U8076 (N_8076,N_4320,N_2815);
and U8077 (N_8077,N_3446,N_2682);
nand U8078 (N_8078,N_788,N_4193);
or U8079 (N_8079,N_2298,N_1678);
or U8080 (N_8080,N_3204,N_2470);
or U8081 (N_8081,N_2017,N_3206);
and U8082 (N_8082,N_978,N_2914);
xnor U8083 (N_8083,N_1537,N_4048);
xnor U8084 (N_8084,N_4797,N_4036);
nor U8085 (N_8085,N_2862,N_4074);
nor U8086 (N_8086,N_1223,N_2479);
nor U8087 (N_8087,N_2847,N_2449);
and U8088 (N_8088,N_1960,N_4715);
or U8089 (N_8089,N_2508,N_3824);
and U8090 (N_8090,N_829,N_1221);
and U8091 (N_8091,N_1523,N_2627);
nand U8092 (N_8092,N_3404,N_3140);
nand U8093 (N_8093,N_4988,N_248);
nor U8094 (N_8094,N_1002,N_2127);
or U8095 (N_8095,N_2560,N_2910);
nor U8096 (N_8096,N_3339,N_2677);
and U8097 (N_8097,N_38,N_3011);
nand U8098 (N_8098,N_3245,N_3530);
nand U8099 (N_8099,N_3926,N_3855);
nand U8100 (N_8100,N_1786,N_4141);
and U8101 (N_8101,N_4931,N_1003);
nor U8102 (N_8102,N_920,N_2673);
nand U8103 (N_8103,N_4452,N_4455);
and U8104 (N_8104,N_2827,N_2680);
and U8105 (N_8105,N_4691,N_4208);
nor U8106 (N_8106,N_1273,N_2938);
and U8107 (N_8107,N_1386,N_2607);
nor U8108 (N_8108,N_2442,N_3000);
and U8109 (N_8109,N_2719,N_2010);
xnor U8110 (N_8110,N_2562,N_4902);
xnor U8111 (N_8111,N_3635,N_4159);
nor U8112 (N_8112,N_3341,N_4392);
or U8113 (N_8113,N_4126,N_2701);
and U8114 (N_8114,N_4908,N_4014);
and U8115 (N_8115,N_2552,N_2935);
nor U8116 (N_8116,N_4619,N_3113);
nor U8117 (N_8117,N_1885,N_1773);
or U8118 (N_8118,N_2490,N_2688);
or U8119 (N_8119,N_4901,N_166);
nor U8120 (N_8120,N_2550,N_2867);
and U8121 (N_8121,N_1685,N_2902);
xor U8122 (N_8122,N_418,N_973);
nand U8123 (N_8123,N_3007,N_1904);
nand U8124 (N_8124,N_3154,N_4905);
nor U8125 (N_8125,N_3537,N_538);
and U8126 (N_8126,N_815,N_3301);
xnor U8127 (N_8127,N_3513,N_3064);
or U8128 (N_8128,N_3550,N_4247);
or U8129 (N_8129,N_1863,N_332);
nand U8130 (N_8130,N_2345,N_4632);
and U8131 (N_8131,N_3447,N_1182);
nand U8132 (N_8132,N_1945,N_1888);
or U8133 (N_8133,N_873,N_4651);
or U8134 (N_8134,N_4772,N_3380);
or U8135 (N_8135,N_4078,N_1883);
and U8136 (N_8136,N_4426,N_4776);
or U8137 (N_8137,N_1344,N_7);
xor U8138 (N_8138,N_1691,N_4802);
and U8139 (N_8139,N_2877,N_1452);
nand U8140 (N_8140,N_3247,N_532);
nand U8141 (N_8141,N_3111,N_4333);
and U8142 (N_8142,N_2529,N_1530);
nor U8143 (N_8143,N_1333,N_1031);
nor U8144 (N_8144,N_1825,N_2309);
nor U8145 (N_8145,N_3997,N_1759);
or U8146 (N_8146,N_246,N_3957);
nor U8147 (N_8147,N_4780,N_4237);
nor U8148 (N_8148,N_207,N_1598);
or U8149 (N_8149,N_2657,N_2946);
and U8150 (N_8150,N_4114,N_2824);
or U8151 (N_8151,N_2811,N_2189);
nor U8152 (N_8152,N_3377,N_224);
or U8153 (N_8153,N_3630,N_1263);
nand U8154 (N_8154,N_4468,N_4490);
nand U8155 (N_8155,N_3605,N_2676);
and U8156 (N_8156,N_3734,N_598);
or U8157 (N_8157,N_2150,N_2776);
nand U8158 (N_8158,N_4426,N_4280);
and U8159 (N_8159,N_2751,N_1411);
and U8160 (N_8160,N_4359,N_3366);
and U8161 (N_8161,N_4704,N_988);
or U8162 (N_8162,N_2045,N_1573);
nand U8163 (N_8163,N_2041,N_4102);
nor U8164 (N_8164,N_890,N_803);
nor U8165 (N_8165,N_3223,N_3741);
or U8166 (N_8166,N_3804,N_1729);
nand U8167 (N_8167,N_3874,N_2516);
and U8168 (N_8168,N_56,N_2766);
nand U8169 (N_8169,N_2317,N_113);
and U8170 (N_8170,N_4173,N_3137);
nor U8171 (N_8171,N_2807,N_1325);
and U8172 (N_8172,N_879,N_507);
or U8173 (N_8173,N_3142,N_4718);
and U8174 (N_8174,N_4755,N_752);
or U8175 (N_8175,N_3865,N_2248);
and U8176 (N_8176,N_3952,N_3861);
nor U8177 (N_8177,N_331,N_2417);
nor U8178 (N_8178,N_2302,N_3081);
or U8179 (N_8179,N_1365,N_3471);
or U8180 (N_8180,N_853,N_2955);
nor U8181 (N_8181,N_2566,N_3239);
nand U8182 (N_8182,N_305,N_3414);
and U8183 (N_8183,N_4491,N_3147);
nor U8184 (N_8184,N_1033,N_2096);
and U8185 (N_8185,N_4596,N_1391);
nor U8186 (N_8186,N_1848,N_1399);
and U8187 (N_8187,N_1282,N_3263);
xor U8188 (N_8188,N_573,N_4933);
or U8189 (N_8189,N_3412,N_3249);
xor U8190 (N_8190,N_4423,N_2494);
and U8191 (N_8191,N_3923,N_3496);
nor U8192 (N_8192,N_2275,N_1841);
xnor U8193 (N_8193,N_988,N_3311);
or U8194 (N_8194,N_2754,N_3496);
nand U8195 (N_8195,N_1364,N_2711);
nand U8196 (N_8196,N_2067,N_26);
nor U8197 (N_8197,N_4187,N_2436);
nand U8198 (N_8198,N_1304,N_4230);
nand U8199 (N_8199,N_3100,N_1911);
or U8200 (N_8200,N_1458,N_3606);
nor U8201 (N_8201,N_219,N_4866);
nand U8202 (N_8202,N_1574,N_319);
or U8203 (N_8203,N_1553,N_2407);
and U8204 (N_8204,N_4504,N_3290);
nor U8205 (N_8205,N_187,N_1041);
or U8206 (N_8206,N_3604,N_1344);
nor U8207 (N_8207,N_2184,N_208);
or U8208 (N_8208,N_292,N_2586);
xor U8209 (N_8209,N_1046,N_1784);
nor U8210 (N_8210,N_813,N_3884);
or U8211 (N_8211,N_2191,N_1112);
and U8212 (N_8212,N_1245,N_86);
nand U8213 (N_8213,N_3841,N_710);
nand U8214 (N_8214,N_4856,N_2259);
or U8215 (N_8215,N_3727,N_2205);
and U8216 (N_8216,N_2901,N_881);
nor U8217 (N_8217,N_3935,N_2919);
nor U8218 (N_8218,N_2032,N_4258);
nor U8219 (N_8219,N_4444,N_732);
and U8220 (N_8220,N_453,N_3185);
and U8221 (N_8221,N_4729,N_3089);
or U8222 (N_8222,N_213,N_3037);
or U8223 (N_8223,N_2233,N_4943);
and U8224 (N_8224,N_3650,N_3289);
nor U8225 (N_8225,N_1023,N_4370);
and U8226 (N_8226,N_4358,N_4894);
nand U8227 (N_8227,N_2387,N_3904);
or U8228 (N_8228,N_265,N_1971);
nand U8229 (N_8229,N_2850,N_1452);
and U8230 (N_8230,N_2520,N_1274);
or U8231 (N_8231,N_765,N_3599);
and U8232 (N_8232,N_2601,N_889);
and U8233 (N_8233,N_1635,N_788);
or U8234 (N_8234,N_2686,N_865);
and U8235 (N_8235,N_2908,N_1600);
and U8236 (N_8236,N_4473,N_4189);
nand U8237 (N_8237,N_4767,N_3953);
nand U8238 (N_8238,N_2529,N_4200);
or U8239 (N_8239,N_3676,N_3738);
and U8240 (N_8240,N_2745,N_4700);
nor U8241 (N_8241,N_4884,N_4864);
and U8242 (N_8242,N_4675,N_4433);
and U8243 (N_8243,N_3167,N_2908);
and U8244 (N_8244,N_3895,N_2201);
and U8245 (N_8245,N_613,N_396);
xor U8246 (N_8246,N_3148,N_2838);
or U8247 (N_8247,N_3057,N_3431);
nor U8248 (N_8248,N_2980,N_2371);
or U8249 (N_8249,N_486,N_4972);
nand U8250 (N_8250,N_3252,N_3354);
nor U8251 (N_8251,N_789,N_1761);
or U8252 (N_8252,N_1268,N_4990);
and U8253 (N_8253,N_4629,N_4032);
nand U8254 (N_8254,N_4614,N_4661);
nor U8255 (N_8255,N_790,N_2251);
or U8256 (N_8256,N_661,N_331);
and U8257 (N_8257,N_1712,N_806);
nor U8258 (N_8258,N_3249,N_2163);
xor U8259 (N_8259,N_4904,N_1659);
xor U8260 (N_8260,N_3558,N_1393);
nor U8261 (N_8261,N_2942,N_1204);
nor U8262 (N_8262,N_848,N_4917);
or U8263 (N_8263,N_458,N_1271);
xor U8264 (N_8264,N_2874,N_3951);
or U8265 (N_8265,N_95,N_2469);
and U8266 (N_8266,N_4671,N_1131);
nand U8267 (N_8267,N_2681,N_3713);
xnor U8268 (N_8268,N_514,N_1899);
nor U8269 (N_8269,N_1021,N_2256);
or U8270 (N_8270,N_3307,N_3195);
nor U8271 (N_8271,N_1143,N_808);
nand U8272 (N_8272,N_3790,N_2359);
nor U8273 (N_8273,N_1134,N_4548);
and U8274 (N_8274,N_2991,N_4791);
or U8275 (N_8275,N_4519,N_3803);
nand U8276 (N_8276,N_4568,N_4357);
and U8277 (N_8277,N_2461,N_2577);
nand U8278 (N_8278,N_4189,N_3987);
and U8279 (N_8279,N_3528,N_4453);
nand U8280 (N_8280,N_1659,N_4249);
or U8281 (N_8281,N_946,N_3383);
nand U8282 (N_8282,N_3404,N_2836);
or U8283 (N_8283,N_1982,N_2852);
and U8284 (N_8284,N_2387,N_4912);
or U8285 (N_8285,N_416,N_3100);
nand U8286 (N_8286,N_664,N_1545);
or U8287 (N_8287,N_4525,N_552);
xnor U8288 (N_8288,N_1303,N_353);
and U8289 (N_8289,N_143,N_1299);
and U8290 (N_8290,N_3698,N_4320);
nand U8291 (N_8291,N_2379,N_1673);
and U8292 (N_8292,N_2652,N_1147);
or U8293 (N_8293,N_2468,N_4855);
or U8294 (N_8294,N_2519,N_535);
xnor U8295 (N_8295,N_1742,N_45);
nor U8296 (N_8296,N_4866,N_3976);
nand U8297 (N_8297,N_1386,N_1094);
or U8298 (N_8298,N_2657,N_2854);
and U8299 (N_8299,N_3138,N_3307);
or U8300 (N_8300,N_3821,N_2490);
or U8301 (N_8301,N_4574,N_2909);
nand U8302 (N_8302,N_405,N_778);
nor U8303 (N_8303,N_727,N_2728);
xnor U8304 (N_8304,N_2349,N_3624);
nor U8305 (N_8305,N_4245,N_2238);
and U8306 (N_8306,N_3932,N_263);
and U8307 (N_8307,N_4230,N_3188);
or U8308 (N_8308,N_1629,N_474);
nand U8309 (N_8309,N_3192,N_3320);
or U8310 (N_8310,N_3085,N_3179);
nor U8311 (N_8311,N_1319,N_4677);
or U8312 (N_8312,N_4456,N_1943);
or U8313 (N_8313,N_2849,N_3179);
nor U8314 (N_8314,N_4182,N_4410);
nor U8315 (N_8315,N_3307,N_4882);
or U8316 (N_8316,N_2682,N_738);
nor U8317 (N_8317,N_2752,N_3124);
and U8318 (N_8318,N_2082,N_1458);
and U8319 (N_8319,N_1132,N_1874);
or U8320 (N_8320,N_3490,N_834);
or U8321 (N_8321,N_2101,N_2052);
nand U8322 (N_8322,N_2105,N_1825);
xnor U8323 (N_8323,N_590,N_3660);
or U8324 (N_8324,N_4723,N_3979);
nand U8325 (N_8325,N_573,N_4113);
and U8326 (N_8326,N_4529,N_3413);
and U8327 (N_8327,N_2827,N_3176);
and U8328 (N_8328,N_2517,N_3646);
or U8329 (N_8329,N_2979,N_1596);
or U8330 (N_8330,N_1238,N_3074);
nor U8331 (N_8331,N_1971,N_783);
or U8332 (N_8332,N_1066,N_3659);
and U8333 (N_8333,N_2762,N_4138);
xnor U8334 (N_8334,N_2830,N_3558);
nand U8335 (N_8335,N_3737,N_2024);
nor U8336 (N_8336,N_3609,N_2295);
and U8337 (N_8337,N_1253,N_4689);
and U8338 (N_8338,N_2369,N_4570);
and U8339 (N_8339,N_1759,N_4715);
xor U8340 (N_8340,N_1709,N_2715);
and U8341 (N_8341,N_1474,N_3660);
and U8342 (N_8342,N_2089,N_723);
or U8343 (N_8343,N_2072,N_2933);
nand U8344 (N_8344,N_1851,N_4594);
nand U8345 (N_8345,N_3609,N_1399);
or U8346 (N_8346,N_4108,N_1429);
nand U8347 (N_8347,N_1708,N_201);
xnor U8348 (N_8348,N_3754,N_654);
or U8349 (N_8349,N_2870,N_853);
or U8350 (N_8350,N_4769,N_3298);
nand U8351 (N_8351,N_4564,N_722);
nand U8352 (N_8352,N_4698,N_4567);
or U8353 (N_8353,N_3265,N_2321);
nand U8354 (N_8354,N_421,N_2773);
xnor U8355 (N_8355,N_1675,N_4821);
nand U8356 (N_8356,N_306,N_4273);
nand U8357 (N_8357,N_4293,N_3618);
nor U8358 (N_8358,N_4542,N_3828);
nand U8359 (N_8359,N_3993,N_5);
and U8360 (N_8360,N_3619,N_792);
and U8361 (N_8361,N_1388,N_822);
and U8362 (N_8362,N_1942,N_1220);
nand U8363 (N_8363,N_2657,N_4987);
nand U8364 (N_8364,N_375,N_1601);
and U8365 (N_8365,N_4096,N_4250);
and U8366 (N_8366,N_2305,N_259);
and U8367 (N_8367,N_3066,N_4362);
nor U8368 (N_8368,N_3615,N_4349);
and U8369 (N_8369,N_4615,N_4914);
or U8370 (N_8370,N_4282,N_4367);
nor U8371 (N_8371,N_124,N_1364);
nand U8372 (N_8372,N_449,N_1855);
or U8373 (N_8373,N_4761,N_4415);
xnor U8374 (N_8374,N_4781,N_2981);
xnor U8375 (N_8375,N_4374,N_4117);
or U8376 (N_8376,N_1993,N_3889);
nand U8377 (N_8377,N_1244,N_2116);
or U8378 (N_8378,N_2970,N_1676);
nor U8379 (N_8379,N_483,N_1651);
xor U8380 (N_8380,N_1774,N_2587);
nand U8381 (N_8381,N_1240,N_2483);
nand U8382 (N_8382,N_3419,N_2550);
or U8383 (N_8383,N_2266,N_1741);
and U8384 (N_8384,N_4214,N_577);
nand U8385 (N_8385,N_2426,N_3971);
nor U8386 (N_8386,N_4625,N_1086);
xnor U8387 (N_8387,N_1325,N_3730);
nand U8388 (N_8388,N_2089,N_190);
nand U8389 (N_8389,N_1231,N_2067);
and U8390 (N_8390,N_4192,N_1126);
nor U8391 (N_8391,N_2626,N_2494);
or U8392 (N_8392,N_2111,N_89);
nor U8393 (N_8393,N_3195,N_2786);
nor U8394 (N_8394,N_3169,N_4738);
xor U8395 (N_8395,N_1709,N_4418);
nand U8396 (N_8396,N_3766,N_4485);
or U8397 (N_8397,N_1914,N_2488);
and U8398 (N_8398,N_843,N_4668);
nor U8399 (N_8399,N_675,N_1274);
nor U8400 (N_8400,N_248,N_2766);
or U8401 (N_8401,N_2805,N_160);
or U8402 (N_8402,N_627,N_1340);
nor U8403 (N_8403,N_439,N_3372);
nor U8404 (N_8404,N_3908,N_3640);
nand U8405 (N_8405,N_3498,N_1195);
nor U8406 (N_8406,N_696,N_2893);
and U8407 (N_8407,N_2539,N_4812);
xor U8408 (N_8408,N_1535,N_403);
nor U8409 (N_8409,N_1281,N_3228);
and U8410 (N_8410,N_4106,N_2311);
xor U8411 (N_8411,N_3642,N_3434);
nand U8412 (N_8412,N_76,N_4680);
and U8413 (N_8413,N_1317,N_576);
nand U8414 (N_8414,N_1596,N_2624);
nor U8415 (N_8415,N_4845,N_484);
and U8416 (N_8416,N_2918,N_41);
nand U8417 (N_8417,N_2517,N_2074);
nand U8418 (N_8418,N_4805,N_2025);
nor U8419 (N_8419,N_3975,N_441);
nand U8420 (N_8420,N_1323,N_2298);
nand U8421 (N_8421,N_3269,N_191);
nand U8422 (N_8422,N_3855,N_1834);
and U8423 (N_8423,N_4416,N_92);
or U8424 (N_8424,N_2259,N_3442);
nor U8425 (N_8425,N_3293,N_315);
and U8426 (N_8426,N_470,N_1439);
nand U8427 (N_8427,N_1722,N_2497);
or U8428 (N_8428,N_295,N_35);
nor U8429 (N_8429,N_1646,N_2830);
xor U8430 (N_8430,N_4459,N_1030);
nand U8431 (N_8431,N_4000,N_1111);
nor U8432 (N_8432,N_3962,N_3806);
nor U8433 (N_8433,N_941,N_1460);
and U8434 (N_8434,N_3738,N_62);
and U8435 (N_8435,N_1192,N_1783);
and U8436 (N_8436,N_2023,N_4530);
nand U8437 (N_8437,N_4258,N_117);
and U8438 (N_8438,N_4412,N_611);
nor U8439 (N_8439,N_2326,N_2143);
nand U8440 (N_8440,N_1381,N_1037);
nor U8441 (N_8441,N_3152,N_892);
or U8442 (N_8442,N_3955,N_2102);
nor U8443 (N_8443,N_1370,N_1001);
nor U8444 (N_8444,N_4771,N_4242);
and U8445 (N_8445,N_2042,N_2443);
or U8446 (N_8446,N_125,N_1125);
and U8447 (N_8447,N_2210,N_4647);
nand U8448 (N_8448,N_942,N_3527);
and U8449 (N_8449,N_4930,N_3671);
and U8450 (N_8450,N_3907,N_1308);
and U8451 (N_8451,N_2867,N_4342);
or U8452 (N_8452,N_3154,N_1355);
nand U8453 (N_8453,N_4356,N_4084);
nand U8454 (N_8454,N_3724,N_2862);
and U8455 (N_8455,N_1314,N_2733);
and U8456 (N_8456,N_1598,N_111);
nor U8457 (N_8457,N_1370,N_2540);
nor U8458 (N_8458,N_2359,N_2982);
xor U8459 (N_8459,N_925,N_832);
or U8460 (N_8460,N_4058,N_113);
and U8461 (N_8461,N_4509,N_1023);
and U8462 (N_8462,N_1582,N_4393);
nor U8463 (N_8463,N_3631,N_3648);
nor U8464 (N_8464,N_987,N_685);
and U8465 (N_8465,N_1118,N_3769);
nand U8466 (N_8466,N_2321,N_1044);
and U8467 (N_8467,N_3017,N_3983);
nand U8468 (N_8468,N_4121,N_1376);
nor U8469 (N_8469,N_2341,N_3129);
and U8470 (N_8470,N_2173,N_398);
xnor U8471 (N_8471,N_1359,N_2760);
nor U8472 (N_8472,N_456,N_3205);
xnor U8473 (N_8473,N_2383,N_2807);
nand U8474 (N_8474,N_3866,N_4684);
xnor U8475 (N_8475,N_1137,N_382);
or U8476 (N_8476,N_2249,N_2815);
nor U8477 (N_8477,N_4934,N_3404);
nor U8478 (N_8478,N_4857,N_1676);
or U8479 (N_8479,N_4676,N_134);
or U8480 (N_8480,N_905,N_1240);
nand U8481 (N_8481,N_4732,N_716);
nor U8482 (N_8482,N_4269,N_2063);
xnor U8483 (N_8483,N_477,N_3641);
nand U8484 (N_8484,N_4994,N_387);
or U8485 (N_8485,N_1227,N_3669);
nand U8486 (N_8486,N_4019,N_863);
nor U8487 (N_8487,N_2389,N_948);
nand U8488 (N_8488,N_3456,N_4235);
nand U8489 (N_8489,N_2028,N_2634);
or U8490 (N_8490,N_557,N_1298);
and U8491 (N_8491,N_1752,N_2874);
nand U8492 (N_8492,N_1957,N_4139);
nand U8493 (N_8493,N_367,N_96);
nand U8494 (N_8494,N_3805,N_3526);
nand U8495 (N_8495,N_1862,N_3572);
or U8496 (N_8496,N_4812,N_1304);
or U8497 (N_8497,N_1302,N_4486);
or U8498 (N_8498,N_1208,N_2520);
and U8499 (N_8499,N_1688,N_584);
nor U8500 (N_8500,N_1956,N_4431);
nand U8501 (N_8501,N_59,N_1042);
or U8502 (N_8502,N_3216,N_2034);
and U8503 (N_8503,N_3566,N_4370);
or U8504 (N_8504,N_4984,N_2142);
nor U8505 (N_8505,N_3989,N_1791);
nor U8506 (N_8506,N_934,N_2619);
nand U8507 (N_8507,N_19,N_328);
nand U8508 (N_8508,N_842,N_922);
and U8509 (N_8509,N_3967,N_1335);
and U8510 (N_8510,N_30,N_2222);
and U8511 (N_8511,N_1006,N_986);
nand U8512 (N_8512,N_3795,N_1409);
and U8513 (N_8513,N_2067,N_2442);
and U8514 (N_8514,N_3723,N_2117);
and U8515 (N_8515,N_3657,N_4619);
nand U8516 (N_8516,N_2370,N_1033);
or U8517 (N_8517,N_1936,N_1750);
or U8518 (N_8518,N_450,N_3000);
nand U8519 (N_8519,N_1227,N_2996);
or U8520 (N_8520,N_2903,N_1310);
or U8521 (N_8521,N_4382,N_3216);
or U8522 (N_8522,N_1728,N_2677);
nand U8523 (N_8523,N_857,N_4204);
and U8524 (N_8524,N_505,N_4270);
and U8525 (N_8525,N_2272,N_2892);
or U8526 (N_8526,N_1188,N_4697);
and U8527 (N_8527,N_1990,N_2431);
or U8528 (N_8528,N_4092,N_655);
nand U8529 (N_8529,N_2128,N_3026);
nor U8530 (N_8530,N_4982,N_1371);
nand U8531 (N_8531,N_816,N_3261);
nand U8532 (N_8532,N_4717,N_1165);
nor U8533 (N_8533,N_1920,N_660);
nor U8534 (N_8534,N_1202,N_872);
and U8535 (N_8535,N_4391,N_1641);
nor U8536 (N_8536,N_1831,N_2604);
nor U8537 (N_8537,N_4483,N_1431);
and U8538 (N_8538,N_4347,N_598);
and U8539 (N_8539,N_2990,N_4787);
or U8540 (N_8540,N_1235,N_4571);
and U8541 (N_8541,N_2274,N_3914);
nand U8542 (N_8542,N_1993,N_235);
or U8543 (N_8543,N_1331,N_3966);
nand U8544 (N_8544,N_2353,N_1108);
nor U8545 (N_8545,N_4381,N_2056);
nand U8546 (N_8546,N_911,N_3995);
and U8547 (N_8547,N_4068,N_1329);
and U8548 (N_8548,N_1126,N_1524);
nand U8549 (N_8549,N_3652,N_2800);
xnor U8550 (N_8550,N_11,N_3392);
and U8551 (N_8551,N_801,N_3090);
xor U8552 (N_8552,N_1103,N_136);
and U8553 (N_8553,N_3267,N_1761);
or U8554 (N_8554,N_1506,N_3146);
xnor U8555 (N_8555,N_1600,N_1183);
nand U8556 (N_8556,N_2276,N_4345);
nand U8557 (N_8557,N_2222,N_2245);
nand U8558 (N_8558,N_3605,N_2536);
nand U8559 (N_8559,N_2498,N_4404);
or U8560 (N_8560,N_1112,N_751);
nor U8561 (N_8561,N_3344,N_3694);
nand U8562 (N_8562,N_1203,N_2589);
and U8563 (N_8563,N_619,N_4256);
or U8564 (N_8564,N_4861,N_1963);
and U8565 (N_8565,N_1324,N_543);
xor U8566 (N_8566,N_688,N_1734);
and U8567 (N_8567,N_4229,N_4411);
or U8568 (N_8568,N_4204,N_3429);
nor U8569 (N_8569,N_3084,N_824);
xor U8570 (N_8570,N_871,N_3604);
or U8571 (N_8571,N_547,N_3206);
and U8572 (N_8572,N_3180,N_1173);
and U8573 (N_8573,N_2701,N_2453);
and U8574 (N_8574,N_3397,N_807);
xor U8575 (N_8575,N_2652,N_4761);
nand U8576 (N_8576,N_4974,N_879);
nand U8577 (N_8577,N_987,N_1286);
and U8578 (N_8578,N_809,N_542);
and U8579 (N_8579,N_4508,N_1615);
nor U8580 (N_8580,N_1636,N_2587);
nor U8581 (N_8581,N_284,N_3723);
nand U8582 (N_8582,N_3954,N_85);
nand U8583 (N_8583,N_189,N_1519);
or U8584 (N_8584,N_4798,N_2332);
nand U8585 (N_8585,N_889,N_1384);
and U8586 (N_8586,N_1855,N_659);
nand U8587 (N_8587,N_1061,N_4262);
or U8588 (N_8588,N_630,N_1894);
and U8589 (N_8589,N_3401,N_3059);
nor U8590 (N_8590,N_1798,N_3661);
nand U8591 (N_8591,N_2249,N_3170);
nor U8592 (N_8592,N_193,N_4649);
and U8593 (N_8593,N_4662,N_2352);
nor U8594 (N_8594,N_4088,N_282);
xor U8595 (N_8595,N_266,N_2030);
or U8596 (N_8596,N_962,N_1252);
nor U8597 (N_8597,N_3060,N_161);
and U8598 (N_8598,N_2092,N_4226);
nand U8599 (N_8599,N_4738,N_4281);
xnor U8600 (N_8600,N_1239,N_3630);
or U8601 (N_8601,N_3339,N_3790);
and U8602 (N_8602,N_4873,N_774);
and U8603 (N_8603,N_2578,N_2250);
nand U8604 (N_8604,N_3594,N_4508);
nand U8605 (N_8605,N_3971,N_2776);
nand U8606 (N_8606,N_4854,N_2193);
nand U8607 (N_8607,N_1473,N_509);
or U8608 (N_8608,N_4941,N_4662);
xnor U8609 (N_8609,N_2676,N_1086);
nor U8610 (N_8610,N_4174,N_4763);
nand U8611 (N_8611,N_2882,N_1679);
xnor U8612 (N_8612,N_343,N_4267);
xor U8613 (N_8613,N_1429,N_2462);
nand U8614 (N_8614,N_4127,N_4568);
xor U8615 (N_8615,N_1136,N_3858);
and U8616 (N_8616,N_4645,N_1802);
or U8617 (N_8617,N_2482,N_558);
xor U8618 (N_8618,N_49,N_4354);
xor U8619 (N_8619,N_2461,N_3405);
nor U8620 (N_8620,N_794,N_709);
nor U8621 (N_8621,N_2522,N_828);
or U8622 (N_8622,N_2001,N_2571);
and U8623 (N_8623,N_4672,N_4309);
or U8624 (N_8624,N_2134,N_231);
nand U8625 (N_8625,N_1167,N_2278);
and U8626 (N_8626,N_3082,N_2112);
or U8627 (N_8627,N_3804,N_2228);
and U8628 (N_8628,N_962,N_1044);
and U8629 (N_8629,N_569,N_3650);
or U8630 (N_8630,N_2099,N_496);
nand U8631 (N_8631,N_1003,N_3790);
nor U8632 (N_8632,N_4125,N_2681);
and U8633 (N_8633,N_1671,N_1981);
nand U8634 (N_8634,N_89,N_3102);
and U8635 (N_8635,N_1439,N_4069);
or U8636 (N_8636,N_2403,N_3987);
or U8637 (N_8637,N_444,N_4148);
or U8638 (N_8638,N_3707,N_2673);
and U8639 (N_8639,N_3234,N_3201);
or U8640 (N_8640,N_3581,N_2839);
or U8641 (N_8641,N_4232,N_4278);
or U8642 (N_8642,N_282,N_4270);
nand U8643 (N_8643,N_624,N_830);
and U8644 (N_8644,N_1313,N_1412);
xor U8645 (N_8645,N_36,N_312);
or U8646 (N_8646,N_3571,N_2801);
and U8647 (N_8647,N_1022,N_954);
xor U8648 (N_8648,N_4761,N_4191);
and U8649 (N_8649,N_3247,N_759);
nor U8650 (N_8650,N_705,N_166);
nand U8651 (N_8651,N_4976,N_2842);
xor U8652 (N_8652,N_3822,N_2667);
nand U8653 (N_8653,N_4703,N_3889);
or U8654 (N_8654,N_4004,N_2724);
and U8655 (N_8655,N_2459,N_2727);
and U8656 (N_8656,N_4436,N_3825);
and U8657 (N_8657,N_4642,N_3808);
and U8658 (N_8658,N_4230,N_100);
nor U8659 (N_8659,N_2252,N_2727);
and U8660 (N_8660,N_1596,N_3109);
nor U8661 (N_8661,N_4338,N_4018);
nand U8662 (N_8662,N_2967,N_4428);
nand U8663 (N_8663,N_3869,N_4693);
and U8664 (N_8664,N_4604,N_1759);
and U8665 (N_8665,N_1647,N_4054);
and U8666 (N_8666,N_3274,N_3371);
xnor U8667 (N_8667,N_2330,N_4666);
and U8668 (N_8668,N_2249,N_1895);
nor U8669 (N_8669,N_1664,N_3771);
or U8670 (N_8670,N_3270,N_3565);
xnor U8671 (N_8671,N_1826,N_1846);
nor U8672 (N_8672,N_3093,N_2904);
xnor U8673 (N_8673,N_4253,N_2819);
nor U8674 (N_8674,N_2987,N_4995);
nand U8675 (N_8675,N_4717,N_3719);
nor U8676 (N_8676,N_4612,N_3673);
nor U8677 (N_8677,N_1302,N_3652);
nor U8678 (N_8678,N_1219,N_1956);
and U8679 (N_8679,N_3412,N_2335);
nand U8680 (N_8680,N_1679,N_4958);
and U8681 (N_8681,N_649,N_4188);
nand U8682 (N_8682,N_1062,N_2683);
or U8683 (N_8683,N_151,N_2137);
xnor U8684 (N_8684,N_4071,N_3518);
and U8685 (N_8685,N_788,N_2967);
or U8686 (N_8686,N_4416,N_3661);
or U8687 (N_8687,N_81,N_3731);
nand U8688 (N_8688,N_2529,N_1905);
nor U8689 (N_8689,N_2718,N_2906);
nand U8690 (N_8690,N_4149,N_1518);
and U8691 (N_8691,N_4493,N_74);
and U8692 (N_8692,N_4474,N_2746);
xor U8693 (N_8693,N_2864,N_1705);
and U8694 (N_8694,N_1472,N_660);
and U8695 (N_8695,N_4521,N_4735);
nand U8696 (N_8696,N_325,N_2240);
and U8697 (N_8697,N_921,N_3607);
and U8698 (N_8698,N_3340,N_1243);
or U8699 (N_8699,N_1373,N_1152);
or U8700 (N_8700,N_1972,N_3644);
nor U8701 (N_8701,N_4138,N_2193);
xnor U8702 (N_8702,N_4051,N_1436);
nand U8703 (N_8703,N_2937,N_726);
xnor U8704 (N_8704,N_2472,N_3094);
nor U8705 (N_8705,N_3282,N_4620);
or U8706 (N_8706,N_219,N_2450);
nand U8707 (N_8707,N_2287,N_3245);
or U8708 (N_8708,N_879,N_1752);
and U8709 (N_8709,N_2169,N_1064);
and U8710 (N_8710,N_60,N_4384);
xor U8711 (N_8711,N_2126,N_694);
nor U8712 (N_8712,N_3153,N_1073);
nor U8713 (N_8713,N_814,N_446);
nand U8714 (N_8714,N_2561,N_3612);
or U8715 (N_8715,N_4341,N_3371);
and U8716 (N_8716,N_1101,N_1152);
nand U8717 (N_8717,N_3599,N_4695);
and U8718 (N_8718,N_3766,N_3567);
xnor U8719 (N_8719,N_1628,N_4777);
nor U8720 (N_8720,N_836,N_921);
nor U8721 (N_8721,N_101,N_4658);
nand U8722 (N_8722,N_2502,N_3969);
and U8723 (N_8723,N_2425,N_3960);
or U8724 (N_8724,N_1044,N_2621);
xnor U8725 (N_8725,N_2801,N_4703);
or U8726 (N_8726,N_4759,N_3717);
and U8727 (N_8727,N_4244,N_3016);
nand U8728 (N_8728,N_3609,N_4009);
and U8729 (N_8729,N_2270,N_1424);
or U8730 (N_8730,N_4446,N_1060);
nand U8731 (N_8731,N_3618,N_3332);
nand U8732 (N_8732,N_4902,N_3850);
nor U8733 (N_8733,N_3479,N_437);
or U8734 (N_8734,N_227,N_264);
and U8735 (N_8735,N_2508,N_2503);
nand U8736 (N_8736,N_2294,N_711);
and U8737 (N_8737,N_1238,N_3738);
nor U8738 (N_8738,N_614,N_1069);
and U8739 (N_8739,N_4450,N_2844);
nand U8740 (N_8740,N_4946,N_3531);
and U8741 (N_8741,N_2185,N_2843);
nand U8742 (N_8742,N_3501,N_1450);
nand U8743 (N_8743,N_1488,N_514);
and U8744 (N_8744,N_583,N_3111);
or U8745 (N_8745,N_4625,N_3910);
nor U8746 (N_8746,N_1649,N_384);
nand U8747 (N_8747,N_1588,N_650);
and U8748 (N_8748,N_1708,N_920);
xnor U8749 (N_8749,N_1492,N_3743);
nand U8750 (N_8750,N_2629,N_2183);
nand U8751 (N_8751,N_3406,N_35);
nand U8752 (N_8752,N_2792,N_1842);
or U8753 (N_8753,N_2044,N_2877);
and U8754 (N_8754,N_2393,N_2654);
and U8755 (N_8755,N_452,N_3096);
nor U8756 (N_8756,N_3476,N_2926);
nor U8757 (N_8757,N_825,N_418);
nor U8758 (N_8758,N_4577,N_1624);
nor U8759 (N_8759,N_4592,N_3659);
xnor U8760 (N_8760,N_1300,N_4230);
nand U8761 (N_8761,N_3550,N_4028);
nand U8762 (N_8762,N_773,N_1203);
nor U8763 (N_8763,N_4485,N_2023);
and U8764 (N_8764,N_2457,N_2701);
and U8765 (N_8765,N_3201,N_2997);
nand U8766 (N_8766,N_1067,N_4931);
or U8767 (N_8767,N_3014,N_1585);
nor U8768 (N_8768,N_2735,N_1090);
or U8769 (N_8769,N_3697,N_2209);
nand U8770 (N_8770,N_3603,N_1840);
nand U8771 (N_8771,N_169,N_2588);
nand U8772 (N_8772,N_2345,N_2890);
and U8773 (N_8773,N_2111,N_2596);
xor U8774 (N_8774,N_1178,N_723);
and U8775 (N_8775,N_4139,N_2387);
and U8776 (N_8776,N_3238,N_4361);
or U8777 (N_8777,N_1553,N_1284);
nand U8778 (N_8778,N_818,N_1489);
nand U8779 (N_8779,N_3104,N_52);
or U8780 (N_8780,N_2005,N_1530);
or U8781 (N_8781,N_686,N_2292);
and U8782 (N_8782,N_2636,N_2051);
or U8783 (N_8783,N_761,N_4337);
and U8784 (N_8784,N_598,N_4245);
nor U8785 (N_8785,N_1329,N_3948);
or U8786 (N_8786,N_686,N_4921);
nand U8787 (N_8787,N_911,N_268);
xnor U8788 (N_8788,N_3628,N_4351);
nand U8789 (N_8789,N_3271,N_2842);
nor U8790 (N_8790,N_4577,N_50);
or U8791 (N_8791,N_1695,N_4477);
or U8792 (N_8792,N_4590,N_763);
or U8793 (N_8793,N_465,N_3791);
nand U8794 (N_8794,N_54,N_1179);
and U8795 (N_8795,N_3817,N_3897);
xnor U8796 (N_8796,N_1940,N_3333);
or U8797 (N_8797,N_3588,N_1612);
nor U8798 (N_8798,N_2567,N_785);
nand U8799 (N_8799,N_38,N_2031);
nor U8800 (N_8800,N_2077,N_4844);
and U8801 (N_8801,N_3708,N_666);
nand U8802 (N_8802,N_2991,N_589);
nand U8803 (N_8803,N_3141,N_3532);
nand U8804 (N_8804,N_823,N_2863);
or U8805 (N_8805,N_4180,N_4892);
and U8806 (N_8806,N_2082,N_115);
xor U8807 (N_8807,N_924,N_1544);
and U8808 (N_8808,N_2938,N_14);
or U8809 (N_8809,N_184,N_4272);
nor U8810 (N_8810,N_805,N_532);
nor U8811 (N_8811,N_1488,N_3501);
nand U8812 (N_8812,N_783,N_4100);
xnor U8813 (N_8813,N_2620,N_3846);
or U8814 (N_8814,N_816,N_4367);
or U8815 (N_8815,N_4877,N_4482);
nand U8816 (N_8816,N_3314,N_4737);
or U8817 (N_8817,N_4365,N_4726);
xnor U8818 (N_8818,N_1804,N_4664);
and U8819 (N_8819,N_3382,N_808);
nand U8820 (N_8820,N_2036,N_2831);
nor U8821 (N_8821,N_2158,N_4728);
or U8822 (N_8822,N_347,N_910);
and U8823 (N_8823,N_777,N_2916);
or U8824 (N_8824,N_3588,N_1584);
and U8825 (N_8825,N_1688,N_708);
nand U8826 (N_8826,N_4067,N_1270);
and U8827 (N_8827,N_3469,N_438);
nor U8828 (N_8828,N_1567,N_4807);
xor U8829 (N_8829,N_4652,N_2242);
or U8830 (N_8830,N_3834,N_2490);
or U8831 (N_8831,N_4138,N_2667);
or U8832 (N_8832,N_849,N_1090);
nor U8833 (N_8833,N_3250,N_4417);
and U8834 (N_8834,N_3518,N_2268);
or U8835 (N_8835,N_4212,N_2395);
nand U8836 (N_8836,N_3017,N_1409);
nor U8837 (N_8837,N_2124,N_1373);
xor U8838 (N_8838,N_1801,N_2356);
nand U8839 (N_8839,N_527,N_3751);
nand U8840 (N_8840,N_1573,N_372);
or U8841 (N_8841,N_2621,N_3747);
xor U8842 (N_8842,N_3759,N_4898);
or U8843 (N_8843,N_2561,N_649);
and U8844 (N_8844,N_719,N_2681);
nor U8845 (N_8845,N_3962,N_3404);
nor U8846 (N_8846,N_4853,N_2624);
or U8847 (N_8847,N_712,N_1329);
or U8848 (N_8848,N_2739,N_3932);
or U8849 (N_8849,N_2473,N_4312);
and U8850 (N_8850,N_1625,N_24);
xnor U8851 (N_8851,N_2544,N_438);
or U8852 (N_8852,N_1734,N_844);
and U8853 (N_8853,N_3789,N_2227);
xnor U8854 (N_8854,N_2218,N_3227);
nor U8855 (N_8855,N_3120,N_2922);
and U8856 (N_8856,N_2123,N_1669);
nor U8857 (N_8857,N_3554,N_541);
nor U8858 (N_8858,N_1936,N_829);
and U8859 (N_8859,N_2819,N_2741);
nor U8860 (N_8860,N_4232,N_2186);
nand U8861 (N_8861,N_187,N_3982);
or U8862 (N_8862,N_224,N_1409);
nor U8863 (N_8863,N_1434,N_2593);
nor U8864 (N_8864,N_2965,N_2055);
xor U8865 (N_8865,N_994,N_752);
or U8866 (N_8866,N_444,N_26);
nor U8867 (N_8867,N_3329,N_3772);
nor U8868 (N_8868,N_1417,N_680);
nand U8869 (N_8869,N_3370,N_4596);
nor U8870 (N_8870,N_1371,N_564);
nor U8871 (N_8871,N_2818,N_3616);
xnor U8872 (N_8872,N_1255,N_691);
nor U8873 (N_8873,N_3042,N_1164);
nor U8874 (N_8874,N_3824,N_100);
nand U8875 (N_8875,N_2706,N_1909);
and U8876 (N_8876,N_4934,N_703);
or U8877 (N_8877,N_905,N_1434);
nor U8878 (N_8878,N_4855,N_4650);
and U8879 (N_8879,N_4572,N_720);
nor U8880 (N_8880,N_4362,N_512);
and U8881 (N_8881,N_722,N_1159);
and U8882 (N_8882,N_4674,N_2497);
nand U8883 (N_8883,N_3659,N_1336);
and U8884 (N_8884,N_2376,N_1542);
nor U8885 (N_8885,N_2468,N_3876);
or U8886 (N_8886,N_4278,N_433);
and U8887 (N_8887,N_1697,N_4567);
xnor U8888 (N_8888,N_3118,N_2661);
nand U8889 (N_8889,N_4582,N_3971);
nand U8890 (N_8890,N_1300,N_3265);
and U8891 (N_8891,N_2010,N_295);
or U8892 (N_8892,N_3931,N_4052);
nand U8893 (N_8893,N_1094,N_4875);
and U8894 (N_8894,N_4946,N_2901);
nor U8895 (N_8895,N_1909,N_2721);
and U8896 (N_8896,N_1999,N_4114);
nand U8897 (N_8897,N_3405,N_4656);
or U8898 (N_8898,N_4743,N_2779);
nand U8899 (N_8899,N_216,N_188);
nand U8900 (N_8900,N_1109,N_609);
and U8901 (N_8901,N_3010,N_3725);
and U8902 (N_8902,N_2952,N_2758);
or U8903 (N_8903,N_2769,N_2428);
nor U8904 (N_8904,N_2989,N_2475);
or U8905 (N_8905,N_3557,N_1694);
and U8906 (N_8906,N_4297,N_4693);
and U8907 (N_8907,N_2578,N_464);
and U8908 (N_8908,N_1293,N_1925);
or U8909 (N_8909,N_2821,N_1805);
or U8910 (N_8910,N_3569,N_4382);
or U8911 (N_8911,N_1356,N_2574);
nor U8912 (N_8912,N_1571,N_4776);
or U8913 (N_8913,N_746,N_2957);
nand U8914 (N_8914,N_924,N_2502);
nand U8915 (N_8915,N_4936,N_3383);
and U8916 (N_8916,N_3959,N_4152);
or U8917 (N_8917,N_1532,N_4606);
nor U8918 (N_8918,N_2137,N_1707);
and U8919 (N_8919,N_3204,N_3160);
xnor U8920 (N_8920,N_1705,N_1885);
xnor U8921 (N_8921,N_2772,N_1415);
or U8922 (N_8922,N_1508,N_4646);
nor U8923 (N_8923,N_2739,N_4718);
nor U8924 (N_8924,N_653,N_3414);
and U8925 (N_8925,N_2983,N_1631);
or U8926 (N_8926,N_2835,N_4993);
and U8927 (N_8927,N_300,N_718);
nand U8928 (N_8928,N_3545,N_4966);
and U8929 (N_8929,N_2289,N_1585);
or U8930 (N_8930,N_2880,N_4434);
nor U8931 (N_8931,N_3155,N_832);
nand U8932 (N_8932,N_2983,N_2605);
and U8933 (N_8933,N_986,N_4443);
and U8934 (N_8934,N_581,N_1338);
nand U8935 (N_8935,N_721,N_1156);
or U8936 (N_8936,N_3122,N_2531);
and U8937 (N_8937,N_2002,N_2236);
and U8938 (N_8938,N_24,N_3952);
nand U8939 (N_8939,N_1374,N_687);
xnor U8940 (N_8940,N_66,N_380);
or U8941 (N_8941,N_3710,N_4407);
nand U8942 (N_8942,N_247,N_3852);
and U8943 (N_8943,N_189,N_3943);
nand U8944 (N_8944,N_2663,N_4400);
nor U8945 (N_8945,N_3447,N_151);
nand U8946 (N_8946,N_634,N_1604);
nand U8947 (N_8947,N_3360,N_1972);
or U8948 (N_8948,N_562,N_156);
nor U8949 (N_8949,N_2033,N_1567);
nand U8950 (N_8950,N_1374,N_2571);
nand U8951 (N_8951,N_2994,N_2955);
nand U8952 (N_8952,N_3134,N_3019);
and U8953 (N_8953,N_4240,N_2068);
or U8954 (N_8954,N_3928,N_1951);
nand U8955 (N_8955,N_1977,N_3731);
nor U8956 (N_8956,N_1254,N_4852);
nor U8957 (N_8957,N_350,N_1286);
and U8958 (N_8958,N_3146,N_2888);
or U8959 (N_8959,N_1267,N_2532);
or U8960 (N_8960,N_4835,N_487);
and U8961 (N_8961,N_4126,N_824);
xor U8962 (N_8962,N_3218,N_4518);
and U8963 (N_8963,N_2651,N_2766);
nor U8964 (N_8964,N_3017,N_754);
and U8965 (N_8965,N_651,N_44);
and U8966 (N_8966,N_533,N_18);
or U8967 (N_8967,N_4267,N_3410);
and U8968 (N_8968,N_2359,N_1720);
or U8969 (N_8969,N_3392,N_2735);
or U8970 (N_8970,N_4907,N_4524);
nor U8971 (N_8971,N_4323,N_4812);
nand U8972 (N_8972,N_4175,N_1995);
and U8973 (N_8973,N_4957,N_3703);
and U8974 (N_8974,N_2752,N_3589);
nand U8975 (N_8975,N_3341,N_1750);
nor U8976 (N_8976,N_4933,N_4848);
nand U8977 (N_8977,N_2499,N_2172);
nand U8978 (N_8978,N_3957,N_3091);
and U8979 (N_8979,N_250,N_1521);
and U8980 (N_8980,N_3303,N_1353);
nand U8981 (N_8981,N_630,N_1923);
and U8982 (N_8982,N_32,N_1803);
or U8983 (N_8983,N_3442,N_1637);
nand U8984 (N_8984,N_588,N_3442);
nand U8985 (N_8985,N_4301,N_464);
or U8986 (N_8986,N_3144,N_4960);
or U8987 (N_8987,N_3893,N_4840);
nand U8988 (N_8988,N_2567,N_522);
nand U8989 (N_8989,N_883,N_1832);
nor U8990 (N_8990,N_1621,N_3680);
nor U8991 (N_8991,N_3357,N_2576);
nand U8992 (N_8992,N_2816,N_2048);
or U8993 (N_8993,N_4392,N_3054);
nor U8994 (N_8994,N_4725,N_4384);
and U8995 (N_8995,N_1082,N_3785);
nand U8996 (N_8996,N_1714,N_431);
nand U8997 (N_8997,N_1328,N_2354);
nand U8998 (N_8998,N_741,N_1851);
nor U8999 (N_8999,N_37,N_331);
and U9000 (N_9000,N_417,N_3227);
nor U9001 (N_9001,N_2562,N_302);
nor U9002 (N_9002,N_121,N_473);
nor U9003 (N_9003,N_1619,N_4079);
nand U9004 (N_9004,N_1085,N_2699);
nor U9005 (N_9005,N_4752,N_2286);
or U9006 (N_9006,N_4686,N_3011);
nand U9007 (N_9007,N_1708,N_4247);
nand U9008 (N_9008,N_3301,N_3423);
or U9009 (N_9009,N_119,N_4161);
nor U9010 (N_9010,N_3146,N_4419);
nor U9011 (N_9011,N_876,N_1220);
nor U9012 (N_9012,N_1632,N_3126);
or U9013 (N_9013,N_2945,N_3687);
nor U9014 (N_9014,N_4109,N_174);
or U9015 (N_9015,N_1435,N_4847);
and U9016 (N_9016,N_1139,N_777);
or U9017 (N_9017,N_2104,N_707);
and U9018 (N_9018,N_2772,N_2100);
and U9019 (N_9019,N_4655,N_4301);
nand U9020 (N_9020,N_4287,N_4846);
or U9021 (N_9021,N_2338,N_823);
and U9022 (N_9022,N_4095,N_1670);
and U9023 (N_9023,N_3190,N_1714);
and U9024 (N_9024,N_1712,N_4104);
and U9025 (N_9025,N_630,N_1569);
nand U9026 (N_9026,N_486,N_4115);
nor U9027 (N_9027,N_464,N_463);
or U9028 (N_9028,N_4899,N_3862);
nand U9029 (N_9029,N_3263,N_2222);
and U9030 (N_9030,N_4451,N_736);
xnor U9031 (N_9031,N_311,N_2593);
or U9032 (N_9032,N_4348,N_3824);
nor U9033 (N_9033,N_1317,N_672);
or U9034 (N_9034,N_1556,N_1552);
or U9035 (N_9035,N_258,N_3118);
or U9036 (N_9036,N_555,N_4726);
nor U9037 (N_9037,N_2685,N_2608);
xor U9038 (N_9038,N_2173,N_4127);
or U9039 (N_9039,N_553,N_1211);
or U9040 (N_9040,N_3604,N_957);
or U9041 (N_9041,N_3536,N_552);
and U9042 (N_9042,N_2403,N_3145);
or U9043 (N_9043,N_4932,N_3236);
nor U9044 (N_9044,N_1980,N_3202);
or U9045 (N_9045,N_354,N_2396);
nor U9046 (N_9046,N_2992,N_2728);
nand U9047 (N_9047,N_174,N_987);
nor U9048 (N_9048,N_2772,N_1031);
nor U9049 (N_9049,N_4885,N_2230);
and U9050 (N_9050,N_1040,N_2105);
and U9051 (N_9051,N_9,N_871);
nor U9052 (N_9052,N_854,N_2846);
or U9053 (N_9053,N_1644,N_564);
and U9054 (N_9054,N_2224,N_2019);
xor U9055 (N_9055,N_3094,N_4552);
and U9056 (N_9056,N_4706,N_2054);
nand U9057 (N_9057,N_4818,N_1020);
nor U9058 (N_9058,N_4914,N_124);
nor U9059 (N_9059,N_1053,N_495);
and U9060 (N_9060,N_2871,N_4901);
nor U9061 (N_9061,N_3946,N_61);
and U9062 (N_9062,N_721,N_1107);
or U9063 (N_9063,N_4912,N_3755);
and U9064 (N_9064,N_2709,N_2435);
nand U9065 (N_9065,N_1642,N_624);
nor U9066 (N_9066,N_3262,N_3477);
and U9067 (N_9067,N_2381,N_243);
nor U9068 (N_9068,N_2196,N_797);
nor U9069 (N_9069,N_1489,N_2687);
and U9070 (N_9070,N_4304,N_4855);
nand U9071 (N_9071,N_3251,N_2724);
and U9072 (N_9072,N_1043,N_1964);
or U9073 (N_9073,N_2658,N_4984);
nand U9074 (N_9074,N_2483,N_1073);
xor U9075 (N_9075,N_4302,N_1008);
nor U9076 (N_9076,N_3733,N_4315);
nand U9077 (N_9077,N_3957,N_3981);
and U9078 (N_9078,N_735,N_3199);
and U9079 (N_9079,N_4478,N_40);
or U9080 (N_9080,N_770,N_1844);
nand U9081 (N_9081,N_3409,N_3794);
xor U9082 (N_9082,N_1747,N_4743);
xnor U9083 (N_9083,N_2970,N_415);
nand U9084 (N_9084,N_1727,N_2764);
nor U9085 (N_9085,N_2394,N_2495);
nand U9086 (N_9086,N_97,N_2187);
xnor U9087 (N_9087,N_4081,N_4458);
nor U9088 (N_9088,N_4921,N_3717);
nand U9089 (N_9089,N_1457,N_70);
nand U9090 (N_9090,N_1208,N_1772);
nand U9091 (N_9091,N_4625,N_206);
or U9092 (N_9092,N_1534,N_645);
xor U9093 (N_9093,N_1077,N_2682);
nand U9094 (N_9094,N_1128,N_2821);
nand U9095 (N_9095,N_4275,N_4285);
nand U9096 (N_9096,N_4709,N_4192);
xor U9097 (N_9097,N_946,N_3880);
xnor U9098 (N_9098,N_4557,N_325);
nor U9099 (N_9099,N_1420,N_4802);
nand U9100 (N_9100,N_4832,N_2214);
or U9101 (N_9101,N_987,N_2546);
nor U9102 (N_9102,N_3927,N_1251);
or U9103 (N_9103,N_1581,N_975);
nor U9104 (N_9104,N_1886,N_1043);
nand U9105 (N_9105,N_2150,N_4718);
xnor U9106 (N_9106,N_3005,N_2382);
nand U9107 (N_9107,N_4983,N_140);
and U9108 (N_9108,N_3051,N_4230);
and U9109 (N_9109,N_1343,N_4230);
nand U9110 (N_9110,N_1794,N_4099);
and U9111 (N_9111,N_2425,N_3920);
and U9112 (N_9112,N_1859,N_650);
nor U9113 (N_9113,N_2209,N_3730);
xnor U9114 (N_9114,N_4690,N_3211);
nor U9115 (N_9115,N_2964,N_357);
and U9116 (N_9116,N_3362,N_3463);
and U9117 (N_9117,N_3906,N_290);
nand U9118 (N_9118,N_2684,N_2421);
nor U9119 (N_9119,N_1940,N_1007);
nand U9120 (N_9120,N_1442,N_2604);
or U9121 (N_9121,N_4567,N_3220);
nand U9122 (N_9122,N_4910,N_4240);
and U9123 (N_9123,N_1130,N_3294);
or U9124 (N_9124,N_2084,N_1827);
nand U9125 (N_9125,N_3732,N_3253);
nor U9126 (N_9126,N_3701,N_4863);
or U9127 (N_9127,N_805,N_4036);
nand U9128 (N_9128,N_3917,N_849);
nor U9129 (N_9129,N_3951,N_3872);
nor U9130 (N_9130,N_1865,N_1549);
nand U9131 (N_9131,N_3597,N_70);
or U9132 (N_9132,N_2861,N_843);
nor U9133 (N_9133,N_2109,N_2046);
nand U9134 (N_9134,N_1551,N_3753);
or U9135 (N_9135,N_4637,N_2733);
xnor U9136 (N_9136,N_2539,N_2840);
nand U9137 (N_9137,N_646,N_1140);
nor U9138 (N_9138,N_4633,N_246);
and U9139 (N_9139,N_1228,N_2266);
and U9140 (N_9140,N_3045,N_3955);
nand U9141 (N_9141,N_2212,N_1973);
nand U9142 (N_9142,N_3028,N_4428);
or U9143 (N_9143,N_648,N_2129);
or U9144 (N_9144,N_840,N_408);
nand U9145 (N_9145,N_2722,N_924);
or U9146 (N_9146,N_1585,N_4333);
or U9147 (N_9147,N_4579,N_1537);
or U9148 (N_9148,N_1234,N_1755);
and U9149 (N_9149,N_2473,N_1475);
nor U9150 (N_9150,N_4535,N_1825);
or U9151 (N_9151,N_4729,N_3035);
and U9152 (N_9152,N_2395,N_2674);
xnor U9153 (N_9153,N_544,N_1414);
nor U9154 (N_9154,N_3185,N_2770);
nand U9155 (N_9155,N_555,N_245);
nand U9156 (N_9156,N_2281,N_4890);
or U9157 (N_9157,N_3271,N_2466);
nand U9158 (N_9158,N_4009,N_1291);
or U9159 (N_9159,N_14,N_2287);
and U9160 (N_9160,N_738,N_4903);
nor U9161 (N_9161,N_553,N_2511);
nor U9162 (N_9162,N_1340,N_4120);
or U9163 (N_9163,N_1940,N_625);
and U9164 (N_9164,N_1338,N_3086);
nor U9165 (N_9165,N_4838,N_4688);
and U9166 (N_9166,N_3294,N_1684);
and U9167 (N_9167,N_4132,N_1623);
or U9168 (N_9168,N_4618,N_4621);
nand U9169 (N_9169,N_2048,N_1330);
and U9170 (N_9170,N_1,N_3355);
and U9171 (N_9171,N_4215,N_1901);
and U9172 (N_9172,N_4196,N_2425);
nand U9173 (N_9173,N_1302,N_1466);
nand U9174 (N_9174,N_1040,N_4690);
or U9175 (N_9175,N_295,N_2795);
and U9176 (N_9176,N_2974,N_1919);
or U9177 (N_9177,N_976,N_1570);
nand U9178 (N_9178,N_1065,N_3656);
nor U9179 (N_9179,N_2839,N_2455);
nand U9180 (N_9180,N_1027,N_158);
or U9181 (N_9181,N_675,N_2163);
and U9182 (N_9182,N_3969,N_3008);
and U9183 (N_9183,N_547,N_2903);
nor U9184 (N_9184,N_3945,N_3426);
xnor U9185 (N_9185,N_4337,N_441);
or U9186 (N_9186,N_889,N_3880);
nand U9187 (N_9187,N_281,N_1380);
nor U9188 (N_9188,N_594,N_1057);
and U9189 (N_9189,N_2778,N_647);
and U9190 (N_9190,N_3623,N_4981);
xnor U9191 (N_9191,N_1267,N_4468);
or U9192 (N_9192,N_3345,N_1238);
nor U9193 (N_9193,N_1715,N_1322);
nand U9194 (N_9194,N_3526,N_3949);
nor U9195 (N_9195,N_2360,N_2141);
nand U9196 (N_9196,N_2940,N_2835);
and U9197 (N_9197,N_2012,N_3320);
and U9198 (N_9198,N_1465,N_4569);
nor U9199 (N_9199,N_4645,N_4261);
and U9200 (N_9200,N_1505,N_1973);
and U9201 (N_9201,N_1403,N_2682);
or U9202 (N_9202,N_4937,N_4104);
or U9203 (N_9203,N_1344,N_3413);
or U9204 (N_9204,N_1745,N_721);
and U9205 (N_9205,N_1118,N_922);
xnor U9206 (N_9206,N_3285,N_417);
nand U9207 (N_9207,N_2673,N_3939);
nand U9208 (N_9208,N_2284,N_4296);
and U9209 (N_9209,N_1632,N_164);
or U9210 (N_9210,N_2093,N_3005);
nand U9211 (N_9211,N_4197,N_2838);
nand U9212 (N_9212,N_4027,N_893);
nor U9213 (N_9213,N_3908,N_3274);
or U9214 (N_9214,N_3259,N_4386);
or U9215 (N_9215,N_4091,N_3513);
or U9216 (N_9216,N_320,N_1360);
nor U9217 (N_9217,N_403,N_4196);
and U9218 (N_9218,N_3259,N_1173);
nor U9219 (N_9219,N_4578,N_1527);
nand U9220 (N_9220,N_423,N_2953);
nand U9221 (N_9221,N_1545,N_2052);
and U9222 (N_9222,N_2345,N_1262);
nand U9223 (N_9223,N_29,N_2982);
nor U9224 (N_9224,N_2742,N_1778);
nor U9225 (N_9225,N_4419,N_3669);
or U9226 (N_9226,N_1696,N_3423);
and U9227 (N_9227,N_2463,N_4102);
nand U9228 (N_9228,N_3669,N_1675);
nand U9229 (N_9229,N_3578,N_2317);
nand U9230 (N_9230,N_1963,N_2770);
xnor U9231 (N_9231,N_2594,N_2216);
or U9232 (N_9232,N_4670,N_3243);
or U9233 (N_9233,N_4551,N_2869);
nand U9234 (N_9234,N_4462,N_4559);
and U9235 (N_9235,N_3192,N_1156);
nand U9236 (N_9236,N_1378,N_3233);
and U9237 (N_9237,N_168,N_1318);
xor U9238 (N_9238,N_3616,N_3577);
and U9239 (N_9239,N_2028,N_715);
nand U9240 (N_9240,N_4240,N_4660);
nand U9241 (N_9241,N_3377,N_1340);
nand U9242 (N_9242,N_1014,N_2356);
and U9243 (N_9243,N_3814,N_4714);
nor U9244 (N_9244,N_3400,N_414);
xor U9245 (N_9245,N_2217,N_4177);
and U9246 (N_9246,N_4263,N_208);
or U9247 (N_9247,N_2426,N_1911);
and U9248 (N_9248,N_4369,N_1961);
nand U9249 (N_9249,N_1186,N_3075);
nor U9250 (N_9250,N_525,N_259);
or U9251 (N_9251,N_821,N_3314);
and U9252 (N_9252,N_3928,N_4782);
nor U9253 (N_9253,N_2545,N_599);
and U9254 (N_9254,N_4268,N_1830);
and U9255 (N_9255,N_3508,N_4691);
nand U9256 (N_9256,N_330,N_2026);
nand U9257 (N_9257,N_4282,N_713);
nand U9258 (N_9258,N_2895,N_637);
xnor U9259 (N_9259,N_4228,N_3555);
xnor U9260 (N_9260,N_38,N_1564);
nand U9261 (N_9261,N_502,N_817);
and U9262 (N_9262,N_4799,N_1534);
and U9263 (N_9263,N_3721,N_2326);
nor U9264 (N_9264,N_1350,N_1899);
nor U9265 (N_9265,N_2266,N_1942);
nand U9266 (N_9266,N_421,N_2061);
nor U9267 (N_9267,N_407,N_4009);
nor U9268 (N_9268,N_148,N_4930);
nand U9269 (N_9269,N_3315,N_1482);
nor U9270 (N_9270,N_2039,N_3848);
xor U9271 (N_9271,N_2948,N_2746);
and U9272 (N_9272,N_1,N_614);
xor U9273 (N_9273,N_2913,N_3570);
and U9274 (N_9274,N_1786,N_3356);
nor U9275 (N_9275,N_2536,N_2999);
nor U9276 (N_9276,N_4380,N_3715);
or U9277 (N_9277,N_3359,N_2591);
or U9278 (N_9278,N_4888,N_151);
nor U9279 (N_9279,N_4183,N_2308);
and U9280 (N_9280,N_631,N_2324);
or U9281 (N_9281,N_700,N_2764);
and U9282 (N_9282,N_3923,N_398);
nor U9283 (N_9283,N_4770,N_2623);
nand U9284 (N_9284,N_3510,N_3144);
or U9285 (N_9285,N_607,N_496);
or U9286 (N_9286,N_4564,N_3961);
or U9287 (N_9287,N_1491,N_4779);
and U9288 (N_9288,N_1433,N_2001);
or U9289 (N_9289,N_2177,N_3085);
xnor U9290 (N_9290,N_3666,N_4750);
nand U9291 (N_9291,N_878,N_4959);
or U9292 (N_9292,N_442,N_2933);
nand U9293 (N_9293,N_3542,N_2732);
and U9294 (N_9294,N_142,N_4008);
and U9295 (N_9295,N_608,N_3686);
or U9296 (N_9296,N_967,N_2542);
and U9297 (N_9297,N_130,N_3675);
or U9298 (N_9298,N_1906,N_195);
and U9299 (N_9299,N_2914,N_1138);
nand U9300 (N_9300,N_1629,N_500);
or U9301 (N_9301,N_2282,N_4237);
and U9302 (N_9302,N_1489,N_1174);
or U9303 (N_9303,N_1314,N_3229);
or U9304 (N_9304,N_4128,N_1195);
and U9305 (N_9305,N_1779,N_2362);
or U9306 (N_9306,N_3188,N_1953);
and U9307 (N_9307,N_2474,N_4259);
and U9308 (N_9308,N_2352,N_1159);
or U9309 (N_9309,N_4615,N_4926);
and U9310 (N_9310,N_1071,N_4395);
or U9311 (N_9311,N_1208,N_1743);
or U9312 (N_9312,N_1058,N_3547);
or U9313 (N_9313,N_729,N_3317);
nor U9314 (N_9314,N_2195,N_3990);
and U9315 (N_9315,N_3354,N_619);
xnor U9316 (N_9316,N_1006,N_2265);
xnor U9317 (N_9317,N_4975,N_1495);
nand U9318 (N_9318,N_1937,N_1418);
and U9319 (N_9319,N_3939,N_4103);
or U9320 (N_9320,N_1554,N_2951);
and U9321 (N_9321,N_4395,N_3574);
xnor U9322 (N_9322,N_4218,N_3511);
nor U9323 (N_9323,N_73,N_3213);
and U9324 (N_9324,N_2464,N_4409);
or U9325 (N_9325,N_61,N_747);
nand U9326 (N_9326,N_10,N_2369);
nor U9327 (N_9327,N_799,N_2023);
xnor U9328 (N_9328,N_4155,N_2512);
and U9329 (N_9329,N_1612,N_368);
xor U9330 (N_9330,N_2116,N_3625);
nand U9331 (N_9331,N_38,N_3683);
nand U9332 (N_9332,N_2531,N_1112);
or U9333 (N_9333,N_837,N_3596);
or U9334 (N_9334,N_3438,N_1222);
or U9335 (N_9335,N_4453,N_4783);
nand U9336 (N_9336,N_890,N_3938);
nand U9337 (N_9337,N_1706,N_4927);
or U9338 (N_9338,N_207,N_657);
nor U9339 (N_9339,N_3952,N_485);
nor U9340 (N_9340,N_1176,N_2400);
nor U9341 (N_9341,N_1219,N_2083);
and U9342 (N_9342,N_3202,N_2914);
and U9343 (N_9343,N_3951,N_177);
nor U9344 (N_9344,N_1466,N_372);
nand U9345 (N_9345,N_4150,N_41);
nand U9346 (N_9346,N_1870,N_303);
nand U9347 (N_9347,N_2634,N_4325);
nand U9348 (N_9348,N_3178,N_4627);
nand U9349 (N_9349,N_964,N_503);
and U9350 (N_9350,N_2583,N_1628);
and U9351 (N_9351,N_4218,N_3356);
or U9352 (N_9352,N_1928,N_4109);
xnor U9353 (N_9353,N_4545,N_4351);
or U9354 (N_9354,N_672,N_4323);
nor U9355 (N_9355,N_1531,N_1803);
and U9356 (N_9356,N_4291,N_3141);
or U9357 (N_9357,N_4869,N_4561);
xor U9358 (N_9358,N_3897,N_790);
nor U9359 (N_9359,N_3427,N_1279);
or U9360 (N_9360,N_4098,N_911);
and U9361 (N_9361,N_4622,N_3565);
nand U9362 (N_9362,N_3935,N_4766);
nand U9363 (N_9363,N_2456,N_1727);
nor U9364 (N_9364,N_928,N_3923);
nand U9365 (N_9365,N_3249,N_4251);
or U9366 (N_9366,N_3953,N_1502);
and U9367 (N_9367,N_1160,N_4957);
nor U9368 (N_9368,N_366,N_4609);
nor U9369 (N_9369,N_2244,N_2264);
or U9370 (N_9370,N_2816,N_299);
xor U9371 (N_9371,N_738,N_4434);
xor U9372 (N_9372,N_416,N_319);
or U9373 (N_9373,N_2850,N_4695);
nor U9374 (N_9374,N_2879,N_397);
xor U9375 (N_9375,N_3057,N_2254);
nand U9376 (N_9376,N_3041,N_1507);
nor U9377 (N_9377,N_4641,N_1423);
nor U9378 (N_9378,N_1235,N_2606);
or U9379 (N_9379,N_1325,N_612);
or U9380 (N_9380,N_1818,N_117);
nand U9381 (N_9381,N_465,N_3000);
and U9382 (N_9382,N_171,N_4239);
nor U9383 (N_9383,N_2437,N_2377);
xnor U9384 (N_9384,N_38,N_2619);
and U9385 (N_9385,N_1673,N_1859);
nand U9386 (N_9386,N_4866,N_3660);
and U9387 (N_9387,N_1132,N_1248);
nor U9388 (N_9388,N_490,N_2215);
nand U9389 (N_9389,N_4344,N_3177);
nand U9390 (N_9390,N_3839,N_1046);
and U9391 (N_9391,N_373,N_4659);
or U9392 (N_9392,N_1457,N_3981);
nor U9393 (N_9393,N_1732,N_2569);
xnor U9394 (N_9394,N_2720,N_2115);
or U9395 (N_9395,N_424,N_4352);
nor U9396 (N_9396,N_97,N_2298);
and U9397 (N_9397,N_1117,N_1219);
or U9398 (N_9398,N_4763,N_4014);
and U9399 (N_9399,N_3266,N_3558);
nand U9400 (N_9400,N_3791,N_4868);
nor U9401 (N_9401,N_2701,N_1833);
xor U9402 (N_9402,N_1213,N_1821);
nand U9403 (N_9403,N_4050,N_3869);
nand U9404 (N_9404,N_3317,N_388);
nor U9405 (N_9405,N_1443,N_1409);
nand U9406 (N_9406,N_48,N_166);
nand U9407 (N_9407,N_4378,N_4851);
or U9408 (N_9408,N_1522,N_1867);
nor U9409 (N_9409,N_3395,N_2418);
nand U9410 (N_9410,N_1974,N_451);
nor U9411 (N_9411,N_2951,N_14);
or U9412 (N_9412,N_2151,N_4303);
and U9413 (N_9413,N_4561,N_2475);
and U9414 (N_9414,N_2307,N_1095);
nor U9415 (N_9415,N_3512,N_2813);
nand U9416 (N_9416,N_2919,N_4474);
xor U9417 (N_9417,N_2069,N_2594);
and U9418 (N_9418,N_1632,N_1335);
nor U9419 (N_9419,N_4938,N_1161);
nand U9420 (N_9420,N_686,N_1077);
nand U9421 (N_9421,N_4456,N_506);
and U9422 (N_9422,N_1285,N_1746);
and U9423 (N_9423,N_2072,N_1521);
nand U9424 (N_9424,N_1083,N_4471);
or U9425 (N_9425,N_3204,N_1565);
nand U9426 (N_9426,N_2369,N_1080);
xnor U9427 (N_9427,N_4468,N_2407);
nand U9428 (N_9428,N_1056,N_2339);
nor U9429 (N_9429,N_3712,N_4483);
or U9430 (N_9430,N_3175,N_4159);
and U9431 (N_9431,N_2298,N_3255);
and U9432 (N_9432,N_3885,N_156);
nand U9433 (N_9433,N_3034,N_820);
xor U9434 (N_9434,N_3691,N_1482);
or U9435 (N_9435,N_4093,N_127);
nand U9436 (N_9436,N_1929,N_1870);
and U9437 (N_9437,N_3837,N_1716);
or U9438 (N_9438,N_305,N_995);
nand U9439 (N_9439,N_204,N_4279);
or U9440 (N_9440,N_4005,N_4605);
nand U9441 (N_9441,N_184,N_3932);
and U9442 (N_9442,N_144,N_4862);
and U9443 (N_9443,N_2004,N_1292);
nand U9444 (N_9444,N_3097,N_3073);
or U9445 (N_9445,N_939,N_586);
xor U9446 (N_9446,N_1953,N_81);
xnor U9447 (N_9447,N_1758,N_2236);
or U9448 (N_9448,N_3705,N_1133);
and U9449 (N_9449,N_3541,N_1729);
nor U9450 (N_9450,N_668,N_724);
and U9451 (N_9451,N_667,N_3547);
nand U9452 (N_9452,N_4827,N_3630);
nand U9453 (N_9453,N_2803,N_574);
nor U9454 (N_9454,N_312,N_2789);
nand U9455 (N_9455,N_4326,N_4124);
nor U9456 (N_9456,N_444,N_531);
nor U9457 (N_9457,N_159,N_3276);
and U9458 (N_9458,N_2740,N_2169);
and U9459 (N_9459,N_1116,N_1568);
nand U9460 (N_9460,N_3376,N_3776);
nor U9461 (N_9461,N_4682,N_3612);
or U9462 (N_9462,N_4012,N_956);
nor U9463 (N_9463,N_2090,N_186);
nor U9464 (N_9464,N_3002,N_4270);
nor U9465 (N_9465,N_2571,N_2060);
and U9466 (N_9466,N_3679,N_1837);
or U9467 (N_9467,N_1827,N_864);
nor U9468 (N_9468,N_4609,N_3292);
nor U9469 (N_9469,N_4256,N_4808);
nor U9470 (N_9470,N_3304,N_4087);
and U9471 (N_9471,N_4219,N_4628);
nor U9472 (N_9472,N_1378,N_3213);
nor U9473 (N_9473,N_2173,N_3096);
or U9474 (N_9474,N_4750,N_4237);
nor U9475 (N_9475,N_1684,N_586);
and U9476 (N_9476,N_1954,N_4271);
and U9477 (N_9477,N_368,N_1864);
nand U9478 (N_9478,N_2482,N_4972);
or U9479 (N_9479,N_2578,N_1180);
nor U9480 (N_9480,N_155,N_4862);
and U9481 (N_9481,N_4385,N_3905);
nand U9482 (N_9482,N_4749,N_1680);
or U9483 (N_9483,N_2581,N_4363);
nor U9484 (N_9484,N_879,N_4209);
or U9485 (N_9485,N_1419,N_3879);
nand U9486 (N_9486,N_3328,N_494);
nor U9487 (N_9487,N_4209,N_2842);
and U9488 (N_9488,N_2927,N_719);
nor U9489 (N_9489,N_3921,N_4908);
nand U9490 (N_9490,N_4476,N_4201);
and U9491 (N_9491,N_3617,N_4247);
or U9492 (N_9492,N_1064,N_1981);
nor U9493 (N_9493,N_1782,N_2864);
xor U9494 (N_9494,N_630,N_1248);
nor U9495 (N_9495,N_1610,N_3820);
xnor U9496 (N_9496,N_2601,N_1960);
and U9497 (N_9497,N_1259,N_91);
nor U9498 (N_9498,N_1475,N_4708);
and U9499 (N_9499,N_3459,N_3778);
and U9500 (N_9500,N_2342,N_715);
nor U9501 (N_9501,N_4974,N_4184);
or U9502 (N_9502,N_2499,N_2856);
and U9503 (N_9503,N_1665,N_1154);
and U9504 (N_9504,N_4428,N_7);
or U9505 (N_9505,N_558,N_3710);
or U9506 (N_9506,N_691,N_3203);
nor U9507 (N_9507,N_3855,N_3040);
or U9508 (N_9508,N_2270,N_3567);
and U9509 (N_9509,N_3391,N_4992);
or U9510 (N_9510,N_1440,N_325);
or U9511 (N_9511,N_1868,N_1617);
nor U9512 (N_9512,N_1215,N_2675);
nand U9513 (N_9513,N_3470,N_4820);
nand U9514 (N_9514,N_547,N_726);
nand U9515 (N_9515,N_2968,N_3815);
and U9516 (N_9516,N_3241,N_2172);
or U9517 (N_9517,N_3747,N_1364);
xnor U9518 (N_9518,N_2655,N_1059);
and U9519 (N_9519,N_3989,N_2527);
or U9520 (N_9520,N_1078,N_3773);
nor U9521 (N_9521,N_2785,N_2572);
and U9522 (N_9522,N_1488,N_4552);
or U9523 (N_9523,N_4112,N_1185);
nand U9524 (N_9524,N_1201,N_990);
nor U9525 (N_9525,N_3549,N_1026);
nor U9526 (N_9526,N_2166,N_4750);
nand U9527 (N_9527,N_2071,N_3499);
xnor U9528 (N_9528,N_3179,N_1128);
nand U9529 (N_9529,N_2933,N_2941);
and U9530 (N_9530,N_4977,N_429);
nor U9531 (N_9531,N_3736,N_1812);
xnor U9532 (N_9532,N_3444,N_309);
and U9533 (N_9533,N_1318,N_567);
nor U9534 (N_9534,N_1082,N_727);
nand U9535 (N_9535,N_1577,N_2086);
nand U9536 (N_9536,N_3791,N_2705);
nor U9537 (N_9537,N_2358,N_3413);
or U9538 (N_9538,N_4921,N_4649);
xnor U9539 (N_9539,N_2145,N_2778);
nor U9540 (N_9540,N_4786,N_4236);
nand U9541 (N_9541,N_1248,N_821);
and U9542 (N_9542,N_3088,N_703);
or U9543 (N_9543,N_2066,N_3858);
nor U9544 (N_9544,N_2667,N_1708);
nor U9545 (N_9545,N_1787,N_3087);
and U9546 (N_9546,N_437,N_4425);
nor U9547 (N_9547,N_2799,N_2121);
and U9548 (N_9548,N_3664,N_2700);
nand U9549 (N_9549,N_4702,N_836);
xnor U9550 (N_9550,N_1372,N_2377);
nand U9551 (N_9551,N_2937,N_3221);
nand U9552 (N_9552,N_2605,N_2862);
and U9553 (N_9553,N_1717,N_1121);
and U9554 (N_9554,N_2878,N_3798);
or U9555 (N_9555,N_2917,N_2986);
and U9556 (N_9556,N_1478,N_3759);
nand U9557 (N_9557,N_1296,N_1714);
nand U9558 (N_9558,N_1857,N_4566);
nor U9559 (N_9559,N_2057,N_255);
or U9560 (N_9560,N_4753,N_1563);
nand U9561 (N_9561,N_4300,N_2207);
nor U9562 (N_9562,N_884,N_1704);
or U9563 (N_9563,N_1430,N_3315);
xor U9564 (N_9564,N_934,N_4756);
nor U9565 (N_9565,N_2931,N_3437);
nor U9566 (N_9566,N_3559,N_3796);
or U9567 (N_9567,N_2024,N_3872);
nor U9568 (N_9568,N_2461,N_2617);
or U9569 (N_9569,N_2848,N_3592);
nor U9570 (N_9570,N_4852,N_913);
and U9571 (N_9571,N_1937,N_1344);
nor U9572 (N_9572,N_3208,N_4694);
nor U9573 (N_9573,N_2061,N_209);
nand U9574 (N_9574,N_2575,N_3569);
or U9575 (N_9575,N_140,N_1324);
nor U9576 (N_9576,N_2351,N_2985);
nand U9577 (N_9577,N_1341,N_3275);
nand U9578 (N_9578,N_4614,N_167);
or U9579 (N_9579,N_3053,N_4792);
nor U9580 (N_9580,N_1475,N_644);
nor U9581 (N_9581,N_2931,N_3919);
nor U9582 (N_9582,N_3722,N_4360);
nor U9583 (N_9583,N_2441,N_938);
or U9584 (N_9584,N_450,N_1741);
nor U9585 (N_9585,N_2031,N_835);
nand U9586 (N_9586,N_3485,N_4605);
or U9587 (N_9587,N_4583,N_1087);
xnor U9588 (N_9588,N_1022,N_4476);
nor U9589 (N_9589,N_1881,N_4430);
nor U9590 (N_9590,N_4569,N_3018);
nand U9591 (N_9591,N_4045,N_1485);
and U9592 (N_9592,N_1807,N_1145);
xor U9593 (N_9593,N_17,N_2986);
nand U9594 (N_9594,N_2193,N_4464);
nand U9595 (N_9595,N_2044,N_2538);
nor U9596 (N_9596,N_3133,N_989);
and U9597 (N_9597,N_783,N_4761);
and U9598 (N_9598,N_3196,N_3213);
and U9599 (N_9599,N_3716,N_2329);
and U9600 (N_9600,N_143,N_1295);
or U9601 (N_9601,N_2082,N_3839);
and U9602 (N_9602,N_235,N_3865);
or U9603 (N_9603,N_4472,N_4431);
and U9604 (N_9604,N_1236,N_1865);
nand U9605 (N_9605,N_3094,N_4295);
or U9606 (N_9606,N_206,N_30);
and U9607 (N_9607,N_3975,N_928);
nand U9608 (N_9608,N_468,N_3318);
or U9609 (N_9609,N_792,N_2123);
nor U9610 (N_9610,N_983,N_81);
nor U9611 (N_9611,N_1811,N_598);
or U9612 (N_9612,N_4193,N_1839);
or U9613 (N_9613,N_3566,N_4604);
nand U9614 (N_9614,N_4653,N_3216);
nand U9615 (N_9615,N_1907,N_2152);
nand U9616 (N_9616,N_1937,N_4362);
nand U9617 (N_9617,N_683,N_1615);
nand U9618 (N_9618,N_4930,N_4644);
and U9619 (N_9619,N_1670,N_987);
or U9620 (N_9620,N_3386,N_729);
nand U9621 (N_9621,N_4049,N_3312);
nor U9622 (N_9622,N_424,N_4170);
and U9623 (N_9623,N_926,N_1761);
or U9624 (N_9624,N_3045,N_2672);
xor U9625 (N_9625,N_3278,N_3376);
nand U9626 (N_9626,N_4020,N_2765);
nor U9627 (N_9627,N_943,N_1978);
or U9628 (N_9628,N_3132,N_4897);
nor U9629 (N_9629,N_3137,N_1136);
xnor U9630 (N_9630,N_1368,N_2107);
nand U9631 (N_9631,N_1247,N_2476);
and U9632 (N_9632,N_3778,N_2214);
xor U9633 (N_9633,N_1908,N_2892);
nand U9634 (N_9634,N_344,N_2073);
and U9635 (N_9635,N_2607,N_3786);
nand U9636 (N_9636,N_119,N_4450);
or U9637 (N_9637,N_4187,N_3143);
nor U9638 (N_9638,N_1752,N_3776);
or U9639 (N_9639,N_143,N_3675);
or U9640 (N_9640,N_4272,N_1933);
nor U9641 (N_9641,N_1752,N_544);
nor U9642 (N_9642,N_4836,N_1087);
or U9643 (N_9643,N_4523,N_4667);
xor U9644 (N_9644,N_3504,N_3062);
nand U9645 (N_9645,N_2990,N_1568);
nand U9646 (N_9646,N_4826,N_2772);
nand U9647 (N_9647,N_1307,N_2545);
or U9648 (N_9648,N_4305,N_4965);
or U9649 (N_9649,N_3876,N_3480);
nand U9650 (N_9650,N_2964,N_1257);
nor U9651 (N_9651,N_1521,N_2918);
nand U9652 (N_9652,N_3464,N_4725);
and U9653 (N_9653,N_468,N_1610);
and U9654 (N_9654,N_3037,N_637);
nor U9655 (N_9655,N_900,N_27);
nand U9656 (N_9656,N_1762,N_4188);
or U9657 (N_9657,N_316,N_999);
and U9658 (N_9658,N_259,N_150);
nand U9659 (N_9659,N_1958,N_2366);
nor U9660 (N_9660,N_706,N_3156);
nand U9661 (N_9661,N_2480,N_2074);
nor U9662 (N_9662,N_2233,N_2275);
nor U9663 (N_9663,N_3344,N_4135);
or U9664 (N_9664,N_2842,N_4060);
nor U9665 (N_9665,N_1271,N_3399);
xnor U9666 (N_9666,N_1594,N_4000);
nand U9667 (N_9667,N_2614,N_1181);
nor U9668 (N_9668,N_2668,N_364);
xnor U9669 (N_9669,N_4994,N_3744);
nand U9670 (N_9670,N_1104,N_2264);
nand U9671 (N_9671,N_812,N_1904);
and U9672 (N_9672,N_3945,N_3745);
and U9673 (N_9673,N_3227,N_2649);
nand U9674 (N_9674,N_2504,N_29);
nand U9675 (N_9675,N_3079,N_1383);
or U9676 (N_9676,N_4327,N_794);
and U9677 (N_9677,N_503,N_934);
nor U9678 (N_9678,N_4957,N_3450);
and U9679 (N_9679,N_1479,N_425);
nand U9680 (N_9680,N_4189,N_3494);
or U9681 (N_9681,N_1278,N_1340);
nor U9682 (N_9682,N_2499,N_4082);
xnor U9683 (N_9683,N_3939,N_4661);
or U9684 (N_9684,N_2279,N_2691);
or U9685 (N_9685,N_378,N_4138);
nand U9686 (N_9686,N_682,N_3397);
nor U9687 (N_9687,N_3832,N_552);
nor U9688 (N_9688,N_1620,N_807);
or U9689 (N_9689,N_1873,N_3608);
or U9690 (N_9690,N_809,N_4664);
nand U9691 (N_9691,N_4495,N_2322);
nand U9692 (N_9692,N_177,N_3114);
xor U9693 (N_9693,N_502,N_2845);
nor U9694 (N_9694,N_2321,N_323);
xor U9695 (N_9695,N_4881,N_1435);
nor U9696 (N_9696,N_3650,N_3050);
and U9697 (N_9697,N_2425,N_1868);
nand U9698 (N_9698,N_863,N_1936);
and U9699 (N_9699,N_1666,N_2695);
nor U9700 (N_9700,N_286,N_1552);
xnor U9701 (N_9701,N_4777,N_1858);
or U9702 (N_9702,N_1696,N_4673);
xor U9703 (N_9703,N_4835,N_3104);
nor U9704 (N_9704,N_3576,N_2073);
nand U9705 (N_9705,N_72,N_1841);
xnor U9706 (N_9706,N_4141,N_4473);
or U9707 (N_9707,N_2650,N_4022);
nand U9708 (N_9708,N_1870,N_955);
nor U9709 (N_9709,N_439,N_2322);
and U9710 (N_9710,N_4826,N_3750);
nor U9711 (N_9711,N_2712,N_3467);
and U9712 (N_9712,N_639,N_1593);
or U9713 (N_9713,N_1707,N_1048);
nor U9714 (N_9714,N_3050,N_4569);
nor U9715 (N_9715,N_174,N_3227);
or U9716 (N_9716,N_256,N_2862);
nor U9717 (N_9717,N_1483,N_3243);
nor U9718 (N_9718,N_2936,N_3468);
nor U9719 (N_9719,N_4175,N_1513);
nand U9720 (N_9720,N_96,N_312);
xnor U9721 (N_9721,N_279,N_216);
or U9722 (N_9722,N_1545,N_4826);
nand U9723 (N_9723,N_238,N_580);
or U9724 (N_9724,N_195,N_3577);
nor U9725 (N_9725,N_265,N_2876);
or U9726 (N_9726,N_287,N_684);
nor U9727 (N_9727,N_4682,N_2900);
xor U9728 (N_9728,N_3370,N_55);
and U9729 (N_9729,N_4284,N_2984);
or U9730 (N_9730,N_2012,N_4214);
nor U9731 (N_9731,N_3912,N_955);
xnor U9732 (N_9732,N_3066,N_561);
and U9733 (N_9733,N_2441,N_4604);
nor U9734 (N_9734,N_2319,N_997);
nand U9735 (N_9735,N_2651,N_372);
nor U9736 (N_9736,N_3726,N_511);
nor U9737 (N_9737,N_4594,N_4260);
nor U9738 (N_9738,N_2236,N_4096);
nor U9739 (N_9739,N_1234,N_3801);
nor U9740 (N_9740,N_2302,N_542);
nand U9741 (N_9741,N_4009,N_2826);
nor U9742 (N_9742,N_4035,N_1092);
xor U9743 (N_9743,N_2383,N_4293);
nand U9744 (N_9744,N_382,N_845);
nor U9745 (N_9745,N_2213,N_2984);
nand U9746 (N_9746,N_4439,N_84);
and U9747 (N_9747,N_3246,N_1539);
and U9748 (N_9748,N_104,N_4165);
xor U9749 (N_9749,N_1101,N_4784);
nand U9750 (N_9750,N_860,N_4704);
or U9751 (N_9751,N_1873,N_917);
and U9752 (N_9752,N_3479,N_2476);
nor U9753 (N_9753,N_636,N_2679);
nor U9754 (N_9754,N_3312,N_608);
nand U9755 (N_9755,N_1925,N_2957);
xor U9756 (N_9756,N_1911,N_4070);
or U9757 (N_9757,N_4397,N_2986);
or U9758 (N_9758,N_93,N_4719);
or U9759 (N_9759,N_1853,N_3419);
or U9760 (N_9760,N_1790,N_441);
and U9761 (N_9761,N_4714,N_4765);
nand U9762 (N_9762,N_82,N_971);
and U9763 (N_9763,N_1690,N_4819);
nand U9764 (N_9764,N_746,N_2058);
and U9765 (N_9765,N_4423,N_4535);
nor U9766 (N_9766,N_3086,N_636);
nand U9767 (N_9767,N_1887,N_3935);
and U9768 (N_9768,N_4892,N_410);
nand U9769 (N_9769,N_2249,N_970);
and U9770 (N_9770,N_4033,N_1666);
and U9771 (N_9771,N_4131,N_4788);
nor U9772 (N_9772,N_4856,N_3228);
and U9773 (N_9773,N_1086,N_1319);
nor U9774 (N_9774,N_1451,N_2385);
or U9775 (N_9775,N_3543,N_1407);
nand U9776 (N_9776,N_3109,N_352);
xor U9777 (N_9777,N_3915,N_697);
nand U9778 (N_9778,N_2831,N_4430);
and U9779 (N_9779,N_4371,N_2758);
and U9780 (N_9780,N_2063,N_4177);
and U9781 (N_9781,N_3243,N_4474);
and U9782 (N_9782,N_1790,N_3874);
nor U9783 (N_9783,N_3067,N_3387);
or U9784 (N_9784,N_3270,N_3079);
and U9785 (N_9785,N_3297,N_2554);
or U9786 (N_9786,N_232,N_1391);
and U9787 (N_9787,N_3925,N_4281);
and U9788 (N_9788,N_4047,N_1875);
xnor U9789 (N_9789,N_619,N_2098);
nand U9790 (N_9790,N_1464,N_4533);
or U9791 (N_9791,N_2068,N_723);
xor U9792 (N_9792,N_4174,N_2026);
nand U9793 (N_9793,N_3954,N_3178);
and U9794 (N_9794,N_3296,N_1472);
xnor U9795 (N_9795,N_4816,N_4891);
nand U9796 (N_9796,N_1782,N_1335);
nand U9797 (N_9797,N_174,N_805);
and U9798 (N_9798,N_2850,N_3201);
nand U9799 (N_9799,N_1677,N_3415);
or U9800 (N_9800,N_2130,N_3387);
nor U9801 (N_9801,N_1483,N_1735);
nor U9802 (N_9802,N_2430,N_2455);
nand U9803 (N_9803,N_4782,N_1996);
and U9804 (N_9804,N_1820,N_2451);
or U9805 (N_9805,N_3142,N_2215);
nand U9806 (N_9806,N_4260,N_2947);
or U9807 (N_9807,N_3087,N_4950);
and U9808 (N_9808,N_1429,N_2843);
nor U9809 (N_9809,N_1055,N_525);
nor U9810 (N_9810,N_3210,N_2933);
xnor U9811 (N_9811,N_2752,N_2289);
nor U9812 (N_9812,N_2299,N_4164);
nand U9813 (N_9813,N_2090,N_1236);
and U9814 (N_9814,N_1608,N_4981);
or U9815 (N_9815,N_1704,N_1446);
nand U9816 (N_9816,N_4551,N_4734);
or U9817 (N_9817,N_830,N_2876);
nand U9818 (N_9818,N_2581,N_2228);
nand U9819 (N_9819,N_4837,N_768);
xor U9820 (N_9820,N_4184,N_4427);
or U9821 (N_9821,N_4083,N_3772);
nor U9822 (N_9822,N_3356,N_921);
nand U9823 (N_9823,N_1395,N_180);
nand U9824 (N_9824,N_1115,N_1781);
or U9825 (N_9825,N_2761,N_2961);
nor U9826 (N_9826,N_3443,N_982);
or U9827 (N_9827,N_3137,N_3654);
and U9828 (N_9828,N_1245,N_3643);
nor U9829 (N_9829,N_2602,N_3134);
and U9830 (N_9830,N_478,N_1154);
xor U9831 (N_9831,N_1926,N_3102);
and U9832 (N_9832,N_811,N_2500);
and U9833 (N_9833,N_1358,N_2306);
and U9834 (N_9834,N_1051,N_1415);
nand U9835 (N_9835,N_3517,N_3354);
and U9836 (N_9836,N_964,N_3355);
or U9837 (N_9837,N_4571,N_4474);
or U9838 (N_9838,N_4563,N_220);
and U9839 (N_9839,N_1637,N_3025);
or U9840 (N_9840,N_3281,N_621);
xnor U9841 (N_9841,N_1276,N_3621);
nand U9842 (N_9842,N_4753,N_4007);
xnor U9843 (N_9843,N_372,N_3778);
or U9844 (N_9844,N_3404,N_4667);
and U9845 (N_9845,N_3750,N_1342);
xnor U9846 (N_9846,N_4625,N_1526);
or U9847 (N_9847,N_3113,N_4737);
nor U9848 (N_9848,N_1829,N_50);
or U9849 (N_9849,N_75,N_2908);
nor U9850 (N_9850,N_1779,N_286);
nor U9851 (N_9851,N_2326,N_3563);
or U9852 (N_9852,N_4077,N_3984);
and U9853 (N_9853,N_3669,N_4704);
nor U9854 (N_9854,N_3067,N_1656);
or U9855 (N_9855,N_2628,N_3529);
and U9856 (N_9856,N_607,N_2168);
or U9857 (N_9857,N_2335,N_1409);
nand U9858 (N_9858,N_1294,N_2214);
and U9859 (N_9859,N_1182,N_3376);
nand U9860 (N_9860,N_956,N_258);
and U9861 (N_9861,N_1008,N_1221);
nand U9862 (N_9862,N_1184,N_3195);
nor U9863 (N_9863,N_3431,N_919);
and U9864 (N_9864,N_4935,N_4255);
nand U9865 (N_9865,N_4098,N_4877);
xnor U9866 (N_9866,N_1719,N_956);
or U9867 (N_9867,N_4452,N_3119);
and U9868 (N_9868,N_1705,N_1642);
nor U9869 (N_9869,N_1255,N_2827);
xnor U9870 (N_9870,N_220,N_2872);
and U9871 (N_9871,N_3834,N_42);
nand U9872 (N_9872,N_2403,N_3229);
xnor U9873 (N_9873,N_2018,N_1495);
nor U9874 (N_9874,N_4139,N_769);
nor U9875 (N_9875,N_2815,N_1955);
and U9876 (N_9876,N_2039,N_3445);
nand U9877 (N_9877,N_4639,N_1810);
or U9878 (N_9878,N_1989,N_2269);
or U9879 (N_9879,N_3887,N_162);
xor U9880 (N_9880,N_4180,N_3797);
or U9881 (N_9881,N_3525,N_606);
nor U9882 (N_9882,N_1571,N_3011);
nand U9883 (N_9883,N_2627,N_1275);
and U9884 (N_9884,N_2455,N_4273);
nand U9885 (N_9885,N_1052,N_3607);
nor U9886 (N_9886,N_3661,N_3918);
nand U9887 (N_9887,N_1706,N_1462);
xnor U9888 (N_9888,N_2385,N_3595);
and U9889 (N_9889,N_3247,N_1036);
nor U9890 (N_9890,N_2491,N_4267);
or U9891 (N_9891,N_4106,N_1346);
nand U9892 (N_9892,N_3875,N_1922);
xnor U9893 (N_9893,N_2763,N_88);
and U9894 (N_9894,N_3459,N_4412);
nor U9895 (N_9895,N_1357,N_4948);
xnor U9896 (N_9896,N_2847,N_2842);
and U9897 (N_9897,N_413,N_1067);
nor U9898 (N_9898,N_3908,N_2650);
or U9899 (N_9899,N_4536,N_4131);
and U9900 (N_9900,N_4776,N_1623);
nor U9901 (N_9901,N_4185,N_3670);
or U9902 (N_9902,N_1847,N_4017);
nor U9903 (N_9903,N_390,N_539);
nor U9904 (N_9904,N_1493,N_2272);
nand U9905 (N_9905,N_1146,N_1742);
and U9906 (N_9906,N_4001,N_3984);
and U9907 (N_9907,N_2901,N_4056);
or U9908 (N_9908,N_1279,N_3099);
or U9909 (N_9909,N_2696,N_542);
nor U9910 (N_9910,N_2247,N_3734);
nand U9911 (N_9911,N_2525,N_362);
and U9912 (N_9912,N_3024,N_695);
and U9913 (N_9913,N_3177,N_4124);
nand U9914 (N_9914,N_4386,N_2555);
and U9915 (N_9915,N_1879,N_1855);
nand U9916 (N_9916,N_1634,N_1838);
and U9917 (N_9917,N_1059,N_3701);
nor U9918 (N_9918,N_2297,N_4376);
nor U9919 (N_9919,N_3875,N_2630);
or U9920 (N_9920,N_1996,N_4237);
nor U9921 (N_9921,N_1805,N_2025);
nor U9922 (N_9922,N_1361,N_1488);
nand U9923 (N_9923,N_3034,N_1184);
nand U9924 (N_9924,N_4012,N_292);
or U9925 (N_9925,N_2682,N_1619);
or U9926 (N_9926,N_2303,N_4986);
nand U9927 (N_9927,N_437,N_490);
and U9928 (N_9928,N_1710,N_1251);
or U9929 (N_9929,N_48,N_2895);
nor U9930 (N_9930,N_2761,N_2686);
nand U9931 (N_9931,N_1005,N_828);
or U9932 (N_9932,N_1898,N_4474);
nor U9933 (N_9933,N_1246,N_3947);
or U9934 (N_9934,N_3133,N_2337);
and U9935 (N_9935,N_1410,N_1329);
or U9936 (N_9936,N_322,N_4525);
xnor U9937 (N_9937,N_1921,N_3147);
or U9938 (N_9938,N_4054,N_2094);
nand U9939 (N_9939,N_1183,N_463);
and U9940 (N_9940,N_3308,N_57);
or U9941 (N_9941,N_3779,N_4074);
nand U9942 (N_9942,N_3655,N_3801);
xor U9943 (N_9943,N_1101,N_743);
nor U9944 (N_9944,N_1487,N_4802);
xnor U9945 (N_9945,N_2441,N_1632);
or U9946 (N_9946,N_3669,N_4579);
nor U9947 (N_9947,N_875,N_3118);
nor U9948 (N_9948,N_3243,N_3353);
and U9949 (N_9949,N_3291,N_2720);
or U9950 (N_9950,N_1856,N_1878);
xnor U9951 (N_9951,N_4267,N_4858);
nand U9952 (N_9952,N_1515,N_520);
and U9953 (N_9953,N_555,N_1318);
xnor U9954 (N_9954,N_700,N_1323);
nor U9955 (N_9955,N_4791,N_4982);
nand U9956 (N_9956,N_1416,N_193);
nand U9957 (N_9957,N_2097,N_4976);
nor U9958 (N_9958,N_4162,N_772);
nor U9959 (N_9959,N_838,N_2495);
xor U9960 (N_9960,N_4054,N_1509);
nand U9961 (N_9961,N_3670,N_3342);
xnor U9962 (N_9962,N_661,N_658);
and U9963 (N_9963,N_2815,N_3349);
xnor U9964 (N_9964,N_2833,N_1066);
xor U9965 (N_9965,N_3043,N_3731);
nand U9966 (N_9966,N_1079,N_3730);
or U9967 (N_9967,N_2173,N_1501);
and U9968 (N_9968,N_1624,N_3416);
xnor U9969 (N_9969,N_4135,N_160);
nand U9970 (N_9970,N_1278,N_4368);
nor U9971 (N_9971,N_3263,N_4721);
nand U9972 (N_9972,N_59,N_2910);
nor U9973 (N_9973,N_961,N_4720);
or U9974 (N_9974,N_3253,N_980);
nor U9975 (N_9975,N_3098,N_4347);
and U9976 (N_9976,N_855,N_1690);
xnor U9977 (N_9977,N_3825,N_2803);
nand U9978 (N_9978,N_467,N_3091);
or U9979 (N_9979,N_418,N_4427);
xnor U9980 (N_9980,N_2139,N_2949);
nand U9981 (N_9981,N_544,N_756);
nor U9982 (N_9982,N_4939,N_1245);
nor U9983 (N_9983,N_771,N_3622);
nor U9984 (N_9984,N_2378,N_4705);
or U9985 (N_9985,N_4699,N_3098);
nand U9986 (N_9986,N_2787,N_4295);
and U9987 (N_9987,N_4418,N_302);
and U9988 (N_9988,N_2904,N_1875);
or U9989 (N_9989,N_2197,N_2389);
or U9990 (N_9990,N_4165,N_1986);
and U9991 (N_9991,N_3921,N_3196);
or U9992 (N_9992,N_4758,N_3469);
nand U9993 (N_9993,N_103,N_3808);
and U9994 (N_9994,N_4077,N_1912);
and U9995 (N_9995,N_4737,N_3595);
nand U9996 (N_9996,N_2507,N_1388);
nand U9997 (N_9997,N_4778,N_2421);
nand U9998 (N_9998,N_3775,N_2687);
or U9999 (N_9999,N_3298,N_749);
or U10000 (N_10000,N_5822,N_7301);
nor U10001 (N_10001,N_6925,N_6372);
nor U10002 (N_10002,N_7171,N_9643);
xor U10003 (N_10003,N_7765,N_8579);
nand U10004 (N_10004,N_7569,N_8935);
nor U10005 (N_10005,N_6983,N_8005);
nor U10006 (N_10006,N_8233,N_9740);
and U10007 (N_10007,N_7878,N_8326);
or U10008 (N_10008,N_7063,N_6554);
nor U10009 (N_10009,N_9066,N_6246);
nor U10010 (N_10010,N_6706,N_6031);
xnor U10011 (N_10011,N_8716,N_6596);
nor U10012 (N_10012,N_5975,N_8495);
nand U10013 (N_10013,N_9328,N_9473);
nor U10014 (N_10014,N_8130,N_5853);
and U10015 (N_10015,N_7648,N_8477);
and U10016 (N_10016,N_9685,N_8010);
and U10017 (N_10017,N_9539,N_7131);
and U10018 (N_10018,N_5068,N_7120);
or U10019 (N_10019,N_7520,N_5575);
xnor U10020 (N_10020,N_5484,N_9981);
or U10021 (N_10021,N_6006,N_7393);
or U10022 (N_10022,N_6923,N_6858);
xnor U10023 (N_10023,N_9576,N_9480);
nor U10024 (N_10024,N_6690,N_5685);
xnor U10025 (N_10025,N_7904,N_9912);
nand U10026 (N_10026,N_5706,N_6829);
nand U10027 (N_10027,N_6151,N_5608);
nor U10028 (N_10028,N_5127,N_9761);
nand U10029 (N_10029,N_9925,N_8550);
and U10030 (N_10030,N_6254,N_8877);
or U10031 (N_10031,N_8372,N_8041);
nor U10032 (N_10032,N_9963,N_7481);
and U10033 (N_10033,N_7855,N_5360);
xor U10034 (N_10034,N_9383,N_8581);
and U10035 (N_10035,N_9844,N_9851);
nor U10036 (N_10036,N_7564,N_8172);
nor U10037 (N_10037,N_9217,N_8216);
xnor U10038 (N_10038,N_9107,N_9563);
nand U10039 (N_10039,N_8588,N_5411);
or U10040 (N_10040,N_7159,N_5747);
and U10041 (N_10041,N_7157,N_7138);
or U10042 (N_10042,N_7141,N_8297);
nand U10043 (N_10043,N_5114,N_7795);
nand U10044 (N_10044,N_9838,N_6806);
nand U10045 (N_10045,N_5789,N_7805);
nor U10046 (N_10046,N_8841,N_6675);
or U10047 (N_10047,N_6497,N_9406);
nand U10048 (N_10048,N_9397,N_8292);
and U10049 (N_10049,N_6307,N_7100);
xnor U10050 (N_10050,N_9693,N_7761);
nand U10051 (N_10051,N_9195,N_6998);
and U10052 (N_10052,N_5536,N_9171);
and U10053 (N_10053,N_9750,N_8534);
nand U10054 (N_10054,N_7209,N_8764);
or U10055 (N_10055,N_5204,N_8440);
nor U10056 (N_10056,N_5546,N_6038);
nor U10057 (N_10057,N_9163,N_7351);
xor U10058 (N_10058,N_6849,N_6773);
and U10059 (N_10059,N_8093,N_5303);
nand U10060 (N_10060,N_8171,N_6518);
and U10061 (N_10061,N_6244,N_6326);
or U10062 (N_10062,N_7501,N_8976);
and U10063 (N_10063,N_9276,N_5585);
or U10064 (N_10064,N_9306,N_9641);
and U10065 (N_10065,N_8343,N_5967);
nor U10066 (N_10066,N_5728,N_7265);
and U10067 (N_10067,N_5952,N_8502);
or U10068 (N_10068,N_8702,N_9338);
or U10069 (N_10069,N_7626,N_9979);
or U10070 (N_10070,N_9872,N_7934);
or U10071 (N_10071,N_9274,N_7468);
nor U10072 (N_10072,N_9772,N_9803);
nand U10073 (N_10073,N_9719,N_9067);
and U10074 (N_10074,N_7603,N_7877);
and U10075 (N_10075,N_8760,N_6471);
or U10076 (N_10076,N_9653,N_8142);
nor U10077 (N_10077,N_7798,N_7740);
xor U10078 (N_10078,N_8674,N_9123);
and U10079 (N_10079,N_9879,N_6229);
nand U10080 (N_10080,N_6939,N_9029);
nor U10081 (N_10081,N_7197,N_6561);
nand U10082 (N_10082,N_9672,N_8788);
and U10083 (N_10083,N_8373,N_9799);
nor U10084 (N_10084,N_9021,N_7738);
or U10085 (N_10085,N_5383,N_6959);
or U10086 (N_10086,N_7349,N_8057);
and U10087 (N_10087,N_7443,N_8724);
and U10088 (N_10088,N_8254,N_8955);
nor U10089 (N_10089,N_9285,N_8381);
nor U10090 (N_10090,N_5920,N_6450);
and U10091 (N_10091,N_8409,N_9730);
and U10092 (N_10092,N_8246,N_5026);
nor U10093 (N_10093,N_5462,N_5556);
xnor U10094 (N_10094,N_5046,N_7371);
nor U10095 (N_10095,N_7010,N_7021);
and U10096 (N_10096,N_9253,N_8896);
nor U10097 (N_10097,N_6490,N_6402);
xnor U10098 (N_10098,N_8457,N_6435);
nand U10099 (N_10099,N_9119,N_7514);
nor U10100 (N_10100,N_5309,N_8344);
nand U10101 (N_10101,N_7561,N_9692);
and U10102 (N_10102,N_5380,N_9177);
nand U10103 (N_10103,N_9402,N_7772);
or U10104 (N_10104,N_9261,N_9807);
nand U10105 (N_10105,N_8771,N_8277);
nor U10106 (N_10106,N_9828,N_8979);
or U10107 (N_10107,N_5979,N_8094);
or U10108 (N_10108,N_5085,N_6902);
nand U10109 (N_10109,N_6569,N_5033);
nor U10110 (N_10110,N_9512,N_8134);
nand U10111 (N_10111,N_8736,N_8335);
nand U10112 (N_10112,N_5633,N_7774);
nand U10113 (N_10113,N_8643,N_5671);
nor U10114 (N_10114,N_8739,N_9068);
and U10115 (N_10115,N_8837,N_7224);
nor U10116 (N_10116,N_9348,N_6651);
xnor U10117 (N_10117,N_6404,N_6265);
or U10118 (N_10118,N_9428,N_6092);
or U10119 (N_10119,N_5404,N_8988);
nand U10120 (N_10120,N_7181,N_6528);
nand U10121 (N_10121,N_5661,N_6467);
xor U10122 (N_10122,N_5646,N_5654);
nand U10123 (N_10123,N_8571,N_7353);
xor U10124 (N_10124,N_8671,N_8719);
or U10125 (N_10125,N_6974,N_5888);
nand U10126 (N_10126,N_7567,N_8384);
or U10127 (N_10127,N_8291,N_5637);
or U10128 (N_10128,N_6687,N_8198);
or U10129 (N_10129,N_7293,N_9247);
nor U10130 (N_10130,N_9291,N_6332);
nor U10131 (N_10131,N_5369,N_8076);
nand U10132 (N_10132,N_7009,N_5140);
or U10133 (N_10133,N_7463,N_5149);
or U10134 (N_10134,N_5902,N_5651);
or U10135 (N_10135,N_6711,N_5418);
nor U10136 (N_10136,N_7883,N_9836);
or U10137 (N_10137,N_8921,N_8572);
and U10138 (N_10138,N_9630,N_7145);
nor U10139 (N_10139,N_5817,N_7426);
or U10140 (N_10140,N_7433,N_8302);
nand U10141 (N_10141,N_7756,N_9548);
nor U10142 (N_10142,N_6146,N_6012);
and U10143 (N_10143,N_6411,N_5222);
nor U10144 (N_10144,N_5214,N_5399);
or U10145 (N_10145,N_5820,N_8023);
nor U10146 (N_10146,N_7226,N_9051);
and U10147 (N_10147,N_8079,N_8768);
xor U10148 (N_10148,N_9041,N_5010);
and U10149 (N_10149,N_8690,N_9189);
nand U10150 (N_10150,N_5577,N_9266);
nor U10151 (N_10151,N_6514,N_8648);
and U10152 (N_10152,N_9385,N_5228);
and U10153 (N_10153,N_6501,N_8725);
or U10154 (N_10154,N_7018,N_5537);
or U10155 (N_10155,N_5761,N_9040);
or U10156 (N_10156,N_8063,N_8073);
or U10157 (N_10157,N_7870,N_9495);
nor U10158 (N_10158,N_8106,N_6359);
or U10159 (N_10159,N_9074,N_9454);
xor U10160 (N_10160,N_5273,N_5672);
and U10161 (N_10161,N_7415,N_5494);
and U10162 (N_10162,N_5514,N_5843);
nor U10163 (N_10163,N_6734,N_7834);
nor U10164 (N_10164,N_9701,N_9344);
and U10165 (N_10165,N_8267,N_5131);
and U10166 (N_10166,N_9880,N_6118);
nor U10167 (N_10167,N_7671,N_8242);
xor U10168 (N_10168,N_6061,N_7339);
or U10169 (N_10169,N_5417,N_9377);
or U10170 (N_10170,N_5885,N_5864);
nor U10171 (N_10171,N_6907,N_8308);
nand U10172 (N_10172,N_7030,N_8113);
nand U10173 (N_10173,N_7780,N_7162);
nand U10174 (N_10174,N_8109,N_8226);
nand U10175 (N_10175,N_7135,N_6245);
nor U10176 (N_10176,N_5136,N_7322);
or U10177 (N_10177,N_7178,N_7570);
xnor U10178 (N_10178,N_5258,N_7698);
and U10179 (N_10179,N_5301,N_5879);
xnor U10180 (N_10180,N_6294,N_5251);
and U10181 (N_10181,N_7900,N_6540);
nand U10182 (N_10182,N_5117,N_8673);
nand U10183 (N_10183,N_5862,N_5054);
nand U10184 (N_10184,N_7440,N_5091);
and U10185 (N_10185,N_6367,N_8784);
nand U10186 (N_10186,N_6495,N_6105);
or U10187 (N_10187,N_7649,N_7260);
and U10188 (N_10188,N_8456,N_8783);
nand U10189 (N_10189,N_7139,N_8249);
xnor U10190 (N_10190,N_9976,N_5996);
or U10191 (N_10191,N_5682,N_6016);
nor U10192 (N_10192,N_9901,N_5423);
xnor U10193 (N_10193,N_8666,N_8547);
and U10194 (N_10194,N_6476,N_7627);
and U10195 (N_10195,N_9884,N_6050);
nor U10196 (N_10196,N_8580,N_8053);
or U10197 (N_10197,N_6887,N_8863);
and U10198 (N_10198,N_5825,N_7860);
and U10199 (N_10199,N_5976,N_9094);
nor U10200 (N_10200,N_9547,N_7960);
nand U10201 (N_10201,N_5405,N_8668);
and U10202 (N_10202,N_5074,N_5437);
nor U10203 (N_10203,N_9149,N_9581);
or U10204 (N_10204,N_7625,N_5406);
nand U10205 (N_10205,N_7238,N_7523);
xnor U10206 (N_10206,N_9129,N_9759);
or U10207 (N_10207,N_8622,N_9399);
nor U10208 (N_10208,N_6594,N_5611);
or U10209 (N_10209,N_7189,N_6795);
and U10210 (N_10210,N_9343,N_9382);
xnor U10211 (N_10211,N_9042,N_8876);
or U10212 (N_10212,N_5714,N_6761);
or U10213 (N_10213,N_5689,N_6396);
or U10214 (N_10214,N_5259,N_5006);
xnor U10215 (N_10215,N_9505,N_7168);
or U10216 (N_10216,N_5512,N_8072);
and U10217 (N_10217,N_5015,N_7993);
and U10218 (N_10218,N_6340,N_8872);
nor U10219 (N_10219,N_5012,N_6606);
and U10220 (N_10220,N_9452,N_7070);
and U10221 (N_10221,N_5754,N_8592);
nor U10222 (N_10222,N_7650,N_9560);
xnor U10223 (N_10223,N_9668,N_7243);
nand U10224 (N_10224,N_9186,N_9591);
or U10225 (N_10225,N_5819,N_7111);
nand U10226 (N_10226,N_6710,N_6169);
and U10227 (N_10227,N_6364,N_7801);
nor U10228 (N_10228,N_5076,N_6993);
or U10229 (N_10229,N_9112,N_7092);
nand U10230 (N_10230,N_7644,N_7606);
or U10231 (N_10231,N_5098,N_5891);
and U10232 (N_10232,N_5687,N_5184);
or U10233 (N_10233,N_9419,N_6756);
or U10234 (N_10234,N_8818,N_9064);
xor U10235 (N_10235,N_5543,N_6778);
nand U10236 (N_10236,N_8660,N_6022);
nand U10237 (N_10237,N_9284,N_8555);
or U10238 (N_10238,N_5688,N_5381);
and U10239 (N_10239,N_5529,N_7390);
xor U10240 (N_10240,N_6285,N_6878);
and U10241 (N_10241,N_6978,N_7673);
nor U10242 (N_10242,N_9648,N_5660);
xnor U10243 (N_10243,N_8672,N_6004);
nand U10244 (N_10244,N_5275,N_8449);
or U10245 (N_10245,N_7205,N_6349);
nand U10246 (N_10246,N_5621,N_5223);
nand U10247 (N_10247,N_6830,N_5827);
nand U10248 (N_10248,N_7953,N_8746);
and U10249 (N_10249,N_6231,N_8484);
nand U10250 (N_10250,N_8039,N_8982);
nand U10251 (N_10251,N_5846,N_6701);
nand U10252 (N_10252,N_8032,N_7096);
and U10253 (N_10253,N_6366,N_6927);
nand U10254 (N_10254,N_5315,N_5851);
and U10255 (N_10255,N_9026,N_9546);
nand U10256 (N_10256,N_5513,N_8756);
nand U10257 (N_10257,N_9786,N_6815);
nor U10258 (N_10258,N_8404,N_9554);
or U10259 (N_10259,N_6931,N_6929);
nand U10260 (N_10260,N_9613,N_9680);
nand U10261 (N_10261,N_5778,N_5833);
nor U10262 (N_10262,N_8853,N_6236);
or U10263 (N_10263,N_9824,N_5558);
nor U10264 (N_10264,N_5370,N_6781);
and U10265 (N_10265,N_6719,N_9293);
xnor U10266 (N_10266,N_5440,N_6228);
nand U10267 (N_10267,N_7763,N_5898);
xnor U10268 (N_10268,N_6434,N_7762);
or U10269 (N_10269,N_8481,N_7277);
and U10270 (N_10270,N_6992,N_8252);
or U10271 (N_10271,N_5872,N_5348);
and U10272 (N_10272,N_6309,N_9037);
and U10273 (N_10273,N_9661,N_6324);
xor U10274 (N_10274,N_9278,N_5697);
and U10275 (N_10275,N_6030,N_9651);
and U10276 (N_10276,N_6593,N_8358);
or U10277 (N_10277,N_7640,N_7326);
nand U10278 (N_10278,N_6913,N_7641);
or U10279 (N_10279,N_9566,N_6612);
nand U10280 (N_10280,N_5784,N_8900);
or U10281 (N_10281,N_9489,N_8488);
xor U10282 (N_10282,N_5663,N_8575);
nand U10283 (N_10283,N_6323,N_7896);
nor U10284 (N_10284,N_6345,N_5670);
nand U10285 (N_10285,N_7005,N_7058);
xnor U10286 (N_10286,N_7931,N_7613);
or U10287 (N_10287,N_7519,N_5524);
and U10288 (N_10288,N_5984,N_7656);
or U10289 (N_10289,N_8993,N_6712);
and U10290 (N_10290,N_6592,N_9118);
or U10291 (N_10291,N_6237,N_7084);
nand U10292 (N_10292,N_8578,N_7620);
nor U10293 (N_10293,N_8056,N_7566);
nor U10294 (N_10294,N_5506,N_5354);
and U10295 (N_10295,N_6667,N_6219);
xnor U10296 (N_10296,N_6032,N_5106);
and U10297 (N_10297,N_7492,N_6808);
xnor U10298 (N_10298,N_6104,N_6224);
or U10299 (N_10299,N_5187,N_7269);
xnor U10300 (N_10300,N_6338,N_5634);
or U10301 (N_10301,N_7786,N_7331);
or U10302 (N_10302,N_8914,N_5464);
nor U10303 (N_10303,N_7592,N_6763);
and U10304 (N_10304,N_6972,N_8593);
nand U10305 (N_10305,N_5375,N_7861);
nand U10306 (N_10306,N_5238,N_6744);
nand U10307 (N_10307,N_6871,N_6089);
nor U10308 (N_10308,N_5248,N_8854);
nand U10309 (N_10309,N_8100,N_5014);
or U10310 (N_10310,N_9430,N_8688);
nand U10311 (N_10311,N_7305,N_8713);
nor U10312 (N_10312,N_8433,N_6011);
or U10313 (N_10313,N_8087,N_6314);
nand U10314 (N_10314,N_8884,N_6835);
or U10315 (N_10315,N_9022,N_7513);
nor U10316 (N_10316,N_5812,N_6156);
and U10317 (N_10317,N_8611,N_9366);
and U10318 (N_10318,N_8891,N_5834);
nor U10319 (N_10319,N_6602,N_6197);
nor U10320 (N_10320,N_6652,N_7548);
and U10321 (N_10321,N_5451,N_6117);
nand U10322 (N_10322,N_8882,N_9146);
nand U10323 (N_10323,N_9852,N_8238);
nor U10324 (N_10324,N_7716,N_7515);
and U10325 (N_10325,N_7085,N_5069);
and U10326 (N_10326,N_7347,N_5174);
xor U10327 (N_10327,N_9464,N_5769);
nand U10328 (N_10328,N_8930,N_6910);
nor U10329 (N_10329,N_5202,N_5804);
nand U10330 (N_10330,N_5636,N_9075);
nand U10331 (N_10331,N_8647,N_8392);
nor U10332 (N_10332,N_7605,N_5983);
and U10333 (N_10333,N_8257,N_7137);
nor U10334 (N_10334,N_6933,N_6318);
nor U10335 (N_10335,N_9705,N_6376);
nand U10336 (N_10336,N_5582,N_8119);
nand U10337 (N_10337,N_9928,N_8926);
and U10338 (N_10338,N_6132,N_9466);
or U10339 (N_10339,N_5393,N_6512);
nand U10340 (N_10340,N_5058,N_5141);
or U10341 (N_10341,N_9179,N_7253);
or U10342 (N_10342,N_5622,N_6258);
xnor U10343 (N_10343,N_7066,N_6759);
and U10344 (N_10344,N_8019,N_9131);
or U10345 (N_10345,N_5762,N_5528);
and U10346 (N_10346,N_9919,N_6915);
xnor U10347 (N_10347,N_6377,N_6157);
nand U10348 (N_10348,N_6166,N_6948);
xor U10349 (N_10349,N_6426,N_9506);
nand U10350 (N_10350,N_6387,N_9762);
and U10351 (N_10351,N_6867,N_9360);
and U10352 (N_10352,N_7289,N_7571);
nand U10353 (N_10353,N_6358,N_7509);
and U10354 (N_10354,N_6056,N_7543);
xor U10355 (N_10355,N_8312,N_7027);
and U10356 (N_10356,N_6715,N_6670);
and U10357 (N_10357,N_5592,N_5286);
or U10358 (N_10358,N_7424,N_7242);
nand U10359 (N_10359,N_7779,N_5110);
and U10360 (N_10360,N_7741,N_6393);
nand U10361 (N_10361,N_8351,N_5908);
or U10362 (N_10362,N_8002,N_8469);
nor U10363 (N_10363,N_7858,N_6453);
or U10364 (N_10364,N_9053,N_7955);
or U10365 (N_10365,N_5379,N_7402);
or U10366 (N_10366,N_9472,N_5549);
nand U10367 (N_10367,N_6587,N_6304);
nand U10368 (N_10368,N_8086,N_7928);
xor U10369 (N_10369,N_8188,N_9335);
or U10370 (N_10370,N_6429,N_7484);
and U10371 (N_10371,N_9126,N_5180);
nor U10372 (N_10372,N_5596,N_5764);
or U10373 (N_10373,N_5758,N_8551);
nand U10374 (N_10374,N_9633,N_6053);
nand U10375 (N_10375,N_8868,N_5115);
or U10376 (N_10376,N_5426,N_6582);
and U10377 (N_10377,N_5724,N_6639);
nor U10378 (N_10378,N_6834,N_9756);
nand U10379 (N_10379,N_8175,N_5037);
and U10380 (N_10380,N_7156,N_6538);
or U10381 (N_10381,N_9393,N_6215);
xor U10382 (N_10382,N_6873,N_5378);
nor U10383 (N_10383,N_5619,N_6519);
or U10384 (N_10384,N_8330,N_7436);
or U10385 (N_10385,N_9455,N_8055);
nor U10386 (N_10386,N_9272,N_5224);
nor U10387 (N_10387,N_6638,N_9818);
and U10388 (N_10388,N_8465,N_8374);
or U10389 (N_10389,N_7479,N_5385);
nor U10390 (N_10390,N_8888,N_7488);
nor U10391 (N_10391,N_6264,N_7752);
and U10392 (N_10392,N_8275,N_9173);
xnor U10393 (N_10393,N_5624,N_8968);
xnor U10394 (N_10394,N_5516,N_5583);
and U10395 (N_10395,N_9805,N_8043);
nand U10396 (N_10396,N_7701,N_8097);
nand U10397 (N_10397,N_6328,N_5145);
nand U10398 (N_10398,N_5161,N_7236);
and U10399 (N_10399,N_5992,N_7867);
nor U10400 (N_10400,N_9557,N_7787);
or U10401 (N_10401,N_9116,N_6418);
or U10402 (N_10402,N_8696,N_6783);
or U10403 (N_10403,N_6828,N_8064);
nor U10404 (N_10404,N_8443,N_8516);
and U10405 (N_10405,N_9984,N_5221);
nand U10406 (N_10406,N_8947,N_5230);
nand U10407 (N_10407,N_8667,N_5120);
nor U10408 (N_10408,N_5072,N_9535);
or U10409 (N_10409,N_9739,N_5295);
and U10410 (N_10410,N_6447,N_9302);
nor U10411 (N_10411,N_5032,N_5531);
nor U10412 (N_10412,N_6472,N_5613);
nor U10413 (N_10413,N_9114,N_8468);
nor U10414 (N_10414,N_7366,N_7706);
nand U10415 (N_10415,N_9649,N_5580);
nand U10416 (N_10416,N_5774,N_6613);
nand U10417 (N_10417,N_8273,N_9746);
or U10418 (N_10418,N_5065,N_7689);
and U10419 (N_10419,N_7694,N_8627);
and U10420 (N_10420,N_9604,N_8451);
or U10421 (N_10421,N_7327,N_8981);
nand U10422 (N_10422,N_7401,N_9590);
nor U10423 (N_10423,N_8345,N_7106);
nor U10424 (N_10424,N_8977,N_8809);
nor U10425 (N_10425,N_7225,N_6239);
nor U10426 (N_10426,N_5288,N_9660);
nand U10427 (N_10427,N_6257,N_7237);
nor U10428 (N_10428,N_5859,N_6449);
and U10429 (N_10429,N_8923,N_6293);
and U10430 (N_10430,N_9570,N_7099);
or U10431 (N_10431,N_5433,N_9665);
nand U10432 (N_10432,N_9446,N_6421);
nand U10433 (N_10433,N_8313,N_7345);
nand U10434 (N_10434,N_8281,N_7288);
xor U10435 (N_10435,N_8124,N_9374);
and U10436 (N_10436,N_8804,N_5374);
nand U10437 (N_10437,N_9626,N_6746);
nor U10438 (N_10438,N_6253,N_7060);
nor U10439 (N_10439,N_6242,N_8943);
nor U10440 (N_10440,N_6570,N_8807);
nor U10441 (N_10441,N_8911,N_7945);
nor U10442 (N_10442,N_9589,N_5217);
and U10443 (N_10443,N_6339,N_8974);
xor U10444 (N_10444,N_6352,N_9038);
nand U10445 (N_10445,N_8399,N_7802);
nand U10446 (N_10446,N_9704,N_5461);
nor U10447 (N_10447,N_8211,N_8733);
nor U10448 (N_10448,N_6713,N_5605);
nor U10449 (N_10449,N_5331,N_8522);
xor U10450 (N_10450,N_8410,N_7491);
nand U10451 (N_10451,N_6041,N_6702);
or U10452 (N_10452,N_8180,N_5503);
nor U10453 (N_10453,N_7538,N_6775);
and U10454 (N_10454,N_5290,N_5403);
nor U10455 (N_10455,N_6508,N_7300);
nor U10456 (N_10456,N_5617,N_6850);
and U10457 (N_10457,N_7483,N_6020);
or U10458 (N_10458,N_8792,N_9615);
and U10459 (N_10459,N_9178,N_9375);
nor U10460 (N_10460,N_9445,N_6862);
xnor U10461 (N_10461,N_9155,N_8241);
nor U10462 (N_10462,N_9175,N_9013);
or U10463 (N_10463,N_8245,N_6462);
nand U10464 (N_10464,N_6378,N_5750);
or U10465 (N_10465,N_8544,N_7328);
and U10466 (N_10466,N_6628,N_5828);
or U10467 (N_10467,N_8081,N_8274);
nand U10468 (N_10468,N_5082,N_8220);
nor U10469 (N_10469,N_7185,N_8678);
and U10470 (N_10470,N_9198,N_7464);
nand U10471 (N_10471,N_7874,N_5708);
and U10472 (N_10472,N_8046,N_6704);
nand U10473 (N_10473,N_7586,N_8560);
and U10474 (N_10474,N_6438,N_8118);
nand U10475 (N_10475,N_6357,N_9150);
nand U10476 (N_10476,N_8029,N_7791);
and U10477 (N_10477,N_7524,N_5802);
or U10478 (N_10478,N_6654,N_8607);
nor U10479 (N_10479,N_6319,N_9502);
nand U10480 (N_10480,N_7800,N_9597);
or U10481 (N_10481,N_6938,N_5738);
nor U10482 (N_10482,N_9248,N_8787);
or U10483 (N_10483,N_7518,N_8624);
or U10484 (N_10484,N_8475,N_7034);
nand U10485 (N_10485,N_5680,N_8362);
and U10486 (N_10486,N_7266,N_9656);
and U10487 (N_10487,N_5126,N_7490);
nand U10488 (N_10488,N_9136,N_9915);
nor U10489 (N_10489,N_7582,N_8820);
nand U10490 (N_10490,N_6875,N_7664);
nor U10491 (N_10491,N_6233,N_9227);
nand U10492 (N_10492,N_7635,N_7580);
xor U10493 (N_10493,N_9237,N_7685);
or U10494 (N_10494,N_5903,N_7405);
or U10495 (N_10495,N_8621,N_8428);
nor U10496 (N_10496,N_7202,N_7578);
and U10497 (N_10497,N_5121,N_9349);
or U10498 (N_10498,N_8377,N_8963);
nand U10499 (N_10499,N_8682,N_8411);
nor U10500 (N_10500,N_6548,N_8918);
and U10501 (N_10501,N_6909,N_6240);
nand U10502 (N_10502,N_7816,N_9065);
nand U10503 (N_10503,N_9931,N_6070);
xor U10504 (N_10504,N_5739,N_9048);
or U10505 (N_10505,N_5988,N_9236);
or U10506 (N_10506,N_9716,N_7248);
nor U10507 (N_10507,N_8367,N_9695);
nor U10508 (N_10508,N_5919,N_7647);
nand U10509 (N_10509,N_5087,N_9577);
or U10510 (N_10510,N_6180,N_7645);
or U10511 (N_10511,N_7367,N_8722);
nand U10512 (N_10512,N_7444,N_9642);
nor U10513 (N_10513,N_5876,N_6174);
nand U10514 (N_10514,N_9970,N_7544);
and U10515 (N_10515,N_5735,N_9708);
and U10516 (N_10516,N_9271,N_7485);
nand U10517 (N_10517,N_5355,N_9376);
or U10518 (N_10518,N_7051,N_9133);
nand U10519 (N_10519,N_5541,N_7105);
and U10520 (N_10520,N_8303,N_6260);
nand U10521 (N_10521,N_9994,N_5994);
or U10522 (N_10522,N_7746,N_5377);
nor U10523 (N_10523,N_9254,N_8638);
nor U10524 (N_10524,N_5321,N_6102);
nand U10525 (N_10525,N_5137,N_5029);
or U10526 (N_10526,N_7677,N_9120);
xnor U10527 (N_10527,N_8442,N_5499);
and U10528 (N_10528,N_6975,N_7452);
nor U10529 (N_10529,N_8375,N_6057);
or U10530 (N_10530,N_8288,N_5573);
and U10531 (N_10531,N_8224,N_6172);
xnor U10532 (N_10532,N_6111,N_6386);
xor U10533 (N_10533,N_9965,N_8887);
or U10534 (N_10534,N_5244,N_8342);
and U10535 (N_10535,N_9501,N_7359);
nor U10536 (N_10536,N_9456,N_7743);
and U10537 (N_10537,N_8957,N_8718);
nor U10538 (N_10538,N_8685,N_5718);
nand U10539 (N_10539,N_6475,N_8363);
or U10540 (N_10540,N_5476,N_8557);
nor U10541 (N_10541,N_8024,N_9610);
nor U10542 (N_10542,N_8054,N_8431);
nand U10543 (N_10543,N_5119,N_8800);
nor U10544 (N_10544,N_5160,N_8531);
nand U10545 (N_10545,N_9532,N_6230);
xnor U10546 (N_10546,N_5757,N_9381);
nand U10547 (N_10547,N_6097,N_6441);
nand U10548 (N_10548,N_7807,N_9905);
and U10549 (N_10549,N_8289,N_9077);
nand U10550 (N_10550,N_8686,N_6069);
or U10551 (N_10551,N_6621,N_7019);
nor U10552 (N_10552,N_7227,N_9487);
nand U10553 (N_10553,N_8825,N_7336);
or U10554 (N_10554,N_8324,N_6185);
nor U10555 (N_10555,N_9043,N_7398);
nand U10556 (N_10556,N_7587,N_7192);
nor U10557 (N_10557,N_7136,N_8759);
nand U10558 (N_10558,N_7091,N_7132);
nor U10559 (N_10559,N_8992,N_5239);
and U10560 (N_10560,N_5135,N_7957);
nand U10561 (N_10561,N_8852,N_9004);
nor U10562 (N_10562,N_8390,N_9900);
nor U10563 (N_10563,N_9010,N_6967);
and U10564 (N_10564,N_9488,N_8806);
nor U10565 (N_10565,N_5387,N_8341);
and U10566 (N_10566,N_6940,N_8000);
and U10567 (N_10567,N_8239,N_5045);
nor U10568 (N_10568,N_5460,N_6688);
nand U10569 (N_10569,N_8170,N_5597);
nand U10570 (N_10570,N_9717,N_8675);
and U10571 (N_10571,N_5061,N_5568);
xnor U10572 (N_10572,N_7041,N_9491);
nand U10573 (N_10573,N_9974,N_8697);
and U10574 (N_10574,N_8114,N_6433);
nand U10575 (N_10575,N_8649,N_5727);
xor U10576 (N_10576,N_6881,N_8121);
xnor U10577 (N_10577,N_5914,N_6901);
or U10578 (N_10578,N_8355,N_5416);
or U10579 (N_10579,N_7254,N_5409);
nand U10580 (N_10580,N_8867,N_9494);
and U10581 (N_10581,N_6585,N_8949);
or U10582 (N_10582,N_7476,N_8145);
and U10583 (N_10583,N_8898,N_8664);
nand U10584 (N_10584,N_8741,N_6296);
nand U10585 (N_10585,N_5686,N_5553);
nor U10586 (N_10586,N_7061,N_5742);
nor U10587 (N_10587,N_9682,N_9176);
or U10588 (N_10588,N_7856,N_6459);
nor U10589 (N_10589,N_6177,N_6695);
and U10590 (N_10590,N_9474,N_5760);
or U10591 (N_10591,N_7375,N_9517);
nor U10592 (N_10592,N_6969,N_7451);
nor U10593 (N_10593,N_9798,N_5857);
nor U10594 (N_10594,N_8727,N_6511);
xnor U10595 (N_10595,N_7221,N_6154);
and U10596 (N_10596,N_6678,N_9996);
nor U10597 (N_10597,N_5001,N_6179);
xor U10598 (N_10598,N_5265,N_9952);
nor U10599 (N_10599,N_6204,N_8670);
or U10600 (N_10600,N_5518,N_7907);
and U10601 (N_10601,N_8708,N_8129);
nor U10602 (N_10602,N_5849,N_7094);
and U10603 (N_10603,N_8083,N_7072);
nand U10604 (N_10604,N_5951,N_6019);
and U10605 (N_10605,N_8479,N_5427);
nor U10606 (N_10606,N_8951,N_8447);
nor U10607 (N_10607,N_5629,N_5326);
and U10608 (N_10608,N_8194,N_9203);
or U10609 (N_10609,N_5143,N_7639);
and U10610 (N_10610,N_8796,N_7862);
nor U10611 (N_10611,N_9005,N_7596);
xor U10612 (N_10612,N_5188,N_7913);
nor U10613 (N_10613,N_5591,N_6039);
and U10614 (N_10614,N_7325,N_6281);
and U10615 (N_10615,N_7245,N_8600);
nand U10616 (N_10616,N_5658,N_8791);
nand U10617 (N_10617,N_5269,N_5765);
and U10618 (N_10618,N_5028,N_6664);
or U10619 (N_10619,N_7196,N_5723);
nand U10620 (N_10620,N_6899,N_7822);
xnor U10621 (N_10621,N_6741,N_7275);
nand U10622 (N_10622,N_9072,N_9619);
nor U10623 (N_10623,N_7332,N_7865);
and U10624 (N_10624,N_6048,N_7611);
xnor U10625 (N_10625,N_8153,N_7442);
or U10626 (N_10626,N_6524,N_9518);
and U10627 (N_10627,N_5521,N_9972);
xnor U10628 (N_10628,N_9569,N_6860);
xor U10629 (N_10629,N_9082,N_6786);
nor U10630 (N_10630,N_8545,N_6208);
or U10631 (N_10631,N_7175,N_8017);
nor U10632 (N_10632,N_9507,N_6591);
and U10633 (N_10633,N_8623,N_9684);
or U10634 (N_10634,N_8606,N_7702);
or U10635 (N_10635,N_5152,N_8378);
and U10636 (N_10636,N_7109,N_7340);
nand U10637 (N_10637,N_5716,N_7059);
nand U10638 (N_10638,N_7542,N_8511);
and U10639 (N_10639,N_8208,N_9054);
nand U10640 (N_10640,N_9796,N_9967);
or U10641 (N_10641,N_7024,N_9538);
nand U10642 (N_10642,N_8790,N_6175);
and U10643 (N_10643,N_8635,N_9424);
nor U10644 (N_10644,N_6008,N_7153);
and U10645 (N_10645,N_7583,N_5197);
nor U10646 (N_10646,N_6216,N_8230);
or U10647 (N_10647,N_7049,N_7246);
or U10648 (N_10648,N_7046,N_7204);
nor U10649 (N_10649,N_8892,N_5628);
nand U10650 (N_10650,N_9251,N_7872);
or U10651 (N_10651,N_7962,N_7247);
and U10652 (N_10652,N_9137,N_8128);
and U10653 (N_10653,N_6921,N_9442);
nor U10654 (N_10654,N_9891,N_8350);
nand U10655 (N_10655,N_8098,N_6313);
or U10656 (N_10656,N_8307,N_6633);
nand U10657 (N_10657,N_8474,N_9056);
nand U10658 (N_10658,N_7597,N_8902);
xor U10659 (N_10659,N_7158,N_6080);
nor U10660 (N_10660,N_8315,N_9835);
and U10661 (N_10661,N_6001,N_6481);
and U10662 (N_10662,N_9329,N_6517);
or U10663 (N_10663,N_6757,N_9006);
nor U10664 (N_10664,N_6370,N_6770);
xnor U10665 (N_10665,N_5896,N_5593);
nor U10666 (N_10666,N_8813,N_6752);
and U10667 (N_10667,N_8812,N_6297);
nor U10668 (N_10668,N_5093,N_6412);
nand U10669 (N_10669,N_9543,N_9460);
or U10670 (N_10670,N_9827,N_7956);
nand U10671 (N_10671,N_8190,N_8207);
nor U10672 (N_10672,N_7403,N_7556);
and U10673 (N_10673,N_5071,N_9541);
nand U10674 (N_10674,N_7577,N_9034);
and U10675 (N_10675,N_5367,N_7337);
or U10676 (N_10676,N_7517,N_6696);
xor U10677 (N_10677,N_8317,N_6700);
nand U10678 (N_10678,N_8223,N_9011);
nor U10679 (N_10679,N_9544,N_9748);
or U10680 (N_10680,N_8543,N_6788);
nor U10681 (N_10681,N_7078,N_6300);
and U10682 (N_10682,N_7886,N_8014);
or U10683 (N_10683,N_8753,N_7675);
xnor U10684 (N_10684,N_6533,N_7825);
and U10685 (N_10685,N_7552,N_9448);
nand U10686 (N_10686,N_9192,N_5799);
or U10687 (N_10687,N_9386,N_6745);
and U10688 (N_10688,N_6085,N_8931);
nand U10689 (N_10689,N_6692,N_7095);
and U10690 (N_10690,N_6970,N_5547);
xnor U10691 (N_10691,N_5973,N_7952);
or U10692 (N_10692,N_7231,N_5737);
or U10693 (N_10693,N_7549,N_6999);
nor U10694 (N_10694,N_8989,N_5296);
and U10695 (N_10695,N_8613,N_6241);
nand U10696 (N_10696,N_9421,N_7575);
nand U10697 (N_10697,N_6238,N_5011);
nor U10698 (N_10698,N_5559,N_5702);
nor U10699 (N_10699,N_5457,N_9727);
and U10700 (N_10700,N_6730,N_6482);
nand U10701 (N_10701,N_9999,N_7222);
and U10702 (N_10702,N_6095,N_9595);
xor U10703 (N_10703,N_9154,N_9212);
nor U10704 (N_10704,N_5995,N_9890);
nand U10705 (N_10705,N_6708,N_5133);
nor U10706 (N_10706,N_7194,N_6790);
and U10707 (N_10707,N_8004,N_5007);
or U10708 (N_10708,N_5806,N_8031);
nor U10709 (N_10709,N_6405,N_6990);
nor U10710 (N_10710,N_5479,N_9788);
and U10711 (N_10711,N_8371,N_9971);
or U10712 (N_10712,N_6355,N_8585);
and U10713 (N_10713,N_5725,N_7739);
nor U10714 (N_10714,N_5644,N_7880);
nor U10715 (N_10715,N_7125,N_9108);
nand U10716 (N_10716,N_7417,N_6575);
and U10717 (N_10717,N_8107,N_5112);
nor U10718 (N_10718,N_7083,N_6748);
nor U10719 (N_10719,N_8770,N_6547);
and U10720 (N_10720,N_6637,N_6013);
nand U10721 (N_10721,N_7352,N_8501);
and U10722 (N_10722,N_9061,N_9568);
nor U10723 (N_10723,N_7420,N_9134);
nand U10724 (N_10724,N_6749,N_6306);
nand U10725 (N_10725,N_6573,N_5240);
nand U10726 (N_10726,N_7127,N_6941);
xor U10727 (N_10727,N_6947,N_5047);
nand U10728 (N_10728,N_6584,N_7511);
nand U10729 (N_10729,N_7917,N_6735);
nor U10730 (N_10730,N_8049,N_5083);
xor U10731 (N_10731,N_8895,N_5563);
nand U10732 (N_10732,N_8821,N_7888);
nor U10733 (N_10733,N_8785,N_9841);
nor U10734 (N_10734,N_9700,N_9132);
and U10735 (N_10735,N_5740,N_9092);
nor U10736 (N_10736,N_5871,N_8972);
or U10737 (N_10737,N_6133,N_7642);
or U10738 (N_10738,N_8521,N_5542);
and U10739 (N_10739,N_8235,N_5618);
nand U10740 (N_10740,N_6017,N_9032);
nor U10741 (N_10741,N_5165,N_9819);
and U10742 (N_10742,N_9802,N_8933);
nor U10743 (N_10743,N_9427,N_8255);
nand U10744 (N_10744,N_5816,N_9936);
and U10745 (N_10745,N_8284,N_5477);
or U10746 (N_10746,N_7612,N_9681);
nor U10747 (N_10747,N_6200,N_5057);
and U10748 (N_10748,N_5510,N_7755);
or U10749 (N_10749,N_8349,N_9564);
nor U10750 (N_10750,N_6619,N_5408);
or U10751 (N_10751,N_6337,N_5700);
or U10752 (N_10752,N_9470,N_9316);
nand U10753 (N_10753,N_7983,N_9558);
and U10754 (N_10754,N_5900,N_9755);
or U10755 (N_10755,N_7885,N_6109);
nor U10756 (N_10756,N_5807,N_7206);
nor U10757 (N_10757,N_9317,N_7615);
and U10758 (N_10758,N_6996,N_8540);
nand U10759 (N_10759,N_9534,N_6379);
nor U10760 (N_10760,N_5268,N_8590);
nor U10761 (N_10761,N_7697,N_7719);
nand U10762 (N_10762,N_8774,N_5002);
and U10763 (N_10763,N_5060,N_6108);
and U10764 (N_10764,N_8651,N_6489);
nor U10765 (N_10765,N_6496,N_5966);
nand U10766 (N_10766,N_7400,N_5795);
or U10767 (N_10767,N_8322,N_9057);
nor U10768 (N_10768,N_5253,N_8824);
nor U10769 (N_10769,N_6427,N_9015);
xnor U10770 (N_10770,N_6851,N_8346);
or U10771 (N_10771,N_8386,N_5566);
and U10772 (N_10772,N_9751,N_7164);
and U10773 (N_10773,N_9714,N_6900);
nand U10774 (N_10774,N_7600,N_8493);
nand U10775 (N_10775,N_5175,N_5345);
nand U10776 (N_10776,N_5449,N_6731);
nor U10777 (N_10777,N_7462,N_7176);
and U10778 (N_10778,N_5927,N_7811);
nand U10779 (N_10779,N_5587,N_7695);
nor U10780 (N_10780,N_6375,N_7866);
nand U10781 (N_10781,N_5319,N_5436);
xnor U10782 (N_10782,N_9493,N_5489);
nand U10783 (N_10783,N_8706,N_7284);
nand U10784 (N_10784,N_8498,N_7922);
nand U10785 (N_10785,N_6420,N_8583);
xor U10786 (N_10786,N_8889,N_7943);
or U10787 (N_10787,N_8881,N_8287);
nand U10788 (N_10788,N_6768,N_9097);
or U10789 (N_10789,N_8620,N_5299);
and U10790 (N_10790,N_8184,N_7918);
nand U10791 (N_10791,N_8470,N_7280);
and U10792 (N_10792,N_9395,N_9255);
and U10793 (N_10793,N_8090,N_7946);
or U10794 (N_10794,N_9339,N_5459);
nand U10795 (N_10795,N_9143,N_8779);
nor U10796 (N_10796,N_8582,N_8368);
xnor U10797 (N_10797,N_7470,N_5870);
and U10798 (N_10798,N_8953,N_5419);
or U10799 (N_10799,N_6812,N_8460);
nand U10800 (N_10800,N_6333,N_8051);
or U10801 (N_10801,N_9215,N_5666);
nand U10802 (N_10802,N_8050,N_7806);
nand U10803 (N_10803,N_5407,N_9698);
and U10804 (N_10804,N_6966,N_7734);
nand U10805 (N_10805,N_7446,N_8243);
nor U10806 (N_10806,N_9895,N_8871);
and U10807 (N_10807,N_7854,N_5347);
or U10808 (N_10808,N_9946,N_8848);
nand U10809 (N_10809,N_8290,N_8641);
nor U10810 (N_10810,N_7599,N_7050);
nor U10811 (N_10811,N_6794,N_9101);
nand U10812 (N_10812,N_5653,N_7412);
and U10813 (N_10813,N_7012,N_5731);
and U10814 (N_10814,N_5284,N_8732);
nand U10815 (N_10815,N_6443,N_6513);
or U10816 (N_10816,N_5867,N_7941);
and U10817 (N_10817,N_9565,N_5313);
or U10818 (N_10818,N_5570,N_8151);
nor U10819 (N_10819,N_9103,N_8486);
or U10820 (N_10820,N_9596,N_6818);
xnor U10821 (N_10821,N_7559,N_9440);
and U10822 (N_10822,N_6650,N_9767);
and U10823 (N_10823,N_9843,N_7392);
and U10824 (N_10824,N_5226,N_8808);
nor U10825 (N_10825,N_6558,N_7693);
and U10826 (N_10826,N_7186,N_8573);
and U10827 (N_10827,N_7844,N_5540);
or U10828 (N_10828,N_7379,N_9858);
nand U10829 (N_10829,N_7144,N_8500);
and U10830 (N_10830,N_9707,N_9551);
and U10831 (N_10831,N_9162,N_5948);
xor U10832 (N_10832,N_9127,N_5236);
xnor U10833 (N_10833,N_5698,N_8997);
xor U10834 (N_10834,N_5598,N_5013);
xor U10835 (N_10835,N_6627,N_6350);
or U10836 (N_10836,N_5768,N_7986);
and U10837 (N_10837,N_5800,N_6494);
nor U10838 (N_10838,N_6390,N_8826);
nand U10839 (N_10839,N_7256,N_8975);
or U10840 (N_10840,N_8062,N_6590);
xnor U10841 (N_10841,N_5535,N_9545);
nand U10842 (N_10842,N_9000,N_8886);
or U10843 (N_10843,N_9415,N_6303);
or U10844 (N_10844,N_6291,N_6466);
or U10845 (N_10845,N_5445,N_8329);
xnor U10846 (N_10846,N_7128,N_6155);
nand U10847 (N_10847,N_7422,N_9416);
or U10848 (N_10848,N_8817,N_5003);
nor U10849 (N_10849,N_7751,N_8723);
and U10850 (N_10850,N_7250,N_6461);
and U10851 (N_10851,N_9733,N_5192);
nand U10852 (N_10852,N_8952,N_5157);
or U10853 (N_10853,N_7813,N_7029);
xnor U10854 (N_10854,N_7381,N_6526);
and U10855 (N_10855,N_7211,N_5392);
and U10856 (N_10856,N_5108,N_7829);
and U10857 (N_10857,N_6782,N_6113);
and U10858 (N_10858,N_6943,N_9069);
and U10859 (N_10859,N_8616,N_8954);
nor U10860 (N_10860,N_8757,N_7679);
or U10861 (N_10861,N_9726,N_7151);
or U10862 (N_10862,N_7546,N_5164);
or U10863 (N_10863,N_8636,N_8676);
nor U10864 (N_10864,N_6852,N_7966);
or U10865 (N_10865,N_7313,N_6822);
and U10866 (N_10866,N_6955,N_7608);
nand U10867 (N_10867,N_6980,N_7948);
and U10868 (N_10868,N_7233,N_8709);
and U10869 (N_10869,N_7908,N_7155);
and U10870 (N_10870,N_9909,N_5206);
and U10871 (N_10871,N_9396,N_8744);
or U10872 (N_10872,N_7419,N_9854);
or U10873 (N_10873,N_5322,N_6994);
nor U10874 (N_10874,N_6148,N_6126);
nand U10875 (N_10875,N_8295,N_5982);
and U10876 (N_10876,N_6810,N_6525);
xor U10877 (N_10877,N_6577,N_6617);
nand U10878 (N_10878,N_7977,N_5398);
and U10879 (N_10879,N_5854,N_7274);
nor U10880 (N_10880,N_9208,N_9467);
or U10881 (N_10881,N_6062,N_8519);
nand U10882 (N_10882,N_6787,N_9260);
or U10883 (N_10883,N_5280,N_5292);
nand U10884 (N_10884,N_6100,N_9690);
and U10885 (N_10885,N_7062,N_8937);
or U10886 (N_10886,N_6595,N_8253);
and U10887 (N_10887,N_7465,N_8503);
and U10888 (N_10888,N_5017,N_5250);
and U10889 (N_10889,N_6823,N_6896);
or U10890 (N_10890,N_9139,N_9635);
or U10891 (N_10891,N_9457,N_5205);
nor U10892 (N_10892,N_7174,N_5277);
nand U10893 (N_10893,N_7617,N_5732);
xor U10894 (N_10894,N_5572,N_9697);
nand U10895 (N_10895,N_5930,N_9235);
nor U10896 (N_10896,N_5562,N_7851);
nor U10897 (N_10897,N_5610,N_8506);
nor U10898 (N_10898,N_8144,N_8994);
and U10899 (N_10899,N_8461,N_5147);
and U10900 (N_10900,N_5989,N_6610);
nand U10901 (N_10901,N_5018,N_6874);
and U10902 (N_10902,N_5642,N_5554);
nand U10903 (N_10903,N_5042,N_7475);
nand U10904 (N_10904,N_7631,N_6152);
or U10905 (N_10905,N_9945,N_8296);
and U10906 (N_10906,N_6793,N_5229);
or U10907 (N_10907,N_8735,N_8138);
nor U10908 (N_10908,N_7429,N_9045);
nand U10909 (N_10909,N_6160,N_9476);
and U10910 (N_10910,N_5929,N_9332);
and U10911 (N_10911,N_6579,N_6416);
and U10912 (N_10912,N_9058,N_5895);
nand U10913 (N_10913,N_7396,N_9993);
and U10914 (N_10914,N_5210,N_7792);
nor U10915 (N_10915,N_9405,N_5023);
nor U10916 (N_10916,N_5467,N_5420);
nand U10917 (N_10917,N_9670,N_7439);
and U10918 (N_10918,N_7220,N_6284);
nor U10919 (N_10919,N_6989,N_7935);
nand U10920 (N_10920,N_6824,N_5830);
nor U10921 (N_10921,N_6499,N_8268);
nor U10922 (N_10922,N_5987,N_7992);
or U10923 (N_10923,N_6722,N_8011);
and U10924 (N_10924,N_6381,N_8610);
or U10925 (N_10925,N_8266,N_6164);
or U10926 (N_10926,N_5466,N_6564);
and U10927 (N_10927,N_7754,N_5158);
and U10928 (N_10928,N_7177,N_5486);
nor U10929 (N_10929,N_5545,N_7657);
or U10930 (N_10930,N_7730,N_8398);
nand U10931 (N_10931,N_7537,N_5144);
and U10932 (N_10932,N_7102,N_9888);
nand U10933 (N_10933,N_9696,N_9423);
and U10934 (N_10934,N_9413,N_9962);
nand U10935 (N_10935,N_5971,N_5040);
or U10936 (N_10936,N_5086,N_8476);
nand U10937 (N_10937,N_7785,N_8438);
xor U10938 (N_10938,N_9378,N_7594);
nor U10939 (N_10939,N_9809,N_9763);
xor U10940 (N_10940,N_8173,N_7496);
xor U10941 (N_10941,N_6424,N_7771);
or U10942 (N_10942,N_7116,N_6912);
nor U10943 (N_10943,N_5446,N_8910);
nor U10944 (N_10944,N_6469,N_8512);
nor U10945 (N_10945,N_9957,N_8878);
and U10946 (N_10946,N_7410,N_8405);
nor U10947 (N_10947,N_8629,N_9017);
and U10948 (N_10948,N_9318,N_6454);
nor U10949 (N_10949,N_7748,N_5576);
nor U10950 (N_10950,N_7358,N_9327);
or U10951 (N_10951,N_6739,N_9571);
nor U10952 (N_10952,N_9262,N_7773);
and U10953 (N_10953,N_6483,N_5520);
or U10954 (N_10954,N_6308,N_5659);
nor U10955 (N_10955,N_5211,N_5468);
nand U10956 (N_10956,N_5623,N_7374);
or U10957 (N_10957,N_5325,N_8206);
nand U10958 (N_10958,N_8962,N_6403);
or U10959 (N_10959,N_6161,N_6191);
nand U10960 (N_10960,N_5883,N_8969);
and U10961 (N_10961,N_7411,N_9609);
or U10962 (N_10962,N_6176,N_6553);
xor U10963 (N_10963,N_6883,N_6043);
or U10964 (N_10964,N_6478,N_6934);
nor U10965 (N_10965,N_7271,N_9599);
nor U10966 (N_10966,N_9683,N_7273);
nor U10967 (N_10967,N_5038,N_6452);
nand U10968 (N_10968,N_5850,N_9897);
nor U10969 (N_10969,N_5151,N_6330);
nor U10970 (N_10970,N_6854,N_7721);
or U10971 (N_10971,N_5845,N_5304);
or U10972 (N_10972,N_7123,N_6877);
nor U10973 (N_10973,N_8731,N_7290);
nor U10974 (N_10974,N_9793,N_9677);
and U10975 (N_10975,N_8530,N_8434);
nand U10976 (N_10976,N_6329,N_7361);
nor U10977 (N_10977,N_6819,N_8932);
nor U10978 (N_10978,N_6184,N_9744);
and U10979 (N_10979,N_9794,N_5215);
or U10980 (N_10980,N_7602,N_7910);
or U10981 (N_10981,N_6448,N_9625);
nor U10982 (N_10982,N_9815,N_7930);
nor U10983 (N_10983,N_9124,N_9354);
nand U10984 (N_10984,N_8558,N_7516);
nand U10985 (N_10985,N_7067,N_7112);
or U10986 (N_10986,N_7199,N_8003);
and U10987 (N_10987,N_8376,N_6353);
xnor U10988 (N_10988,N_9121,N_8331);
nor U10989 (N_10989,N_9359,N_5557);
and U10990 (N_10990,N_9832,N_8899);
or U10991 (N_10991,N_7453,N_9232);
and U10992 (N_10992,N_5208,N_6220);
and U10993 (N_10993,N_6305,N_5170);
and U10994 (N_10994,N_6315,N_8379);
nand U10995 (N_10995,N_5954,N_5771);
nor U10996 (N_10996,N_8646,N_9369);
nor U10997 (N_10997,N_5522,N_6531);
or U10998 (N_10998,N_6397,N_7621);
or U10999 (N_10999,N_6071,N_8393);
nand U11000 (N_11000,N_8185,N_8747);
nor U11001 (N_11001,N_9046,N_8728);
nor U11002 (N_11002,N_7529,N_7777);
nor U11003 (N_11003,N_8402,N_6723);
and U11004 (N_11004,N_9871,N_8836);
nand U11005 (N_11005,N_8857,N_9652);
nand U11006 (N_11006,N_8248,N_5111);
nor U11007 (N_11007,N_8096,N_7363);
and U11008 (N_11008,N_5138,N_7404);
nor U11009 (N_11009,N_6831,N_9322);
nand U11010 (N_11010,N_6897,N_9429);
or U11011 (N_11011,N_6799,N_6535);
nand U11012 (N_11012,N_7015,N_7704);
nor U11013 (N_11013,N_9238,N_7604);
or U11014 (N_11014,N_8586,N_9602);
or U11015 (N_11015,N_8464,N_5102);
and U11016 (N_11016,N_9439,N_6262);
nand U11017 (N_11017,N_5836,N_9846);
or U11018 (N_11018,N_6181,N_6282);
nand U11019 (N_11019,N_8361,N_6373);
nor U11020 (N_11020,N_9640,N_7857);
nand U11021 (N_11021,N_7006,N_8944);
and U11022 (N_11022,N_5777,N_6616);
nor U11023 (N_11023,N_5829,N_8482);
nor U11024 (N_11024,N_9307,N_6764);
and U11025 (N_11025,N_9270,N_7218);
nor U11026 (N_11026,N_7982,N_6572);
nor U11027 (N_11027,N_7971,N_6811);
nor U11028 (N_11028,N_7497,N_7134);
nor U11029 (N_11029,N_9865,N_6455);
nand U11030 (N_11030,N_8258,N_7002);
and U11031 (N_11031,N_8525,N_7382);
nand U11032 (N_11032,N_5049,N_5508);
nand U11033 (N_11033,N_6709,N_6743);
and U11034 (N_11034,N_9973,N_8859);
nand U11035 (N_11035,N_8152,N_5109);
or U11036 (N_11036,N_8839,N_8637);
and U11037 (N_11037,N_5574,N_9365);
and U11038 (N_11038,N_5154,N_5649);
and U11039 (N_11039,N_5025,N_7809);
nor U11040 (N_11040,N_9161,N_5711);
nand U11041 (N_11041,N_5438,N_9249);
and U11042 (N_11042,N_6302,N_9292);
nor U11043 (N_11043,N_5835,N_7778);
nand U11044 (N_11044,N_8518,N_7376);
nor U11045 (N_11045,N_5455,N_6052);
or U11046 (N_11046,N_7425,N_8123);
xnor U11047 (N_11047,N_9449,N_8922);
and U11048 (N_11048,N_8901,N_6771);
nand U11049 (N_11049,N_9471,N_8231);
and U11050 (N_11050,N_8452,N_5359);
or U11051 (N_11051,N_6930,N_9469);
nand U11052 (N_11052,N_9842,N_7539);
nor U11053 (N_11053,N_6114,N_6630);
nand U11054 (N_11054,N_9933,N_5183);
nor U11055 (N_11055,N_6653,N_7119);
nand U11056 (N_11056,N_8092,N_8644);
and U11057 (N_11057,N_9263,N_9001);
nor U11058 (N_11058,N_5198,N_5641);
nor U11059 (N_11059,N_5218,N_9863);
and U11060 (N_11060,N_5342,N_6210);
and U11061 (N_11061,N_8189,N_9658);
xor U11062 (N_11062,N_6733,N_7214);
xnor U11063 (N_11063,N_8959,N_7423);
or U11064 (N_11064,N_6608,N_6033);
nand U11065 (N_11065,N_9499,N_5099);
or U11066 (N_11066,N_7406,N_5317);
nor U11067 (N_11067,N_8958,N_5130);
or U11068 (N_11068,N_9958,N_7107);
and U11069 (N_11069,N_8681,N_9906);
nor U11070 (N_11070,N_6385,N_6870);
nand U11071 (N_11071,N_5602,N_8654);
and U11072 (N_11072,N_6079,N_8042);
nand U11073 (N_11073,N_8541,N_6280);
or U11074 (N_11074,N_5262,N_7818);
nand U11075 (N_11075,N_6189,N_8941);
nor U11076 (N_11076,N_5794,N_9932);
and U11077 (N_11077,N_9461,N_9436);
and U11078 (N_11078,N_7793,N_5386);
or U11079 (N_11079,N_5308,N_8775);
or U11080 (N_11080,N_7799,N_6103);
and U11081 (N_11081,N_5339,N_7487);
nor U11082 (N_11082,N_8707,N_8761);
nor U11083 (N_11083,N_6703,N_5473);
nand U11084 (N_11084,N_9776,N_8909);
nor U11085 (N_11085,N_6864,N_8745);
nor U11086 (N_11086,N_6259,N_7262);
nor U11087 (N_11087,N_6919,N_8608);
or U11088 (N_11088,N_8279,N_6738);
or U11089 (N_11089,N_6446,N_9621);
xnor U11090 (N_11090,N_7110,N_5921);
xnor U11091 (N_11091,N_9496,N_9414);
and U11092 (N_11092,N_7011,N_6680);
or U11093 (N_11093,N_8508,N_5335);
and U11094 (N_11094,N_7690,N_8698);
or U11095 (N_11095,N_9141,N_8847);
or U11096 (N_11096,N_6178,N_7660);
or U11097 (N_11097,N_5254,N_5861);
nor U11098 (N_11098,N_7576,N_9738);
nor U11099 (N_11099,N_8327,N_9820);
and U11100 (N_11100,N_6368,N_7810);
xnor U11101 (N_11101,N_8893,N_5382);
or U11102 (N_11102,N_9218,N_8765);
nor U11103 (N_11103,N_7146,N_8357);
nand U11104 (N_11104,N_5329,N_6686);
nand U11105 (N_11105,N_8515,N_8018);
nor U11106 (N_11106,N_7920,N_6521);
and U11107 (N_11107,N_7531,N_7682);
nor U11108 (N_11108,N_8169,N_9202);
nand U11109 (N_11109,N_9781,N_6187);
and U11110 (N_11110,N_5941,N_5783);
nand U11111 (N_11111,N_8485,N_8221);
xnor U11112 (N_11112,N_9514,N_8880);
and U11113 (N_11113,N_9503,N_6503);
nor U11114 (N_11114,N_7217,N_6506);
nor U11115 (N_11115,N_7942,N_5852);
or U11116 (N_11116,N_6186,N_7348);
xor U11117 (N_11117,N_6551,N_5863);
xnor U11118 (N_11118,N_5956,N_7921);
or U11119 (N_11119,N_5901,N_7309);
and U11120 (N_11120,N_8684,N_6646);
or U11121 (N_11121,N_6150,N_5333);
nand U11122 (N_11122,N_6044,N_7565);
and U11123 (N_11123,N_5235,N_6977);
and U11124 (N_11124,N_7241,N_6159);
and U11125 (N_11125,N_7782,N_9220);
and U11126 (N_11126,N_6785,N_8680);
xor U11127 (N_11127,N_7590,N_8276);
or U11128 (N_11128,N_5075,N_6589);
or U11129 (N_11129,N_9156,N_6135);
nor U11130 (N_11130,N_5821,N_5318);
nor U11131 (N_11131,N_7454,N_7728);
nor U11132 (N_11132,N_6868,N_9245);
or U11133 (N_11133,N_8562,N_9929);
nand U11134 (N_11134,N_9959,N_9998);
or U11135 (N_11135,N_7630,N_9087);
nor U11136 (N_11136,N_8566,N_6163);
xor U11137 (N_11137,N_6601,N_5500);
and U11138 (N_11138,N_5397,N_9234);
nand U11139 (N_11139,N_6301,N_7040);
xnor U11140 (N_11140,N_6973,N_7666);
nand U11141 (N_11141,N_5565,N_9256);
and U11142 (N_11142,N_9334,N_5431);
nand U11143 (N_11143,N_7459,N_5194);
nor U11144 (N_11144,N_5848,N_6288);
and U11145 (N_11145,N_5813,N_9187);
and U11146 (N_11146,N_6736,N_6068);
nand U11147 (N_11147,N_9550,N_5650);
nor U11148 (N_11148,N_5255,N_7916);
and U11149 (N_11149,N_9295,N_6289);
xnor U11150 (N_11150,N_9089,N_9732);
or U11151 (N_11151,N_5823,N_9702);
and U11152 (N_11152,N_8694,N_6755);
or U11153 (N_11153,N_5478,N_5798);
nor U11154 (N_11154,N_7692,N_7551);
nand U11155 (N_11155,N_6221,N_7812);
or U11156 (N_11156,N_7143,N_7628);
nor U11157 (N_11157,N_8236,N_5539);
or U11158 (N_11158,N_5736,N_5880);
nor U11159 (N_11159,N_9917,N_6277);
or U11160 (N_11160,N_8364,N_9221);
or U11161 (N_11161,N_9258,N_8422);
nor U11162 (N_11162,N_6422,N_9533);
nor U11163 (N_11163,N_8021,N_5719);
nand U11164 (N_11164,N_9991,N_5341);
or U11165 (N_11165,N_6882,N_5155);
nand U11166 (N_11166,N_8869,N_6225);
or U11167 (N_11167,N_6772,N_9071);
xnor U11168 (N_11168,N_9280,N_7263);
or U11169 (N_11169,N_5869,N_7223);
and U11170 (N_11170,N_8466,N_7623);
nand U11171 (N_11171,N_8655,N_9233);
and U11172 (N_11172,N_5627,N_8196);
or U11173 (N_11173,N_9508,N_7879);
nor U11174 (N_11174,N_7687,N_6195);
and U11175 (N_11175,N_6065,N_6344);
and U11176 (N_11176,N_5078,N_6903);
and U11177 (N_11177,N_7506,N_7749);
nand U11178 (N_11178,N_8286,N_6051);
and U11179 (N_11179,N_6351,N_8401);
nand U11180 (N_11180,N_6944,N_8987);
and U11181 (N_11181,N_7840,N_7075);
nor U11182 (N_11182,N_7261,N_7598);
xor U11183 (N_11183,N_8729,N_8293);
xnor U11184 (N_11184,N_5450,N_9079);
xor U11185 (N_11185,N_5447,N_5527);
nand U11186 (N_11186,N_8587,N_5788);
or U11187 (N_11187,N_9371,N_6855);
and U11188 (N_11188,N_8272,N_5931);
nand U11189 (N_11189,N_6663,N_8125);
nand U11190 (N_11190,N_6059,N_6182);
and U11191 (N_11191,N_9606,N_6891);
or U11192 (N_11192,N_6123,N_7098);
or U11193 (N_11193,N_9745,N_6737);
nor U11194 (N_11194,N_6384,N_8524);
or U11195 (N_11195,N_8782,N_9025);
nand U11196 (N_11196,N_6074,N_6322);
or U11197 (N_11197,N_8391,N_8903);
or U11198 (N_11198,N_9110,N_8070);
and U11199 (N_11199,N_6342,N_7037);
nand U11200 (N_11200,N_6791,N_7827);
nand U11201 (N_11201,N_9125,N_9978);
and U11202 (N_11202,N_8009,N_5067);
nand U11203 (N_11203,N_8044,N_6382);
or U11204 (N_11204,N_5664,N_5675);
and U11205 (N_11205,N_6798,N_7669);
and U11206 (N_11206,N_5291,N_6769);
or U11207 (N_11207,N_9345,N_5371);
and U11208 (N_11208,N_5356,N_6131);
xor U11209 (N_11209,N_9655,N_8007);
xnor U11210 (N_11210,N_6408,N_9939);
nand U11211 (N_11211,N_6905,N_5297);
xnor U11212 (N_11212,N_9822,N_7183);
and U11213 (N_11213,N_5681,N_9213);
nor U11214 (N_11214,N_5691,N_9081);
nor U11215 (N_11215,N_6486,N_5063);
or U11216 (N_11216,N_9223,N_9833);
or U11217 (N_11217,N_6659,N_7350);
and U11218 (N_11218,N_7691,N_6895);
and U11219 (N_11219,N_5044,N_8321);
nand U11220 (N_11220,N_9196,N_5134);
and U11221 (N_11221,N_9892,N_8160);
and U11222 (N_11222,N_9553,N_5946);
nor U11223 (N_11223,N_7318,N_5561);
nor U11224 (N_11224,N_5842,N_6740);
and U11225 (N_11225,N_6649,N_5974);
nor U11226 (N_11226,N_5050,N_6981);
and U11227 (N_11227,N_5599,N_9885);
nor U11228 (N_11228,N_8758,N_6985);
nand U11229 (N_11229,N_6023,N_8492);
nand U11230 (N_11230,N_5721,N_8095);
and U11231 (N_11231,N_9319,N_8720);
or U11232 (N_11232,N_6614,N_8154);
or U11233 (N_11233,N_9356,N_5662);
and U11234 (N_11234,N_7893,N_5168);
nand U11235 (N_11235,N_9960,N_7726);
nor U11236 (N_11236,N_8102,N_6599);
nand U11237 (N_11237,N_9666,N_9777);
and U11238 (N_11238,N_7663,N_5751);
and U11239 (N_11239,N_9504,N_7572);
nor U11240 (N_11240,N_8328,N_6642);
and U11241 (N_11241,N_8794,N_7996);
or U11242 (N_11242,N_9647,N_9014);
nand U11243 (N_11243,N_7149,N_5809);
nand U11244 (N_11244,N_9304,N_5237);
nor U11245 (N_11245,N_7317,N_7184);
and U11246 (N_11246,N_8127,N_6268);
nor U11247 (N_11247,N_9731,N_7013);
and U11248 (N_11248,N_6805,N_5705);
and U11249 (N_11249,N_8489,N_9484);
or U11250 (N_11250,N_9814,N_8640);
or U11251 (N_11251,N_7775,N_7828);
or U11252 (N_11252,N_5963,N_7368);
or U11253 (N_11253,N_5792,N_9801);
nand U11254 (N_11254,N_9400,N_7308);
nor U11255 (N_11255,N_9770,N_5780);
or U11256 (N_11256,N_7869,N_9490);
or U11257 (N_11257,N_8133,N_8455);
nand U11258 (N_11258,N_5312,N_8653);
or U11259 (N_11259,N_8165,N_7287);
xnor U11260 (N_11260,N_6615,N_9115);
and U11261 (N_11261,N_8412,N_8509);
and U11262 (N_11262,N_7999,N_5865);
nor U11263 (N_11263,N_6336,N_5746);
and U11264 (N_11264,N_8986,N_6183);
xnor U11265 (N_11265,N_6714,N_9225);
nor U11266 (N_11266,N_8844,N_6957);
nor U11267 (N_11267,N_6145,N_7557);
nand U11268 (N_11268,N_6036,N_9426);
and U11269 (N_11269,N_6299,N_5276);
nand U11270 (N_11270,N_9433,N_7732);
nand U11271 (N_11271,N_9783,N_8115);
nor U11272 (N_11272,N_7377,N_7503);
or U11273 (N_11273,N_7147,N_6717);
nand U11274 (N_11274,N_6444,N_9368);
nor U11275 (N_11275,N_7389,N_6362);
or U11276 (N_11276,N_5986,N_9398);
xnor U11277 (N_11277,N_8264,N_9182);
or U11278 (N_11278,N_6436,N_8270);
nand U11279 (N_11279,N_9016,N_9598);
nand U11280 (N_11280,N_9575,N_5483);
or U11281 (N_11281,N_6168,N_5997);
or U11282 (N_11282,N_6605,N_5912);
and U11283 (N_11283,N_7093,N_5667);
nor U11284 (N_11284,N_6005,N_6842);
or U11285 (N_11285,N_7847,N_8325);
nand U11286 (N_11286,N_5841,N_7821);
and U11287 (N_11287,N_9747,N_8427);
nand U11288 (N_11288,N_9782,N_8780);
nand U11289 (N_11289,N_6726,N_6214);
nand U11290 (N_11290,N_8755,N_9883);
and U11291 (N_11291,N_5090,N_9008);
xnor U11292 (N_11292,N_5225,N_5635);
xor U11293 (N_11293,N_8347,N_5693);
or U11294 (N_11294,N_5043,N_8591);
and U11295 (N_11295,N_6127,N_9882);
nor U11296 (N_11296,N_8904,N_7074);
nand U11297 (N_11297,N_5191,N_8832);
nand U11298 (N_11298,N_7923,N_7048);
nor U11299 (N_11299,N_6124,N_7354);
or U11300 (N_11300,N_6346,N_5957);
nand U11301 (N_11301,N_7979,N_8299);
nand U11302 (N_11302,N_9811,N_5507);
xnor U11303 (N_11303,N_9388,N_7508);
nand U11304 (N_11304,N_6986,N_8677);
nor U11305 (N_11305,N_9331,N_5766);
and U11306 (N_11306,N_9675,N_6766);
nand U11307 (N_11307,N_9664,N_9095);
or U11308 (N_11308,N_9555,N_5350);
nand U11309 (N_11309,N_9191,N_6848);
and U11310 (N_11310,N_8149,N_9216);
and U11311 (N_11311,N_9333,N_5665);
or U11312 (N_11312,N_8058,N_7460);
and U11313 (N_11313,N_6162,N_7909);
or U11314 (N_11314,N_7808,N_6027);
and U11315 (N_11315,N_7906,N_9244);
nor U11316 (N_11316,N_6846,N_7169);
and U11317 (N_11317,N_5781,N_5928);
nor U11318 (N_11318,N_9241,N_6295);
or U11319 (N_11319,N_9997,N_5630);
or U11320 (N_11320,N_9324,N_7703);
nand U11321 (N_11321,N_6859,N_5481);
nor U11322 (N_11322,N_8159,N_5560);
or U11323 (N_11323,N_6936,N_6493);
and U11324 (N_11324,N_5752,N_5311);
or U11325 (N_11325,N_8426,N_7912);
nand U11326 (N_11326,N_6872,N_7545);
nor U11327 (N_11327,N_9531,N_8229);
or U11328 (N_11328,N_6076,N_5009);
and U11329 (N_11329,N_6952,N_5657);
nand U11330 (N_11330,N_9211,N_6689);
nor U11331 (N_11331,N_7035,N_6211);
nor U11332 (N_11332,N_9346,N_9100);
xor U11333 (N_11333,N_7257,N_7278);
nor U11334 (N_11334,N_8920,N_6203);
xor U11335 (N_11335,N_8353,N_8047);
and U11336 (N_11336,N_9617,N_7581);
nor U11337 (N_11337,N_6205,N_9869);
nor U11338 (N_11338,N_8625,N_8035);
or U11339 (N_11339,N_9588,N_6817);
nor U11340 (N_11340,N_5958,N_6171);
or U11341 (N_11341,N_9839,N_5640);
nor U11342 (N_11342,N_8569,N_7547);
and U11343 (N_11343,N_6965,N_7984);
or U11344 (N_11344,N_7950,N_5679);
nand U11345 (N_11345,N_9321,N_8453);
and U11346 (N_11346,N_9468,N_9091);
or U11347 (N_11347,N_5073,N_7889);
xnor U11348 (N_11348,N_7228,N_7541);
and U11349 (N_11349,N_9711,N_5200);
and U11350 (N_11350,N_8861,N_7148);
and U11351 (N_11351,N_9007,N_9673);
or U11352 (N_11352,N_9511,N_7683);
nand U11353 (N_11353,N_9033,N_9450);
and U11354 (N_11354,N_6138,N_9341);
nand U11355 (N_11355,N_7817,N_6327);
nand U11356 (N_11356,N_8209,N_6192);
xor U11357 (N_11357,N_9724,N_9023);
nor U11358 (N_11358,N_5101,N_9582);
nand U11359 (N_11359,N_7949,N_9771);
nor U11360 (N_11360,N_5652,N_5425);
and U11361 (N_11361,N_9391,N_6979);
nand U11362 (N_11362,N_9955,N_6122);
nand U11363 (N_11363,N_6470,N_5337);
nor U11364 (N_11364,N_7676,N_7725);
nand U11365 (N_11365,N_7622,N_5055);
nand U11366 (N_11366,N_7286,N_9447);
and U11367 (N_11367,N_7434,N_8991);
or U11368 (N_11368,N_8700,N_8703);
nand U11369 (N_11369,N_6047,N_6861);
nand U11370 (N_11370,N_8599,N_7959);
xnor U11371 (N_11371,N_7670,N_7187);
or U11372 (N_11372,N_6255,N_6801);
nand U11373 (N_11373,N_8425,N_8549);
nand U11374 (N_11374,N_7560,N_8789);
nand U11375 (N_11375,N_6252,N_9898);
nor U11376 (N_11376,N_8084,N_6414);
nor U11377 (N_11377,N_9172,N_9084);
nand U11378 (N_11378,N_8077,N_7212);
or U11379 (N_11379,N_7610,N_8305);
and U11380 (N_11380,N_9969,N_6543);
or U11381 (N_11381,N_5968,N_7850);
or U11382 (N_11382,N_5252,N_7472);
xnor U11383 (N_11383,N_8834,N_9927);
and U11384 (N_11384,N_6243,N_9521);
and U11385 (N_11385,N_7270,N_5797);
and U11386 (N_11386,N_6266,N_5601);
nor U11387 (N_11387,N_6212,N_5490);
and U11388 (N_11388,N_8103,N_9592);
nand U11389 (N_11389,N_5316,N_5874);
or U11390 (N_11390,N_5056,N_5796);
nor U11391 (N_11391,N_5103,N_9174);
nand U11392 (N_11392,N_8323,N_8862);
nand U11393 (N_11393,N_5492,N_6413);
or U11394 (N_11394,N_8897,N_9222);
nand U11395 (N_11395,N_5749,N_9515);
nor U11396 (N_11396,N_8618,N_7372);
nand U11397 (N_11397,N_5550,N_6316);
and U11398 (N_11398,N_5787,N_7388);
nor U11399 (N_11399,N_7905,N_8858);
nor U11400 (N_11400,N_8797,N_8163);
and U11401 (N_11401,N_5515,N_8337);
and U11402 (N_11402,N_6298,N_5395);
xor U11403 (N_11403,N_9812,N_6018);
nand U11404 (N_11404,N_9432,N_6643);
nand U11405 (N_11405,N_9950,N_8089);
or U11406 (N_11406,N_9062,N_8314);
nor U11407 (N_11407,N_8396,N_7014);
nor U11408 (N_11408,N_5505,N_7859);
nor U11409 (N_11409,N_8883,N_6945);
nand U11410 (N_11410,N_8609,N_6964);
nor U11411 (N_11411,N_7008,N_9485);
nand U11412 (N_11412,N_8283,N_7087);
or U11413 (N_11413,N_8752,N_7926);
and U11414 (N_11414,N_5095,N_7634);
xnor U11415 (N_11415,N_8915,N_6458);
nand U11416 (N_11416,N_8601,N_9438);
nor U11417 (N_11417,N_7080,N_7655);
or U11418 (N_11418,N_6666,N_5638);
nor U11419 (N_11419,N_6622,N_5181);
and U11420 (N_11420,N_9646,N_7295);
nor U11421 (N_11421,N_6153,N_5234);
nand U11422 (N_11422,N_9526,N_8567);
nor U11423 (N_11423,N_8298,N_5785);
nor U11424 (N_11424,N_6463,N_5256);
nand U11425 (N_11425,N_9070,N_8429);
or U11426 (N_11426,N_5710,N_9736);
or U11427 (N_11427,N_8065,N_5917);
or U11428 (N_11428,N_9778,N_8827);
or U11429 (N_11429,N_6460,N_6625);
xnor U11430 (N_11430,N_6644,N_5844);
and U11431 (N_11431,N_8628,N_9676);
nand U11432 (N_11432,N_7672,N_6120);
nor U11433 (N_11433,N_8421,N_7705);
nand U11434 (N_11434,N_6137,N_7251);
nand U11435 (N_11435,N_7891,N_6661);
nor U11436 (N_11436,N_9169,N_8022);
and U11437 (N_11437,N_9903,N_9451);
nor U11438 (N_11438,N_6826,N_6248);
nand U11439 (N_11439,N_5113,N_5270);
xor U11440 (N_11440,N_5189,N_7383);
nand U11441 (N_11441,N_9297,N_8966);
and U11442 (N_11442,N_8984,N_9709);
nor U11443 (N_11443,N_9209,N_5953);
and U11444 (N_11444,N_5480,N_5428);
nand U11445 (N_11445,N_9052,N_5589);
xor U11446 (N_11446,N_8158,N_6857);
nor U11447 (N_11447,N_7315,N_8025);
and U11448 (N_11448,N_5361,N_9837);
or U11449 (N_11449,N_5019,N_8798);
or U11450 (N_11450,N_6498,N_6202);
or U11451 (N_11451,N_5939,N_9951);
and U11452 (N_11452,N_9031,N_7259);
or U11453 (N_11453,N_9298,N_8748);
and U11454 (N_11454,N_9320,N_5612);
nor U11455 (N_11455,N_6487,N_6488);
nor U11456 (N_11456,N_8430,N_8403);
and U11457 (N_11457,N_9954,N_5264);
or U11458 (N_11458,N_9769,N_7686);
nand U11459 (N_11459,N_9930,N_5364);
and U11460 (N_11460,N_8537,N_9076);
or U11461 (N_11461,N_6227,N_6840);
nor U11462 (N_11462,N_6400,N_7055);
or U11463 (N_11463,N_7299,N_6911);
and U11464 (N_11464,N_6423,N_9510);
nand U11465 (N_11465,N_7026,N_6971);
and U11466 (N_11466,N_7333,N_5323);
and U11467 (N_11467,N_7077,N_9758);
and U11468 (N_11468,N_8116,N_7043);
or U11469 (N_11469,N_9310,N_7126);
or U11470 (N_11470,N_5444,N_8418);
or U11471 (N_11471,N_6419,N_5227);
or U11472 (N_11472,N_7279,N_9942);
xnor U11473 (N_11473,N_6609,N_5647);
xor U11474 (N_11474,N_9184,N_6209);
and U11475 (N_11475,N_8483,N_7255);
nand U11476 (N_11476,N_6583,N_6010);
or U11477 (N_11477,N_9059,N_5219);
nand U11478 (N_11478,N_7940,N_8013);
or U11479 (N_11479,N_8849,N_6635);
nor U11480 (N_11480,N_9003,N_7324);
or U11481 (N_11481,N_6129,N_9362);
nand U11482 (N_11482,N_9009,N_5925);
nand U11483 (N_11483,N_7387,N_7482);
or U11484 (N_11484,N_5538,N_5584);
xor U11485 (N_11485,N_5839,N_5855);
and U11486 (N_11486,N_5123,N_5089);
or U11487 (N_11487,N_9825,N_6007);
and U11488 (N_11488,N_5943,N_7903);
or U11489 (N_11489,N_7654,N_8333);
or U11490 (N_11490,N_6507,N_8692);
nand U11491 (N_11491,N_9524,N_7249);
and U11492 (N_11492,N_6371,N_7579);
nor U11493 (N_11493,N_6807,N_9104);
and U11494 (N_11494,N_6029,N_6002);
or U11495 (N_11495,N_9913,N_9632);
nor U11496 (N_11496,N_7969,N_7555);
nand U11497 (N_11497,N_8634,N_6398);
nor U11498 (N_11498,N_8068,N_6961);
nand U11499 (N_11499,N_8162,N_7711);
nand U11500 (N_11500,N_9275,N_7213);
nor U11501 (N_11501,N_9556,N_6655);
nor U11502 (N_11502,N_6922,N_7480);
nand U11503 (N_11503,N_6958,N_5782);
nand U11504 (N_11504,N_5169,N_9611);
nand U11505 (N_11505,N_6656,N_9305);
xnor U11506 (N_11506,N_5826,N_7958);
nor U11507 (N_11507,N_8645,N_6415);
or U11508 (N_11508,N_9194,N_5772);
and U11509 (N_11509,N_8141,N_7843);
nor U11510 (N_11510,N_5456,N_7988);
nor U11511 (N_11511,N_8071,N_6750);
nand U11512 (N_11512,N_9401,N_7562);
or U11513 (N_11513,N_5977,N_8998);
and U11514 (N_11514,N_9407,N_9689);
nor U11515 (N_11515,N_6167,N_7990);
nand U11516 (N_11516,N_8214,N_8778);
and U11517 (N_11517,N_9372,N_9483);
xnor U11518 (N_11518,N_7421,N_7838);
or U11519 (N_11519,N_8526,N_6951);
and U11520 (N_11520,N_5471,N_7215);
and U11521 (N_11521,N_9230,N_5294);
and U11522 (N_11522,N_7688,N_8080);
nand U11523 (N_11523,N_8548,N_6473);
nand U11524 (N_11524,N_6520,N_7849);
nand U11525 (N_11525,N_7972,N_7824);
nor U11526 (N_11526,N_8202,N_6232);
or U11527 (N_11527,N_7455,N_6015);
or U11528 (N_11528,N_5801,N_9144);
nand U11529 (N_11529,N_6037,N_5936);
nor U11530 (N_11530,N_9982,N_5909);
nor U11531 (N_11531,N_7784,N_9479);
and U11532 (N_11532,N_7033,N_8413);
nor U11533 (N_11533,N_9246,N_6629);
nand U11534 (N_11534,N_9390,N_5692);
nand U11535 (N_11535,N_9290,N_6884);
nand U11536 (N_11536,N_6550,N_7003);
xnor U11537 (N_11537,N_8510,N_9312);
nand U11538 (N_11538,N_6544,N_5053);
or U11539 (N_11539,N_6287,N_9725);
nand U11540 (N_11540,N_9411,N_5469);
and U11541 (N_11541,N_9200,N_8823);
nor U11542 (N_11542,N_6926,N_7767);
xor U11543 (N_11543,N_9785,N_9158);
or U11544 (N_11544,N_9914,N_5300);
and U11545 (N_11545,N_8320,N_7527);
and U11546 (N_11546,N_7674,N_7161);
or U11547 (N_11547,N_9347,N_7239);
nor U11548 (N_11548,N_9340,N_5441);
nor U11549 (N_11549,N_9185,N_8439);
xor U11550 (N_11550,N_8553,N_8665);
nor U11551 (N_11551,N_7414,N_7198);
nor U11552 (N_11552,N_5430,N_5249);
xnor U11553 (N_11553,N_8980,N_9308);
or U11554 (N_11554,N_5344,N_7884);
xor U11555 (N_11555,N_9834,N_6437);
or U11556 (N_11556,N_5207,N_5424);
nand U11557 (N_11557,N_9574,N_8282);
and U11558 (N_11558,N_6523,N_9088);
nor U11559 (N_11559,N_9453,N_6196);
and U11560 (N_11560,N_9645,N_6096);
or U11561 (N_11561,N_6468,N_9165);
or U11562 (N_11562,N_9513,N_9947);
nor U11563 (N_11563,N_8619,N_9573);
nor U11564 (N_11564,N_5519,N_8850);
nor U11565 (N_11565,N_9183,N_9201);
nor U11566 (N_11566,N_7895,N_5443);
xor U11567 (N_11567,N_9985,N_5717);
nand U11568 (N_11568,N_9638,N_6087);
or U11569 (N_11569,N_9373,N_8340);
or U11570 (N_11570,N_8091,N_9299);
and U11571 (N_11571,N_6890,N_5281);
nor U11572 (N_11572,N_6222,N_6892);
nor U11573 (N_11573,N_6758,N_6440);
xnor U11574 (N_11574,N_9757,N_5020);
nor U11575 (N_11575,N_9330,N_9691);
and U11576 (N_11576,N_5470,N_8860);
or U11577 (N_11577,N_9636,N_7232);
nand U11578 (N_11578,N_5129,N_7757);
nand U11579 (N_11579,N_8015,N_8642);
and U11580 (N_11580,N_6762,N_7200);
nand U11581 (N_11581,N_6682,N_7512);
nand U11582 (N_11582,N_7089,N_5257);
or U11583 (N_11583,N_8890,N_6509);
and U11584 (N_11584,N_8630,N_9654);
and U11585 (N_11585,N_8126,N_7057);
or U11586 (N_11586,N_8631,N_7201);
nor U11587 (N_11587,N_8099,N_9478);
nor U11588 (N_11588,N_5196,N_9536);
or U11589 (N_11589,N_7031,N_8996);
or U11590 (N_11590,N_5603,N_8866);
nor U11591 (N_11591,N_9650,N_8913);
nor U11592 (N_11592,N_7651,N_5146);
nor U11593 (N_11593,N_8919,N_6914);
or U11594 (N_11594,N_5052,N_8444);
xor U11595 (N_11595,N_8069,N_5704);
nand U11596 (N_11596,N_6279,N_6779);
or U11597 (N_11597,N_6392,N_5279);
nand U11598 (N_11598,N_9907,N_5159);
nor U11599 (N_11599,N_8310,N_6201);
and U11600 (N_11600,N_7848,N_8205);
nand U11601 (N_11601,N_5786,N_5336);
or U11602 (N_11602,N_8192,N_8360);
nand U11603 (N_11603,N_8514,N_5972);
nand U11604 (N_11604,N_6658,N_8244);
or U11605 (N_11605,N_6249,N_6401);
nor U11606 (N_11606,N_8227,N_5320);
nor U11607 (N_11607,N_8513,N_8906);
or U11608 (N_11608,N_6556,N_6082);
nor U11609 (N_11609,N_5729,N_9355);
nor U11610 (N_11610,N_8132,N_7370);
nand U11611 (N_11611,N_7835,N_7589);
nor U11612 (N_11612,N_9303,N_6410);
and U11613 (N_11613,N_7493,N_9861);
and U11614 (N_11614,N_8754,N_6904);
and U11615 (N_11615,N_9674,N_7471);
xnor U11616 (N_11616,N_5858,N_8104);
nand U11617 (N_11617,N_5832,N_5673);
nand U11618 (N_11618,N_8605,N_6843);
and U11619 (N_11619,N_7297,N_5245);
nor U11620 (N_11620,N_8136,N_6640);
and U11621 (N_11621,N_5324,N_7747);
nor U11622 (N_11622,N_5394,N_8294);
nor U11623 (N_11623,N_6698,N_8336);
nor U11624 (N_11624,N_7873,N_5571);
nand U11625 (N_11625,N_9279,N_9663);
nand U11626 (N_11626,N_6491,N_8234);
nor U11627 (N_11627,N_6724,N_7729);
nand U11628 (N_11628,N_9117,N_7585);
and U11629 (N_11629,N_6389,N_6290);
or U11630 (N_11630,N_7409,N_5334);
and U11631 (N_11631,N_8527,N_7207);
or U11632 (N_11632,N_9784,N_6112);
nand U11633 (N_11633,N_6369,N_6853);
nand U11634 (N_11634,N_7681,N_8985);
or U11635 (N_11635,N_9239,N_5922);
and U11636 (N_11636,N_9525,N_5306);
nand U11637 (N_11637,N_8435,N_9147);
xnor U11638 (N_11638,N_5128,N_8961);
nor U11639 (N_11639,N_9728,N_7486);
and U11640 (N_11640,N_9657,N_7839);
or U11641 (N_11641,N_6866,N_9392);
and U11642 (N_11642,N_5429,N_7759);
nand U11643 (N_11643,N_9686,N_7068);
nor U11644 (N_11644,N_8917,N_6067);
and U11645 (N_11645,N_5186,N_5517);
and U11646 (N_11646,N_8432,N_5690);
and U11647 (N_11647,N_5701,N_8416);
xor U11648 (N_11648,N_8570,N_7121);
and U11649 (N_11649,N_7090,N_8078);
nand U11650 (N_11650,N_9710,N_9463);
nor U11651 (N_11651,N_6869,N_6705);
nand U11652 (N_11652,N_6275,N_6607);
nand U11653 (N_11653,N_7568,N_9264);
nor U11654 (N_11654,N_6066,N_8546);
or U11655 (N_11655,N_7282,N_9817);
xor U11656 (N_11656,N_5934,N_8339);
and U11657 (N_11657,N_5458,N_8304);
nand U11658 (N_11658,N_5059,N_6334);
or U11659 (N_11659,N_7088,N_9265);
nor U11660 (N_11660,N_7742,N_9206);
and U11661 (N_11661,N_8034,N_6837);
nand U11662 (N_11662,N_9301,N_5485);
xnor U11663 (N_11663,N_9412,N_9166);
and U11664 (N_11664,N_7268,N_7071);
and U11665 (N_11665,N_5088,N_8176);
and U11666 (N_11666,N_7343,N_7430);
and U11667 (N_11667,N_9987,N_7831);
nor U11668 (N_11668,N_6598,N_9718);
xnor U11669 (N_11669,N_7845,N_8799);
nor U11670 (N_11670,N_6796,N_9444);
and U11671 (N_11671,N_8699,N_9878);
and U11672 (N_11672,N_7150,N_7790);
and U11673 (N_11673,N_6054,N_6119);
or U11674 (N_11674,N_8285,N_7897);
xnor U11675 (N_11675,N_9420,N_5241);
or U11676 (N_11676,N_9269,N_8380);
nand U11677 (N_11677,N_8689,N_8950);
or U11678 (N_11678,N_9226,N_6962);
or U11679 (N_11679,N_5639,N_8316);
or U11680 (N_11680,N_8155,N_8366);
nand U11681 (N_11681,N_7447,N_7504);
and U11682 (N_11682,N_7007,N_9934);
and U11683 (N_11683,N_5564,N_5594);
nor U11684 (N_11684,N_8715,N_7272);
or U11685 (N_11685,N_8178,N_9923);
nor U11686 (N_11686,N_7498,N_9516);
nand U11687 (N_11687,N_9940,N_6198);
or U11688 (N_11688,N_5373,N_5625);
nand U11689 (N_11689,N_5005,N_5388);
and U11690 (N_11690,N_6464,N_6325);
nor U11691 (N_11691,N_6699,N_9561);
and U11692 (N_11692,N_9953,N_9283);
xor U11693 (N_11693,N_8870,N_5465);
nand U11694 (N_11694,N_8166,N_9864);
and U11695 (N_11695,N_5298,N_6273);
and U11696 (N_11696,N_9868,N_8710);
or U11697 (N_11697,N_5940,N_6560);
and U11698 (N_11698,N_5287,N_9792);
nor U11699 (N_11699,N_6046,N_9181);
nand U11700 (N_11700,N_5171,N_7965);
nand U11701 (N_11701,N_8574,N_5763);
and U11702 (N_11702,N_7285,N_9787);
or U11703 (N_11703,N_8612,N_9723);
and U11704 (N_11704,N_5274,N_6839);
xor U11705 (N_11705,N_5439,N_8334);
or U11706 (N_11706,N_5104,N_9337);
and U11707 (N_11707,N_9099,N_5866);
xnor U11708 (N_11708,N_6668,N_8533);
or U11709 (N_11709,N_7964,N_9605);
and U11710 (N_11710,N_5978,N_7525);
or U11711 (N_11711,N_8542,N_7291);
or U11712 (N_11712,N_6343,N_8338);
and U11713 (N_11713,N_6190,N_8354);
nor U11714 (N_11714,N_5156,N_5677);
nand U11715 (N_11715,N_6522,N_6173);
nor U11716 (N_11716,N_7408,N_8840);
nor U11717 (N_11717,N_8204,N_6317);
nand U11718 (N_11718,N_6542,N_6147);
nand U11719 (N_11719,N_8309,N_6632);
and U11720 (N_11720,N_8598,N_6399);
and U11721 (N_11721,N_8929,N_5488);
or U11722 (N_11722,N_6442,N_8704);
nand U11723 (N_11723,N_5873,N_8006);
nor U11724 (N_11724,N_8406,N_5753);
and U11725 (N_11725,N_5945,N_6546);
nand U11726 (N_11726,N_7911,N_8250);
or U11727 (N_11727,N_5890,N_9250);
xnor U11728 (N_11728,N_6395,N_8111);
and U11729 (N_11729,N_8394,N_6072);
nand U11730 (N_11730,N_8389,N_7710);
and U11731 (N_11731,N_5837,N_5036);
nor U11732 (N_11732,N_5212,N_6217);
xor U11733 (N_11733,N_5363,N_7373);
nor U11734 (N_11734,N_5935,N_6484);
nor U11735 (N_11735,N_8088,N_6107);
xor U11736 (N_11736,N_7180,N_6662);
xor U11737 (N_11737,N_6188,N_9631);
xnor U11738 (N_11738,N_8712,N_7629);
or U11739 (N_11739,N_9294,N_7875);
nor U11740 (N_11740,N_9106,N_9085);
or U11741 (N_11741,N_7188,N_9911);
nor U11742 (N_11742,N_5413,N_7616);
nor U11743 (N_11743,N_7532,N_6045);
nor U11744 (N_11744,N_9764,N_7973);
xnor U11745 (N_11745,N_8213,N_6206);
nand U11746 (N_11746,N_5877,N_9667);
nor U11747 (N_11747,N_9199,N_5899);
nor U11748 (N_11748,N_7264,N_5626);
or U11749 (N_11749,N_8164,N_5884);
nor U11750 (N_11750,N_7142,N_7441);
and U11751 (N_11751,N_5016,N_8939);
or U11752 (N_11752,N_9961,N_9462);
nor U11753 (N_11753,N_8186,N_6347);
xnor U11754 (N_11754,N_9712,N_6090);
and U11755 (N_11755,N_5166,N_7661);
or U11756 (N_11756,N_9168,N_5856);
or U11757 (N_11757,N_7283,N_7882);
or U11758 (N_11758,N_5302,N_5096);
nand U11759 (N_11759,N_5793,N_7445);
or U11760 (N_11760,N_6394,N_8187);
nand U11761 (N_11761,N_8174,N_5588);
and U11762 (N_11762,N_5548,N_8942);
nor U11763 (N_11763,N_7823,N_8027);
nor U11764 (N_11764,N_7500,N_7025);
and U11765 (N_11765,N_7536,N_8691);
nor U11766 (N_11766,N_6432,N_7659);
nand U11767 (N_11767,N_9477,N_7998);
xnor U11768 (N_11768,N_8596,N_7191);
xor U11769 (N_11769,N_5182,N_8740);
nand U11770 (N_11770,N_8777,N_6697);
nor U11771 (N_11771,N_6645,N_9086);
or U11772 (N_11772,N_8875,N_6335);
xor U11773 (N_11773,N_8146,N_8669);
xnor U11774 (N_11774,N_6932,N_7360);
or U11775 (N_11775,N_6272,N_9323);
nor U11776 (N_11776,N_7715,N_5453);
nor U11777 (N_11777,N_8831,N_8232);
nand U11778 (N_11778,N_7170,N_9289);
and U11779 (N_11779,N_9808,N_6250);
nand U11780 (N_11780,N_7428,N_9594);
or U11781 (N_11781,N_5696,N_9219);
nor U11782 (N_11782,N_7076,N_9893);
or U11783 (N_11783,N_8075,N_7563);
nor U11784 (N_11784,N_9679,N_7714);
nor U11785 (N_11785,N_8408,N_9853);
xor U11786 (N_11786,N_6356,N_7981);
nor U11787 (N_11787,N_9669,N_5713);
or U11788 (N_11788,N_7129,N_7494);
nand U11789 (N_11789,N_8423,N_5913);
nand U11790 (N_11790,N_8714,N_6073);
or U11791 (N_11791,N_8215,N_8773);
and U11792 (N_11792,N_8762,N_5683);
nand U11793 (N_11793,N_5950,N_6920);
nand U11794 (N_11794,N_9078,N_8278);
xor U11795 (N_11795,N_9313,N_5414);
nand U11796 (N_11796,N_9363,N_9434);
nor U11797 (N_11797,N_5695,N_6672);
nand U11798 (N_11798,N_8838,N_9336);
nand U11799 (N_11799,N_8210,N_8490);
xor U11800 (N_11800,N_6194,N_6950);
and U11801 (N_11801,N_5915,N_8256);
nor U11802 (N_11802,N_6863,N_7355);
and U11803 (N_11803,N_7081,N_6576);
and U11804 (N_11804,N_8856,N_8507);
or U11805 (N_11805,N_5051,N_8842);
or U11806 (N_11806,N_6685,N_9151);
or U11807 (N_11807,N_8436,N_8085);
and U11808 (N_11808,N_9519,N_5942);
or U11809 (N_11809,N_6732,N_8652);
and U11810 (N_11810,N_9924,N_7166);
xor U11811 (N_11811,N_9481,N_6847);
nand U11812 (N_11812,N_6751,N_5907);
nand U11813 (N_11813,N_5401,N_5620);
or U11814 (N_11814,N_9500,N_5726);
nor U11815 (N_11815,N_7837,N_5600);
nand U11816 (N_11816,N_8262,N_6827);
or U11817 (N_11817,N_8964,N_5118);
nor U11818 (N_11818,N_7240,N_7720);
nor U11819 (N_11819,N_5818,N_9047);
nor U11820 (N_11820,N_8815,N_9703);
nor U11821 (N_11821,N_5776,N_7022);
and U11822 (N_11822,N_7234,N_7700);
or U11823 (N_11823,N_7830,N_8020);
nand U11824 (N_11824,N_5289,N_5495);
and U11825 (N_11825,N_8148,N_8563);
nor U11826 (N_11826,N_6270,N_6567);
and U11827 (N_11827,N_5079,N_9902);
or U11828 (N_11828,N_8971,N_7892);
and U11829 (N_11829,N_9694,N_6800);
and U11830 (N_11830,N_5770,N_6836);
nor U11831 (N_11831,N_7768,N_8026);
nand U11832 (N_11832,N_6928,N_9840);
and U11833 (N_11833,N_8956,N_8218);
or U11834 (N_11834,N_6144,N_9210);
nand U11835 (N_11835,N_6094,N_6348);
nand U11836 (N_11836,N_9435,N_5669);
and U11837 (N_11837,N_9243,N_8934);
nor U11838 (N_11838,N_6527,N_5590);
or U11839 (N_11839,N_7122,N_7311);
nor U11840 (N_11840,N_5616,N_8687);
or U11841 (N_11841,N_8225,N_8156);
nor U11842 (N_11842,N_7991,N_5756);
or U11843 (N_11843,N_9096,N_7987);
nor U11844 (N_11844,N_8750,N_8200);
nor U11845 (N_11845,N_9458,N_8927);
or U11846 (N_11846,N_7467,N_7832);
and U11847 (N_11847,N_7047,N_8499);
and U11848 (N_11848,N_7871,N_7435);
nand U11849 (N_11849,N_7298,N_7510);
nor U11850 (N_11850,N_8382,N_7160);
or U11851 (N_11851,N_9859,N_7165);
nor U11852 (N_11852,N_7776,N_9847);
and U11853 (N_11853,N_9093,N_8417);
nand U11854 (N_11854,N_6586,N_9935);
and U11855 (N_11855,N_5791,N_5293);
nand U11856 (N_11856,N_9867,N_7267);
xnor U11857 (N_11857,N_9282,N_5720);
or U11858 (N_11858,N_5523,N_9459);
xnor U11859 (N_11859,N_5305,N_9721);
nor U11860 (N_11860,N_5502,N_6673);
nor U11861 (N_11861,N_8576,N_9379);
and U11862 (N_11862,N_6445,N_6128);
xor U11863 (N_11863,N_9586,N_6391);
or U11864 (N_11864,N_9800,N_9160);
nand U11865 (N_11865,N_6618,N_9083);
and U11866 (N_11866,N_8658,N_5707);
nand U11867 (N_11867,N_7258,N_8117);
xor U11868 (N_11868,N_5368,N_6681);
nand U11869 (N_11869,N_6115,N_5066);
nand U11870 (N_11870,N_6516,N_8059);
and U11871 (N_11871,N_7499,N_9148);
nand U11872 (N_11872,N_6261,N_7179);
nand U11873 (N_11873,N_6754,N_7321);
and U11874 (N_11874,N_7505,N_5694);
nor U11875 (N_11875,N_8851,N_7193);
or U11876 (N_11876,N_7853,N_8995);
nor U11877 (N_11877,N_7815,N_9995);
nand U11878 (N_11878,N_5944,N_6130);
nand U11879 (N_11879,N_7399,N_7341);
or U11880 (N_11880,N_7045,N_7936);
xor U11881 (N_11881,N_8260,N_7104);
or U11882 (N_11882,N_6968,N_7970);
nand U11883 (N_11883,N_7356,N_9475);
nand U11884 (N_11884,N_9706,N_9314);
nor U11885 (N_11885,N_6529,N_6765);
nor U11886 (N_11886,N_8584,N_9549);
or U11887 (N_11887,N_9983,N_8199);
nor U11888 (N_11888,N_8946,N_9943);
or U11889 (N_11889,N_9795,N_5609);
or U11890 (N_11890,N_8663,N_6935);
and U11891 (N_11891,N_8201,N_9735);
nand U11892 (N_11892,N_5242,N_5327);
nor U11893 (N_11893,N_8348,N_7976);
or U11894 (N_11894,N_6949,N_6320);
or U11895 (N_11895,N_7588,N_5645);
nor U11896 (N_11896,N_9138,N_5567);
nand U11897 (N_11897,N_8737,N_7978);
nand U11898 (N_11898,N_8212,N_9618);
nand U11899 (N_11899,N_9228,N_5906);
and U11900 (N_11900,N_5201,N_8948);
or U11901 (N_11901,N_6792,N_6906);
and U11902 (N_11902,N_8816,N_8905);
xnor U11903 (N_11903,N_8864,N_6976);
nand U11904 (N_11904,N_8577,N_9715);
or U11905 (N_11905,N_6813,N_5340);
or U11906 (N_11906,N_5604,N_9622);
nor U11907 (N_11907,N_6597,N_7618);
or U11908 (N_11908,N_8157,N_8873);
or U11909 (N_11909,N_6545,N_9873);
nor U11910 (N_11910,N_5744,N_9080);
nor U11911 (N_11911,N_8532,N_8450);
nand U11912 (N_11912,N_7004,N_5412);
or U11913 (N_11913,N_6235,N_7574);
nand U11914 (N_11914,N_5190,N_8318);
and U11915 (N_11915,N_6480,N_7668);
nand U11916 (N_11916,N_7097,N_5743);
nand U11917 (N_11917,N_9687,N_6274);
nor U11918 (N_11918,N_8632,N_8251);
nor U11919 (N_11919,N_5260,N_6341);
or U11920 (N_11920,N_7624,N_5918);
nand U11921 (N_11921,N_5497,N_9562);
nand U11922 (N_11922,N_6477,N_8967);
or U11923 (N_11923,N_9153,N_7296);
nor U11924 (N_11924,N_8112,N_7495);
nand U11925 (N_11925,N_6457,N_8030);
or U11926 (N_11926,N_7899,N_6286);
and U11927 (N_11927,N_7294,N_7281);
nor U11928 (N_11928,N_7219,N_7770);
or U11929 (N_11929,N_6626,N_9540);
nor U11930 (N_11930,N_9813,N_6388);
nor U11931 (N_11931,N_7173,N_9342);
nand U11932 (N_11932,N_7413,N_6865);
and U11933 (N_11933,N_6136,N_9688);
and U11934 (N_11934,N_8561,N_5209);
nand U11935 (N_11935,N_7320,N_7963);
and U11936 (N_11936,N_8505,N_7407);
or U11937 (N_11937,N_8936,N_7330);
xor U11938 (N_11938,N_8830,N_8772);
xor U11939 (N_11939,N_9829,N_7929);
nor U11940 (N_11940,N_6982,N_5153);
or U11941 (N_11941,N_8843,N_7039);
or U11942 (N_11942,N_5990,N_6532);
and U11943 (N_11943,N_7736,N_5926);
or U11944 (N_11944,N_5533,N_9734);
nand U11945 (N_11945,N_5703,N_6312);
and U11946 (N_11946,N_6003,N_8161);
or U11947 (N_11947,N_8445,N_6574);
xnor U11948 (N_11948,N_9214,N_5139);
nand U11949 (N_11949,N_5614,N_6716);
nand U11950 (N_11950,N_7937,N_9027);
xor U11951 (N_11951,N_5343,N_6451);
and U11952 (N_11952,N_8319,N_7783);
or U11953 (N_11953,N_9063,N_9644);
xor U11954 (N_11954,N_7842,N_8182);
or U11955 (N_11955,N_7760,N_9729);
and U11956 (N_11956,N_7044,N_8907);
xnor U11957 (N_11957,N_6213,N_6064);
and U11958 (N_11958,N_7890,N_6620);
and U11959 (N_11959,N_9207,N_7708);
and U11960 (N_11960,N_5246,N_8016);
and U11961 (N_11961,N_5232,N_6603);
nor U11962 (N_11962,N_7781,N_9542);
nand U11963 (N_11963,N_7038,N_9267);
nand U11964 (N_11964,N_6841,N_9326);
nor U11965 (N_11965,N_8835,N_9850);
xor U11966 (N_11966,N_6674,N_5893);
nand U11967 (N_11967,N_8383,N_7450);
or U11968 (N_11968,N_5472,N_9593);
nand U11969 (N_11969,N_7344,N_8565);
and U11970 (N_11970,N_5261,N_5452);
and U11971 (N_11971,N_8828,N_9380);
and U11972 (N_11972,N_9603,N_7713);
xor U11973 (N_11973,N_7530,N_7968);
or U11974 (N_11974,N_9530,N_5372);
and U11975 (N_11975,N_8556,N_7124);
nand U11976 (N_11976,N_7230,N_5463);
nand U11977 (N_11977,N_9281,N_6226);
nand U11978 (N_11978,N_8424,N_8595);
nand U11979 (N_11979,N_8167,N_6946);
or U11980 (N_11980,N_8805,N_6984);
and U11981 (N_11981,N_6953,N_7431);
xor U11982 (N_11982,N_6292,N_8538);
nor U11983 (N_11983,N_8140,N_6988);
or U11984 (N_11984,N_6581,N_9968);
and U11985 (N_11985,N_7073,N_9797);
nor U11986 (N_11986,N_6924,N_8793);
and U11987 (N_11987,N_9296,N_9926);
nand U11988 (N_11988,N_7397,N_5203);
nor U11989 (N_11989,N_9580,N_8147);
nand U11990 (N_11990,N_9831,N_6430);
nor U11991 (N_11991,N_9749,N_7997);
or U11992 (N_11992,N_9309,N_6049);
nor U11993 (N_11993,N_8040,N_6893);
nor U11994 (N_11994,N_6256,N_5034);
nor U11995 (N_11995,N_7733,N_5167);
or U11996 (N_11996,N_5496,N_5882);
or U11997 (N_11997,N_7820,N_5498);
nand U11998 (N_11998,N_8365,N_5892);
nand U11999 (N_11999,N_6110,N_7507);
or U12000 (N_12000,N_9193,N_6677);
xnor U12001 (N_12001,N_6888,N_8626);
nand U12002 (N_12002,N_6802,N_9145);
nor U12003 (N_12003,N_5712,N_9862);
nor U12004 (N_12004,N_5961,N_9585);
nand U12005 (N_12005,N_8061,N_6832);
or U12006 (N_12006,N_5179,N_6728);
and U12007 (N_12007,N_6660,N_9790);
and U12008 (N_12008,N_9190,N_8960);
nor U12009 (N_12009,N_9584,N_6425);
or U12010 (N_12010,N_6776,N_7876);
nand U12011 (N_12011,N_9361,N_6580);
and U12012 (N_12012,N_5173,N_7766);
xnor U12013 (N_12013,N_9109,N_8137);
or U12014 (N_12014,N_7108,N_5434);
or U12015 (N_12015,N_8395,N_6588);
or U12016 (N_12016,N_9273,N_6331);
and U12017 (N_12017,N_6578,N_8717);
and U12018 (N_12018,N_8415,N_6165);
nor U12019 (N_12019,N_5122,N_6942);
and U12020 (N_12020,N_6321,N_5632);
or U12021 (N_12021,N_8763,N_7652);
nand U12022 (N_12022,N_7335,N_8743);
xnor U12023 (N_12023,N_8045,N_7473);
or U12024 (N_12024,N_8529,N_9578);
or U12025 (N_12025,N_8865,N_9300);
or U12026 (N_12026,N_5172,N_7868);
xor U12027 (N_12027,N_8120,N_7334);
and U12028 (N_12028,N_8786,N_9020);
or U12029 (N_12029,N_7887,N_7103);
nand U12030 (N_12030,N_7306,N_6040);
nor U12031 (N_12031,N_6876,N_7056);
nand U12032 (N_12032,N_7919,N_7614);
and U12033 (N_12033,N_9389,N_8240);
nor U12034 (N_12034,N_6555,N_6693);
nand U12035 (N_12035,N_9242,N_6760);
nor U12036 (N_12036,N_8369,N_5715);
nand U12037 (N_12037,N_6456,N_8822);
nand U12038 (N_12038,N_9616,N_7980);
and U12039 (N_12039,N_7558,N_9699);
and U12040 (N_12040,N_9552,N_8564);
nand U12041 (N_12041,N_6055,N_5035);
and U12042 (N_12042,N_5332,N_9157);
nand U12043 (N_12043,N_9350,N_5722);
nor U12044 (N_12044,N_9394,N_7130);
and U12045 (N_12045,N_9090,N_9403);
nor U12046 (N_12046,N_6140,N_7395);
nor U12047 (N_12047,N_7521,N_9231);
nor U12048 (N_12048,N_7316,N_6825);
xnor U12049 (N_12049,N_8301,N_6354);
nand U12050 (N_12050,N_6223,N_5838);
and U12051 (N_12051,N_9492,N_5886);
or U12052 (N_12052,N_6937,N_6908);
or U12053 (N_12053,N_5755,N_8916);
and U12054 (N_12054,N_8594,N_7115);
xor U12055 (N_12055,N_6694,N_7735);
nand U12056 (N_12056,N_6479,N_7881);
or U12057 (N_12057,N_5534,N_6568);
xnor U12058 (N_12058,N_7432,N_7609);
nand U12059 (N_12059,N_5077,N_5448);
nand U12060 (N_12060,N_9845,N_8028);
nand U12061 (N_12061,N_8795,N_7082);
nand U12062 (N_12062,N_6106,N_5442);
nor U12063 (N_12063,N_8970,N_5551);
nand U12064 (N_12064,N_9899,N_6885);
or U12065 (N_12065,N_7065,N_9977);
nor U12066 (N_12066,N_9922,N_7210);
or U12067 (N_12067,N_7307,N_6707);
nor U12068 (N_12068,N_7133,N_9409);
nor U12069 (N_12069,N_5390,N_8306);
or U12070 (N_12070,N_9830,N_6789);
and U12071 (N_12071,N_5000,N_7384);
nand U12072 (N_12072,N_7362,N_7310);
nand U12073 (N_12073,N_7017,N_7385);
or U12074 (N_12074,N_7994,N_6125);
or U12075 (N_12075,N_9404,N_7744);
nand U12076 (N_12076,N_7437,N_9810);
or U12077 (N_12077,N_9741,N_8662);
or U12078 (N_12078,N_5185,N_9992);
xor U12079 (N_12079,N_7724,N_6963);
and U12080 (N_12080,N_5526,N_5263);
and U12081 (N_12081,N_9159,N_8067);
xor U12082 (N_12082,N_5366,N_8222);
and U12083 (N_12083,N_5004,N_9164);
or U12084 (N_12084,N_7456,N_7864);
or U12085 (N_12085,N_6916,N_9848);
or U12086 (N_12086,N_5924,N_7637);
or U12087 (N_12087,N_6099,N_7593);
and U12088 (N_12088,N_5923,N_6557);
nand U12089 (N_12089,N_6729,N_5643);
nor U12090 (N_12090,N_8101,N_8437);
nand U12091 (N_12091,N_8846,N_5162);
or U12092 (N_12092,N_5767,N_7064);
nand U12093 (N_12093,N_8589,N_8983);
and U12094 (N_12094,N_7833,N_6780);
nand U12095 (N_12095,N_8965,N_5875);
and U12096 (N_12096,N_9806,N_7118);
nand U12097 (N_12097,N_9856,N_9949);
xnor U12098 (N_12098,N_9662,N_9886);
nor U12099 (N_12099,N_7553,N_7653);
xor U12100 (N_12100,N_5525,N_7292);
nand U12101 (N_12101,N_5105,N_8473);
xnor U12102 (N_12102,N_8265,N_5894);
nand U12103 (N_12103,N_6777,N_6889);
or U12104 (N_12104,N_6563,N_6636);
nor U12105 (N_12105,N_7591,N_6009);
nand U12106 (N_12106,N_7163,N_9608);
nor U12107 (N_12107,N_9766,N_5176);
or U12108 (N_12108,N_8705,N_7028);
and U12109 (N_12109,N_5532,N_9167);
or U12110 (N_12110,N_9826,N_8650);
nand U12111 (N_12111,N_7540,N_6365);
nand U12112 (N_12112,N_7418,N_9410);
or U12113 (N_12113,N_7636,N_9559);
nor U12114 (N_12114,N_6234,N_7814);
xor U12115 (N_12115,N_9018,N_7502);
nor U12116 (N_12116,N_8912,N_7172);
and U12117 (N_12117,N_7939,N_9268);
or U12118 (N_12118,N_9486,N_5435);
nor U12119 (N_12119,N_8855,N_5730);
or U12120 (N_12120,N_6604,N_9612);
nor U12121 (N_12121,N_6886,N_9128);
nand U12122 (N_12122,N_6631,N_9431);
nor U12123 (N_12123,N_5352,N_8332);
or U12124 (N_12124,N_6809,N_5932);
nand U12125 (N_12125,N_6536,N_7638);
or U12126 (N_12126,N_6611,N_9030);
nand U12127 (N_12127,N_6844,N_9135);
or U12128 (N_12128,N_7737,N_5389);
or U12129 (N_12129,N_7804,N_9634);
nor U12130 (N_12130,N_9877,N_5421);
nor U12131 (N_12131,N_8259,N_5810);
and U12132 (N_12132,N_5904,N_8074);
or U12133 (N_12133,N_6727,N_9768);
or U12134 (N_12134,N_7190,N_9780);
and U12135 (N_12135,N_8924,N_8462);
xor U12136 (N_12136,N_5474,N_9049);
and U12137 (N_12137,N_9887,N_5116);
nand U12138 (N_12138,N_6207,N_7323);
and U12139 (N_12139,N_9941,N_6406);
xnor U12140 (N_12140,N_5674,N_5310);
xnor U12141 (N_12141,N_6539,N_9894);
and U12142 (N_12142,N_6026,N_5391);
nor U12143 (N_12143,N_5216,N_7054);
and U12144 (N_12144,N_7944,N_5779);
nand U12145 (N_12145,N_9259,N_9224);
and U12146 (N_12146,N_8749,N_9752);
nor U12147 (N_12147,N_5062,N_6559);
or U12148 (N_12148,N_6431,N_8385);
nor U12149 (N_12149,N_6510,N_6251);
nor U12150 (N_12150,N_9866,N_9002);
and U12151 (N_12151,N_5970,N_8504);
and U12152 (N_12152,N_6995,N_5124);
or U12153 (N_12153,N_9816,N_8721);
nor U12154 (N_12154,N_6838,N_5648);
and U12155 (N_12155,N_5824,N_9789);
nand U12156 (N_12156,N_7789,N_8108);
and U12157 (N_12157,N_8833,N_8300);
or U12158 (N_12158,N_9804,N_5328);
nor U12159 (N_12159,N_6042,N_5933);
nand U12160 (N_12160,N_5338,N_5271);
nor U12161 (N_12161,N_7448,N_9364);
and U12162 (N_12162,N_9024,N_9288);
nand U12163 (N_12163,N_8388,N_9111);
xnor U12164 (N_12164,N_7727,N_7101);
nand U12165 (N_12165,N_6502,N_9152);
and U12166 (N_12166,N_9889,N_5938);
nand U12167 (N_12167,N_5581,N_7550);
nor U12168 (N_12168,N_9624,N_6081);
nor U12169 (N_12169,N_9579,N_6623);
nand U12170 (N_12170,N_8001,N_9422);
xnor U12171 (N_12171,N_5432,N_7252);
and U12172 (N_12172,N_9315,N_6718);
nor U12173 (N_12173,N_6691,N_9639);
nor U12174 (N_12174,N_9607,N_7001);
or U12175 (N_12175,N_9050,N_6562);
nand U12176 (N_12176,N_5980,N_8730);
and U12177 (N_12177,N_7535,N_8945);
nor U12178 (N_12178,N_8701,N_9387);
nand U12179 (N_12179,N_9629,N_7731);
or U12180 (N_12180,N_5491,N_6856);
and U12181 (N_12181,N_7841,N_8523);
nand U12182 (N_12182,N_6549,N_7975);
nand U12183 (N_12183,N_5070,N_9760);
or U12184 (N_12184,N_8467,N_7554);
nor U12185 (N_12185,N_6665,N_5805);
nor U12186 (N_12186,N_5803,N_7380);
or U12187 (N_12187,N_8397,N_8801);
xor U12188 (N_12188,N_5351,N_6093);
and U12189 (N_12189,N_7461,N_9989);
and U12190 (N_12190,N_6720,N_9614);
or U12191 (N_12191,N_9823,N_7607);
or U12192 (N_12192,N_7667,N_6571);
nor U12193 (N_12193,N_8776,N_6500);
nor U12194 (N_12194,N_5493,N_5655);
or U12195 (N_12195,N_7114,N_8012);
nand U12196 (N_12196,N_9140,N_7680);
or U12197 (N_12197,N_9904,N_8280);
or U12198 (N_12198,N_8767,N_5231);
or U12199 (N_12199,N_6088,N_5699);
nor U12200 (N_12200,N_7416,N_6721);
and U12201 (N_12201,N_9742,N_8131);
or U12202 (N_12202,N_6894,N_8261);
nand U12203 (N_12203,N_5247,N_9252);
nor U12204 (N_12204,N_5964,N_7796);
nand U12205 (N_12205,N_5163,N_9073);
and U12206 (N_12206,N_5709,N_6218);
nand U12207 (N_12207,N_7314,N_7662);
nor U12208 (N_12208,N_7723,N_8568);
nand U12209 (N_12209,N_8602,N_7794);
nor U12210 (N_12210,N_6485,N_8414);
or U12211 (N_12211,N_8973,N_5267);
or U12212 (N_12212,N_7573,N_7933);
or U12213 (N_12213,N_8520,N_7974);
and U12214 (N_12214,N_8271,N_7458);
or U12215 (N_12215,N_9113,N_7528);
or U12216 (N_12216,N_6121,N_8614);
or U12217 (N_12217,N_7633,N_9188);
and U12218 (N_12218,N_5668,N_8217);
nor U12219 (N_12219,N_8247,N_9529);
xor U12220 (N_12220,N_7069,N_5840);
or U12221 (N_12221,N_7394,N_5080);
and U12222 (N_12222,N_8810,N_6360);
and U12223 (N_12223,N_7023,N_6380);
nor U12224 (N_12224,N_5384,N_8179);
nor U12225 (N_12225,N_7632,N_6820);
and U12226 (N_12226,N_5741,N_7584);
xnor U12227 (N_12227,N_9990,N_7707);
and U12228 (N_12228,N_7438,N_6439);
nor U12229 (N_12229,N_8237,N_5897);
nor U12230 (N_12230,N_5353,N_5081);
nand U12231 (N_12231,N_7898,N_7391);
and U12232 (N_12232,N_6269,N_7758);
or U12233 (N_12233,N_7086,N_9678);
and U12234 (N_12234,N_5962,N_9659);
nand U12235 (N_12235,N_7182,N_9860);
and U12236 (N_12236,N_6534,N_9896);
nand U12237 (N_12237,N_9918,N_7932);
xnor U12238 (N_12238,N_9357,N_7302);
and U12239 (N_12239,N_5330,N_7619);
xor U12240 (N_12240,N_5733,N_8441);
and U12241 (N_12241,N_6879,N_7717);
nand U12242 (N_12242,N_7478,N_8048);
and U12243 (N_12243,N_5376,N_6407);
and U12244 (N_12244,N_9240,N_9170);
nor U12245 (N_12245,N_5911,N_6383);
nand U12246 (N_12246,N_6158,N_7665);
or U12247 (N_12247,N_9130,N_7989);
nor U12248 (N_12248,N_9876,N_9875);
and U12249 (N_12249,N_9583,N_5949);
nand U12250 (N_12250,N_7803,N_5960);
xnor U12251 (N_12251,N_8536,N_9197);
nand U12252 (N_12252,N_8925,N_5969);
and U12253 (N_12253,N_8168,N_6078);
or U12254 (N_12254,N_5039,N_7951);
or U12255 (N_12255,N_7750,N_6684);
or U12256 (N_12256,N_5358,N_7053);
nand U12257 (N_12257,N_6537,N_9352);
nand U12258 (N_12258,N_8802,N_6515);
nand U12259 (N_12259,N_6804,N_5008);
nor U12260 (N_12260,N_9791,N_5415);
or U12261 (N_12261,N_8311,N_6267);
or U12262 (N_12262,N_7722,N_7745);
nand U12263 (N_12263,N_5362,N_6063);
nor U12264 (N_12264,N_8656,N_5916);
nor U12265 (N_12265,N_5030,N_8811);
nor U12266 (N_12266,N_7477,N_8387);
and U12267 (N_12267,N_8999,N_6530);
xnor U12268 (N_12268,N_7938,N_9105);
and U12269 (N_12269,N_6742,N_8082);
and U12270 (N_12270,N_8066,N_6960);
nand U12271 (N_12271,N_5125,N_7117);
nand U12272 (N_12272,N_9437,N_9743);
or U12273 (N_12273,N_5220,N_8661);
nor U12274 (N_12274,N_9370,N_8554);
or U12275 (N_12275,N_6565,N_6276);
nand U12276 (N_12276,N_8269,N_6091);
xnor U12277 (N_12277,N_6917,N_6541);
and U12278 (N_12278,N_9287,N_8819);
and U12279 (N_12279,N_8400,N_8604);
nor U12280 (N_12280,N_9849,N_6193);
nand U12281 (N_12281,N_7203,N_5266);
or U12282 (N_12282,N_5027,N_7304);
nand U12283 (N_12283,N_5847,N_8359);
nor U12284 (N_12284,N_5759,N_5595);
nor U12285 (N_12285,N_9916,N_8060);
xor U12286 (N_12286,N_7466,N_9180);
and U12287 (N_12287,N_6797,N_9443);
or U12288 (N_12288,N_5815,N_8008);
or U12289 (N_12289,N_9623,N_5084);
and U12290 (N_12290,N_6634,N_9528);
nand U12291 (N_12291,N_8617,N_5107);
nor U12292 (N_12292,N_9821,N_5402);
and U12293 (N_12293,N_8615,N_7113);
and U12294 (N_12294,N_8193,N_7753);
or U12295 (N_12295,N_6465,N_5993);
xnor U12296 (N_12296,N_5881,N_7826);
nor U12297 (N_12297,N_5178,N_5048);
nand U12298 (N_12298,N_7489,N_6767);
or U12299 (N_12299,N_9720,N_8480);
and U12300 (N_12300,N_6647,N_7365);
or U12301 (N_12301,N_9572,N_7684);
nor U12302 (N_12302,N_8052,N_7469);
nor U12303 (N_12303,N_7985,N_9509);
xor U12304 (N_12304,N_6898,N_5808);
nand U12305 (N_12305,N_5544,N_8197);
nand U12306 (N_12306,N_8352,N_8633);
xnor U12307 (N_12307,N_9637,N_9921);
xor U12308 (N_12308,N_8143,N_6075);
and U12309 (N_12309,N_7718,N_5285);
nand U12310 (N_12310,N_7601,N_6084);
xnor U12311 (N_12311,N_7154,N_5278);
xnor U12312 (N_12312,N_9956,N_6753);
or U12313 (N_12313,N_9325,N_6014);
nor U12314 (N_12314,N_6058,N_7000);
nor U12315 (N_12315,N_9587,N_6845);
nor U12316 (N_12316,N_8734,N_7819);
nand U12317 (N_12317,N_8738,N_6098);
xnor U12318 (N_12318,N_6803,N_6816);
or U12319 (N_12319,N_5676,N_5985);
or U12320 (N_12320,N_8356,N_7378);
or U12321 (N_12321,N_6880,N_9881);
nor U12322 (N_12322,N_7852,N_6671);
nand U12323 (N_12323,N_7457,N_7595);
and U12324 (N_12324,N_7915,N_7342);
and U12325 (N_12325,N_8894,N_5307);
and U12326 (N_12326,N_5243,N_6247);
nand U12327 (N_12327,N_5142,N_7902);
nor U12328 (N_12328,N_5734,N_6997);
and U12329 (N_12329,N_5631,N_5097);
nand U12330 (N_12330,N_5606,N_7042);
and U12331 (N_12331,N_8711,N_7369);
nand U12332 (N_12332,N_9737,N_6083);
xor U12333 (N_12333,N_9910,N_6086);
nand U12334 (N_12334,N_9779,N_5656);
nor U12335 (N_12335,N_5814,N_7533);
xnor U12336 (N_12336,N_7863,N_8203);
nor U12337 (N_12337,N_9204,N_5400);
nor U12338 (N_12338,N_7338,N_8879);
or U12339 (N_12339,N_8033,N_5910);
xnor U12340 (N_12340,N_7140,N_6504);
nand U12341 (N_12341,N_8978,N_6028);
and U12342 (N_12342,N_9035,N_9713);
and U12343 (N_12343,N_7329,N_7678);
xor U12344 (N_12344,N_6833,N_9537);
nor U12345 (N_12345,N_7386,N_8539);
and U12346 (N_12346,N_8135,N_5410);
or U12347 (N_12347,N_5150,N_5947);
nand U12348 (N_12348,N_9060,N_6149);
and U12349 (N_12349,N_5346,N_8803);
or U12350 (N_12350,N_5357,N_5509);
xnor U12351 (N_12351,N_5889,N_6566);
xnor U12352 (N_12352,N_5272,N_8657);
or U12353 (N_12353,N_6170,N_9039);
and U12354 (N_12354,N_8814,N_9988);
nand U12355 (N_12355,N_5775,N_5748);
nor U12356 (N_12356,N_9497,N_6648);
nand U12357 (N_12357,N_6821,N_8552);
and U12358 (N_12358,N_7526,N_9964);
nand U12359 (N_12359,N_8845,N_8726);
nor U12360 (N_12360,N_6263,N_9019);
or U12361 (N_12361,N_6283,N_5283);
or U12362 (N_12362,N_5349,N_8496);
or U12363 (N_12363,N_6814,N_8597);
and U12364 (N_12364,N_8751,N_6987);
xnor U12365 (N_12365,N_5790,N_7235);
nor U12366 (N_12366,N_5487,N_6725);
or U12367 (N_12367,N_8472,N_5092);
nor U12368 (N_12368,N_9601,N_6363);
xor U12369 (N_12369,N_6143,N_9482);
or U12370 (N_12370,N_5100,N_9498);
nor U12371 (N_12371,N_9122,N_9520);
or U12372 (N_12372,N_7846,N_6310);
nand U12373 (N_12373,N_8874,N_8769);
nand U12374 (N_12374,N_9773,N_6035);
or U12375 (N_12375,N_9765,N_5314);
nand U12376 (N_12376,N_5552,N_9774);
xnor U12377 (N_12377,N_9028,N_7788);
xor U12378 (N_12378,N_9408,N_5094);
nor U12379 (N_12379,N_9098,N_5193);
xor U12380 (N_12380,N_8419,N_7449);
or U12381 (N_12381,N_5905,N_8742);
and U12382 (N_12382,N_5684,N_8263);
nand U12383 (N_12383,N_9036,N_6956);
nand U12384 (N_12384,N_8517,N_7427);
and U12385 (N_12385,N_7712,N_9754);
and U12386 (N_12386,N_7534,N_8639);
nor U12387 (N_12387,N_7079,N_7036);
xor U12388 (N_12388,N_8454,N_8990);
nor U12389 (N_12389,N_8781,N_7474);
nor U12390 (N_12390,N_7319,N_7699);
nand U12391 (N_12391,N_8938,N_5132);
and U12392 (N_12392,N_9257,N_9417);
nor U12393 (N_12393,N_8219,N_5454);
and U12394 (N_12394,N_8370,N_6641);
and U12395 (N_12395,N_6021,N_6918);
or U12396 (N_12396,N_9286,N_5887);
and U12397 (N_12397,N_5148,N_9358);
nand U12398 (N_12398,N_6025,N_6474);
and U12399 (N_12399,N_5868,N_5615);
and U12400 (N_12400,N_7646,N_7303);
nand U12401 (N_12401,N_8195,N_9775);
or U12402 (N_12402,N_5530,N_9523);
xnor U12403 (N_12403,N_5586,N_5022);
nor U12404 (N_12404,N_9418,N_6000);
nor U12405 (N_12405,N_9628,N_5998);
or U12406 (N_12406,N_5745,N_7914);
nor U12407 (N_12407,N_9465,N_9753);
nor U12408 (N_12408,N_9367,N_7961);
or U12409 (N_12409,N_9567,N_5773);
and U12410 (N_12410,N_5504,N_8150);
nand U12411 (N_12411,N_6676,N_6683);
or U12412 (N_12412,N_9012,N_5422);
or U12413 (N_12413,N_9277,N_8535);
nand U12414 (N_12414,N_8603,N_5831);
and U12415 (N_12415,N_5365,N_5041);
nor U12416 (N_12416,N_7208,N_6024);
nor U12417 (N_12417,N_6101,N_7020);
xor U12418 (N_12418,N_5811,N_5031);
nand U12419 (N_12419,N_8559,N_7276);
and U12420 (N_12420,N_5991,N_6492);
nand U12421 (N_12421,N_8448,N_5965);
nand U12422 (N_12422,N_8659,N_9527);
or U12423 (N_12423,N_9920,N_7167);
and U12424 (N_12424,N_5555,N_7244);
and U12425 (N_12425,N_7797,N_8940);
or U12426 (N_12426,N_8928,N_8037);
or U12427 (N_12427,N_6409,N_6991);
nor U12428 (N_12428,N_5511,N_6747);
or U12429 (N_12429,N_7927,N_9857);
nand U12430 (N_12430,N_7769,N_9441);
xor U12431 (N_12431,N_6116,N_8228);
nor U12432 (N_12432,N_5233,N_6669);
and U12433 (N_12433,N_8695,N_6077);
nand U12434 (N_12434,N_7709,N_8038);
nor U12435 (N_12435,N_5282,N_8693);
and U12436 (N_12436,N_9351,N_8528);
or U12437 (N_12437,N_8177,N_7925);
xnor U12438 (N_12438,N_8183,N_8491);
or U12439 (N_12439,N_7357,N_7954);
nor U12440 (N_12440,N_8829,N_6060);
nand U12441 (N_12441,N_8478,N_6374);
and U12442 (N_12442,N_8110,N_9311);
or U12443 (N_12443,N_7016,N_9975);
xnor U12444 (N_12444,N_8181,N_7658);
nor U12445 (N_12445,N_5195,N_9874);
or U12446 (N_12446,N_6774,N_7195);
or U12447 (N_12447,N_9938,N_5501);
nor U12448 (N_12448,N_8459,N_5213);
or U12449 (N_12449,N_5937,N_8420);
and U12450 (N_12450,N_6278,N_9205);
nor U12451 (N_12451,N_7522,N_8036);
nand U12452 (N_12452,N_9384,N_9627);
nor U12453 (N_12453,N_9908,N_7764);
and U12454 (N_12454,N_8122,N_5678);
nand U12455 (N_12455,N_7924,N_6142);
and U12456 (N_12456,N_7901,N_8105);
or U12457 (N_12457,N_5579,N_5064);
nor U12458 (N_12458,N_5999,N_6552);
nand U12459 (N_12459,N_6311,N_8471);
and U12460 (N_12460,N_9966,N_6505);
or U12461 (N_12461,N_9229,N_8139);
nand U12462 (N_12462,N_6954,N_6199);
and U12463 (N_12463,N_8683,N_9044);
nor U12464 (N_12464,N_5981,N_7643);
and U12465 (N_12465,N_9620,N_7152);
and U12466 (N_12466,N_8494,N_7312);
nor U12467 (N_12467,N_6624,N_7947);
nor U12468 (N_12468,N_9522,N_7216);
and U12469 (N_12469,N_8191,N_8446);
nor U12470 (N_12470,N_9055,N_9671);
nor U12471 (N_12471,N_8463,N_7894);
nor U12472 (N_12472,N_9425,N_5482);
nand U12473 (N_12473,N_6361,N_5396);
nor U12474 (N_12474,N_9855,N_7364);
or U12475 (N_12475,N_6657,N_6271);
nand U12476 (N_12476,N_9980,N_6784);
nand U12477 (N_12477,N_9722,N_6417);
nor U12478 (N_12478,N_6428,N_6141);
nand U12479 (N_12479,N_8497,N_9944);
xor U12480 (N_12480,N_5024,N_5578);
nand U12481 (N_12481,N_5569,N_9948);
nor U12482 (N_12482,N_8487,N_9600);
nand U12483 (N_12483,N_5607,N_6139);
and U12484 (N_12484,N_8407,N_5959);
nand U12485 (N_12485,N_9353,N_6679);
nor U12486 (N_12486,N_9870,N_9986);
nand U12487 (N_12487,N_7696,N_7967);
and U12488 (N_12488,N_6034,N_9142);
nand U12489 (N_12489,N_8679,N_5475);
xor U12490 (N_12490,N_5860,N_9937);
or U12491 (N_12491,N_8766,N_7032);
and U12492 (N_12492,N_5021,N_5199);
nor U12493 (N_12493,N_7346,N_9102);
or U12494 (N_12494,N_5177,N_7995);
and U12495 (N_12495,N_6600,N_6134);
and U12496 (N_12496,N_8908,N_7229);
nand U12497 (N_12497,N_5878,N_5955);
nor U12498 (N_12498,N_7052,N_8885);
or U12499 (N_12499,N_7836,N_8458);
and U12500 (N_12500,N_8681,N_5547);
and U12501 (N_12501,N_7485,N_8425);
nor U12502 (N_12502,N_8407,N_8967);
or U12503 (N_12503,N_6302,N_6069);
or U12504 (N_12504,N_7048,N_8929);
or U12505 (N_12505,N_5131,N_5765);
and U12506 (N_12506,N_6691,N_5741);
nand U12507 (N_12507,N_9982,N_5301);
xor U12508 (N_12508,N_9421,N_8293);
and U12509 (N_12509,N_5804,N_8759);
nor U12510 (N_12510,N_8071,N_8537);
and U12511 (N_12511,N_5635,N_8818);
xor U12512 (N_12512,N_7958,N_5385);
and U12513 (N_12513,N_8724,N_7718);
xnor U12514 (N_12514,N_7015,N_5183);
nor U12515 (N_12515,N_5135,N_7392);
or U12516 (N_12516,N_6473,N_9848);
or U12517 (N_12517,N_9142,N_7624);
or U12518 (N_12518,N_5494,N_8172);
nand U12519 (N_12519,N_5893,N_5448);
nand U12520 (N_12520,N_9928,N_9665);
nor U12521 (N_12521,N_5429,N_7527);
xnor U12522 (N_12522,N_8531,N_7824);
or U12523 (N_12523,N_8494,N_9626);
xor U12524 (N_12524,N_6254,N_5519);
nand U12525 (N_12525,N_7336,N_9479);
or U12526 (N_12526,N_9982,N_7854);
nor U12527 (N_12527,N_5644,N_7094);
nor U12528 (N_12528,N_8591,N_7250);
and U12529 (N_12529,N_8745,N_6974);
nor U12530 (N_12530,N_8317,N_8727);
nand U12531 (N_12531,N_5732,N_6275);
nand U12532 (N_12532,N_8121,N_8572);
nand U12533 (N_12533,N_5183,N_5813);
nor U12534 (N_12534,N_8847,N_9374);
and U12535 (N_12535,N_8251,N_7246);
nand U12536 (N_12536,N_7182,N_9925);
nand U12537 (N_12537,N_9872,N_8115);
or U12538 (N_12538,N_5270,N_9345);
and U12539 (N_12539,N_5014,N_5678);
and U12540 (N_12540,N_7428,N_6434);
nor U12541 (N_12541,N_7283,N_6352);
and U12542 (N_12542,N_7874,N_6168);
and U12543 (N_12543,N_6710,N_6327);
or U12544 (N_12544,N_7317,N_6124);
or U12545 (N_12545,N_9845,N_7550);
and U12546 (N_12546,N_9932,N_9044);
or U12547 (N_12547,N_6564,N_9089);
or U12548 (N_12548,N_5475,N_8648);
xnor U12549 (N_12549,N_9765,N_9778);
nand U12550 (N_12550,N_9858,N_8596);
and U12551 (N_12551,N_7859,N_9313);
and U12552 (N_12552,N_7737,N_8051);
or U12553 (N_12553,N_6934,N_9479);
and U12554 (N_12554,N_7536,N_7235);
nor U12555 (N_12555,N_5023,N_6894);
nor U12556 (N_12556,N_6224,N_7306);
nor U12557 (N_12557,N_9974,N_5794);
and U12558 (N_12558,N_9464,N_8519);
or U12559 (N_12559,N_8986,N_9358);
or U12560 (N_12560,N_6048,N_8368);
xor U12561 (N_12561,N_9551,N_6845);
xor U12562 (N_12562,N_5827,N_7998);
nor U12563 (N_12563,N_7681,N_8728);
nor U12564 (N_12564,N_8023,N_8960);
and U12565 (N_12565,N_7208,N_6189);
and U12566 (N_12566,N_6250,N_8315);
and U12567 (N_12567,N_5675,N_9685);
nand U12568 (N_12568,N_7683,N_7110);
and U12569 (N_12569,N_6381,N_8848);
or U12570 (N_12570,N_6122,N_9594);
nor U12571 (N_12571,N_5001,N_7264);
or U12572 (N_12572,N_7341,N_8998);
xor U12573 (N_12573,N_8961,N_8091);
nand U12574 (N_12574,N_9838,N_7271);
nor U12575 (N_12575,N_5634,N_5744);
nand U12576 (N_12576,N_5729,N_5003);
nor U12577 (N_12577,N_9783,N_9697);
or U12578 (N_12578,N_7482,N_7803);
nand U12579 (N_12579,N_8412,N_9397);
xor U12580 (N_12580,N_7359,N_6131);
or U12581 (N_12581,N_5822,N_8294);
and U12582 (N_12582,N_7639,N_7655);
nand U12583 (N_12583,N_7236,N_9003);
and U12584 (N_12584,N_5775,N_7802);
or U12585 (N_12585,N_8512,N_7458);
xor U12586 (N_12586,N_9761,N_5886);
nor U12587 (N_12587,N_5472,N_6313);
nand U12588 (N_12588,N_8475,N_8648);
or U12589 (N_12589,N_6134,N_5641);
or U12590 (N_12590,N_5981,N_8937);
xor U12591 (N_12591,N_9290,N_5374);
and U12592 (N_12592,N_9317,N_5913);
or U12593 (N_12593,N_7929,N_6304);
xnor U12594 (N_12594,N_6975,N_5007);
and U12595 (N_12595,N_7696,N_9969);
and U12596 (N_12596,N_5845,N_7914);
or U12597 (N_12597,N_8622,N_7545);
nand U12598 (N_12598,N_7431,N_6106);
and U12599 (N_12599,N_9560,N_7172);
nor U12600 (N_12600,N_9911,N_5380);
nand U12601 (N_12601,N_7078,N_9658);
and U12602 (N_12602,N_8250,N_6959);
nor U12603 (N_12603,N_8210,N_7114);
and U12604 (N_12604,N_7143,N_6538);
or U12605 (N_12605,N_8503,N_6236);
or U12606 (N_12606,N_6998,N_6779);
nand U12607 (N_12607,N_7215,N_7955);
nor U12608 (N_12608,N_6352,N_6363);
or U12609 (N_12609,N_8994,N_8862);
or U12610 (N_12610,N_5678,N_7338);
xor U12611 (N_12611,N_7643,N_8812);
nand U12612 (N_12612,N_5069,N_9623);
nor U12613 (N_12613,N_6678,N_5635);
or U12614 (N_12614,N_6540,N_8084);
nor U12615 (N_12615,N_6596,N_7643);
and U12616 (N_12616,N_6388,N_6474);
and U12617 (N_12617,N_8866,N_5773);
or U12618 (N_12618,N_8004,N_5076);
and U12619 (N_12619,N_8772,N_9877);
or U12620 (N_12620,N_9358,N_9671);
nand U12621 (N_12621,N_5842,N_5508);
nor U12622 (N_12622,N_8826,N_5254);
xnor U12623 (N_12623,N_9463,N_7826);
or U12624 (N_12624,N_9265,N_9864);
xor U12625 (N_12625,N_5308,N_6773);
nor U12626 (N_12626,N_8422,N_6815);
or U12627 (N_12627,N_5635,N_8929);
nand U12628 (N_12628,N_7799,N_9883);
and U12629 (N_12629,N_8889,N_5535);
and U12630 (N_12630,N_7213,N_7593);
nor U12631 (N_12631,N_9712,N_7898);
xor U12632 (N_12632,N_7517,N_6585);
or U12633 (N_12633,N_6035,N_5355);
nand U12634 (N_12634,N_6280,N_9220);
nor U12635 (N_12635,N_8338,N_9864);
xnor U12636 (N_12636,N_6629,N_6451);
nand U12637 (N_12637,N_5227,N_7322);
or U12638 (N_12638,N_6691,N_8986);
or U12639 (N_12639,N_8224,N_9376);
nor U12640 (N_12640,N_7028,N_7531);
nor U12641 (N_12641,N_7205,N_7996);
and U12642 (N_12642,N_6787,N_7231);
nor U12643 (N_12643,N_8596,N_9814);
nor U12644 (N_12644,N_9275,N_6574);
and U12645 (N_12645,N_8030,N_6205);
and U12646 (N_12646,N_5843,N_6507);
xnor U12647 (N_12647,N_5781,N_5120);
and U12648 (N_12648,N_6039,N_6196);
and U12649 (N_12649,N_8949,N_8187);
nand U12650 (N_12650,N_5566,N_8319);
nor U12651 (N_12651,N_6814,N_7552);
xor U12652 (N_12652,N_7089,N_9513);
or U12653 (N_12653,N_5881,N_5051);
or U12654 (N_12654,N_5201,N_7863);
xnor U12655 (N_12655,N_9175,N_7480);
and U12656 (N_12656,N_7072,N_6713);
xnor U12657 (N_12657,N_7229,N_5983);
or U12658 (N_12658,N_7031,N_7402);
nor U12659 (N_12659,N_8089,N_9498);
or U12660 (N_12660,N_8880,N_5191);
nor U12661 (N_12661,N_9653,N_7844);
nand U12662 (N_12662,N_5806,N_8639);
or U12663 (N_12663,N_5773,N_8674);
and U12664 (N_12664,N_9137,N_7716);
and U12665 (N_12665,N_6773,N_5125);
and U12666 (N_12666,N_6146,N_5083);
nor U12667 (N_12667,N_6799,N_8039);
and U12668 (N_12668,N_7751,N_8781);
nor U12669 (N_12669,N_6038,N_9810);
nor U12670 (N_12670,N_8493,N_6001);
nand U12671 (N_12671,N_8350,N_7877);
xnor U12672 (N_12672,N_5760,N_6203);
and U12673 (N_12673,N_7543,N_6951);
nor U12674 (N_12674,N_8896,N_7302);
nor U12675 (N_12675,N_5902,N_7748);
nand U12676 (N_12676,N_7138,N_5976);
nand U12677 (N_12677,N_5033,N_7913);
xnor U12678 (N_12678,N_8249,N_5442);
nand U12679 (N_12679,N_6668,N_9928);
nand U12680 (N_12680,N_9007,N_8233);
or U12681 (N_12681,N_8598,N_9241);
xnor U12682 (N_12682,N_7991,N_5102);
nand U12683 (N_12683,N_5872,N_5660);
nor U12684 (N_12684,N_7548,N_7323);
and U12685 (N_12685,N_9559,N_6615);
and U12686 (N_12686,N_6649,N_7940);
xor U12687 (N_12687,N_8571,N_8477);
nand U12688 (N_12688,N_6462,N_7541);
nor U12689 (N_12689,N_5355,N_8211);
or U12690 (N_12690,N_6964,N_6220);
and U12691 (N_12691,N_7526,N_7541);
nand U12692 (N_12692,N_9832,N_5647);
nor U12693 (N_12693,N_8873,N_9451);
nand U12694 (N_12694,N_7007,N_9421);
nor U12695 (N_12695,N_8178,N_8403);
or U12696 (N_12696,N_9956,N_9284);
nor U12697 (N_12697,N_7605,N_6736);
and U12698 (N_12698,N_6719,N_9333);
xor U12699 (N_12699,N_5066,N_5752);
xnor U12700 (N_12700,N_7913,N_6894);
nand U12701 (N_12701,N_7146,N_9716);
or U12702 (N_12702,N_7881,N_8985);
or U12703 (N_12703,N_7347,N_7053);
xor U12704 (N_12704,N_9964,N_5273);
xor U12705 (N_12705,N_9356,N_6785);
and U12706 (N_12706,N_5806,N_9913);
or U12707 (N_12707,N_7155,N_9990);
and U12708 (N_12708,N_5920,N_5459);
nand U12709 (N_12709,N_5518,N_7806);
or U12710 (N_12710,N_5909,N_5424);
nor U12711 (N_12711,N_5665,N_9650);
and U12712 (N_12712,N_8136,N_6830);
xor U12713 (N_12713,N_9559,N_9356);
and U12714 (N_12714,N_9505,N_9389);
nor U12715 (N_12715,N_7455,N_7278);
and U12716 (N_12716,N_5833,N_8382);
nor U12717 (N_12717,N_9612,N_8056);
nand U12718 (N_12718,N_6485,N_7397);
and U12719 (N_12719,N_9385,N_9441);
and U12720 (N_12720,N_6315,N_6323);
or U12721 (N_12721,N_8913,N_6240);
xnor U12722 (N_12722,N_8480,N_8798);
xnor U12723 (N_12723,N_7770,N_7329);
nand U12724 (N_12724,N_9350,N_8108);
nor U12725 (N_12725,N_5762,N_6020);
and U12726 (N_12726,N_6677,N_6800);
nand U12727 (N_12727,N_7560,N_8888);
nand U12728 (N_12728,N_7571,N_8370);
xor U12729 (N_12729,N_6382,N_5385);
or U12730 (N_12730,N_5968,N_6021);
or U12731 (N_12731,N_7741,N_5287);
or U12732 (N_12732,N_6483,N_9641);
nor U12733 (N_12733,N_7021,N_9615);
nor U12734 (N_12734,N_6836,N_9969);
or U12735 (N_12735,N_9075,N_6450);
nor U12736 (N_12736,N_6756,N_6880);
or U12737 (N_12737,N_8783,N_9441);
and U12738 (N_12738,N_7322,N_5968);
xor U12739 (N_12739,N_6430,N_7978);
and U12740 (N_12740,N_7432,N_9554);
and U12741 (N_12741,N_9712,N_8329);
and U12742 (N_12742,N_7349,N_6107);
or U12743 (N_12743,N_9136,N_7665);
and U12744 (N_12744,N_5632,N_6352);
or U12745 (N_12745,N_7871,N_7768);
nor U12746 (N_12746,N_6106,N_5574);
nor U12747 (N_12747,N_9956,N_7590);
nand U12748 (N_12748,N_8996,N_5236);
and U12749 (N_12749,N_6288,N_7705);
or U12750 (N_12750,N_7019,N_5116);
nand U12751 (N_12751,N_5299,N_9394);
nor U12752 (N_12752,N_6852,N_5547);
nor U12753 (N_12753,N_9204,N_8473);
nand U12754 (N_12754,N_6693,N_9655);
nor U12755 (N_12755,N_6257,N_5882);
or U12756 (N_12756,N_7880,N_6233);
or U12757 (N_12757,N_9111,N_6188);
xnor U12758 (N_12758,N_7516,N_6726);
and U12759 (N_12759,N_9376,N_8103);
or U12760 (N_12760,N_7234,N_5214);
or U12761 (N_12761,N_6247,N_8248);
or U12762 (N_12762,N_9491,N_9471);
nor U12763 (N_12763,N_6902,N_7526);
and U12764 (N_12764,N_5407,N_5792);
and U12765 (N_12765,N_8610,N_6000);
or U12766 (N_12766,N_8760,N_9605);
nand U12767 (N_12767,N_9083,N_6426);
or U12768 (N_12768,N_7040,N_6275);
or U12769 (N_12769,N_6947,N_9116);
or U12770 (N_12770,N_5563,N_5378);
or U12771 (N_12771,N_7766,N_6518);
or U12772 (N_12772,N_5897,N_8902);
or U12773 (N_12773,N_9047,N_8499);
and U12774 (N_12774,N_5864,N_5348);
nor U12775 (N_12775,N_8614,N_6294);
nand U12776 (N_12776,N_5306,N_7883);
and U12777 (N_12777,N_9243,N_6086);
xnor U12778 (N_12778,N_6932,N_9067);
or U12779 (N_12779,N_6875,N_5889);
nor U12780 (N_12780,N_7342,N_5853);
nand U12781 (N_12781,N_5644,N_6153);
nand U12782 (N_12782,N_7373,N_6641);
nor U12783 (N_12783,N_7529,N_5349);
nand U12784 (N_12784,N_8925,N_5249);
and U12785 (N_12785,N_5396,N_9120);
nand U12786 (N_12786,N_7360,N_8839);
or U12787 (N_12787,N_9730,N_6112);
and U12788 (N_12788,N_6039,N_5526);
and U12789 (N_12789,N_9978,N_8219);
and U12790 (N_12790,N_7099,N_6877);
nand U12791 (N_12791,N_6217,N_7425);
nand U12792 (N_12792,N_6665,N_8568);
nand U12793 (N_12793,N_7970,N_7646);
and U12794 (N_12794,N_6928,N_6185);
xnor U12795 (N_12795,N_5219,N_5244);
and U12796 (N_12796,N_7441,N_6035);
xnor U12797 (N_12797,N_9675,N_6986);
and U12798 (N_12798,N_7716,N_9649);
or U12799 (N_12799,N_8735,N_5950);
or U12800 (N_12800,N_6543,N_7457);
xnor U12801 (N_12801,N_7353,N_9819);
or U12802 (N_12802,N_9560,N_5773);
or U12803 (N_12803,N_7080,N_5293);
xnor U12804 (N_12804,N_9358,N_6190);
and U12805 (N_12805,N_9482,N_6357);
nand U12806 (N_12806,N_7784,N_8582);
nor U12807 (N_12807,N_5026,N_9329);
or U12808 (N_12808,N_7781,N_6527);
or U12809 (N_12809,N_9094,N_5217);
and U12810 (N_12810,N_7090,N_5510);
nor U12811 (N_12811,N_7936,N_6510);
nand U12812 (N_12812,N_5223,N_9319);
nand U12813 (N_12813,N_9135,N_9057);
or U12814 (N_12814,N_9037,N_7541);
nand U12815 (N_12815,N_9296,N_8074);
xor U12816 (N_12816,N_7791,N_7632);
and U12817 (N_12817,N_5720,N_7746);
nand U12818 (N_12818,N_7657,N_6115);
nand U12819 (N_12819,N_5442,N_8971);
or U12820 (N_12820,N_6915,N_9202);
nand U12821 (N_12821,N_7001,N_6239);
or U12822 (N_12822,N_7795,N_7947);
nand U12823 (N_12823,N_8453,N_6484);
and U12824 (N_12824,N_5888,N_8908);
and U12825 (N_12825,N_5252,N_9950);
or U12826 (N_12826,N_5235,N_8843);
nand U12827 (N_12827,N_6886,N_7616);
xnor U12828 (N_12828,N_8016,N_7755);
and U12829 (N_12829,N_6062,N_8382);
or U12830 (N_12830,N_7355,N_5273);
and U12831 (N_12831,N_6002,N_7959);
nand U12832 (N_12832,N_5778,N_8087);
or U12833 (N_12833,N_5471,N_6148);
xnor U12834 (N_12834,N_8216,N_6038);
nand U12835 (N_12835,N_8088,N_6637);
nor U12836 (N_12836,N_7788,N_9081);
or U12837 (N_12837,N_6301,N_6036);
and U12838 (N_12838,N_9014,N_7557);
or U12839 (N_12839,N_9746,N_6005);
nor U12840 (N_12840,N_7677,N_5516);
or U12841 (N_12841,N_5007,N_6457);
nor U12842 (N_12842,N_7285,N_9806);
and U12843 (N_12843,N_7478,N_9849);
nor U12844 (N_12844,N_9755,N_8834);
and U12845 (N_12845,N_5368,N_9715);
nand U12846 (N_12846,N_6826,N_7584);
and U12847 (N_12847,N_6349,N_7295);
nand U12848 (N_12848,N_6435,N_7498);
and U12849 (N_12849,N_7020,N_9138);
nor U12850 (N_12850,N_8795,N_5628);
or U12851 (N_12851,N_6279,N_9525);
or U12852 (N_12852,N_8803,N_9428);
or U12853 (N_12853,N_7140,N_7400);
xnor U12854 (N_12854,N_5538,N_8950);
xor U12855 (N_12855,N_9994,N_9204);
and U12856 (N_12856,N_5052,N_7529);
nand U12857 (N_12857,N_7096,N_6840);
and U12858 (N_12858,N_6302,N_8899);
nand U12859 (N_12859,N_7880,N_6068);
nor U12860 (N_12860,N_7094,N_8557);
nor U12861 (N_12861,N_5477,N_5077);
nand U12862 (N_12862,N_7028,N_8984);
xor U12863 (N_12863,N_9665,N_5722);
xor U12864 (N_12864,N_6386,N_5346);
nand U12865 (N_12865,N_5787,N_8877);
and U12866 (N_12866,N_8697,N_8414);
nand U12867 (N_12867,N_8691,N_9192);
and U12868 (N_12868,N_6448,N_5233);
nor U12869 (N_12869,N_6946,N_7925);
and U12870 (N_12870,N_5551,N_8177);
and U12871 (N_12871,N_6193,N_9490);
nand U12872 (N_12872,N_9709,N_5154);
nand U12873 (N_12873,N_6439,N_5761);
nand U12874 (N_12874,N_8001,N_5713);
nor U12875 (N_12875,N_8768,N_9944);
or U12876 (N_12876,N_6868,N_8694);
nand U12877 (N_12877,N_8040,N_6294);
nand U12878 (N_12878,N_5047,N_5050);
and U12879 (N_12879,N_5916,N_7465);
nor U12880 (N_12880,N_7811,N_9281);
and U12881 (N_12881,N_6352,N_9854);
nand U12882 (N_12882,N_8463,N_9179);
nand U12883 (N_12883,N_6235,N_6848);
nand U12884 (N_12884,N_9691,N_5021);
nor U12885 (N_12885,N_5182,N_6731);
nor U12886 (N_12886,N_9753,N_6822);
nor U12887 (N_12887,N_8463,N_6536);
or U12888 (N_12888,N_8096,N_9521);
and U12889 (N_12889,N_9709,N_8853);
nor U12890 (N_12890,N_7161,N_5178);
and U12891 (N_12891,N_9072,N_5808);
or U12892 (N_12892,N_6904,N_7582);
nor U12893 (N_12893,N_7542,N_9000);
nor U12894 (N_12894,N_9698,N_7529);
xnor U12895 (N_12895,N_8683,N_5611);
and U12896 (N_12896,N_6297,N_8611);
and U12897 (N_12897,N_5099,N_9837);
or U12898 (N_12898,N_9415,N_9809);
or U12899 (N_12899,N_5603,N_5533);
nor U12900 (N_12900,N_7169,N_8211);
and U12901 (N_12901,N_9475,N_6764);
nor U12902 (N_12902,N_8862,N_9541);
and U12903 (N_12903,N_8108,N_9388);
nor U12904 (N_12904,N_7380,N_6425);
or U12905 (N_12905,N_5150,N_7328);
nor U12906 (N_12906,N_5884,N_9625);
nor U12907 (N_12907,N_6648,N_7193);
and U12908 (N_12908,N_7744,N_5374);
nor U12909 (N_12909,N_7304,N_8099);
or U12910 (N_12910,N_7808,N_7374);
nand U12911 (N_12911,N_7718,N_5935);
nor U12912 (N_12912,N_9979,N_7288);
nand U12913 (N_12913,N_8141,N_8252);
nor U12914 (N_12914,N_7404,N_8213);
and U12915 (N_12915,N_8757,N_8387);
nor U12916 (N_12916,N_7340,N_6220);
nor U12917 (N_12917,N_6976,N_5880);
and U12918 (N_12918,N_8654,N_8570);
nand U12919 (N_12919,N_9230,N_6061);
nor U12920 (N_12920,N_8278,N_8354);
nor U12921 (N_12921,N_6487,N_5991);
or U12922 (N_12922,N_6189,N_5059);
nand U12923 (N_12923,N_6111,N_7103);
or U12924 (N_12924,N_7056,N_9762);
nor U12925 (N_12925,N_9866,N_5267);
and U12926 (N_12926,N_5111,N_8478);
and U12927 (N_12927,N_7033,N_6502);
or U12928 (N_12928,N_5500,N_7991);
nor U12929 (N_12929,N_6929,N_8947);
or U12930 (N_12930,N_9390,N_8531);
and U12931 (N_12931,N_5420,N_9335);
nor U12932 (N_12932,N_8687,N_5106);
nor U12933 (N_12933,N_8791,N_7503);
nand U12934 (N_12934,N_6965,N_8112);
nor U12935 (N_12935,N_8661,N_9777);
xnor U12936 (N_12936,N_8313,N_6684);
xnor U12937 (N_12937,N_8491,N_7743);
nor U12938 (N_12938,N_6286,N_7144);
nor U12939 (N_12939,N_5388,N_7210);
nand U12940 (N_12940,N_6298,N_9338);
and U12941 (N_12941,N_5554,N_9854);
and U12942 (N_12942,N_7801,N_6603);
and U12943 (N_12943,N_7003,N_5833);
nand U12944 (N_12944,N_9920,N_6267);
or U12945 (N_12945,N_9953,N_8726);
nor U12946 (N_12946,N_5795,N_9100);
or U12947 (N_12947,N_9207,N_5418);
xnor U12948 (N_12948,N_6348,N_7814);
nand U12949 (N_12949,N_6035,N_7309);
and U12950 (N_12950,N_8115,N_6112);
nor U12951 (N_12951,N_7617,N_5691);
or U12952 (N_12952,N_5632,N_9455);
and U12953 (N_12953,N_8925,N_7219);
nand U12954 (N_12954,N_9956,N_5439);
or U12955 (N_12955,N_9814,N_9393);
nand U12956 (N_12956,N_6673,N_9619);
or U12957 (N_12957,N_7605,N_7748);
or U12958 (N_12958,N_5222,N_5752);
nand U12959 (N_12959,N_6965,N_7165);
or U12960 (N_12960,N_9691,N_8495);
nand U12961 (N_12961,N_6550,N_8585);
nor U12962 (N_12962,N_5890,N_5340);
xor U12963 (N_12963,N_9027,N_9890);
nand U12964 (N_12964,N_8404,N_7515);
and U12965 (N_12965,N_6422,N_8692);
nor U12966 (N_12966,N_8609,N_5209);
xor U12967 (N_12967,N_9281,N_6592);
or U12968 (N_12968,N_5501,N_8446);
or U12969 (N_12969,N_7419,N_9175);
nand U12970 (N_12970,N_6631,N_5582);
nand U12971 (N_12971,N_5203,N_5550);
and U12972 (N_12972,N_8000,N_6573);
nand U12973 (N_12973,N_8908,N_7969);
or U12974 (N_12974,N_7436,N_9547);
nor U12975 (N_12975,N_7145,N_5936);
nand U12976 (N_12976,N_5266,N_9836);
and U12977 (N_12977,N_5871,N_5487);
xnor U12978 (N_12978,N_6305,N_7507);
nand U12979 (N_12979,N_5174,N_6394);
or U12980 (N_12980,N_8980,N_6440);
nand U12981 (N_12981,N_7025,N_9109);
and U12982 (N_12982,N_5889,N_7437);
and U12983 (N_12983,N_5196,N_6884);
xnor U12984 (N_12984,N_9644,N_6203);
nor U12985 (N_12985,N_5864,N_8193);
nor U12986 (N_12986,N_8241,N_7761);
nor U12987 (N_12987,N_9799,N_9838);
nor U12988 (N_12988,N_8596,N_7767);
or U12989 (N_12989,N_9833,N_7900);
nand U12990 (N_12990,N_7408,N_6894);
xor U12991 (N_12991,N_7814,N_7524);
nor U12992 (N_12992,N_5401,N_8801);
and U12993 (N_12993,N_7416,N_9245);
or U12994 (N_12994,N_8055,N_9439);
or U12995 (N_12995,N_6832,N_9823);
nor U12996 (N_12996,N_5592,N_6636);
nand U12997 (N_12997,N_7529,N_6851);
nor U12998 (N_12998,N_8431,N_7038);
nand U12999 (N_12999,N_6086,N_5170);
or U13000 (N_13000,N_5356,N_5380);
or U13001 (N_13001,N_7016,N_6597);
or U13002 (N_13002,N_6982,N_6022);
or U13003 (N_13003,N_9249,N_6754);
xor U13004 (N_13004,N_9388,N_5323);
nand U13005 (N_13005,N_8778,N_9245);
nor U13006 (N_13006,N_7692,N_5419);
or U13007 (N_13007,N_7661,N_6008);
nor U13008 (N_13008,N_7950,N_9037);
nand U13009 (N_13009,N_7011,N_9775);
nand U13010 (N_13010,N_6271,N_5133);
nor U13011 (N_13011,N_6069,N_8953);
nor U13012 (N_13012,N_8822,N_7056);
nand U13013 (N_13013,N_8922,N_5200);
nand U13014 (N_13014,N_5798,N_8741);
nand U13015 (N_13015,N_9122,N_5511);
nand U13016 (N_13016,N_7230,N_6996);
nor U13017 (N_13017,N_9360,N_6767);
nand U13018 (N_13018,N_9275,N_8050);
nand U13019 (N_13019,N_6114,N_9863);
and U13020 (N_13020,N_7269,N_7514);
or U13021 (N_13021,N_9845,N_9257);
nor U13022 (N_13022,N_6143,N_5364);
xnor U13023 (N_13023,N_5567,N_8378);
or U13024 (N_13024,N_7354,N_7468);
nand U13025 (N_13025,N_6967,N_7613);
or U13026 (N_13026,N_7594,N_7258);
xor U13027 (N_13027,N_7255,N_8324);
or U13028 (N_13028,N_5348,N_7435);
nand U13029 (N_13029,N_6345,N_7230);
or U13030 (N_13030,N_5343,N_6811);
nor U13031 (N_13031,N_5017,N_5662);
and U13032 (N_13032,N_6269,N_6449);
or U13033 (N_13033,N_8840,N_8395);
nor U13034 (N_13034,N_9639,N_6938);
nor U13035 (N_13035,N_5927,N_5471);
or U13036 (N_13036,N_7930,N_6743);
nor U13037 (N_13037,N_7617,N_5436);
or U13038 (N_13038,N_8100,N_6397);
nand U13039 (N_13039,N_5771,N_7018);
nor U13040 (N_13040,N_8227,N_7928);
nor U13041 (N_13041,N_7337,N_8584);
and U13042 (N_13042,N_5216,N_5378);
nor U13043 (N_13043,N_6326,N_7106);
nand U13044 (N_13044,N_9514,N_8298);
nor U13045 (N_13045,N_9205,N_8908);
nor U13046 (N_13046,N_8990,N_6239);
and U13047 (N_13047,N_9965,N_5206);
and U13048 (N_13048,N_8866,N_7608);
nand U13049 (N_13049,N_5672,N_7002);
or U13050 (N_13050,N_9591,N_9973);
and U13051 (N_13051,N_7022,N_5945);
nand U13052 (N_13052,N_7869,N_8374);
xor U13053 (N_13053,N_6153,N_5580);
nand U13054 (N_13054,N_8262,N_9970);
and U13055 (N_13055,N_5624,N_6064);
nor U13056 (N_13056,N_9956,N_9830);
and U13057 (N_13057,N_9567,N_9152);
nand U13058 (N_13058,N_6995,N_8222);
or U13059 (N_13059,N_9257,N_6962);
nor U13060 (N_13060,N_5753,N_6063);
xor U13061 (N_13061,N_7623,N_7557);
or U13062 (N_13062,N_7906,N_7851);
or U13063 (N_13063,N_9872,N_6972);
nor U13064 (N_13064,N_6091,N_6727);
and U13065 (N_13065,N_7856,N_5919);
and U13066 (N_13066,N_6297,N_5831);
and U13067 (N_13067,N_8066,N_6142);
xor U13068 (N_13068,N_9165,N_9780);
xnor U13069 (N_13069,N_8486,N_7936);
nor U13070 (N_13070,N_5777,N_5869);
nand U13071 (N_13071,N_7019,N_5369);
nand U13072 (N_13072,N_7430,N_9196);
or U13073 (N_13073,N_6768,N_8360);
nand U13074 (N_13074,N_9414,N_7148);
or U13075 (N_13075,N_7125,N_6772);
nor U13076 (N_13076,N_6363,N_7905);
nand U13077 (N_13077,N_9965,N_6493);
nand U13078 (N_13078,N_7509,N_5557);
or U13079 (N_13079,N_6226,N_9863);
or U13080 (N_13080,N_9952,N_7555);
nand U13081 (N_13081,N_9813,N_8403);
nand U13082 (N_13082,N_8822,N_7471);
nand U13083 (N_13083,N_7149,N_5702);
nand U13084 (N_13084,N_7987,N_7164);
nand U13085 (N_13085,N_7086,N_7867);
nor U13086 (N_13086,N_5334,N_6427);
nor U13087 (N_13087,N_8483,N_8148);
or U13088 (N_13088,N_7017,N_6946);
xor U13089 (N_13089,N_7637,N_5124);
or U13090 (N_13090,N_8553,N_5014);
and U13091 (N_13091,N_7220,N_5927);
nor U13092 (N_13092,N_7897,N_5606);
and U13093 (N_13093,N_8418,N_6731);
nor U13094 (N_13094,N_9743,N_9825);
nand U13095 (N_13095,N_7733,N_7553);
xnor U13096 (N_13096,N_7358,N_5534);
nand U13097 (N_13097,N_7410,N_8429);
xnor U13098 (N_13098,N_5497,N_7601);
and U13099 (N_13099,N_8982,N_5418);
nor U13100 (N_13100,N_6454,N_7195);
nor U13101 (N_13101,N_6414,N_5747);
nand U13102 (N_13102,N_9957,N_8947);
and U13103 (N_13103,N_8827,N_7216);
nand U13104 (N_13104,N_5408,N_5727);
xor U13105 (N_13105,N_6829,N_9735);
or U13106 (N_13106,N_9882,N_7419);
and U13107 (N_13107,N_9148,N_8721);
nor U13108 (N_13108,N_8010,N_7476);
and U13109 (N_13109,N_5311,N_7811);
or U13110 (N_13110,N_9813,N_9109);
nor U13111 (N_13111,N_9109,N_9825);
and U13112 (N_13112,N_7782,N_8178);
nand U13113 (N_13113,N_9752,N_7701);
nand U13114 (N_13114,N_7332,N_8399);
and U13115 (N_13115,N_9293,N_5877);
nor U13116 (N_13116,N_5289,N_7671);
nor U13117 (N_13117,N_6479,N_8745);
or U13118 (N_13118,N_5576,N_9787);
or U13119 (N_13119,N_5647,N_9399);
or U13120 (N_13120,N_8897,N_7306);
and U13121 (N_13121,N_6539,N_7285);
or U13122 (N_13122,N_5347,N_8939);
or U13123 (N_13123,N_6897,N_9149);
and U13124 (N_13124,N_9339,N_5952);
xnor U13125 (N_13125,N_9797,N_7077);
or U13126 (N_13126,N_7545,N_9780);
or U13127 (N_13127,N_9352,N_7797);
nor U13128 (N_13128,N_8961,N_5391);
nand U13129 (N_13129,N_5911,N_7734);
and U13130 (N_13130,N_5526,N_6416);
xor U13131 (N_13131,N_6413,N_6505);
nand U13132 (N_13132,N_7362,N_8602);
nand U13133 (N_13133,N_5002,N_5423);
and U13134 (N_13134,N_9442,N_6863);
xor U13135 (N_13135,N_7161,N_8883);
nor U13136 (N_13136,N_5807,N_9010);
and U13137 (N_13137,N_7183,N_8582);
nand U13138 (N_13138,N_8581,N_9545);
nor U13139 (N_13139,N_7473,N_8665);
nand U13140 (N_13140,N_5245,N_8492);
nor U13141 (N_13141,N_6846,N_5890);
and U13142 (N_13142,N_9295,N_9293);
nor U13143 (N_13143,N_5372,N_7222);
nor U13144 (N_13144,N_9888,N_7120);
nor U13145 (N_13145,N_6753,N_5349);
nor U13146 (N_13146,N_6101,N_6622);
or U13147 (N_13147,N_6360,N_8194);
and U13148 (N_13148,N_9263,N_6971);
xnor U13149 (N_13149,N_8247,N_5179);
or U13150 (N_13150,N_7907,N_6666);
nor U13151 (N_13151,N_7893,N_6482);
nor U13152 (N_13152,N_9779,N_7545);
or U13153 (N_13153,N_6103,N_7706);
or U13154 (N_13154,N_5910,N_5159);
or U13155 (N_13155,N_8652,N_6711);
and U13156 (N_13156,N_7382,N_8671);
nand U13157 (N_13157,N_6179,N_8030);
nor U13158 (N_13158,N_6829,N_7943);
nand U13159 (N_13159,N_9155,N_6440);
or U13160 (N_13160,N_5983,N_7976);
or U13161 (N_13161,N_9954,N_5200);
or U13162 (N_13162,N_9731,N_7922);
nor U13163 (N_13163,N_5746,N_8485);
nand U13164 (N_13164,N_9738,N_6342);
xor U13165 (N_13165,N_9084,N_7913);
or U13166 (N_13166,N_9980,N_6540);
or U13167 (N_13167,N_5347,N_6422);
or U13168 (N_13168,N_7638,N_9125);
or U13169 (N_13169,N_5478,N_9681);
or U13170 (N_13170,N_6425,N_5340);
and U13171 (N_13171,N_5877,N_5448);
or U13172 (N_13172,N_9567,N_5387);
and U13173 (N_13173,N_7653,N_6304);
nand U13174 (N_13174,N_9842,N_8986);
or U13175 (N_13175,N_5161,N_8129);
nand U13176 (N_13176,N_6154,N_5765);
xor U13177 (N_13177,N_7686,N_5570);
and U13178 (N_13178,N_6722,N_7517);
xnor U13179 (N_13179,N_5432,N_8082);
nand U13180 (N_13180,N_5114,N_6963);
nor U13181 (N_13181,N_9868,N_9291);
nor U13182 (N_13182,N_8054,N_9763);
nor U13183 (N_13183,N_9848,N_8024);
or U13184 (N_13184,N_7674,N_6047);
or U13185 (N_13185,N_6049,N_7750);
or U13186 (N_13186,N_6141,N_6325);
xor U13187 (N_13187,N_7593,N_5110);
and U13188 (N_13188,N_9757,N_9912);
xnor U13189 (N_13189,N_6575,N_8550);
nor U13190 (N_13190,N_9898,N_9944);
xnor U13191 (N_13191,N_6405,N_7271);
nand U13192 (N_13192,N_7800,N_9386);
nand U13193 (N_13193,N_8592,N_5380);
nor U13194 (N_13194,N_5478,N_7853);
nand U13195 (N_13195,N_7750,N_9320);
nor U13196 (N_13196,N_8853,N_7364);
or U13197 (N_13197,N_6768,N_6763);
and U13198 (N_13198,N_8830,N_5207);
and U13199 (N_13199,N_5141,N_9965);
nor U13200 (N_13200,N_6731,N_7047);
nand U13201 (N_13201,N_6693,N_5754);
and U13202 (N_13202,N_7553,N_9763);
nand U13203 (N_13203,N_5035,N_5154);
nand U13204 (N_13204,N_5186,N_5734);
or U13205 (N_13205,N_7327,N_6921);
nor U13206 (N_13206,N_7914,N_6348);
and U13207 (N_13207,N_9444,N_9673);
or U13208 (N_13208,N_8501,N_9265);
or U13209 (N_13209,N_6513,N_8466);
and U13210 (N_13210,N_7776,N_7946);
xor U13211 (N_13211,N_7721,N_9043);
or U13212 (N_13212,N_6303,N_8053);
and U13213 (N_13213,N_9278,N_7723);
nor U13214 (N_13214,N_8667,N_8738);
or U13215 (N_13215,N_6131,N_9744);
nor U13216 (N_13216,N_6382,N_5656);
nand U13217 (N_13217,N_8252,N_9893);
or U13218 (N_13218,N_5921,N_6879);
or U13219 (N_13219,N_6871,N_6876);
xnor U13220 (N_13220,N_9177,N_8367);
nor U13221 (N_13221,N_5544,N_5852);
and U13222 (N_13222,N_6562,N_8904);
or U13223 (N_13223,N_7308,N_8889);
nor U13224 (N_13224,N_6152,N_5698);
or U13225 (N_13225,N_7934,N_6652);
nor U13226 (N_13226,N_7320,N_9980);
and U13227 (N_13227,N_9019,N_8249);
xor U13228 (N_13228,N_5262,N_8594);
or U13229 (N_13229,N_6830,N_7963);
and U13230 (N_13230,N_7544,N_5725);
nand U13231 (N_13231,N_7780,N_8928);
or U13232 (N_13232,N_6542,N_7529);
or U13233 (N_13233,N_6930,N_6641);
xor U13234 (N_13234,N_5603,N_8745);
or U13235 (N_13235,N_9765,N_8357);
xnor U13236 (N_13236,N_7373,N_5024);
nor U13237 (N_13237,N_7083,N_5232);
xor U13238 (N_13238,N_7061,N_7742);
or U13239 (N_13239,N_7344,N_7515);
and U13240 (N_13240,N_6215,N_6920);
and U13241 (N_13241,N_8482,N_5503);
and U13242 (N_13242,N_6291,N_5646);
nand U13243 (N_13243,N_9844,N_8084);
and U13244 (N_13244,N_9378,N_5869);
or U13245 (N_13245,N_8862,N_9145);
or U13246 (N_13246,N_6816,N_5674);
and U13247 (N_13247,N_7621,N_9006);
and U13248 (N_13248,N_5266,N_9844);
or U13249 (N_13249,N_6026,N_9138);
and U13250 (N_13250,N_7880,N_6814);
and U13251 (N_13251,N_5808,N_7191);
nand U13252 (N_13252,N_9950,N_9235);
nand U13253 (N_13253,N_6892,N_6427);
and U13254 (N_13254,N_7781,N_5937);
nand U13255 (N_13255,N_6174,N_6267);
nor U13256 (N_13256,N_9089,N_6444);
nor U13257 (N_13257,N_8578,N_9703);
nand U13258 (N_13258,N_7914,N_9649);
nor U13259 (N_13259,N_6592,N_7240);
nor U13260 (N_13260,N_7433,N_9782);
nor U13261 (N_13261,N_5509,N_8692);
and U13262 (N_13262,N_5829,N_7004);
and U13263 (N_13263,N_7025,N_7434);
and U13264 (N_13264,N_6965,N_8725);
nor U13265 (N_13265,N_6498,N_6137);
and U13266 (N_13266,N_6729,N_8510);
or U13267 (N_13267,N_9992,N_6622);
nand U13268 (N_13268,N_9173,N_7858);
nand U13269 (N_13269,N_9001,N_9451);
or U13270 (N_13270,N_5953,N_6633);
nand U13271 (N_13271,N_9169,N_7839);
xor U13272 (N_13272,N_7035,N_7450);
or U13273 (N_13273,N_5925,N_5268);
and U13274 (N_13274,N_9799,N_5399);
and U13275 (N_13275,N_7049,N_5383);
nand U13276 (N_13276,N_8589,N_7085);
nor U13277 (N_13277,N_5539,N_8513);
nor U13278 (N_13278,N_9940,N_5865);
and U13279 (N_13279,N_9502,N_9511);
and U13280 (N_13280,N_5958,N_8273);
xnor U13281 (N_13281,N_7770,N_5958);
and U13282 (N_13282,N_9920,N_9757);
nor U13283 (N_13283,N_9633,N_7981);
nand U13284 (N_13284,N_5042,N_6469);
nor U13285 (N_13285,N_5438,N_7715);
or U13286 (N_13286,N_8969,N_7661);
and U13287 (N_13287,N_8360,N_5145);
nand U13288 (N_13288,N_6073,N_6208);
xor U13289 (N_13289,N_9978,N_6817);
nand U13290 (N_13290,N_9189,N_7025);
xor U13291 (N_13291,N_9263,N_6949);
or U13292 (N_13292,N_6938,N_5433);
xnor U13293 (N_13293,N_9560,N_5263);
or U13294 (N_13294,N_9685,N_9226);
nand U13295 (N_13295,N_5727,N_6988);
and U13296 (N_13296,N_7996,N_5828);
and U13297 (N_13297,N_7182,N_5799);
nand U13298 (N_13298,N_7924,N_8597);
or U13299 (N_13299,N_7712,N_8340);
nand U13300 (N_13300,N_6209,N_9368);
or U13301 (N_13301,N_5335,N_6422);
nand U13302 (N_13302,N_8702,N_9512);
nand U13303 (N_13303,N_6226,N_6445);
or U13304 (N_13304,N_8637,N_6267);
nand U13305 (N_13305,N_9506,N_9513);
or U13306 (N_13306,N_6112,N_7165);
nand U13307 (N_13307,N_7364,N_6999);
or U13308 (N_13308,N_9334,N_5720);
xnor U13309 (N_13309,N_8464,N_6501);
and U13310 (N_13310,N_9782,N_7389);
or U13311 (N_13311,N_5992,N_8411);
and U13312 (N_13312,N_7927,N_7433);
nand U13313 (N_13313,N_8786,N_5282);
or U13314 (N_13314,N_7740,N_5928);
nor U13315 (N_13315,N_9046,N_7277);
xor U13316 (N_13316,N_7317,N_7328);
nor U13317 (N_13317,N_7864,N_6271);
or U13318 (N_13318,N_8881,N_9960);
nor U13319 (N_13319,N_7080,N_5505);
nor U13320 (N_13320,N_9874,N_5015);
and U13321 (N_13321,N_5735,N_5784);
and U13322 (N_13322,N_5408,N_7613);
and U13323 (N_13323,N_8361,N_6792);
nor U13324 (N_13324,N_7435,N_5262);
or U13325 (N_13325,N_8986,N_7372);
and U13326 (N_13326,N_8408,N_9495);
nor U13327 (N_13327,N_5929,N_5528);
and U13328 (N_13328,N_8383,N_8514);
and U13329 (N_13329,N_7561,N_7077);
nand U13330 (N_13330,N_6106,N_5052);
and U13331 (N_13331,N_8887,N_8815);
nand U13332 (N_13332,N_6351,N_7727);
xor U13333 (N_13333,N_6175,N_7967);
xnor U13334 (N_13334,N_6309,N_6236);
nand U13335 (N_13335,N_5211,N_6703);
or U13336 (N_13336,N_5616,N_5885);
or U13337 (N_13337,N_5213,N_6041);
and U13338 (N_13338,N_8767,N_6840);
nand U13339 (N_13339,N_5005,N_9553);
or U13340 (N_13340,N_9382,N_6027);
xnor U13341 (N_13341,N_6924,N_5473);
and U13342 (N_13342,N_6993,N_5662);
or U13343 (N_13343,N_8559,N_6173);
and U13344 (N_13344,N_5774,N_7896);
nor U13345 (N_13345,N_6607,N_6596);
nor U13346 (N_13346,N_8626,N_8826);
nor U13347 (N_13347,N_5876,N_7425);
and U13348 (N_13348,N_8526,N_9588);
or U13349 (N_13349,N_6765,N_7124);
nor U13350 (N_13350,N_9930,N_8083);
nand U13351 (N_13351,N_9077,N_6038);
and U13352 (N_13352,N_8663,N_9601);
nand U13353 (N_13353,N_8878,N_8349);
and U13354 (N_13354,N_8952,N_9444);
xor U13355 (N_13355,N_7258,N_5887);
or U13356 (N_13356,N_5816,N_8401);
and U13357 (N_13357,N_5131,N_8556);
nor U13358 (N_13358,N_5538,N_9698);
nand U13359 (N_13359,N_9171,N_7698);
or U13360 (N_13360,N_6444,N_7360);
and U13361 (N_13361,N_6742,N_8034);
or U13362 (N_13362,N_6358,N_9737);
nand U13363 (N_13363,N_7693,N_9837);
nand U13364 (N_13364,N_5282,N_7216);
and U13365 (N_13365,N_8847,N_5729);
nand U13366 (N_13366,N_6875,N_8459);
and U13367 (N_13367,N_9246,N_9642);
xor U13368 (N_13368,N_9816,N_6082);
nand U13369 (N_13369,N_9891,N_9698);
and U13370 (N_13370,N_8561,N_5551);
and U13371 (N_13371,N_5079,N_5999);
nor U13372 (N_13372,N_7835,N_6934);
and U13373 (N_13373,N_9969,N_5590);
or U13374 (N_13374,N_8982,N_8783);
nor U13375 (N_13375,N_7837,N_5254);
and U13376 (N_13376,N_6668,N_9828);
nor U13377 (N_13377,N_9146,N_8806);
or U13378 (N_13378,N_5608,N_8636);
or U13379 (N_13379,N_7116,N_8320);
or U13380 (N_13380,N_7829,N_5789);
or U13381 (N_13381,N_6267,N_6155);
nor U13382 (N_13382,N_5349,N_9497);
nand U13383 (N_13383,N_5757,N_9813);
or U13384 (N_13384,N_8779,N_9490);
or U13385 (N_13385,N_5498,N_9543);
nor U13386 (N_13386,N_6170,N_8182);
or U13387 (N_13387,N_5856,N_5631);
and U13388 (N_13388,N_6768,N_9559);
and U13389 (N_13389,N_9012,N_5955);
xor U13390 (N_13390,N_8458,N_6404);
or U13391 (N_13391,N_6337,N_5607);
nor U13392 (N_13392,N_8607,N_6416);
nand U13393 (N_13393,N_5231,N_6553);
and U13394 (N_13394,N_9249,N_5743);
or U13395 (N_13395,N_7612,N_6428);
and U13396 (N_13396,N_9690,N_5204);
or U13397 (N_13397,N_5978,N_7709);
or U13398 (N_13398,N_9669,N_7345);
xnor U13399 (N_13399,N_9845,N_8071);
and U13400 (N_13400,N_5748,N_9765);
nor U13401 (N_13401,N_8079,N_8929);
xnor U13402 (N_13402,N_6152,N_7784);
and U13403 (N_13403,N_5571,N_8192);
or U13404 (N_13404,N_7611,N_6348);
and U13405 (N_13405,N_7141,N_7763);
nand U13406 (N_13406,N_7353,N_5435);
nand U13407 (N_13407,N_7862,N_7024);
and U13408 (N_13408,N_9740,N_7165);
nand U13409 (N_13409,N_7529,N_8258);
and U13410 (N_13410,N_6534,N_5723);
and U13411 (N_13411,N_5445,N_7244);
xnor U13412 (N_13412,N_7185,N_6039);
nor U13413 (N_13413,N_6699,N_9476);
or U13414 (N_13414,N_6632,N_9065);
and U13415 (N_13415,N_5230,N_7265);
nand U13416 (N_13416,N_7437,N_5327);
nor U13417 (N_13417,N_8882,N_9834);
nand U13418 (N_13418,N_6278,N_6259);
or U13419 (N_13419,N_6740,N_6975);
nand U13420 (N_13420,N_5566,N_5970);
nor U13421 (N_13421,N_6976,N_9989);
and U13422 (N_13422,N_7217,N_5545);
and U13423 (N_13423,N_9869,N_9522);
and U13424 (N_13424,N_5266,N_7844);
nand U13425 (N_13425,N_9156,N_7582);
nand U13426 (N_13426,N_7383,N_8908);
and U13427 (N_13427,N_7795,N_5011);
or U13428 (N_13428,N_8064,N_5096);
nand U13429 (N_13429,N_6191,N_5337);
nor U13430 (N_13430,N_5940,N_6484);
and U13431 (N_13431,N_5996,N_7023);
nand U13432 (N_13432,N_9622,N_7717);
or U13433 (N_13433,N_7251,N_7512);
nor U13434 (N_13434,N_9955,N_7968);
nand U13435 (N_13435,N_7280,N_6646);
nand U13436 (N_13436,N_7915,N_6738);
and U13437 (N_13437,N_9129,N_7802);
or U13438 (N_13438,N_9489,N_5886);
nand U13439 (N_13439,N_6888,N_8293);
nor U13440 (N_13440,N_7474,N_5009);
nor U13441 (N_13441,N_9834,N_9936);
nor U13442 (N_13442,N_9238,N_5928);
nor U13443 (N_13443,N_7690,N_5152);
or U13444 (N_13444,N_5938,N_5363);
or U13445 (N_13445,N_7604,N_8324);
nor U13446 (N_13446,N_5474,N_9038);
and U13447 (N_13447,N_5068,N_5553);
nor U13448 (N_13448,N_7509,N_9166);
or U13449 (N_13449,N_5061,N_8443);
or U13450 (N_13450,N_7967,N_8006);
or U13451 (N_13451,N_8946,N_5420);
or U13452 (N_13452,N_5661,N_8111);
nor U13453 (N_13453,N_5576,N_7980);
nand U13454 (N_13454,N_6972,N_6234);
or U13455 (N_13455,N_8246,N_7026);
nor U13456 (N_13456,N_5230,N_5501);
nor U13457 (N_13457,N_6486,N_5511);
xnor U13458 (N_13458,N_8671,N_9382);
and U13459 (N_13459,N_9330,N_6336);
nand U13460 (N_13460,N_9735,N_7427);
nand U13461 (N_13461,N_6521,N_7613);
nor U13462 (N_13462,N_6887,N_8120);
nand U13463 (N_13463,N_7279,N_7268);
nand U13464 (N_13464,N_5129,N_9706);
xor U13465 (N_13465,N_8032,N_5063);
and U13466 (N_13466,N_9449,N_5111);
nor U13467 (N_13467,N_7160,N_7784);
nand U13468 (N_13468,N_9056,N_8667);
nand U13469 (N_13469,N_6951,N_5403);
xor U13470 (N_13470,N_6836,N_7572);
and U13471 (N_13471,N_9486,N_5917);
xnor U13472 (N_13472,N_9531,N_8292);
nor U13473 (N_13473,N_7194,N_5023);
or U13474 (N_13474,N_8329,N_8153);
and U13475 (N_13475,N_7332,N_8249);
and U13476 (N_13476,N_8130,N_5901);
nor U13477 (N_13477,N_7774,N_8062);
nor U13478 (N_13478,N_9102,N_6538);
nand U13479 (N_13479,N_6935,N_5269);
or U13480 (N_13480,N_8289,N_6622);
and U13481 (N_13481,N_5572,N_9521);
nand U13482 (N_13482,N_8634,N_5321);
nor U13483 (N_13483,N_6500,N_5536);
nor U13484 (N_13484,N_5773,N_9809);
nor U13485 (N_13485,N_5173,N_9602);
or U13486 (N_13486,N_5760,N_9073);
nand U13487 (N_13487,N_5784,N_7096);
and U13488 (N_13488,N_8119,N_7547);
nand U13489 (N_13489,N_8175,N_7625);
nor U13490 (N_13490,N_9991,N_5858);
or U13491 (N_13491,N_6574,N_9503);
or U13492 (N_13492,N_5346,N_6129);
or U13493 (N_13493,N_5498,N_8510);
nor U13494 (N_13494,N_5865,N_5665);
or U13495 (N_13495,N_7865,N_7290);
and U13496 (N_13496,N_7325,N_9796);
nand U13497 (N_13497,N_6774,N_6937);
or U13498 (N_13498,N_8807,N_6378);
and U13499 (N_13499,N_8706,N_6600);
and U13500 (N_13500,N_6477,N_6287);
nand U13501 (N_13501,N_7280,N_6825);
or U13502 (N_13502,N_8894,N_7079);
and U13503 (N_13503,N_8295,N_8982);
nor U13504 (N_13504,N_8658,N_6709);
nor U13505 (N_13505,N_8915,N_7639);
xor U13506 (N_13506,N_9239,N_7625);
and U13507 (N_13507,N_6617,N_9577);
or U13508 (N_13508,N_8547,N_5172);
and U13509 (N_13509,N_5331,N_5388);
nor U13510 (N_13510,N_6203,N_8647);
nand U13511 (N_13511,N_9900,N_9987);
nand U13512 (N_13512,N_8028,N_5740);
nand U13513 (N_13513,N_9569,N_6214);
and U13514 (N_13514,N_8826,N_9796);
nand U13515 (N_13515,N_5684,N_9708);
nor U13516 (N_13516,N_5583,N_8218);
and U13517 (N_13517,N_6331,N_5038);
and U13518 (N_13518,N_7966,N_6384);
nand U13519 (N_13519,N_7519,N_8197);
nand U13520 (N_13520,N_7212,N_6195);
xor U13521 (N_13521,N_5436,N_5801);
nor U13522 (N_13522,N_6401,N_8497);
xnor U13523 (N_13523,N_5953,N_9779);
nor U13524 (N_13524,N_5763,N_7868);
nand U13525 (N_13525,N_8535,N_5716);
or U13526 (N_13526,N_5349,N_5711);
nand U13527 (N_13527,N_5346,N_6094);
xor U13528 (N_13528,N_8693,N_8226);
and U13529 (N_13529,N_7218,N_9808);
or U13530 (N_13530,N_5026,N_6028);
nand U13531 (N_13531,N_6118,N_8896);
nand U13532 (N_13532,N_5213,N_7680);
or U13533 (N_13533,N_5985,N_9671);
nand U13534 (N_13534,N_9985,N_7849);
nor U13535 (N_13535,N_8828,N_9518);
or U13536 (N_13536,N_8156,N_7808);
nor U13537 (N_13537,N_5848,N_6759);
and U13538 (N_13538,N_7385,N_8898);
xnor U13539 (N_13539,N_6542,N_9465);
nor U13540 (N_13540,N_5108,N_5775);
nand U13541 (N_13541,N_5460,N_6271);
nor U13542 (N_13542,N_6340,N_7925);
nor U13543 (N_13543,N_7014,N_9535);
and U13544 (N_13544,N_5853,N_9576);
and U13545 (N_13545,N_8987,N_5483);
or U13546 (N_13546,N_6176,N_7508);
or U13547 (N_13547,N_5169,N_8716);
nor U13548 (N_13548,N_5286,N_8599);
nor U13549 (N_13549,N_8784,N_5169);
nor U13550 (N_13550,N_7046,N_9231);
nand U13551 (N_13551,N_7067,N_7900);
or U13552 (N_13552,N_6530,N_9721);
nor U13553 (N_13553,N_8703,N_5720);
or U13554 (N_13554,N_5914,N_5155);
xnor U13555 (N_13555,N_8004,N_5615);
nor U13556 (N_13556,N_6443,N_5147);
and U13557 (N_13557,N_5698,N_8576);
nor U13558 (N_13558,N_5673,N_6196);
and U13559 (N_13559,N_8746,N_5291);
nand U13560 (N_13560,N_5027,N_6399);
and U13561 (N_13561,N_5645,N_5896);
and U13562 (N_13562,N_5023,N_8766);
nor U13563 (N_13563,N_9444,N_7379);
and U13564 (N_13564,N_6187,N_8495);
or U13565 (N_13565,N_5467,N_8605);
nand U13566 (N_13566,N_6551,N_8494);
or U13567 (N_13567,N_8395,N_8938);
nand U13568 (N_13568,N_9679,N_9519);
nor U13569 (N_13569,N_8280,N_7018);
and U13570 (N_13570,N_5736,N_5192);
and U13571 (N_13571,N_6166,N_7671);
or U13572 (N_13572,N_9896,N_6830);
xor U13573 (N_13573,N_8417,N_7891);
nor U13574 (N_13574,N_6840,N_9377);
or U13575 (N_13575,N_7600,N_6040);
xor U13576 (N_13576,N_9552,N_9499);
nor U13577 (N_13577,N_6943,N_7624);
or U13578 (N_13578,N_9230,N_9830);
nand U13579 (N_13579,N_7760,N_9067);
nor U13580 (N_13580,N_7603,N_5361);
or U13581 (N_13581,N_9917,N_6909);
nor U13582 (N_13582,N_7781,N_7205);
xor U13583 (N_13583,N_5607,N_8470);
xor U13584 (N_13584,N_6714,N_5553);
nand U13585 (N_13585,N_9284,N_8487);
or U13586 (N_13586,N_9708,N_7775);
nand U13587 (N_13587,N_8844,N_5166);
xor U13588 (N_13588,N_6358,N_5908);
nor U13589 (N_13589,N_7176,N_7535);
nor U13590 (N_13590,N_7881,N_7372);
or U13591 (N_13591,N_8737,N_9288);
nand U13592 (N_13592,N_6645,N_7751);
nand U13593 (N_13593,N_6041,N_7611);
nand U13594 (N_13594,N_8575,N_8294);
nor U13595 (N_13595,N_9892,N_8002);
or U13596 (N_13596,N_5237,N_5012);
and U13597 (N_13597,N_6973,N_8239);
or U13598 (N_13598,N_6702,N_7424);
or U13599 (N_13599,N_9292,N_6964);
nor U13600 (N_13600,N_8695,N_5747);
nand U13601 (N_13601,N_7834,N_8892);
or U13602 (N_13602,N_7490,N_6719);
nand U13603 (N_13603,N_5547,N_7673);
or U13604 (N_13604,N_7403,N_6858);
and U13605 (N_13605,N_7434,N_9230);
nand U13606 (N_13606,N_8083,N_7751);
and U13607 (N_13607,N_6800,N_5645);
nand U13608 (N_13608,N_5098,N_7399);
and U13609 (N_13609,N_5734,N_8079);
and U13610 (N_13610,N_6098,N_5231);
or U13611 (N_13611,N_6270,N_6898);
or U13612 (N_13612,N_6629,N_5302);
nor U13613 (N_13613,N_9532,N_6299);
nand U13614 (N_13614,N_8425,N_8796);
or U13615 (N_13615,N_5521,N_8924);
or U13616 (N_13616,N_5488,N_8116);
or U13617 (N_13617,N_9238,N_8465);
and U13618 (N_13618,N_7778,N_8185);
nand U13619 (N_13619,N_9976,N_6037);
nor U13620 (N_13620,N_8819,N_8755);
nor U13621 (N_13621,N_6556,N_9122);
nor U13622 (N_13622,N_9706,N_9323);
and U13623 (N_13623,N_9377,N_8750);
nand U13624 (N_13624,N_9684,N_8786);
or U13625 (N_13625,N_5536,N_7476);
nor U13626 (N_13626,N_8916,N_6005);
nand U13627 (N_13627,N_5319,N_7444);
nand U13628 (N_13628,N_9321,N_7421);
or U13629 (N_13629,N_8187,N_9489);
or U13630 (N_13630,N_7085,N_6298);
xor U13631 (N_13631,N_7259,N_8013);
and U13632 (N_13632,N_7642,N_5345);
and U13633 (N_13633,N_8075,N_9729);
or U13634 (N_13634,N_8422,N_9633);
nor U13635 (N_13635,N_8925,N_5128);
nor U13636 (N_13636,N_8168,N_9331);
or U13637 (N_13637,N_6486,N_6612);
nor U13638 (N_13638,N_8050,N_7386);
or U13639 (N_13639,N_8119,N_7606);
nor U13640 (N_13640,N_6781,N_5675);
xnor U13641 (N_13641,N_9390,N_8780);
nor U13642 (N_13642,N_6159,N_7449);
or U13643 (N_13643,N_8014,N_8573);
or U13644 (N_13644,N_7304,N_6921);
nor U13645 (N_13645,N_9510,N_6430);
nor U13646 (N_13646,N_9445,N_5544);
and U13647 (N_13647,N_6394,N_5553);
nor U13648 (N_13648,N_6633,N_6362);
and U13649 (N_13649,N_8964,N_8808);
and U13650 (N_13650,N_6501,N_9663);
nor U13651 (N_13651,N_7194,N_9421);
xor U13652 (N_13652,N_5435,N_8091);
and U13653 (N_13653,N_8187,N_9739);
or U13654 (N_13654,N_9535,N_9493);
or U13655 (N_13655,N_8681,N_5741);
nor U13656 (N_13656,N_6104,N_6115);
and U13657 (N_13657,N_7096,N_7072);
xor U13658 (N_13658,N_9086,N_9495);
nor U13659 (N_13659,N_5575,N_8580);
nor U13660 (N_13660,N_6122,N_6135);
nor U13661 (N_13661,N_9555,N_6149);
nor U13662 (N_13662,N_5557,N_9751);
nand U13663 (N_13663,N_9080,N_8179);
nor U13664 (N_13664,N_5740,N_9271);
nor U13665 (N_13665,N_5973,N_8150);
nand U13666 (N_13666,N_8078,N_6744);
and U13667 (N_13667,N_5205,N_6812);
or U13668 (N_13668,N_9958,N_9184);
nor U13669 (N_13669,N_8359,N_8222);
or U13670 (N_13670,N_9459,N_5206);
xor U13671 (N_13671,N_6584,N_6610);
and U13672 (N_13672,N_7689,N_9586);
nand U13673 (N_13673,N_7764,N_9463);
nor U13674 (N_13674,N_5562,N_6587);
and U13675 (N_13675,N_9160,N_7858);
nor U13676 (N_13676,N_9500,N_7297);
or U13677 (N_13677,N_6019,N_7864);
nor U13678 (N_13678,N_6209,N_5151);
or U13679 (N_13679,N_6263,N_9296);
or U13680 (N_13680,N_5731,N_5554);
or U13681 (N_13681,N_7110,N_7666);
and U13682 (N_13682,N_8794,N_7005);
nand U13683 (N_13683,N_6430,N_5736);
or U13684 (N_13684,N_7829,N_8303);
and U13685 (N_13685,N_9660,N_6632);
nand U13686 (N_13686,N_9778,N_6265);
and U13687 (N_13687,N_8582,N_8758);
xnor U13688 (N_13688,N_7791,N_9709);
or U13689 (N_13689,N_9593,N_9109);
nor U13690 (N_13690,N_8813,N_5966);
nand U13691 (N_13691,N_5428,N_9072);
nor U13692 (N_13692,N_9564,N_5647);
xor U13693 (N_13693,N_7646,N_6878);
or U13694 (N_13694,N_5711,N_5202);
or U13695 (N_13695,N_6957,N_6583);
nand U13696 (N_13696,N_5973,N_6933);
nor U13697 (N_13697,N_7633,N_9248);
xnor U13698 (N_13698,N_7090,N_9784);
or U13699 (N_13699,N_5526,N_8821);
nor U13700 (N_13700,N_7785,N_5114);
and U13701 (N_13701,N_7253,N_7180);
nand U13702 (N_13702,N_5844,N_5572);
nand U13703 (N_13703,N_7719,N_7981);
nand U13704 (N_13704,N_8442,N_5738);
and U13705 (N_13705,N_6329,N_9879);
or U13706 (N_13706,N_7423,N_9125);
nor U13707 (N_13707,N_7166,N_7272);
nor U13708 (N_13708,N_8303,N_5885);
xor U13709 (N_13709,N_6380,N_9114);
or U13710 (N_13710,N_5710,N_5397);
nor U13711 (N_13711,N_5416,N_5167);
and U13712 (N_13712,N_5999,N_5242);
or U13713 (N_13713,N_9316,N_5028);
and U13714 (N_13714,N_8569,N_6563);
xnor U13715 (N_13715,N_7346,N_8905);
and U13716 (N_13716,N_6666,N_9382);
xnor U13717 (N_13717,N_9354,N_5896);
nand U13718 (N_13718,N_6428,N_9026);
or U13719 (N_13719,N_9186,N_8880);
xnor U13720 (N_13720,N_9309,N_5087);
or U13721 (N_13721,N_6686,N_8457);
nand U13722 (N_13722,N_8640,N_7504);
or U13723 (N_13723,N_7334,N_9520);
and U13724 (N_13724,N_9154,N_8951);
or U13725 (N_13725,N_5922,N_8640);
nor U13726 (N_13726,N_9196,N_9156);
nor U13727 (N_13727,N_5075,N_8516);
nor U13728 (N_13728,N_7230,N_6571);
or U13729 (N_13729,N_7634,N_7952);
or U13730 (N_13730,N_6403,N_9426);
and U13731 (N_13731,N_6123,N_6310);
or U13732 (N_13732,N_5393,N_7734);
nor U13733 (N_13733,N_7123,N_5231);
nand U13734 (N_13734,N_9955,N_5363);
and U13735 (N_13735,N_5657,N_8591);
nand U13736 (N_13736,N_6565,N_7198);
nand U13737 (N_13737,N_9747,N_9091);
and U13738 (N_13738,N_6189,N_7669);
nand U13739 (N_13739,N_9856,N_9835);
xor U13740 (N_13740,N_5589,N_9225);
nand U13741 (N_13741,N_9033,N_7434);
nand U13742 (N_13742,N_5017,N_9104);
nand U13743 (N_13743,N_8552,N_7942);
or U13744 (N_13744,N_9979,N_6464);
or U13745 (N_13745,N_7277,N_7267);
nor U13746 (N_13746,N_7895,N_9849);
or U13747 (N_13747,N_7852,N_7060);
nor U13748 (N_13748,N_7241,N_6039);
or U13749 (N_13749,N_8517,N_5125);
and U13750 (N_13750,N_7685,N_7530);
or U13751 (N_13751,N_9527,N_8112);
nor U13752 (N_13752,N_8209,N_8583);
or U13753 (N_13753,N_8917,N_5349);
nand U13754 (N_13754,N_5039,N_9693);
and U13755 (N_13755,N_8663,N_7149);
or U13756 (N_13756,N_6984,N_6638);
and U13757 (N_13757,N_8096,N_9524);
or U13758 (N_13758,N_8294,N_8697);
and U13759 (N_13759,N_9911,N_9073);
or U13760 (N_13760,N_6696,N_8492);
nor U13761 (N_13761,N_6894,N_9452);
and U13762 (N_13762,N_7674,N_7704);
or U13763 (N_13763,N_9089,N_8169);
or U13764 (N_13764,N_8916,N_6381);
or U13765 (N_13765,N_7588,N_5273);
or U13766 (N_13766,N_8245,N_8724);
nand U13767 (N_13767,N_9255,N_5349);
xnor U13768 (N_13768,N_7357,N_6508);
and U13769 (N_13769,N_6606,N_9898);
xnor U13770 (N_13770,N_5451,N_6759);
and U13771 (N_13771,N_9337,N_8547);
nand U13772 (N_13772,N_7361,N_9788);
or U13773 (N_13773,N_7766,N_7114);
or U13774 (N_13774,N_8873,N_8781);
or U13775 (N_13775,N_5835,N_8035);
nand U13776 (N_13776,N_7968,N_9712);
and U13777 (N_13777,N_5492,N_7555);
nand U13778 (N_13778,N_6926,N_6379);
nor U13779 (N_13779,N_8657,N_7605);
and U13780 (N_13780,N_6386,N_9657);
and U13781 (N_13781,N_6351,N_6484);
nand U13782 (N_13782,N_5257,N_8624);
and U13783 (N_13783,N_6816,N_6648);
and U13784 (N_13784,N_8101,N_7969);
and U13785 (N_13785,N_8880,N_6866);
nand U13786 (N_13786,N_9951,N_7674);
nor U13787 (N_13787,N_7705,N_7872);
or U13788 (N_13788,N_6993,N_6624);
nand U13789 (N_13789,N_8072,N_6224);
nor U13790 (N_13790,N_5523,N_8143);
or U13791 (N_13791,N_5652,N_8387);
nand U13792 (N_13792,N_8496,N_6317);
or U13793 (N_13793,N_6268,N_9475);
and U13794 (N_13794,N_9728,N_9753);
nor U13795 (N_13795,N_5823,N_6376);
or U13796 (N_13796,N_5580,N_5728);
xnor U13797 (N_13797,N_7232,N_8462);
or U13798 (N_13798,N_7292,N_7256);
nor U13799 (N_13799,N_5646,N_5771);
or U13800 (N_13800,N_5095,N_8544);
or U13801 (N_13801,N_5585,N_6997);
or U13802 (N_13802,N_6361,N_8504);
and U13803 (N_13803,N_8160,N_8041);
or U13804 (N_13804,N_7531,N_5581);
or U13805 (N_13805,N_6145,N_5930);
and U13806 (N_13806,N_9849,N_5591);
nor U13807 (N_13807,N_8362,N_7967);
nand U13808 (N_13808,N_8827,N_8950);
xnor U13809 (N_13809,N_9690,N_6472);
nor U13810 (N_13810,N_9952,N_5942);
or U13811 (N_13811,N_7013,N_5229);
and U13812 (N_13812,N_6942,N_6190);
nand U13813 (N_13813,N_6498,N_9859);
nand U13814 (N_13814,N_6008,N_6952);
nand U13815 (N_13815,N_7175,N_7200);
and U13816 (N_13816,N_7093,N_9777);
nand U13817 (N_13817,N_9234,N_6572);
or U13818 (N_13818,N_8894,N_6541);
or U13819 (N_13819,N_7191,N_7642);
or U13820 (N_13820,N_8945,N_9991);
or U13821 (N_13821,N_7353,N_9994);
nor U13822 (N_13822,N_9851,N_9075);
or U13823 (N_13823,N_8863,N_6647);
or U13824 (N_13824,N_6139,N_6833);
nor U13825 (N_13825,N_9905,N_6936);
and U13826 (N_13826,N_9994,N_9003);
nand U13827 (N_13827,N_8647,N_5725);
xnor U13828 (N_13828,N_9787,N_7725);
or U13829 (N_13829,N_8701,N_6965);
nor U13830 (N_13830,N_9054,N_9210);
and U13831 (N_13831,N_8879,N_5185);
nand U13832 (N_13832,N_6749,N_8170);
or U13833 (N_13833,N_9056,N_6170);
nand U13834 (N_13834,N_8362,N_7630);
xor U13835 (N_13835,N_9459,N_9117);
nor U13836 (N_13836,N_9489,N_9144);
and U13837 (N_13837,N_6747,N_6361);
nor U13838 (N_13838,N_8599,N_9322);
nand U13839 (N_13839,N_7886,N_8870);
nor U13840 (N_13840,N_6804,N_5698);
nand U13841 (N_13841,N_5894,N_7432);
and U13842 (N_13842,N_8677,N_5186);
nand U13843 (N_13843,N_5053,N_9507);
nor U13844 (N_13844,N_6490,N_7751);
or U13845 (N_13845,N_7901,N_6517);
and U13846 (N_13846,N_7523,N_8947);
and U13847 (N_13847,N_7933,N_7568);
xor U13848 (N_13848,N_9888,N_8093);
nand U13849 (N_13849,N_6922,N_5499);
and U13850 (N_13850,N_7863,N_7856);
and U13851 (N_13851,N_9564,N_9218);
and U13852 (N_13852,N_7821,N_6190);
and U13853 (N_13853,N_5855,N_8045);
nand U13854 (N_13854,N_5071,N_9786);
or U13855 (N_13855,N_6434,N_5978);
nand U13856 (N_13856,N_5904,N_5797);
nand U13857 (N_13857,N_5086,N_8181);
or U13858 (N_13858,N_8324,N_6245);
xnor U13859 (N_13859,N_9382,N_9110);
xnor U13860 (N_13860,N_5650,N_7680);
nor U13861 (N_13861,N_5079,N_9118);
and U13862 (N_13862,N_7795,N_9266);
and U13863 (N_13863,N_7362,N_9214);
or U13864 (N_13864,N_5984,N_5199);
nand U13865 (N_13865,N_9875,N_8910);
or U13866 (N_13866,N_7919,N_5330);
nor U13867 (N_13867,N_6265,N_5950);
nand U13868 (N_13868,N_9569,N_5562);
nand U13869 (N_13869,N_6955,N_5337);
or U13870 (N_13870,N_9339,N_8638);
or U13871 (N_13871,N_6410,N_5822);
and U13872 (N_13872,N_8476,N_9794);
xnor U13873 (N_13873,N_5602,N_7882);
xor U13874 (N_13874,N_6837,N_7086);
or U13875 (N_13875,N_8631,N_8364);
or U13876 (N_13876,N_6252,N_5547);
nor U13877 (N_13877,N_5048,N_9246);
nand U13878 (N_13878,N_9832,N_5444);
xnor U13879 (N_13879,N_6809,N_9585);
nand U13880 (N_13880,N_7885,N_7842);
xor U13881 (N_13881,N_8618,N_9413);
or U13882 (N_13882,N_5604,N_8514);
or U13883 (N_13883,N_9720,N_6988);
and U13884 (N_13884,N_6788,N_9067);
and U13885 (N_13885,N_6566,N_7972);
and U13886 (N_13886,N_6349,N_6102);
or U13887 (N_13887,N_8741,N_5093);
or U13888 (N_13888,N_7339,N_6756);
nand U13889 (N_13889,N_9494,N_6652);
and U13890 (N_13890,N_5990,N_7520);
or U13891 (N_13891,N_6467,N_7579);
and U13892 (N_13892,N_7491,N_9534);
nand U13893 (N_13893,N_8131,N_8064);
nor U13894 (N_13894,N_5810,N_9489);
or U13895 (N_13895,N_7291,N_5570);
xnor U13896 (N_13896,N_8516,N_9182);
nand U13897 (N_13897,N_6497,N_8314);
xnor U13898 (N_13898,N_5262,N_9762);
xor U13899 (N_13899,N_7274,N_6214);
or U13900 (N_13900,N_5733,N_8098);
or U13901 (N_13901,N_7428,N_6345);
nor U13902 (N_13902,N_5828,N_5689);
nor U13903 (N_13903,N_8864,N_9462);
nor U13904 (N_13904,N_6663,N_5690);
nor U13905 (N_13905,N_7129,N_6341);
or U13906 (N_13906,N_9824,N_8942);
and U13907 (N_13907,N_7054,N_9360);
nand U13908 (N_13908,N_8545,N_5942);
or U13909 (N_13909,N_6704,N_5017);
or U13910 (N_13910,N_7732,N_9079);
nor U13911 (N_13911,N_7885,N_6466);
xor U13912 (N_13912,N_7877,N_6947);
nand U13913 (N_13913,N_5381,N_5664);
nor U13914 (N_13914,N_5116,N_8532);
and U13915 (N_13915,N_9362,N_9574);
nand U13916 (N_13916,N_9768,N_6241);
nor U13917 (N_13917,N_7336,N_9433);
nor U13918 (N_13918,N_9161,N_5781);
and U13919 (N_13919,N_6360,N_7553);
or U13920 (N_13920,N_5380,N_7438);
nand U13921 (N_13921,N_7474,N_9349);
nand U13922 (N_13922,N_6523,N_6982);
and U13923 (N_13923,N_7319,N_6801);
and U13924 (N_13924,N_5059,N_5831);
or U13925 (N_13925,N_6368,N_5376);
and U13926 (N_13926,N_7947,N_9635);
nor U13927 (N_13927,N_7141,N_5972);
xor U13928 (N_13928,N_7493,N_8731);
and U13929 (N_13929,N_9338,N_9940);
nand U13930 (N_13930,N_8542,N_6306);
nor U13931 (N_13931,N_7638,N_8462);
nand U13932 (N_13932,N_9086,N_5102);
or U13933 (N_13933,N_9457,N_5142);
nor U13934 (N_13934,N_6574,N_7613);
xnor U13935 (N_13935,N_8590,N_5706);
nand U13936 (N_13936,N_7577,N_7325);
or U13937 (N_13937,N_9860,N_5912);
nor U13938 (N_13938,N_6671,N_5402);
or U13939 (N_13939,N_5613,N_5711);
nor U13940 (N_13940,N_7088,N_9706);
nand U13941 (N_13941,N_8566,N_5759);
and U13942 (N_13942,N_6251,N_5490);
xnor U13943 (N_13943,N_6431,N_6849);
or U13944 (N_13944,N_6585,N_6324);
and U13945 (N_13945,N_6024,N_5505);
xnor U13946 (N_13946,N_7309,N_9012);
or U13947 (N_13947,N_6545,N_5895);
xnor U13948 (N_13948,N_7342,N_7078);
nor U13949 (N_13949,N_9946,N_6571);
nand U13950 (N_13950,N_6086,N_6052);
nor U13951 (N_13951,N_7402,N_8893);
xor U13952 (N_13952,N_5150,N_8781);
nand U13953 (N_13953,N_9015,N_8070);
or U13954 (N_13954,N_6589,N_6325);
and U13955 (N_13955,N_9352,N_9807);
and U13956 (N_13956,N_7951,N_7664);
or U13957 (N_13957,N_8848,N_8653);
nor U13958 (N_13958,N_6944,N_5632);
or U13959 (N_13959,N_8653,N_6380);
xor U13960 (N_13960,N_8325,N_8868);
nor U13961 (N_13961,N_6266,N_9266);
and U13962 (N_13962,N_8536,N_6756);
and U13963 (N_13963,N_7952,N_8173);
nand U13964 (N_13964,N_8112,N_6947);
and U13965 (N_13965,N_8579,N_8410);
and U13966 (N_13966,N_6095,N_6171);
nor U13967 (N_13967,N_6206,N_9678);
xor U13968 (N_13968,N_6138,N_9622);
and U13969 (N_13969,N_5863,N_8034);
nand U13970 (N_13970,N_7070,N_5098);
and U13971 (N_13971,N_9203,N_8105);
nand U13972 (N_13972,N_8455,N_7931);
or U13973 (N_13973,N_9931,N_5578);
nor U13974 (N_13974,N_8032,N_6124);
xnor U13975 (N_13975,N_9247,N_5989);
nor U13976 (N_13976,N_8109,N_9472);
or U13977 (N_13977,N_5884,N_6845);
or U13978 (N_13978,N_8836,N_7099);
nand U13979 (N_13979,N_8255,N_8351);
xnor U13980 (N_13980,N_7441,N_7373);
nor U13981 (N_13981,N_9486,N_6186);
xor U13982 (N_13982,N_8621,N_9601);
nand U13983 (N_13983,N_5127,N_7115);
or U13984 (N_13984,N_7150,N_8870);
nand U13985 (N_13985,N_8970,N_9549);
nand U13986 (N_13986,N_9078,N_6074);
xnor U13987 (N_13987,N_8893,N_9575);
or U13988 (N_13988,N_6623,N_8534);
and U13989 (N_13989,N_8938,N_6338);
xnor U13990 (N_13990,N_7480,N_7095);
nand U13991 (N_13991,N_5213,N_9573);
or U13992 (N_13992,N_5638,N_5512);
nor U13993 (N_13993,N_5129,N_5060);
and U13994 (N_13994,N_8427,N_7890);
nor U13995 (N_13995,N_7568,N_8264);
xor U13996 (N_13996,N_5023,N_5568);
nor U13997 (N_13997,N_9950,N_9853);
nor U13998 (N_13998,N_9980,N_7011);
or U13999 (N_13999,N_6049,N_8687);
and U14000 (N_14000,N_6604,N_7646);
nand U14001 (N_14001,N_7879,N_6757);
nand U14002 (N_14002,N_6043,N_8718);
nor U14003 (N_14003,N_6751,N_8351);
nand U14004 (N_14004,N_8645,N_8539);
nor U14005 (N_14005,N_5821,N_6363);
xnor U14006 (N_14006,N_9696,N_7295);
or U14007 (N_14007,N_6363,N_6377);
nor U14008 (N_14008,N_7307,N_7134);
nand U14009 (N_14009,N_7725,N_8347);
or U14010 (N_14010,N_9743,N_6477);
nand U14011 (N_14011,N_8924,N_5468);
and U14012 (N_14012,N_6196,N_6895);
nor U14013 (N_14013,N_8395,N_7612);
and U14014 (N_14014,N_8458,N_9075);
xnor U14015 (N_14015,N_7761,N_9228);
nor U14016 (N_14016,N_6642,N_8204);
nor U14017 (N_14017,N_7455,N_8030);
xnor U14018 (N_14018,N_5186,N_6963);
and U14019 (N_14019,N_9637,N_7481);
or U14020 (N_14020,N_6090,N_7975);
or U14021 (N_14021,N_6231,N_7533);
or U14022 (N_14022,N_6595,N_5782);
or U14023 (N_14023,N_7237,N_8918);
and U14024 (N_14024,N_7040,N_9391);
or U14025 (N_14025,N_9635,N_6217);
nor U14026 (N_14026,N_9055,N_9636);
or U14027 (N_14027,N_7412,N_8064);
or U14028 (N_14028,N_9831,N_8174);
and U14029 (N_14029,N_6601,N_5868);
nor U14030 (N_14030,N_9194,N_9094);
or U14031 (N_14031,N_7354,N_9738);
nand U14032 (N_14032,N_6572,N_5568);
nor U14033 (N_14033,N_7423,N_8797);
and U14034 (N_14034,N_8696,N_6435);
xor U14035 (N_14035,N_6186,N_5596);
and U14036 (N_14036,N_5787,N_5801);
xor U14037 (N_14037,N_5242,N_8944);
or U14038 (N_14038,N_7404,N_8859);
and U14039 (N_14039,N_9516,N_6400);
nor U14040 (N_14040,N_6162,N_6061);
or U14041 (N_14041,N_6144,N_5058);
xor U14042 (N_14042,N_8119,N_9037);
nor U14043 (N_14043,N_7239,N_6621);
xor U14044 (N_14044,N_6767,N_8918);
nor U14045 (N_14045,N_8147,N_5160);
or U14046 (N_14046,N_5296,N_8734);
or U14047 (N_14047,N_8337,N_9494);
nand U14048 (N_14048,N_9501,N_7572);
xor U14049 (N_14049,N_6257,N_5383);
or U14050 (N_14050,N_5436,N_5321);
or U14051 (N_14051,N_5739,N_9559);
and U14052 (N_14052,N_5171,N_9007);
nand U14053 (N_14053,N_5610,N_7714);
nor U14054 (N_14054,N_9934,N_7423);
nand U14055 (N_14055,N_8267,N_5053);
xor U14056 (N_14056,N_6960,N_5201);
nand U14057 (N_14057,N_6253,N_8895);
xnor U14058 (N_14058,N_9568,N_5830);
and U14059 (N_14059,N_6391,N_9742);
nor U14060 (N_14060,N_5963,N_7118);
xnor U14061 (N_14061,N_7325,N_9814);
or U14062 (N_14062,N_9902,N_9932);
or U14063 (N_14063,N_6083,N_9680);
nor U14064 (N_14064,N_7196,N_7639);
nand U14065 (N_14065,N_6490,N_8379);
xnor U14066 (N_14066,N_7753,N_7211);
and U14067 (N_14067,N_8209,N_9307);
nand U14068 (N_14068,N_5698,N_7561);
nand U14069 (N_14069,N_8808,N_9912);
nand U14070 (N_14070,N_7329,N_7083);
nor U14071 (N_14071,N_7264,N_8814);
or U14072 (N_14072,N_9069,N_6750);
nand U14073 (N_14073,N_6252,N_7438);
or U14074 (N_14074,N_8325,N_6101);
nor U14075 (N_14075,N_6515,N_6198);
xnor U14076 (N_14076,N_7773,N_9692);
xor U14077 (N_14077,N_8423,N_9381);
and U14078 (N_14078,N_6667,N_6258);
nor U14079 (N_14079,N_8904,N_5830);
nand U14080 (N_14080,N_7053,N_7884);
or U14081 (N_14081,N_8557,N_9211);
nor U14082 (N_14082,N_6991,N_9836);
and U14083 (N_14083,N_8363,N_6151);
xnor U14084 (N_14084,N_9676,N_5401);
nand U14085 (N_14085,N_8735,N_6272);
or U14086 (N_14086,N_9990,N_9922);
or U14087 (N_14087,N_6452,N_6093);
and U14088 (N_14088,N_7546,N_9802);
xnor U14089 (N_14089,N_8233,N_6620);
and U14090 (N_14090,N_8224,N_7642);
or U14091 (N_14091,N_5612,N_6323);
nor U14092 (N_14092,N_5007,N_5737);
and U14093 (N_14093,N_9001,N_9850);
nand U14094 (N_14094,N_6053,N_9118);
nor U14095 (N_14095,N_6854,N_8527);
nand U14096 (N_14096,N_6791,N_7096);
and U14097 (N_14097,N_5077,N_8333);
and U14098 (N_14098,N_5118,N_9191);
nor U14099 (N_14099,N_5431,N_7012);
and U14100 (N_14100,N_5003,N_9639);
or U14101 (N_14101,N_5700,N_5909);
nor U14102 (N_14102,N_9601,N_9989);
nand U14103 (N_14103,N_6719,N_5068);
and U14104 (N_14104,N_7373,N_5820);
nand U14105 (N_14105,N_7012,N_8390);
nor U14106 (N_14106,N_7358,N_8194);
nand U14107 (N_14107,N_8081,N_9609);
xor U14108 (N_14108,N_5433,N_5601);
nor U14109 (N_14109,N_6717,N_5408);
or U14110 (N_14110,N_7797,N_6266);
and U14111 (N_14111,N_8107,N_5792);
and U14112 (N_14112,N_8969,N_8301);
or U14113 (N_14113,N_8523,N_8021);
nor U14114 (N_14114,N_8712,N_7026);
or U14115 (N_14115,N_9291,N_8925);
and U14116 (N_14116,N_9361,N_8889);
nand U14117 (N_14117,N_9223,N_6107);
or U14118 (N_14118,N_8505,N_8085);
nand U14119 (N_14119,N_8933,N_8551);
nor U14120 (N_14120,N_7244,N_7718);
nor U14121 (N_14121,N_8644,N_7624);
or U14122 (N_14122,N_5258,N_6939);
nand U14123 (N_14123,N_6039,N_8327);
and U14124 (N_14124,N_9279,N_5357);
or U14125 (N_14125,N_8124,N_5651);
nor U14126 (N_14126,N_6799,N_9408);
nand U14127 (N_14127,N_6930,N_5862);
and U14128 (N_14128,N_7540,N_7236);
or U14129 (N_14129,N_6397,N_7790);
nor U14130 (N_14130,N_7665,N_8146);
and U14131 (N_14131,N_8859,N_6039);
xnor U14132 (N_14132,N_5756,N_7902);
and U14133 (N_14133,N_9128,N_6309);
and U14134 (N_14134,N_7979,N_5215);
or U14135 (N_14135,N_7238,N_8655);
and U14136 (N_14136,N_7142,N_7685);
and U14137 (N_14137,N_6979,N_6216);
or U14138 (N_14138,N_6750,N_8558);
xor U14139 (N_14139,N_7376,N_5667);
nand U14140 (N_14140,N_9725,N_9819);
nand U14141 (N_14141,N_8121,N_7250);
nor U14142 (N_14142,N_5647,N_5739);
xnor U14143 (N_14143,N_5376,N_8497);
or U14144 (N_14144,N_7816,N_9275);
nand U14145 (N_14145,N_7832,N_6256);
xnor U14146 (N_14146,N_8417,N_7201);
nand U14147 (N_14147,N_5826,N_6327);
nor U14148 (N_14148,N_7895,N_5211);
xnor U14149 (N_14149,N_7434,N_6308);
or U14150 (N_14150,N_5030,N_9106);
or U14151 (N_14151,N_7539,N_9162);
and U14152 (N_14152,N_5651,N_9141);
nor U14153 (N_14153,N_6030,N_9624);
nand U14154 (N_14154,N_5474,N_5032);
and U14155 (N_14155,N_9664,N_6737);
xnor U14156 (N_14156,N_8762,N_9206);
nand U14157 (N_14157,N_6668,N_6993);
nor U14158 (N_14158,N_6062,N_8127);
nor U14159 (N_14159,N_9532,N_7389);
xnor U14160 (N_14160,N_8333,N_7732);
xor U14161 (N_14161,N_8951,N_8929);
and U14162 (N_14162,N_7890,N_6575);
nor U14163 (N_14163,N_8422,N_5844);
nand U14164 (N_14164,N_7895,N_9876);
and U14165 (N_14165,N_7113,N_7507);
xor U14166 (N_14166,N_7956,N_7598);
nand U14167 (N_14167,N_6569,N_5664);
and U14168 (N_14168,N_7228,N_9370);
nand U14169 (N_14169,N_6278,N_8506);
nand U14170 (N_14170,N_5667,N_8964);
or U14171 (N_14171,N_9956,N_8564);
and U14172 (N_14172,N_7246,N_8466);
and U14173 (N_14173,N_9287,N_7072);
nor U14174 (N_14174,N_5313,N_9791);
or U14175 (N_14175,N_9593,N_7467);
nor U14176 (N_14176,N_8444,N_9272);
nand U14177 (N_14177,N_9159,N_6569);
nand U14178 (N_14178,N_9569,N_8057);
or U14179 (N_14179,N_9266,N_8770);
nand U14180 (N_14180,N_7512,N_7486);
and U14181 (N_14181,N_6063,N_8960);
or U14182 (N_14182,N_8826,N_8286);
nand U14183 (N_14183,N_5429,N_6428);
nor U14184 (N_14184,N_9510,N_9726);
and U14185 (N_14185,N_7240,N_6175);
nand U14186 (N_14186,N_9014,N_8034);
nand U14187 (N_14187,N_6753,N_8865);
xnor U14188 (N_14188,N_7734,N_8606);
xor U14189 (N_14189,N_6456,N_7122);
or U14190 (N_14190,N_5682,N_7758);
nor U14191 (N_14191,N_9679,N_9169);
nor U14192 (N_14192,N_7221,N_8991);
nor U14193 (N_14193,N_6469,N_6679);
and U14194 (N_14194,N_5846,N_7573);
and U14195 (N_14195,N_8894,N_5931);
and U14196 (N_14196,N_8433,N_6620);
and U14197 (N_14197,N_7428,N_5247);
or U14198 (N_14198,N_5202,N_8021);
and U14199 (N_14199,N_6838,N_6240);
nand U14200 (N_14200,N_6858,N_6963);
nand U14201 (N_14201,N_6433,N_8437);
or U14202 (N_14202,N_6884,N_5597);
and U14203 (N_14203,N_9628,N_9583);
nand U14204 (N_14204,N_9085,N_9139);
xor U14205 (N_14205,N_7958,N_9878);
xor U14206 (N_14206,N_6791,N_7356);
nand U14207 (N_14207,N_5324,N_8653);
nor U14208 (N_14208,N_5674,N_7534);
xor U14209 (N_14209,N_9011,N_6183);
or U14210 (N_14210,N_7789,N_5702);
and U14211 (N_14211,N_7129,N_6027);
nand U14212 (N_14212,N_6367,N_5953);
or U14213 (N_14213,N_6309,N_5418);
and U14214 (N_14214,N_6768,N_9589);
and U14215 (N_14215,N_6043,N_7325);
xnor U14216 (N_14216,N_7570,N_5953);
nor U14217 (N_14217,N_7659,N_7147);
and U14218 (N_14218,N_6343,N_7150);
and U14219 (N_14219,N_6867,N_8003);
and U14220 (N_14220,N_5688,N_8080);
nor U14221 (N_14221,N_5547,N_9952);
xor U14222 (N_14222,N_5682,N_8733);
nand U14223 (N_14223,N_6255,N_5123);
and U14224 (N_14224,N_8465,N_6830);
and U14225 (N_14225,N_9340,N_9947);
or U14226 (N_14226,N_8735,N_5572);
or U14227 (N_14227,N_5226,N_8834);
nand U14228 (N_14228,N_6136,N_9069);
or U14229 (N_14229,N_5717,N_5661);
or U14230 (N_14230,N_9800,N_5486);
or U14231 (N_14231,N_8389,N_6545);
and U14232 (N_14232,N_9973,N_7699);
nor U14233 (N_14233,N_5818,N_8245);
nor U14234 (N_14234,N_9565,N_6522);
nand U14235 (N_14235,N_8375,N_7488);
xor U14236 (N_14236,N_5933,N_7138);
xor U14237 (N_14237,N_6025,N_6666);
nor U14238 (N_14238,N_6354,N_6068);
or U14239 (N_14239,N_5103,N_7390);
nand U14240 (N_14240,N_5233,N_6117);
nor U14241 (N_14241,N_6114,N_9003);
or U14242 (N_14242,N_6493,N_5307);
nand U14243 (N_14243,N_8047,N_8801);
or U14244 (N_14244,N_8391,N_6002);
nor U14245 (N_14245,N_5835,N_5998);
nand U14246 (N_14246,N_5849,N_6844);
xor U14247 (N_14247,N_8518,N_8682);
or U14248 (N_14248,N_8477,N_8622);
and U14249 (N_14249,N_6816,N_9895);
nor U14250 (N_14250,N_8887,N_6764);
xnor U14251 (N_14251,N_7583,N_9656);
and U14252 (N_14252,N_7981,N_9782);
or U14253 (N_14253,N_9721,N_9070);
xnor U14254 (N_14254,N_6596,N_8742);
and U14255 (N_14255,N_8463,N_7924);
and U14256 (N_14256,N_8252,N_5772);
nor U14257 (N_14257,N_8365,N_5802);
xnor U14258 (N_14258,N_6494,N_5899);
and U14259 (N_14259,N_6179,N_5526);
nor U14260 (N_14260,N_6039,N_7379);
and U14261 (N_14261,N_6847,N_6439);
and U14262 (N_14262,N_7129,N_6357);
xor U14263 (N_14263,N_6034,N_7581);
and U14264 (N_14264,N_8327,N_6820);
or U14265 (N_14265,N_6285,N_6656);
nand U14266 (N_14266,N_7005,N_7705);
nand U14267 (N_14267,N_6533,N_7089);
nand U14268 (N_14268,N_8763,N_9282);
and U14269 (N_14269,N_9344,N_6593);
nand U14270 (N_14270,N_9342,N_7713);
nor U14271 (N_14271,N_5482,N_7966);
nor U14272 (N_14272,N_7595,N_8280);
or U14273 (N_14273,N_9170,N_7146);
and U14274 (N_14274,N_5681,N_9368);
nor U14275 (N_14275,N_6399,N_7475);
nor U14276 (N_14276,N_5659,N_6911);
and U14277 (N_14277,N_6984,N_7353);
and U14278 (N_14278,N_5334,N_6417);
or U14279 (N_14279,N_5364,N_6792);
nand U14280 (N_14280,N_5743,N_9863);
nand U14281 (N_14281,N_5440,N_5055);
nand U14282 (N_14282,N_8837,N_5054);
nor U14283 (N_14283,N_5979,N_8590);
and U14284 (N_14284,N_7796,N_9634);
nand U14285 (N_14285,N_7728,N_5680);
and U14286 (N_14286,N_7482,N_6404);
xnor U14287 (N_14287,N_5150,N_7208);
xor U14288 (N_14288,N_6084,N_5540);
and U14289 (N_14289,N_7577,N_5153);
nor U14290 (N_14290,N_8430,N_5529);
and U14291 (N_14291,N_6142,N_7449);
xor U14292 (N_14292,N_9591,N_9982);
nand U14293 (N_14293,N_5595,N_9955);
nor U14294 (N_14294,N_8367,N_6575);
and U14295 (N_14295,N_9861,N_9812);
nor U14296 (N_14296,N_8734,N_5189);
or U14297 (N_14297,N_5150,N_5132);
nand U14298 (N_14298,N_5595,N_6288);
and U14299 (N_14299,N_6678,N_5923);
nor U14300 (N_14300,N_7685,N_7866);
nor U14301 (N_14301,N_5600,N_5606);
nor U14302 (N_14302,N_8717,N_7808);
nand U14303 (N_14303,N_8541,N_5320);
nand U14304 (N_14304,N_5865,N_5141);
and U14305 (N_14305,N_6746,N_7748);
and U14306 (N_14306,N_5959,N_5755);
nand U14307 (N_14307,N_5476,N_5116);
nor U14308 (N_14308,N_6503,N_9646);
nor U14309 (N_14309,N_5018,N_5501);
nor U14310 (N_14310,N_6594,N_5602);
nor U14311 (N_14311,N_8768,N_5268);
nor U14312 (N_14312,N_8237,N_8552);
nand U14313 (N_14313,N_6815,N_7628);
nand U14314 (N_14314,N_9521,N_6428);
nand U14315 (N_14315,N_5217,N_5175);
nand U14316 (N_14316,N_6860,N_8213);
nand U14317 (N_14317,N_6442,N_9266);
nor U14318 (N_14318,N_7528,N_7695);
nor U14319 (N_14319,N_6285,N_8196);
nand U14320 (N_14320,N_7416,N_8841);
nand U14321 (N_14321,N_9792,N_6958);
and U14322 (N_14322,N_8511,N_5430);
nor U14323 (N_14323,N_8818,N_9619);
nor U14324 (N_14324,N_8730,N_8530);
nand U14325 (N_14325,N_5764,N_7259);
and U14326 (N_14326,N_7553,N_7367);
nand U14327 (N_14327,N_9168,N_6698);
or U14328 (N_14328,N_5524,N_8885);
or U14329 (N_14329,N_6756,N_5826);
or U14330 (N_14330,N_8822,N_9921);
or U14331 (N_14331,N_6184,N_5786);
xor U14332 (N_14332,N_7314,N_8633);
and U14333 (N_14333,N_5829,N_8892);
or U14334 (N_14334,N_6542,N_9572);
nor U14335 (N_14335,N_9931,N_8391);
or U14336 (N_14336,N_9490,N_8338);
or U14337 (N_14337,N_9014,N_7225);
and U14338 (N_14338,N_9092,N_7862);
and U14339 (N_14339,N_8963,N_9597);
nor U14340 (N_14340,N_6200,N_8934);
nand U14341 (N_14341,N_5663,N_6590);
or U14342 (N_14342,N_8629,N_8786);
or U14343 (N_14343,N_7602,N_9329);
and U14344 (N_14344,N_8040,N_8956);
nand U14345 (N_14345,N_9204,N_9908);
and U14346 (N_14346,N_8432,N_9547);
nand U14347 (N_14347,N_8966,N_5070);
nand U14348 (N_14348,N_5000,N_8284);
and U14349 (N_14349,N_6093,N_9234);
or U14350 (N_14350,N_9873,N_6251);
and U14351 (N_14351,N_9488,N_5703);
and U14352 (N_14352,N_8575,N_9812);
or U14353 (N_14353,N_6634,N_9842);
nor U14354 (N_14354,N_8378,N_7398);
nand U14355 (N_14355,N_7942,N_9875);
or U14356 (N_14356,N_9645,N_6624);
and U14357 (N_14357,N_8957,N_7730);
and U14358 (N_14358,N_6367,N_7229);
nor U14359 (N_14359,N_6402,N_8394);
nor U14360 (N_14360,N_9232,N_5332);
nor U14361 (N_14361,N_8383,N_8660);
and U14362 (N_14362,N_7247,N_7366);
xnor U14363 (N_14363,N_8704,N_6702);
and U14364 (N_14364,N_7752,N_9208);
and U14365 (N_14365,N_8534,N_6645);
and U14366 (N_14366,N_8115,N_5469);
nor U14367 (N_14367,N_5814,N_6801);
and U14368 (N_14368,N_6639,N_9330);
or U14369 (N_14369,N_7745,N_9924);
nand U14370 (N_14370,N_6223,N_5922);
nand U14371 (N_14371,N_5809,N_6234);
nand U14372 (N_14372,N_8048,N_5164);
nor U14373 (N_14373,N_6497,N_7828);
nor U14374 (N_14374,N_8246,N_9631);
nor U14375 (N_14375,N_8937,N_9272);
nor U14376 (N_14376,N_8233,N_8008);
nand U14377 (N_14377,N_5092,N_5530);
nor U14378 (N_14378,N_5325,N_5629);
nand U14379 (N_14379,N_8053,N_8195);
xnor U14380 (N_14380,N_7210,N_5594);
or U14381 (N_14381,N_5697,N_6976);
xnor U14382 (N_14382,N_5970,N_8167);
or U14383 (N_14383,N_8725,N_7830);
nor U14384 (N_14384,N_9222,N_8256);
or U14385 (N_14385,N_7538,N_6987);
or U14386 (N_14386,N_8535,N_5154);
or U14387 (N_14387,N_9035,N_8096);
or U14388 (N_14388,N_7457,N_7246);
xnor U14389 (N_14389,N_6209,N_5477);
nor U14390 (N_14390,N_8077,N_9373);
nor U14391 (N_14391,N_6452,N_6337);
and U14392 (N_14392,N_9459,N_7488);
nand U14393 (N_14393,N_8496,N_9498);
or U14394 (N_14394,N_8461,N_9738);
nor U14395 (N_14395,N_7761,N_6600);
nor U14396 (N_14396,N_7382,N_5697);
nor U14397 (N_14397,N_7900,N_6052);
xnor U14398 (N_14398,N_9504,N_9571);
nand U14399 (N_14399,N_7738,N_8342);
or U14400 (N_14400,N_8472,N_8451);
or U14401 (N_14401,N_6165,N_6987);
xnor U14402 (N_14402,N_8098,N_9621);
or U14403 (N_14403,N_6512,N_7723);
or U14404 (N_14404,N_7401,N_7907);
nor U14405 (N_14405,N_7351,N_8715);
nor U14406 (N_14406,N_5821,N_8427);
or U14407 (N_14407,N_8756,N_5822);
xor U14408 (N_14408,N_8129,N_8599);
and U14409 (N_14409,N_8004,N_6164);
or U14410 (N_14410,N_8433,N_6854);
or U14411 (N_14411,N_7655,N_5244);
and U14412 (N_14412,N_6685,N_9222);
xor U14413 (N_14413,N_9357,N_5347);
nor U14414 (N_14414,N_8037,N_8177);
or U14415 (N_14415,N_6721,N_8531);
or U14416 (N_14416,N_7670,N_9456);
nor U14417 (N_14417,N_9250,N_6435);
nor U14418 (N_14418,N_7416,N_7105);
nor U14419 (N_14419,N_5485,N_9219);
nor U14420 (N_14420,N_8070,N_6127);
and U14421 (N_14421,N_6460,N_8041);
or U14422 (N_14422,N_8957,N_8598);
and U14423 (N_14423,N_5994,N_8283);
nor U14424 (N_14424,N_9802,N_6379);
nor U14425 (N_14425,N_5196,N_7748);
or U14426 (N_14426,N_7433,N_8124);
and U14427 (N_14427,N_5498,N_7191);
nor U14428 (N_14428,N_9463,N_6281);
and U14429 (N_14429,N_8304,N_6818);
and U14430 (N_14430,N_7284,N_7676);
and U14431 (N_14431,N_7016,N_6174);
or U14432 (N_14432,N_8434,N_7534);
xnor U14433 (N_14433,N_7178,N_8313);
nand U14434 (N_14434,N_5661,N_5174);
or U14435 (N_14435,N_9540,N_8474);
and U14436 (N_14436,N_7301,N_7185);
nand U14437 (N_14437,N_5140,N_5311);
nand U14438 (N_14438,N_9523,N_8617);
and U14439 (N_14439,N_9167,N_5805);
nor U14440 (N_14440,N_9422,N_6526);
and U14441 (N_14441,N_7394,N_9172);
and U14442 (N_14442,N_5913,N_6580);
xnor U14443 (N_14443,N_8268,N_6121);
and U14444 (N_14444,N_5536,N_7369);
and U14445 (N_14445,N_8556,N_7373);
or U14446 (N_14446,N_8431,N_9736);
nor U14447 (N_14447,N_7355,N_9265);
and U14448 (N_14448,N_5877,N_8814);
or U14449 (N_14449,N_9286,N_6503);
xor U14450 (N_14450,N_7309,N_6663);
nor U14451 (N_14451,N_9480,N_8337);
nor U14452 (N_14452,N_9720,N_5241);
or U14453 (N_14453,N_9542,N_7123);
nor U14454 (N_14454,N_8426,N_7793);
nor U14455 (N_14455,N_5760,N_7795);
nand U14456 (N_14456,N_7749,N_8845);
nor U14457 (N_14457,N_8449,N_6628);
or U14458 (N_14458,N_6887,N_9774);
and U14459 (N_14459,N_8681,N_8876);
xor U14460 (N_14460,N_9475,N_6766);
or U14461 (N_14461,N_5386,N_6976);
nor U14462 (N_14462,N_7538,N_8862);
and U14463 (N_14463,N_9278,N_6047);
nor U14464 (N_14464,N_5235,N_6452);
nor U14465 (N_14465,N_9884,N_8930);
nor U14466 (N_14466,N_7726,N_5739);
and U14467 (N_14467,N_6546,N_5267);
and U14468 (N_14468,N_6943,N_7963);
nand U14469 (N_14469,N_9443,N_5203);
nand U14470 (N_14470,N_6803,N_8771);
nand U14471 (N_14471,N_9214,N_8396);
nand U14472 (N_14472,N_5125,N_9622);
nand U14473 (N_14473,N_6226,N_7665);
nor U14474 (N_14474,N_9793,N_6743);
and U14475 (N_14475,N_6131,N_8461);
and U14476 (N_14476,N_6739,N_9134);
or U14477 (N_14477,N_9657,N_7145);
and U14478 (N_14478,N_5168,N_9379);
nor U14479 (N_14479,N_9670,N_5097);
xor U14480 (N_14480,N_5993,N_6119);
and U14481 (N_14481,N_8104,N_8662);
and U14482 (N_14482,N_9802,N_5770);
nand U14483 (N_14483,N_8222,N_9562);
and U14484 (N_14484,N_8081,N_5766);
nor U14485 (N_14485,N_9748,N_9456);
nand U14486 (N_14486,N_8277,N_8850);
and U14487 (N_14487,N_7826,N_7677);
or U14488 (N_14488,N_8657,N_5534);
xnor U14489 (N_14489,N_9408,N_6822);
or U14490 (N_14490,N_9253,N_5092);
nor U14491 (N_14491,N_6162,N_6291);
nor U14492 (N_14492,N_9448,N_9159);
or U14493 (N_14493,N_6577,N_8297);
xnor U14494 (N_14494,N_6992,N_7260);
nand U14495 (N_14495,N_7513,N_5376);
nand U14496 (N_14496,N_9559,N_8591);
and U14497 (N_14497,N_7438,N_8021);
or U14498 (N_14498,N_8898,N_7981);
nand U14499 (N_14499,N_6087,N_8400);
and U14500 (N_14500,N_7652,N_6988);
nand U14501 (N_14501,N_9347,N_5016);
nand U14502 (N_14502,N_7374,N_7530);
xor U14503 (N_14503,N_6740,N_6460);
or U14504 (N_14504,N_7661,N_5711);
or U14505 (N_14505,N_5698,N_9622);
xnor U14506 (N_14506,N_6155,N_5280);
xnor U14507 (N_14507,N_5666,N_5085);
nor U14508 (N_14508,N_5291,N_8920);
and U14509 (N_14509,N_6029,N_7426);
and U14510 (N_14510,N_9279,N_8269);
or U14511 (N_14511,N_5842,N_7485);
nor U14512 (N_14512,N_8634,N_6931);
xnor U14513 (N_14513,N_7012,N_5768);
or U14514 (N_14514,N_8401,N_9318);
or U14515 (N_14515,N_7285,N_5731);
nand U14516 (N_14516,N_7577,N_8312);
or U14517 (N_14517,N_5360,N_8495);
nor U14518 (N_14518,N_9475,N_8416);
and U14519 (N_14519,N_8754,N_6130);
nand U14520 (N_14520,N_5333,N_6147);
and U14521 (N_14521,N_5644,N_7602);
xnor U14522 (N_14522,N_9202,N_5230);
or U14523 (N_14523,N_8306,N_7090);
nand U14524 (N_14524,N_5385,N_7914);
nor U14525 (N_14525,N_8640,N_8687);
xor U14526 (N_14526,N_5490,N_7655);
or U14527 (N_14527,N_8336,N_6816);
or U14528 (N_14528,N_7247,N_9253);
nor U14529 (N_14529,N_7304,N_5047);
and U14530 (N_14530,N_5351,N_9907);
xor U14531 (N_14531,N_9715,N_9370);
or U14532 (N_14532,N_8316,N_7148);
or U14533 (N_14533,N_6033,N_8819);
nor U14534 (N_14534,N_8344,N_6184);
nand U14535 (N_14535,N_5044,N_8763);
nor U14536 (N_14536,N_6179,N_9657);
or U14537 (N_14537,N_6618,N_9501);
nor U14538 (N_14538,N_7549,N_7739);
and U14539 (N_14539,N_6565,N_8570);
nand U14540 (N_14540,N_6914,N_7652);
nand U14541 (N_14541,N_5492,N_9846);
xnor U14542 (N_14542,N_7876,N_5946);
xor U14543 (N_14543,N_9505,N_9011);
nand U14544 (N_14544,N_8035,N_5303);
and U14545 (N_14545,N_7444,N_5588);
xor U14546 (N_14546,N_9214,N_7069);
or U14547 (N_14547,N_5373,N_7839);
nand U14548 (N_14548,N_8285,N_7841);
or U14549 (N_14549,N_5792,N_7132);
or U14550 (N_14550,N_5051,N_8038);
nor U14551 (N_14551,N_6723,N_8468);
nor U14552 (N_14552,N_9295,N_8847);
nor U14553 (N_14553,N_9632,N_6902);
xor U14554 (N_14554,N_5456,N_7116);
and U14555 (N_14555,N_9131,N_6424);
and U14556 (N_14556,N_9359,N_6616);
nand U14557 (N_14557,N_6919,N_6950);
and U14558 (N_14558,N_8662,N_5962);
or U14559 (N_14559,N_7388,N_7493);
nor U14560 (N_14560,N_6499,N_6404);
or U14561 (N_14561,N_8267,N_5310);
or U14562 (N_14562,N_7047,N_8949);
or U14563 (N_14563,N_7519,N_7909);
nand U14564 (N_14564,N_7883,N_5822);
xnor U14565 (N_14565,N_8294,N_9672);
nand U14566 (N_14566,N_7749,N_9147);
nor U14567 (N_14567,N_7895,N_5231);
nand U14568 (N_14568,N_6384,N_7534);
nor U14569 (N_14569,N_9294,N_9440);
or U14570 (N_14570,N_8583,N_5887);
or U14571 (N_14571,N_9579,N_5435);
nand U14572 (N_14572,N_9843,N_6382);
or U14573 (N_14573,N_5341,N_8093);
xor U14574 (N_14574,N_5630,N_6828);
nand U14575 (N_14575,N_7423,N_6260);
or U14576 (N_14576,N_5059,N_8120);
or U14577 (N_14577,N_5080,N_5381);
nand U14578 (N_14578,N_9360,N_7915);
and U14579 (N_14579,N_9791,N_8937);
nor U14580 (N_14580,N_8648,N_8686);
nor U14581 (N_14581,N_6660,N_7244);
and U14582 (N_14582,N_6996,N_6842);
nand U14583 (N_14583,N_8512,N_5679);
or U14584 (N_14584,N_6604,N_6805);
nor U14585 (N_14585,N_5713,N_7564);
nor U14586 (N_14586,N_7756,N_6581);
or U14587 (N_14587,N_6642,N_5678);
and U14588 (N_14588,N_6493,N_5712);
or U14589 (N_14589,N_8264,N_7433);
nor U14590 (N_14590,N_8760,N_5252);
and U14591 (N_14591,N_7564,N_7699);
or U14592 (N_14592,N_6672,N_9757);
xnor U14593 (N_14593,N_7595,N_5811);
nor U14594 (N_14594,N_6565,N_5353);
nor U14595 (N_14595,N_6112,N_7937);
and U14596 (N_14596,N_8824,N_8810);
nand U14597 (N_14597,N_8042,N_7379);
xor U14598 (N_14598,N_7873,N_5526);
and U14599 (N_14599,N_7189,N_5114);
nand U14600 (N_14600,N_7403,N_7081);
nand U14601 (N_14601,N_7903,N_6580);
and U14602 (N_14602,N_9850,N_9808);
and U14603 (N_14603,N_5065,N_9151);
nor U14604 (N_14604,N_8432,N_6795);
nor U14605 (N_14605,N_9311,N_9234);
or U14606 (N_14606,N_7321,N_8231);
nand U14607 (N_14607,N_6569,N_6836);
or U14608 (N_14608,N_9229,N_5553);
nand U14609 (N_14609,N_9390,N_9301);
nand U14610 (N_14610,N_6014,N_8405);
and U14611 (N_14611,N_6945,N_5295);
nor U14612 (N_14612,N_7506,N_5494);
and U14613 (N_14613,N_9238,N_7358);
nand U14614 (N_14614,N_8572,N_5877);
and U14615 (N_14615,N_6947,N_5820);
nand U14616 (N_14616,N_8480,N_7602);
nor U14617 (N_14617,N_5953,N_9838);
xnor U14618 (N_14618,N_9036,N_5968);
xor U14619 (N_14619,N_5949,N_5390);
nor U14620 (N_14620,N_6228,N_5327);
and U14621 (N_14621,N_7922,N_7735);
xor U14622 (N_14622,N_7534,N_6827);
or U14623 (N_14623,N_8572,N_6377);
xnor U14624 (N_14624,N_9949,N_7092);
and U14625 (N_14625,N_9443,N_8674);
and U14626 (N_14626,N_6035,N_7184);
nand U14627 (N_14627,N_5014,N_9828);
xnor U14628 (N_14628,N_8142,N_8921);
or U14629 (N_14629,N_9772,N_8103);
and U14630 (N_14630,N_8439,N_9541);
nor U14631 (N_14631,N_7002,N_9185);
or U14632 (N_14632,N_8963,N_8840);
or U14633 (N_14633,N_8596,N_9722);
and U14634 (N_14634,N_8491,N_8587);
nor U14635 (N_14635,N_7634,N_6305);
nor U14636 (N_14636,N_7045,N_9281);
nand U14637 (N_14637,N_6823,N_7734);
nor U14638 (N_14638,N_5139,N_7754);
or U14639 (N_14639,N_8164,N_9739);
xor U14640 (N_14640,N_6368,N_9693);
or U14641 (N_14641,N_6340,N_6009);
or U14642 (N_14642,N_7918,N_7034);
xnor U14643 (N_14643,N_8512,N_7369);
nor U14644 (N_14644,N_8186,N_9558);
nand U14645 (N_14645,N_5224,N_9720);
xnor U14646 (N_14646,N_8956,N_8858);
nand U14647 (N_14647,N_6823,N_9100);
or U14648 (N_14648,N_7859,N_5854);
nand U14649 (N_14649,N_8610,N_6417);
or U14650 (N_14650,N_6004,N_7209);
or U14651 (N_14651,N_8470,N_9806);
and U14652 (N_14652,N_8540,N_8095);
xnor U14653 (N_14653,N_6856,N_5968);
and U14654 (N_14654,N_9087,N_8090);
nand U14655 (N_14655,N_6363,N_8354);
or U14656 (N_14656,N_5748,N_5149);
or U14657 (N_14657,N_9021,N_5061);
nand U14658 (N_14658,N_6304,N_5976);
xor U14659 (N_14659,N_8079,N_5490);
or U14660 (N_14660,N_7911,N_9423);
nand U14661 (N_14661,N_9037,N_9212);
nand U14662 (N_14662,N_5242,N_5815);
or U14663 (N_14663,N_5381,N_6891);
nand U14664 (N_14664,N_6548,N_7818);
nor U14665 (N_14665,N_6820,N_8772);
nor U14666 (N_14666,N_8936,N_5103);
and U14667 (N_14667,N_5232,N_9555);
or U14668 (N_14668,N_8174,N_6028);
or U14669 (N_14669,N_9912,N_9060);
nand U14670 (N_14670,N_6705,N_9012);
and U14671 (N_14671,N_6690,N_7497);
and U14672 (N_14672,N_7209,N_7897);
nand U14673 (N_14673,N_5235,N_5918);
and U14674 (N_14674,N_7764,N_9445);
or U14675 (N_14675,N_7705,N_6910);
and U14676 (N_14676,N_8508,N_8413);
nand U14677 (N_14677,N_8591,N_6622);
or U14678 (N_14678,N_7541,N_5670);
nand U14679 (N_14679,N_8941,N_7056);
nor U14680 (N_14680,N_7018,N_5023);
nand U14681 (N_14681,N_5537,N_9472);
nor U14682 (N_14682,N_7673,N_5731);
nand U14683 (N_14683,N_6847,N_8234);
nand U14684 (N_14684,N_7560,N_8637);
and U14685 (N_14685,N_9706,N_9426);
nand U14686 (N_14686,N_8779,N_5008);
xor U14687 (N_14687,N_8430,N_6015);
nor U14688 (N_14688,N_5986,N_6959);
nor U14689 (N_14689,N_7945,N_6783);
xor U14690 (N_14690,N_5868,N_5203);
nand U14691 (N_14691,N_6659,N_5498);
and U14692 (N_14692,N_7827,N_6383);
xnor U14693 (N_14693,N_5040,N_8807);
and U14694 (N_14694,N_5919,N_6305);
nor U14695 (N_14695,N_8049,N_7884);
nand U14696 (N_14696,N_6724,N_6618);
or U14697 (N_14697,N_5724,N_8531);
and U14698 (N_14698,N_6257,N_6781);
or U14699 (N_14699,N_6991,N_8205);
or U14700 (N_14700,N_9700,N_8155);
nand U14701 (N_14701,N_7102,N_6535);
nor U14702 (N_14702,N_6598,N_8981);
or U14703 (N_14703,N_9544,N_5024);
nor U14704 (N_14704,N_5636,N_9379);
xnor U14705 (N_14705,N_8202,N_7752);
or U14706 (N_14706,N_7295,N_6141);
xnor U14707 (N_14707,N_9483,N_5818);
xnor U14708 (N_14708,N_8405,N_6847);
or U14709 (N_14709,N_7201,N_6792);
nor U14710 (N_14710,N_6478,N_5828);
nand U14711 (N_14711,N_8426,N_9029);
or U14712 (N_14712,N_6048,N_8853);
nand U14713 (N_14713,N_5691,N_5235);
nor U14714 (N_14714,N_5369,N_6941);
nor U14715 (N_14715,N_7680,N_9636);
xnor U14716 (N_14716,N_9868,N_9011);
and U14717 (N_14717,N_9820,N_7531);
nor U14718 (N_14718,N_6723,N_7214);
and U14719 (N_14719,N_8349,N_9032);
or U14720 (N_14720,N_7451,N_9876);
and U14721 (N_14721,N_8409,N_6648);
xnor U14722 (N_14722,N_6181,N_8981);
nand U14723 (N_14723,N_6486,N_9266);
or U14724 (N_14724,N_9715,N_8985);
or U14725 (N_14725,N_5646,N_9221);
nand U14726 (N_14726,N_9818,N_6350);
nand U14727 (N_14727,N_6828,N_9589);
nor U14728 (N_14728,N_7770,N_7441);
or U14729 (N_14729,N_8608,N_5690);
or U14730 (N_14730,N_7575,N_5620);
xnor U14731 (N_14731,N_5698,N_9890);
and U14732 (N_14732,N_6069,N_7060);
and U14733 (N_14733,N_8599,N_9973);
xor U14734 (N_14734,N_7237,N_8914);
or U14735 (N_14735,N_5015,N_5476);
nor U14736 (N_14736,N_7357,N_7167);
nand U14737 (N_14737,N_7694,N_6530);
and U14738 (N_14738,N_8647,N_8373);
nor U14739 (N_14739,N_8225,N_6014);
nand U14740 (N_14740,N_6619,N_5672);
xnor U14741 (N_14741,N_9553,N_9385);
nor U14742 (N_14742,N_8222,N_6539);
and U14743 (N_14743,N_9548,N_9465);
or U14744 (N_14744,N_9794,N_9772);
nor U14745 (N_14745,N_5920,N_6589);
and U14746 (N_14746,N_5875,N_8890);
nand U14747 (N_14747,N_9939,N_8547);
nor U14748 (N_14748,N_6869,N_5328);
and U14749 (N_14749,N_5850,N_7224);
nand U14750 (N_14750,N_7488,N_7680);
nor U14751 (N_14751,N_8569,N_8270);
and U14752 (N_14752,N_7430,N_9941);
nand U14753 (N_14753,N_6334,N_7438);
or U14754 (N_14754,N_5408,N_8996);
nand U14755 (N_14755,N_5854,N_7229);
nor U14756 (N_14756,N_5687,N_7672);
or U14757 (N_14757,N_8003,N_5596);
xor U14758 (N_14758,N_6412,N_8329);
nor U14759 (N_14759,N_7488,N_5720);
xnor U14760 (N_14760,N_7841,N_5204);
nor U14761 (N_14761,N_5775,N_5494);
or U14762 (N_14762,N_9950,N_8790);
or U14763 (N_14763,N_8218,N_9292);
or U14764 (N_14764,N_8199,N_7039);
nand U14765 (N_14765,N_8520,N_6665);
nand U14766 (N_14766,N_6834,N_5178);
nand U14767 (N_14767,N_6327,N_6631);
and U14768 (N_14768,N_6825,N_9237);
nor U14769 (N_14769,N_8744,N_9540);
nor U14770 (N_14770,N_8449,N_9074);
nor U14771 (N_14771,N_8688,N_8343);
nand U14772 (N_14772,N_6422,N_5024);
nor U14773 (N_14773,N_9139,N_6007);
and U14774 (N_14774,N_7528,N_7079);
xnor U14775 (N_14775,N_5890,N_7540);
nor U14776 (N_14776,N_5058,N_6054);
or U14777 (N_14777,N_5322,N_5308);
or U14778 (N_14778,N_7881,N_9517);
nor U14779 (N_14779,N_5664,N_6683);
or U14780 (N_14780,N_5704,N_9931);
nand U14781 (N_14781,N_9596,N_9732);
nand U14782 (N_14782,N_6708,N_8820);
nand U14783 (N_14783,N_8124,N_9798);
nand U14784 (N_14784,N_8667,N_7703);
nor U14785 (N_14785,N_9925,N_5737);
nand U14786 (N_14786,N_7363,N_6538);
nand U14787 (N_14787,N_5506,N_5128);
nand U14788 (N_14788,N_9774,N_6171);
and U14789 (N_14789,N_6411,N_9463);
nand U14790 (N_14790,N_8518,N_9700);
and U14791 (N_14791,N_5874,N_8809);
nor U14792 (N_14792,N_8720,N_5367);
and U14793 (N_14793,N_7096,N_7157);
nor U14794 (N_14794,N_7442,N_9266);
nor U14795 (N_14795,N_5694,N_8524);
nor U14796 (N_14796,N_9129,N_7853);
or U14797 (N_14797,N_8972,N_6006);
and U14798 (N_14798,N_6977,N_6736);
and U14799 (N_14799,N_6442,N_5074);
or U14800 (N_14800,N_5781,N_7184);
or U14801 (N_14801,N_6627,N_7485);
or U14802 (N_14802,N_8838,N_6770);
nor U14803 (N_14803,N_5907,N_6657);
xnor U14804 (N_14804,N_8977,N_9031);
xor U14805 (N_14805,N_8769,N_6677);
xnor U14806 (N_14806,N_5739,N_8428);
nand U14807 (N_14807,N_6614,N_9157);
nand U14808 (N_14808,N_9266,N_8670);
nor U14809 (N_14809,N_9880,N_6748);
nand U14810 (N_14810,N_9620,N_6151);
nand U14811 (N_14811,N_7873,N_7505);
nand U14812 (N_14812,N_5848,N_6327);
nand U14813 (N_14813,N_8530,N_6548);
and U14814 (N_14814,N_7057,N_8709);
and U14815 (N_14815,N_5132,N_6344);
and U14816 (N_14816,N_8502,N_7611);
nand U14817 (N_14817,N_9623,N_8991);
nor U14818 (N_14818,N_7870,N_9504);
xor U14819 (N_14819,N_8568,N_5666);
and U14820 (N_14820,N_9975,N_9945);
and U14821 (N_14821,N_7584,N_7760);
nand U14822 (N_14822,N_8156,N_7077);
and U14823 (N_14823,N_8327,N_6518);
or U14824 (N_14824,N_9129,N_9717);
and U14825 (N_14825,N_5128,N_7531);
nor U14826 (N_14826,N_6872,N_6198);
or U14827 (N_14827,N_7410,N_7767);
nand U14828 (N_14828,N_7646,N_5349);
nand U14829 (N_14829,N_7719,N_7555);
and U14830 (N_14830,N_6077,N_7462);
or U14831 (N_14831,N_9476,N_7131);
or U14832 (N_14832,N_8952,N_9234);
and U14833 (N_14833,N_7564,N_7537);
nor U14834 (N_14834,N_8761,N_7415);
nor U14835 (N_14835,N_8333,N_7074);
nor U14836 (N_14836,N_8319,N_5781);
nor U14837 (N_14837,N_5729,N_6290);
xor U14838 (N_14838,N_8478,N_5320);
nor U14839 (N_14839,N_6563,N_9050);
and U14840 (N_14840,N_6907,N_7277);
or U14841 (N_14841,N_9178,N_7837);
nor U14842 (N_14842,N_6634,N_8882);
and U14843 (N_14843,N_6944,N_9080);
xnor U14844 (N_14844,N_7455,N_6302);
nand U14845 (N_14845,N_9653,N_9854);
nor U14846 (N_14846,N_6145,N_7885);
nand U14847 (N_14847,N_8268,N_7121);
nand U14848 (N_14848,N_8678,N_6399);
nor U14849 (N_14849,N_5692,N_8477);
nor U14850 (N_14850,N_7765,N_8201);
xnor U14851 (N_14851,N_5920,N_8870);
xor U14852 (N_14852,N_6857,N_5501);
nand U14853 (N_14853,N_7822,N_7047);
and U14854 (N_14854,N_8721,N_8757);
nor U14855 (N_14855,N_5701,N_9152);
or U14856 (N_14856,N_5265,N_9755);
and U14857 (N_14857,N_8117,N_9456);
xnor U14858 (N_14858,N_9407,N_5278);
and U14859 (N_14859,N_9685,N_7284);
and U14860 (N_14860,N_7115,N_8112);
nand U14861 (N_14861,N_9653,N_8408);
nand U14862 (N_14862,N_9404,N_8010);
or U14863 (N_14863,N_5442,N_5961);
xor U14864 (N_14864,N_5535,N_8281);
and U14865 (N_14865,N_8348,N_6168);
nor U14866 (N_14866,N_7646,N_9478);
nor U14867 (N_14867,N_6712,N_8703);
nor U14868 (N_14868,N_5120,N_8000);
nand U14869 (N_14869,N_5272,N_8973);
and U14870 (N_14870,N_7614,N_9133);
nor U14871 (N_14871,N_8395,N_8381);
nand U14872 (N_14872,N_7893,N_5032);
nand U14873 (N_14873,N_9136,N_5035);
nor U14874 (N_14874,N_8808,N_6379);
nand U14875 (N_14875,N_8214,N_5614);
and U14876 (N_14876,N_6067,N_8858);
nand U14877 (N_14877,N_5067,N_9209);
nand U14878 (N_14878,N_5208,N_7160);
or U14879 (N_14879,N_7205,N_7914);
nand U14880 (N_14880,N_5264,N_5102);
or U14881 (N_14881,N_7754,N_9854);
or U14882 (N_14882,N_5181,N_7733);
nor U14883 (N_14883,N_6715,N_7876);
nor U14884 (N_14884,N_8640,N_9008);
xnor U14885 (N_14885,N_7623,N_8359);
nor U14886 (N_14886,N_6873,N_6795);
nand U14887 (N_14887,N_8311,N_6336);
xor U14888 (N_14888,N_9497,N_9591);
nand U14889 (N_14889,N_8684,N_5832);
nor U14890 (N_14890,N_8265,N_6136);
nand U14891 (N_14891,N_9835,N_8660);
or U14892 (N_14892,N_8524,N_9946);
nor U14893 (N_14893,N_8774,N_8157);
or U14894 (N_14894,N_8334,N_5954);
nor U14895 (N_14895,N_6231,N_6646);
nand U14896 (N_14896,N_5316,N_8353);
and U14897 (N_14897,N_9053,N_6228);
and U14898 (N_14898,N_5062,N_7643);
xnor U14899 (N_14899,N_7957,N_5710);
or U14900 (N_14900,N_8031,N_6513);
nor U14901 (N_14901,N_6811,N_7591);
nand U14902 (N_14902,N_7205,N_9448);
or U14903 (N_14903,N_6267,N_6697);
nor U14904 (N_14904,N_5370,N_7929);
nor U14905 (N_14905,N_7306,N_7192);
xor U14906 (N_14906,N_6201,N_5500);
xor U14907 (N_14907,N_9734,N_6593);
or U14908 (N_14908,N_8617,N_6164);
nand U14909 (N_14909,N_5505,N_9981);
and U14910 (N_14910,N_9610,N_8742);
nand U14911 (N_14911,N_5819,N_8389);
or U14912 (N_14912,N_6668,N_6966);
and U14913 (N_14913,N_6486,N_7108);
xnor U14914 (N_14914,N_9491,N_9504);
nor U14915 (N_14915,N_6239,N_9050);
nor U14916 (N_14916,N_5465,N_5957);
or U14917 (N_14917,N_5218,N_8048);
nor U14918 (N_14918,N_8584,N_9695);
or U14919 (N_14919,N_9427,N_7502);
or U14920 (N_14920,N_9236,N_7122);
nor U14921 (N_14921,N_8965,N_7063);
and U14922 (N_14922,N_7859,N_5554);
nor U14923 (N_14923,N_9176,N_9792);
and U14924 (N_14924,N_7847,N_7872);
xor U14925 (N_14925,N_7153,N_6294);
nand U14926 (N_14926,N_9955,N_8244);
nand U14927 (N_14927,N_7731,N_8495);
nand U14928 (N_14928,N_6606,N_5261);
nand U14929 (N_14929,N_5662,N_7139);
nand U14930 (N_14930,N_9687,N_7969);
or U14931 (N_14931,N_6515,N_7922);
nand U14932 (N_14932,N_7043,N_5192);
or U14933 (N_14933,N_7220,N_5694);
and U14934 (N_14934,N_7975,N_8209);
and U14935 (N_14935,N_7835,N_5209);
nand U14936 (N_14936,N_8057,N_9680);
or U14937 (N_14937,N_7320,N_8614);
nor U14938 (N_14938,N_6398,N_7041);
nor U14939 (N_14939,N_6687,N_5893);
and U14940 (N_14940,N_7538,N_5086);
nor U14941 (N_14941,N_6583,N_5177);
xnor U14942 (N_14942,N_9043,N_9823);
or U14943 (N_14943,N_5273,N_7795);
xor U14944 (N_14944,N_7553,N_9622);
or U14945 (N_14945,N_8010,N_5948);
and U14946 (N_14946,N_7908,N_9943);
and U14947 (N_14947,N_5275,N_9725);
and U14948 (N_14948,N_9617,N_5891);
or U14949 (N_14949,N_7549,N_6927);
or U14950 (N_14950,N_5370,N_9908);
xor U14951 (N_14951,N_9487,N_8020);
or U14952 (N_14952,N_5483,N_5707);
or U14953 (N_14953,N_8590,N_8417);
and U14954 (N_14954,N_7476,N_9231);
and U14955 (N_14955,N_8224,N_6868);
nand U14956 (N_14956,N_8473,N_9971);
nand U14957 (N_14957,N_8458,N_9516);
and U14958 (N_14958,N_5659,N_5409);
nand U14959 (N_14959,N_9076,N_6470);
xor U14960 (N_14960,N_5286,N_7355);
and U14961 (N_14961,N_9090,N_8197);
nor U14962 (N_14962,N_6076,N_5181);
or U14963 (N_14963,N_8635,N_6414);
and U14964 (N_14964,N_5854,N_9718);
xnor U14965 (N_14965,N_6871,N_8616);
nand U14966 (N_14966,N_6495,N_8231);
nand U14967 (N_14967,N_5685,N_9146);
xnor U14968 (N_14968,N_6013,N_7685);
nand U14969 (N_14969,N_9445,N_6869);
or U14970 (N_14970,N_9072,N_8445);
and U14971 (N_14971,N_5901,N_5137);
nor U14972 (N_14972,N_6736,N_8724);
or U14973 (N_14973,N_9856,N_9426);
and U14974 (N_14974,N_5080,N_9257);
or U14975 (N_14975,N_7218,N_9116);
and U14976 (N_14976,N_6130,N_8894);
or U14977 (N_14977,N_5869,N_7891);
nand U14978 (N_14978,N_7892,N_6231);
or U14979 (N_14979,N_8922,N_6989);
and U14980 (N_14980,N_9886,N_9990);
or U14981 (N_14981,N_5347,N_9902);
or U14982 (N_14982,N_6390,N_5981);
or U14983 (N_14983,N_9712,N_9872);
and U14984 (N_14984,N_5313,N_9470);
and U14985 (N_14985,N_5643,N_7438);
or U14986 (N_14986,N_6336,N_6343);
nor U14987 (N_14987,N_6475,N_8399);
nand U14988 (N_14988,N_7711,N_8457);
nand U14989 (N_14989,N_9865,N_7684);
nor U14990 (N_14990,N_5926,N_7017);
nor U14991 (N_14991,N_7100,N_8324);
nand U14992 (N_14992,N_6316,N_6852);
xor U14993 (N_14993,N_6102,N_6195);
nor U14994 (N_14994,N_5897,N_5174);
nor U14995 (N_14995,N_8058,N_9668);
and U14996 (N_14996,N_7500,N_7211);
nor U14997 (N_14997,N_8883,N_6003);
and U14998 (N_14998,N_7305,N_6491);
and U14999 (N_14999,N_9632,N_9726);
nand U15000 (N_15000,N_12602,N_12676);
or U15001 (N_15001,N_10825,N_12485);
nor U15002 (N_15002,N_10301,N_13181);
nor U15003 (N_15003,N_13264,N_11503);
and U15004 (N_15004,N_11032,N_14515);
nand U15005 (N_15005,N_11436,N_11019);
nand U15006 (N_15006,N_10818,N_14664);
nand U15007 (N_15007,N_10789,N_12193);
nor U15008 (N_15008,N_10277,N_13759);
nand U15009 (N_15009,N_10320,N_13184);
and U15010 (N_15010,N_10365,N_11544);
nand U15011 (N_15011,N_14186,N_12731);
xor U15012 (N_15012,N_13337,N_14798);
nor U15013 (N_15013,N_12996,N_13857);
nand U15014 (N_15014,N_10890,N_10337);
and U15015 (N_15015,N_11721,N_14998);
and U15016 (N_15016,N_10898,N_14674);
nor U15017 (N_15017,N_13458,N_11123);
nand U15018 (N_15018,N_11796,N_10918);
xnor U15019 (N_15019,N_12131,N_13074);
nor U15020 (N_15020,N_13794,N_12237);
nand U15021 (N_15021,N_10116,N_10043);
nor U15022 (N_15022,N_12951,N_13037);
or U15023 (N_15023,N_13599,N_11568);
nand U15024 (N_15024,N_14169,N_10517);
and U15025 (N_15025,N_14468,N_10374);
nor U15026 (N_15026,N_11667,N_14181);
nor U15027 (N_15027,N_12266,N_10091);
and U15028 (N_15028,N_12055,N_10456);
and U15029 (N_15029,N_11697,N_14842);
and U15030 (N_15030,N_10744,N_14005);
nor U15031 (N_15031,N_14087,N_10336);
nand U15032 (N_15032,N_14710,N_12248);
xnor U15033 (N_15033,N_10634,N_10390);
and U15034 (N_15034,N_10798,N_13790);
nand U15035 (N_15035,N_13633,N_10975);
or U15036 (N_15036,N_12197,N_12021);
and U15037 (N_15037,N_11818,N_14292);
and U15038 (N_15038,N_14766,N_13110);
nand U15039 (N_15039,N_10536,N_12574);
nor U15040 (N_15040,N_13832,N_13654);
or U15041 (N_15041,N_12110,N_12019);
or U15042 (N_15042,N_11006,N_10075);
or U15043 (N_15043,N_11399,N_10308);
nand U15044 (N_15044,N_12842,N_11749);
xor U15045 (N_15045,N_11491,N_10197);
nor U15046 (N_15046,N_11541,N_10815);
nor U15047 (N_15047,N_13365,N_10626);
nand U15048 (N_15048,N_13341,N_10196);
nor U15049 (N_15049,N_11695,N_10567);
nand U15050 (N_15050,N_12910,N_10787);
or U15051 (N_15051,N_11404,N_10707);
and U15052 (N_15052,N_11204,N_10375);
xor U15053 (N_15053,N_14273,N_11737);
nor U15054 (N_15054,N_13168,N_13994);
nand U15055 (N_15055,N_10096,N_14801);
or U15056 (N_15056,N_11165,N_10486);
nand U15057 (N_15057,N_14265,N_14979);
nor U15058 (N_15058,N_13896,N_14111);
or U15059 (N_15059,N_11186,N_12453);
or U15060 (N_15060,N_14696,N_12064);
and U15061 (N_15061,N_13714,N_13262);
xnor U15062 (N_15062,N_11470,N_13908);
and U15063 (N_15063,N_10505,N_10441);
xnor U15064 (N_15064,N_12807,N_13787);
or U15065 (N_15065,N_12076,N_11292);
and U15066 (N_15066,N_13851,N_14883);
and U15067 (N_15067,N_13156,N_13313);
and U15068 (N_15068,N_12413,N_11400);
or U15069 (N_15069,N_12551,N_10560);
nand U15070 (N_15070,N_14506,N_10589);
nor U15071 (N_15071,N_10514,N_10912);
nor U15072 (N_15072,N_12457,N_10880);
or U15073 (N_15073,N_14619,N_10957);
nand U15074 (N_15074,N_12588,N_10125);
and U15075 (N_15075,N_14828,N_10235);
and U15076 (N_15076,N_14419,N_11587);
xnor U15077 (N_15077,N_10034,N_11702);
nor U15078 (N_15078,N_11993,N_14253);
or U15079 (N_15079,N_10916,N_14933);
and U15080 (N_15080,N_13981,N_14239);
xor U15081 (N_15081,N_10548,N_11335);
and U15082 (N_15082,N_14759,N_14035);
nor U15083 (N_15083,N_10284,N_13568);
nor U15084 (N_15084,N_12834,N_13311);
and U15085 (N_15085,N_13656,N_10528);
nor U15086 (N_15086,N_10325,N_14874);
or U15087 (N_15087,N_10379,N_14505);
or U15088 (N_15088,N_11874,N_11857);
xnor U15089 (N_15089,N_10478,N_14475);
nand U15090 (N_15090,N_13531,N_14106);
and U15091 (N_15091,N_11090,N_10758);
xor U15092 (N_15092,N_11862,N_12865);
or U15093 (N_15093,N_11246,N_10018);
nor U15094 (N_15094,N_10198,N_14437);
and U15095 (N_15095,N_14852,N_11728);
nand U15096 (N_15096,N_11953,N_12018);
xor U15097 (N_15097,N_14754,N_13558);
xor U15098 (N_15098,N_12729,N_11287);
and U15099 (N_15099,N_13040,N_10129);
or U15100 (N_15100,N_13866,N_12326);
nor U15101 (N_15101,N_10977,N_13067);
or U15102 (N_15102,N_11301,N_10350);
or U15103 (N_15103,N_13248,N_14415);
nor U15104 (N_15104,N_12959,N_14802);
xor U15105 (N_15105,N_14909,N_13758);
nand U15106 (N_15106,N_14302,N_14393);
nand U15107 (N_15107,N_14446,N_11093);
and U15108 (N_15108,N_13527,N_12356);
nor U15109 (N_15109,N_12200,N_13068);
nand U15110 (N_15110,N_13647,N_12709);
or U15111 (N_15111,N_11917,N_13629);
nor U15112 (N_15112,N_13782,N_14136);
or U15113 (N_15113,N_12500,N_14637);
nand U15114 (N_15114,N_12247,N_12930);
and U15115 (N_15115,N_14806,N_11699);
nand U15116 (N_15116,N_14075,N_10780);
and U15117 (N_15117,N_12624,N_11227);
nand U15118 (N_15118,N_11632,N_13487);
or U15119 (N_15119,N_12803,N_13336);
nor U15120 (N_15120,N_10743,N_11440);
nand U15121 (N_15121,N_13906,N_14693);
xor U15122 (N_15122,N_14584,N_13998);
xnor U15123 (N_15123,N_11560,N_11378);
xor U15124 (N_15124,N_10396,N_10387);
and U15125 (N_15125,N_14790,N_10426);
nor U15126 (N_15126,N_11866,N_12404);
nand U15127 (N_15127,N_14433,N_14764);
xnor U15128 (N_15128,N_12726,N_13000);
or U15129 (N_15129,N_11886,N_12875);
xor U15130 (N_15130,N_12094,N_10570);
and U15131 (N_15131,N_13669,N_14250);
nor U15132 (N_15132,N_13569,N_13444);
nor U15133 (N_15133,N_14590,N_11974);
or U15134 (N_15134,N_12394,N_14055);
xnor U15135 (N_15135,N_10158,N_13742);
and U15136 (N_15136,N_10946,N_14886);
nand U15137 (N_15137,N_10013,N_12030);
and U15138 (N_15138,N_10439,N_13975);
and U15139 (N_15139,N_12320,N_13333);
or U15140 (N_15140,N_13206,N_11091);
nor U15141 (N_15141,N_10835,N_14315);
nor U15142 (N_15142,N_13466,N_10940);
or U15143 (N_15143,N_14521,N_13301);
or U15144 (N_15144,N_11778,N_10612);
or U15145 (N_15145,N_12994,N_13355);
nand U15146 (N_15146,N_12324,N_10399);
nor U15147 (N_15147,N_12416,N_10296);
and U15148 (N_15148,N_12614,N_13592);
nor U15149 (N_15149,N_14752,N_11173);
nand U15150 (N_15150,N_10554,N_11213);
nor U15151 (N_15151,N_11466,N_12153);
xor U15152 (N_15152,N_13504,N_10856);
xor U15153 (N_15153,N_12056,N_11014);
nor U15154 (N_15154,N_14684,N_12950);
nand U15155 (N_15155,N_14480,N_14881);
nor U15156 (N_15156,N_11820,N_11623);
nor U15157 (N_15157,N_11340,N_12516);
nor U15158 (N_15158,N_12881,N_13370);
nor U15159 (N_15159,N_10370,N_14227);
nand U15160 (N_15160,N_12621,N_11633);
and U15161 (N_15161,N_11475,N_13549);
and U15162 (N_15162,N_12114,N_12700);
or U15163 (N_15163,N_13800,N_12623);
xnor U15164 (N_15164,N_10925,N_13026);
nor U15165 (N_15165,N_14348,N_12043);
or U15166 (N_15166,N_14533,N_12484);
nor U15167 (N_15167,N_13218,N_14202);
xnor U15168 (N_15168,N_10913,N_13563);
nand U15169 (N_15169,N_14960,N_14918);
and U15170 (N_15170,N_14225,N_10144);
nor U15171 (N_15171,N_10850,N_10683);
nand U15172 (N_15172,N_11498,N_14695);
or U15173 (N_15173,N_10828,N_13401);
nand U15174 (N_15174,N_11952,N_12366);
or U15175 (N_15175,N_11525,N_11407);
nor U15176 (N_15176,N_13543,N_14819);
nor U15177 (N_15177,N_11561,N_13318);
nand U15178 (N_15178,N_10706,N_14527);
nand U15179 (N_15179,N_12308,N_12313);
or U15180 (N_15180,N_11469,N_10045);
nor U15181 (N_15181,N_13115,N_14992);
nand U15182 (N_15182,N_10385,N_12222);
and U15183 (N_15183,N_10924,N_13415);
or U15184 (N_15184,N_13544,N_14681);
nor U15185 (N_15185,N_12282,N_13095);
nor U15186 (N_15186,N_13547,N_12900);
or U15187 (N_15187,N_13047,N_13471);
nor U15188 (N_15188,N_10412,N_12204);
and U15189 (N_15189,N_11085,N_13565);
nor U15190 (N_15190,N_11700,N_12605);
xor U15191 (N_15191,N_13863,N_12735);
nor U15192 (N_15192,N_10165,N_12987);
nand U15193 (N_15193,N_12782,N_13472);
nor U15194 (N_15194,N_13161,N_14373);
or U15195 (N_15195,N_11524,N_13587);
and U15196 (N_15196,N_13798,N_12948);
nor U15197 (N_15197,N_14548,N_11488);
and U15198 (N_15198,N_10113,N_11338);
nor U15199 (N_15199,N_14885,N_10564);
and U15200 (N_15200,N_10061,N_13757);
and U15201 (N_15201,N_10872,N_10493);
nand U15202 (N_15202,N_12963,N_11427);
nor U15203 (N_15203,N_14479,N_10137);
and U15204 (N_15204,N_13071,N_11539);
or U15205 (N_15205,N_10782,N_10998);
nor U15206 (N_15206,N_10696,N_12788);
nor U15207 (N_15207,N_12058,N_11076);
nand U15208 (N_15208,N_11550,N_10413);
or U15209 (N_15209,N_13140,N_11883);
xor U15210 (N_15210,N_10182,N_10215);
or U15211 (N_15211,N_14723,N_10652);
nor U15212 (N_15212,N_10981,N_11356);
nor U15213 (N_15213,N_14103,N_12130);
and U15214 (N_15214,N_14204,N_11757);
nor U15215 (N_15215,N_12396,N_13093);
nand U15216 (N_15216,N_11806,N_13588);
nand U15217 (N_15217,N_13123,N_11562);
nand U15218 (N_15218,N_10476,N_11709);
xnor U15219 (N_15219,N_11433,N_13578);
nand U15220 (N_15220,N_12942,N_10565);
or U15221 (N_15221,N_13993,N_14534);
and U15222 (N_15222,N_11864,N_14875);
and U15223 (N_15223,N_13202,N_13810);
nand U15224 (N_15224,N_13836,N_11104);
or U15225 (N_15225,N_11169,N_10359);
and U15226 (N_15226,N_14335,N_10660);
xnor U15227 (N_15227,N_14755,N_10575);
or U15228 (N_15228,N_12649,N_13303);
or U15229 (N_15229,N_12613,N_13422);
and U15230 (N_15230,N_10057,N_12395);
nor U15231 (N_15231,N_12669,N_11055);
nand U15232 (N_15232,N_13246,N_14525);
or U15233 (N_15233,N_13505,N_13923);
nand U15234 (N_15234,N_10067,N_12111);
nand U15235 (N_15235,N_14203,N_11109);
and U15236 (N_15236,N_12784,N_12220);
nand U15237 (N_15237,N_14474,N_10069);
nand U15238 (N_15238,N_11008,N_10468);
or U15239 (N_15239,N_10952,N_11652);
and U15240 (N_15240,N_11997,N_13723);
nor U15241 (N_15241,N_14063,N_10467);
or U15242 (N_15242,N_14467,N_11659);
nand U15243 (N_15243,N_11431,N_14542);
nand U15244 (N_15244,N_14295,N_10894);
and U15245 (N_15245,N_13024,N_11175);
nand U15246 (N_15246,N_10771,N_10039);
or U15247 (N_15247,N_14568,N_12651);
xor U15248 (N_15248,N_11484,N_11372);
nand U15249 (N_15249,N_13372,N_13885);
and U15250 (N_15250,N_11178,N_13006);
nor U15251 (N_15251,N_12552,N_12117);
nand U15252 (N_15252,N_11973,N_10553);
nand U15253 (N_15253,N_12540,N_12372);
nor U15254 (N_15254,N_14700,N_10557);
and U15255 (N_15255,N_13524,N_14473);
nor U15256 (N_15256,N_10742,N_11374);
or U15257 (N_15257,N_12003,N_10207);
or U15258 (N_15258,N_10122,N_10900);
or U15259 (N_15259,N_13175,N_11596);
nor U15260 (N_15260,N_13295,N_13671);
or U15261 (N_15261,N_13449,N_12607);
nor U15262 (N_15262,N_12302,N_10563);
and U15263 (N_15263,N_12468,N_13771);
or U15264 (N_15264,N_12670,N_11506);
nand U15265 (N_15265,N_10171,N_10990);
xnor U15266 (N_15266,N_13745,N_14043);
nand U15267 (N_15267,N_13883,N_10623);
nor U15268 (N_15268,N_12126,N_11441);
nand U15269 (N_15269,N_12228,N_13595);
or U15270 (N_15270,N_12754,N_13116);
or U15271 (N_15271,N_10275,N_13838);
or U15272 (N_15272,N_13721,N_14914);
and U15273 (N_15273,N_12686,N_12344);
and U15274 (N_15274,N_14299,N_10697);
nor U15275 (N_15275,N_12381,N_14247);
and U15276 (N_15276,N_12305,N_11447);
or U15277 (N_15277,N_12433,N_14685);
xnor U15278 (N_15278,N_13497,N_10710);
nor U15279 (N_15279,N_14785,N_13465);
and U15280 (N_15280,N_10269,N_11305);
or U15281 (N_15281,N_12147,N_12749);
and U15282 (N_15282,N_14839,N_10840);
xnor U15283 (N_15283,N_12217,N_13991);
nor U15284 (N_15284,N_12504,N_13436);
or U15285 (N_15285,N_13682,N_10504);
xor U15286 (N_15286,N_13921,N_11859);
nand U15287 (N_15287,N_13394,N_14236);
nand U15288 (N_15288,N_11226,N_11815);
and U15289 (N_15289,N_10741,N_12045);
or U15290 (N_15290,N_13048,N_11987);
xnor U15291 (N_15291,N_10844,N_11144);
and U15292 (N_15292,N_14466,N_10735);
or U15293 (N_15293,N_13166,N_12891);
nand U15294 (N_15294,N_11369,N_11830);
or U15295 (N_15295,N_14330,N_11795);
or U15296 (N_15296,N_12949,N_10152);
and U15297 (N_15297,N_13747,N_11681);
and U15298 (N_15298,N_13102,N_11120);
nor U15299 (N_15299,N_11328,N_12690);
and U15300 (N_15300,N_13183,N_10721);
and U15301 (N_15301,N_10323,N_13634);
or U15302 (N_15302,N_14276,N_11159);
and U15303 (N_15303,N_13983,N_10958);
nand U15304 (N_15304,N_12838,N_13260);
or U15305 (N_15305,N_13482,N_10666);
nand U15306 (N_15306,N_12233,N_14789);
nand U15307 (N_15307,N_10498,N_11999);
nand U15308 (N_15308,N_12663,N_10988);
nand U15309 (N_15309,N_13240,N_10826);
nand U15310 (N_15310,N_11527,N_12107);
nor U15311 (N_15311,N_11312,N_12447);
nor U15312 (N_15312,N_10531,N_14758);
nor U15313 (N_15313,N_12177,N_13462);
and U15314 (N_15314,N_12420,N_14301);
xor U15315 (N_15315,N_13731,N_11950);
xor U15316 (N_15316,N_11239,N_14425);
or U15317 (N_15317,N_10944,N_10436);
nor U15318 (N_15318,N_10876,N_14104);
xor U15319 (N_15319,N_13045,N_14317);
and U15320 (N_15320,N_14160,N_13391);
or U15321 (N_15321,N_11708,N_11496);
and U15322 (N_15322,N_13580,N_11835);
nor U15323 (N_15323,N_11260,N_10264);
nand U15324 (N_15324,N_11182,N_13608);
and U15325 (N_15325,N_14318,N_10598);
or U15326 (N_15326,N_10962,N_13271);
xnor U15327 (N_15327,N_11478,N_13703);
xor U15328 (N_15328,N_12243,N_12713);
or U15329 (N_15329,N_13502,N_14701);
or U15330 (N_15330,N_14683,N_14650);
nor U15331 (N_15331,N_11210,N_13511);
nor U15332 (N_15332,N_11222,N_14793);
or U15333 (N_15333,N_13384,N_12819);
nand U15334 (N_15334,N_10280,N_11278);
xor U15335 (N_15335,N_10328,N_13638);
nand U15336 (N_15336,N_10725,N_13276);
nand U15337 (N_15337,N_11654,N_14694);
and U15338 (N_15338,N_11131,N_13261);
xor U15339 (N_15339,N_11445,N_14131);
or U15340 (N_15340,N_10321,N_11900);
or U15341 (N_15341,N_10020,N_14632);
and U15342 (N_15342,N_10542,N_10964);
and U15343 (N_15343,N_14528,N_12833);
nor U15344 (N_15344,N_12901,N_13281);
xor U15345 (N_15345,N_11978,N_12898);
xor U15346 (N_15346,N_12231,N_12980);
and U15347 (N_15347,N_10042,N_10012);
xor U15348 (N_15348,N_13591,N_11912);
nand U15349 (N_15349,N_12093,N_10714);
nand U15350 (N_15350,N_14189,N_12345);
xnor U15351 (N_15351,N_10140,N_11664);
nor U15352 (N_15352,N_10146,N_11809);
and U15353 (N_15353,N_10678,N_13488);
or U15354 (N_15354,N_10543,N_14195);
xnor U15355 (N_15355,N_10620,N_10906);
nand U15356 (N_15356,N_13010,N_10812);
and U15357 (N_15357,N_12734,N_12975);
nand U15358 (N_15358,N_14529,N_12645);
nor U15359 (N_15359,N_14155,N_12641);
nand U15360 (N_15360,N_13722,N_14384);
xor U15361 (N_15361,N_10480,N_14690);
and U15362 (N_15362,N_14635,N_11471);
nor U15363 (N_15363,N_10720,N_13196);
xnor U15364 (N_15364,N_12124,N_11313);
nand U15365 (N_15365,N_12268,N_10577);
or U15366 (N_15366,N_11773,N_11208);
nor U15367 (N_15367,N_10041,N_14228);
and U15368 (N_15368,N_10785,N_10407);
and U15369 (N_15369,N_12657,N_11483);
nand U15370 (N_15370,N_14128,N_13913);
xor U15371 (N_15371,N_12772,N_11983);
or U15372 (N_15372,N_12992,N_11281);
nand U15373 (N_15373,N_14064,N_11603);
and U15374 (N_15374,N_13702,N_11710);
and U15375 (N_15375,N_12956,N_11121);
nor U15376 (N_15376,N_14894,N_12099);
or U15377 (N_15377,N_12284,N_12276);
xor U15378 (N_15378,N_13572,N_13508);
or U15379 (N_15379,N_14329,N_10667);
and U15380 (N_15380,N_14321,N_14185);
or U15381 (N_15381,N_12488,N_14198);
and U15382 (N_15382,N_10992,N_11600);
nand U15383 (N_15383,N_10353,N_10929);
or U15384 (N_15384,N_13424,N_14543);
and U15385 (N_15385,N_11873,N_12493);
xnor U15386 (N_15386,N_11095,N_12740);
and U15387 (N_15387,N_14059,N_14497);
nand U15388 (N_15388,N_13817,N_14622);
and U15389 (N_15389,N_13938,N_12102);
nand U15390 (N_15390,N_13766,N_10932);
or U15391 (N_15391,N_10950,N_14919);
nand U15392 (N_15392,N_11489,N_10052);
or U15393 (N_15393,N_11578,N_11412);
or U15394 (N_15394,N_11976,N_11345);
nor U15395 (N_15395,N_10130,N_10283);
nand U15396 (N_15396,N_12499,N_13789);
nand U15397 (N_15397,N_10217,N_11966);
nand U15398 (N_15398,N_14956,N_11609);
or U15399 (N_15399,N_10689,N_11612);
or U15400 (N_15400,N_12636,N_11535);
nand U15401 (N_15401,N_12962,N_13856);
nor U15402 (N_15402,N_14818,N_12523);
and U15403 (N_15403,N_10679,N_12139);
nor U15404 (N_15404,N_12870,N_10600);
or U15405 (N_15405,N_13641,N_11669);
and U15406 (N_15406,N_11396,N_10201);
xor U15407 (N_15407,N_11156,N_12068);
nor U15408 (N_15408,N_13808,N_11885);
and U15409 (N_15409,N_13089,N_12989);
and U15410 (N_15410,N_10873,N_13850);
or U15411 (N_15411,N_13139,N_14478);
nand U15412 (N_15412,N_13957,N_11683);
and U15413 (N_15413,N_12696,N_12584);
nor U15414 (N_15414,N_14296,N_10243);
or U15415 (N_15415,N_13680,N_14322);
nand U15416 (N_15416,N_10286,N_13418);
or U15417 (N_15417,N_13410,N_10066);
and U15418 (N_15418,N_10529,N_10796);
nor U15419 (N_15419,N_14149,N_10764);
nor U15420 (N_15420,N_12839,N_10444);
or U15421 (N_15421,N_13389,N_14021);
nor U15422 (N_15422,N_12351,N_11636);
or U15423 (N_15423,N_13230,N_13953);
and U15424 (N_15424,N_12764,N_11180);
xor U15425 (N_15425,N_11843,N_13007);
and U15426 (N_15426,N_14165,N_11563);
and U15427 (N_15427,N_11254,N_14953);
nor U15428 (N_15428,N_12042,N_11041);
xor U15429 (N_15429,N_11311,N_13978);
nor U15430 (N_15430,N_11429,N_11833);
nor U15431 (N_15431,N_14815,N_10699);
nor U15432 (N_15432,N_11136,N_10266);
nand U15433 (N_15433,N_14341,N_13486);
or U15434 (N_15434,N_13576,N_11291);
or U15435 (N_15435,N_11988,N_11884);
nor U15436 (N_15436,N_14441,N_13090);
and U15437 (N_15437,N_12961,N_12059);
or U15438 (N_15438,N_12186,N_14491);
nor U15439 (N_15439,N_13642,N_13852);
and U15440 (N_15440,N_14938,N_12378);
nand U15441 (N_15441,N_13297,N_11893);
or U15442 (N_15442,N_13092,N_12203);
or U15443 (N_15443,N_12467,N_14609);
nor U15444 (N_15444,N_11847,N_11585);
and U15445 (N_15445,N_12511,N_10040);
nand U15446 (N_15446,N_12312,N_12244);
nand U15447 (N_15447,N_14540,N_11331);
or U15448 (N_15448,N_12022,N_11255);
nand U15449 (N_15449,N_14015,N_11161);
nand U15450 (N_15450,N_10085,N_10842);
nand U15451 (N_15451,N_14680,N_14193);
nor U15452 (N_15452,N_14625,N_12048);
nor U15453 (N_15453,N_14887,N_11420);
and U15454 (N_15454,N_14036,N_10915);
nand U15455 (N_15455,N_12896,N_10378);
or U15456 (N_15456,N_11098,N_12125);
nor U15457 (N_15457,N_12608,N_10586);
and U15458 (N_15458,N_10227,N_14636);
nand U15459 (N_15459,N_13491,N_13227);
and U15460 (N_15460,N_11490,N_14878);
nand U15461 (N_15461,N_12857,N_11696);
xor U15462 (N_15462,N_14237,N_11268);
and U15463 (N_15463,N_14923,N_12520);
and U15464 (N_15464,N_14174,N_10142);
and U15465 (N_15465,N_12791,N_12465);
nand U15466 (N_15466,N_13562,N_11863);
nand U15467 (N_15467,N_14932,N_12423);
nor U15468 (N_15468,N_14371,N_12937);
or U15469 (N_15469,N_10050,N_14518);
nor U15470 (N_15470,N_11867,N_11364);
or U15471 (N_15471,N_12677,N_14688);
and U15472 (N_15472,N_11942,N_14001);
nor U15473 (N_15473,N_10401,N_11515);
nand U15474 (N_15474,N_11051,N_13872);
and U15475 (N_15475,N_13995,N_10884);
and U15476 (N_15476,N_10003,N_11354);
nor U15477 (N_15477,N_10719,N_11367);
xor U15478 (N_15478,N_14066,N_12770);
or U15479 (N_15479,N_14969,N_13507);
or U15480 (N_15480,N_14325,N_12928);
xor U15481 (N_15481,N_12432,N_11125);
and U15482 (N_15482,N_14269,N_14423);
or U15483 (N_15483,N_11235,N_13103);
and U15484 (N_15484,N_10619,N_11230);
nand U15485 (N_15485,N_13478,N_13335);
or U15486 (N_15486,N_10596,N_11054);
or U15487 (N_15487,N_12474,N_14304);
and U15488 (N_15488,N_12884,N_13075);
and U15489 (N_15489,N_13645,N_11564);
or U15490 (N_15490,N_11837,N_10341);
or U15491 (N_15491,N_12814,N_14895);
or U15492 (N_15492,N_13453,N_13083);
nand U15493 (N_15493,N_10416,N_14630);
or U15494 (N_15494,N_12682,N_11639);
nand U15495 (N_15495,N_10819,N_11157);
nand U15496 (N_15496,N_11145,N_14134);
nor U15497 (N_15497,N_14153,N_14487);
nor U15498 (N_15498,N_11238,N_12346);
nor U15499 (N_15499,N_13972,N_12851);
nand U15500 (N_15500,N_14510,N_10597);
nand U15501 (N_15501,N_12831,N_11615);
xor U15502 (N_15502,N_13120,N_11872);
and U15503 (N_15503,N_11456,N_14554);
or U15504 (N_15504,N_10675,N_10099);
or U15505 (N_15505,N_13209,N_12914);
or U15506 (N_15506,N_10588,N_10604);
and U15507 (N_15507,N_12750,N_12001);
nor U15508 (N_15508,N_12066,N_14868);
nor U15509 (N_15509,N_12615,N_10834);
nor U15510 (N_15510,N_14597,N_11823);
or U15511 (N_15511,N_14342,N_12620);
and U15512 (N_15512,N_14392,N_12477);
nand U15513 (N_15513,N_13738,N_14871);
and U15514 (N_15514,N_10354,N_11772);
or U15515 (N_15515,N_12049,N_14337);
xnor U15516 (N_15516,N_14140,N_10222);
or U15517 (N_15517,N_14180,N_11124);
nor U15518 (N_15518,N_10110,N_12417);
or U15519 (N_15519,N_13124,N_14070);
and U15520 (N_15520,N_14970,N_12004);
xor U15521 (N_15521,N_13039,N_13306);
or U15522 (N_15522,N_11870,N_13443);
or U15523 (N_15523,N_14118,N_11185);
nand U15524 (N_15524,N_11207,N_10298);
and U15525 (N_15525,N_10591,N_12370);
nand U15526 (N_15526,N_11651,N_10105);
and U15527 (N_15527,N_14424,N_14613);
and U15528 (N_15528,N_13695,N_11516);
or U15529 (N_15529,N_10822,N_13583);
and U15530 (N_15530,N_13613,N_12585);
and U15531 (N_15531,N_12932,N_11298);
nand U15532 (N_15532,N_13518,N_10102);
nor U15533 (N_15533,N_10271,N_10767);
nand U15534 (N_15534,N_12448,N_12972);
nor U15535 (N_15535,N_11579,N_12733);
xnor U15536 (N_15536,N_14983,N_12011);
and U15537 (N_15537,N_14137,N_13773);
nor U15538 (N_15538,N_14799,N_14499);
nand U15539 (N_15539,N_13383,N_10492);
xnor U15540 (N_15540,N_12269,N_11522);
nor U15541 (N_15541,N_10161,N_13661);
xor U15542 (N_15542,N_12280,N_11330);
nor U15543 (N_15543,N_10968,N_11194);
and U15544 (N_15544,N_11951,N_14737);
nor U15545 (N_15545,N_11723,N_13690);
nand U15546 (N_15546,N_14667,N_14138);
nor U15547 (N_15547,N_12472,N_12539);
nand U15548 (N_15548,N_13250,N_14804);
nor U15549 (N_15549,N_10829,N_14280);
nor U15550 (N_15550,N_13687,N_13428);
nand U15551 (N_15551,N_12554,N_13893);
or U15552 (N_15552,N_13898,N_10705);
nand U15553 (N_15553,N_13490,N_14279);
nor U15554 (N_15554,N_11865,N_11070);
and U15555 (N_15555,N_12919,N_12478);
nand U15556 (N_15556,N_12707,N_10738);
nor U15557 (N_15557,N_12783,N_13445);
and U15558 (N_15558,N_14570,N_13901);
nor U15559 (N_15559,N_12297,N_13996);
xnor U15560 (N_15560,N_12999,N_14746);
and U15561 (N_15561,N_14009,N_11996);
or U15562 (N_15562,N_12306,N_14944);
and U15563 (N_15563,N_12384,N_14549);
nor U15564 (N_15564,N_10332,N_10348);
nand U15565 (N_15565,N_14172,N_14863);
nand U15566 (N_15566,N_12368,N_12410);
nand U15567 (N_15567,N_12033,N_13655);
or U15568 (N_15568,N_13910,N_13429);
or U15569 (N_15569,N_12323,N_11146);
or U15570 (N_15570,N_14774,N_10797);
or U15571 (N_15571,N_11595,N_10510);
nand U15572 (N_15572,N_10527,N_13322);
nor U15573 (N_15573,N_10587,N_10870);
nand U15574 (N_15574,N_13939,N_12333);
nand U15575 (N_15575,N_12113,N_14282);
nor U15576 (N_15576,N_13697,N_10300);
nand U15577 (N_15577,N_13662,N_10392);
or U15578 (N_15578,N_10035,N_11919);
and U15579 (N_15579,N_12051,N_12595);
nor U15580 (N_15580,N_11258,N_10804);
and U15581 (N_15581,N_11743,N_10205);
or U15582 (N_15582,N_14547,N_10595);
and U15583 (N_15583,N_10053,N_11619);
and U15584 (N_15584,N_11129,N_13788);
nand U15585 (N_15585,N_12031,N_11353);
or U15586 (N_15586,N_12242,N_10745);
nor U15587 (N_15587,N_10004,N_13551);
or U15588 (N_15588,N_13698,N_10212);
or U15589 (N_15589,N_13216,N_12568);
nand U15590 (N_15590,N_10766,N_11554);
nand U15591 (N_15591,N_14776,N_12328);
nand U15592 (N_15592,N_11922,N_14130);
or U15593 (N_15593,N_12918,N_10326);
and U15594 (N_15594,N_10814,N_14713);
nand U15595 (N_15595,N_14052,N_14283);
and U15596 (N_15596,N_10827,N_12893);
or U15597 (N_15597,N_13498,N_14906);
nand U15598 (N_15598,N_14810,N_13288);
nor U15599 (N_15599,N_11388,N_14663);
nand U15600 (N_15600,N_10083,N_11137);
xor U15601 (N_15601,N_12562,N_13275);
nand U15602 (N_15602,N_13719,N_12255);
xor U15603 (N_15603,N_11703,N_11622);
or U15604 (N_15604,N_10724,N_13078);
or U15605 (N_15605,N_11058,N_14911);
or U15606 (N_15606,N_13686,N_13559);
and U15607 (N_15607,N_14360,N_13734);
nand U15608 (N_15608,N_12872,N_11798);
or U15609 (N_15609,N_10005,N_10036);
or U15610 (N_15610,N_10693,N_13830);
nor U15611 (N_15611,N_14205,N_13426);
and U15612 (N_15612,N_13631,N_11450);
xor U15613 (N_15613,N_14083,N_13512);
nor U15614 (N_15614,N_12260,N_11994);
and U15615 (N_15615,N_11678,N_11326);
nor U15616 (N_15616,N_10629,N_14612);
and U15617 (N_15617,N_13709,N_12721);
and U15618 (N_15618,N_12024,N_12506);
xor U15619 (N_15619,N_12142,N_14175);
nand U15620 (N_15620,N_11393,N_12032);
xor U15621 (N_15621,N_14712,N_14004);
nor U15622 (N_15622,N_10226,N_14346);
or U15623 (N_15623,N_11075,N_10680);
or U15624 (N_15624,N_14472,N_11009);
nor U15625 (N_15625,N_12192,N_13154);
nand U15626 (N_15626,N_14387,N_12874);
nor U15627 (N_15627,N_12451,N_10806);
and U15628 (N_15628,N_12548,N_10511);
and U15629 (N_15629,N_13736,N_14589);
xor U15630 (N_15630,N_13653,N_10657);
and U15631 (N_15631,N_12671,N_13287);
or U15632 (N_15632,N_12737,N_12081);
nor U15633 (N_15633,N_14638,N_11944);
nor U15634 (N_15634,N_10233,N_13345);
nor U15635 (N_15635,N_13891,N_11567);
nand U15636 (N_15636,N_13769,N_10824);
nor U15637 (N_15637,N_12867,N_14076);
or U15638 (N_15638,N_10791,N_11959);
or U15639 (N_15639,N_11897,N_13413);
nor U15640 (N_15640,N_13151,N_14270);
nor U15641 (N_15641,N_12611,N_14560);
nand U15642 (N_15642,N_12424,N_14320);
nand U15643 (N_15643,N_10109,N_10853);
nor U15644 (N_15644,N_11279,N_13265);
nand U15645 (N_15645,N_14879,N_14767);
xnor U15646 (N_15646,N_10241,N_13762);
or U15647 (N_15647,N_11546,N_13622);
nand U15648 (N_15648,N_11333,N_14892);
or U15649 (N_15649,N_14224,N_11673);
nand U15650 (N_15650,N_11716,N_13146);
nor U15651 (N_15651,N_10362,N_10103);
and U15652 (N_15652,N_11474,N_13214);
nor U15653 (N_15653,N_14047,N_13464);
nand U15654 (N_15654,N_11134,N_11106);
or U15655 (N_15655,N_14272,N_12067);
nand U15656 (N_15656,N_12541,N_11571);
nor U15657 (N_15657,N_13877,N_13052);
nand U15658 (N_15658,N_12062,N_10369);
or U15659 (N_15659,N_14846,N_12070);
nand U15660 (N_15660,N_11626,N_12905);
and U15661 (N_15661,N_10624,N_13085);
and U15662 (N_15662,N_10263,N_12245);
nand U15663 (N_15663,N_10994,N_13548);
xnor U15664 (N_15664,N_13793,N_13446);
and U15665 (N_15665,N_11671,N_14297);
nand U15666 (N_15666,N_13887,N_13658);
nand U15667 (N_15667,N_14856,N_11979);
nor U15668 (N_15668,N_14380,N_13648);
xor U15669 (N_15669,N_13849,N_14388);
nand U15670 (N_15670,N_11302,N_14105);
nor U15671 (N_15671,N_14401,N_11824);
nor U15672 (N_15672,N_11602,N_12489);
and U15673 (N_15673,N_13679,N_14686);
nand U15674 (N_15674,N_14691,N_11435);
nor U15675 (N_15675,N_12643,N_11143);
and U15676 (N_15676,N_11437,N_10482);
nand U15677 (N_15677,N_14069,N_10613);
or U15678 (N_15678,N_14305,N_12145);
nor U15679 (N_15679,N_11586,N_11628);
and U15680 (N_15680,N_13603,N_12039);
nand U15681 (N_15681,N_14903,N_11637);
nand U15682 (N_15682,N_13784,N_12570);
nand U15683 (N_15683,N_10418,N_11034);
nor U15684 (N_15684,N_10891,N_12763);
nand U15685 (N_15685,N_12510,N_12743);
nor U15686 (N_15686,N_11380,N_14459);
nor U15687 (N_15687,N_11370,N_13070);
nor U15688 (N_15688,N_12213,N_11196);
nand U15689 (N_15689,N_10376,N_14967);
nor U15690 (N_15690,N_14857,N_11599);
or U15691 (N_15691,N_14882,N_10162);
nor U15692 (N_15692,N_12252,N_10843);
xor U15693 (N_15693,N_10866,N_11386);
and U15694 (N_15694,N_13025,N_12409);
nand U15695 (N_15695,N_11443,N_10219);
nor U15696 (N_15696,N_14800,N_11690);
nand U15697 (N_15697,N_13495,N_13468);
xor U15698 (N_15698,N_14908,N_10360);
nor U15699 (N_15699,N_10545,N_13777);
xor U15700 (N_15700,N_11905,N_11842);
or U15701 (N_15701,N_14937,N_11839);
or U15702 (N_15702,N_10461,N_12089);
nand U15703 (N_15703,N_14026,N_13134);
nand U15704 (N_15704,N_14351,N_13621);
or U15705 (N_15705,N_12446,N_11223);
nor U15706 (N_15706,N_13949,N_10127);
xnor U15707 (N_15707,N_12199,N_13894);
nand U15708 (N_15708,N_12702,N_13253);
nor U15709 (N_15709,N_10234,N_10000);
nor U15710 (N_15710,N_11368,N_13959);
and U15711 (N_15711,N_10867,N_13827);
nand U15712 (N_15712,N_13280,N_12586);
nand U15713 (N_15713,N_14948,N_11765);
and U15714 (N_15714,N_14725,N_12128);
or U15715 (N_15715,N_13735,N_10753);
or U15716 (N_15716,N_11739,N_14074);
and U15717 (N_15717,N_14234,N_14794);
nor U15718 (N_15718,N_13833,N_12286);
and U15719 (N_15719,N_14849,N_12985);
and U15720 (N_15720,N_11547,N_10400);
nor U15721 (N_15721,N_11980,N_12503);
and U15722 (N_15722,N_14571,N_13061);
nor U15723 (N_15723,N_13598,N_11566);
nand U15724 (N_15724,N_14999,N_13169);
or U15725 (N_15725,N_10863,N_13865);
nand U15726 (N_15726,N_14017,N_13257);
nand U15727 (N_15727,N_12134,N_12096);
and U15728 (N_15728,N_14158,N_11191);
nand U15729 (N_15729,N_12382,N_13188);
nor U15730 (N_15730,N_12227,N_10421);
nor U15731 (N_15731,N_13448,N_11214);
and U15732 (N_15732,N_11409,N_14408);
and U15733 (N_15733,N_14343,N_14913);
xnor U15734 (N_15734,N_13831,N_11903);
and U15735 (N_15735,N_11881,N_12388);
or U15736 (N_15736,N_14706,N_14604);
and U15737 (N_15737,N_14383,N_13792);
xnor U15738 (N_15738,N_13605,N_14094);
or U15739 (N_15739,N_13617,N_11663);
nor U15740 (N_15740,N_14258,N_13909);
nand U15741 (N_15741,N_10763,N_10897);
and U15742 (N_15742,N_11860,N_11221);
and U15743 (N_15743,N_12978,N_13900);
nor U15744 (N_15744,N_10572,N_12148);
nand U15745 (N_15745,N_14010,N_12841);
nor U15746 (N_15746,N_11117,N_13290);
nand U15747 (N_15747,N_13924,N_11249);
and U15748 (N_15748,N_12941,N_14699);
and U15749 (N_15749,N_13944,N_11738);
and U15750 (N_15750,N_11896,N_12798);
nor U15751 (N_15751,N_12494,N_13828);
nor U15752 (N_15752,N_11295,N_11391);
xor U15753 (N_15753,N_10701,N_14440);
or U15754 (N_15754,N_14455,N_14575);
nand U15755 (N_15755,N_10593,N_14217);
or U15756 (N_15756,N_12778,N_14194);
or U15757 (N_15757,N_11115,N_14141);
and U15758 (N_15758,N_11029,N_13752);
nor U15759 (N_15759,N_11421,N_11479);
and U15760 (N_15760,N_10658,N_14773);
and U15761 (N_15761,N_14422,N_13097);
and U15762 (N_15762,N_12576,N_14867);
xor U15763 (N_15763,N_10849,N_10164);
nor U15764 (N_15764,N_10631,N_12164);
xnor U15765 (N_15765,N_12979,N_10908);
and U15766 (N_15766,N_12973,N_12983);
nand U15767 (N_15767,N_11620,N_11211);
nor U15768 (N_15768,N_10008,N_11376);
nand U15769 (N_15769,N_13876,N_11608);
nor U15770 (N_15770,N_11151,N_10537);
nand U15771 (N_15771,N_12211,N_10709);
and U15772 (N_15772,N_10355,N_12512);
and U15773 (N_15773,N_13594,N_10513);
nor U15774 (N_15774,N_11819,N_14756);
nand U15775 (N_15775,N_12355,N_10015);
or U15776 (N_15776,N_10185,N_11969);
and U15777 (N_15777,N_12256,N_10917);
nand U15778 (N_15778,N_13726,N_10055);
or U15779 (N_15779,N_13767,N_14935);
nand U15780 (N_15780,N_12761,N_14257);
and U15781 (N_15781,N_14655,N_12086);
xor U15782 (N_15782,N_11110,N_13739);
and U15783 (N_15783,N_13612,N_11152);
and U15784 (N_15784,N_14537,N_13038);
nand U15785 (N_15785,N_13423,N_14053);
nor U15786 (N_15786,N_13266,N_10154);
xor U15787 (N_15787,N_10088,N_12358);
and U15788 (N_15788,N_11731,N_13969);
xor U15789 (N_15789,N_10966,N_11717);
nand U15790 (N_15790,N_10726,N_10892);
and U15791 (N_15791,N_12325,N_14985);
or U15792 (N_15792,N_13904,N_14670);
nand U15793 (N_15793,N_13082,N_13441);
and U15794 (N_15794,N_12082,N_11844);
nand U15795 (N_15795,N_11149,N_14729);
nor U15796 (N_15796,N_14662,N_10547);
and U15797 (N_15797,N_10868,N_10752);
or U15798 (N_15798,N_10691,N_14552);
nand U15799 (N_15799,N_13207,N_10100);
nor U15800 (N_15800,N_12542,N_14741);
xnor U15801 (N_15801,N_10106,N_10265);
or U15802 (N_15802,N_14620,N_10831);
and U15803 (N_15803,N_14492,N_13812);
and U15804 (N_15804,N_11377,N_13172);
xor U15805 (N_15805,N_12466,N_12261);
and U15806 (N_15806,N_14353,N_12112);
or U15807 (N_15807,N_12040,N_10192);
and U15808 (N_15808,N_11583,N_13732);
and U15809 (N_15809,N_14097,N_11706);
nand U15810 (N_15810,N_11790,N_13254);
nand U15811 (N_15811,N_12887,N_14145);
or U15812 (N_15812,N_13017,N_12505);
and U15813 (N_15813,N_13925,N_11614);
or U15814 (N_15814,N_10295,N_14458);
xor U15815 (N_15815,N_11444,N_13606);
or U15816 (N_15816,N_10751,N_10452);
xnor U15817 (N_15817,N_12687,N_11111);
nor U15818 (N_15818,N_10685,N_12387);
xor U15819 (N_15819,N_14949,N_13571);
and U15820 (N_15820,N_12861,N_10524);
nand U15821 (N_15821,N_11589,N_10420);
and U15822 (N_15822,N_12373,N_14200);
or U15823 (N_15823,N_14934,N_10779);
and U15824 (N_15824,N_13197,N_14223);
xnor U15825 (N_15825,N_13225,N_14024);
or U15826 (N_15826,N_13853,N_10449);
nor U15827 (N_15827,N_10703,N_10647);
and U15828 (N_15828,N_12953,N_13982);
and U15829 (N_15829,N_13348,N_11655);
nor U15830 (N_15830,N_14545,N_10474);
or U15831 (N_15831,N_13432,N_12846);
nor U15832 (N_15832,N_14816,N_13241);
xnor U15833 (N_15833,N_12514,N_14557);
or U15834 (N_15834,N_14486,N_11855);
nand U15835 (N_15835,N_14738,N_11200);
or U15836 (N_15836,N_13870,N_11220);
nor U15837 (N_15837,N_10971,N_14796);
nor U15838 (N_15838,N_14157,N_11635);
nand U15839 (N_15839,N_13203,N_13343);
and U15840 (N_15840,N_10084,N_11879);
nor U15841 (N_15841,N_13004,N_11390);
xnor U15842 (N_15842,N_10475,N_14287);
and U15843 (N_15843,N_14000,N_11318);
and U15844 (N_15844,N_12794,N_12795);
nand U15845 (N_15845,N_13258,N_11403);
nand U15846 (N_15846,N_10821,N_11346);
and U15847 (N_15847,N_11582,N_10139);
nand U15848 (N_15848,N_14290,N_11748);
nor U15849 (N_15849,N_10718,N_12906);
nand U15850 (N_15850,N_10902,N_10969);
or U15851 (N_15851,N_13963,N_12716);
or U15852 (N_15852,N_12296,N_13778);
nor U15853 (N_15853,N_10509,N_14212);
nand U15854 (N_15854,N_12640,N_10611);
or U15855 (N_15855,N_11718,N_11943);
or U15856 (N_15856,N_10087,N_12801);
and U15857 (N_15857,N_10342,N_10089);
nand U15858 (N_15858,N_13164,N_13226);
nand U15859 (N_15859,N_12426,N_10193);
or U15860 (N_15860,N_12158,N_14962);
nor U15861 (N_15861,N_11518,N_10082);
and U15862 (N_15862,N_11341,N_12832);
nor U15863 (N_15863,N_14435,N_11216);
and U15864 (N_15864,N_13427,N_14566);
or U15865 (N_15865,N_13117,N_12224);
nor U15866 (N_15866,N_10315,N_11457);
and U15867 (N_15867,N_13219,N_13050);
nand U15868 (N_15868,N_12087,N_13920);
nor U15869 (N_15869,N_10566,N_11895);
and U15870 (N_15870,N_12769,N_14262);
nand U15871 (N_15871,N_10970,N_14954);
nand U15872 (N_15872,N_13421,N_10221);
or U15873 (N_15873,N_12728,N_10017);
and U15874 (N_15874,N_14556,N_11365);
nor U15875 (N_15875,N_12273,N_14661);
nor U15876 (N_15876,N_10389,N_11666);
or U15877 (N_15877,N_13905,N_11711);
or U15878 (N_15878,N_13347,N_11607);
or U15879 (N_15879,N_13077,N_13515);
or U15880 (N_15880,N_10851,N_13317);
or U15881 (N_15881,N_12597,N_10367);
and U15882 (N_15882,N_10259,N_11929);
nand U15883 (N_15883,N_11397,N_13846);
and U15884 (N_15884,N_12265,N_11043);
nor U15885 (N_15885,N_12405,N_14271);
and U15886 (N_15886,N_12108,N_11876);
and U15887 (N_15887,N_13111,N_11359);
or U15888 (N_15888,N_14166,N_10188);
nand U15889 (N_15889,N_14993,N_11551);
or U15890 (N_15890,N_14964,N_10244);
and U15891 (N_15891,N_13382,N_11494);
or U15892 (N_15892,N_14942,N_13269);
or U15893 (N_15893,N_14940,N_12712);
nand U15894 (N_15894,N_10216,N_12698);
and U15895 (N_15895,N_13664,N_11851);
nor U15896 (N_15896,N_11304,N_11155);
nor U15897 (N_15897,N_13834,N_14600);
or U15898 (N_15898,N_14078,N_10002);
or U15899 (N_15899,N_14012,N_11428);
and U15900 (N_15900,N_12618,N_12491);
nand U15901 (N_15901,N_12817,N_11362);
nor U15902 (N_15902,N_13774,N_14901);
or U15903 (N_15903,N_12027,N_13014);
and U15904 (N_15904,N_14994,N_10672);
xor U15905 (N_15905,N_14788,N_13016);
nor U15906 (N_15906,N_13032,N_11657);
xor U15907 (N_15907,N_10145,N_14671);
and U15908 (N_15908,N_11116,N_12281);
nor U15909 (N_15909,N_11910,N_11598);
nor U15910 (N_15910,N_11375,N_13167);
nand U15911 (N_15911,N_13727,N_11529);
nand U15912 (N_15912,N_13574,N_13087);
nand U15913 (N_15913,N_11010,N_10024);
xor U15914 (N_15914,N_10191,N_11102);
or U15915 (N_15915,N_13278,N_11073);
nor U15916 (N_15916,N_13399,N_14829);
or U15917 (N_15917,N_14394,N_13779);
or U15918 (N_15918,N_14328,N_10772);
nor U15919 (N_15919,N_14838,N_14958);
and U15920 (N_15920,N_12479,N_10788);
nand U15921 (N_15921,N_11459,N_10261);
or U15922 (N_15922,N_10424,N_13970);
nand U15923 (N_15923,N_14925,N_11468);
nand U15924 (N_15924,N_14439,N_13400);
or U15925 (N_15925,N_10538,N_12666);
or U15926 (N_15926,N_11510,N_14432);
nand U15927 (N_15927,N_13509,N_14098);
nor U15928 (N_15928,N_13520,N_12079);
and U15929 (N_15929,N_13375,N_10803);
or U15930 (N_15930,N_12440,N_13955);
nor U15931 (N_15931,N_12871,N_14574);
nand U15932 (N_15932,N_14657,N_10487);
xnor U15933 (N_15933,N_12780,N_11840);
nand U15934 (N_15934,N_14602,N_11972);
or U15935 (N_15935,N_14143,N_10526);
nor U15936 (N_15936,N_12673,N_12779);
or U15937 (N_15937,N_13326,N_11691);
nor U15938 (N_15938,N_10458,N_14643);
and U15939 (N_15939,N_14761,N_10433);
or U15940 (N_15940,N_14168,N_13820);
xnor U15941 (N_15941,N_14233,N_12715);
or U15942 (N_15942,N_14711,N_10608);
xor U15943 (N_15943,N_12216,N_13191);
nand U15944 (N_15944,N_11565,N_14567);
and U15945 (N_15945,N_10147,N_13525);
or U15946 (N_15946,N_11193,N_10073);
or U15947 (N_15947,N_12701,N_13080);
nor U15948 (N_15948,N_13869,N_12210);
and U15949 (N_15949,N_13430,N_11786);
nor U15950 (N_15950,N_14708,N_10989);
xor U15951 (N_15951,N_11925,N_10584);
nor U15952 (N_15952,N_12830,N_13056);
nor U15953 (N_15953,N_12547,N_11753);
or U15954 (N_15954,N_12338,N_10568);
and U15955 (N_15955,N_11661,N_13456);
nand U15956 (N_15956,N_14079,N_13473);
and U15957 (N_15957,N_11181,N_12283);
and U15958 (N_15958,N_10669,N_10578);
nand U15959 (N_15959,N_13084,N_10179);
or U15960 (N_15960,N_10304,N_10617);
or U15961 (N_15961,N_13296,N_10322);
nor U15962 (N_15962,N_10515,N_10190);
or U15963 (N_15963,N_10762,N_14489);
nand U15964 (N_15964,N_12853,N_13816);
nor U15965 (N_15965,N_10953,N_10134);
and U15966 (N_15966,N_12679,N_10781);
or U15967 (N_15967,N_14581,N_13460);
or U15968 (N_15968,N_10157,N_11088);
nand U15969 (N_15969,N_11742,N_13021);
and U15970 (N_15970,N_11831,N_14062);
nand U15971 (N_15971,N_13228,N_13122);
or U15972 (N_15972,N_13023,N_10931);
nand U15973 (N_15973,N_14411,N_12025);
nor U15974 (N_15974,N_11788,N_12307);
xor U15975 (N_15975,N_14434,N_10654);
nor U15976 (N_15976,N_12202,N_13210);
and U15977 (N_15977,N_13712,N_13187);
nor U15978 (N_15978,N_14354,N_10737);
nand U15979 (N_15979,N_13159,N_14209);
or U15980 (N_15980,N_14382,N_10951);
or U15981 (N_15981,N_12159,N_14679);
nand U15982 (N_15982,N_12418,N_12376);
or U15983 (N_15983,N_10408,N_14583);
nand U15984 (N_15984,N_12289,N_14263);
nand U15985 (N_15985,N_14349,N_13404);
nor U15986 (N_15986,N_10761,N_12431);
nand U15987 (N_15987,N_11768,N_11273);
nand U15988 (N_15988,N_14500,N_12844);
nor U15989 (N_15989,N_12873,N_10616);
nand U15990 (N_15990,N_12492,N_13932);
nand U15991 (N_15991,N_14254,N_13799);
nand U15992 (N_15992,N_12522,N_10255);
or U15993 (N_15993,N_14631,N_11068);
and U15994 (N_15994,N_13395,N_11956);
nand U15995 (N_15995,N_12925,N_14235);
nor U15996 (N_15996,N_13935,N_12929);
or U15997 (N_15997,N_14081,N_12741);
or U15998 (N_15998,N_14634,N_13890);
or U15999 (N_15999,N_12993,N_13818);
or U16000 (N_16000,N_13435,N_13358);
and U16001 (N_16001,N_10274,N_10533);
or U16002 (N_16002,N_12184,N_11446);
nand U16003 (N_16003,N_12469,N_10676);
or U16004 (N_16004,N_13967,N_11458);
or U16005 (N_16005,N_10544,N_10463);
and U16006 (N_16006,N_12984,N_13340);
xor U16007 (N_16007,N_12829,N_13554);
or U16008 (N_16008,N_11940,N_13055);
or U16009 (N_16009,N_11247,N_11746);
xor U16010 (N_16010,N_13157,N_14678);
nand U16011 (N_16011,N_11036,N_11549);
and U16012 (N_16012,N_11958,N_11924);
nand U16013 (N_16013,N_10793,N_11224);
or U16014 (N_16014,N_11688,N_13911);
or U16015 (N_16015,N_10128,N_10333);
xor U16016 (N_16016,N_13439,N_14184);
or U16017 (N_16017,N_13353,N_14872);
and U16018 (N_16018,N_10502,N_14082);
or U16019 (N_16019,N_13755,N_13649);
nand U16020 (N_16020,N_11141,N_13194);
nand U16021 (N_16021,N_12835,N_11715);
nor U16022 (N_16022,N_12742,N_13378);
or U16023 (N_16023,N_14398,N_11770);
and U16024 (N_16024,N_10756,N_14811);
xnor U16025 (N_16025,N_14256,N_10895);
nand U16026 (N_16026,N_11045,N_12101);
nand U16027 (N_16027,N_10535,N_14482);
and U16028 (N_16028,N_12169,N_11913);
and U16029 (N_16029,N_13454,N_14451);
nor U16030 (N_16030,N_13079,N_14390);
nor U16031 (N_16031,N_13030,N_14285);
nand U16032 (N_16032,N_12982,N_10344);
nand U16033 (N_16033,N_12654,N_14014);
nor U16034 (N_16034,N_11321,N_13284);
nor U16035 (N_16035,N_11096,N_11781);
and U16036 (N_16036,N_12012,N_11570);
and U16037 (N_16037,N_10671,N_13871);
or U16038 (N_16038,N_14485,N_14211);
nand U16039 (N_16039,N_13121,N_11923);
nand U16040 (N_16040,N_14190,N_12892);
or U16041 (N_16041,N_12073,N_12797);
and U16042 (N_16042,N_10942,N_13663);
and U16043 (N_16043,N_13344,N_11004);
and U16044 (N_16044,N_12882,N_11303);
nand U16045 (N_16045,N_10311,N_13501);
and U16046 (N_16046,N_14539,N_13043);
nor U16047 (N_16047,N_14073,N_12777);
nand U16048 (N_16048,N_14006,N_10610);
or U16049 (N_16049,N_14436,N_10251);
nor U16050 (N_16050,N_13628,N_14444);
or U16051 (N_16051,N_10080,N_13874);
or U16052 (N_16052,N_14361,N_11170);
nor U16053 (N_16053,N_14456,N_13614);
or U16054 (N_16054,N_13903,N_14988);
or U16055 (N_16055,N_12804,N_13535);
nor U16056 (N_16056,N_11856,N_10877);
or U16057 (N_16057,N_11858,N_10605);
nand U16058 (N_16058,N_13980,N_14862);
xor U16059 (N_16059,N_12863,N_13630);
xor U16060 (N_16060,N_13069,N_10278);
nand U16061 (N_16061,N_10607,N_13285);
or U16062 (N_16062,N_12434,N_14018);
nand U16063 (N_16063,N_12078,N_11118);
nor U16064 (N_16064,N_10580,N_14880);
or U16065 (N_16065,N_12894,N_12363);
xnor U16066 (N_16066,N_13153,N_11849);
nand U16067 (N_16067,N_11520,N_11947);
nand U16068 (N_16068,N_12530,N_14504);
nor U16069 (N_16069,N_14139,N_12098);
or U16070 (N_16070,N_10151,N_12852);
and U16071 (N_16071,N_12334,N_13922);
nand U16072 (N_16072,N_11028,N_14413);
and U16073 (N_16073,N_13182,N_11360);
nand U16074 (N_16074,N_12219,N_13546);
or U16075 (N_16075,N_12944,N_12519);
nor U16076 (N_16076,N_14963,N_13066);
nor U16077 (N_16077,N_14102,N_13968);
nor U16078 (N_16078,N_13539,N_10051);
nor U16079 (N_16079,N_11735,N_13530);
or U16080 (N_16080,N_14668,N_14623);
nand U16081 (N_16081,N_14833,N_13802);
and U16082 (N_16082,N_12866,N_10339);
and U16083 (N_16083,N_12013,N_10628);
and U16084 (N_16084,N_12845,N_13596);
nor U16085 (N_16085,N_12538,N_12253);
and U16086 (N_16086,N_11060,N_12391);
nor U16087 (N_16087,N_10974,N_12719);
or U16088 (N_16088,N_10180,N_12357);
nand U16089 (N_16089,N_10414,N_13756);
nor U16090 (N_16090,N_12196,N_11653);
nand U16091 (N_16091,N_14676,N_12746);
and U16092 (N_16092,N_14007,N_11613);
and U16093 (N_16093,N_13141,N_12425);
nand U16094 (N_16094,N_13319,N_10921);
nor U16095 (N_16095,N_14660,N_14417);
and U16096 (N_16096,N_12934,N_12524);
nand U16097 (N_16097,N_14391,N_10343);
and U16098 (N_16098,N_13496,N_13749);
or U16099 (N_16099,N_10327,N_10852);
nand U16100 (N_16100,N_11285,N_12725);
or U16101 (N_16101,N_11701,N_10288);
xnor U16102 (N_16102,N_12668,N_14171);
and U16103 (N_16103,N_14517,N_10976);
nand U16104 (N_16104,N_13211,N_14587);
nand U16105 (N_16105,N_14812,N_11071);
xor U16106 (N_16106,N_12091,N_14641);
nand U16107 (N_16107,N_10576,N_10603);
or U16108 (N_16108,N_13627,N_12974);
nor U16109 (N_16109,N_14364,N_12183);
or U16110 (N_16110,N_14431,N_12816);
xnor U16111 (N_16111,N_10027,N_11113);
nand U16112 (N_16112,N_10911,N_10176);
and U16113 (N_16113,N_12229,N_14976);
nor U16114 (N_16114,N_10945,N_12566);
and U16115 (N_16115,N_14450,N_11430);
xor U16116 (N_16116,N_13740,N_11887);
xor U16117 (N_16117,N_12811,N_10434);
or U16118 (N_16118,N_10777,N_14363);
or U16119 (N_16119,N_11119,N_12257);
and U16120 (N_16120,N_10077,N_10717);
and U16121 (N_16121,N_11741,N_11556);
or U16122 (N_16122,N_11347,N_14721);
nand U16123 (N_16123,N_13291,N_10111);
nor U16124 (N_16124,N_14161,N_13476);
nor U16125 (N_16125,N_13881,N_12069);
and U16126 (N_16126,N_10809,N_13540);
and U16127 (N_16127,N_12249,N_13705);
nand U16128 (N_16128,N_13943,N_12902);
nand U16129 (N_16129,N_11031,N_14718);
nand U16130 (N_16130,N_10178,N_13867);
nor U16131 (N_16131,N_13493,N_12294);
and U16132 (N_16132,N_12856,N_13352);
xor U16133 (N_16133,N_10409,N_10996);
nor U16134 (N_16134,N_10117,N_12888);
and U16135 (N_16135,N_13693,N_11945);
xnor U16136 (N_16136,N_12459,N_12470);
xnor U16137 (N_16137,N_12143,N_13483);
or U16138 (N_16138,N_13065,N_11593);
and U16139 (N_16139,N_11827,N_11005);
nor U16140 (N_16140,N_12427,N_14260);
and U16141 (N_16141,N_11500,N_14460);
and U16142 (N_16142,N_13760,N_13713);
and U16143 (N_16143,N_10324,N_14598);
nor U16144 (N_16144,N_11920,N_12336);
nand U16145 (N_16145,N_11130,N_10285);
nand U16146 (N_16146,N_10183,N_11288);
or U16147 (N_16147,N_14199,N_13013);
xor U16148 (N_16148,N_10464,N_12072);
nand U16149 (N_16149,N_13864,N_12806);
nand U16150 (N_16150,N_11898,N_11240);
and U16151 (N_16151,N_14763,N_12010);
or U16152 (N_16152,N_11344,N_12293);
or U16153 (N_16153,N_11704,N_13155);
nor U16154 (N_16154,N_11782,N_14427);
nor U16155 (N_16155,N_11452,N_10023);
and U16156 (N_16156,N_12337,N_10708);
and U16157 (N_16157,N_12515,N_11206);
or U16158 (N_16158,N_12342,N_10163);
nand U16159 (N_16159,N_10279,N_11992);
nand U16160 (N_16160,N_12174,N_10747);
nand U16161 (N_16161,N_10247,N_14822);
and U16162 (N_16162,N_13744,N_14936);
nor U16163 (N_16163,N_13717,N_10448);
and U16164 (N_16164,N_14192,N_14926);
and U16165 (N_16165,N_14220,N_11531);
nand U16166 (N_16166,N_11499,N_13051);
and U16167 (N_16167,N_12365,N_12267);
nand U16168 (N_16168,N_12582,N_11415);
or U16169 (N_16169,N_14293,N_14559);
and U16170 (N_16170,N_13575,N_10858);
nor U16171 (N_16171,N_14208,N_12115);
xor U16172 (N_16172,N_14042,N_10386);
and U16173 (N_16173,N_13708,N_14369);
or U16174 (N_16174,N_14978,N_13561);
nor U16175 (N_16175,N_11792,N_11337);
nand U16176 (N_16176,N_11939,N_11007);
nor U16177 (N_16177,N_10282,N_11686);
or U16178 (N_16178,N_11852,N_10290);
nand U16179 (N_16179,N_12745,N_14350);
or U16180 (N_16180,N_10559,N_13309);
and U16181 (N_16181,N_12037,N_11538);
or U16182 (N_16182,N_12343,N_11315);
xor U16183 (N_16183,N_14781,N_12931);
or U16184 (N_16184,N_12710,N_13623);
xor U16185 (N_16185,N_14569,N_11630);
or U16186 (N_16186,N_10398,N_14704);
and U16187 (N_16187,N_14331,N_11713);
nor U16188 (N_16188,N_13147,N_10358);
or U16189 (N_16189,N_10046,N_10431);
or U16190 (N_16190,N_13474,N_11283);
or U16191 (N_16191,N_11543,N_12521);
nor U16192 (N_16192,N_10189,N_12238);
nor U16193 (N_16193,N_13683,N_11675);
or U16194 (N_16194,N_13710,N_10388);
nand U16195 (N_16195,N_13104,N_10483);
or U16196 (N_16196,N_10313,N_10428);
nor U16197 (N_16197,N_13243,N_13582);
xnor U16198 (N_16198,N_12544,N_10984);
and U16199 (N_16199,N_14897,N_12303);
nor U16200 (N_16200,N_13447,N_14240);
and U16201 (N_16201,N_11163,N_12390);
or U16202 (N_16202,N_14267,N_12160);
nor U16203 (N_16203,N_12658,N_11714);
nand U16204 (N_16204,N_12454,N_13463);
or U16205 (N_16205,N_11552,N_11928);
nor U16206 (N_16206,N_11660,N_10466);
and U16207 (N_16207,N_11899,N_14779);
and U16208 (N_16208,N_13620,N_10453);
nand U16209 (N_16209,N_12714,N_12627);
nor U16210 (N_16210,N_10769,N_10270);
or U16211 (N_16211,N_11371,N_12912);
or U16212 (N_16212,N_14553,N_10347);
and U16213 (N_16213,N_10340,N_12622);
xnor U16214 (N_16214,N_14022,N_13215);
nor U16215 (N_16215,N_14490,N_14621);
and U16216 (N_16216,N_13914,N_14243);
and U16217 (N_16217,N_13163,N_12647);
nor U16218 (N_16218,N_13387,N_14982);
or U16219 (N_16219,N_12371,N_10973);
nor U16220 (N_16220,N_13034,N_13009);
nor U16221 (N_16221,N_11975,N_14917);
and U16222 (N_16222,N_13733,N_11002);
and U16223 (N_16223,N_12940,N_10518);
nand U16224 (N_16224,N_10638,N_10579);
nor U16225 (N_16225,N_12361,N_12854);
or U16226 (N_16226,N_11411,N_12667);
xor U16227 (N_16227,N_10847,N_14751);
and U16228 (N_16228,N_13977,N_14218);
nand U16229 (N_16229,N_12380,N_12475);
nor U16230 (N_16230,N_10881,N_10673);
and U16231 (N_16231,N_12935,N_11189);
or U16232 (N_16232,N_14421,N_11584);
or U16233 (N_16233,N_14266,N_12646);
and U16234 (N_16234,N_12407,N_10792);
and U16235 (N_16235,N_11107,N_10060);
nor U16236 (N_16236,N_10248,N_12501);
xor U16237 (N_16237,N_13300,N_13480);
or U16238 (N_16238,N_13636,N_14011);
and U16239 (N_16239,N_12053,N_14020);
or U16240 (N_16240,N_12691,N_13960);
or U16241 (N_16241,N_14188,N_14986);
nor U16242 (N_16242,N_12421,N_11789);
nor U16243 (N_16243,N_12014,N_10031);
nand U16244 (N_16244,N_14578,N_12408);
or U16245 (N_16245,N_14037,N_12660);
or U16246 (N_16246,N_13342,N_13534);
and U16247 (N_16247,N_11179,N_10038);
xnor U16248 (N_16248,N_12569,N_12815);
nand U16249 (N_16249,N_13989,N_12933);
xnor U16250 (N_16250,N_12692,N_11257);
and U16251 (N_16251,N_10384,N_10445);
nor U16252 (N_16252,N_13419,N_12864);
nand U16253 (N_16253,N_13008,N_14735);
or U16254 (N_16254,N_10143,N_13728);
and U16255 (N_16255,N_13997,N_10037);
and U16256 (N_16256,N_10729,N_12198);
xnor U16257 (N_16257,N_12633,N_10755);
nor U16258 (N_16258,N_10213,N_13610);
xor U16259 (N_16259,N_14745,N_13537);
xnor U16260 (N_16260,N_11906,N_12038);
nand U16261 (N_16261,N_11521,N_13469);
and U16262 (N_16262,N_10869,N_11965);
xnor U16263 (N_16263,N_12201,N_13328);
nor U16264 (N_16264,N_13130,N_14041);
nor U16265 (N_16265,N_11252,N_10302);
or U16266 (N_16266,N_14716,N_10090);
nand U16267 (N_16267,N_11812,N_12065);
or U16268 (N_16268,N_13748,N_10817);
nand U16269 (N_16269,N_13815,N_12684);
and U16270 (N_16270,N_10086,N_12270);
nand U16271 (N_16271,N_11198,N_12299);
and U16272 (N_16272,N_10268,N_10888);
nand U16273 (N_16273,N_10430,N_13251);
nor U16274 (N_16274,N_11989,N_12046);
nand U16275 (N_16275,N_11573,N_14445);
or U16276 (N_16276,N_11890,N_10641);
or U16277 (N_16277,N_13555,N_14167);
nand U16278 (N_16278,N_13018,N_14120);
or U16279 (N_16279,N_14333,N_11454);
nand U16280 (N_16280,N_13385,N_13751);
nor U16281 (N_16281,N_13607,N_10808);
xor U16282 (N_16282,N_10250,N_10485);
and U16283 (N_16283,N_13239,N_14898);
nand U16284 (N_16284,N_13459,N_12549);
or U16285 (N_16285,N_14927,N_12002);
and U16286 (N_16286,N_14115,N_13988);
and U16287 (N_16287,N_11381,N_13484);
or U16288 (N_16288,N_10602,N_11100);
xor U16289 (N_16289,N_10650,N_13964);
and U16290 (N_16290,N_11930,N_11164);
nand U16291 (N_16291,N_12028,N_10135);
nand U16292 (N_16292,N_14522,N_11426);
nor U16293 (N_16293,N_12768,N_12969);
nor U16294 (N_16294,N_14268,N_10739);
or U16295 (N_16295,N_13062,N_10317);
or U16296 (N_16296,N_11293,N_10963);
nand U16297 (N_16297,N_10245,N_12758);
and U16298 (N_16298,N_13609,N_14252);
and U16299 (N_16299,N_11199,N_10155);
and U16300 (N_16300,N_13235,N_13158);
nand U16301 (N_16301,N_13011,N_11808);
and U16302 (N_16302,N_12557,N_12631);
or U16303 (N_16303,N_14503,N_12771);
nand U16304 (N_16304,N_14511,N_13310);
and U16305 (N_16305,N_14300,N_10859);
nand U16306 (N_16306,N_10795,N_10639);
nand U16307 (N_16307,N_12097,N_13492);
and U16308 (N_16308,N_13624,N_14065);
and U16309 (N_16309,N_12695,N_10746);
or U16310 (N_16310,N_12279,N_10582);
nor U16311 (N_16311,N_14823,N_11306);
xnor U16312 (N_16312,N_10258,N_11487);
nor U16313 (N_16313,N_12311,N_14617);
xnor U16314 (N_16314,N_13811,N_12757);
nand U16315 (N_16315,N_13926,N_14743);
nor U16316 (N_16316,N_13213,N_11771);
or U16317 (N_16317,N_13809,N_11829);
nor U16318 (N_16318,N_13396,N_10549);
nor U16319 (N_16319,N_14627,N_11322);
or U16320 (N_16320,N_12971,N_11299);
and U16321 (N_16321,N_10943,N_11559);
and U16322 (N_16322,N_14981,N_14122);
or U16323 (N_16323,N_10108,N_14327);
or U16324 (N_16324,N_13570,N_10731);
and U16325 (N_16325,N_14900,N_10686);
or U16326 (N_16326,N_14264,N_12239);
xnor U16327 (N_16327,N_14719,N_14563);
nand U16328 (N_16328,N_12913,N_10555);
nor U16329 (N_16329,N_10063,N_11074);
nand U16330 (N_16330,N_10236,N_13350);
nor U16331 (N_16331,N_12862,N_11810);
nor U16332 (N_16332,N_12809,N_12606);
nor U16333 (N_16333,N_11272,N_10702);
and U16334 (N_16334,N_11270,N_14365);
nor U16335 (N_16335,N_13718,N_13765);
xor U16336 (N_16336,N_11275,N_13369);
and U16337 (N_16337,N_11526,N_11631);
or U16338 (N_16338,N_10167,N_13334);
or U16339 (N_16339,N_13895,N_14724);
or U16340 (N_16340,N_10025,N_13374);
and U16341 (N_16341,N_14896,N_12587);
nand U16342 (N_16342,N_13173,N_12868);
nor U16343 (N_16343,N_13770,N_11745);
nor U16344 (N_16344,N_12437,N_13371);
nor U16345 (N_16345,N_12246,N_11209);
xor U16346 (N_16346,N_12403,N_11383);
and U16347 (N_16347,N_13283,N_13041);
and U16348 (N_16348,N_12880,N_12495);
or U16349 (N_16349,N_13772,N_12047);
or U16350 (N_16350,N_12855,N_14057);
or U16351 (N_16351,N_11732,N_10098);
or U16352 (N_16352,N_12071,N_10889);
nor U16353 (N_16353,N_14593,N_12890);
or U16354 (N_16354,N_11308,N_10200);
xor U16355 (N_16355,N_10540,N_11641);
or U16356 (N_16356,N_14984,N_11405);
xor U16357 (N_16357,N_10256,N_12321);
or U16358 (N_16358,N_10500,N_12796);
and U16359 (N_16359,N_11648,N_13990);
and U16360 (N_16360,N_13841,N_12133);
nand U16361 (N_16361,N_11998,N_11679);
nor U16362 (N_16362,N_10232,N_13657);
nand U16363 (N_16363,N_14966,N_12825);
or U16364 (N_16364,N_10469,N_13643);
nor U16365 (N_16365,N_11672,N_11932);
or U16366 (N_16366,N_14357,N_11398);
and U16367 (N_16367,N_10303,N_10816);
nand U16368 (N_16368,N_12360,N_13958);
nand U16369 (N_16369,N_11907,N_14564);
or U16370 (N_16370,N_14742,N_11986);
nand U16371 (N_16371,N_10262,N_12400);
nand U16372 (N_16372,N_12722,N_10186);
or U16373 (N_16373,N_14865,N_14132);
nand U16374 (N_16374,N_13200,N_12732);
or U16375 (N_16375,N_11822,N_11135);
and U16376 (N_16376,N_11114,N_11509);
nand U16377 (N_16377,N_11187,N_11838);
nand U16378 (N_16378,N_14400,N_10512);
nand U16379 (N_16379,N_13042,N_10901);
nor U16380 (N_16380,N_10534,N_13665);
xor U16381 (N_16381,N_13233,N_13715);
and U16382 (N_16382,N_11756,N_13560);
and U16383 (N_16383,N_14231,N_11933);
nor U16384 (N_16384,N_13564,N_10985);
nand U16385 (N_16385,N_13346,N_10095);
nand U16386 (N_16386,N_11265,N_11133);
nor U16387 (N_16387,N_10202,N_11590);
or U16388 (N_16388,N_13868,N_14626);
nand U16389 (N_16389,N_12044,N_10460);
and U16390 (N_16390,N_13785,N_11061);
nand U16391 (N_16391,N_12708,N_11472);
xnor U16392 (N_16392,N_12480,N_13406);
nand U16393 (N_16393,N_10904,N_12818);
or U16394 (N_16394,N_12545,N_13514);
or U16395 (N_16395,N_14226,N_13094);
or U16396 (N_16396,N_14902,N_14399);
nor U16397 (N_16397,N_13950,N_12171);
nand U16398 (N_16398,N_11232,N_10184);
or U16399 (N_16399,N_12290,N_11140);
or U16400 (N_16400,N_12481,N_10065);
nand U16401 (N_16401,N_12946,N_11894);
or U16402 (N_16402,N_11558,N_14116);
nor U16403 (N_16403,N_12291,N_13224);
xnor U16404 (N_16404,N_10664,N_11511);
or U16405 (N_16405,N_12718,N_11946);
nand U16406 (N_16406,N_14726,N_13659);
or U16407 (N_16407,N_11203,N_11464);
nor U16408 (N_16408,N_14345,N_14633);
nor U16409 (N_16409,N_11282,N_14541);
and U16410 (N_16410,N_14910,N_11229);
xor U16411 (N_16411,N_12009,N_14274);
and U16412 (N_16412,N_12088,N_13402);
and U16413 (N_16413,N_10044,N_12883);
nor U16414 (N_16414,N_14736,N_11037);
nor U16415 (N_16415,N_13843,N_10677);
or U16416 (N_16416,N_14170,N_11050);
nor U16417 (N_16417,N_10156,N_14207);
nand U16418 (N_16418,N_13590,N_13860);
xnor U16419 (N_16419,N_11555,N_14853);
or U16420 (N_16420,N_13367,N_13688);
nor U16421 (N_16421,N_10094,N_14298);
and U16422 (N_16422,N_14844,N_14303);
and U16423 (N_16423,N_13954,N_10377);
nor U16424 (N_16424,N_14717,N_14284);
and U16425 (N_16425,N_11057,N_14040);
nor U16426 (N_16426,N_14249,N_10334);
or U16427 (N_16427,N_11042,N_11423);
or U16428 (N_16428,N_11846,N_13899);
nand U16429 (N_16429,N_13349,N_11047);
and U16430 (N_16430,N_13912,N_10733);
and U16431 (N_16431,N_11127,N_12264);
and U16432 (N_16432,N_14163,N_11038);
and U16433 (N_16433,N_10681,N_13503);
nor U16434 (N_16434,N_13244,N_11734);
and U16435 (N_16435,N_10187,N_13884);
or U16436 (N_16436,N_13701,N_13170);
or U16437 (N_16437,N_12828,N_10794);
and U16438 (N_16438,N_13057,N_10630);
xnor U16439 (N_16439,N_14309,N_13936);
or U16440 (N_16440,N_14997,N_11350);
or U16441 (N_16441,N_14888,N_12939);
nand U16442 (N_16442,N_12444,N_12507);
nand U16443 (N_16443,N_12558,N_10489);
xor U16444 (N_16444,N_12167,N_12188);
or U16445 (N_16445,N_11677,N_11638);
nor U16446 (N_16446,N_12490,N_14101);
nor U16447 (N_16447,N_10635,N_10228);
and U16448 (N_16448,N_13150,N_11023);
and U16449 (N_16449,N_11251,N_14023);
nor U16450 (N_16450,N_11767,N_14123);
and U16451 (N_16451,N_12375,N_10802);
and U16452 (N_16452,N_13299,N_14151);
nor U16453 (N_16453,N_12172,N_12672);
or U16454 (N_16454,N_14973,N_11366);
nor U16455 (N_16455,N_10805,N_11334);
and U16456 (N_16456,N_10960,N_14899);
or U16457 (N_16457,N_14201,N_10081);
and U16458 (N_16458,N_12886,N_14077);
or U16459 (N_16459,N_11793,N_13091);
nand U16460 (N_16460,N_14438,N_13797);
xor U16461 (N_16461,N_12889,N_11581);
nor U16462 (N_16462,N_14628,N_12120);
xnor U16463 (N_16463,N_12155,N_12122);
nor U16464 (N_16464,N_10033,N_14027);
nor U16465 (N_16465,N_10854,N_11572);
nand U16466 (N_16466,N_11358,N_12129);
nand U16467 (N_16467,N_11548,N_14658);
or U16468 (N_16468,N_10240,N_12596);
nor U16469 (N_16469,N_14443,N_12799);
and U16470 (N_16470,N_14941,N_12836);
or U16471 (N_16471,N_10356,N_14376);
nor U16472 (N_16472,N_14447,N_13101);
nand U16473 (N_16473,N_13289,N_12661);
nand U16474 (N_16474,N_12823,N_10422);
nand U16475 (N_16475,N_13666,N_10865);
or U16476 (N_16476,N_10734,N_13854);
nor U16477 (N_16477,N_12927,N_10926);
and U16478 (N_16478,N_13601,N_10120);
nand U16479 (N_16479,N_10754,N_10218);
nand U16480 (N_16480,N_13457,N_10651);
nor U16481 (N_16481,N_10455,N_14313);
and U16482 (N_16482,N_12036,N_12215);
xnor U16483 (N_16483,N_12625,N_14091);
and U16484 (N_16484,N_12577,N_10860);
nand U16485 (N_16485,N_12422,N_13847);
or U16486 (N_16486,N_13046,N_12785);
and U16487 (N_16487,N_10450,N_13933);
nand U16488 (N_16488,N_12580,N_13315);
and U16489 (N_16489,N_14753,N_13195);
or U16490 (N_16490,N_13338,N_14048);
xor U16491 (N_16491,N_12331,N_10272);
nor U16492 (N_16492,N_14148,N_13160);
or U16493 (N_16493,N_10848,N_14029);
or U16494 (N_16494,N_10550,N_11336);
and U16495 (N_16495,N_13725,N_13072);
and U16496 (N_16496,N_11046,N_11276);
nor U16497 (N_16497,N_11722,N_10009);
nand U16498 (N_16498,N_10209,N_10079);
and U16499 (N_16499,N_14426,N_10309);
and U16500 (N_16500,N_14546,N_13999);
and U16501 (N_16501,N_13741,N_12705);
nand U16502 (N_16502,N_13363,N_14442);
nand U16503 (N_16503,N_13022,N_11261);
and U16504 (N_16504,N_13381,N_14770);
nand U16505 (N_16505,N_14608,N_10800);
nor U16506 (N_16506,N_10473,N_10583);
nand U16507 (N_16507,N_14565,N_10674);
and U16508 (N_16508,N_10124,N_14601);
nor U16509 (N_16509,N_12600,N_11647);
nor U16510 (N_16510,N_11797,N_11517);
and U16511 (N_16511,N_10437,N_14025);
or U16512 (N_16512,N_11253,N_10556);
and U16513 (N_16513,N_10936,N_11234);
xnor U16514 (N_16514,N_12727,N_14030);
nor U16515 (N_16515,N_10861,N_10501);
and U16516 (N_16516,N_12990,N_14286);
or U16517 (N_16517,N_13185,N_13848);
or U16518 (N_16518,N_10740,N_14033);
and U16519 (N_16519,N_13805,N_11084);
and U16520 (N_16520,N_10254,N_14470);
nor U16521 (N_16521,N_12050,N_13263);
and U16522 (N_16522,N_13692,N_14127);
or U16523 (N_16523,N_10909,N_14912);
or U16524 (N_16524,N_13951,N_14959);
xnor U16525 (N_16525,N_13461,N_14428);
nand U16526 (N_16526,N_12379,N_13366);
nor U16527 (N_16527,N_13012,N_13390);
or U16528 (N_16528,N_10357,N_10937);
nand U16529 (N_16529,N_11719,N_13015);
nor U16530 (N_16530,N_14196,N_14777);
or U16531 (N_16531,N_10760,N_11212);
or U16532 (N_16532,N_13545,N_12571);
or U16533 (N_16533,N_10574,N_11201);
nor U16534 (N_16534,N_11627,N_13304);
xor U16535 (N_16535,N_12751,N_10774);
nand U16536 (N_16536,N_12166,N_11026);
and U16537 (N_16537,N_11453,N_10058);
and U16538 (N_16538,N_12327,N_12920);
or U16539 (N_16539,N_12438,N_14596);
or U16540 (N_16540,N_13431,N_10249);
nand U16541 (N_16541,N_12502,N_14164);
or U16542 (N_16542,N_10019,N_12968);
nand U16543 (N_16543,N_10592,N_11508);
and U16544 (N_16544,N_14928,N_11747);
or U16545 (N_16545,N_12776,N_10007);
nor U16546 (N_16546,N_14765,N_11680);
nor U16547 (N_16547,N_14536,N_12016);
and U16548 (N_16548,N_11574,N_14289);
nand U16549 (N_16549,N_11481,N_13475);
nand U16550 (N_16550,N_12240,N_10993);
or U16551 (N_16551,N_14845,N_13917);
nor U16552 (N_16552,N_10775,N_14648);
nand U16553 (N_16553,N_11432,N_12609);
or U16554 (N_16554,N_14703,N_14448);
and U16555 (N_16555,N_10521,N_13133);
nor U16556 (N_16556,N_10687,N_11395);
nand U16557 (N_16557,N_13746,N_11097);
or U16558 (N_16558,N_10331,N_12730);
and U16559 (N_16559,N_13814,N_13523);
and U16560 (N_16560,N_10078,N_12858);
nand U16561 (N_16561,N_10886,N_13807);
or U16562 (N_16562,N_14385,N_14762);
or U16563 (N_16563,N_12483,N_13201);
or U16564 (N_16564,N_10811,N_11592);
nand U16565 (N_16565,N_13407,N_10242);
nand U16566 (N_16566,N_11086,N_13743);
nand U16567 (N_16567,N_14210,N_11926);
or U16568 (N_16568,N_13268,N_10169);
nor U16569 (N_16569,N_10520,N_14187);
and U16570 (N_16570,N_14117,N_10029);
nor U16571 (N_16571,N_13632,N_13538);
and U16572 (N_16572,N_10141,N_11418);
nand U16573 (N_16573,N_10770,N_13129);
nor U16574 (N_16574,N_10148,N_14847);
and U16575 (N_16575,N_13247,N_11462);
or U16576 (N_16576,N_11343,N_14085);
xnor U16577 (N_16577,N_10472,N_14722);
nor U16578 (N_16578,N_10273,N_12525);
or U16579 (N_16579,N_12205,N_11103);
nor U16580 (N_16580,N_12964,N_12617);
nor U16581 (N_16581,N_11108,N_10646);
and U16582 (N_16582,N_11656,N_14768);
and U16583 (N_16583,N_14003,N_12579);
nand U16584 (N_16584,N_14312,N_13764);
or U16585 (N_16585,N_14310,N_14142);
nor U16586 (N_16586,N_14381,N_10590);
nor U16587 (N_16587,N_13059,N_11266);
and U16588 (N_16588,N_10071,N_10329);
nand U16589 (N_16589,N_12802,N_10194);
and U16590 (N_16590,N_12314,N_10933);
nor U16591 (N_16591,N_12634,N_14769);
nor U16592 (N_16592,N_13529,N_12402);
nand U16593 (N_16593,N_10406,N_10965);
xor U16594 (N_16594,N_13108,N_14338);
nand U16595 (N_16595,N_13135,N_11977);
and U16596 (N_16596,N_10022,N_14866);
nor U16597 (N_16597,N_12724,N_13223);
or U16598 (N_16598,N_13114,N_11177);
or U16599 (N_16599,N_14805,N_13500);
and U16600 (N_16600,N_10907,N_10338);
nor U16601 (N_16601,N_13553,N_11836);
nor U16602 (N_16602,N_14248,N_11537);
nand U16603 (N_16603,N_11277,N_14731);
nor U16604 (N_16604,N_12753,N_12464);
nor U16605 (N_16605,N_12665,N_10016);
nor U16606 (N_16606,N_13186,N_14028);
and U16607 (N_16607,N_12429,N_13602);
nor U16608 (N_16608,N_13861,N_12824);
nor U16609 (N_16609,N_12509,N_10150);
or U16610 (N_16610,N_11955,N_14646);
or U16611 (N_16611,N_14152,N_11814);
and U16612 (N_16612,N_13058,N_13420);
or U16613 (N_16613,N_13440,N_11799);
and U16614 (N_16614,N_14238,N_13878);
or U16615 (N_16615,N_12923,N_13063);
and U16616 (N_16616,N_12106,N_14113);
and U16617 (N_16617,N_14606,N_11730);
nand U16618 (N_16618,N_10552,N_13916);
nor U16619 (N_16619,N_14715,N_14095);
and U16620 (N_16620,N_13393,N_10757);
and U16621 (N_16621,N_10896,N_10394);
and U16622 (N_16622,N_11674,N_12550);
and U16623 (N_16623,N_10778,N_14108);
nand U16624 (N_16624,N_14347,N_10621);
nand U16625 (N_16625,N_14068,N_14501);
and U16626 (N_16626,N_12897,N_13403);
nor U16627 (N_16627,N_11231,N_14356);
and U16628 (N_16628,N_10571,N_10123);
and U16629 (N_16629,N_14576,N_14477);
nand U16630 (N_16630,N_14586,N_11962);
xnor U16631 (N_16631,N_13293,N_14308);
or U16632 (N_16632,N_12639,N_13706);
nor U16633 (N_16633,N_13377,N_11964);
nor U16634 (N_16634,N_12787,N_11267);
and U16635 (N_16635,N_11401,N_10168);
nand U16636 (N_16636,N_10006,N_12471);
and U16637 (N_16637,N_11493,N_10107);
xnor U16638 (N_16638,N_12706,N_14255);
nor U16639 (N_16639,N_11082,N_10435);
nor U16640 (N_16640,N_13359,N_10879);
nand U16641 (N_16641,N_10935,N_12508);
nor U16642 (N_16642,N_11785,N_11355);
nand U16643 (N_16643,N_12650,N_11935);
and U16644 (N_16644,N_10419,N_11868);
nand U16645 (N_16645,N_11237,N_11750);
nor U16646 (N_16646,N_14508,N_12398);
nor U16647 (N_16647,N_10291,N_10364);
xnor U16648 (N_16648,N_14649,N_12821);
or U16649 (N_16649,N_10068,N_13716);
nand U16650 (N_16650,N_12341,N_13780);
nor U16651 (N_16651,N_10177,N_14836);
or U16652 (N_16652,N_14050,N_13302);
and U16653 (N_16653,N_12034,N_10668);
nor U16654 (N_16654,N_12288,N_12601);
nor U16655 (N_16655,N_12680,N_11053);
or U16656 (N_16656,N_12786,N_10594);
and U16657 (N_16657,N_12258,N_10614);
nand U16658 (N_16658,N_11724,N_14826);
or U16659 (N_16659,N_12300,N_11825);
xor U16660 (N_16660,N_12826,N_13364);
and U16661 (N_16661,N_13144,N_13837);
nor U16662 (N_16662,N_11693,N_12146);
nand U16663 (N_16663,N_12329,N_12711);
nand U16664 (N_16664,N_11775,N_13176);
nor U16665 (N_16665,N_10954,N_10115);
nor U16666 (N_16666,N_14760,N_13567);
or U16667 (N_16667,N_11995,N_14016);
xor U16668 (N_16668,N_14368,N_13199);
and U16669 (N_16669,N_13616,N_12063);
nand U16670 (N_16670,N_13930,N_13675);
xor U16671 (N_16671,N_11269,N_12077);
nand U16672 (N_16672,N_13450,N_11451);
nor U16673 (N_16673,N_12005,N_12986);
nand U16674 (N_16674,N_10318,N_12406);
nor U16675 (N_16675,N_13532,N_13892);
or U16676 (N_16676,N_12352,N_14403);
nand U16677 (N_16677,N_10059,N_10072);
or U16678 (N_16678,N_13330,N_11284);
nor U16679 (N_16679,N_12085,N_14056);
xor U16680 (N_16680,N_10405,N_12017);
or U16681 (N_16681,N_12655,N_12156);
xnor U16682 (N_16682,N_12347,N_13481);
nand U16683 (N_16683,N_12135,N_10497);
nor U16684 (N_16684,N_12704,N_11957);
nand U16685 (N_16685,N_13044,N_10836);
nand U16686 (N_16686,N_10021,N_12157);
or U16687 (N_16687,N_13737,N_12194);
nand U16688 (N_16688,N_11271,N_12214);
or U16689 (N_16689,N_14971,N_11725);
xnor U16690 (N_16690,N_11908,N_13803);
or U16691 (N_16691,N_14950,N_10170);
xnor U16692 (N_16692,N_11402,N_11624);
or U16693 (N_16693,N_13236,N_12518);
and U16694 (N_16694,N_13149,N_11534);
nand U16695 (N_16695,N_12813,N_11779);
and U16696 (N_16696,N_11332,N_14562);
and U16697 (N_16697,N_11387,N_14803);
and U16698 (N_16698,N_14595,N_11325);
nand U16699 (N_16699,N_12847,N_14820);
xnor U16700 (N_16700,N_11003,N_11099);
and U16701 (N_16701,N_12583,N_13761);
or U16702 (N_16702,N_11419,N_13776);
and U16703 (N_16703,N_10930,N_14339);
nor U16704 (N_16704,N_11878,N_10810);
and U16705 (N_16705,N_13522,N_13405);
or U16706 (N_16706,N_13550,N_12301);
and U16707 (N_16707,N_11934,N_13229);
nand U16708 (N_16708,N_14682,N_14747);
or U16709 (N_16709,N_13707,N_12659);
nand U16710 (N_16710,N_14483,N_14904);
nor U16711 (N_16711,N_13768,N_12926);
nand U16712 (N_16712,N_12827,N_12616);
and U16713 (N_16713,N_12354,N_12251);
and U16714 (N_16714,N_10712,N_13060);
nand U16715 (N_16715,N_12178,N_14407);
xor U16716 (N_16716,N_14809,N_14980);
nand U16717 (N_16717,N_12837,N_11351);
nor U16718 (N_16718,N_11382,N_14965);
nor U16719 (N_16719,N_13597,N_14780);
or U16720 (N_16720,N_13029,N_10632);
and U16721 (N_16721,N_13049,N_10982);
nand U16722 (N_16722,N_12304,N_12678);
and U16723 (N_16723,N_13411,N_12546);
or U16724 (N_16724,N_13506,N_14498);
nand U16725 (N_16725,N_13256,N_11643);
or U16726 (N_16726,N_11634,N_10633);
or U16727 (N_16727,N_12316,N_14389);
nor U16728 (N_16728,N_12435,N_14072);
or U16729 (N_16729,N_13477,N_11941);
or U16730 (N_16730,N_11482,N_11434);
nand U16731 (N_16731,N_13934,N_14476);
or U16732 (N_16732,N_10479,N_10293);
and U16733 (N_16733,N_11064,N_11968);
and U16734 (N_16734,N_11384,N_13437);
and U16735 (N_16735,N_14129,N_10887);
and U16736 (N_16736,N_10028,N_14645);
or U16737 (N_16737,N_11394,N_11323);
nand U16738 (N_16738,N_12138,N_11869);
nand U16739 (N_16739,N_12473,N_12527);
nor U16740 (N_16740,N_10292,N_11262);
nor U16741 (N_16741,N_11066,N_12460);
nor U16742 (N_16742,N_12026,N_11642);
nand U16743 (N_16743,N_12144,N_11760);
nand U16744 (N_16744,N_12061,N_10287);
and U16745 (N_16745,N_11063,N_11780);
and U16746 (N_16746,N_12497,N_12236);
nor U16747 (N_16747,N_13821,N_11914);
and U16748 (N_16748,N_13667,N_14516);
or U16749 (N_16749,N_11000,N_10101);
or U16750 (N_16750,N_14877,N_10299);
and U16751 (N_16751,N_10979,N_14420);
or U16752 (N_16752,N_13593,N_14929);
nor U16753 (N_16753,N_11300,N_14307);
xor U16754 (N_16754,N_12967,N_13193);
xnor U16755 (N_16755,N_13020,N_11309);
xor U16756 (N_16756,N_10864,N_14939);
or U16757 (N_16757,N_12689,N_11960);
xnor U16758 (N_16758,N_13033,N_13668);
nand U16759 (N_16759,N_13986,N_13208);
nor U16760 (N_16760,N_11707,N_11727);
and U16761 (N_16761,N_10442,N_11069);
nand U16762 (N_16762,N_10692,N_11056);
nand U16763 (N_16763,N_11486,N_11821);
and U16764 (N_16764,N_14179,N_11532);
nand U16765 (N_16765,N_10618,N_14154);
nand U16766 (N_16766,N_11597,N_14370);
and U16767 (N_16767,N_13835,N_11764);
and U16768 (N_16768,N_13494,N_13684);
and U16769 (N_16769,N_12195,N_14889);
and U16770 (N_16770,N_12592,N_14281);
or U16771 (N_16771,N_13376,N_12208);
xor U16772 (N_16772,N_14126,N_13965);
nor U16773 (N_16773,N_14469,N_12109);
nand U16774 (N_16774,N_11142,N_11802);
nor U16775 (N_16775,N_10765,N_10459);
nand U16776 (N_16776,N_14786,N_14775);
nor U16777 (N_16777,N_10432,N_10903);
or U16778 (N_16778,N_12533,N_12057);
nor U16779 (N_16779,N_11744,N_11502);
nor U16780 (N_16780,N_14610,N_12843);
and U16781 (N_16781,N_11274,N_13325);
or U16782 (N_16782,N_10462,N_14961);
and U16783 (N_16783,N_12775,N_14972);
nor U16784 (N_16784,N_10211,N_13408);
nand U16785 (N_16785,N_13312,N_11172);
nand U16786 (N_16786,N_12330,N_11938);
nand U16787 (N_16787,N_10551,N_13152);
nand U16788 (N_16788,N_12793,N_14323);
nand U16789 (N_16789,N_11828,N_10783);
nand U16790 (N_16790,N_11605,N_14813);
and U16791 (N_16791,N_12694,N_13862);
nor U16792 (N_16792,N_12263,N_12449);
nand U16793 (N_16793,N_12450,N_13873);
nor U16794 (N_16794,N_11754,N_10330);
xnor U16795 (N_16795,N_10665,N_11971);
and U16796 (N_16796,N_14178,N_12685);
xor U16797 (N_16797,N_11497,N_11811);
or U16798 (N_16798,N_14864,N_14921);
or U16799 (N_16799,N_14261,N_13035);
nand U16800 (N_16800,N_10411,N_11294);
or U16801 (N_16801,N_11834,N_10403);
nand U16802 (N_16802,N_14653,N_14110);
or U16803 (N_16803,N_14831,N_11406);
nor U16804 (N_16804,N_10939,N_14044);
nor U16805 (N_16805,N_10153,N_13100);
nand U16806 (N_16806,N_11591,N_13171);
and U16807 (N_16807,N_10599,N_12738);
or U16808 (N_16808,N_12207,N_10637);
nand U16809 (N_16809,N_12179,N_12664);
nand U16810 (N_16810,N_11949,N_14702);
and U16811 (N_16811,N_13414,N_14206);
nor U16812 (N_16812,N_13678,N_12907);
or U16813 (N_16813,N_14344,N_12805);
nand U16814 (N_16814,N_10642,N_10656);
and U16815 (N_16815,N_13974,N_10690);
nand U16816 (N_16816,N_10070,N_13646);
nand U16817 (N_16817,N_10857,N_13886);
nor U16818 (N_16818,N_12137,N_10750);
xnor U16819 (N_16819,N_13915,N_10539);
nor U16820 (N_16820,N_12766,N_10643);
and U16821 (N_16821,N_10229,N_10495);
or U16822 (N_16822,N_11875,N_13796);
xor U16823 (N_16823,N_14974,N_14002);
nor U16824 (N_16824,N_11676,N_12287);
and U16825 (N_16825,N_12374,N_14352);
nand U16826 (N_16826,N_10001,N_10307);
or U16827 (N_16827,N_12564,N_10373);
nor U16828 (N_16828,N_11580,N_14672);
nor U16829 (N_16829,N_13730,N_14216);
or U16830 (N_16830,N_10723,N_10830);
nand U16831 (N_16831,N_14463,N_12656);
nor U16832 (N_16832,N_10427,N_13962);
nand U16833 (N_16833,N_11954,N_13489);
and U16834 (N_16834,N_14125,N_10845);
and U16835 (N_16835,N_14947,N_10991);
and U16836 (N_16836,N_13750,N_10049);
and U16837 (N_16837,N_12628,N_14177);
nor U16838 (N_16838,N_13255,N_14840);
nor U16839 (N_16839,N_12362,N_13452);
xor U16840 (N_16840,N_13577,N_12976);
or U16841 (N_16841,N_12936,N_11408);
nand U16842 (N_16842,N_14013,N_12559);
nor U16843 (N_16843,N_12849,N_11871);
nor U16844 (N_16844,N_10260,N_14675);
or U16845 (N_16845,N_12458,N_14579);
or U16846 (N_16846,N_14599,N_14374);
xor U16847 (N_16847,N_12699,N_10225);
and U16848 (N_16848,N_11067,N_11190);
nand U16849 (N_16849,N_12226,N_12383);
or U16850 (N_16850,N_11507,N_13204);
and U16851 (N_16851,N_13858,N_12922);
nand U16852 (N_16852,N_14054,N_10136);
nor U16853 (N_16853,N_10371,N_12105);
nor U16854 (N_16854,N_13179,N_11079);
and U16855 (N_16855,N_12103,N_13220);
nand U16856 (N_16856,N_11425,N_13928);
nand U16857 (N_16857,N_11668,N_12165);
or U16858 (N_16858,N_11816,N_11320);
and U16859 (N_16859,N_12272,N_12744);
nor U16860 (N_16860,N_14092,N_14336);
or U16861 (N_16861,N_14916,N_11122);
or U16862 (N_16862,N_12534,N_12981);
nor U16863 (N_16863,N_11245,N_10465);
or U16864 (N_16864,N_14624,N_10423);
and U16865 (N_16865,N_13670,N_13879);
or U16866 (N_16866,N_10653,N_11882);
and U16867 (N_16867,N_14144,N_11101);
or U16868 (N_16868,N_11241,N_12456);
and U16869 (N_16869,N_11373,N_13579);
and U16870 (N_16870,N_14214,N_12498);
nand U16871 (N_16871,N_11205,N_12581);
nand U16872 (N_16872,N_12662,N_12947);
nor U16873 (N_16873,N_12513,N_12092);
nor U16874 (N_16874,N_12350,N_12630);
and U16875 (N_16875,N_13685,N_13510);
xnor U16876 (N_16876,N_11540,N_13162);
nand U16877 (N_16877,N_10949,N_13178);
and U16878 (N_16878,N_10609,N_14409);
nand U16879 (N_16879,N_13976,N_10948);
xor U16880 (N_16880,N_14386,N_13361);
nor U16881 (N_16881,N_13232,N_12191);
or U16882 (N_16882,N_12162,N_11089);
xor U16883 (N_16883,N_12369,N_10223);
nor U16884 (N_16884,N_13897,N_14673);
nand U16885 (N_16885,N_11800,N_11080);
nor U16886 (N_16886,N_13945,N_11049);
nand U16887 (N_16887,N_13754,N_12723);
or U16888 (N_16888,N_13324,N_13321);
nor U16889 (N_16889,N_10820,N_10659);
xor U16890 (N_16890,N_11024,N_10711);
xnor U16891 (N_16891,N_13528,N_13711);
and U16892 (N_16892,N_10875,N_12332);
nand U16893 (N_16893,N_12790,N_12988);
nand U16894 (N_16894,N_11611,N_14603);
and U16895 (N_16895,N_13919,N_10837);
and U16896 (N_16896,N_14183,N_11645);
and U16897 (N_16897,N_10208,N_13825);
or U16898 (N_16898,N_10516,N_13795);
nand U16899 (N_16899,N_13064,N_10417);
xor U16900 (N_16900,N_14605,N_11970);
nor U16901 (N_16901,N_14990,N_14814);
nand U16902 (N_16902,N_11463,N_11242);
or U16903 (N_16903,N_12278,N_12958);
nor U16904 (N_16904,N_14058,N_11576);
or U16905 (N_16905,N_14146,N_13273);
nand U16906 (N_16906,N_11594,N_12755);
or U16907 (N_16907,N_13781,N_10622);
and U16908 (N_16908,N_10383,N_13221);
or U16909 (N_16909,N_12250,N_13902);
or U16910 (N_16910,N_11841,N_13637);
nor U16911 (N_16911,N_14340,N_11044);
nor U16912 (N_16912,N_14406,N_12693);
nor U16913 (N_16913,N_11891,N_11762);
nand U16914 (N_16914,N_12414,N_10855);
and U16915 (N_16915,N_10397,N_10204);
and U16916 (N_16916,N_10648,N_14100);
nor U16917 (N_16917,N_11316,N_11751);
or U16918 (N_16918,N_14461,N_11492);
or U16919 (N_16919,N_13417,N_10923);
or U16920 (N_16920,N_11310,N_13479);
or U16921 (N_16921,N_11927,N_10922);
xnor U16922 (N_16922,N_14156,N_10114);
or U16923 (N_16923,N_11617,N_10684);
nand U16924 (N_16924,N_11948,N_13286);
nor U16925 (N_16925,N_10238,N_14366);
xnor U16926 (N_16926,N_13918,N_10214);
or U16927 (N_16927,N_14930,N_10048);
nand U16928 (N_16928,N_14294,N_11480);
nor U16929 (N_16929,N_14096,N_11662);
nand U16930 (N_16930,N_10874,N_12916);
or U16931 (N_16931,N_13379,N_13644);
nor U16932 (N_16932,N_11361,N_14665);
nand U16933 (N_16933,N_14614,N_11087);
nor U16934 (N_16934,N_13586,N_10910);
xnor U16935 (N_16935,N_10032,N_14288);
nor U16936 (N_16936,N_12054,N_12908);
and U16937 (N_16937,N_10636,N_12717);
nor U16938 (N_16938,N_11915,N_11244);
nor U16939 (N_16939,N_14031,N_14080);
xor U16940 (N_16940,N_13307,N_10581);
or U16941 (N_16941,N_12876,N_13907);
nand U16942 (N_16942,N_10955,N_14464);
or U16943 (N_16943,N_10871,N_12385);
nand U16944 (N_16944,N_14744,N_11791);
or U16945 (N_16945,N_10174,N_13109);
and U16946 (N_16946,N_11256,N_14481);
and U16947 (N_16947,N_12487,N_13566);
and U16948 (N_16948,N_14709,N_11473);
or U16949 (N_16949,N_10627,N_10928);
and U16950 (N_16950,N_13937,N_12560);
or U16951 (N_16951,N_10440,N_12443);
or U16952 (N_16952,N_12359,N_12455);
and U16953 (N_16953,N_12008,N_13231);
nand U16954 (N_16954,N_13267,N_14572);
or U16955 (N_16955,N_13316,N_13274);
nand U16956 (N_16956,N_12141,N_11916);
nor U16957 (N_16957,N_13720,N_13526);
or U16958 (N_16958,N_11039,N_11644);
and U16959 (N_16959,N_12274,N_12911);
nor U16960 (N_16960,N_13252,N_10625);
nand U16961 (N_16961,N_12150,N_14412);
or U16962 (N_16962,N_14573,N_10281);
or U16963 (N_16963,N_11138,N_13279);
xor U16964 (N_16964,N_11766,N_12952);
nor U16965 (N_16965,N_12295,N_14086);
or U16966 (N_16966,N_10882,N_11461);
or U16967 (N_16967,N_11621,N_11889);
and U16968 (N_16968,N_10862,N_12995);
or U16969 (N_16969,N_10644,N_12591);
xor U16970 (N_16970,N_11519,N_10813);
and U16971 (N_16971,N_14968,N_12015);
and U16972 (N_16972,N_10056,N_14854);
nor U16973 (N_16973,N_13826,N_12221);
and U16974 (N_16974,N_10381,N_14135);
nand U16975 (N_16975,N_10491,N_11545);
nand U16976 (N_16976,N_11072,N_12781);
nor U16977 (N_16977,N_10118,N_13652);
xor U16978 (N_16978,N_13143,N_12023);
xnor U16979 (N_16979,N_14647,N_11202);
and U16980 (N_16980,N_10649,N_12653);
or U16981 (N_16981,N_10368,N_12759);
xor U16982 (N_16982,N_10404,N_14377);
or U16983 (N_16983,N_11414,N_10166);
nor U16984 (N_16984,N_13125,N_13615);
and U16985 (N_16985,N_14159,N_13329);
nor U16986 (N_16986,N_10585,N_12149);
nor U16987 (N_16987,N_11575,N_13177);
nand U16988 (N_16988,N_13409,N_14314);
and U16989 (N_16989,N_10471,N_10410);
nand U16990 (N_16990,N_13650,N_10363);
nand U16991 (N_16991,N_11850,N_12445);
or U16992 (N_16992,N_13119,N_12118);
or U16993 (N_16993,N_14524,N_11807);
and U16994 (N_16994,N_12401,N_11048);
nand U16995 (N_16995,N_14739,N_12526);
or U16996 (N_16996,N_14830,N_10335);
nand U16997 (N_16997,N_10832,N_12556);
nor U16998 (N_16998,N_10919,N_12461);
and U16999 (N_16999,N_10230,N_13985);
and U17000 (N_17000,N_11774,N_12298);
nand U17001 (N_17001,N_11018,N_12364);
and U17002 (N_17002,N_12163,N_10941);
and U17003 (N_17003,N_12619,N_13584);
nand U17004 (N_17004,N_13696,N_10558);
xnor U17005 (N_17005,N_14884,N_11389);
and U17006 (N_17006,N_12957,N_14222);
and U17007 (N_17007,N_14652,N_14876);
or U17008 (N_17008,N_10133,N_13031);
xnor U17009 (N_17009,N_13581,N_14837);
or U17010 (N_17010,N_13112,N_13217);
xnor U17011 (N_17011,N_11160,N_11016);
and U17012 (N_17012,N_14859,N_12080);
nand U17013 (N_17013,N_14229,N_12185);
and U17014 (N_17014,N_12254,N_12590);
and U17015 (N_17015,N_10615,N_12966);
and U17016 (N_17016,N_12924,N_10833);
and U17017 (N_17017,N_12476,N_10395);
or U17018 (N_17018,N_12136,N_11259);
and U17019 (N_17019,N_10748,N_10541);
nor U17020 (N_17020,N_13987,N_11861);
nand U17021 (N_17021,N_10569,N_11467);
nand U17022 (N_17022,N_10047,N_10883);
nor U17023 (N_17023,N_13984,N_11339);
nor U17024 (N_17024,N_13368,N_10503);
xnor U17025 (N_17025,N_12463,N_14046);
and U17026 (N_17026,N_11991,N_10663);
or U17027 (N_17027,N_12638,N_10312);
nor U17028 (N_17028,N_12397,N_14215);
nor U17029 (N_17029,N_12991,N_10231);
and U17030 (N_17030,N_10967,N_10670);
and U17031 (N_17031,N_14825,N_13386);
nand U17032 (N_17032,N_14038,N_11692);
nand U17033 (N_17033,N_10160,N_11684);
and U17034 (N_17034,N_10956,N_11219);
or U17035 (N_17035,N_13470,N_14561);
nor U17036 (N_17036,N_12859,N_11263);
nor U17037 (N_17037,N_14642,N_13753);
and U17038 (N_17038,N_14099,N_11348);
and U17039 (N_17039,N_11307,N_11601);
or U17040 (N_17040,N_14734,N_12637);
nand U17041 (N_17041,N_13245,N_14858);
and U17042 (N_17042,N_11030,N_14493);
or U17043 (N_17043,N_11317,N_13174);
xor U17044 (N_17044,N_10203,N_13357);
xnor U17045 (N_17045,N_11787,N_11455);
and U17046 (N_17046,N_14689,N_12104);
nor U17047 (N_17047,N_11625,N_14677);
nor U17048 (N_17048,N_13699,N_14049);
and U17049 (N_17049,N_12675,N_12090);
nand U17050 (N_17050,N_12895,N_10074);
and U17051 (N_17051,N_14405,N_11981);
or U17052 (N_17052,N_11512,N_14324);
and U17053 (N_17053,N_10064,N_13106);
nor U17054 (N_17054,N_11606,N_14150);
and U17055 (N_17055,N_10159,N_14749);
and U17056 (N_17056,N_13942,N_10496);
nand U17057 (N_17057,N_10682,N_14538);
nand U17058 (N_17058,N_10893,N_11015);
nand U17059 (N_17059,N_14449,N_14991);
nand U17060 (N_17060,N_12161,N_11319);
nor U17061 (N_17061,N_10841,N_10838);
nor U17062 (N_17062,N_13840,N_11438);
or U17063 (N_17063,N_13611,N_11783);
xor U17064 (N_17064,N_13005,N_14835);
and U17065 (N_17065,N_14640,N_14355);
xnor U17066 (N_17066,N_10801,N_14727);
nor U17067 (N_17067,N_11040,N_10477);
and U17068 (N_17068,N_13142,N_13308);
or U17069 (N_17069,N_10920,N_10393);
nor U17070 (N_17070,N_13086,N_10276);
and U17071 (N_17071,N_11670,N_12555);
or U17072 (N_17072,N_14577,N_13801);
nor U17073 (N_17073,N_14326,N_12536);
or U17074 (N_17074,N_12322,N_11092);
xor U17075 (N_17075,N_13416,N_14378);
nand U17076 (N_17076,N_11197,N_10987);
or U17077 (N_17077,N_11148,N_11557);
nand U17078 (N_17078,N_14396,N_10905);
and U17079 (N_17079,N_10314,N_13822);
xnor U17080 (N_17080,N_11357,N_14714);
nand U17081 (N_17081,N_14841,N_12774);
nor U17082 (N_17082,N_13927,N_13521);
and U17083 (N_17083,N_13222,N_12367);
nor U17084 (N_17084,N_12095,N_11112);
and U17085 (N_17085,N_12535,N_10730);
and U17086 (N_17086,N_13677,N_11225);
xor U17087 (N_17087,N_12878,N_12140);
nor U17088 (N_17088,N_11705,N_11228);
nand U17089 (N_17089,N_13002,N_14656);
or U17090 (N_17090,N_11880,N_10728);
nand U17091 (N_17091,N_10119,N_10488);
xor U17092 (N_17092,N_11083,N_12209);
nor U17093 (N_17093,N_14246,N_12760);
nand U17094 (N_17094,N_11888,N_14848);
nand U17095 (N_17095,N_11685,N_10688);
or U17096 (N_17096,N_12412,N_11848);
nor U17097 (N_17097,N_14496,N_14639);
nor U17098 (N_17098,N_12041,N_10112);
nand U17099 (N_17099,N_11937,N_13205);
nor U17100 (N_17100,N_13786,N_14644);
and U17101 (N_17101,N_14987,N_11327);
nand U17102 (N_17102,N_13940,N_13556);
xnor U17103 (N_17103,N_14654,N_11505);
and U17104 (N_17104,N_10716,N_14523);
and U17105 (N_17105,N_11465,N_10030);
or U17106 (N_17106,N_11513,N_12885);
nand U17107 (N_17107,N_10267,N_13516);
nand U17108 (N_17108,N_11689,N_12271);
or U17109 (N_17109,N_11982,N_13689);
or U17110 (N_17110,N_12035,N_14471);
and U17111 (N_17111,N_14502,N_12083);
or U17112 (N_17112,N_12235,N_10508);
nand U17113 (N_17113,N_14824,N_13242);
and U17114 (N_17114,N_14808,N_13704);
nand U17115 (N_17115,N_13259,N_10562);
xor U17116 (N_17116,N_13542,N_13234);
or U17117 (N_17117,N_11530,N_10470);
nand U17118 (N_17118,N_13804,N_10790);
and U17119 (N_17119,N_14616,N_10494);
nor U17120 (N_17120,N_13880,N_12436);
and U17121 (N_17121,N_10121,N_13533);
and U17122 (N_17122,N_12339,N_12869);
or U17123 (N_17123,N_14416,N_13585);
nor U17124 (N_17124,N_10076,N_11289);
nor U17125 (N_17125,N_13081,N_12904);
or U17126 (N_17126,N_14311,N_13113);
and U17127 (N_17127,N_12697,N_10447);
and U17128 (N_17128,N_12632,N_11845);
or U17129 (N_17129,N_11020,N_13339);
and U17130 (N_17130,N_14873,N_12955);
or U17131 (N_17131,N_10799,N_14850);
nor U17132 (N_17132,N_10961,N_14121);
nand U17133 (N_17133,N_12720,N_13824);
and U17134 (N_17134,N_11477,N_10655);
nor U17135 (N_17135,N_14834,N_14358);
xnor U17136 (N_17136,N_12393,N_13700);
nor U17137 (N_17137,N_12800,N_13327);
xor U17138 (N_17138,N_10784,N_14585);
or U17139 (N_17139,N_14807,N_12181);
or U17140 (N_17140,N_11629,N_14241);
xor U17141 (N_17141,N_13589,N_14008);
or U17142 (N_17142,N_12292,N_11536);
nand U17143 (N_17143,N_11813,N_10305);
nor U17144 (N_17144,N_13783,N_13356);
and U17145 (N_17145,N_12612,N_13839);
nand U17146 (N_17146,N_12573,N_13270);
xnor U17147 (N_17147,N_10713,N_13467);
and U17148 (N_17148,N_10983,N_10927);
and U17149 (N_17149,N_11902,N_11528);
xnor U17150 (N_17150,N_11682,N_11264);
and U17151 (N_17151,N_10999,N_14733);
xnor U17152 (N_17152,N_11755,N_14707);
nand U17153 (N_17153,N_11416,N_11665);
and U17154 (N_17154,N_12392,N_10938);
nand U17155 (N_17155,N_14922,N_10415);
xor U17156 (N_17156,N_10525,N_12565);
nor U17157 (N_17157,N_13499,N_12173);
nand U17158 (N_17158,N_14544,N_14232);
xnor U17159 (N_17159,N_10054,N_14588);
nor U17160 (N_17160,N_13003,N_14905);
nand U17161 (N_17161,N_10997,N_11077);
or U17162 (N_17162,N_14795,N_11021);
nand U17163 (N_17163,N_11342,N_14787);
and U17164 (N_17164,N_12349,N_13442);
or U17165 (N_17165,N_10768,N_13681);
nor U17166 (N_17166,N_12589,N_12626);
nand U17167 (N_17167,N_14219,N_14772);
nor U17168 (N_17168,N_13362,N_12879);
and U17169 (N_17169,N_12773,N_13651);
nand U17170 (N_17170,N_10097,N_11017);
nand U17171 (N_17171,N_11911,N_11013);
xor U17172 (N_17172,N_14513,N_12635);
xor U17173 (N_17173,N_11033,N_12212);
xor U17174 (N_17174,N_11698,N_14147);
nand U17175 (N_17175,N_14230,N_10175);
nor U17176 (N_17176,N_10173,N_13806);
nand U17177 (N_17177,N_10306,N_12860);
nand U17178 (N_17178,N_10361,N_12603);
and U17179 (N_17179,N_13763,N_11280);
nand U17180 (N_17180,N_13676,N_14666);
or U17181 (N_17181,N_10014,N_14182);
nor U17182 (N_17182,N_13888,N_10446);
nand U17183 (N_17183,N_13249,N_13131);
nor U17184 (N_17184,N_14870,N_12377);
xnor U17185 (N_17185,N_14728,N_10319);
and U17186 (N_17186,N_12572,N_10986);
nand U17187 (N_17187,N_12756,N_12598);
xnor U17188 (N_17188,N_11776,N_14797);
xor U17189 (N_17189,N_10523,N_14611);
nor U17190 (N_17190,N_14943,N_12528);
nand U17191 (N_17191,N_13694,N_13956);
nand U17192 (N_17192,N_13054,N_14931);
and U17193 (N_17193,N_10914,N_13691);
or U17194 (N_17194,N_11694,N_12938);
and U17195 (N_17195,N_11094,N_14045);
and U17196 (N_17196,N_11184,N_14114);
or U17197 (N_17197,N_11174,N_10257);
nor U17198 (N_17198,N_11442,N_10601);
or U17199 (N_17199,N_14484,N_12241);
and U17200 (N_17200,N_12736,N_10773);
or U17201 (N_17201,N_12176,N_14306);
or U17202 (N_17202,N_14890,N_12762);
nor U17203 (N_17203,N_13961,N_10104);
or U17204 (N_17204,N_11604,N_14740);
xor U17205 (N_17205,N_14891,N_13791);
nand U17206 (N_17206,N_11154,N_11078);
nor U17207 (N_17207,N_11035,N_11290);
nand U17208 (N_17208,N_10126,N_14221);
nand U17209 (N_17209,N_13076,N_13126);
and U17210 (N_17210,N_13189,N_11413);
or U17211 (N_17211,N_11286,N_13724);
or U17212 (N_17212,N_14034,N_11062);
xor U17213 (N_17213,N_12275,N_10429);
nor U17214 (N_17214,N_14507,N_13619);
xnor U17215 (N_17215,N_11918,N_12765);
nor U17216 (N_17216,N_12335,N_11495);
and U17217 (N_17217,N_10366,N_14367);
or U17218 (N_17218,N_12644,N_11854);
and U17219 (N_17219,N_13635,N_13844);
or U17220 (N_17220,N_12132,N_14550);
nor U17221 (N_17221,N_12020,N_14861);
nor U17222 (N_17222,N_10776,N_11805);
nand U17223 (N_17223,N_10181,N_11349);
or U17224 (N_17224,N_12543,N_14977);
nor U17225 (N_17225,N_14093,N_14176);
and U17226 (N_17226,N_14591,N_14778);
or U17227 (N_17227,N_12683,N_12567);
nand U17228 (N_17228,N_10351,N_13292);
xnor U17229 (N_17229,N_11569,N_11243);
or U17230 (N_17230,N_13842,N_14580);
and U17231 (N_17231,N_11147,N_13573);
and U17232 (N_17232,N_11712,N_14607);
nand U17233 (N_17233,N_12348,N_11736);
or U17234 (N_17234,N_10093,N_10380);
or U17235 (N_17235,N_11176,N_14402);
xor U17236 (N_17236,N_13180,N_10391);
and U17237 (N_17237,N_10972,N_10239);
or U17238 (N_17238,N_13660,N_13107);
or U17239 (N_17239,N_12441,N_10149);
nand U17240 (N_17240,N_12848,N_11233);
nor U17241 (N_17241,N_11921,N_14514);
and U17242 (N_17242,N_14109,N_12943);
nand U17243 (N_17243,N_14452,N_10749);
nand U17244 (N_17244,N_13729,N_11126);
or U17245 (N_17245,N_14495,N_12180);
nand U17246 (N_17246,N_12430,N_12442);
and U17247 (N_17247,N_14551,N_13238);
and U17248 (N_17248,N_13314,N_12652);
nand U17249 (N_17249,N_13845,N_14618);
nor U17250 (N_17250,N_12575,N_14869);
or U17251 (N_17251,N_14061,N_13165);
nand U17252 (N_17252,N_11162,N_14410);
nor U17253 (N_17253,N_11392,N_13433);
nor U17254 (N_17254,N_13380,N_11501);
nand U17255 (N_17255,N_10823,N_12419);
or U17256 (N_17256,N_14893,N_11758);
nand U17257 (N_17257,N_10352,N_12820);
xnor U17258 (N_17258,N_11027,N_12075);
nand U17259 (N_17259,N_11687,N_12792);
nor U17260 (N_17260,N_13036,N_14291);
nand U17261 (N_17261,N_10026,N_11012);
or U17262 (N_17262,N_12496,N_11171);
nor U17263 (N_17263,N_13519,N_11832);
or U17264 (N_17264,N_13105,N_14705);
nand U17265 (N_17265,N_13829,N_13425);
nor U17266 (N_17266,N_10732,N_12532);
nor U17267 (N_17267,N_14783,N_11649);
and U17268 (N_17268,N_13941,N_11729);
xnor U17269 (N_17269,N_11901,N_14453);
nor U17270 (N_17270,N_10522,N_12531);
and U17271 (N_17271,N_12340,N_13128);
nand U17272 (N_17272,N_11990,N_10885);
and U17273 (N_17273,N_10694,N_11985);
xor U17274 (N_17274,N_12810,N_11167);
nand U17275 (N_17275,N_12000,N_14245);
and U17276 (N_17276,N_14920,N_13192);
or U17277 (N_17277,N_10606,N_10700);
or U17278 (N_17278,N_13557,N_13001);
or U17279 (N_17279,N_10246,N_14379);
and U17280 (N_17280,N_10546,N_14843);
and U17281 (N_17281,N_12084,N_11542);
nand U17282 (N_17282,N_12909,N_10661);
nand U17283 (N_17283,N_12415,N_10532);
nand U17284 (N_17284,N_12593,N_11967);
or U17285 (N_17285,N_11065,N_12127);
nor U17286 (N_17286,N_10839,N_14090);
or U17287 (N_17287,N_14532,N_10759);
nor U17288 (N_17288,N_14067,N_10640);
and U17289 (N_17289,N_14757,N_12052);
and U17290 (N_17290,N_14594,N_12517);
or U17291 (N_17291,N_10316,N_11105);
nand U17292 (N_17292,N_13027,N_10662);
nand U17293 (N_17293,N_10199,N_14946);
nand U17294 (N_17294,N_12808,N_10451);
nand U17295 (N_17295,N_11794,N_12168);
and U17296 (N_17296,N_12970,N_12747);
nand U17297 (N_17297,N_13132,N_12789);
or U17298 (N_17298,N_14924,N_13397);
and U17299 (N_17299,N_14071,N_12452);
xnor U17300 (N_17300,N_12318,N_12553);
or U17301 (N_17301,N_12029,N_14531);
nand U17302 (N_17302,N_14251,N_10253);
or U17303 (N_17303,N_14784,N_10252);
and U17304 (N_17304,N_11460,N_14558);
and U17305 (N_17305,N_12642,N_12152);
xor U17306 (N_17306,N_10878,N_13882);
or U17307 (N_17307,N_11410,N_13282);
and U17308 (N_17308,N_12277,N_12123);
and U17309 (N_17309,N_13992,N_13019);
or U17310 (N_17310,N_13948,N_14851);
nand U17311 (N_17311,N_13952,N_14032);
and U17312 (N_17312,N_13398,N_13626);
or U17313 (N_17313,N_12462,N_12259);
nor U17314 (N_17314,N_12386,N_14414);
nor U17315 (N_17315,N_14259,N_12945);
nand U17316 (N_17316,N_10995,N_14404);
and U17317 (N_17317,N_12121,N_12389);
and U17318 (N_17318,N_14494,N_11892);
or U17319 (N_17319,N_11324,N_13855);
and U17320 (N_17320,N_10573,N_14957);
nor U17321 (N_17321,N_13819,N_13360);
or U17322 (N_17322,N_12594,N_11363);
nor U17323 (N_17323,N_11616,N_11514);
nor U17324 (N_17324,N_14698,N_10138);
or U17325 (N_17325,N_13138,N_14039);
and U17326 (N_17326,N_10345,N_11961);
nor U17327 (N_17327,N_10934,N_14278);
and U17328 (N_17328,N_14692,N_13947);
nand U17329 (N_17329,N_11215,N_12681);
and U17330 (N_17330,N_10899,N_13277);
nor U17331 (N_17331,N_12812,N_14687);
nand U17332 (N_17332,N_10722,N_10454);
and U17333 (N_17333,N_12116,N_14133);
nor U17334 (N_17334,N_12767,N_10481);
or U17335 (N_17335,N_12752,N_14277);
and U17336 (N_17336,N_14112,N_12319);
nor U17337 (N_17337,N_11188,N_12074);
nor U17338 (N_17338,N_14915,N_11001);
xor U17339 (N_17339,N_12486,N_13438);
xor U17340 (N_17340,N_14860,N_11448);
and U17341 (N_17341,N_10294,N_12309);
nor U17342 (N_17342,N_14084,N_11763);
or U17343 (N_17343,N_12977,N_11769);
nand U17344 (N_17344,N_13455,N_10715);
and U17345 (N_17345,N_10978,N_13929);
or U17346 (N_17346,N_11759,N_12537);
or U17347 (N_17347,N_10645,N_14362);
nand U17348 (N_17348,N_11640,N_11183);
nand U17349 (N_17349,N_11236,N_14669);
or U17350 (N_17350,N_10507,N_10959);
or U17351 (N_17351,N_12599,N_14162);
xor U17352 (N_17352,N_11417,N_13889);
or U17353 (N_17353,N_14629,N_11158);
or U17354 (N_17354,N_10237,N_12119);
nor U17355 (N_17355,N_10695,N_11726);
or U17356 (N_17356,N_14319,N_13775);
or U17357 (N_17357,N_14197,N_11153);
and U17358 (N_17358,N_13517,N_14955);
nor U17359 (N_17359,N_13272,N_13813);
and U17360 (N_17360,N_10727,N_13118);
or U17361 (N_17361,N_14907,N_12218);
nor U17362 (N_17362,N_11132,N_13098);
nor U17363 (N_17363,N_11658,N_10519);
xor U17364 (N_17364,N_12223,N_12232);
or U17365 (N_17365,N_13931,N_12921);
nand U17366 (N_17366,N_14316,N_10010);
nand U17367 (N_17367,N_12954,N_14748);
nor U17368 (N_17368,N_11650,N_11385);
nand U17369 (N_17369,N_13823,N_14989);
or U17370 (N_17370,N_13451,N_14771);
nand U17371 (N_17371,N_13536,N_10704);
nor U17372 (N_17372,N_11646,N_14782);
and U17373 (N_17373,N_11826,N_12688);
or U17374 (N_17374,N_11610,N_11439);
and U17375 (N_17375,N_10457,N_11166);
or U17376 (N_17376,N_13323,N_10172);
nand U17377 (N_17377,N_10092,N_13332);
or U17378 (N_17378,N_10506,N_10786);
nand U17379 (N_17379,N_14088,N_10402);
and U17380 (N_17380,N_10131,N_14397);
and U17381 (N_17381,N_14821,N_11379);
and U17382 (N_17382,N_13237,N_10220);
and U17383 (N_17383,N_14817,N_11752);
or U17384 (N_17384,N_13552,N_12230);
or U17385 (N_17385,N_11931,N_10561);
or U17386 (N_17386,N_13541,N_14430);
nor U17387 (N_17387,N_11139,N_12739);
nand U17388 (N_17388,N_11248,N_13513);
nor U17389 (N_17389,N_14519,N_10980);
and U17390 (N_17390,N_14535,N_13088);
nand U17391 (N_17391,N_14530,N_10499);
nand U17392 (N_17392,N_12262,N_13136);
xnor U17393 (N_17393,N_10210,N_13331);
nand U17394 (N_17394,N_12187,N_14975);
nand U17395 (N_17395,N_12411,N_13859);
nor U17396 (N_17396,N_14512,N_13373);
xnor U17397 (N_17397,N_14395,N_10132);
and U17398 (N_17398,N_11853,N_13294);
and U17399 (N_17399,N_12154,N_12965);
and U17400 (N_17400,N_14582,N_11803);
and U17401 (N_17401,N_12629,N_14996);
and U17402 (N_17402,N_11449,N_11553);
nand U17403 (N_17403,N_14124,N_11784);
and U17404 (N_17404,N_14730,N_12563);
and U17405 (N_17405,N_10349,N_11817);
nor U17406 (N_17406,N_13672,N_12428);
or U17407 (N_17407,N_12561,N_11192);
and U17408 (N_17408,N_10807,N_14359);
nand U17409 (N_17409,N_14089,N_14462);
xor U17410 (N_17410,N_13190,N_11297);
nor U17411 (N_17411,N_11217,N_13145);
nor U17412 (N_17412,N_13392,N_12285);
nand U17413 (N_17413,N_13298,N_14465);
or U17414 (N_17414,N_10736,N_12225);
nor U17415 (N_17415,N_12917,N_12877);
xnor U17416 (N_17416,N_11733,N_14375);
or U17417 (N_17417,N_14509,N_12310);
nor U17418 (N_17418,N_11588,N_14454);
or U17419 (N_17419,N_11909,N_13979);
xor U17420 (N_17420,N_13198,N_11485);
nand U17421 (N_17421,N_13966,N_14651);
and U17422 (N_17422,N_13412,N_11250);
or U17423 (N_17423,N_12822,N_12578);
and U17424 (N_17424,N_14244,N_10297);
nor U17425 (N_17425,N_11022,N_10846);
nor U17426 (N_17426,N_12007,N_11504);
and U17427 (N_17427,N_13674,N_13137);
nand U17428 (N_17428,N_11422,N_13640);
and U17429 (N_17429,N_10062,N_12703);
and U17430 (N_17430,N_12151,N_11476);
nand U17431 (N_17431,N_10947,N_13600);
nand U17432 (N_17432,N_14732,N_14488);
or U17433 (N_17433,N_13673,N_12610);
nor U17434 (N_17434,N_12317,N_10425);
or U17435 (N_17435,N_12353,N_13434);
or U17436 (N_17436,N_14526,N_13096);
nor U17437 (N_17437,N_14791,N_10224);
and U17438 (N_17438,N_11801,N_14372);
and U17439 (N_17439,N_11128,N_13485);
or U17440 (N_17440,N_11963,N_14275);
nor U17441 (N_17441,N_14995,N_14418);
nor U17442 (N_17442,N_11081,N_14750);
nand U17443 (N_17443,N_10195,N_11025);
nand U17444 (N_17444,N_14555,N_12006);
nand U17445 (N_17445,N_13148,N_12903);
nor U17446 (N_17446,N_13127,N_14213);
or U17447 (N_17447,N_14951,N_11804);
and U17448 (N_17448,N_14945,N_14242);
xor U17449 (N_17449,N_11936,N_11424);
and U17450 (N_17450,N_13639,N_14792);
nand U17451 (N_17451,N_10289,N_11523);
and U17452 (N_17452,N_12604,N_10206);
or U17453 (N_17453,N_13946,N_13212);
nand U17454 (N_17454,N_12998,N_14592);
and U17455 (N_17455,N_14615,N_14659);
xor U17456 (N_17456,N_12206,N_12748);
nor U17457 (N_17457,N_14952,N_13099);
or U17458 (N_17458,N_13604,N_12899);
nor U17459 (N_17459,N_13028,N_14457);
xnor U17460 (N_17460,N_12189,N_13973);
nor U17461 (N_17461,N_14119,N_13320);
and U17462 (N_17462,N_10382,N_13618);
and U17463 (N_17463,N_14520,N_13053);
nand U17464 (N_17464,N_13625,N_10484);
nand U17465 (N_17465,N_14332,N_12170);
nand U17466 (N_17466,N_14173,N_10443);
and U17467 (N_17467,N_13971,N_10698);
or U17468 (N_17468,N_12850,N_10346);
xnor U17469 (N_17469,N_10490,N_13073);
or U17470 (N_17470,N_12915,N_11877);
nand U17471 (N_17471,N_12439,N_12182);
nand U17472 (N_17472,N_11168,N_12315);
nand U17473 (N_17473,N_11059,N_12960);
nand U17474 (N_17474,N_14720,N_11296);
nor U17475 (N_17475,N_12234,N_11218);
nor U17476 (N_17476,N_11195,N_11533);
xnor U17477 (N_17477,N_11577,N_11720);
nand U17478 (N_17478,N_11329,N_13388);
xnor U17479 (N_17479,N_10372,N_12100);
nor U17480 (N_17480,N_14429,N_12399);
or U17481 (N_17481,N_14334,N_14827);
nor U17482 (N_17482,N_12674,N_11314);
or U17483 (N_17483,N_12190,N_10530);
nand U17484 (N_17484,N_12529,N_10310);
and U17485 (N_17485,N_12175,N_14019);
nor U17486 (N_17486,N_12840,N_10438);
or U17487 (N_17487,N_14697,N_10011);
or U17488 (N_17488,N_14191,N_11150);
nor U17489 (N_17489,N_12648,N_14832);
or U17490 (N_17490,N_12997,N_14051);
nor U17491 (N_17491,N_11777,N_14107);
nand U17492 (N_17492,N_11052,N_11761);
or U17493 (N_17493,N_13875,N_11352);
xnor U17494 (N_17494,N_11011,N_14060);
and U17495 (N_17495,N_12482,N_11904);
or U17496 (N_17496,N_11984,N_13351);
or U17497 (N_17497,N_12060,N_11618);
nor U17498 (N_17498,N_14855,N_13354);
nor U17499 (N_17499,N_13305,N_11740);
and U17500 (N_17500,N_13447,N_11360);
and U17501 (N_17501,N_14732,N_10767);
nand U17502 (N_17502,N_12893,N_14236);
nand U17503 (N_17503,N_12024,N_10728);
and U17504 (N_17504,N_10011,N_14341);
nor U17505 (N_17505,N_14023,N_13678);
nand U17506 (N_17506,N_14903,N_13015);
nor U17507 (N_17507,N_11062,N_11193);
or U17508 (N_17508,N_11777,N_11130);
and U17509 (N_17509,N_12270,N_13788);
or U17510 (N_17510,N_11771,N_13893);
nand U17511 (N_17511,N_11251,N_11540);
nor U17512 (N_17512,N_10254,N_11206);
and U17513 (N_17513,N_12971,N_10403);
nand U17514 (N_17514,N_11967,N_13378);
nor U17515 (N_17515,N_10421,N_11428);
or U17516 (N_17516,N_11971,N_10240);
nor U17517 (N_17517,N_13421,N_10565);
nor U17518 (N_17518,N_11171,N_12223);
nor U17519 (N_17519,N_13440,N_11029);
nand U17520 (N_17520,N_11996,N_11703);
or U17521 (N_17521,N_11290,N_12277);
and U17522 (N_17522,N_10571,N_12029);
nor U17523 (N_17523,N_12776,N_13693);
or U17524 (N_17524,N_14001,N_11699);
or U17525 (N_17525,N_11702,N_13479);
or U17526 (N_17526,N_10820,N_13202);
nand U17527 (N_17527,N_13165,N_13669);
or U17528 (N_17528,N_10730,N_13260);
and U17529 (N_17529,N_13944,N_13421);
xnor U17530 (N_17530,N_12287,N_12209);
or U17531 (N_17531,N_12949,N_13360);
xor U17532 (N_17532,N_11635,N_10479);
or U17533 (N_17533,N_12105,N_12689);
nand U17534 (N_17534,N_13433,N_10091);
nand U17535 (N_17535,N_13024,N_14244);
and U17536 (N_17536,N_11349,N_13158);
and U17537 (N_17537,N_10640,N_14064);
nor U17538 (N_17538,N_11818,N_11067);
or U17539 (N_17539,N_11593,N_10414);
and U17540 (N_17540,N_13847,N_12118);
or U17541 (N_17541,N_11108,N_11937);
and U17542 (N_17542,N_14440,N_10504);
or U17543 (N_17543,N_13042,N_14116);
nand U17544 (N_17544,N_12584,N_14929);
or U17545 (N_17545,N_12207,N_10575);
nor U17546 (N_17546,N_10508,N_13368);
and U17547 (N_17547,N_11272,N_13840);
and U17548 (N_17548,N_12398,N_13973);
and U17549 (N_17549,N_10770,N_12643);
and U17550 (N_17550,N_12763,N_12802);
nand U17551 (N_17551,N_10239,N_12904);
nand U17552 (N_17552,N_12289,N_12547);
xor U17553 (N_17553,N_11589,N_14678);
and U17554 (N_17554,N_13819,N_11284);
or U17555 (N_17555,N_10160,N_14466);
nor U17556 (N_17556,N_14021,N_10611);
or U17557 (N_17557,N_13158,N_13782);
nand U17558 (N_17558,N_10164,N_11126);
nor U17559 (N_17559,N_12189,N_11637);
or U17560 (N_17560,N_10822,N_13085);
or U17561 (N_17561,N_10853,N_12319);
nor U17562 (N_17562,N_13027,N_12673);
nand U17563 (N_17563,N_13606,N_10347);
nor U17564 (N_17564,N_12276,N_11203);
and U17565 (N_17565,N_12966,N_10407);
nand U17566 (N_17566,N_10120,N_11207);
nand U17567 (N_17567,N_12258,N_14467);
nor U17568 (N_17568,N_10703,N_13661);
nand U17569 (N_17569,N_13974,N_13219);
nand U17570 (N_17570,N_10613,N_12346);
nand U17571 (N_17571,N_14344,N_14791);
or U17572 (N_17572,N_13063,N_10697);
or U17573 (N_17573,N_11483,N_13323);
or U17574 (N_17574,N_10063,N_11480);
or U17575 (N_17575,N_12227,N_11918);
nor U17576 (N_17576,N_12948,N_12609);
nand U17577 (N_17577,N_10941,N_11473);
nand U17578 (N_17578,N_12452,N_13098);
nor U17579 (N_17579,N_13941,N_13807);
nor U17580 (N_17580,N_14306,N_10420);
nor U17581 (N_17581,N_10774,N_12862);
or U17582 (N_17582,N_11098,N_12303);
nor U17583 (N_17583,N_11311,N_11505);
nor U17584 (N_17584,N_10877,N_10147);
nor U17585 (N_17585,N_13173,N_10018);
and U17586 (N_17586,N_14396,N_11210);
nor U17587 (N_17587,N_14517,N_11362);
nor U17588 (N_17588,N_10485,N_14853);
or U17589 (N_17589,N_14579,N_12248);
or U17590 (N_17590,N_13952,N_11163);
and U17591 (N_17591,N_10240,N_10468);
nor U17592 (N_17592,N_13837,N_11981);
or U17593 (N_17593,N_10906,N_13961);
nor U17594 (N_17594,N_14805,N_12929);
and U17595 (N_17595,N_11034,N_10337);
or U17596 (N_17596,N_10043,N_10770);
nand U17597 (N_17597,N_10952,N_12745);
nor U17598 (N_17598,N_12745,N_12491);
and U17599 (N_17599,N_12408,N_14953);
or U17600 (N_17600,N_13143,N_10885);
nor U17601 (N_17601,N_13673,N_14292);
or U17602 (N_17602,N_13343,N_10074);
xnor U17603 (N_17603,N_11855,N_12107);
nor U17604 (N_17604,N_11311,N_14290);
and U17605 (N_17605,N_10628,N_10081);
nor U17606 (N_17606,N_14754,N_12745);
nand U17607 (N_17607,N_12671,N_14125);
and U17608 (N_17608,N_14254,N_12783);
or U17609 (N_17609,N_14951,N_11778);
nor U17610 (N_17610,N_13333,N_10586);
and U17611 (N_17611,N_13385,N_14521);
nor U17612 (N_17612,N_13252,N_13550);
or U17613 (N_17613,N_14572,N_10052);
and U17614 (N_17614,N_10855,N_13186);
xnor U17615 (N_17615,N_14204,N_14248);
nor U17616 (N_17616,N_13889,N_11866);
nand U17617 (N_17617,N_12062,N_13226);
nand U17618 (N_17618,N_12830,N_13344);
or U17619 (N_17619,N_12666,N_12094);
nor U17620 (N_17620,N_12246,N_14212);
and U17621 (N_17621,N_13878,N_12889);
or U17622 (N_17622,N_14220,N_13163);
nand U17623 (N_17623,N_12004,N_11779);
or U17624 (N_17624,N_10085,N_12477);
nand U17625 (N_17625,N_12447,N_12817);
nor U17626 (N_17626,N_11362,N_13213);
xnor U17627 (N_17627,N_14724,N_11883);
nor U17628 (N_17628,N_12910,N_11429);
or U17629 (N_17629,N_13603,N_13045);
nor U17630 (N_17630,N_13482,N_12630);
xnor U17631 (N_17631,N_14150,N_14022);
or U17632 (N_17632,N_12862,N_11540);
or U17633 (N_17633,N_12412,N_12512);
nand U17634 (N_17634,N_14022,N_11986);
and U17635 (N_17635,N_14136,N_14293);
nand U17636 (N_17636,N_11896,N_10590);
nand U17637 (N_17637,N_10908,N_13426);
and U17638 (N_17638,N_13204,N_12533);
nand U17639 (N_17639,N_14864,N_12920);
xnor U17640 (N_17640,N_10613,N_13132);
and U17641 (N_17641,N_12517,N_13666);
nand U17642 (N_17642,N_14891,N_13175);
or U17643 (N_17643,N_14424,N_10659);
and U17644 (N_17644,N_10575,N_12586);
nor U17645 (N_17645,N_14415,N_11708);
xnor U17646 (N_17646,N_10985,N_11561);
and U17647 (N_17647,N_10168,N_10066);
and U17648 (N_17648,N_11510,N_11588);
or U17649 (N_17649,N_14893,N_11688);
nand U17650 (N_17650,N_12115,N_10238);
or U17651 (N_17651,N_10408,N_12778);
xnor U17652 (N_17652,N_14085,N_12836);
or U17653 (N_17653,N_10048,N_10172);
and U17654 (N_17654,N_12293,N_12740);
nand U17655 (N_17655,N_13167,N_11587);
or U17656 (N_17656,N_10467,N_10460);
nand U17657 (N_17657,N_14169,N_12498);
nand U17658 (N_17658,N_14783,N_14706);
and U17659 (N_17659,N_12871,N_12063);
or U17660 (N_17660,N_10792,N_14084);
nand U17661 (N_17661,N_10611,N_14938);
and U17662 (N_17662,N_13471,N_14062);
nor U17663 (N_17663,N_11241,N_13323);
or U17664 (N_17664,N_10361,N_14582);
or U17665 (N_17665,N_10475,N_12422);
or U17666 (N_17666,N_11623,N_13534);
and U17667 (N_17667,N_11285,N_10763);
and U17668 (N_17668,N_13485,N_11734);
or U17669 (N_17669,N_13595,N_13738);
nand U17670 (N_17670,N_12836,N_10271);
or U17671 (N_17671,N_10721,N_12835);
nand U17672 (N_17672,N_10857,N_13873);
or U17673 (N_17673,N_11748,N_13907);
and U17674 (N_17674,N_14480,N_10269);
nand U17675 (N_17675,N_10280,N_10462);
nand U17676 (N_17676,N_13320,N_11764);
nand U17677 (N_17677,N_12552,N_13035);
nor U17678 (N_17678,N_11298,N_14980);
nand U17679 (N_17679,N_11662,N_10389);
nor U17680 (N_17680,N_12183,N_12028);
nor U17681 (N_17681,N_13950,N_11896);
xor U17682 (N_17682,N_11938,N_14158);
xor U17683 (N_17683,N_11409,N_10022);
or U17684 (N_17684,N_11549,N_12429);
nand U17685 (N_17685,N_13976,N_12965);
xor U17686 (N_17686,N_10162,N_12643);
or U17687 (N_17687,N_11400,N_14794);
xor U17688 (N_17688,N_10394,N_11452);
nor U17689 (N_17689,N_12961,N_12278);
nor U17690 (N_17690,N_13752,N_12729);
and U17691 (N_17691,N_11309,N_10845);
xnor U17692 (N_17692,N_13903,N_10694);
or U17693 (N_17693,N_13943,N_10495);
or U17694 (N_17694,N_13308,N_12709);
and U17695 (N_17695,N_11726,N_11535);
nand U17696 (N_17696,N_12539,N_11318);
or U17697 (N_17697,N_10405,N_10562);
xnor U17698 (N_17698,N_13257,N_12503);
or U17699 (N_17699,N_12453,N_13580);
or U17700 (N_17700,N_13583,N_10767);
and U17701 (N_17701,N_13042,N_12829);
or U17702 (N_17702,N_12629,N_10977);
nand U17703 (N_17703,N_12152,N_13865);
and U17704 (N_17704,N_14932,N_13503);
nor U17705 (N_17705,N_10903,N_12636);
and U17706 (N_17706,N_11341,N_12382);
nand U17707 (N_17707,N_14608,N_14871);
nor U17708 (N_17708,N_10746,N_11306);
or U17709 (N_17709,N_13675,N_14881);
nor U17710 (N_17710,N_13292,N_14424);
and U17711 (N_17711,N_13954,N_10001);
nand U17712 (N_17712,N_12337,N_12408);
nand U17713 (N_17713,N_12658,N_12327);
and U17714 (N_17714,N_14990,N_14128);
xor U17715 (N_17715,N_13871,N_13601);
and U17716 (N_17716,N_10250,N_10104);
xor U17717 (N_17717,N_14063,N_13210);
nand U17718 (N_17718,N_13833,N_11858);
nor U17719 (N_17719,N_14539,N_10290);
and U17720 (N_17720,N_14900,N_11233);
nand U17721 (N_17721,N_13234,N_14898);
nor U17722 (N_17722,N_12278,N_14236);
xnor U17723 (N_17723,N_13582,N_14468);
nand U17724 (N_17724,N_11344,N_13624);
nor U17725 (N_17725,N_11808,N_11305);
nor U17726 (N_17726,N_14480,N_11182);
xor U17727 (N_17727,N_13167,N_14869);
and U17728 (N_17728,N_14779,N_14162);
or U17729 (N_17729,N_14447,N_12597);
and U17730 (N_17730,N_10802,N_10118);
nand U17731 (N_17731,N_10547,N_10644);
or U17732 (N_17732,N_12894,N_14075);
and U17733 (N_17733,N_10903,N_12446);
and U17734 (N_17734,N_12048,N_10228);
or U17735 (N_17735,N_14126,N_13814);
nor U17736 (N_17736,N_11103,N_10321);
and U17737 (N_17737,N_12376,N_13865);
nand U17738 (N_17738,N_14918,N_14006);
nand U17739 (N_17739,N_11576,N_13493);
and U17740 (N_17740,N_13955,N_11946);
and U17741 (N_17741,N_12049,N_13845);
nand U17742 (N_17742,N_14326,N_14068);
and U17743 (N_17743,N_14923,N_12369);
xor U17744 (N_17744,N_10700,N_14335);
nand U17745 (N_17745,N_14227,N_12163);
or U17746 (N_17746,N_11946,N_12012);
or U17747 (N_17747,N_12899,N_10930);
and U17748 (N_17748,N_14981,N_10085);
nand U17749 (N_17749,N_11866,N_13805);
xnor U17750 (N_17750,N_11634,N_13495);
and U17751 (N_17751,N_14069,N_12427);
xnor U17752 (N_17752,N_14655,N_14423);
nor U17753 (N_17753,N_11346,N_11087);
and U17754 (N_17754,N_14748,N_14872);
or U17755 (N_17755,N_14139,N_13666);
nor U17756 (N_17756,N_12304,N_14789);
or U17757 (N_17757,N_11923,N_11184);
and U17758 (N_17758,N_10519,N_13726);
or U17759 (N_17759,N_11294,N_14118);
nand U17760 (N_17760,N_11620,N_13170);
nor U17761 (N_17761,N_13282,N_10308);
nand U17762 (N_17762,N_12675,N_12228);
nand U17763 (N_17763,N_13800,N_11190);
and U17764 (N_17764,N_13740,N_10060);
xor U17765 (N_17765,N_14061,N_10856);
xnor U17766 (N_17766,N_11035,N_14334);
or U17767 (N_17767,N_13821,N_10864);
nand U17768 (N_17768,N_11650,N_11734);
and U17769 (N_17769,N_14519,N_13460);
or U17770 (N_17770,N_14411,N_13237);
nand U17771 (N_17771,N_14841,N_12653);
nand U17772 (N_17772,N_13834,N_10447);
nand U17773 (N_17773,N_13056,N_14184);
and U17774 (N_17774,N_12297,N_10630);
nor U17775 (N_17775,N_11181,N_10332);
nor U17776 (N_17776,N_12210,N_10962);
and U17777 (N_17777,N_12180,N_14208);
or U17778 (N_17778,N_14871,N_14527);
nor U17779 (N_17779,N_10978,N_12639);
or U17780 (N_17780,N_12218,N_11248);
and U17781 (N_17781,N_14709,N_12484);
xnor U17782 (N_17782,N_11344,N_10536);
and U17783 (N_17783,N_10991,N_12573);
or U17784 (N_17784,N_14283,N_13879);
and U17785 (N_17785,N_10380,N_13522);
and U17786 (N_17786,N_12290,N_12942);
or U17787 (N_17787,N_13533,N_13942);
nor U17788 (N_17788,N_14236,N_14936);
or U17789 (N_17789,N_14911,N_12233);
nor U17790 (N_17790,N_11925,N_14768);
nor U17791 (N_17791,N_11880,N_10273);
nor U17792 (N_17792,N_11352,N_14013);
and U17793 (N_17793,N_12151,N_11004);
nand U17794 (N_17794,N_11620,N_13321);
nand U17795 (N_17795,N_12120,N_12341);
or U17796 (N_17796,N_11490,N_10037);
xnor U17797 (N_17797,N_11046,N_12503);
nand U17798 (N_17798,N_11449,N_10055);
nand U17799 (N_17799,N_10361,N_14677);
or U17800 (N_17800,N_14785,N_13559);
nand U17801 (N_17801,N_13969,N_14639);
nor U17802 (N_17802,N_13170,N_13571);
and U17803 (N_17803,N_14992,N_11514);
nand U17804 (N_17804,N_10184,N_13636);
nor U17805 (N_17805,N_14056,N_12240);
and U17806 (N_17806,N_13864,N_11927);
nor U17807 (N_17807,N_14496,N_11262);
nand U17808 (N_17808,N_11300,N_14951);
nand U17809 (N_17809,N_11606,N_10396);
nor U17810 (N_17810,N_12775,N_10712);
nor U17811 (N_17811,N_10569,N_12619);
nor U17812 (N_17812,N_11163,N_11292);
nand U17813 (N_17813,N_12043,N_11594);
or U17814 (N_17814,N_12150,N_10872);
or U17815 (N_17815,N_11966,N_14136);
nand U17816 (N_17816,N_12573,N_11697);
or U17817 (N_17817,N_14085,N_11684);
and U17818 (N_17818,N_10182,N_13979);
nand U17819 (N_17819,N_14956,N_14368);
nor U17820 (N_17820,N_12837,N_12640);
or U17821 (N_17821,N_12759,N_13866);
nand U17822 (N_17822,N_10182,N_11057);
and U17823 (N_17823,N_11697,N_14974);
and U17824 (N_17824,N_10262,N_13122);
and U17825 (N_17825,N_14225,N_10684);
xor U17826 (N_17826,N_14257,N_11237);
or U17827 (N_17827,N_11351,N_14152);
nor U17828 (N_17828,N_13000,N_12187);
or U17829 (N_17829,N_12429,N_13414);
xnor U17830 (N_17830,N_11942,N_14747);
or U17831 (N_17831,N_14113,N_13134);
nor U17832 (N_17832,N_10356,N_11795);
nand U17833 (N_17833,N_14873,N_13938);
or U17834 (N_17834,N_11856,N_12852);
xor U17835 (N_17835,N_14437,N_14521);
and U17836 (N_17836,N_14256,N_12176);
nor U17837 (N_17837,N_11252,N_13707);
nor U17838 (N_17838,N_12433,N_10414);
xor U17839 (N_17839,N_11257,N_13791);
nand U17840 (N_17840,N_13840,N_13383);
or U17841 (N_17841,N_10833,N_13595);
or U17842 (N_17842,N_11599,N_11192);
xnor U17843 (N_17843,N_10715,N_11694);
nor U17844 (N_17844,N_12804,N_12258);
xor U17845 (N_17845,N_12995,N_13987);
or U17846 (N_17846,N_11474,N_13565);
nand U17847 (N_17847,N_12307,N_10204);
xnor U17848 (N_17848,N_11760,N_13461);
nor U17849 (N_17849,N_10636,N_13252);
nand U17850 (N_17850,N_10558,N_14563);
nand U17851 (N_17851,N_14758,N_10983);
or U17852 (N_17852,N_10678,N_13189);
xor U17853 (N_17853,N_14071,N_11466);
nor U17854 (N_17854,N_14564,N_12656);
xor U17855 (N_17855,N_10987,N_13885);
nor U17856 (N_17856,N_10482,N_13251);
nor U17857 (N_17857,N_13503,N_13108);
nor U17858 (N_17858,N_13802,N_12387);
xnor U17859 (N_17859,N_11993,N_14983);
nand U17860 (N_17860,N_12696,N_14290);
nand U17861 (N_17861,N_14089,N_10285);
nand U17862 (N_17862,N_14747,N_10962);
or U17863 (N_17863,N_10515,N_10358);
and U17864 (N_17864,N_12552,N_13366);
nand U17865 (N_17865,N_10530,N_13356);
nand U17866 (N_17866,N_11049,N_12931);
and U17867 (N_17867,N_13748,N_14878);
and U17868 (N_17868,N_14708,N_13753);
nand U17869 (N_17869,N_12834,N_13883);
nand U17870 (N_17870,N_10686,N_13729);
and U17871 (N_17871,N_11645,N_13485);
nand U17872 (N_17872,N_11611,N_13151);
and U17873 (N_17873,N_11699,N_11703);
and U17874 (N_17874,N_11708,N_12197);
nor U17875 (N_17875,N_10911,N_14896);
or U17876 (N_17876,N_13085,N_10780);
nand U17877 (N_17877,N_10352,N_12550);
and U17878 (N_17878,N_12403,N_12597);
or U17879 (N_17879,N_14028,N_10148);
or U17880 (N_17880,N_14010,N_14450);
or U17881 (N_17881,N_10059,N_13515);
or U17882 (N_17882,N_10675,N_12559);
and U17883 (N_17883,N_10539,N_10794);
nand U17884 (N_17884,N_11202,N_11547);
nor U17885 (N_17885,N_12320,N_14530);
nor U17886 (N_17886,N_12254,N_11724);
nor U17887 (N_17887,N_13625,N_10632);
xor U17888 (N_17888,N_14131,N_14408);
nand U17889 (N_17889,N_10712,N_13334);
and U17890 (N_17890,N_11675,N_14988);
nand U17891 (N_17891,N_14747,N_11937);
or U17892 (N_17892,N_10110,N_12874);
or U17893 (N_17893,N_14522,N_11707);
nand U17894 (N_17894,N_12468,N_10636);
xor U17895 (N_17895,N_13894,N_12957);
and U17896 (N_17896,N_10977,N_13188);
or U17897 (N_17897,N_11058,N_10134);
and U17898 (N_17898,N_12028,N_10611);
nand U17899 (N_17899,N_12944,N_11264);
and U17900 (N_17900,N_10886,N_10651);
nor U17901 (N_17901,N_13221,N_12437);
and U17902 (N_17902,N_14066,N_10490);
or U17903 (N_17903,N_11435,N_11969);
and U17904 (N_17904,N_13055,N_13778);
nand U17905 (N_17905,N_11995,N_12084);
nand U17906 (N_17906,N_11781,N_14202);
nor U17907 (N_17907,N_13160,N_12647);
or U17908 (N_17908,N_11633,N_14413);
nor U17909 (N_17909,N_12566,N_11756);
nor U17910 (N_17910,N_12452,N_12915);
or U17911 (N_17911,N_14969,N_10961);
and U17912 (N_17912,N_13159,N_14658);
or U17913 (N_17913,N_14305,N_13403);
and U17914 (N_17914,N_14282,N_12130);
or U17915 (N_17915,N_11265,N_12410);
nor U17916 (N_17916,N_13551,N_10809);
nor U17917 (N_17917,N_11268,N_10358);
or U17918 (N_17918,N_14396,N_13363);
or U17919 (N_17919,N_12719,N_11538);
nand U17920 (N_17920,N_12593,N_11149);
nand U17921 (N_17921,N_10500,N_12748);
and U17922 (N_17922,N_12273,N_10545);
nor U17923 (N_17923,N_11162,N_14152);
and U17924 (N_17924,N_11565,N_14617);
or U17925 (N_17925,N_12046,N_10516);
or U17926 (N_17926,N_13708,N_10704);
or U17927 (N_17927,N_14041,N_10339);
nor U17928 (N_17928,N_14446,N_14633);
or U17929 (N_17929,N_13478,N_13560);
nor U17930 (N_17930,N_14643,N_12070);
xnor U17931 (N_17931,N_11159,N_12483);
xor U17932 (N_17932,N_10570,N_10779);
nor U17933 (N_17933,N_11339,N_12602);
or U17934 (N_17934,N_13668,N_11175);
nand U17935 (N_17935,N_11957,N_11699);
or U17936 (N_17936,N_11266,N_13345);
xnor U17937 (N_17937,N_10558,N_11849);
and U17938 (N_17938,N_12653,N_13214);
nor U17939 (N_17939,N_12961,N_10940);
xor U17940 (N_17940,N_12745,N_12939);
or U17941 (N_17941,N_12408,N_11731);
xor U17942 (N_17942,N_12408,N_12530);
nor U17943 (N_17943,N_14798,N_13884);
nor U17944 (N_17944,N_10593,N_14061);
and U17945 (N_17945,N_11076,N_14168);
or U17946 (N_17946,N_10108,N_13626);
nand U17947 (N_17947,N_13891,N_11099);
and U17948 (N_17948,N_11689,N_10427);
nand U17949 (N_17949,N_14430,N_12942);
nor U17950 (N_17950,N_10752,N_10419);
or U17951 (N_17951,N_13874,N_11547);
and U17952 (N_17952,N_10120,N_14592);
nor U17953 (N_17953,N_11990,N_13677);
nand U17954 (N_17954,N_10358,N_10470);
nor U17955 (N_17955,N_11411,N_13786);
nor U17956 (N_17956,N_12656,N_12396);
nand U17957 (N_17957,N_10223,N_10153);
or U17958 (N_17958,N_12248,N_12332);
nor U17959 (N_17959,N_11307,N_11244);
or U17960 (N_17960,N_13228,N_11635);
nor U17961 (N_17961,N_13442,N_10688);
and U17962 (N_17962,N_14120,N_13660);
xor U17963 (N_17963,N_12649,N_10677);
nand U17964 (N_17964,N_10128,N_13915);
nand U17965 (N_17965,N_12974,N_13507);
nor U17966 (N_17966,N_13256,N_11063);
or U17967 (N_17967,N_14705,N_13529);
and U17968 (N_17968,N_10424,N_10438);
xor U17969 (N_17969,N_13370,N_11980);
nor U17970 (N_17970,N_12910,N_11374);
and U17971 (N_17971,N_12428,N_12794);
nor U17972 (N_17972,N_12973,N_13868);
or U17973 (N_17973,N_12372,N_11463);
and U17974 (N_17974,N_10868,N_12536);
nand U17975 (N_17975,N_11586,N_12136);
or U17976 (N_17976,N_13121,N_10687);
xnor U17977 (N_17977,N_14855,N_14164);
and U17978 (N_17978,N_10091,N_11610);
or U17979 (N_17979,N_12661,N_12724);
nor U17980 (N_17980,N_12166,N_11609);
nand U17981 (N_17981,N_13417,N_14192);
or U17982 (N_17982,N_14918,N_12343);
and U17983 (N_17983,N_12303,N_13352);
nand U17984 (N_17984,N_10051,N_14520);
or U17985 (N_17985,N_12343,N_14245);
nor U17986 (N_17986,N_11787,N_10012);
and U17987 (N_17987,N_13886,N_11658);
and U17988 (N_17988,N_10757,N_14694);
nor U17989 (N_17989,N_13151,N_10920);
nand U17990 (N_17990,N_14254,N_13584);
or U17991 (N_17991,N_13837,N_12044);
xnor U17992 (N_17992,N_12601,N_11693);
nor U17993 (N_17993,N_11759,N_10042);
or U17994 (N_17994,N_10127,N_14165);
or U17995 (N_17995,N_11160,N_14176);
and U17996 (N_17996,N_11533,N_11861);
and U17997 (N_17997,N_14588,N_12842);
nor U17998 (N_17998,N_10772,N_14628);
and U17999 (N_17999,N_14264,N_14075);
or U18000 (N_18000,N_14828,N_13300);
nand U18001 (N_18001,N_13003,N_13385);
xor U18002 (N_18002,N_10434,N_11580);
nor U18003 (N_18003,N_13046,N_13956);
and U18004 (N_18004,N_12507,N_12107);
nand U18005 (N_18005,N_14846,N_13168);
xnor U18006 (N_18006,N_11520,N_12757);
or U18007 (N_18007,N_14480,N_13601);
and U18008 (N_18008,N_13420,N_10137);
nor U18009 (N_18009,N_11427,N_13921);
nand U18010 (N_18010,N_11891,N_12732);
or U18011 (N_18011,N_12892,N_13172);
and U18012 (N_18012,N_14000,N_13802);
nor U18013 (N_18013,N_14569,N_10375);
or U18014 (N_18014,N_13383,N_13453);
and U18015 (N_18015,N_13740,N_14140);
nor U18016 (N_18016,N_13323,N_14423);
and U18017 (N_18017,N_14208,N_14377);
or U18018 (N_18018,N_10272,N_10994);
and U18019 (N_18019,N_10483,N_13756);
and U18020 (N_18020,N_14239,N_13854);
or U18021 (N_18021,N_13932,N_13505);
or U18022 (N_18022,N_13518,N_13870);
nand U18023 (N_18023,N_12071,N_14872);
nand U18024 (N_18024,N_12968,N_11347);
and U18025 (N_18025,N_13235,N_10719);
and U18026 (N_18026,N_13483,N_14720);
or U18027 (N_18027,N_12818,N_13519);
nor U18028 (N_18028,N_11321,N_11704);
nor U18029 (N_18029,N_11221,N_13502);
and U18030 (N_18030,N_13869,N_13228);
nor U18031 (N_18031,N_12129,N_14940);
nor U18032 (N_18032,N_11647,N_12689);
xnor U18033 (N_18033,N_12757,N_11135);
nor U18034 (N_18034,N_14315,N_14984);
and U18035 (N_18035,N_10087,N_12617);
and U18036 (N_18036,N_11463,N_11866);
nand U18037 (N_18037,N_11357,N_13650);
nand U18038 (N_18038,N_10784,N_12868);
nand U18039 (N_18039,N_13420,N_10752);
nand U18040 (N_18040,N_11082,N_10821);
and U18041 (N_18041,N_14894,N_10973);
nor U18042 (N_18042,N_10388,N_11748);
or U18043 (N_18043,N_11351,N_14959);
and U18044 (N_18044,N_13601,N_10155);
and U18045 (N_18045,N_13220,N_11223);
nand U18046 (N_18046,N_13909,N_12373);
or U18047 (N_18047,N_14065,N_11556);
or U18048 (N_18048,N_10575,N_12096);
and U18049 (N_18049,N_13744,N_10728);
and U18050 (N_18050,N_12038,N_12329);
nand U18051 (N_18051,N_14311,N_11693);
nand U18052 (N_18052,N_14332,N_14984);
and U18053 (N_18053,N_13287,N_10536);
xor U18054 (N_18054,N_14849,N_14838);
nor U18055 (N_18055,N_10301,N_12902);
nor U18056 (N_18056,N_11662,N_12222);
and U18057 (N_18057,N_14127,N_14242);
or U18058 (N_18058,N_10527,N_10431);
xor U18059 (N_18059,N_12096,N_13178);
nand U18060 (N_18060,N_10281,N_13768);
xnor U18061 (N_18061,N_10433,N_10878);
nand U18062 (N_18062,N_10999,N_13446);
xnor U18063 (N_18063,N_14050,N_12911);
nor U18064 (N_18064,N_10688,N_10546);
nor U18065 (N_18065,N_13382,N_11007);
xor U18066 (N_18066,N_10997,N_10093);
or U18067 (N_18067,N_10499,N_13843);
nand U18068 (N_18068,N_12724,N_13381);
xnor U18069 (N_18069,N_12996,N_11477);
and U18070 (N_18070,N_10413,N_12435);
nor U18071 (N_18071,N_10646,N_10113);
nand U18072 (N_18072,N_11550,N_14533);
nor U18073 (N_18073,N_10785,N_13501);
nor U18074 (N_18074,N_10688,N_14517);
and U18075 (N_18075,N_12063,N_13285);
and U18076 (N_18076,N_12693,N_11869);
nor U18077 (N_18077,N_10096,N_12194);
nor U18078 (N_18078,N_13102,N_12223);
and U18079 (N_18079,N_11799,N_13535);
xnor U18080 (N_18080,N_14687,N_10818);
nand U18081 (N_18081,N_14956,N_13944);
nor U18082 (N_18082,N_12652,N_14381);
nand U18083 (N_18083,N_13424,N_11134);
or U18084 (N_18084,N_13709,N_10950);
nor U18085 (N_18085,N_10811,N_11576);
and U18086 (N_18086,N_14234,N_13529);
or U18087 (N_18087,N_12649,N_11620);
nand U18088 (N_18088,N_10642,N_11887);
and U18089 (N_18089,N_13654,N_10487);
and U18090 (N_18090,N_10284,N_12882);
and U18091 (N_18091,N_13133,N_12824);
and U18092 (N_18092,N_14296,N_14841);
nor U18093 (N_18093,N_13373,N_14489);
or U18094 (N_18094,N_11584,N_10233);
nor U18095 (N_18095,N_13368,N_11851);
nor U18096 (N_18096,N_14246,N_12676);
nand U18097 (N_18097,N_12017,N_13758);
nand U18098 (N_18098,N_14299,N_12182);
or U18099 (N_18099,N_12558,N_11911);
or U18100 (N_18100,N_13641,N_12872);
nand U18101 (N_18101,N_14774,N_12003);
xor U18102 (N_18102,N_13809,N_14571);
or U18103 (N_18103,N_10071,N_12569);
nand U18104 (N_18104,N_11869,N_14928);
nand U18105 (N_18105,N_11146,N_10576);
and U18106 (N_18106,N_12237,N_12793);
or U18107 (N_18107,N_13542,N_10541);
nor U18108 (N_18108,N_12357,N_10628);
nand U18109 (N_18109,N_12884,N_11253);
xor U18110 (N_18110,N_10076,N_12601);
nor U18111 (N_18111,N_13725,N_13319);
nand U18112 (N_18112,N_11204,N_12229);
and U18113 (N_18113,N_13388,N_10490);
and U18114 (N_18114,N_13468,N_12414);
and U18115 (N_18115,N_10457,N_14639);
nor U18116 (N_18116,N_13906,N_11259);
and U18117 (N_18117,N_10053,N_14281);
nor U18118 (N_18118,N_11202,N_13028);
nor U18119 (N_18119,N_11516,N_11229);
nand U18120 (N_18120,N_14733,N_14921);
and U18121 (N_18121,N_11504,N_14218);
nor U18122 (N_18122,N_12613,N_10669);
nor U18123 (N_18123,N_12538,N_13639);
nor U18124 (N_18124,N_12703,N_12753);
nand U18125 (N_18125,N_12945,N_13855);
nor U18126 (N_18126,N_11183,N_12587);
or U18127 (N_18127,N_13408,N_13445);
nand U18128 (N_18128,N_12260,N_11533);
nand U18129 (N_18129,N_13048,N_13747);
or U18130 (N_18130,N_11200,N_14645);
or U18131 (N_18131,N_12818,N_12171);
xnor U18132 (N_18132,N_14132,N_13079);
and U18133 (N_18133,N_13305,N_14848);
and U18134 (N_18134,N_11055,N_14947);
and U18135 (N_18135,N_11994,N_12083);
nor U18136 (N_18136,N_10960,N_11237);
and U18137 (N_18137,N_10079,N_10491);
xnor U18138 (N_18138,N_13154,N_11601);
xor U18139 (N_18139,N_11261,N_10636);
nand U18140 (N_18140,N_12656,N_14118);
and U18141 (N_18141,N_12566,N_12575);
and U18142 (N_18142,N_13891,N_12646);
nand U18143 (N_18143,N_12137,N_10860);
nor U18144 (N_18144,N_13969,N_14665);
nand U18145 (N_18145,N_14610,N_10893);
or U18146 (N_18146,N_10992,N_12851);
or U18147 (N_18147,N_13610,N_11279);
or U18148 (N_18148,N_13337,N_14206);
or U18149 (N_18149,N_12594,N_10888);
nor U18150 (N_18150,N_13444,N_14206);
nand U18151 (N_18151,N_12189,N_12054);
nor U18152 (N_18152,N_13195,N_12744);
and U18153 (N_18153,N_14152,N_10806);
and U18154 (N_18154,N_11962,N_13008);
or U18155 (N_18155,N_11622,N_14492);
nand U18156 (N_18156,N_10196,N_12415);
nand U18157 (N_18157,N_10946,N_13861);
nand U18158 (N_18158,N_13326,N_12998);
or U18159 (N_18159,N_14064,N_14495);
or U18160 (N_18160,N_12670,N_13350);
and U18161 (N_18161,N_14259,N_11966);
nand U18162 (N_18162,N_11853,N_10893);
or U18163 (N_18163,N_12463,N_13782);
nor U18164 (N_18164,N_12061,N_13993);
or U18165 (N_18165,N_14784,N_13344);
nor U18166 (N_18166,N_14584,N_14905);
and U18167 (N_18167,N_11444,N_12836);
xor U18168 (N_18168,N_11570,N_10518);
nor U18169 (N_18169,N_13586,N_10661);
xnor U18170 (N_18170,N_10168,N_10925);
or U18171 (N_18171,N_13647,N_11473);
and U18172 (N_18172,N_14226,N_13161);
nand U18173 (N_18173,N_10871,N_13410);
or U18174 (N_18174,N_14049,N_14376);
and U18175 (N_18175,N_12538,N_11408);
and U18176 (N_18176,N_14783,N_13325);
xor U18177 (N_18177,N_10081,N_11800);
or U18178 (N_18178,N_14170,N_13755);
xor U18179 (N_18179,N_11321,N_12590);
and U18180 (N_18180,N_14075,N_14234);
nor U18181 (N_18181,N_10319,N_14471);
xnor U18182 (N_18182,N_11564,N_13145);
or U18183 (N_18183,N_10110,N_12549);
nor U18184 (N_18184,N_13866,N_12604);
and U18185 (N_18185,N_14785,N_14551);
nand U18186 (N_18186,N_10094,N_14494);
or U18187 (N_18187,N_14312,N_10344);
xnor U18188 (N_18188,N_12565,N_10235);
nand U18189 (N_18189,N_14514,N_12692);
or U18190 (N_18190,N_14543,N_10938);
and U18191 (N_18191,N_12792,N_11567);
and U18192 (N_18192,N_13843,N_14417);
or U18193 (N_18193,N_14538,N_13725);
and U18194 (N_18194,N_13233,N_13396);
nor U18195 (N_18195,N_10598,N_10366);
or U18196 (N_18196,N_12708,N_13438);
or U18197 (N_18197,N_10178,N_10626);
nor U18198 (N_18198,N_11435,N_10626);
nor U18199 (N_18199,N_10462,N_10386);
nand U18200 (N_18200,N_11495,N_12710);
and U18201 (N_18201,N_13784,N_11939);
and U18202 (N_18202,N_14868,N_14931);
or U18203 (N_18203,N_10852,N_10020);
and U18204 (N_18204,N_10854,N_14083);
nand U18205 (N_18205,N_13958,N_12129);
and U18206 (N_18206,N_14280,N_14505);
and U18207 (N_18207,N_10269,N_12361);
nand U18208 (N_18208,N_13725,N_14435);
nand U18209 (N_18209,N_10255,N_13612);
or U18210 (N_18210,N_10923,N_10230);
nor U18211 (N_18211,N_14948,N_14460);
and U18212 (N_18212,N_10621,N_10245);
and U18213 (N_18213,N_12428,N_11832);
and U18214 (N_18214,N_13183,N_10094);
or U18215 (N_18215,N_13724,N_12363);
xor U18216 (N_18216,N_12480,N_13738);
and U18217 (N_18217,N_10631,N_12809);
nor U18218 (N_18218,N_11016,N_13895);
xor U18219 (N_18219,N_14767,N_11699);
and U18220 (N_18220,N_10895,N_10595);
and U18221 (N_18221,N_11859,N_13650);
and U18222 (N_18222,N_11669,N_12428);
or U18223 (N_18223,N_10625,N_10416);
and U18224 (N_18224,N_12458,N_12508);
nand U18225 (N_18225,N_14453,N_14280);
nand U18226 (N_18226,N_13704,N_11785);
and U18227 (N_18227,N_12995,N_13877);
nand U18228 (N_18228,N_10821,N_12973);
nor U18229 (N_18229,N_14919,N_11473);
nand U18230 (N_18230,N_10868,N_12199);
and U18231 (N_18231,N_10790,N_11508);
or U18232 (N_18232,N_14231,N_10544);
nand U18233 (N_18233,N_10407,N_14352);
nor U18234 (N_18234,N_12952,N_14575);
or U18235 (N_18235,N_14548,N_14866);
and U18236 (N_18236,N_12552,N_14398);
nand U18237 (N_18237,N_10098,N_12646);
or U18238 (N_18238,N_10695,N_13139);
nor U18239 (N_18239,N_12017,N_12569);
and U18240 (N_18240,N_12315,N_11845);
xor U18241 (N_18241,N_14743,N_14754);
nand U18242 (N_18242,N_13913,N_10855);
and U18243 (N_18243,N_14739,N_13892);
nand U18244 (N_18244,N_14843,N_12902);
nor U18245 (N_18245,N_11874,N_10291);
nand U18246 (N_18246,N_10890,N_13855);
or U18247 (N_18247,N_11466,N_12955);
and U18248 (N_18248,N_11628,N_10492);
or U18249 (N_18249,N_13705,N_13899);
and U18250 (N_18250,N_12115,N_13485);
and U18251 (N_18251,N_11219,N_13842);
nor U18252 (N_18252,N_10836,N_11963);
nand U18253 (N_18253,N_11671,N_14057);
or U18254 (N_18254,N_11768,N_12563);
xnor U18255 (N_18255,N_12473,N_11586);
nand U18256 (N_18256,N_12850,N_10269);
nor U18257 (N_18257,N_11409,N_10987);
xor U18258 (N_18258,N_10368,N_11537);
nor U18259 (N_18259,N_14160,N_10158);
nor U18260 (N_18260,N_13985,N_14076);
and U18261 (N_18261,N_11550,N_13851);
nor U18262 (N_18262,N_14041,N_12443);
and U18263 (N_18263,N_12169,N_14916);
xnor U18264 (N_18264,N_11494,N_10103);
and U18265 (N_18265,N_14390,N_14372);
nor U18266 (N_18266,N_12572,N_11086);
nand U18267 (N_18267,N_13561,N_13938);
nand U18268 (N_18268,N_10311,N_10889);
or U18269 (N_18269,N_14588,N_13946);
and U18270 (N_18270,N_13729,N_13670);
or U18271 (N_18271,N_12586,N_13211);
and U18272 (N_18272,N_10372,N_10932);
nand U18273 (N_18273,N_11751,N_12118);
or U18274 (N_18274,N_11435,N_13371);
nor U18275 (N_18275,N_13345,N_10222);
nor U18276 (N_18276,N_11979,N_13990);
nor U18277 (N_18277,N_11726,N_11602);
xnor U18278 (N_18278,N_12381,N_10604);
or U18279 (N_18279,N_13624,N_14936);
and U18280 (N_18280,N_14413,N_14154);
and U18281 (N_18281,N_11459,N_14692);
nand U18282 (N_18282,N_11528,N_13174);
and U18283 (N_18283,N_13640,N_10795);
nor U18284 (N_18284,N_11389,N_14121);
and U18285 (N_18285,N_13835,N_13811);
or U18286 (N_18286,N_10044,N_10633);
nand U18287 (N_18287,N_12972,N_14860);
or U18288 (N_18288,N_13804,N_12076);
or U18289 (N_18289,N_12601,N_12362);
or U18290 (N_18290,N_10316,N_13998);
nor U18291 (N_18291,N_11728,N_12894);
xor U18292 (N_18292,N_12494,N_13042);
or U18293 (N_18293,N_12312,N_10618);
or U18294 (N_18294,N_14469,N_10978);
nor U18295 (N_18295,N_13776,N_12508);
and U18296 (N_18296,N_13544,N_14053);
nand U18297 (N_18297,N_11761,N_10468);
and U18298 (N_18298,N_14814,N_10937);
nand U18299 (N_18299,N_11232,N_13005);
and U18300 (N_18300,N_10277,N_10214);
nor U18301 (N_18301,N_13628,N_14098);
nand U18302 (N_18302,N_11832,N_11396);
nand U18303 (N_18303,N_11841,N_11205);
and U18304 (N_18304,N_10410,N_13597);
and U18305 (N_18305,N_14957,N_14572);
nor U18306 (N_18306,N_11147,N_10480);
nand U18307 (N_18307,N_12156,N_12793);
nor U18308 (N_18308,N_11683,N_10733);
xor U18309 (N_18309,N_10771,N_12728);
nand U18310 (N_18310,N_12980,N_10915);
xor U18311 (N_18311,N_13729,N_10685);
xnor U18312 (N_18312,N_12753,N_10808);
xor U18313 (N_18313,N_10840,N_12397);
or U18314 (N_18314,N_14193,N_10312);
or U18315 (N_18315,N_14167,N_14224);
xor U18316 (N_18316,N_11666,N_10875);
xnor U18317 (N_18317,N_11021,N_10305);
nor U18318 (N_18318,N_14882,N_12060);
and U18319 (N_18319,N_11760,N_10093);
nand U18320 (N_18320,N_14788,N_11848);
nor U18321 (N_18321,N_10367,N_10293);
nor U18322 (N_18322,N_13457,N_11608);
and U18323 (N_18323,N_13963,N_10884);
nand U18324 (N_18324,N_12128,N_14535);
xnor U18325 (N_18325,N_13843,N_12213);
nor U18326 (N_18326,N_12039,N_14156);
xor U18327 (N_18327,N_10118,N_11853);
or U18328 (N_18328,N_11011,N_14117);
or U18329 (N_18329,N_10930,N_12444);
nand U18330 (N_18330,N_14266,N_12293);
nor U18331 (N_18331,N_11180,N_14189);
or U18332 (N_18332,N_13051,N_14194);
and U18333 (N_18333,N_13785,N_10680);
nand U18334 (N_18334,N_10432,N_10210);
or U18335 (N_18335,N_11626,N_10661);
nand U18336 (N_18336,N_13179,N_13961);
nor U18337 (N_18337,N_10194,N_12873);
nor U18338 (N_18338,N_13935,N_13710);
or U18339 (N_18339,N_14724,N_14526);
xnor U18340 (N_18340,N_12136,N_11168);
nand U18341 (N_18341,N_12041,N_14732);
nor U18342 (N_18342,N_12134,N_10693);
or U18343 (N_18343,N_13216,N_10179);
xor U18344 (N_18344,N_10453,N_12975);
nor U18345 (N_18345,N_12752,N_13544);
or U18346 (N_18346,N_14240,N_10962);
nor U18347 (N_18347,N_14921,N_12812);
nand U18348 (N_18348,N_11970,N_11248);
and U18349 (N_18349,N_11832,N_10304);
nor U18350 (N_18350,N_14344,N_14659);
xor U18351 (N_18351,N_11918,N_10482);
nand U18352 (N_18352,N_11251,N_12524);
and U18353 (N_18353,N_12593,N_13375);
nor U18354 (N_18354,N_14378,N_12241);
nand U18355 (N_18355,N_10396,N_12843);
nand U18356 (N_18356,N_13873,N_10431);
nor U18357 (N_18357,N_14736,N_12609);
and U18358 (N_18358,N_14434,N_10703);
xnor U18359 (N_18359,N_14448,N_12266);
or U18360 (N_18360,N_11800,N_14910);
xor U18361 (N_18361,N_12130,N_11301);
xnor U18362 (N_18362,N_10845,N_13920);
nand U18363 (N_18363,N_14596,N_14747);
or U18364 (N_18364,N_13272,N_12065);
and U18365 (N_18365,N_14944,N_10835);
xor U18366 (N_18366,N_11910,N_12703);
and U18367 (N_18367,N_13658,N_11645);
nor U18368 (N_18368,N_13327,N_11426);
and U18369 (N_18369,N_11101,N_13822);
nor U18370 (N_18370,N_10636,N_12932);
or U18371 (N_18371,N_13261,N_11649);
or U18372 (N_18372,N_14987,N_11723);
or U18373 (N_18373,N_13941,N_12520);
or U18374 (N_18374,N_12482,N_10089);
xnor U18375 (N_18375,N_10100,N_11549);
nor U18376 (N_18376,N_12340,N_14343);
or U18377 (N_18377,N_13014,N_11337);
nor U18378 (N_18378,N_12177,N_12004);
nor U18379 (N_18379,N_12131,N_10421);
nand U18380 (N_18380,N_11660,N_12240);
or U18381 (N_18381,N_14217,N_12838);
and U18382 (N_18382,N_14072,N_14326);
nor U18383 (N_18383,N_10013,N_12561);
nor U18384 (N_18384,N_11605,N_12466);
and U18385 (N_18385,N_13537,N_10788);
xnor U18386 (N_18386,N_14740,N_12947);
nor U18387 (N_18387,N_11514,N_10255);
and U18388 (N_18388,N_13486,N_10258);
nand U18389 (N_18389,N_14507,N_10266);
nor U18390 (N_18390,N_11394,N_12557);
xor U18391 (N_18391,N_14459,N_10609);
nand U18392 (N_18392,N_12168,N_14856);
nand U18393 (N_18393,N_11468,N_12013);
nor U18394 (N_18394,N_12384,N_12308);
nand U18395 (N_18395,N_14206,N_11188);
and U18396 (N_18396,N_14405,N_10800);
and U18397 (N_18397,N_13197,N_11166);
nor U18398 (N_18398,N_10714,N_12943);
or U18399 (N_18399,N_14538,N_14210);
and U18400 (N_18400,N_11060,N_14788);
xor U18401 (N_18401,N_11336,N_10558);
and U18402 (N_18402,N_10270,N_14541);
xnor U18403 (N_18403,N_11488,N_14403);
or U18404 (N_18404,N_12993,N_12458);
nor U18405 (N_18405,N_14667,N_11394);
nand U18406 (N_18406,N_14000,N_14174);
nor U18407 (N_18407,N_13328,N_14115);
nand U18408 (N_18408,N_10313,N_13097);
nor U18409 (N_18409,N_11450,N_12662);
or U18410 (N_18410,N_12500,N_12339);
nor U18411 (N_18411,N_13382,N_10332);
and U18412 (N_18412,N_13400,N_14985);
nand U18413 (N_18413,N_12979,N_12674);
nand U18414 (N_18414,N_12265,N_12776);
nor U18415 (N_18415,N_13050,N_12640);
and U18416 (N_18416,N_14525,N_11423);
nor U18417 (N_18417,N_12654,N_14005);
nor U18418 (N_18418,N_13218,N_14885);
and U18419 (N_18419,N_11014,N_12666);
nor U18420 (N_18420,N_10145,N_12958);
xor U18421 (N_18421,N_14000,N_11637);
nor U18422 (N_18422,N_11077,N_13255);
or U18423 (N_18423,N_11632,N_14876);
or U18424 (N_18424,N_13486,N_13863);
or U18425 (N_18425,N_14508,N_13559);
nor U18426 (N_18426,N_10604,N_13825);
nand U18427 (N_18427,N_11005,N_14231);
or U18428 (N_18428,N_10110,N_10450);
nor U18429 (N_18429,N_10159,N_12593);
nand U18430 (N_18430,N_14426,N_14910);
and U18431 (N_18431,N_12111,N_10923);
and U18432 (N_18432,N_13898,N_10538);
or U18433 (N_18433,N_11254,N_11379);
nor U18434 (N_18434,N_14937,N_12618);
nand U18435 (N_18435,N_12913,N_12078);
and U18436 (N_18436,N_12359,N_11310);
and U18437 (N_18437,N_14073,N_14245);
or U18438 (N_18438,N_14278,N_12028);
nor U18439 (N_18439,N_14162,N_14349);
or U18440 (N_18440,N_10971,N_14503);
or U18441 (N_18441,N_13137,N_13072);
nand U18442 (N_18442,N_13389,N_10808);
or U18443 (N_18443,N_14970,N_14206);
nand U18444 (N_18444,N_12834,N_14927);
or U18445 (N_18445,N_12422,N_13060);
and U18446 (N_18446,N_12552,N_12586);
or U18447 (N_18447,N_13882,N_13580);
or U18448 (N_18448,N_11220,N_13381);
nor U18449 (N_18449,N_13723,N_12708);
and U18450 (N_18450,N_13132,N_11062);
nor U18451 (N_18451,N_12401,N_14456);
xor U18452 (N_18452,N_11052,N_12428);
nand U18453 (N_18453,N_11659,N_14837);
and U18454 (N_18454,N_11463,N_13051);
xor U18455 (N_18455,N_11869,N_13995);
and U18456 (N_18456,N_13824,N_13035);
and U18457 (N_18457,N_11800,N_14955);
nor U18458 (N_18458,N_11456,N_10381);
or U18459 (N_18459,N_13979,N_14969);
and U18460 (N_18460,N_10693,N_13862);
xnor U18461 (N_18461,N_13532,N_13897);
and U18462 (N_18462,N_10429,N_10380);
and U18463 (N_18463,N_12856,N_10021);
nand U18464 (N_18464,N_13953,N_11550);
or U18465 (N_18465,N_10977,N_12561);
nor U18466 (N_18466,N_12095,N_12622);
or U18467 (N_18467,N_10721,N_11456);
and U18468 (N_18468,N_11195,N_10978);
and U18469 (N_18469,N_11054,N_10047);
or U18470 (N_18470,N_11457,N_10973);
and U18471 (N_18471,N_13477,N_14756);
nand U18472 (N_18472,N_13476,N_11666);
and U18473 (N_18473,N_10498,N_13743);
nand U18474 (N_18474,N_14010,N_12228);
xnor U18475 (N_18475,N_13121,N_13779);
nor U18476 (N_18476,N_13259,N_14885);
and U18477 (N_18477,N_14385,N_10719);
or U18478 (N_18478,N_10452,N_13461);
nor U18479 (N_18479,N_10416,N_10038);
or U18480 (N_18480,N_12479,N_14988);
or U18481 (N_18481,N_13346,N_13584);
nand U18482 (N_18482,N_11997,N_14423);
or U18483 (N_18483,N_10441,N_13185);
and U18484 (N_18484,N_14403,N_14473);
nand U18485 (N_18485,N_13598,N_12954);
xnor U18486 (N_18486,N_12609,N_12233);
or U18487 (N_18487,N_10886,N_11790);
nor U18488 (N_18488,N_10385,N_13044);
nor U18489 (N_18489,N_12103,N_14831);
and U18490 (N_18490,N_13905,N_11559);
or U18491 (N_18491,N_12853,N_11166);
and U18492 (N_18492,N_11151,N_12565);
and U18493 (N_18493,N_11938,N_12885);
xor U18494 (N_18494,N_11090,N_12149);
nand U18495 (N_18495,N_13334,N_13516);
and U18496 (N_18496,N_14506,N_11023);
nand U18497 (N_18497,N_11996,N_13924);
or U18498 (N_18498,N_12138,N_11285);
and U18499 (N_18499,N_10804,N_11799);
and U18500 (N_18500,N_10165,N_14552);
nand U18501 (N_18501,N_13591,N_14130);
and U18502 (N_18502,N_14104,N_12999);
or U18503 (N_18503,N_11480,N_11665);
nand U18504 (N_18504,N_10487,N_13400);
nand U18505 (N_18505,N_11221,N_13591);
or U18506 (N_18506,N_12856,N_13135);
xnor U18507 (N_18507,N_14258,N_13383);
or U18508 (N_18508,N_13598,N_11020);
xnor U18509 (N_18509,N_14353,N_14508);
nand U18510 (N_18510,N_13635,N_14016);
or U18511 (N_18511,N_10061,N_10714);
or U18512 (N_18512,N_11507,N_14234);
and U18513 (N_18513,N_14045,N_12080);
or U18514 (N_18514,N_12895,N_13190);
nand U18515 (N_18515,N_14499,N_10739);
xnor U18516 (N_18516,N_13967,N_13063);
nand U18517 (N_18517,N_11733,N_14801);
or U18518 (N_18518,N_11985,N_11087);
nand U18519 (N_18519,N_11768,N_10418);
or U18520 (N_18520,N_11589,N_13064);
and U18521 (N_18521,N_11333,N_12573);
or U18522 (N_18522,N_12147,N_11248);
or U18523 (N_18523,N_12622,N_10688);
xor U18524 (N_18524,N_13817,N_14564);
or U18525 (N_18525,N_14742,N_12671);
and U18526 (N_18526,N_10356,N_13355);
nor U18527 (N_18527,N_13015,N_10480);
xnor U18528 (N_18528,N_13673,N_12701);
and U18529 (N_18529,N_13523,N_12159);
and U18530 (N_18530,N_11182,N_14355);
or U18531 (N_18531,N_12765,N_12819);
or U18532 (N_18532,N_14312,N_13809);
or U18533 (N_18533,N_10091,N_12548);
or U18534 (N_18534,N_11946,N_10616);
or U18535 (N_18535,N_13861,N_12897);
nand U18536 (N_18536,N_13134,N_12789);
or U18537 (N_18537,N_13558,N_11278);
nand U18538 (N_18538,N_14208,N_12196);
xnor U18539 (N_18539,N_14383,N_13666);
nand U18540 (N_18540,N_14546,N_13342);
nor U18541 (N_18541,N_10911,N_14181);
nand U18542 (N_18542,N_11796,N_14163);
nor U18543 (N_18543,N_10839,N_10153);
nor U18544 (N_18544,N_11369,N_11608);
or U18545 (N_18545,N_10372,N_12369);
or U18546 (N_18546,N_14939,N_13977);
or U18547 (N_18547,N_14116,N_13789);
nor U18548 (N_18548,N_13297,N_14443);
and U18549 (N_18549,N_14627,N_12981);
nand U18550 (N_18550,N_14110,N_12349);
nor U18551 (N_18551,N_13704,N_11726);
or U18552 (N_18552,N_10771,N_14412);
and U18553 (N_18553,N_11639,N_11177);
nor U18554 (N_18554,N_11368,N_13003);
nand U18555 (N_18555,N_10719,N_14950);
nor U18556 (N_18556,N_13897,N_13889);
and U18557 (N_18557,N_12765,N_13964);
or U18558 (N_18558,N_12362,N_13923);
nand U18559 (N_18559,N_11025,N_11859);
nand U18560 (N_18560,N_12460,N_13763);
and U18561 (N_18561,N_13963,N_12173);
nand U18562 (N_18562,N_14536,N_11682);
nor U18563 (N_18563,N_12247,N_14754);
and U18564 (N_18564,N_13851,N_12829);
nand U18565 (N_18565,N_10848,N_14660);
and U18566 (N_18566,N_10607,N_10174);
nor U18567 (N_18567,N_11775,N_13879);
or U18568 (N_18568,N_11365,N_10320);
nand U18569 (N_18569,N_14085,N_13273);
nor U18570 (N_18570,N_14574,N_12713);
nand U18571 (N_18571,N_10216,N_10347);
nand U18572 (N_18572,N_13085,N_14542);
and U18573 (N_18573,N_11159,N_12376);
xnor U18574 (N_18574,N_13776,N_11604);
nor U18575 (N_18575,N_14928,N_10348);
or U18576 (N_18576,N_14870,N_10480);
and U18577 (N_18577,N_11884,N_12351);
or U18578 (N_18578,N_14714,N_13988);
xor U18579 (N_18579,N_12224,N_13999);
nor U18580 (N_18580,N_13588,N_11956);
nand U18581 (N_18581,N_12699,N_14571);
or U18582 (N_18582,N_12804,N_13601);
or U18583 (N_18583,N_11773,N_12308);
nand U18584 (N_18584,N_13210,N_13339);
xor U18585 (N_18585,N_11203,N_10726);
xnor U18586 (N_18586,N_13364,N_13959);
and U18587 (N_18587,N_11705,N_12085);
and U18588 (N_18588,N_14208,N_13043);
or U18589 (N_18589,N_12593,N_12129);
or U18590 (N_18590,N_10739,N_12077);
and U18591 (N_18591,N_12607,N_12291);
nand U18592 (N_18592,N_14614,N_10656);
nand U18593 (N_18593,N_10517,N_13120);
nor U18594 (N_18594,N_12575,N_11971);
nand U18595 (N_18595,N_10555,N_10809);
and U18596 (N_18596,N_11877,N_13676);
nand U18597 (N_18597,N_11157,N_14784);
and U18598 (N_18598,N_10922,N_14070);
nand U18599 (N_18599,N_14125,N_14181);
or U18600 (N_18600,N_13700,N_14374);
and U18601 (N_18601,N_12510,N_14567);
and U18602 (N_18602,N_12248,N_11973);
and U18603 (N_18603,N_14511,N_13535);
or U18604 (N_18604,N_10477,N_13217);
and U18605 (N_18605,N_10701,N_14733);
and U18606 (N_18606,N_11313,N_12746);
nand U18607 (N_18607,N_14240,N_10535);
nand U18608 (N_18608,N_11881,N_12639);
nor U18609 (N_18609,N_10172,N_10770);
nor U18610 (N_18610,N_10295,N_10433);
and U18611 (N_18611,N_14200,N_11824);
and U18612 (N_18612,N_13354,N_11283);
nor U18613 (N_18613,N_12349,N_10789);
nand U18614 (N_18614,N_14594,N_12898);
or U18615 (N_18615,N_14330,N_13562);
nand U18616 (N_18616,N_10195,N_13470);
xor U18617 (N_18617,N_13469,N_13172);
or U18618 (N_18618,N_13097,N_12401);
and U18619 (N_18619,N_10873,N_12081);
nand U18620 (N_18620,N_14553,N_14436);
nor U18621 (N_18621,N_13201,N_12523);
and U18622 (N_18622,N_12505,N_14482);
or U18623 (N_18623,N_14485,N_10781);
nand U18624 (N_18624,N_10475,N_12441);
or U18625 (N_18625,N_10710,N_11703);
or U18626 (N_18626,N_11599,N_11968);
nand U18627 (N_18627,N_14710,N_13249);
nand U18628 (N_18628,N_13381,N_10397);
xnor U18629 (N_18629,N_14721,N_11864);
nand U18630 (N_18630,N_10350,N_14498);
or U18631 (N_18631,N_12361,N_11177);
or U18632 (N_18632,N_10900,N_10254);
and U18633 (N_18633,N_14129,N_11337);
nand U18634 (N_18634,N_11657,N_11803);
nor U18635 (N_18635,N_14727,N_13466);
or U18636 (N_18636,N_10943,N_12938);
nor U18637 (N_18637,N_11467,N_13394);
xor U18638 (N_18638,N_12892,N_12108);
nand U18639 (N_18639,N_13255,N_13918);
or U18640 (N_18640,N_13317,N_11594);
or U18641 (N_18641,N_10842,N_13792);
nor U18642 (N_18642,N_10707,N_11196);
nand U18643 (N_18643,N_11298,N_10914);
nor U18644 (N_18644,N_10641,N_13775);
and U18645 (N_18645,N_13773,N_11252);
nand U18646 (N_18646,N_10870,N_14362);
and U18647 (N_18647,N_10184,N_14043);
or U18648 (N_18648,N_12133,N_13544);
nor U18649 (N_18649,N_11223,N_11502);
nand U18650 (N_18650,N_13365,N_11476);
nand U18651 (N_18651,N_13261,N_11185);
nand U18652 (N_18652,N_13570,N_10645);
nor U18653 (N_18653,N_12245,N_11985);
or U18654 (N_18654,N_10613,N_13666);
or U18655 (N_18655,N_13896,N_10622);
and U18656 (N_18656,N_14346,N_10739);
nor U18657 (N_18657,N_14784,N_11131);
nor U18658 (N_18658,N_14222,N_11869);
nor U18659 (N_18659,N_12320,N_11971);
or U18660 (N_18660,N_14025,N_13559);
nor U18661 (N_18661,N_13731,N_10270);
or U18662 (N_18662,N_12049,N_10214);
or U18663 (N_18663,N_11644,N_13600);
nor U18664 (N_18664,N_10986,N_14780);
and U18665 (N_18665,N_10341,N_13797);
and U18666 (N_18666,N_14060,N_12163);
nor U18667 (N_18667,N_10493,N_10334);
nor U18668 (N_18668,N_11378,N_12564);
and U18669 (N_18669,N_10238,N_10725);
nand U18670 (N_18670,N_10423,N_13282);
nand U18671 (N_18671,N_14365,N_10008);
and U18672 (N_18672,N_10447,N_12049);
nand U18673 (N_18673,N_12271,N_12292);
or U18674 (N_18674,N_13551,N_12106);
nand U18675 (N_18675,N_14182,N_12978);
or U18676 (N_18676,N_11203,N_13969);
or U18677 (N_18677,N_12191,N_13769);
or U18678 (N_18678,N_12804,N_11593);
xnor U18679 (N_18679,N_12184,N_12407);
nand U18680 (N_18680,N_12283,N_13678);
nand U18681 (N_18681,N_13973,N_12902);
or U18682 (N_18682,N_11643,N_14499);
or U18683 (N_18683,N_13874,N_11913);
nand U18684 (N_18684,N_12132,N_13436);
or U18685 (N_18685,N_13484,N_13420);
xor U18686 (N_18686,N_12259,N_14531);
xor U18687 (N_18687,N_10634,N_14610);
nor U18688 (N_18688,N_10204,N_14984);
or U18689 (N_18689,N_12645,N_14623);
and U18690 (N_18690,N_13488,N_12130);
nand U18691 (N_18691,N_11367,N_13004);
nor U18692 (N_18692,N_12437,N_14753);
nor U18693 (N_18693,N_14238,N_14154);
xnor U18694 (N_18694,N_13501,N_13846);
nor U18695 (N_18695,N_13400,N_10132);
nand U18696 (N_18696,N_12241,N_11732);
or U18697 (N_18697,N_14209,N_11750);
and U18698 (N_18698,N_14240,N_14121);
nor U18699 (N_18699,N_11186,N_11129);
xor U18700 (N_18700,N_11014,N_12957);
nor U18701 (N_18701,N_13818,N_12684);
nor U18702 (N_18702,N_12701,N_13042);
nor U18703 (N_18703,N_13992,N_11525);
or U18704 (N_18704,N_13254,N_13211);
nand U18705 (N_18705,N_13058,N_10238);
and U18706 (N_18706,N_12441,N_13309);
and U18707 (N_18707,N_10558,N_10079);
and U18708 (N_18708,N_10421,N_14295);
nand U18709 (N_18709,N_10446,N_12293);
nor U18710 (N_18710,N_10980,N_12544);
xor U18711 (N_18711,N_14604,N_11112);
nand U18712 (N_18712,N_11718,N_10488);
and U18713 (N_18713,N_11391,N_14984);
nand U18714 (N_18714,N_14627,N_10969);
nand U18715 (N_18715,N_11854,N_14549);
nor U18716 (N_18716,N_11027,N_14272);
nor U18717 (N_18717,N_14158,N_14692);
or U18718 (N_18718,N_13388,N_10682);
nor U18719 (N_18719,N_14203,N_14311);
and U18720 (N_18720,N_11769,N_12990);
xnor U18721 (N_18721,N_13695,N_13908);
xor U18722 (N_18722,N_12658,N_10070);
nand U18723 (N_18723,N_11843,N_12547);
nand U18724 (N_18724,N_12466,N_11725);
nand U18725 (N_18725,N_13504,N_10298);
or U18726 (N_18726,N_14831,N_14362);
and U18727 (N_18727,N_12325,N_14511);
or U18728 (N_18728,N_11028,N_10612);
nor U18729 (N_18729,N_14106,N_10819);
xor U18730 (N_18730,N_12698,N_10868);
and U18731 (N_18731,N_12041,N_11817);
or U18732 (N_18732,N_14152,N_12438);
and U18733 (N_18733,N_14545,N_10441);
nor U18734 (N_18734,N_10896,N_10263);
nand U18735 (N_18735,N_11406,N_14750);
or U18736 (N_18736,N_11857,N_14767);
or U18737 (N_18737,N_12908,N_12505);
nand U18738 (N_18738,N_12656,N_10063);
nor U18739 (N_18739,N_12349,N_11983);
nor U18740 (N_18740,N_13150,N_10564);
or U18741 (N_18741,N_13716,N_12604);
nand U18742 (N_18742,N_12714,N_12307);
and U18743 (N_18743,N_10101,N_12398);
or U18744 (N_18744,N_14596,N_10443);
nand U18745 (N_18745,N_12772,N_11564);
and U18746 (N_18746,N_13143,N_12131);
and U18747 (N_18747,N_14399,N_11508);
nand U18748 (N_18748,N_12414,N_14641);
nor U18749 (N_18749,N_12744,N_14487);
or U18750 (N_18750,N_11211,N_13996);
or U18751 (N_18751,N_12027,N_10492);
or U18752 (N_18752,N_14029,N_12519);
nand U18753 (N_18753,N_14250,N_14670);
xnor U18754 (N_18754,N_14677,N_12334);
xnor U18755 (N_18755,N_11154,N_14152);
nor U18756 (N_18756,N_14010,N_11379);
nand U18757 (N_18757,N_12878,N_13984);
or U18758 (N_18758,N_13184,N_12593);
nor U18759 (N_18759,N_13932,N_10058);
and U18760 (N_18760,N_14559,N_13136);
and U18761 (N_18761,N_11286,N_13933);
or U18762 (N_18762,N_14705,N_12285);
nand U18763 (N_18763,N_12909,N_10810);
or U18764 (N_18764,N_13900,N_14025);
nor U18765 (N_18765,N_14016,N_14259);
nor U18766 (N_18766,N_10251,N_14796);
nor U18767 (N_18767,N_12869,N_13074);
and U18768 (N_18768,N_13499,N_13768);
nand U18769 (N_18769,N_11311,N_13922);
nor U18770 (N_18770,N_13390,N_13578);
and U18771 (N_18771,N_12966,N_14003);
or U18772 (N_18772,N_11614,N_10350);
nor U18773 (N_18773,N_14730,N_14705);
or U18774 (N_18774,N_12301,N_13385);
nor U18775 (N_18775,N_12409,N_14711);
and U18776 (N_18776,N_14232,N_14839);
xnor U18777 (N_18777,N_13639,N_14438);
nand U18778 (N_18778,N_10355,N_12872);
nand U18779 (N_18779,N_12066,N_12954);
nor U18780 (N_18780,N_13976,N_14903);
nor U18781 (N_18781,N_12249,N_14904);
or U18782 (N_18782,N_13945,N_13983);
nor U18783 (N_18783,N_14134,N_11860);
xnor U18784 (N_18784,N_12633,N_12243);
nor U18785 (N_18785,N_13465,N_13670);
or U18786 (N_18786,N_14301,N_11747);
nor U18787 (N_18787,N_13758,N_14045);
nand U18788 (N_18788,N_12612,N_12889);
xnor U18789 (N_18789,N_13898,N_10913);
and U18790 (N_18790,N_13258,N_10033);
nand U18791 (N_18791,N_12081,N_11219);
nand U18792 (N_18792,N_14143,N_11925);
and U18793 (N_18793,N_13053,N_12373);
xnor U18794 (N_18794,N_13340,N_10073);
or U18795 (N_18795,N_11710,N_12222);
xnor U18796 (N_18796,N_14185,N_11076);
or U18797 (N_18797,N_11400,N_11411);
or U18798 (N_18798,N_14820,N_14944);
or U18799 (N_18799,N_10724,N_11593);
or U18800 (N_18800,N_13601,N_14805);
and U18801 (N_18801,N_13826,N_14845);
or U18802 (N_18802,N_11285,N_10407);
nand U18803 (N_18803,N_14159,N_13734);
nand U18804 (N_18804,N_13698,N_10904);
nand U18805 (N_18805,N_11963,N_10000);
nor U18806 (N_18806,N_14287,N_12096);
nor U18807 (N_18807,N_12372,N_14323);
nor U18808 (N_18808,N_10720,N_14308);
or U18809 (N_18809,N_13122,N_14455);
or U18810 (N_18810,N_10049,N_12849);
and U18811 (N_18811,N_10334,N_10415);
nand U18812 (N_18812,N_10919,N_14235);
nor U18813 (N_18813,N_12782,N_14909);
or U18814 (N_18814,N_13010,N_10370);
and U18815 (N_18815,N_11009,N_13457);
and U18816 (N_18816,N_14869,N_13555);
and U18817 (N_18817,N_13890,N_11089);
nand U18818 (N_18818,N_13909,N_10890);
nor U18819 (N_18819,N_10477,N_11153);
xnor U18820 (N_18820,N_14036,N_11272);
and U18821 (N_18821,N_10224,N_13590);
and U18822 (N_18822,N_12888,N_10936);
xnor U18823 (N_18823,N_14249,N_12114);
or U18824 (N_18824,N_12477,N_12533);
nand U18825 (N_18825,N_14129,N_12683);
or U18826 (N_18826,N_13577,N_12313);
or U18827 (N_18827,N_14985,N_10610);
or U18828 (N_18828,N_12597,N_13974);
and U18829 (N_18829,N_11362,N_12592);
or U18830 (N_18830,N_11273,N_12910);
nand U18831 (N_18831,N_13300,N_11530);
or U18832 (N_18832,N_11804,N_10421);
nand U18833 (N_18833,N_10427,N_14113);
nand U18834 (N_18834,N_14694,N_10431);
nor U18835 (N_18835,N_14296,N_11197);
or U18836 (N_18836,N_12152,N_11969);
or U18837 (N_18837,N_12657,N_14086);
and U18838 (N_18838,N_13449,N_11384);
nor U18839 (N_18839,N_13773,N_11219);
nand U18840 (N_18840,N_14905,N_13421);
and U18841 (N_18841,N_12689,N_11423);
or U18842 (N_18842,N_13868,N_10812);
or U18843 (N_18843,N_14677,N_12488);
nand U18844 (N_18844,N_12627,N_10116);
or U18845 (N_18845,N_14844,N_12844);
nand U18846 (N_18846,N_10609,N_13402);
nand U18847 (N_18847,N_13154,N_11690);
xnor U18848 (N_18848,N_14645,N_12884);
nor U18849 (N_18849,N_10906,N_12571);
xor U18850 (N_18850,N_12888,N_10931);
and U18851 (N_18851,N_13896,N_12753);
nor U18852 (N_18852,N_13427,N_10557);
nand U18853 (N_18853,N_11190,N_14264);
and U18854 (N_18854,N_13020,N_14040);
nor U18855 (N_18855,N_12810,N_12665);
nor U18856 (N_18856,N_10361,N_10286);
nor U18857 (N_18857,N_11303,N_11862);
nor U18858 (N_18858,N_12402,N_13198);
or U18859 (N_18859,N_14599,N_13961);
and U18860 (N_18860,N_14030,N_12734);
or U18861 (N_18861,N_11866,N_14795);
and U18862 (N_18862,N_13932,N_11355);
nor U18863 (N_18863,N_11138,N_10769);
nor U18864 (N_18864,N_14522,N_11409);
or U18865 (N_18865,N_12415,N_11845);
nor U18866 (N_18866,N_11985,N_14799);
nand U18867 (N_18867,N_14822,N_13293);
and U18868 (N_18868,N_10440,N_11929);
xor U18869 (N_18869,N_14525,N_13294);
and U18870 (N_18870,N_12531,N_12358);
nor U18871 (N_18871,N_10542,N_11962);
and U18872 (N_18872,N_13001,N_13614);
nor U18873 (N_18873,N_14502,N_13154);
and U18874 (N_18874,N_13718,N_13239);
xnor U18875 (N_18875,N_13715,N_10678);
or U18876 (N_18876,N_13274,N_12775);
xnor U18877 (N_18877,N_14696,N_11025);
nor U18878 (N_18878,N_14095,N_13222);
nand U18879 (N_18879,N_10733,N_11761);
and U18880 (N_18880,N_11442,N_12273);
or U18881 (N_18881,N_14751,N_14255);
nor U18882 (N_18882,N_10981,N_14887);
nor U18883 (N_18883,N_11098,N_12494);
nor U18884 (N_18884,N_11818,N_11960);
xor U18885 (N_18885,N_11376,N_10630);
nor U18886 (N_18886,N_11864,N_12346);
or U18887 (N_18887,N_12665,N_14562);
nand U18888 (N_18888,N_14383,N_14055);
xor U18889 (N_18889,N_13417,N_10319);
nor U18890 (N_18890,N_14929,N_12565);
xnor U18891 (N_18891,N_11470,N_11574);
and U18892 (N_18892,N_11429,N_10580);
or U18893 (N_18893,N_14715,N_13498);
nand U18894 (N_18894,N_10966,N_12419);
nor U18895 (N_18895,N_11185,N_12552);
and U18896 (N_18896,N_13307,N_13781);
nand U18897 (N_18897,N_11912,N_10986);
and U18898 (N_18898,N_14592,N_14537);
nor U18899 (N_18899,N_13692,N_14394);
nand U18900 (N_18900,N_14136,N_13136);
xnor U18901 (N_18901,N_12991,N_13775);
and U18902 (N_18902,N_13314,N_14837);
or U18903 (N_18903,N_14810,N_13586);
and U18904 (N_18904,N_11796,N_10430);
and U18905 (N_18905,N_11032,N_11655);
and U18906 (N_18906,N_12818,N_11999);
and U18907 (N_18907,N_10015,N_10588);
nand U18908 (N_18908,N_11620,N_12131);
and U18909 (N_18909,N_11276,N_13648);
and U18910 (N_18910,N_13351,N_10166);
nor U18911 (N_18911,N_12073,N_11109);
xnor U18912 (N_18912,N_13955,N_10722);
nor U18913 (N_18913,N_13683,N_14344);
nor U18914 (N_18914,N_13646,N_13491);
or U18915 (N_18915,N_13282,N_10825);
nand U18916 (N_18916,N_14667,N_12758);
nor U18917 (N_18917,N_11724,N_14587);
nor U18918 (N_18918,N_12663,N_10676);
nand U18919 (N_18919,N_10932,N_12510);
or U18920 (N_18920,N_14601,N_14229);
or U18921 (N_18921,N_12915,N_10431);
nand U18922 (N_18922,N_14197,N_12086);
and U18923 (N_18923,N_13712,N_11133);
xnor U18924 (N_18924,N_10087,N_11872);
nor U18925 (N_18925,N_13446,N_12272);
nand U18926 (N_18926,N_12447,N_11237);
and U18927 (N_18927,N_13111,N_11057);
xor U18928 (N_18928,N_11742,N_14364);
and U18929 (N_18929,N_10402,N_11973);
or U18930 (N_18930,N_12198,N_13927);
nor U18931 (N_18931,N_11320,N_12130);
xor U18932 (N_18932,N_14135,N_11348);
nand U18933 (N_18933,N_11802,N_13167);
nor U18934 (N_18934,N_10116,N_13556);
nand U18935 (N_18935,N_14773,N_11633);
and U18936 (N_18936,N_11336,N_11128);
nor U18937 (N_18937,N_11456,N_14478);
xnor U18938 (N_18938,N_13998,N_13378);
nand U18939 (N_18939,N_11909,N_11093);
xnor U18940 (N_18940,N_12786,N_13932);
xnor U18941 (N_18941,N_13165,N_12048);
nor U18942 (N_18942,N_14558,N_10917);
nor U18943 (N_18943,N_14283,N_10437);
and U18944 (N_18944,N_11025,N_14937);
or U18945 (N_18945,N_12459,N_11046);
nand U18946 (N_18946,N_12636,N_13544);
or U18947 (N_18947,N_12298,N_10273);
or U18948 (N_18948,N_12695,N_14705);
and U18949 (N_18949,N_14436,N_12774);
and U18950 (N_18950,N_14155,N_11054);
nand U18951 (N_18951,N_13270,N_12943);
nand U18952 (N_18952,N_10917,N_11651);
nand U18953 (N_18953,N_11013,N_13625);
nand U18954 (N_18954,N_14959,N_11926);
and U18955 (N_18955,N_14083,N_10644);
and U18956 (N_18956,N_10020,N_10083);
and U18957 (N_18957,N_11586,N_14891);
and U18958 (N_18958,N_12592,N_14672);
or U18959 (N_18959,N_13427,N_14975);
nand U18960 (N_18960,N_11359,N_11681);
and U18961 (N_18961,N_13342,N_11915);
and U18962 (N_18962,N_13290,N_11397);
xnor U18963 (N_18963,N_14917,N_10196);
or U18964 (N_18964,N_11626,N_10880);
nor U18965 (N_18965,N_14410,N_10258);
nand U18966 (N_18966,N_12046,N_14852);
and U18967 (N_18967,N_12040,N_11120);
and U18968 (N_18968,N_13084,N_13014);
nand U18969 (N_18969,N_14997,N_10994);
xor U18970 (N_18970,N_11819,N_11181);
xor U18971 (N_18971,N_13056,N_11131);
nand U18972 (N_18972,N_12505,N_10024);
nand U18973 (N_18973,N_11791,N_11429);
and U18974 (N_18974,N_10794,N_14143);
or U18975 (N_18975,N_14582,N_14438);
and U18976 (N_18976,N_11817,N_11426);
xor U18977 (N_18977,N_13508,N_11362);
and U18978 (N_18978,N_11178,N_13795);
nand U18979 (N_18979,N_12567,N_13356);
nand U18980 (N_18980,N_13201,N_13444);
nand U18981 (N_18981,N_14163,N_12603);
or U18982 (N_18982,N_13246,N_10925);
or U18983 (N_18983,N_14744,N_11625);
and U18984 (N_18984,N_12226,N_12536);
or U18985 (N_18985,N_14126,N_11831);
nor U18986 (N_18986,N_11189,N_10890);
nor U18987 (N_18987,N_14594,N_12339);
nor U18988 (N_18988,N_11258,N_12640);
nand U18989 (N_18989,N_13112,N_11916);
nand U18990 (N_18990,N_11415,N_14604);
and U18991 (N_18991,N_10167,N_14813);
nor U18992 (N_18992,N_11755,N_10902);
and U18993 (N_18993,N_10098,N_13243);
and U18994 (N_18994,N_13251,N_11582);
nand U18995 (N_18995,N_13908,N_13440);
and U18996 (N_18996,N_14796,N_14861);
xor U18997 (N_18997,N_10416,N_10707);
or U18998 (N_18998,N_14414,N_12863);
nand U18999 (N_18999,N_10968,N_14019);
nor U19000 (N_19000,N_11690,N_13322);
nand U19001 (N_19001,N_13383,N_13250);
nand U19002 (N_19002,N_13582,N_10929);
nand U19003 (N_19003,N_11836,N_14696);
xnor U19004 (N_19004,N_11258,N_12335);
nand U19005 (N_19005,N_14369,N_13895);
nand U19006 (N_19006,N_11242,N_10573);
or U19007 (N_19007,N_11432,N_13584);
or U19008 (N_19008,N_14815,N_10017);
and U19009 (N_19009,N_13492,N_14205);
or U19010 (N_19010,N_14857,N_13080);
and U19011 (N_19011,N_14860,N_10630);
or U19012 (N_19012,N_13426,N_10547);
and U19013 (N_19013,N_13249,N_14276);
nor U19014 (N_19014,N_12247,N_14309);
and U19015 (N_19015,N_11429,N_12592);
or U19016 (N_19016,N_12118,N_12569);
xor U19017 (N_19017,N_11257,N_13559);
xnor U19018 (N_19018,N_13091,N_12119);
xor U19019 (N_19019,N_12724,N_14254);
or U19020 (N_19020,N_10197,N_12389);
nand U19021 (N_19021,N_13733,N_10483);
and U19022 (N_19022,N_12185,N_13947);
nand U19023 (N_19023,N_12717,N_13945);
or U19024 (N_19024,N_11361,N_13357);
nand U19025 (N_19025,N_10520,N_11992);
nand U19026 (N_19026,N_14766,N_10292);
and U19027 (N_19027,N_10726,N_10356);
or U19028 (N_19028,N_11975,N_14455);
nor U19029 (N_19029,N_11853,N_12173);
and U19030 (N_19030,N_11251,N_13963);
and U19031 (N_19031,N_12256,N_14628);
xnor U19032 (N_19032,N_13050,N_12773);
and U19033 (N_19033,N_11001,N_11239);
nor U19034 (N_19034,N_12019,N_11415);
nand U19035 (N_19035,N_10651,N_11911);
nor U19036 (N_19036,N_13348,N_10962);
and U19037 (N_19037,N_14053,N_10639);
nand U19038 (N_19038,N_14941,N_13097);
nand U19039 (N_19039,N_14001,N_14195);
nand U19040 (N_19040,N_10735,N_10914);
or U19041 (N_19041,N_11019,N_11097);
nand U19042 (N_19042,N_12708,N_13376);
and U19043 (N_19043,N_10083,N_13919);
nor U19044 (N_19044,N_10869,N_11648);
nand U19045 (N_19045,N_14020,N_13107);
nor U19046 (N_19046,N_11178,N_12013);
nor U19047 (N_19047,N_13557,N_13377);
nor U19048 (N_19048,N_13678,N_14731);
nand U19049 (N_19049,N_12155,N_11260);
nor U19050 (N_19050,N_12173,N_12571);
nor U19051 (N_19051,N_14045,N_11530);
or U19052 (N_19052,N_10614,N_13648);
and U19053 (N_19053,N_10926,N_12515);
and U19054 (N_19054,N_14776,N_12100);
xnor U19055 (N_19055,N_12926,N_13703);
nand U19056 (N_19056,N_10086,N_10804);
xor U19057 (N_19057,N_13753,N_14399);
nor U19058 (N_19058,N_12224,N_11635);
and U19059 (N_19059,N_10362,N_12130);
nor U19060 (N_19060,N_13549,N_12534);
xor U19061 (N_19061,N_10244,N_11772);
nand U19062 (N_19062,N_13429,N_12203);
and U19063 (N_19063,N_14264,N_11473);
or U19064 (N_19064,N_11763,N_10006);
nor U19065 (N_19065,N_10116,N_13773);
nor U19066 (N_19066,N_10055,N_13172);
nor U19067 (N_19067,N_12644,N_14106);
xor U19068 (N_19068,N_11877,N_14527);
or U19069 (N_19069,N_13364,N_14026);
nand U19070 (N_19070,N_14601,N_10877);
or U19071 (N_19071,N_14311,N_13533);
nand U19072 (N_19072,N_10992,N_11051);
or U19073 (N_19073,N_10411,N_11425);
nor U19074 (N_19074,N_10655,N_14362);
or U19075 (N_19075,N_14170,N_11110);
nand U19076 (N_19076,N_11950,N_10954);
nor U19077 (N_19077,N_12344,N_11444);
xor U19078 (N_19078,N_12117,N_14221);
or U19079 (N_19079,N_14065,N_12428);
and U19080 (N_19080,N_14362,N_12276);
xor U19081 (N_19081,N_13740,N_13220);
and U19082 (N_19082,N_10197,N_11976);
or U19083 (N_19083,N_10270,N_14691);
nor U19084 (N_19084,N_10596,N_13950);
and U19085 (N_19085,N_14514,N_12666);
nor U19086 (N_19086,N_14327,N_14108);
and U19087 (N_19087,N_10819,N_13616);
and U19088 (N_19088,N_12206,N_12162);
nand U19089 (N_19089,N_11570,N_10968);
or U19090 (N_19090,N_14531,N_12158);
nand U19091 (N_19091,N_10771,N_10332);
xnor U19092 (N_19092,N_11865,N_11006);
and U19093 (N_19093,N_14532,N_12413);
nor U19094 (N_19094,N_12569,N_12404);
or U19095 (N_19095,N_12207,N_13086);
xor U19096 (N_19096,N_14948,N_10280);
and U19097 (N_19097,N_11059,N_11485);
and U19098 (N_19098,N_11060,N_10994);
or U19099 (N_19099,N_12514,N_14813);
nor U19100 (N_19100,N_10555,N_12014);
or U19101 (N_19101,N_12614,N_10379);
nor U19102 (N_19102,N_10584,N_11010);
nand U19103 (N_19103,N_11749,N_12440);
or U19104 (N_19104,N_13498,N_12866);
and U19105 (N_19105,N_10661,N_11335);
nor U19106 (N_19106,N_10604,N_10797);
nand U19107 (N_19107,N_14112,N_10448);
or U19108 (N_19108,N_14241,N_10560);
and U19109 (N_19109,N_10600,N_11623);
nor U19110 (N_19110,N_14519,N_13605);
or U19111 (N_19111,N_14456,N_12519);
nor U19112 (N_19112,N_11921,N_12996);
and U19113 (N_19113,N_13483,N_12256);
or U19114 (N_19114,N_10179,N_11431);
xor U19115 (N_19115,N_10457,N_12865);
or U19116 (N_19116,N_12344,N_11990);
nand U19117 (N_19117,N_11420,N_11008);
nor U19118 (N_19118,N_13954,N_12385);
xnor U19119 (N_19119,N_10806,N_14920);
nor U19120 (N_19120,N_14385,N_10192);
and U19121 (N_19121,N_11671,N_12203);
nor U19122 (N_19122,N_14576,N_11769);
nor U19123 (N_19123,N_10473,N_13151);
or U19124 (N_19124,N_10470,N_12650);
and U19125 (N_19125,N_13076,N_12202);
and U19126 (N_19126,N_14088,N_11516);
nor U19127 (N_19127,N_14238,N_13247);
nor U19128 (N_19128,N_14364,N_10772);
xnor U19129 (N_19129,N_10677,N_14763);
or U19130 (N_19130,N_13813,N_14454);
or U19131 (N_19131,N_10811,N_14150);
nand U19132 (N_19132,N_11911,N_13836);
or U19133 (N_19133,N_13539,N_12935);
xor U19134 (N_19134,N_12599,N_12781);
nand U19135 (N_19135,N_10280,N_13142);
nand U19136 (N_19136,N_11332,N_14815);
nand U19137 (N_19137,N_11301,N_13465);
nand U19138 (N_19138,N_11684,N_10455);
xor U19139 (N_19139,N_11013,N_13427);
nand U19140 (N_19140,N_11981,N_13591);
and U19141 (N_19141,N_14477,N_10401);
nor U19142 (N_19142,N_10486,N_13755);
xor U19143 (N_19143,N_14840,N_11634);
and U19144 (N_19144,N_11507,N_14005);
and U19145 (N_19145,N_14126,N_10346);
and U19146 (N_19146,N_11032,N_11328);
nor U19147 (N_19147,N_13737,N_13303);
and U19148 (N_19148,N_13404,N_12225);
nor U19149 (N_19149,N_10073,N_10167);
nor U19150 (N_19150,N_11016,N_12779);
nor U19151 (N_19151,N_12867,N_12965);
or U19152 (N_19152,N_10518,N_12000);
nand U19153 (N_19153,N_10758,N_10517);
xnor U19154 (N_19154,N_11720,N_14025);
and U19155 (N_19155,N_13340,N_11656);
and U19156 (N_19156,N_11503,N_11104);
nor U19157 (N_19157,N_14086,N_10300);
or U19158 (N_19158,N_12521,N_11860);
nor U19159 (N_19159,N_10723,N_13320);
or U19160 (N_19160,N_12008,N_11046);
and U19161 (N_19161,N_10169,N_10012);
nor U19162 (N_19162,N_14767,N_12573);
nor U19163 (N_19163,N_13097,N_14194);
xnor U19164 (N_19164,N_11291,N_10851);
nor U19165 (N_19165,N_11414,N_12525);
xnor U19166 (N_19166,N_10062,N_13325);
or U19167 (N_19167,N_11971,N_12461);
or U19168 (N_19168,N_12267,N_11073);
nor U19169 (N_19169,N_14635,N_13387);
or U19170 (N_19170,N_10529,N_10770);
or U19171 (N_19171,N_13263,N_14456);
or U19172 (N_19172,N_11419,N_12561);
nor U19173 (N_19173,N_13495,N_13838);
nor U19174 (N_19174,N_12139,N_11562);
nor U19175 (N_19175,N_10684,N_12691);
nor U19176 (N_19176,N_10724,N_10834);
nor U19177 (N_19177,N_14559,N_14579);
and U19178 (N_19178,N_10993,N_12641);
nand U19179 (N_19179,N_14638,N_14210);
and U19180 (N_19180,N_14211,N_10068);
or U19181 (N_19181,N_13660,N_12303);
nand U19182 (N_19182,N_14927,N_12962);
or U19183 (N_19183,N_13589,N_11619);
or U19184 (N_19184,N_10004,N_14858);
xor U19185 (N_19185,N_13776,N_11239);
nor U19186 (N_19186,N_12983,N_10831);
or U19187 (N_19187,N_12100,N_12730);
nand U19188 (N_19188,N_11756,N_14858);
nor U19189 (N_19189,N_10520,N_13166);
nand U19190 (N_19190,N_11933,N_11109);
nor U19191 (N_19191,N_11210,N_14486);
or U19192 (N_19192,N_11035,N_13766);
or U19193 (N_19193,N_10487,N_11497);
xor U19194 (N_19194,N_11010,N_13243);
nand U19195 (N_19195,N_10598,N_14563);
nand U19196 (N_19196,N_13946,N_13009);
xor U19197 (N_19197,N_14827,N_13415);
or U19198 (N_19198,N_10612,N_13816);
or U19199 (N_19199,N_10287,N_11622);
and U19200 (N_19200,N_12085,N_12592);
or U19201 (N_19201,N_11383,N_12260);
xnor U19202 (N_19202,N_14060,N_11045);
nor U19203 (N_19203,N_13815,N_12332);
and U19204 (N_19204,N_14270,N_10761);
nand U19205 (N_19205,N_12890,N_12109);
nor U19206 (N_19206,N_12306,N_10449);
or U19207 (N_19207,N_12246,N_11177);
nand U19208 (N_19208,N_13250,N_13977);
xor U19209 (N_19209,N_14552,N_14314);
nand U19210 (N_19210,N_11550,N_10816);
and U19211 (N_19211,N_11986,N_11673);
or U19212 (N_19212,N_11802,N_12887);
nor U19213 (N_19213,N_14511,N_11816);
and U19214 (N_19214,N_13514,N_14587);
or U19215 (N_19215,N_13414,N_13350);
nor U19216 (N_19216,N_13736,N_14898);
nand U19217 (N_19217,N_13555,N_12449);
and U19218 (N_19218,N_14422,N_12179);
nand U19219 (N_19219,N_12703,N_13852);
or U19220 (N_19220,N_12475,N_10730);
xnor U19221 (N_19221,N_12292,N_11038);
nand U19222 (N_19222,N_10106,N_14844);
nand U19223 (N_19223,N_13325,N_11217);
nand U19224 (N_19224,N_11441,N_14316);
or U19225 (N_19225,N_11938,N_12977);
or U19226 (N_19226,N_12973,N_13365);
nor U19227 (N_19227,N_11204,N_12279);
xnor U19228 (N_19228,N_12565,N_14279);
nand U19229 (N_19229,N_13029,N_10174);
nand U19230 (N_19230,N_11407,N_11362);
or U19231 (N_19231,N_13399,N_14747);
nand U19232 (N_19232,N_10700,N_13812);
nand U19233 (N_19233,N_14327,N_14540);
nor U19234 (N_19234,N_14200,N_13063);
and U19235 (N_19235,N_13166,N_13267);
nor U19236 (N_19236,N_14980,N_13645);
nand U19237 (N_19237,N_14354,N_14658);
and U19238 (N_19238,N_13031,N_12548);
or U19239 (N_19239,N_14558,N_10941);
xnor U19240 (N_19240,N_10319,N_10775);
and U19241 (N_19241,N_13195,N_13980);
nand U19242 (N_19242,N_12758,N_10519);
nand U19243 (N_19243,N_12192,N_14229);
nand U19244 (N_19244,N_12019,N_10034);
nand U19245 (N_19245,N_14819,N_12823);
nor U19246 (N_19246,N_13960,N_13437);
nand U19247 (N_19247,N_14394,N_11568);
and U19248 (N_19248,N_11550,N_11300);
nand U19249 (N_19249,N_12470,N_13800);
nand U19250 (N_19250,N_11032,N_10963);
nor U19251 (N_19251,N_13946,N_13174);
nand U19252 (N_19252,N_10535,N_13597);
nand U19253 (N_19253,N_10975,N_10278);
and U19254 (N_19254,N_12371,N_13200);
nor U19255 (N_19255,N_12900,N_13484);
and U19256 (N_19256,N_10449,N_14654);
or U19257 (N_19257,N_14574,N_14542);
nand U19258 (N_19258,N_14076,N_14820);
nor U19259 (N_19259,N_12858,N_10086);
nand U19260 (N_19260,N_10932,N_12261);
nand U19261 (N_19261,N_13796,N_14085);
nand U19262 (N_19262,N_14667,N_13210);
nor U19263 (N_19263,N_10156,N_11111);
nor U19264 (N_19264,N_14030,N_11875);
xnor U19265 (N_19265,N_11800,N_10686);
or U19266 (N_19266,N_11870,N_11305);
nor U19267 (N_19267,N_10808,N_14918);
nor U19268 (N_19268,N_14867,N_11664);
and U19269 (N_19269,N_14533,N_10474);
and U19270 (N_19270,N_14247,N_13908);
or U19271 (N_19271,N_11869,N_14064);
or U19272 (N_19272,N_10988,N_12880);
or U19273 (N_19273,N_13045,N_12040);
nand U19274 (N_19274,N_13810,N_14340);
or U19275 (N_19275,N_13122,N_12909);
or U19276 (N_19276,N_13643,N_12817);
nor U19277 (N_19277,N_10182,N_12454);
nand U19278 (N_19278,N_10835,N_12244);
and U19279 (N_19279,N_14644,N_10215);
nand U19280 (N_19280,N_12422,N_10355);
and U19281 (N_19281,N_14204,N_12849);
xnor U19282 (N_19282,N_13836,N_11400);
nor U19283 (N_19283,N_11272,N_14798);
or U19284 (N_19284,N_14836,N_11729);
and U19285 (N_19285,N_10207,N_10937);
and U19286 (N_19286,N_10567,N_11466);
nor U19287 (N_19287,N_11259,N_13819);
nand U19288 (N_19288,N_14205,N_12687);
nand U19289 (N_19289,N_10557,N_13056);
and U19290 (N_19290,N_13461,N_12435);
and U19291 (N_19291,N_13430,N_11167);
or U19292 (N_19292,N_12490,N_14323);
nor U19293 (N_19293,N_12889,N_13087);
nor U19294 (N_19294,N_10374,N_12774);
nor U19295 (N_19295,N_10020,N_13663);
xnor U19296 (N_19296,N_10247,N_14716);
and U19297 (N_19297,N_12549,N_14304);
nand U19298 (N_19298,N_14943,N_12433);
nor U19299 (N_19299,N_13851,N_10308);
nand U19300 (N_19300,N_14279,N_12635);
nand U19301 (N_19301,N_14722,N_14058);
and U19302 (N_19302,N_13203,N_13145);
nand U19303 (N_19303,N_13475,N_11159);
xnor U19304 (N_19304,N_10981,N_11704);
or U19305 (N_19305,N_12470,N_10712);
or U19306 (N_19306,N_10627,N_10679);
nand U19307 (N_19307,N_12593,N_12696);
or U19308 (N_19308,N_11370,N_10006);
nor U19309 (N_19309,N_12757,N_14105);
nor U19310 (N_19310,N_10652,N_12497);
nor U19311 (N_19311,N_12858,N_14047);
xor U19312 (N_19312,N_14578,N_14048);
nand U19313 (N_19313,N_10539,N_12605);
or U19314 (N_19314,N_14134,N_12490);
or U19315 (N_19315,N_11731,N_12463);
xor U19316 (N_19316,N_11854,N_11008);
and U19317 (N_19317,N_10126,N_13421);
nand U19318 (N_19318,N_12663,N_13350);
xnor U19319 (N_19319,N_14783,N_11816);
or U19320 (N_19320,N_14148,N_10997);
xor U19321 (N_19321,N_10665,N_14860);
nand U19322 (N_19322,N_13352,N_14391);
or U19323 (N_19323,N_13075,N_13009);
or U19324 (N_19324,N_12518,N_13440);
and U19325 (N_19325,N_12246,N_14576);
nor U19326 (N_19326,N_11359,N_14900);
or U19327 (N_19327,N_12535,N_12489);
nand U19328 (N_19328,N_12347,N_11127);
nor U19329 (N_19329,N_10442,N_12652);
or U19330 (N_19330,N_12582,N_12089);
nor U19331 (N_19331,N_13308,N_11261);
nor U19332 (N_19332,N_10753,N_10535);
nand U19333 (N_19333,N_14979,N_12906);
nand U19334 (N_19334,N_14707,N_11323);
xnor U19335 (N_19335,N_12465,N_14204);
nor U19336 (N_19336,N_10856,N_11147);
and U19337 (N_19337,N_11886,N_12182);
and U19338 (N_19338,N_10285,N_14780);
nor U19339 (N_19339,N_14998,N_11091);
nand U19340 (N_19340,N_10993,N_12043);
nor U19341 (N_19341,N_11600,N_14112);
or U19342 (N_19342,N_11077,N_11519);
and U19343 (N_19343,N_12113,N_11930);
and U19344 (N_19344,N_10490,N_10903);
nand U19345 (N_19345,N_14449,N_10645);
nor U19346 (N_19346,N_14246,N_12723);
nor U19347 (N_19347,N_10121,N_14445);
and U19348 (N_19348,N_12884,N_10397);
nand U19349 (N_19349,N_12768,N_14604);
and U19350 (N_19350,N_13773,N_10005);
and U19351 (N_19351,N_12956,N_12681);
nand U19352 (N_19352,N_10769,N_14863);
or U19353 (N_19353,N_10074,N_14205);
xor U19354 (N_19354,N_12536,N_13510);
nand U19355 (N_19355,N_13313,N_10781);
nor U19356 (N_19356,N_11978,N_10805);
xnor U19357 (N_19357,N_12001,N_14356);
and U19358 (N_19358,N_13163,N_14229);
nor U19359 (N_19359,N_13931,N_14845);
nor U19360 (N_19360,N_11581,N_11901);
or U19361 (N_19361,N_10722,N_13151);
nand U19362 (N_19362,N_13873,N_14861);
and U19363 (N_19363,N_13888,N_14033);
xor U19364 (N_19364,N_14089,N_14107);
nand U19365 (N_19365,N_11117,N_10230);
and U19366 (N_19366,N_11125,N_14997);
nor U19367 (N_19367,N_14572,N_11313);
and U19368 (N_19368,N_12845,N_14126);
nor U19369 (N_19369,N_11978,N_12957);
nand U19370 (N_19370,N_12502,N_10737);
and U19371 (N_19371,N_12263,N_14153);
nor U19372 (N_19372,N_12784,N_13672);
and U19373 (N_19373,N_12105,N_12734);
nand U19374 (N_19374,N_10489,N_13303);
or U19375 (N_19375,N_14022,N_10897);
nor U19376 (N_19376,N_10499,N_12282);
nor U19377 (N_19377,N_14760,N_11305);
or U19378 (N_19378,N_11039,N_10272);
nor U19379 (N_19379,N_13366,N_14282);
xnor U19380 (N_19380,N_13533,N_10499);
or U19381 (N_19381,N_12076,N_12996);
or U19382 (N_19382,N_13547,N_13109);
nor U19383 (N_19383,N_10152,N_11600);
or U19384 (N_19384,N_14055,N_13329);
nor U19385 (N_19385,N_13310,N_12961);
and U19386 (N_19386,N_10097,N_12217);
or U19387 (N_19387,N_11063,N_14841);
or U19388 (N_19388,N_11080,N_14799);
or U19389 (N_19389,N_13549,N_13579);
and U19390 (N_19390,N_11351,N_13324);
or U19391 (N_19391,N_11902,N_13487);
xor U19392 (N_19392,N_11564,N_13649);
nand U19393 (N_19393,N_12116,N_11913);
and U19394 (N_19394,N_10044,N_11559);
nand U19395 (N_19395,N_12763,N_12660);
nor U19396 (N_19396,N_11912,N_13509);
nand U19397 (N_19397,N_14857,N_13621);
or U19398 (N_19398,N_13465,N_13639);
and U19399 (N_19399,N_13522,N_12879);
or U19400 (N_19400,N_13100,N_10343);
nor U19401 (N_19401,N_11278,N_11297);
nand U19402 (N_19402,N_14986,N_11794);
and U19403 (N_19403,N_12166,N_10569);
and U19404 (N_19404,N_12105,N_11221);
or U19405 (N_19405,N_11508,N_10125);
and U19406 (N_19406,N_11119,N_13102);
or U19407 (N_19407,N_12286,N_13224);
nor U19408 (N_19408,N_11463,N_13648);
or U19409 (N_19409,N_14907,N_13794);
nand U19410 (N_19410,N_12734,N_12704);
nand U19411 (N_19411,N_10425,N_14495);
nor U19412 (N_19412,N_12475,N_12161);
nor U19413 (N_19413,N_11709,N_14148);
and U19414 (N_19414,N_10779,N_14422);
nand U19415 (N_19415,N_14978,N_10884);
nor U19416 (N_19416,N_11594,N_14969);
nor U19417 (N_19417,N_11352,N_14627);
nand U19418 (N_19418,N_11192,N_14710);
nand U19419 (N_19419,N_10707,N_12936);
and U19420 (N_19420,N_12198,N_11462);
xnor U19421 (N_19421,N_13707,N_12933);
nand U19422 (N_19422,N_10785,N_14491);
xnor U19423 (N_19423,N_11795,N_10787);
nand U19424 (N_19424,N_12335,N_12290);
and U19425 (N_19425,N_12845,N_13347);
and U19426 (N_19426,N_14869,N_14472);
or U19427 (N_19427,N_12920,N_14532);
or U19428 (N_19428,N_10235,N_10572);
nor U19429 (N_19429,N_14451,N_10763);
or U19430 (N_19430,N_13702,N_13056);
nand U19431 (N_19431,N_14920,N_10887);
xor U19432 (N_19432,N_14140,N_14325);
or U19433 (N_19433,N_11579,N_13289);
or U19434 (N_19434,N_12235,N_14740);
and U19435 (N_19435,N_12517,N_13454);
xnor U19436 (N_19436,N_13761,N_11149);
and U19437 (N_19437,N_12400,N_11043);
and U19438 (N_19438,N_13683,N_12054);
or U19439 (N_19439,N_13621,N_14078);
nand U19440 (N_19440,N_14059,N_14655);
or U19441 (N_19441,N_13754,N_14652);
nand U19442 (N_19442,N_12250,N_14246);
nor U19443 (N_19443,N_12638,N_14085);
or U19444 (N_19444,N_13305,N_12069);
or U19445 (N_19445,N_12609,N_11450);
or U19446 (N_19446,N_14025,N_10403);
nand U19447 (N_19447,N_13893,N_13417);
or U19448 (N_19448,N_12631,N_11542);
and U19449 (N_19449,N_14583,N_14436);
nor U19450 (N_19450,N_13575,N_10900);
nand U19451 (N_19451,N_12870,N_11507);
or U19452 (N_19452,N_14178,N_13852);
nand U19453 (N_19453,N_13133,N_13907);
or U19454 (N_19454,N_13282,N_14024);
nand U19455 (N_19455,N_14028,N_10669);
and U19456 (N_19456,N_10886,N_14527);
nor U19457 (N_19457,N_13166,N_14538);
and U19458 (N_19458,N_10249,N_11097);
and U19459 (N_19459,N_11868,N_10984);
nor U19460 (N_19460,N_14012,N_13241);
nor U19461 (N_19461,N_10492,N_11129);
nor U19462 (N_19462,N_12589,N_11584);
nor U19463 (N_19463,N_14728,N_12674);
nor U19464 (N_19464,N_11453,N_12767);
or U19465 (N_19465,N_11797,N_13813);
nor U19466 (N_19466,N_10544,N_10106);
and U19467 (N_19467,N_12337,N_12447);
and U19468 (N_19468,N_11459,N_14048);
or U19469 (N_19469,N_14106,N_13021);
nor U19470 (N_19470,N_10328,N_13065);
nand U19471 (N_19471,N_12298,N_11832);
or U19472 (N_19472,N_12677,N_14855);
nor U19473 (N_19473,N_12098,N_11525);
nand U19474 (N_19474,N_10271,N_13222);
or U19475 (N_19475,N_11853,N_13606);
xnor U19476 (N_19476,N_10688,N_13264);
or U19477 (N_19477,N_13984,N_12539);
or U19478 (N_19478,N_11332,N_10422);
nand U19479 (N_19479,N_13679,N_13419);
or U19480 (N_19480,N_13099,N_12581);
and U19481 (N_19481,N_10566,N_13717);
nand U19482 (N_19482,N_11088,N_14077);
nor U19483 (N_19483,N_13815,N_12956);
or U19484 (N_19484,N_13659,N_13761);
and U19485 (N_19485,N_12433,N_12760);
nand U19486 (N_19486,N_14051,N_14227);
or U19487 (N_19487,N_10619,N_13840);
or U19488 (N_19488,N_12654,N_11791);
nand U19489 (N_19489,N_11521,N_14120);
nand U19490 (N_19490,N_10360,N_12839);
nor U19491 (N_19491,N_14124,N_12867);
nand U19492 (N_19492,N_13964,N_13376);
nand U19493 (N_19493,N_11337,N_14243);
or U19494 (N_19494,N_12820,N_11780);
nand U19495 (N_19495,N_12599,N_11270);
and U19496 (N_19496,N_10923,N_10229);
xor U19497 (N_19497,N_12837,N_12390);
and U19498 (N_19498,N_14948,N_12314);
and U19499 (N_19499,N_10578,N_10850);
and U19500 (N_19500,N_10174,N_11346);
nand U19501 (N_19501,N_11656,N_11427);
nor U19502 (N_19502,N_13041,N_12595);
or U19503 (N_19503,N_11601,N_11498);
or U19504 (N_19504,N_11120,N_11387);
nor U19505 (N_19505,N_10233,N_12435);
and U19506 (N_19506,N_13947,N_10912);
nor U19507 (N_19507,N_13457,N_12764);
nor U19508 (N_19508,N_10534,N_12536);
and U19509 (N_19509,N_12826,N_10967);
and U19510 (N_19510,N_14137,N_13715);
or U19511 (N_19511,N_10127,N_14406);
nand U19512 (N_19512,N_13500,N_11901);
and U19513 (N_19513,N_12074,N_14341);
and U19514 (N_19514,N_13998,N_12321);
nor U19515 (N_19515,N_13076,N_14681);
xor U19516 (N_19516,N_11215,N_11951);
or U19517 (N_19517,N_12620,N_13884);
or U19518 (N_19518,N_13393,N_13448);
nor U19519 (N_19519,N_11449,N_14017);
nand U19520 (N_19520,N_11039,N_11973);
and U19521 (N_19521,N_10157,N_11495);
nor U19522 (N_19522,N_12923,N_10771);
nor U19523 (N_19523,N_13552,N_10694);
nand U19524 (N_19524,N_14847,N_10722);
nor U19525 (N_19525,N_11590,N_11288);
and U19526 (N_19526,N_10741,N_12638);
nand U19527 (N_19527,N_12303,N_14720);
xnor U19528 (N_19528,N_12975,N_14063);
and U19529 (N_19529,N_14440,N_13937);
and U19530 (N_19530,N_12728,N_10846);
xor U19531 (N_19531,N_12420,N_10624);
xnor U19532 (N_19532,N_11796,N_14884);
nand U19533 (N_19533,N_14290,N_14477);
nand U19534 (N_19534,N_10758,N_14982);
and U19535 (N_19535,N_10801,N_14072);
xor U19536 (N_19536,N_11409,N_13453);
or U19537 (N_19537,N_11285,N_13979);
or U19538 (N_19538,N_10247,N_10554);
or U19539 (N_19539,N_13945,N_11028);
nor U19540 (N_19540,N_11796,N_10337);
or U19541 (N_19541,N_10611,N_10659);
nand U19542 (N_19542,N_14628,N_12934);
nor U19543 (N_19543,N_12108,N_14880);
or U19544 (N_19544,N_11407,N_14781);
nand U19545 (N_19545,N_14013,N_14414);
nor U19546 (N_19546,N_11702,N_12813);
nor U19547 (N_19547,N_10262,N_11156);
nand U19548 (N_19548,N_13643,N_13563);
nor U19549 (N_19549,N_13434,N_13572);
and U19550 (N_19550,N_12646,N_11205);
and U19551 (N_19551,N_14077,N_12851);
xor U19552 (N_19552,N_11783,N_14535);
and U19553 (N_19553,N_13915,N_10083);
nor U19554 (N_19554,N_14989,N_12140);
nand U19555 (N_19555,N_10626,N_13875);
nor U19556 (N_19556,N_13693,N_10096);
nor U19557 (N_19557,N_13345,N_10263);
or U19558 (N_19558,N_11480,N_11902);
xnor U19559 (N_19559,N_14537,N_13627);
nor U19560 (N_19560,N_10440,N_12588);
or U19561 (N_19561,N_11381,N_11729);
nor U19562 (N_19562,N_14033,N_13253);
nand U19563 (N_19563,N_14740,N_10230);
and U19564 (N_19564,N_10190,N_11355);
nor U19565 (N_19565,N_10059,N_11500);
nand U19566 (N_19566,N_14497,N_11108);
nor U19567 (N_19567,N_14746,N_14529);
and U19568 (N_19568,N_11908,N_13723);
nand U19569 (N_19569,N_11126,N_12151);
nand U19570 (N_19570,N_13977,N_12207);
nand U19571 (N_19571,N_14968,N_11220);
nor U19572 (N_19572,N_14074,N_10722);
or U19573 (N_19573,N_11978,N_11399);
or U19574 (N_19574,N_14647,N_13366);
nor U19575 (N_19575,N_13930,N_12119);
nand U19576 (N_19576,N_14974,N_12557);
and U19577 (N_19577,N_14950,N_11589);
xnor U19578 (N_19578,N_11967,N_10217);
nor U19579 (N_19579,N_14544,N_14813);
and U19580 (N_19580,N_12679,N_12331);
nand U19581 (N_19581,N_10336,N_11754);
nand U19582 (N_19582,N_11866,N_11885);
nand U19583 (N_19583,N_12726,N_10800);
or U19584 (N_19584,N_13050,N_10563);
and U19585 (N_19585,N_14864,N_14000);
and U19586 (N_19586,N_10351,N_11109);
xnor U19587 (N_19587,N_12013,N_11334);
or U19588 (N_19588,N_11605,N_10874);
and U19589 (N_19589,N_11616,N_12591);
nand U19590 (N_19590,N_14165,N_14096);
xor U19591 (N_19591,N_13360,N_10846);
nor U19592 (N_19592,N_12243,N_12436);
nor U19593 (N_19593,N_10712,N_12856);
or U19594 (N_19594,N_10164,N_10046);
nand U19595 (N_19595,N_10585,N_11012);
nand U19596 (N_19596,N_10242,N_11100);
nor U19597 (N_19597,N_11909,N_12006);
or U19598 (N_19598,N_12324,N_14494);
nand U19599 (N_19599,N_13179,N_12980);
or U19600 (N_19600,N_11431,N_10455);
and U19601 (N_19601,N_13844,N_14687);
nor U19602 (N_19602,N_13964,N_11117);
xnor U19603 (N_19603,N_13033,N_12810);
nand U19604 (N_19604,N_12909,N_12399);
nor U19605 (N_19605,N_14991,N_14772);
and U19606 (N_19606,N_12372,N_14178);
or U19607 (N_19607,N_11178,N_14531);
nand U19608 (N_19608,N_11924,N_13656);
or U19609 (N_19609,N_13855,N_13939);
and U19610 (N_19610,N_12034,N_11465);
nor U19611 (N_19611,N_12324,N_11598);
and U19612 (N_19612,N_13596,N_13896);
or U19613 (N_19613,N_12327,N_14128);
and U19614 (N_19614,N_10950,N_14934);
nand U19615 (N_19615,N_11314,N_13212);
or U19616 (N_19616,N_12691,N_12681);
nor U19617 (N_19617,N_12845,N_12030);
nor U19618 (N_19618,N_13823,N_12624);
nand U19619 (N_19619,N_13443,N_13164);
nor U19620 (N_19620,N_11631,N_10559);
xnor U19621 (N_19621,N_13415,N_10855);
and U19622 (N_19622,N_10003,N_12445);
nand U19623 (N_19623,N_12293,N_12933);
and U19624 (N_19624,N_14174,N_14441);
and U19625 (N_19625,N_14257,N_11625);
nand U19626 (N_19626,N_11451,N_13331);
nor U19627 (N_19627,N_10061,N_12670);
or U19628 (N_19628,N_12326,N_13155);
nor U19629 (N_19629,N_11330,N_11548);
xnor U19630 (N_19630,N_13292,N_12423);
nor U19631 (N_19631,N_11202,N_13983);
nand U19632 (N_19632,N_13017,N_13720);
xor U19633 (N_19633,N_14195,N_10569);
and U19634 (N_19634,N_14788,N_11992);
and U19635 (N_19635,N_10783,N_13502);
and U19636 (N_19636,N_13367,N_10388);
nor U19637 (N_19637,N_12603,N_13224);
nand U19638 (N_19638,N_12427,N_11551);
nor U19639 (N_19639,N_14598,N_14055);
and U19640 (N_19640,N_11652,N_12816);
or U19641 (N_19641,N_11189,N_11645);
nor U19642 (N_19642,N_11759,N_12259);
nand U19643 (N_19643,N_10285,N_11340);
or U19644 (N_19644,N_10243,N_11243);
and U19645 (N_19645,N_14945,N_10311);
xor U19646 (N_19646,N_11190,N_11983);
xor U19647 (N_19647,N_12351,N_10570);
and U19648 (N_19648,N_13893,N_12524);
and U19649 (N_19649,N_10318,N_13331);
nand U19650 (N_19650,N_10895,N_14825);
and U19651 (N_19651,N_14213,N_11973);
nor U19652 (N_19652,N_12991,N_14121);
nand U19653 (N_19653,N_12692,N_14509);
or U19654 (N_19654,N_11147,N_13163);
nand U19655 (N_19655,N_11463,N_13839);
and U19656 (N_19656,N_12050,N_13036);
and U19657 (N_19657,N_11187,N_10196);
nand U19658 (N_19658,N_13484,N_10242);
and U19659 (N_19659,N_13315,N_12786);
and U19660 (N_19660,N_13344,N_13311);
nor U19661 (N_19661,N_12891,N_10119);
and U19662 (N_19662,N_14909,N_13293);
or U19663 (N_19663,N_14659,N_14202);
nor U19664 (N_19664,N_10693,N_12666);
nor U19665 (N_19665,N_12547,N_10339);
nor U19666 (N_19666,N_14125,N_10586);
or U19667 (N_19667,N_14769,N_13207);
xnor U19668 (N_19668,N_13884,N_14194);
or U19669 (N_19669,N_12443,N_11114);
and U19670 (N_19670,N_11745,N_12378);
xnor U19671 (N_19671,N_12092,N_14010);
or U19672 (N_19672,N_10273,N_12557);
xnor U19673 (N_19673,N_13733,N_11587);
and U19674 (N_19674,N_14717,N_13086);
nor U19675 (N_19675,N_14610,N_12126);
and U19676 (N_19676,N_12218,N_11382);
or U19677 (N_19677,N_14234,N_14676);
nor U19678 (N_19678,N_12362,N_11006);
or U19679 (N_19679,N_12843,N_13979);
and U19680 (N_19680,N_12027,N_10315);
or U19681 (N_19681,N_13881,N_13659);
nand U19682 (N_19682,N_13839,N_13629);
xor U19683 (N_19683,N_13589,N_11006);
or U19684 (N_19684,N_12856,N_12663);
nand U19685 (N_19685,N_14625,N_10347);
and U19686 (N_19686,N_13340,N_13466);
and U19687 (N_19687,N_13364,N_12280);
xor U19688 (N_19688,N_12656,N_10530);
or U19689 (N_19689,N_10976,N_13905);
nor U19690 (N_19690,N_14243,N_10695);
nand U19691 (N_19691,N_11605,N_13298);
nor U19692 (N_19692,N_13743,N_11990);
and U19693 (N_19693,N_11103,N_10311);
nor U19694 (N_19694,N_11122,N_13229);
nand U19695 (N_19695,N_14972,N_14588);
nand U19696 (N_19696,N_14510,N_10455);
or U19697 (N_19697,N_12284,N_12632);
nor U19698 (N_19698,N_13188,N_10318);
and U19699 (N_19699,N_12165,N_14401);
xnor U19700 (N_19700,N_14774,N_10663);
nand U19701 (N_19701,N_12699,N_14391);
or U19702 (N_19702,N_11270,N_14827);
nand U19703 (N_19703,N_11049,N_13035);
nor U19704 (N_19704,N_10896,N_12683);
or U19705 (N_19705,N_12330,N_14718);
nand U19706 (N_19706,N_13574,N_12795);
nand U19707 (N_19707,N_10957,N_13659);
nand U19708 (N_19708,N_13925,N_11555);
and U19709 (N_19709,N_10369,N_10954);
nand U19710 (N_19710,N_12891,N_13807);
or U19711 (N_19711,N_10609,N_11525);
xor U19712 (N_19712,N_12353,N_10273);
nand U19713 (N_19713,N_12782,N_11688);
and U19714 (N_19714,N_11344,N_10797);
and U19715 (N_19715,N_12829,N_13218);
nand U19716 (N_19716,N_11876,N_11407);
nor U19717 (N_19717,N_13101,N_14989);
nand U19718 (N_19718,N_13403,N_13476);
and U19719 (N_19719,N_11294,N_11061);
nand U19720 (N_19720,N_10885,N_13211);
xnor U19721 (N_19721,N_13394,N_12038);
xor U19722 (N_19722,N_11659,N_11093);
nor U19723 (N_19723,N_13982,N_14203);
or U19724 (N_19724,N_14299,N_12519);
and U19725 (N_19725,N_10744,N_13017);
and U19726 (N_19726,N_10121,N_10529);
or U19727 (N_19727,N_13331,N_11098);
or U19728 (N_19728,N_10514,N_12564);
and U19729 (N_19729,N_12513,N_13577);
xnor U19730 (N_19730,N_10966,N_13001);
nand U19731 (N_19731,N_10677,N_12144);
xor U19732 (N_19732,N_10249,N_14101);
or U19733 (N_19733,N_11455,N_13237);
and U19734 (N_19734,N_10147,N_13292);
nor U19735 (N_19735,N_11667,N_12852);
or U19736 (N_19736,N_13374,N_10358);
and U19737 (N_19737,N_10929,N_13431);
nand U19738 (N_19738,N_13105,N_11862);
nor U19739 (N_19739,N_14607,N_14309);
or U19740 (N_19740,N_14806,N_10389);
and U19741 (N_19741,N_11808,N_13400);
nand U19742 (N_19742,N_13491,N_11724);
nand U19743 (N_19743,N_13263,N_13397);
or U19744 (N_19744,N_13660,N_11868);
and U19745 (N_19745,N_11673,N_13034);
or U19746 (N_19746,N_14984,N_11238);
nor U19747 (N_19747,N_11281,N_14096);
nand U19748 (N_19748,N_10134,N_10486);
nor U19749 (N_19749,N_13887,N_11795);
and U19750 (N_19750,N_12145,N_10936);
or U19751 (N_19751,N_10069,N_11014);
nor U19752 (N_19752,N_12265,N_12523);
or U19753 (N_19753,N_12356,N_13914);
and U19754 (N_19754,N_13278,N_14942);
and U19755 (N_19755,N_14970,N_13237);
or U19756 (N_19756,N_12062,N_10494);
and U19757 (N_19757,N_11737,N_14545);
or U19758 (N_19758,N_10166,N_12479);
and U19759 (N_19759,N_10030,N_11020);
nand U19760 (N_19760,N_11174,N_12912);
or U19761 (N_19761,N_10646,N_13931);
or U19762 (N_19762,N_10164,N_14447);
and U19763 (N_19763,N_14510,N_14420);
nor U19764 (N_19764,N_14848,N_10711);
nand U19765 (N_19765,N_12775,N_10431);
xnor U19766 (N_19766,N_12746,N_14457);
and U19767 (N_19767,N_10004,N_14695);
xor U19768 (N_19768,N_14095,N_12817);
xor U19769 (N_19769,N_13288,N_14050);
nor U19770 (N_19770,N_14083,N_13730);
nor U19771 (N_19771,N_11618,N_13171);
or U19772 (N_19772,N_12015,N_12059);
xor U19773 (N_19773,N_10058,N_11495);
or U19774 (N_19774,N_14056,N_13741);
xor U19775 (N_19775,N_13031,N_10823);
nand U19776 (N_19776,N_14166,N_14499);
nor U19777 (N_19777,N_11993,N_13207);
or U19778 (N_19778,N_14214,N_11126);
and U19779 (N_19779,N_14249,N_10336);
and U19780 (N_19780,N_11426,N_14061);
nor U19781 (N_19781,N_10129,N_11496);
nand U19782 (N_19782,N_11859,N_14567);
or U19783 (N_19783,N_11533,N_10930);
nor U19784 (N_19784,N_13277,N_12666);
nor U19785 (N_19785,N_13863,N_13413);
and U19786 (N_19786,N_12785,N_13709);
nand U19787 (N_19787,N_12199,N_13104);
or U19788 (N_19788,N_14774,N_11523);
nor U19789 (N_19789,N_14431,N_14687);
xnor U19790 (N_19790,N_14491,N_12025);
and U19791 (N_19791,N_14783,N_10051);
nor U19792 (N_19792,N_10007,N_13078);
or U19793 (N_19793,N_10808,N_11324);
or U19794 (N_19794,N_11601,N_11225);
and U19795 (N_19795,N_13816,N_11476);
and U19796 (N_19796,N_12570,N_10004);
and U19797 (N_19797,N_12994,N_14623);
nor U19798 (N_19798,N_13293,N_11936);
nand U19799 (N_19799,N_14519,N_11775);
or U19800 (N_19800,N_12056,N_12969);
nand U19801 (N_19801,N_11071,N_11434);
nand U19802 (N_19802,N_13951,N_10533);
nand U19803 (N_19803,N_14129,N_10310);
nand U19804 (N_19804,N_12873,N_14657);
nand U19805 (N_19805,N_13712,N_10055);
nor U19806 (N_19806,N_11660,N_11526);
xnor U19807 (N_19807,N_11793,N_11745);
nor U19808 (N_19808,N_11210,N_10694);
and U19809 (N_19809,N_12079,N_10514);
nand U19810 (N_19810,N_14503,N_11106);
nand U19811 (N_19811,N_13462,N_11443);
nand U19812 (N_19812,N_11480,N_12276);
nand U19813 (N_19813,N_11221,N_12023);
and U19814 (N_19814,N_13195,N_10736);
nor U19815 (N_19815,N_11736,N_12070);
and U19816 (N_19816,N_10727,N_10508);
or U19817 (N_19817,N_11752,N_12528);
nand U19818 (N_19818,N_13971,N_14531);
or U19819 (N_19819,N_14576,N_12677);
nor U19820 (N_19820,N_10962,N_10465);
or U19821 (N_19821,N_11724,N_12768);
or U19822 (N_19822,N_13164,N_10030);
xnor U19823 (N_19823,N_14951,N_14755);
xor U19824 (N_19824,N_10912,N_14215);
xnor U19825 (N_19825,N_12937,N_10284);
xnor U19826 (N_19826,N_14223,N_13358);
nand U19827 (N_19827,N_13680,N_14366);
or U19828 (N_19828,N_10467,N_12218);
nand U19829 (N_19829,N_10482,N_13270);
nor U19830 (N_19830,N_12252,N_11315);
or U19831 (N_19831,N_14876,N_13002);
nor U19832 (N_19832,N_14696,N_11783);
nand U19833 (N_19833,N_13379,N_10551);
nor U19834 (N_19834,N_12296,N_10342);
nand U19835 (N_19835,N_14188,N_11313);
or U19836 (N_19836,N_13429,N_10719);
and U19837 (N_19837,N_13120,N_14827);
and U19838 (N_19838,N_14946,N_11419);
or U19839 (N_19839,N_14056,N_11334);
and U19840 (N_19840,N_11733,N_10825);
nor U19841 (N_19841,N_10455,N_11004);
or U19842 (N_19842,N_10007,N_14739);
nand U19843 (N_19843,N_12453,N_12063);
and U19844 (N_19844,N_12061,N_14457);
nand U19845 (N_19845,N_12859,N_10351);
and U19846 (N_19846,N_13811,N_14903);
nand U19847 (N_19847,N_10219,N_14814);
or U19848 (N_19848,N_12920,N_14242);
nor U19849 (N_19849,N_12529,N_14253);
and U19850 (N_19850,N_12863,N_11764);
nand U19851 (N_19851,N_14711,N_13937);
nor U19852 (N_19852,N_13881,N_14219);
and U19853 (N_19853,N_13942,N_11488);
nand U19854 (N_19854,N_14980,N_12801);
or U19855 (N_19855,N_11777,N_10165);
or U19856 (N_19856,N_12510,N_12430);
and U19857 (N_19857,N_11754,N_11424);
or U19858 (N_19858,N_11167,N_10914);
nand U19859 (N_19859,N_14834,N_11736);
and U19860 (N_19860,N_10378,N_12668);
nand U19861 (N_19861,N_10439,N_10119);
xnor U19862 (N_19862,N_11166,N_12118);
or U19863 (N_19863,N_14333,N_10032);
and U19864 (N_19864,N_12890,N_14335);
or U19865 (N_19865,N_14130,N_14341);
nand U19866 (N_19866,N_14576,N_10003);
and U19867 (N_19867,N_14868,N_11682);
or U19868 (N_19868,N_11055,N_10678);
and U19869 (N_19869,N_13690,N_14392);
and U19870 (N_19870,N_12645,N_13335);
or U19871 (N_19871,N_14880,N_10074);
nor U19872 (N_19872,N_11397,N_13470);
nor U19873 (N_19873,N_14371,N_10169);
and U19874 (N_19874,N_12807,N_12712);
nand U19875 (N_19875,N_12348,N_12567);
nand U19876 (N_19876,N_14898,N_12748);
or U19877 (N_19877,N_13692,N_12089);
nand U19878 (N_19878,N_10380,N_10522);
or U19879 (N_19879,N_12775,N_13170);
nor U19880 (N_19880,N_10895,N_12011);
and U19881 (N_19881,N_12124,N_14257);
nand U19882 (N_19882,N_10609,N_10587);
and U19883 (N_19883,N_11051,N_10766);
or U19884 (N_19884,N_11484,N_12039);
and U19885 (N_19885,N_11100,N_10429);
or U19886 (N_19886,N_14696,N_11890);
nor U19887 (N_19887,N_14105,N_12744);
or U19888 (N_19888,N_14733,N_14798);
or U19889 (N_19889,N_10256,N_10430);
nand U19890 (N_19890,N_11581,N_13601);
or U19891 (N_19891,N_13513,N_11687);
and U19892 (N_19892,N_10294,N_11084);
and U19893 (N_19893,N_10291,N_11194);
nor U19894 (N_19894,N_12152,N_13873);
or U19895 (N_19895,N_12942,N_11367);
nand U19896 (N_19896,N_13410,N_11646);
and U19897 (N_19897,N_12942,N_13044);
nor U19898 (N_19898,N_10410,N_10151);
and U19899 (N_19899,N_10095,N_10246);
nand U19900 (N_19900,N_11678,N_14179);
xor U19901 (N_19901,N_11793,N_12168);
nand U19902 (N_19902,N_14961,N_14280);
nand U19903 (N_19903,N_13126,N_12200);
and U19904 (N_19904,N_10467,N_11928);
nor U19905 (N_19905,N_13729,N_12688);
nand U19906 (N_19906,N_12111,N_11708);
nand U19907 (N_19907,N_13562,N_14810);
nand U19908 (N_19908,N_11409,N_12070);
and U19909 (N_19909,N_11480,N_11117);
nor U19910 (N_19910,N_11930,N_14060);
nor U19911 (N_19911,N_11091,N_14018);
nor U19912 (N_19912,N_11417,N_10945);
or U19913 (N_19913,N_14232,N_12122);
or U19914 (N_19914,N_13656,N_12672);
or U19915 (N_19915,N_11111,N_12877);
nand U19916 (N_19916,N_11084,N_14854);
xnor U19917 (N_19917,N_14375,N_13981);
or U19918 (N_19918,N_10032,N_10458);
nor U19919 (N_19919,N_14478,N_13713);
nand U19920 (N_19920,N_11611,N_12205);
nand U19921 (N_19921,N_14901,N_12429);
or U19922 (N_19922,N_11657,N_10380);
nor U19923 (N_19923,N_12623,N_12551);
nor U19924 (N_19924,N_11851,N_14346);
nand U19925 (N_19925,N_12071,N_12273);
or U19926 (N_19926,N_11333,N_12098);
or U19927 (N_19927,N_12756,N_12202);
xnor U19928 (N_19928,N_13566,N_10995);
or U19929 (N_19929,N_10100,N_14201);
or U19930 (N_19930,N_13071,N_10178);
and U19931 (N_19931,N_10088,N_11625);
nor U19932 (N_19932,N_11111,N_13142);
nand U19933 (N_19933,N_11489,N_10877);
or U19934 (N_19934,N_10916,N_12004);
and U19935 (N_19935,N_14668,N_13533);
nor U19936 (N_19936,N_12785,N_14575);
and U19937 (N_19937,N_10266,N_12253);
nand U19938 (N_19938,N_11193,N_13240);
nand U19939 (N_19939,N_11930,N_12025);
nand U19940 (N_19940,N_10134,N_12248);
or U19941 (N_19941,N_13066,N_12544);
and U19942 (N_19942,N_11224,N_14086);
nand U19943 (N_19943,N_14491,N_14367);
or U19944 (N_19944,N_10839,N_13911);
or U19945 (N_19945,N_11895,N_10257);
nand U19946 (N_19946,N_11960,N_10233);
and U19947 (N_19947,N_13275,N_10765);
or U19948 (N_19948,N_14237,N_12678);
or U19949 (N_19949,N_10261,N_12397);
xor U19950 (N_19950,N_14728,N_10997);
or U19951 (N_19951,N_12133,N_13638);
xnor U19952 (N_19952,N_12853,N_11968);
nor U19953 (N_19953,N_13724,N_14256);
and U19954 (N_19954,N_12691,N_12036);
or U19955 (N_19955,N_12998,N_12807);
and U19956 (N_19956,N_10023,N_13544);
nor U19957 (N_19957,N_11374,N_14428);
nor U19958 (N_19958,N_13321,N_14414);
or U19959 (N_19959,N_12674,N_12580);
nand U19960 (N_19960,N_11508,N_10727);
or U19961 (N_19961,N_10781,N_13153);
xnor U19962 (N_19962,N_10705,N_12009);
nor U19963 (N_19963,N_12573,N_14993);
and U19964 (N_19964,N_12714,N_14801);
or U19965 (N_19965,N_14315,N_13810);
nand U19966 (N_19966,N_10971,N_12347);
or U19967 (N_19967,N_11813,N_11893);
and U19968 (N_19968,N_12218,N_10124);
or U19969 (N_19969,N_13348,N_14110);
or U19970 (N_19970,N_13112,N_10464);
nand U19971 (N_19971,N_12971,N_10253);
or U19972 (N_19972,N_11492,N_14867);
nand U19973 (N_19973,N_14476,N_11167);
nor U19974 (N_19974,N_14429,N_11199);
or U19975 (N_19975,N_12405,N_10699);
nand U19976 (N_19976,N_13939,N_11821);
and U19977 (N_19977,N_13019,N_14747);
and U19978 (N_19978,N_10497,N_12692);
nor U19979 (N_19979,N_10410,N_10882);
and U19980 (N_19980,N_11534,N_11100);
nor U19981 (N_19981,N_13451,N_11956);
and U19982 (N_19982,N_14813,N_11543);
and U19983 (N_19983,N_10236,N_13773);
nand U19984 (N_19984,N_13522,N_11652);
nor U19985 (N_19985,N_10700,N_14898);
nand U19986 (N_19986,N_14621,N_14674);
xnor U19987 (N_19987,N_13917,N_14740);
and U19988 (N_19988,N_14560,N_13020);
and U19989 (N_19989,N_12232,N_13850);
nand U19990 (N_19990,N_14268,N_10219);
and U19991 (N_19991,N_13425,N_13747);
or U19992 (N_19992,N_11448,N_14184);
nor U19993 (N_19993,N_12095,N_14352);
or U19994 (N_19994,N_10677,N_14470);
or U19995 (N_19995,N_11656,N_13133);
or U19996 (N_19996,N_14612,N_12619);
or U19997 (N_19997,N_10189,N_14188);
and U19998 (N_19998,N_10704,N_11932);
xnor U19999 (N_19999,N_11654,N_14207);
or U20000 (N_20000,N_15159,N_17436);
nand U20001 (N_20001,N_15502,N_18221);
and U20002 (N_20002,N_17938,N_17060);
nor U20003 (N_20003,N_18427,N_16805);
xor U20004 (N_20004,N_18338,N_18849);
and U20005 (N_20005,N_18613,N_15060);
xor U20006 (N_20006,N_16691,N_17552);
xnor U20007 (N_20007,N_17245,N_19691);
nand U20008 (N_20008,N_18994,N_19584);
or U20009 (N_20009,N_17102,N_16948);
nor U20010 (N_20010,N_18708,N_19198);
and U20011 (N_20011,N_16186,N_17007);
and U20012 (N_20012,N_15027,N_18743);
or U20013 (N_20013,N_19719,N_15307);
nand U20014 (N_20014,N_19985,N_17066);
nand U20015 (N_20015,N_16518,N_17501);
xor U20016 (N_20016,N_18906,N_19866);
xnor U20017 (N_20017,N_18079,N_18331);
nand U20018 (N_20018,N_19552,N_19916);
or U20019 (N_20019,N_15311,N_17683);
nor U20020 (N_20020,N_17500,N_18966);
xor U20021 (N_20021,N_17379,N_15294);
and U20022 (N_20022,N_18093,N_18100);
nand U20023 (N_20023,N_19740,N_19476);
and U20024 (N_20024,N_15541,N_17125);
nand U20025 (N_20025,N_16853,N_15017);
or U20026 (N_20026,N_16574,N_17701);
xnor U20027 (N_20027,N_17016,N_15648);
xnor U20028 (N_20028,N_17283,N_15690);
and U20029 (N_20029,N_19255,N_18759);
and U20030 (N_20030,N_18362,N_19055);
and U20031 (N_20031,N_16863,N_16568);
or U20032 (N_20032,N_16940,N_17770);
xor U20033 (N_20033,N_15145,N_19414);
nor U20034 (N_20034,N_15858,N_18929);
or U20035 (N_20035,N_18406,N_17099);
and U20036 (N_20036,N_17837,N_17282);
or U20037 (N_20037,N_18762,N_17289);
nor U20038 (N_20038,N_19309,N_18777);
nand U20039 (N_20039,N_16468,N_18050);
or U20040 (N_20040,N_16992,N_19179);
nor U20041 (N_20041,N_16148,N_17943);
or U20042 (N_20042,N_19714,N_17575);
or U20043 (N_20043,N_16850,N_19911);
nor U20044 (N_20044,N_16273,N_16868);
nand U20045 (N_20045,N_17634,N_15763);
and U20046 (N_20046,N_18810,N_15567);
or U20047 (N_20047,N_16364,N_19791);
and U20048 (N_20048,N_18961,N_16341);
nor U20049 (N_20049,N_18897,N_15594);
and U20050 (N_20050,N_16284,N_16161);
nand U20051 (N_20051,N_16081,N_15949);
and U20052 (N_20052,N_15869,N_18830);
nand U20053 (N_20053,N_18788,N_15891);
or U20054 (N_20054,N_15251,N_15391);
nor U20055 (N_20055,N_19852,N_17692);
nor U20056 (N_20056,N_15987,N_17252);
or U20057 (N_20057,N_19252,N_18108);
and U20058 (N_20058,N_18448,N_18548);
or U20059 (N_20059,N_17285,N_18622);
nor U20060 (N_20060,N_16430,N_18755);
and U20061 (N_20061,N_15736,N_16881);
or U20062 (N_20062,N_17670,N_17337);
and U20063 (N_20063,N_16140,N_15865);
nor U20064 (N_20064,N_15070,N_18518);
xor U20065 (N_20065,N_15523,N_15623);
and U20066 (N_20066,N_15799,N_17246);
nor U20067 (N_20067,N_16956,N_19335);
nor U20068 (N_20068,N_15656,N_16968);
nor U20069 (N_20069,N_17328,N_15163);
nor U20070 (N_20070,N_16860,N_15128);
and U20071 (N_20071,N_18711,N_19104);
nand U20072 (N_20072,N_15469,N_15090);
or U20073 (N_20073,N_18158,N_15722);
nand U20074 (N_20074,N_18761,N_15542);
nor U20075 (N_20075,N_15728,N_19223);
nor U20076 (N_20076,N_15928,N_19537);
or U20077 (N_20077,N_19070,N_15720);
and U20078 (N_20078,N_19380,N_15224);
or U20079 (N_20079,N_16315,N_15993);
nand U20080 (N_20080,N_16587,N_18945);
and U20081 (N_20081,N_18213,N_17493);
nor U20082 (N_20082,N_16517,N_15069);
nor U20083 (N_20083,N_17030,N_19295);
nand U20084 (N_20084,N_17086,N_15777);
xor U20085 (N_20085,N_17696,N_19680);
or U20086 (N_20086,N_16338,N_15545);
nor U20087 (N_20087,N_15016,N_16055);
nand U20088 (N_20088,N_16913,N_18279);
or U20089 (N_20089,N_15305,N_17439);
and U20090 (N_20090,N_19549,N_15535);
nor U20091 (N_20091,N_16293,N_17058);
nor U20092 (N_20092,N_17921,N_15330);
nor U20093 (N_20093,N_19051,N_19043);
nor U20094 (N_20094,N_19455,N_17904);
nor U20095 (N_20095,N_18066,N_15436);
xor U20096 (N_20096,N_19562,N_19162);
nand U20097 (N_20097,N_15936,N_17796);
or U20098 (N_20098,N_19646,N_15909);
nand U20099 (N_20099,N_17843,N_19794);
nand U20100 (N_20100,N_19499,N_18299);
and U20101 (N_20101,N_18935,N_15143);
nor U20102 (N_20102,N_17602,N_16191);
or U20103 (N_20103,N_16447,N_16425);
nor U20104 (N_20104,N_17738,N_19034);
nand U20105 (N_20105,N_18414,N_17841);
nand U20106 (N_20106,N_19609,N_16949);
nor U20107 (N_20107,N_16335,N_19577);
and U20108 (N_20108,N_18956,N_19766);
and U20109 (N_20109,N_15323,N_15931);
or U20110 (N_20110,N_15361,N_16975);
or U20111 (N_20111,N_18292,N_19016);
nand U20112 (N_20112,N_18343,N_17717);
or U20113 (N_20113,N_15009,N_19767);
nand U20114 (N_20114,N_15137,N_18684);
or U20115 (N_20115,N_18582,N_15636);
and U20116 (N_20116,N_18317,N_15024);
or U20117 (N_20117,N_15902,N_18649);
or U20118 (N_20118,N_15446,N_18899);
xnor U20119 (N_20119,N_15908,N_16365);
nor U20120 (N_20120,N_17533,N_18545);
or U20121 (N_20121,N_19156,N_17885);
nor U20122 (N_20122,N_18220,N_16264);
nand U20123 (N_20123,N_16946,N_19385);
nand U20124 (N_20124,N_17234,N_19005);
and U20125 (N_20125,N_16229,N_15553);
nor U20126 (N_20126,N_18655,N_18997);
nor U20127 (N_20127,N_19987,N_19582);
nor U20128 (N_20128,N_16785,N_19910);
or U20129 (N_20129,N_16352,N_16433);
nor U20130 (N_20130,N_18462,N_15444);
nor U20131 (N_20131,N_18578,N_17319);
or U20132 (N_20132,N_17576,N_15832);
nand U20133 (N_20133,N_16446,N_18537);
and U20134 (N_20134,N_15384,N_15876);
and U20135 (N_20135,N_19967,N_17084);
nor U20136 (N_20136,N_19081,N_17806);
nor U20137 (N_20137,N_18699,N_18875);
and U20138 (N_20138,N_15293,N_19298);
nand U20139 (N_20139,N_17599,N_19689);
and U20140 (N_20140,N_17956,N_16379);
or U20141 (N_20141,N_16193,N_18275);
nor U20142 (N_20142,N_19853,N_17476);
or U20143 (N_20143,N_19696,N_16996);
nand U20144 (N_20144,N_16584,N_17868);
or U20145 (N_20145,N_17371,N_18610);
nor U20146 (N_20146,N_15517,N_17179);
or U20147 (N_20147,N_15074,N_16909);
and U20148 (N_20148,N_15829,N_17636);
nand U20149 (N_20149,N_17606,N_18394);
nand U20150 (N_20150,N_17249,N_17341);
nor U20151 (N_20151,N_15455,N_16203);
nor U20152 (N_20152,N_18727,N_19276);
nand U20153 (N_20153,N_19970,N_19573);
nand U20154 (N_20154,N_16632,N_18784);
nor U20155 (N_20155,N_18674,N_18013);
nor U20156 (N_20156,N_18922,N_17094);
and U20157 (N_20157,N_17525,N_15114);
or U20158 (N_20158,N_17356,N_16634);
or U20159 (N_20159,N_17197,N_19367);
nor U20160 (N_20160,N_17464,N_18047);
nor U20161 (N_20161,N_17440,N_16849);
or U20162 (N_20162,N_19876,N_19830);
and U20163 (N_20163,N_19170,N_17235);
and U20164 (N_20164,N_19508,N_15334);
nor U20165 (N_20165,N_16497,N_15061);
and U20166 (N_20166,N_18544,N_17603);
or U20167 (N_20167,N_19381,N_15001);
nor U20168 (N_20168,N_16861,N_16967);
and U20169 (N_20169,N_15055,N_19701);
and U20170 (N_20170,N_15659,N_15248);
or U20171 (N_20171,N_18261,N_15012);
nor U20172 (N_20172,N_19858,N_16945);
nand U20173 (N_20173,N_18511,N_16390);
and U20174 (N_20174,N_16455,N_19002);
nor U20175 (N_20175,N_19810,N_15864);
or U20176 (N_20176,N_16550,N_19079);
nand U20177 (N_20177,N_19195,N_19021);
and U20178 (N_20178,N_18790,N_18197);
and U20179 (N_20179,N_16195,N_15528);
and U20180 (N_20180,N_16917,N_17129);
xnor U20181 (N_20181,N_16136,N_19224);
nor U20182 (N_20182,N_15974,N_16930);
nor U20183 (N_20183,N_19554,N_18744);
nand U20184 (N_20184,N_16276,N_16884);
nand U20185 (N_20185,N_17668,N_19654);
nand U20186 (N_20186,N_19974,N_17159);
or U20187 (N_20187,N_18796,N_18828);
and U20188 (N_20188,N_19069,N_19319);
nand U20189 (N_20189,N_16445,N_18624);
and U20190 (N_20190,N_19752,N_15564);
and U20191 (N_20191,N_15658,N_16932);
or U20192 (N_20192,N_19763,N_19913);
xnor U20193 (N_20193,N_15943,N_15065);
and U20194 (N_20194,N_18071,N_19697);
and U20195 (N_20195,N_15418,N_17357);
nor U20196 (N_20196,N_17975,N_17845);
or U20197 (N_20197,N_19044,N_18065);
nand U20198 (N_20198,N_19474,N_16109);
nor U20199 (N_20199,N_17588,N_19799);
or U20200 (N_20200,N_19468,N_17393);
xnor U20201 (N_20201,N_16586,N_19631);
and U20202 (N_20202,N_15506,N_19387);
and U20203 (N_20203,N_18246,N_18522);
nor U20204 (N_20204,N_19759,N_18164);
or U20205 (N_20205,N_19193,N_17727);
or U20206 (N_20206,N_17992,N_19535);
and U20207 (N_20207,N_19837,N_17279);
or U20208 (N_20208,N_19520,N_17398);
and U20209 (N_20209,N_18516,N_16828);
nand U20210 (N_20210,N_15747,N_18721);
nor U20211 (N_20211,N_16617,N_19174);
and U20212 (N_20212,N_19262,N_17987);
nor U20213 (N_20213,N_19346,N_15106);
or U20214 (N_20214,N_15914,N_18663);
nor U20215 (N_20215,N_16029,N_18532);
nor U20216 (N_20216,N_18098,N_16502);
or U20217 (N_20217,N_19402,N_15835);
and U20218 (N_20218,N_15220,N_17526);
nand U20219 (N_20219,N_16974,N_15649);
nand U20220 (N_20220,N_19265,N_15318);
and U20221 (N_20221,N_18060,N_17230);
nor U20222 (N_20222,N_19730,N_18510);
xnor U20223 (N_20223,N_16259,N_17494);
nand U20224 (N_20224,N_18116,N_15929);
nand U20225 (N_20225,N_19778,N_18948);
nor U20226 (N_20226,N_17029,N_16170);
and U20227 (N_20227,N_17999,N_16258);
nand U20228 (N_20228,N_16399,N_19328);
and U20229 (N_20229,N_19803,N_19976);
nor U20230 (N_20230,N_18854,N_19007);
and U20231 (N_20231,N_16432,N_17240);
and U20232 (N_20232,N_19962,N_16615);
nand U20233 (N_20233,N_17661,N_19798);
xor U20234 (N_20234,N_17678,N_15321);
nand U20235 (N_20235,N_17615,N_18895);
nor U20236 (N_20236,N_18000,N_15996);
nand U20237 (N_20237,N_18440,N_15395);
and U20238 (N_20238,N_16757,N_15838);
or U20239 (N_20239,N_19511,N_16024);
or U20240 (N_20240,N_15295,N_19506);
nor U20241 (N_20241,N_18883,N_15465);
xnor U20242 (N_20242,N_15075,N_16776);
nor U20243 (N_20243,N_18957,N_18823);
nor U20244 (N_20244,N_17188,N_17981);
nand U20245 (N_20245,N_18782,N_17055);
or U20246 (N_20246,N_16746,N_15403);
or U20247 (N_20247,N_15514,N_16278);
nand U20248 (N_20248,N_18153,N_18775);
and U20249 (N_20249,N_15803,N_17384);
and U20250 (N_20250,N_15474,N_17148);
nor U20251 (N_20251,N_15085,N_16891);
and U20252 (N_20252,N_19222,N_19815);
nor U20253 (N_20253,N_18417,N_19294);
and U20254 (N_20254,N_18114,N_15241);
nand U20255 (N_20255,N_18434,N_17189);
and U20256 (N_20256,N_17772,N_15282);
and U20257 (N_20257,N_16743,N_15168);
or U20258 (N_20258,N_19116,N_16799);
or U20259 (N_20259,N_16836,N_17718);
nand U20260 (N_20260,N_18342,N_16534);
or U20261 (N_20261,N_17713,N_15496);
or U20262 (N_20262,N_19140,N_19313);
nor U20263 (N_20263,N_15717,N_18262);
or U20264 (N_20264,N_17009,N_19042);
nand U20265 (N_20265,N_19475,N_19770);
nor U20266 (N_20266,N_15546,N_17182);
nand U20267 (N_20267,N_16825,N_16385);
nand U20268 (N_20268,N_19398,N_18584);
and U20269 (N_20269,N_16200,N_18955);
or U20270 (N_20270,N_17812,N_16609);
or U20271 (N_20271,N_18475,N_19234);
and U20272 (N_20272,N_15771,N_19536);
or U20273 (N_20273,N_17323,N_15245);
and U20274 (N_20274,N_15743,N_19325);
and U20275 (N_20275,N_18175,N_16053);
or U20276 (N_20276,N_15607,N_17829);
nand U20277 (N_20277,N_18436,N_16521);
or U20278 (N_20278,N_16794,N_19529);
and U20279 (N_20279,N_15371,N_15000);
or U20280 (N_20280,N_16784,N_19683);
nand U20281 (N_20281,N_16566,N_15346);
nand U20282 (N_20282,N_19143,N_19039);
xnor U20283 (N_20283,N_16321,N_17155);
and U20284 (N_20284,N_18459,N_19995);
or U20285 (N_20285,N_16249,N_19301);
nand U20286 (N_20286,N_19240,N_15298);
nand U20287 (N_20287,N_18818,N_18631);
xor U20288 (N_20288,N_18628,N_15529);
or U20289 (N_20289,N_17491,N_17831);
xnor U20290 (N_20290,N_15023,N_19210);
nor U20291 (N_20291,N_18590,N_18497);
nor U20292 (N_20292,N_19626,N_16084);
and U20293 (N_20293,N_17733,N_16984);
xnor U20294 (N_20294,N_15152,N_17205);
nand U20295 (N_20295,N_18827,N_17995);
nand U20296 (N_20296,N_16202,N_18264);
nand U20297 (N_20297,N_17656,N_18268);
and U20298 (N_20298,N_19370,N_16947);
nand U20299 (N_20299,N_17305,N_19945);
or U20300 (N_20300,N_17000,N_17378);
or U20301 (N_20301,N_17994,N_18337);
or U20302 (N_20302,N_19659,N_15249);
or U20303 (N_20303,N_17460,N_17586);
and U20304 (N_20304,N_15158,N_15170);
nand U20305 (N_20305,N_19183,N_19273);
nor U20306 (N_20306,N_16520,N_16325);
nand U20307 (N_20307,N_17888,N_17287);
or U20308 (N_20308,N_17939,N_16630);
nor U20309 (N_20309,N_16208,N_17196);
nand U20310 (N_20310,N_19336,N_15811);
or U20311 (N_20311,N_16192,N_16604);
nand U20312 (N_20312,N_18503,N_17359);
nor U20313 (N_20313,N_19338,N_18259);
nor U20314 (N_20314,N_15397,N_18249);
xor U20315 (N_20315,N_16019,N_18964);
and U20316 (N_20316,N_16579,N_17534);
or U20317 (N_20317,N_19544,N_15083);
nor U20318 (N_20318,N_16642,N_15338);
and U20319 (N_20319,N_16725,N_17658);
nor U20320 (N_20320,N_18398,N_18927);
or U20321 (N_20321,N_17783,N_18151);
or U20322 (N_20322,N_15808,N_18633);
nor U20323 (N_20323,N_17451,N_17318);
nand U20324 (N_20324,N_19568,N_19327);
or U20325 (N_20325,N_15831,N_18473);
or U20326 (N_20326,N_17894,N_15316);
nor U20327 (N_20327,N_18531,N_17497);
and U20328 (N_20328,N_16644,N_18075);
nor U20329 (N_20329,N_15466,N_15415);
nor U20330 (N_20330,N_15368,N_16886);
or U20331 (N_20331,N_19726,N_16826);
nor U20332 (N_20332,N_18869,N_16535);
nand U20333 (N_20333,N_19532,N_16857);
or U20334 (N_20334,N_17955,N_15725);
and U20335 (N_20335,N_18974,N_15369);
and U20336 (N_20336,N_15167,N_16572);
or U20337 (N_20337,N_16716,N_17983);
nor U20338 (N_20338,N_18600,N_17489);
or U20339 (N_20339,N_18088,N_19545);
nor U20340 (N_20340,N_18535,N_16532);
and U20341 (N_20341,N_16294,N_17801);
and U20342 (N_20342,N_18657,N_18365);
nand U20343 (N_20343,N_15956,N_15558);
nor U20344 (N_20344,N_19560,N_16303);
nand U20345 (N_20345,N_19997,N_18599);
and U20346 (N_20346,N_16991,N_17262);
nor U20347 (N_20347,N_15605,N_16242);
nand U20348 (N_20348,N_19912,N_15825);
nand U20349 (N_20349,N_18224,N_16134);
and U20350 (N_20350,N_17998,N_15924);
nand U20351 (N_20351,N_19032,N_16966);
nor U20352 (N_20352,N_18193,N_19067);
nand U20353 (N_20353,N_16260,N_15794);
nor U20354 (N_20354,N_16554,N_19119);
and U20355 (N_20355,N_18080,N_18753);
nor U20356 (N_20356,N_18217,N_15288);
and U20357 (N_20357,N_17177,N_15254);
xnor U20358 (N_20358,N_18671,N_18484);
nand U20359 (N_20359,N_17152,N_15157);
and U20360 (N_20360,N_19366,N_17237);
xnor U20361 (N_20361,N_19580,N_17640);
and U20362 (N_20362,N_17502,N_19085);
nor U20363 (N_20363,N_15587,N_15327);
and U20364 (N_20364,N_19509,N_18195);
nand U20365 (N_20365,N_19038,N_18947);
nand U20366 (N_20366,N_17610,N_19317);
or U20367 (N_20367,N_15150,N_19879);
or U20368 (N_20368,N_17157,N_19820);
nand U20369 (N_20369,N_15177,N_18654);
nand U20370 (N_20370,N_17954,N_18551);
nor U20371 (N_20371,N_18768,N_18185);
nor U20372 (N_20372,N_17915,N_17570);
nor U20373 (N_20373,N_15501,N_18402);
nand U20374 (N_20374,N_17834,N_16558);
or U20375 (N_20375,N_17539,N_16684);
or U20376 (N_20376,N_19709,N_16451);
nand U20377 (N_20377,N_18911,N_19331);
nand U20378 (N_20378,N_18144,N_17083);
or U20379 (N_20379,N_18432,N_15774);
or U20380 (N_20380,N_19917,N_16431);
nand U20381 (N_20381,N_18081,N_17677);
nand U20382 (N_20382,N_16553,N_19386);
nand U20383 (N_20383,N_18465,N_18730);
or U20384 (N_20384,N_17273,N_17274);
and U20385 (N_20385,N_17962,N_17721);
nand U20386 (N_20386,N_17798,N_18466);
or U20387 (N_20387,N_15748,N_16500);
xnor U20388 (N_20388,N_16544,N_17551);
xor U20389 (N_20389,N_19284,N_16097);
nand U20390 (N_20390,N_16677,N_15570);
or U20391 (N_20391,N_17932,N_18552);
or U20392 (N_20392,N_15209,N_17232);
and U20393 (N_20393,N_19094,N_17380);
or U20394 (N_20394,N_16829,N_19939);
nand U20395 (N_20395,N_16788,N_19406);
nor U20396 (N_20396,N_18426,N_15189);
nand U20397 (N_20397,N_16704,N_17930);
and U20398 (N_20398,N_16075,N_19419);
nand U20399 (N_20399,N_15745,N_17597);
nor U20400 (N_20400,N_15709,N_19695);
or U20401 (N_20401,N_17141,N_17804);
xnor U20402 (N_20402,N_16792,N_17163);
and U20403 (N_20403,N_16739,N_17216);
xnor U20404 (N_20404,N_18999,N_19883);
nor U20405 (N_20405,N_16406,N_19975);
and U20406 (N_20406,N_15842,N_18526);
nand U20407 (N_20407,N_18919,N_15406);
nand U20408 (N_20408,N_17527,N_18542);
nor U20409 (N_20409,N_19115,N_17174);
or U20410 (N_20410,N_17299,N_16806);
nor U20411 (N_20411,N_18612,N_17920);
nor U20412 (N_20412,N_18991,N_19599);
and U20413 (N_20413,N_16672,N_18120);
or U20414 (N_20414,N_16377,N_16622);
or U20415 (N_20415,N_19286,N_15279);
or U20416 (N_20416,N_19244,N_15979);
nand U20417 (N_20417,N_19458,N_15058);
nor U20418 (N_20418,N_15915,N_17266);
and U20419 (N_20419,N_16943,N_15934);
and U20420 (N_20420,N_19050,N_16707);
nor U20421 (N_20421,N_15989,N_16878);
and U20422 (N_20422,N_17449,N_19379);
nand U20423 (N_20423,N_18393,N_19235);
nor U20424 (N_20424,N_19750,N_18139);
or U20425 (N_20425,N_15022,N_19438);
or U20426 (N_20426,N_18296,N_15103);
and U20427 (N_20427,N_15547,N_16994);
or U20428 (N_20428,N_15440,N_15651);
nor U20429 (N_20429,N_18773,N_15999);
or U20430 (N_20430,N_15376,N_15827);
nor U20431 (N_20431,N_18335,N_15941);
nor U20432 (N_20432,N_16590,N_17420);
and U20433 (N_20433,N_16296,N_16955);
xnor U20434 (N_20434,N_19431,N_16651);
and U20435 (N_20435,N_19624,N_16629);
nand U20436 (N_20436,N_19875,N_16777);
and U20437 (N_20437,N_19469,N_19063);
and U20438 (N_20438,N_15086,N_17479);
or U20439 (N_20439,N_17771,N_19897);
xor U20440 (N_20440,N_19805,N_18996);
xnor U20441 (N_20441,N_16848,N_18178);
and U20442 (N_20442,N_16256,N_18936);
xor U20443 (N_20443,N_15661,N_15664);
or U20444 (N_20444,N_17794,N_17978);
xnor U20445 (N_20445,N_19546,N_16606);
or U20446 (N_20446,N_15856,N_17857);
nand U20447 (N_20447,N_17112,N_15611);
nor U20448 (N_20448,N_19653,N_16220);
nor U20449 (N_20449,N_19772,N_18377);
nor U20450 (N_20450,N_15102,N_19771);
or U20451 (N_20451,N_15612,N_16280);
or U20452 (N_20452,N_19722,N_15120);
and U20453 (N_20453,N_19321,N_15309);
and U20454 (N_20454,N_19444,N_19227);
or U20455 (N_20455,N_18183,N_17556);
nand U20456 (N_20456,N_18306,N_18562);
or U20457 (N_20457,N_19358,N_15809);
or U20458 (N_20458,N_19049,N_16665);
and U20459 (N_20459,N_18634,N_17792);
or U20460 (N_20460,N_16834,N_18585);
xor U20461 (N_20461,N_15166,N_15525);
nand U20462 (N_20462,N_17406,N_15215);
nor U20463 (N_20463,N_16439,N_17859);
nand U20464 (N_20464,N_15954,N_19783);
and U20465 (N_20465,N_16018,N_18791);
nand U20466 (N_20466,N_16981,N_19688);
nor U20467 (N_20467,N_16954,N_16540);
and U20468 (N_20468,N_18764,N_16187);
and U20469 (N_20469,N_19517,N_18437);
or U20470 (N_20470,N_15349,N_19220);
nor U20471 (N_20471,N_16421,N_16453);
nor U20472 (N_20472,N_18980,N_17679);
and U20473 (N_20473,N_16008,N_16837);
nor U20474 (N_20474,N_16907,N_16745);
xor U20475 (N_20475,N_18210,N_16108);
nand U20476 (N_20476,N_15003,N_16982);
nor U20477 (N_20477,N_16659,N_19575);
nor U20478 (N_20478,N_17558,N_18822);
or U20479 (N_20479,N_15814,N_19375);
nor U20480 (N_20480,N_19315,N_16042);
and U20481 (N_20481,N_18346,N_15682);
and U20482 (N_20482,N_19348,N_15396);
nand U20483 (N_20483,N_16887,N_16318);
and U20484 (N_20484,N_18486,N_15151);
or U20485 (N_20485,N_16894,N_17331);
nand U20486 (N_20486,N_15433,N_18982);
or U20487 (N_20487,N_18975,N_17294);
or U20488 (N_20488,N_15961,N_16735);
or U20489 (N_20489,N_17728,N_19863);
xnor U20490 (N_20490,N_19541,N_16027);
nand U20491 (N_20491,N_18920,N_15131);
and U20492 (N_20492,N_17173,N_19919);
nor U20493 (N_20493,N_19718,N_15310);
nor U20494 (N_20494,N_18576,N_15208);
or U20495 (N_20495,N_19944,N_15983);
or U20496 (N_20496,N_16620,N_17788);
and U20497 (N_20497,N_19217,N_19725);
nor U20498 (N_20498,N_18190,N_17893);
nor U20499 (N_20499,N_19168,N_16819);
and U20500 (N_20500,N_17311,N_16218);
or U20501 (N_20501,N_18740,N_16360);
nor U20502 (N_20502,N_16413,N_17405);
nor U20503 (N_20503,N_15853,N_16885);
xor U20504 (N_20504,N_17883,N_17791);
and U20505 (N_20505,N_17040,N_15533);
xor U20506 (N_20506,N_19720,N_15343);
nor U20507 (N_20507,N_18227,N_17079);
nor U20508 (N_20508,N_16787,N_16073);
nand U20509 (N_20509,N_16457,N_19835);
and U20510 (N_20510,N_16667,N_16480);
nor U20511 (N_20511,N_15038,N_16244);
or U20512 (N_20512,N_15951,N_17589);
or U20513 (N_20513,N_19250,N_19848);
and U20514 (N_20514,N_17993,N_17361);
nand U20515 (N_20515,N_17151,N_15320);
and U20516 (N_20516,N_19194,N_15312);
or U20517 (N_20517,N_16526,N_17587);
nor U20518 (N_20518,N_19547,N_16026);
nand U20519 (N_20519,N_18416,N_17210);
or U20520 (N_20520,N_15758,N_17630);
and U20521 (N_20521,N_18811,N_16401);
or U20522 (N_20522,N_16323,N_19542);
or U20523 (N_20523,N_17169,N_18078);
xor U20524 (N_20524,N_15472,N_15358);
and U20525 (N_20525,N_15483,N_18460);
nand U20526 (N_20526,N_16418,N_19112);
and U20527 (N_20527,N_18844,N_17918);
nor U20528 (N_20528,N_15750,N_18735);
nand U20529 (N_20529,N_17469,N_15692);
and U20530 (N_20530,N_15205,N_15485);
xnor U20531 (N_20531,N_15425,N_16899);
or U20532 (N_20532,N_19491,N_19364);
nor U20533 (N_20533,N_17963,N_18378);
or U20534 (N_20534,N_15156,N_18166);
xnor U20535 (N_20535,N_17714,N_15302);
nor U20536 (N_20536,N_17014,N_16513);
nand U20537 (N_20537,N_15590,N_15264);
and U20538 (N_20538,N_15975,N_19644);
nor U20539 (N_20539,N_19617,N_16124);
nand U20540 (N_20540,N_16802,N_19157);
nand U20541 (N_20541,N_18352,N_17213);
nor U20542 (N_20542,N_16876,N_16175);
nand U20543 (N_20543,N_16839,N_19645);
nor U20544 (N_20544,N_15495,N_18457);
and U20545 (N_20545,N_15393,N_15804);
or U20546 (N_20546,N_15147,N_19742);
or U20547 (N_20547,N_15683,N_19389);
or U20548 (N_20548,N_19952,N_17376);
and U20549 (N_20549,N_19272,N_18617);
or U20550 (N_20550,N_17631,N_16015);
nand U20551 (N_20551,N_17832,N_19966);
and U20552 (N_20552,N_15959,N_17542);
nor U20553 (N_20553,N_18469,N_19237);
nand U20554 (N_20554,N_18137,N_16101);
or U20555 (N_20555,N_18238,N_16602);
nor U20556 (N_20556,N_15134,N_15033);
nor U20557 (N_20557,N_17144,N_16065);
nor U20558 (N_20558,N_19337,N_15772);
nor U20559 (N_20559,N_16896,N_17689);
xor U20560 (N_20560,N_19515,N_19957);
or U20561 (N_20561,N_18145,N_19550);
nand U20562 (N_20562,N_15603,N_18222);
or U20563 (N_20563,N_16559,N_17929);
nor U20564 (N_20564,N_18468,N_19590);
nand U20565 (N_20565,N_18165,N_18789);
and U20566 (N_20566,N_19663,N_16492);
nand U20567 (N_20567,N_18133,N_18257);
nor U20568 (N_20568,N_17195,N_17997);
nand U20569 (N_20569,N_18592,N_18739);
or U20570 (N_20570,N_15967,N_19627);
nand U20571 (N_20571,N_17100,N_18129);
nor U20572 (N_20572,N_16494,N_19886);
nand U20573 (N_20573,N_19184,N_17923);
or U20574 (N_20574,N_19581,N_18063);
and U20575 (N_20575,N_16189,N_16944);
nand U20576 (N_20576,N_17719,N_16438);
nor U20577 (N_20577,N_16168,N_16612);
and U20578 (N_20578,N_16804,N_18738);
or U20579 (N_20579,N_15819,N_19190);
or U20580 (N_20580,N_16402,N_15389);
nor U20581 (N_20581,N_15104,N_17785);
or U20582 (N_20582,N_17203,N_17329);
nor U20583 (N_20583,N_19890,N_19451);
or U20584 (N_20584,N_15042,N_17941);
or U20585 (N_20585,N_16726,N_18281);
nor U20586 (N_20586,N_15238,N_16153);
and U20587 (N_20587,N_16942,N_15481);
nor U20588 (N_20588,N_19588,N_16113);
or U20589 (N_20589,N_17712,N_19233);
xnor U20590 (N_20590,N_17022,N_17343);
or U20591 (N_20591,N_17028,N_16624);
nor U20592 (N_20592,N_17207,N_15713);
nand U20593 (N_20593,N_16302,N_18597);
nand U20594 (N_20594,N_15263,N_19466);
xnor U20595 (N_20595,N_17573,N_19949);
nand U20596 (N_20596,N_17777,N_18318);
and U20597 (N_20597,N_19443,N_16772);
and U20598 (N_20598,N_19968,N_15286);
or U20599 (N_20599,N_16288,N_15315);
nor U20600 (N_20600,N_17463,N_16874);
xnor U20601 (N_20601,N_16037,N_15734);
or U20602 (N_20602,N_15600,N_16173);
or U20603 (N_20603,N_19254,N_15015);
and U20604 (N_20604,N_19378,N_15183);
xor U20605 (N_20605,N_16481,N_16950);
xnor U20606 (N_20606,N_19861,N_19323);
nand U20607 (N_20607,N_17908,N_18169);
nand U20608 (N_20608,N_16901,N_15613);
xnor U20609 (N_20609,N_17764,N_16400);
or U20610 (N_20610,N_15828,N_15730);
nor U20611 (N_20611,N_18058,N_16129);
and U20612 (N_20612,N_18181,N_16238);
or U20613 (N_20613,N_17787,N_19182);
or U20614 (N_20614,N_15988,N_19608);
or U20615 (N_20615,N_17548,N_19776);
nand U20616 (N_20616,N_19015,N_15867);
nor U20617 (N_20617,N_15894,N_17700);
or U20618 (N_20618,N_19489,N_16210);
xnor U20619 (N_20619,N_15431,N_19373);
and U20620 (N_20620,N_19339,N_16769);
or U20621 (N_20621,N_19685,N_15887);
and U20622 (N_20622,N_18900,N_18285);
nand U20623 (N_20623,N_15866,N_15490);
nand U20624 (N_20624,N_19922,N_15428);
and U20625 (N_20625,N_19232,N_18767);
nor U20626 (N_20626,N_19180,N_15193);
or U20627 (N_20627,N_19300,N_19228);
and U20628 (N_20628,N_19487,N_15283);
and U20629 (N_20629,N_19258,N_16014);
and U20630 (N_20630,N_15822,N_16374);
or U20631 (N_20631,N_15456,N_16013);
and U20632 (N_20632,N_16697,N_17498);
and U20633 (N_20633,N_18171,N_16753);
and U20634 (N_20634,N_15970,N_15900);
nand U20635 (N_20635,N_19694,N_19022);
nor U20636 (N_20636,N_18177,N_16902);
nor U20637 (N_20637,N_16577,N_18862);
or U20638 (N_20638,N_19822,N_17372);
or U20639 (N_20639,N_17281,N_15359);
nor U20640 (N_20640,N_15551,N_18639);
or U20641 (N_20641,N_18885,N_18490);
or U20642 (N_20642,N_15752,N_16567);
nor U20643 (N_20643,N_18965,N_17503);
nand U20644 (N_20644,N_17818,N_19563);
or U20645 (N_20645,N_16686,N_17089);
nor U20646 (N_20646,N_19500,N_18390);
nand U20647 (N_20647,N_17253,N_15852);
and U20648 (N_20648,N_15257,N_18411);
nand U20649 (N_20649,N_16872,N_18043);
xnor U20650 (N_20650,N_19000,N_16715);
nand U20651 (N_20651,N_16219,N_17291);
nor U20652 (N_20652,N_16443,N_17126);
nor U20653 (N_20653,N_18596,N_19020);
nor U20654 (N_20654,N_19450,N_17856);
nor U20655 (N_20655,N_17957,N_19176);
nor U20656 (N_20656,N_18877,N_17006);
and U20657 (N_20657,N_16529,N_19318);
or U20658 (N_20658,N_15066,N_16796);
nor U20659 (N_20659,N_18121,N_15785);
or U20660 (N_20660,N_15430,N_16618);
nor U20661 (N_20661,N_18867,N_17851);
and U20662 (N_20662,N_17648,N_15379);
and U20663 (N_20663,N_18345,N_15164);
and U20664 (N_20664,N_18229,N_19047);
and U20665 (N_20665,N_15162,N_19757);
nor U20666 (N_20666,N_18189,N_19972);
or U20667 (N_20667,N_17158,N_19817);
nand U20668 (N_20668,N_19440,N_16539);
or U20669 (N_20669,N_17945,N_17482);
nand U20670 (N_20670,N_17363,N_19187);
nor U20671 (N_20671,N_19993,N_19555);
nand U20672 (N_20672,N_18880,N_15515);
nor U20673 (N_20673,N_18741,N_17951);
nor U20674 (N_20674,N_16199,N_18501);
nor U20675 (N_20675,N_15861,N_17773);
or U20676 (N_20676,N_19775,N_17454);
and U20677 (N_20677,N_15741,N_17964);
or U20678 (N_20678,N_16386,N_18508);
or U20679 (N_20679,N_16939,N_18429);
or U20680 (N_20680,N_18204,N_15196);
or U20681 (N_20681,N_17795,N_18626);
and U20682 (N_20682,N_18772,N_16209);
nand U20683 (N_20683,N_18889,N_18757);
nor U20684 (N_20684,N_18408,N_16074);
nor U20685 (N_20685,N_18170,N_15191);
xor U20686 (N_20686,N_16952,N_15693);
or U20687 (N_20687,N_17227,N_16813);
nor U20688 (N_20688,N_19936,N_19743);
and U20689 (N_20689,N_18799,N_15165);
xnor U20690 (N_20690,N_19700,N_19149);
nor U20691 (N_20691,N_19296,N_19519);
or U20692 (N_20692,N_18615,N_17321);
nor U20693 (N_20693,N_17447,N_18424);
xor U20694 (N_20694,N_17461,N_18015);
nand U20695 (N_20695,N_16758,N_17481);
or U20696 (N_20696,N_18215,N_16958);
and U20697 (N_20697,N_16355,N_16407);
and U20698 (N_20698,N_17034,N_15497);
nor U20699 (N_20699,N_19470,N_19229);
or U20700 (N_20700,N_16911,N_19017);
nand U20701 (N_20701,N_17808,N_19887);
and U20702 (N_20702,N_18710,N_19707);
and U20703 (N_20703,N_18418,N_16919);
nand U20704 (N_20704,N_17980,N_16030);
nor U20705 (N_20705,N_16409,N_18125);
nor U20706 (N_20706,N_16951,N_18668);
and U20707 (N_20707,N_17819,N_15443);
nor U20708 (N_20708,N_19559,N_19479);
and U20709 (N_20709,N_19353,N_18766);
nand U20710 (N_20710,N_18491,N_16292);
or U20711 (N_20711,N_16889,N_17023);
nor U20712 (N_20712,N_19903,N_15782);
or U20713 (N_20713,N_18560,N_16660);
and U20714 (N_20714,N_19311,N_16125);
nor U20715 (N_20715,N_16369,N_16456);
or U20716 (N_20716,N_15331,N_18149);
nand U20717 (N_20717,N_16201,N_19120);
and U20718 (N_20718,N_15964,N_18527);
and U20719 (N_20719,N_16733,N_17403);
nand U20720 (N_20720,N_16685,N_17068);
nor U20721 (N_20721,N_19514,N_15841);
or U20722 (N_20722,N_19611,N_19065);
xnor U20723 (N_20723,N_15760,N_17214);
or U20724 (N_20724,N_15672,N_16877);
and U20725 (N_20725,N_16935,N_17635);
or U20726 (N_20726,N_16138,N_17968);
and U20727 (N_20727,N_17039,N_16762);
nand U20728 (N_20728,N_16248,N_16724);
xor U20729 (N_20729,N_19572,N_15932);
or U20730 (N_20730,N_15289,N_18554);
nor U20731 (N_20731,N_15966,N_17850);
nand U20732 (N_20732,N_18478,N_15751);
nor U20733 (N_20733,N_17775,N_17886);
and U20734 (N_20734,N_15020,N_18430);
xnor U20735 (N_20735,N_16150,N_17690);
nand U20736 (N_20736,N_18493,N_15246);
and U20737 (N_20737,N_17643,N_15329);
nor U20738 (N_20738,N_15036,N_15947);
and U20739 (N_20739,N_19134,N_19553);
nor U20740 (N_20740,N_19011,N_15635);
nor U20741 (N_20741,N_18915,N_19831);
nor U20742 (N_20742,N_16204,N_17093);
nor U20743 (N_20743,N_15927,N_17560);
and U20744 (N_20744,N_18888,N_18062);
or U20745 (N_20745,N_18447,N_19128);
or U20746 (N_20746,N_19090,N_18685);
or U20747 (N_20747,N_15685,N_16820);
nand U20748 (N_20748,N_16236,N_18022);
nand U20749 (N_20749,N_17477,N_19906);
xnor U20750 (N_20750,N_17991,N_19283);
xnor U20751 (N_20751,N_17916,N_17082);
xor U20752 (N_20752,N_15792,N_19436);
nand U20753 (N_20753,N_19978,N_18037);
and U20754 (N_20754,N_17762,N_17005);
xor U20755 (N_20755,N_18167,N_17519);
or U20756 (N_20756,N_15487,N_15586);
nor U20757 (N_20757,N_19564,N_19152);
or U20758 (N_20758,N_18632,N_16458);
nor U20759 (N_20759,N_17942,N_18461);
nand U20760 (N_20760,N_18669,N_16106);
nor U20761 (N_20761,N_17699,N_18629);
nand U20762 (N_20762,N_17766,N_19839);
and U20763 (N_20763,N_16808,N_18454);
nor U20764 (N_20764,N_16890,N_18547);
and U20765 (N_20765,N_16688,N_17505);
xor U20766 (N_20766,N_16479,N_16281);
and U20767 (N_20767,N_15079,N_18549);
and U20768 (N_20768,N_18388,N_17649);
nand U20769 (N_20769,N_18371,N_17425);
and U20770 (N_20770,N_15688,N_19230);
nor U20771 (N_20771,N_16510,N_18946);
nand U20772 (N_20772,N_16811,N_18301);
or U20773 (N_20773,N_16345,N_15614);
and U20774 (N_20774,N_19601,N_18085);
or U20775 (N_20775,N_15344,N_18938);
nand U20776 (N_20776,N_18284,N_15424);
nor U20777 (N_20777,N_19684,N_16830);
nand U20778 (N_20778,N_17838,N_15960);
nand U20779 (N_20779,N_17193,N_17971);
nor U20780 (N_20780,N_15364,N_18731);
and U20781 (N_20781,N_15781,N_18715);
xnor U20782 (N_20782,N_17751,N_17156);
nor U20783 (N_20783,N_15034,N_15606);
xor U20784 (N_20784,N_18326,N_17815);
or U20785 (N_20785,N_15646,N_18242);
xnor U20786 (N_20786,N_16061,N_18921);
or U20787 (N_20787,N_15689,N_17435);
or U20788 (N_20788,N_16301,N_17619);
nor U20789 (N_20789,N_17248,N_17127);
and U20790 (N_20790,N_19855,N_18950);
nor U20791 (N_20791,N_19135,N_19257);
or U20792 (N_20792,N_19188,N_16897);
and U20793 (N_20793,N_16595,N_17295);
nand U20794 (N_20794,N_18489,N_15647);
or U20795 (N_20795,N_16600,N_18713);
nand U20796 (N_20796,N_16993,N_16228);
and U20797 (N_20797,N_16484,N_18095);
and U20798 (N_20798,N_16980,N_16927);
and U20799 (N_20799,N_15197,N_15905);
or U20800 (N_20800,N_17741,N_18976);
and U20801 (N_20801,N_19087,N_17685);
xnor U20802 (N_20802,N_16827,N_16334);
and U20803 (N_20803,N_17496,N_17095);
and U20804 (N_20804,N_18941,N_19882);
and U20805 (N_20805,N_17853,N_19452);
nand U20806 (N_20806,N_18676,N_15094);
and U20807 (N_20807,N_18800,N_19478);
and U20808 (N_20808,N_18304,N_16936);
and U20809 (N_20809,N_15783,N_15718);
nand U20810 (N_20810,N_17485,N_16166);
or U20811 (N_20811,N_18819,N_15574);
xnor U20812 (N_20812,N_19503,N_18104);
nor U20813 (N_20813,N_17912,N_18007);
nand U20814 (N_20814,N_18758,N_18648);
xor U20815 (N_20815,N_18487,N_19673);
nor U20816 (N_20816,N_19447,N_15126);
or U20817 (N_20817,N_19415,N_18385);
xnor U20818 (N_20818,N_16298,N_15210);
nand U20819 (N_20819,N_18972,N_16556);
nor U20820 (N_20820,N_15270,N_18272);
nand U20821 (N_20821,N_17826,N_18861);
nand U20822 (N_20822,N_15493,N_18859);
nand U20823 (N_20823,N_17045,N_16021);
nand U20824 (N_20824,N_16317,N_19984);
or U20825 (N_20825,N_16410,N_19100);
nand U20826 (N_20826,N_15447,N_18978);
and U20827 (N_20827,N_15325,N_17784);
and U20828 (N_20828,N_19058,N_19711);
or U20829 (N_20829,N_19592,N_18076);
and U20830 (N_20830,N_16290,N_17302);
and U20831 (N_20831,N_16368,N_18423);
nand U20832 (N_20832,N_16322,N_17187);
nor U20833 (N_20833,N_16313,N_19430);
and U20834 (N_20834,N_15227,N_19484);
nand U20835 (N_20835,N_18808,N_18512);
and U20836 (N_20836,N_19354,N_18198);
nand U20837 (N_20837,N_15721,N_17878);
and U20838 (N_20838,N_15512,N_18857);
xor U20839 (N_20839,N_18971,N_15370);
nor U20840 (N_20840,N_16167,N_19915);
and U20841 (N_20841,N_19155,N_18441);
nor U20842 (N_20842,N_19660,N_18756);
nand U20843 (N_20843,N_16358,N_17550);
nor U20844 (N_20844,N_15460,N_15797);
or U20845 (N_20845,N_17805,N_18192);
and U20846 (N_20846,N_18323,N_17003);
nand U20847 (N_20847,N_18036,N_16469);
or U20848 (N_20848,N_17774,N_19941);
and U20849 (N_20849,N_15715,N_19303);
nor U20850 (N_20850,N_19723,N_16734);
and U20851 (N_20851,N_15139,N_17664);
nand U20852 (N_20852,N_16477,N_18664);
nand U20853 (N_20853,N_16270,N_18298);
xor U20854 (N_20854,N_16929,N_17109);
nand U20855 (N_20855,N_15176,N_15885);
and U20856 (N_20856,N_17882,N_16549);
and U20857 (N_20857,N_17257,N_17760);
or U20858 (N_20858,N_15977,N_17545);
or U20859 (N_20859,N_18557,N_19421);
nand U20860 (N_20860,N_18876,N_18297);
and U20861 (N_20861,N_15076,N_16499);
or U20862 (N_20862,N_16528,N_15073);
nor U20863 (N_20863,N_18004,N_18330);
nand U20864 (N_20864,N_18391,N_18293);
nor U20865 (N_20865,N_15695,N_19538);
nor U20866 (N_20866,N_16361,N_15592);
nor U20867 (N_20867,N_18136,N_19907);
and U20868 (N_20868,N_17535,N_15155);
nand U20869 (N_20869,N_16767,N_17800);
nor U20870 (N_20870,N_19390,N_19821);
nor U20871 (N_20871,N_19892,N_18963);
nand U20872 (N_20872,N_17506,N_15221);
nor U20873 (N_20873,N_16670,N_19635);
or U20874 (N_20874,N_19647,N_15354);
or U20875 (N_20875,N_19840,N_16742);
nand U20876 (N_20876,N_15776,N_19860);
nor U20877 (N_20877,N_17746,N_16164);
nor U20878 (N_20878,N_15834,N_15458);
and U20879 (N_20879,N_15630,N_16731);
nand U20880 (N_20880,N_18712,N_19279);
or U20881 (N_20881,N_17761,N_18369);
nor U20882 (N_20882,N_16375,N_15530);
nand U20883 (N_20883,N_16491,N_18884);
or U20884 (N_20884,N_16326,N_16895);
nor U20885 (N_20885,N_19990,N_18191);
or U20886 (N_20886,N_19350,N_17286);
or U20887 (N_20887,N_19613,N_15500);
nor U20888 (N_20888,N_18270,N_16017);
xor U20889 (N_20889,N_17110,N_16843);
or U20890 (N_20890,N_17473,N_17414);
or U20891 (N_20891,N_18235,N_19595);
nor U20892 (N_20892,N_18184,N_15287);
and U20893 (N_20893,N_19736,N_18570);
nand U20894 (N_20894,N_18207,N_17368);
and U20895 (N_20895,N_16730,N_15339);
xnor U20896 (N_20896,N_17652,N_19448);
nand U20897 (N_20897,N_17293,N_18679);
xor U20898 (N_20898,N_16650,N_18809);
nor U20899 (N_20899,N_15348,N_15985);
nor U20900 (N_20900,N_18606,N_18807);
nor U20901 (N_20901,N_15982,N_19963);
or U20902 (N_20902,N_17088,N_16295);
and U20903 (N_20903,N_19692,N_15419);
or U20904 (N_20904,N_18001,N_16311);
and U20905 (N_20905,N_16165,N_18728);
nand U20906 (N_20906,N_15652,N_17913);
nor U20907 (N_20907,N_16508,N_18951);
and U20908 (N_20908,N_18605,N_18096);
or U20909 (N_20909,N_18896,N_19524);
nor U20910 (N_20910,N_17442,N_19433);
or U20911 (N_20911,N_15919,N_19639);
or U20912 (N_20912,N_19946,N_18973);
nor U20913 (N_20913,N_17090,N_18736);
xor U20914 (N_20914,N_15198,N_18621);
nor U20915 (N_20915,N_15062,N_18820);
nand U20916 (N_20916,N_17967,N_15011);
nor U20917 (N_20917,N_18569,N_15888);
or U20918 (N_20918,N_16389,N_19392);
xor U20919 (N_20919,N_18384,N_18387);
nor U20920 (N_20920,N_17618,N_18494);
nand U20921 (N_20921,N_15780,N_15123);
xnor U20922 (N_20922,N_19148,N_16003);
xnor U20923 (N_20923,N_16127,N_19824);
nor U20924 (N_20924,N_17121,N_18240);
and U20925 (N_20925,N_15340,N_17979);
or U20926 (N_20926,N_16522,N_15252);
nor U20927 (N_20927,N_18134,N_15454);
nor U20928 (N_20928,N_17241,N_16394);
nor U20929 (N_20929,N_17574,N_15178);
nor U20930 (N_20930,N_16217,N_19578);
and U20931 (N_20931,N_18686,N_15297);
and U20932 (N_20932,N_16832,N_15006);
nor U20933 (N_20933,N_18206,N_16263);
and U20934 (N_20934,N_16706,N_15332);
xor U20935 (N_20935,N_16085,N_19299);
nand U20936 (N_20936,N_18420,N_19159);
or U20937 (N_20937,N_17410,N_17212);
and U20938 (N_20938,N_17705,N_17407);
nand U20939 (N_20939,N_19073,N_18031);
nand U20940 (N_20940,N_16773,N_18086);
or U20941 (N_20941,N_19202,N_17639);
and U20942 (N_20942,N_17590,N_16082);
nor U20943 (N_20943,N_19048,N_18325);
nand U20944 (N_20944,N_18188,N_17632);
nand U20945 (N_20945,N_18173,N_18327);
nand U20946 (N_20946,N_17400,N_19030);
or U20947 (N_20947,N_17483,N_19745);
or U20948 (N_20948,N_18020,N_19642);
or U20949 (N_20949,N_18607,N_15477);
or U20950 (N_20950,N_16470,N_19658);
or U20951 (N_20951,N_16475,N_18838);
nand U20952 (N_20952,N_18689,N_18930);
nand U20953 (N_20953,N_18021,N_19095);
xor U20954 (N_20954,N_19488,N_16233);
and U20955 (N_20955,N_15990,N_15753);
nand U20956 (N_20956,N_15489,N_19322);
xnor U20957 (N_20957,N_15939,N_18112);
nand U20958 (N_20958,N_18109,N_16490);
nor U20959 (N_20959,N_17259,N_16563);
nand U20960 (N_20960,N_15414,N_18793);
nor U20961 (N_20961,N_16147,N_19516);
nor U20962 (N_20962,N_15108,N_15958);
or U20963 (N_20963,N_16750,N_17814);
and U20964 (N_20964,N_17052,N_15524);
nor U20965 (N_20965,N_17388,N_19249);
or U20966 (N_20966,N_15097,N_17011);
nor U20967 (N_20967,N_15863,N_19305);
or U20968 (N_20968,N_19154,N_16673);
nor U20969 (N_20969,N_16449,N_16342);
and U20970 (N_20970,N_19746,N_18010);
nand U20971 (N_20971,N_16388,N_19983);
or U20972 (N_20972,N_18704,N_15138);
or U20973 (N_20973,N_19940,N_16120);
nor U20974 (N_20974,N_16524,N_19797);
or U20975 (N_20975,N_18030,N_15423);
nand U20976 (N_20976,N_18614,N_16336);
or U20977 (N_20977,N_17876,N_16454);
and U20978 (N_20978,N_15699,N_17906);
and U20979 (N_20979,N_16020,N_18865);
or U20980 (N_20980,N_19383,N_15633);
xor U20981 (N_20981,N_17769,N_17846);
or U20982 (N_20982,N_19393,N_17555);
and U20983 (N_20983,N_18594,N_16370);
or U20984 (N_20984,N_18528,N_17096);
nor U20985 (N_20985,N_15855,N_18786);
nand U20986 (N_20986,N_18690,N_16133);
or U20987 (N_20987,N_18392,N_16983);
and U20988 (N_20988,N_19241,N_15716);
nor U20989 (N_20989,N_17340,N_18593);
or U20990 (N_20990,N_18083,N_15679);
or U20991 (N_20991,N_19125,N_15723);
xor U20992 (N_20992,N_15796,N_15543);
xnor U20993 (N_20993,N_16174,N_17621);
and U20994 (N_20994,N_18581,N_16599);
nand U20995 (N_20995,N_16795,N_16464);
xnor U20996 (N_20996,N_19896,N_16419);
and U20997 (N_20997,N_16511,N_16001);
xor U20998 (N_20998,N_19376,N_18368);
and U20999 (N_20999,N_15707,N_16194);
and U21000 (N_21000,N_19664,N_15585);
nand U21001 (N_21001,N_18589,N_19028);
nor U21002 (N_21002,N_17367,N_15913);
nor U21003 (N_21003,N_16071,N_16308);
xnor U21004 (N_21004,N_16610,N_17154);
or U21005 (N_21005,N_18105,N_19988);
or U21006 (N_21006,N_17146,N_15795);
nand U21007 (N_21007,N_17443,N_15093);
or U21008 (N_21008,N_16856,N_19634);
or U21009 (N_21009,N_18644,N_16973);
and U21010 (N_21010,N_16460,N_16605);
nor U21011 (N_21011,N_18073,N_16487);
and U21012 (N_21012,N_17131,N_18882);
or U21013 (N_21013,N_15562,N_16363);
and U21014 (N_21014,N_19121,N_16007);
xor U21015 (N_21015,N_15234,N_16119);
nor U21016 (N_21016,N_15088,N_19846);
or U21017 (N_21017,N_18747,N_18271);
and U21018 (N_21018,N_15691,N_19862);
nor U21019 (N_21019,N_15113,N_19877);
nand U21020 (N_21020,N_18174,N_15889);
nor U21021 (N_21021,N_19954,N_19213);
and U21022 (N_21022,N_17296,N_18002);
or U21023 (N_21023,N_19023,N_19908);
and U21024 (N_21024,N_15013,N_15142);
or U21025 (N_21025,N_15849,N_15963);
and U21026 (N_21026,N_16005,N_17499);
and U21027 (N_21027,N_16330,N_18351);
or U21028 (N_21028,N_16493,N_19513);
xnor U21029 (N_21029,N_15035,N_19785);
nand U21030 (N_21030,N_17855,N_17480);
and U21031 (N_21031,N_17472,N_17428);
and U21032 (N_21032,N_18278,N_19754);
nor U21033 (N_21033,N_17465,N_19391);
nor U21034 (N_21034,N_16654,N_19760);
nand U21035 (N_21035,N_17578,N_17284);
and U21036 (N_21036,N_19947,N_16226);
or U21037 (N_21037,N_15925,N_15081);
and U21038 (N_21038,N_15854,N_19172);
and U21039 (N_21039,N_16789,N_17032);
and U21040 (N_21040,N_19171,N_16080);
or U21041 (N_21041,N_18843,N_18651);
xor U21042 (N_21042,N_19456,N_17138);
nand U21043 (N_21043,N_15805,N_18336);
nand U21044 (N_21044,N_19304,N_16551);
nand U21045 (N_21045,N_17143,N_18498);
nor U21046 (N_21046,N_17613,N_16649);
or U21047 (N_21047,N_19585,N_18471);
and U21048 (N_21048,N_15096,N_19731);
xor U21049 (N_21049,N_18103,N_16105);
nand U21050 (N_21050,N_15923,N_19114);
nand U21051 (N_21051,N_19829,N_19288);
or U21052 (N_21052,N_17229,N_17175);
xnor U21053 (N_21053,N_16222,N_19727);
and U21054 (N_21054,N_16145,N_18719);
nor U21055 (N_21055,N_17895,N_17350);
nor U21056 (N_21056,N_19088,N_15190);
nor U21057 (N_21057,N_18694,N_18776);
or U21058 (N_21058,N_16669,N_19089);
and U21059 (N_21059,N_18565,N_19218);
nand U21060 (N_21060,N_17261,N_19716);
and U21061 (N_21061,N_15109,N_17085);
nor U21062 (N_21062,N_18567,N_17251);
nor U21063 (N_21063,N_16069,N_16052);
and U21064 (N_21064,N_19625,N_16472);
nor U21065 (N_21065,N_19219,N_17940);
or U21066 (N_21066,N_18316,N_16261);
or U21067 (N_21067,N_16488,N_17960);
and U21068 (N_21068,N_16920,N_19854);
and U21069 (N_21069,N_18413,N_15812);
and U21070 (N_21070,N_17399,N_15010);
nor U21071 (N_21071,N_19604,N_15896);
nor U21072 (N_21072,N_16565,N_17349);
and U21073 (N_21073,N_18328,N_19998);
nand U21074 (N_21074,N_15539,N_17217);
or U21075 (N_21075,N_19061,N_15018);
nor U21076 (N_21076,N_15642,N_19371);
or U21077 (N_21077,N_15394,N_17817);
and U21078 (N_21078,N_16775,N_17861);
nand U21079 (N_21079,N_16344,N_18864);
nor U21080 (N_21080,N_16576,N_16434);
nor U21081 (N_21081,N_18995,N_15786);
xnor U21082 (N_21082,N_15801,N_17307);
or U21083 (N_21083,N_19955,N_15868);
or U21084 (N_21084,N_15260,N_19748);
and U21085 (N_21085,N_15583,N_18640);
or U21086 (N_21086,N_17221,N_15135);
nor U21087 (N_21087,N_18056,N_16619);
nand U21088 (N_21088,N_17948,N_17637);
or U21089 (N_21089,N_18647,N_19755);
nand U21090 (N_21090,N_19501,N_15080);
nand U21091 (N_21091,N_15655,N_15573);
nor U21092 (N_21092,N_19788,N_15946);
xor U21093 (N_21093,N_19971,N_19208);
and U21094 (N_21094,N_18571,N_16414);
and U21095 (N_21095,N_16266,N_19285);
or U21096 (N_21096,N_17450,N_15372);
nand U21097 (N_21097,N_16593,N_16823);
xor U21098 (N_21098,N_18561,N_17036);
nor U21099 (N_21099,N_19277,N_15488);
nor U21100 (N_21100,N_17687,N_17554);
and U21101 (N_21101,N_18504,N_18623);
or U21102 (N_21102,N_16448,N_15702);
nor U21103 (N_21103,N_16482,N_17049);
nand U21104 (N_21104,N_17614,N_19512);
and U21105 (N_21105,N_15708,N_18163);
nor U21106 (N_21106,N_15994,N_19596);
or U21107 (N_21107,N_18214,N_15223);
and U21108 (N_21108,N_18986,N_18059);
nand U21109 (N_21109,N_18723,N_15670);
nor U21110 (N_21110,N_15516,N_15242);
nand U21111 (N_21111,N_15225,N_18407);
nor U21112 (N_21112,N_17518,N_18749);
nand U21113 (N_21113,N_17183,N_15620);
nand U21114 (N_21114,N_16035,N_16046);
nand U21115 (N_21115,N_15313,N_19477);
nand U21116 (N_21116,N_17802,N_15243);
or U21117 (N_21117,N_16570,N_17601);
nand U21118 (N_21118,N_18933,N_15029);
nor U21119 (N_21119,N_17523,N_16603);
xor U21120 (N_21120,N_19531,N_19046);
and U21121 (N_21121,N_16387,N_15618);
nand U21122 (N_21122,N_19423,N_16512);
and U21123 (N_21123,N_18300,N_15650);
nor U21124 (N_21124,N_19758,N_18160);
nand U21125 (N_21125,N_16694,N_17737);
nand U21126 (N_21126,N_15037,N_17348);
or U21127 (N_21127,N_18340,N_18541);
and U21128 (N_21128,N_15239,N_16038);
nand U21129 (N_21129,N_17292,N_16661);
nor U21130 (N_21130,N_19281,N_18053);
or U21131 (N_21131,N_19842,N_17200);
nand U21132 (N_21132,N_18692,N_16501);
and U21133 (N_21133,N_17870,N_19057);
and U21134 (N_21134,N_15687,N_17584);
nand U21135 (N_21135,N_19269,N_15972);
and U21136 (N_21136,N_16059,N_19843);
nor U21137 (N_21137,N_18928,N_19930);
and U21138 (N_21138,N_19650,N_17269);
or U21139 (N_21139,N_19977,N_19462);
and U21140 (N_21140,N_19888,N_17593);
or U21141 (N_21141,N_16343,N_15314);
or U21142 (N_21142,N_18012,N_19453);
nand U21143 (N_21143,N_15593,N_18724);
nor U21144 (N_21144,N_15426,N_17676);
or U21145 (N_21145,N_17557,N_18403);
or U21146 (N_21146,N_18452,N_19446);
or U21147 (N_21147,N_16810,N_15980);
or U21148 (N_21148,N_18886,N_17919);
nand U21149 (N_21149,N_17462,N_15030);
nor U21150 (N_21150,N_17124,N_15089);
nor U21151 (N_21151,N_15617,N_16756);
or U21152 (N_21152,N_19186,N_17767);
or U21153 (N_21153,N_18645,N_17426);
or U21154 (N_21154,N_15199,N_18525);
nand U21155 (N_21155,N_15696,N_16033);
nand U21156 (N_21156,N_19292,N_19425);
or U21157 (N_21157,N_18914,N_19589);
nand U21158 (N_21158,N_18410,N_18680);
nand U21159 (N_21159,N_18608,N_16987);
nand U21160 (N_21160,N_18356,N_18892);
nor U21161 (N_21161,N_16183,N_17528);
or U21162 (N_21162,N_16009,N_16915);
and U21163 (N_21163,N_19291,N_18295);
and U21164 (N_21164,N_18638,N_18419);
and U21165 (N_21165,N_16818,N_15779);
xnor U21166 (N_21166,N_17278,N_17749);
nor U21167 (N_21167,N_18803,N_17300);
and U21168 (N_21168,N_19865,N_18702);
or U21169 (N_21169,N_19019,N_18670);
and U21170 (N_21170,N_18658,N_15231);
nor U21171 (N_21171,N_15511,N_17667);
xnor U21172 (N_21172,N_15602,N_17415);
and U21173 (N_21173,N_15047,N_15898);
nand U21174 (N_21174,N_15637,N_15051);
nand U21175 (N_21175,N_17768,N_16006);
xnor U21176 (N_21176,N_17911,N_19873);
and U21177 (N_21177,N_19773,N_19928);
or U21178 (N_21178,N_15077,N_18421);
xnor U21179 (N_21179,N_19807,N_17726);
nor U21180 (N_21180,N_19686,N_18835);
nor U21181 (N_21181,N_18360,N_17362);
nand U21182 (N_21182,N_15353,N_17081);
nand U21183 (N_21183,N_15144,N_15398);
and U21184 (N_21184,N_17391,N_19138);
nand U21185 (N_21185,N_18422,N_16054);
and U21186 (N_21186,N_18969,N_15918);
nor U21187 (N_21187,N_15067,N_15112);
nor U21188 (N_21188,N_16239,N_18492);
nor U21189 (N_21189,N_17026,N_19111);
xor U21190 (N_21190,N_19682,N_18729);
nand U21191 (N_21191,N_16403,N_18794);
nand U21192 (N_21192,N_16682,N_18077);
nand U21193 (N_21193,N_19246,N_17790);
nor U21194 (N_21194,N_15317,N_18754);
and U21195 (N_21195,N_17840,N_17653);
or U21196 (N_21196,N_18341,N_16633);
and U21197 (N_21197,N_16705,N_17048);
xnor U21198 (N_21198,N_18243,N_16714);
and U21199 (N_21199,N_17604,N_15824);
and U21200 (N_21200,N_17752,N_19463);
xor U21201 (N_21201,N_18506,N_18244);
or U21202 (N_21202,N_16542,N_17139);
and U21203 (N_21203,N_18399,N_16190);
and U21204 (N_21204,N_19064,N_18208);
nand U21205 (N_21205,N_17702,N_18992);
and U21206 (N_21206,N_16381,N_18180);
nand U21207 (N_21207,N_15768,N_15973);
nand U21208 (N_21208,N_16824,N_19607);
nor U21209 (N_21209,N_18157,N_19287);
nor U21210 (N_21210,N_17467,N_16847);
xor U21211 (N_21211,N_17176,N_18329);
or U21212 (N_21212,N_19958,N_15049);
nand U21213 (N_21213,N_15380,N_19713);
nand U21214 (N_21214,N_15479,N_15666);
nor U21215 (N_21215,N_17168,N_19543);
nand U21216 (N_21216,N_19496,N_15665);
and U21217 (N_21217,N_18357,N_15532);
nor U21218 (N_21218,N_17098,N_19490);
and U21219 (N_21219,N_17582,N_19905);
or U21220 (N_21220,N_18529,N_15357);
nand U21221 (N_21221,N_15899,N_17037);
or U21222 (N_21222,N_15787,N_18523);
nand U21223 (N_21223,N_17457,N_15250);
nand U21224 (N_21224,N_15420,N_17858);
and U21225 (N_21225,N_17996,N_18580);
nor U21226 (N_21226,N_16251,N_17312);
nand U21227 (N_21227,N_19374,N_18354);
or U21228 (N_21228,N_18745,N_18604);
nand U21229 (N_21229,N_17910,N_16585);
nor U21230 (N_21230,N_15639,N_17881);
and U21231 (N_21231,N_18813,N_17914);
nand U21232 (N_21232,N_18563,N_18280);
and U21233 (N_21233,N_16221,N_15698);
nor U21234 (N_21234,N_17657,N_15667);
nor U21235 (N_21235,N_18445,N_17038);
and U21236 (N_21236,N_18159,N_19981);
or U21237 (N_21237,N_16092,N_18874);
nand U21238 (N_21238,N_17459,N_19078);
and U21239 (N_21239,N_16178,N_17448);
and U21240 (N_21240,N_19377,N_16764);
and U21241 (N_21241,N_19734,N_17320);
nor U21242 (N_21242,N_17973,N_17118);
or U21243 (N_21243,N_18202,N_17579);
nand U21244 (N_21244,N_18308,N_16627);
nand U21245 (N_21245,N_18450,N_16578);
xor U21246 (N_21246,N_16275,N_15184);
and U21247 (N_21247,N_19166,N_15968);
or U21248 (N_21248,N_15791,N_16045);
and U21249 (N_21249,N_18363,N_19144);
nand U21250 (N_21250,N_19084,N_16835);
nand U21251 (N_21251,N_19953,N_18347);
or U21252 (N_21252,N_16152,N_15404);
nor U21253 (N_21253,N_18350,N_15738);
xor U21254 (N_21254,N_15214,N_17270);
xnor U21255 (N_21255,N_15971,N_16300);
or U21256 (N_21256,N_17437,N_17432);
nand U21257 (N_21257,N_16028,N_15172);
or U21258 (N_21258,N_18908,N_19933);
and U21259 (N_21259,N_19485,N_16838);
nor U21260 (N_21260,N_15408,N_15948);
nor U21261 (N_21261,N_17313,N_17754);
and U21262 (N_21262,N_18216,N_16965);
nor U21263 (N_21263,N_18200,N_18039);
or U21264 (N_21264,N_19040,N_19900);
nand U21265 (N_21265,N_19384,N_16171);
nand U21266 (N_21266,N_16623,N_17544);
or U21267 (N_21267,N_19675,N_19204);
xnor U21268 (N_21268,N_15278,N_17872);
nor U21269 (N_21269,N_17333,N_18550);
and U21270 (N_21270,N_17988,N_15953);
nor U21271 (N_21271,N_16158,N_19131);
or U21272 (N_21272,N_19014,N_16925);
or U21273 (N_21273,N_17073,N_19147);
and U21274 (N_21274,N_16588,N_18472);
nand U21275 (N_21275,N_18201,N_17335);
nor U21276 (N_21276,N_19938,N_15673);
nor U21277 (N_21277,N_16751,N_19388);
nand U21278 (N_21278,N_18698,N_17577);
nor U21279 (N_21279,N_17047,N_15186);
nor U21280 (N_21280,N_15435,N_17374);
nand U21281 (N_21281,N_15450,N_18863);
nand U21282 (N_21282,N_18733,N_18016);
xnor U21283 (N_21283,N_15461,N_15671);
and U21284 (N_21284,N_18988,N_15439);
xnor U21285 (N_21285,N_15700,N_18480);
xor U21286 (N_21286,N_18442,N_16613);
xnor U21287 (N_21287,N_19893,N_18990);
nand U21288 (N_21288,N_17507,N_17075);
or U21289 (N_21289,N_17644,N_16422);
or U21290 (N_21290,N_19473,N_18771);
or U21291 (N_21291,N_16933,N_17025);
or U21292 (N_21292,N_18912,N_18785);
xor U21293 (N_21293,N_19200,N_18247);
nor U21294 (N_21294,N_17529,N_16582);
and U21295 (N_21295,N_18061,N_15383);
nand U21296 (N_21296,N_17004,N_19961);
nor U21297 (N_21297,N_15146,N_17233);
nand U21298 (N_21298,N_16286,N_17065);
nand U21299 (N_21299,N_17972,N_18521);
nand U21300 (N_21300,N_15880,N_17015);
nor U21301 (N_21301,N_15756,N_15356);
and U21302 (N_21302,N_19181,N_18117);
xor U21303 (N_21303,N_18313,N_17566);
nor U21304 (N_21304,N_16025,N_19638);
or U21305 (N_21305,N_19253,N_19362);
nand U21306 (N_21306,N_16683,N_16812);
or U21307 (N_21307,N_18307,N_18319);
nor U21308 (N_21308,N_16962,N_18852);
nor U21309 (N_21309,N_19706,N_16990);
or U21310 (N_21310,N_16144,N_15136);
nand U21311 (N_21311,N_17327,N_19895);
or U21312 (N_21312,N_19417,N_17268);
nor U21313 (N_21313,N_19401,N_17421);
nand U21314 (N_21314,N_15823,N_16041);
or U21315 (N_21315,N_15850,N_15235);
nand U21316 (N_21316,N_16307,N_16791);
or U21317 (N_21317,N_17418,N_19332);
nor U21318 (N_21318,N_17747,N_15591);
and U21319 (N_21319,N_17180,N_17484);
xnor U21320 (N_21320,N_17108,N_16864);
and U21321 (N_21321,N_17031,N_15438);
and U21322 (N_21322,N_19777,N_16979);
or U21323 (N_21323,N_19175,N_17852);
nand U21324 (N_21324,N_17171,N_15271);
and U21325 (N_21325,N_17308,N_18097);
and U21326 (N_21326,N_18939,N_19932);
xnor U21327 (N_21327,N_15584,N_15883);
or U21328 (N_21328,N_15429,N_16058);
and U21329 (N_21329,N_19329,N_19437);
xor U21330 (N_21330,N_15830,N_19160);
xnor U21331 (N_21331,N_18482,N_19267);
xor U21332 (N_21332,N_19964,N_18234);
nand U21333 (N_21333,N_17947,N_19841);
or U21334 (N_21334,N_17928,N_19141);
and U21335 (N_21335,N_19671,N_18172);
or U21336 (N_21336,N_16157,N_16349);
nor U21337 (N_21337,N_18902,N_19632);
nand U21338 (N_21338,N_19251,N_15045);
xnor U21339 (N_21339,N_19297,N_15597);
or U21340 (N_21340,N_15211,N_17605);
and U21341 (N_21341,N_18998,N_18409);
or U21342 (N_21342,N_16214,N_18709);
or U21343 (N_21343,N_17865,N_17813);
nor U21344 (N_21344,N_18691,N_17409);
nor U21345 (N_21345,N_16822,N_18303);
or U21346 (N_21346,N_15657,N_15374);
and U21347 (N_21347,N_19293,N_15903);
or U21348 (N_21348,N_16316,N_19571);
nand U21349 (N_21349,N_19062,N_19665);
nor U21350 (N_21350,N_18366,N_15552);
xnor U21351 (N_21351,N_17352,N_18245);
nand U21352 (N_21352,N_17353,N_16561);
or U21353 (N_21353,N_17056,N_17043);
and U21354 (N_21354,N_16392,N_19352);
nand U21355 (N_21355,N_18401,N_15063);
nand U21356 (N_21356,N_16507,N_19643);
nand U21357 (N_21357,N_18381,N_16215);
or U21358 (N_21358,N_19075,N_18253);
nor U21359 (N_21359,N_15267,N_18236);
or U21360 (N_21360,N_16583,N_17133);
nor U21361 (N_21361,N_19359,N_15531);
nor U21362 (N_21362,N_19636,N_15536);
and U21363 (N_21363,N_15467,N_19274);
nor U21364 (N_21364,N_16489,N_17799);
or U21365 (N_21365,N_17470,N_15631);
xor U21366 (N_21366,N_19899,N_18858);
nor U21367 (N_21367,N_15921,N_15099);
xnor U21368 (N_21368,N_16070,N_19308);
nand U21369 (N_21369,N_15933,N_18438);
and U21370 (N_21370,N_19278,N_15453);
and U21371 (N_21371,N_16898,N_16023);
nand U21372 (N_21372,N_17724,N_18987);
or U21373 (N_21373,N_15409,N_15122);
xor U21374 (N_21374,N_17734,N_15882);
and U21375 (N_21375,N_18683,N_19076);
and U21376 (N_21376,N_16957,N_16048);
or U21377 (N_21377,N_17757,N_15675);
nand U21378 (N_21378,N_18389,N_18898);
or U21379 (N_21379,N_19416,N_18925);
nand U21380 (N_21380,N_16888,N_15457);
or U21381 (N_21381,N_17092,N_17514);
nand U21382 (N_21382,N_19091,N_15520);
or U21383 (N_21383,N_19460,N_16801);
nand U21384 (N_21384,N_16333,N_19819);
and U21385 (N_21385,N_16115,N_15793);
nor U21386 (N_21386,N_19715,N_18110);
nand U21387 (N_21387,N_19749,N_18873);
or U21388 (N_21388,N_17020,N_19929);
nand U21389 (N_21389,N_17306,N_15098);
and U21390 (N_21390,N_17763,N_19110);
or U21391 (N_21391,N_18404,N_17807);
and U21392 (N_21392,N_15518,N_15192);
nand U21393 (N_21393,N_18960,N_19816);
nor U21394 (N_21394,N_18913,N_15299);
nor U21395 (N_21395,N_17880,N_16527);
nor U21396 (N_21396,N_16252,N_16740);
nand U21397 (N_21397,N_15416,N_17863);
nand U21398 (N_21398,N_17839,N_18697);
nand U21399 (N_21399,N_17513,N_18008);
and U21400 (N_21400,N_16083,N_16206);
nand U21401 (N_21401,N_16137,N_18905);
nor U21402 (N_21402,N_15513,N_17628);
and U21403 (N_21403,N_19165,N_18774);
nand U21404 (N_21404,N_19461,N_16305);
nor U21405 (N_21405,N_17612,N_17389);
nand U21406 (N_21406,N_15802,N_19464);
and U21407 (N_21407,N_19397,N_19280);
nor U21408 (N_21408,N_15851,N_16429);
and U21409 (N_21409,N_17134,N_19424);
nand U21410 (N_21410,N_19031,N_17354);
and U21411 (N_21411,N_18868,N_17224);
and U21412 (N_21412,N_15767,N_17106);
nand U21413 (N_21413,N_16376,N_15402);
nor U21414 (N_21414,N_17622,N_19033);
and U21415 (N_21415,N_18415,N_17382);
or U21416 (N_21416,N_18265,N_19753);
nand U21417 (N_21417,N_15807,N_17275);
or U21418 (N_21418,N_18252,N_19418);
and U21419 (N_21419,N_16875,N_19045);
nor U21420 (N_21420,N_17608,N_16562);
and U21421 (N_21421,N_16763,N_15482);
and U21422 (N_21422,N_17583,N_19526);
and U21423 (N_21423,N_18540,N_16299);
or U21424 (N_21424,N_17347,N_15724);
and U21425 (N_21425,N_16589,N_18814);
and U21426 (N_21426,N_17884,N_19780);
or U21427 (N_21427,N_19207,N_16461);
xnor U21428 (N_21428,N_15233,N_17740);
nand U21429 (N_21429,N_19096,N_15627);
and U21430 (N_21430,N_18673,N_17487);
and U21431 (N_21431,N_19880,N_19242);
or U21432 (N_21432,N_18901,N_16371);
nor U21433 (N_21433,N_17394,N_15634);
or U21434 (N_21434,N_16862,N_16988);
or U21435 (N_21435,N_17111,N_17185);
nor U21436 (N_21436,N_17879,N_15336);
nand U21437 (N_21437,N_15826,N_16067);
nor U21438 (N_21438,N_18106,N_17674);
nor U21439 (N_21439,N_19914,N_17782);
nor U21440 (N_21440,N_16506,N_16471);
or U21441 (N_21441,N_18826,N_19041);
or U21442 (N_21442,N_18038,N_17753);
nand U21443 (N_21443,N_19326,N_17822);
and U21444 (N_21444,N_18687,N_17247);
nand U21445 (N_21445,N_19991,N_15625);
nand U21446 (N_21446,N_15596,N_19872);
or U21447 (N_21447,N_17330,N_15194);
or U21448 (N_21448,N_18040,N_16591);
and U21449 (N_21449,N_18722,N_15232);
nand U21450 (N_21450,N_16653,N_15572);
nor U21451 (N_21451,N_17433,N_18209);
or U21452 (N_21452,N_16094,N_15846);
or U21453 (N_21453,N_15290,N_17190);
nand U21454 (N_21454,N_18742,N_15821);
and U21455 (N_21455,N_18194,N_17164);
nand U21456 (N_21456,N_18856,N_17862);
nand U21457 (N_21457,N_15581,N_18588);
nor U21458 (N_21458,N_16196,N_17646);
nor U21459 (N_21459,N_16072,N_19025);
nand U21460 (N_21460,N_17580,N_18848);
or U21461 (N_21461,N_16900,N_19836);
xnor U21462 (N_21462,N_16536,N_16663);
nand U21463 (N_21463,N_17051,N_18361);
and U21464 (N_21464,N_17303,N_19029);
or U21465 (N_21465,N_17012,N_19641);
or U21466 (N_21466,N_17510,N_16709);
nand U21467 (N_21467,N_15213,N_15992);
nor U21468 (N_21468,N_18127,N_17466);
nand U21469 (N_21469,N_18464,N_15686);
nor U21470 (N_21470,N_15360,N_19891);
xnor U21471 (N_21471,N_19498,N_18968);
or U21472 (N_21472,N_18979,N_18718);
nand U21473 (N_21473,N_18003,N_15207);
nor U21474 (N_21474,N_16093,N_18344);
and U21475 (N_21475,N_19282,N_17304);
or U21476 (N_21476,N_16744,N_15976);
or U21477 (N_21477,N_16207,N_18397);
or U21478 (N_21478,N_15021,N_16036);
nor U21479 (N_21479,N_17101,N_16597);
nor U21480 (N_21480,N_15537,N_19618);
nor U21481 (N_21481,N_15462,N_16703);
and U21482 (N_21482,N_15352,N_15188);
or U21483 (N_21483,N_16814,N_17547);
or U21484 (N_21484,N_19053,N_17641);
or U21485 (N_21485,N_16702,N_15480);
or U21486 (N_21486,N_17703,N_17218);
xor U21487 (N_21487,N_19847,N_18218);
or U21488 (N_21488,N_17866,N_18241);
or U21489 (N_21489,N_16509,N_17310);
or U21490 (N_21490,N_17508,N_17833);
nand U21491 (N_21491,N_16044,N_16718);
and U21492 (N_21492,N_19787,N_17370);
or U21493 (N_21493,N_18122,N_18840);
and U21494 (N_21494,N_17828,N_15206);
xnor U21495 (N_21495,N_16142,N_17789);
and U21496 (N_21496,N_15078,N_17419);
xnor U21497 (N_21497,N_18751,N_15521);
and U21498 (N_21498,N_15681,N_19859);
and U21499 (N_21499,N_17211,N_18507);
nand U21500 (N_21500,N_15204,N_19521);
and U21501 (N_21501,N_17836,N_15072);
or U21502 (N_21502,N_19164,N_16976);
nand U21503 (N_21503,N_15559,N_17827);
nor U21504 (N_21504,N_15272,N_19850);
and U21505 (N_21505,N_16538,N_17594);
or U21506 (N_21506,N_16636,N_15002);
or U21507 (N_21507,N_15555,N_17803);
xor U21508 (N_21508,N_15296,N_15498);
or U21509 (N_21509,N_16126,N_16314);
nor U21510 (N_21510,N_16722,N_17669);
or U21511 (N_21511,N_19101,N_19334);
nor U21512 (N_21512,N_15471,N_17153);
nor U21513 (N_21513,N_15226,N_18894);
nor U21514 (N_21514,N_16289,N_16871);
and U21515 (N_21515,N_18348,N_18084);
nor U21516 (N_21516,N_15092,N_18485);
and U21517 (N_21517,N_19158,N_17385);
nor U21518 (N_21518,N_15276,N_17572);
nor U21519 (N_21519,N_16666,N_16754);
or U21520 (N_21520,N_15560,N_17386);
nor U21521 (N_21521,N_17458,N_17944);
or U21522 (N_21522,N_19610,N_15171);
xnor U21523 (N_21523,N_19163,N_17495);
nand U21524 (N_21524,N_19344,N_16678);
or U21525 (N_21525,N_15054,N_19655);
nand U21526 (N_21526,N_16154,N_18027);
or U21527 (N_21527,N_19594,N_18034);
and U21528 (N_21528,N_15895,N_19472);
nor U21529 (N_21529,N_15920,N_19066);
and U21530 (N_21530,N_16327,N_15154);
nor U21531 (N_21531,N_17568,N_15571);
xnor U21532 (N_21532,N_16552,N_18653);
and U21533 (N_21533,N_18481,N_16928);
and U21534 (N_21534,N_16541,N_19107);
or U21535 (N_21535,N_15599,N_15609);
nand U21536 (N_21536,N_16415,N_16780);
nor U21537 (N_21537,N_19245,N_18839);
xor U21538 (N_21538,N_18161,N_17695);
or U21539 (N_21539,N_19054,N_15522);
nor U21540 (N_21540,N_18795,N_17091);
or U21541 (N_21541,N_15557,N_16514);
or U21542 (N_21542,N_16467,N_16690);
and U21543 (N_21543,N_19614,N_17250);
or U21544 (N_21544,N_18052,N_15046);
nor U21545 (N_21545,N_16999,N_19704);
nor U21546 (N_21546,N_18156,N_19795);
xnor U21547 (N_21547,N_18250,N_15765);
nand U21548 (N_21548,N_16759,N_17927);
nand U21549 (N_21549,N_19703,N_16713);
nor U21550 (N_21550,N_17130,N_19904);
nor U21551 (N_21551,N_18449,N_17478);
nand U21552 (N_21552,N_19921,N_15790);
or U21553 (N_21553,N_19656,N_18302);
or U21554 (N_21554,N_16728,N_15200);
and U21555 (N_21555,N_16155,N_15274);
xnor U21556 (N_21556,N_17334,N_18479);
and U21557 (N_21557,N_17314,N_16247);
xor U21558 (N_21558,N_18603,N_17271);
and U21559 (N_21559,N_18074,N_16515);
nor U21560 (N_21560,N_17243,N_18312);
or U21561 (N_21561,N_17706,N_19483);
nor U21562 (N_21562,N_18616,N_18682);
nor U21563 (N_21563,N_17445,N_18044);
or U21564 (N_21564,N_16131,N_19603);
or U21565 (N_21565,N_17663,N_18695);
nor U21566 (N_21566,N_17854,N_18538);
nor U21567 (N_21567,N_16346,N_16268);
nand U21568 (N_21568,N_15624,N_18962);
nor U21569 (N_21569,N_18017,N_15365);
or U21570 (N_21570,N_19395,N_17326);
or U21571 (N_21571,N_15427,N_17901);
nor U21572 (N_21572,N_15405,N_19035);
xor U21573 (N_21573,N_15544,N_19926);
and U21574 (N_21574,N_17524,N_16883);
or U21575 (N_21575,N_19534,N_18989);
or U21576 (N_21576,N_17625,N_16699);
or U21577 (N_21577,N_17184,N_18373);
nor U21578 (N_21578,N_18146,N_15563);
and U21579 (N_21579,N_16969,N_15527);
nor U21580 (N_21580,N_19838,N_15445);
xor U21581 (N_21581,N_16601,N_19060);
or U21582 (N_21582,N_15839,N_19507);
nor U21583 (N_21583,N_16010,N_15668);
or U21584 (N_21584,N_18952,N_17309);
nor U21585 (N_21585,N_19369,N_15857);
xnor U21586 (N_21586,N_15608,N_16880);
or U21587 (N_21587,N_19630,N_15265);
nor U21588 (N_21588,N_16995,N_19672);
or U21589 (N_21589,N_18855,N_19901);
nor U21590 (N_21590,N_17117,N_18182);
nand U21591 (N_21591,N_17647,N_17725);
nor U21592 (N_21592,N_19289,N_16426);
or U21593 (N_21593,N_18113,N_18564);
or U21594 (N_21594,N_16640,N_16393);
and U21595 (N_21595,N_17730,N_18656);
or U21596 (N_21596,N_18878,N_18026);
nand U21597 (N_21597,N_18023,N_17244);
or U21598 (N_21598,N_15273,N_17874);
nand U21599 (N_21599,N_17402,N_15816);
and U21600 (N_21600,N_15401,N_17720);
or U21601 (N_21601,N_19640,N_16635);
nand U21602 (N_21602,N_18444,N_17192);
and U21603 (N_21603,N_18320,N_15392);
nor U21604 (N_21604,N_17905,N_18509);
nor U21605 (N_21605,N_17684,N_16177);
nand U21606 (N_21606,N_15494,N_19518);
or U21607 (N_21607,N_16240,N_16086);
xor U21608 (N_21608,N_15619,N_19261);
and U21609 (N_21609,N_15459,N_15275);
nor U21610 (N_21610,N_19363,N_18505);
xnor U21611 (N_21611,N_15991,N_18860);
and U21612 (N_21612,N_19003,N_15008);
nand U21613 (N_21613,N_18801,N_17638);
nand U21614 (N_21614,N_17887,N_19434);
xor U21615 (N_21615,N_19994,N_19260);
nor U21616 (N_21616,N_17444,N_15798);
and U21617 (N_21617,N_18123,N_17896);
or U21618 (N_21618,N_15653,N_15761);
and U21619 (N_21619,N_17392,N_15870);
nand U21620 (N_21620,N_15588,N_19225);
nor U21621 (N_21621,N_16096,N_16077);
nand U21622 (N_21622,N_16692,N_16087);
xor U21623 (N_21623,N_16329,N_19449);
and U21624 (N_21624,N_16815,N_16564);
nand U21625 (N_21625,N_17899,N_15095);
or U21626 (N_21626,N_19196,N_19674);
nand U21627 (N_21627,N_15262,N_18661);
nand U21628 (N_21628,N_17793,N_15837);
nor U21629 (N_21629,N_18539,N_18094);
nor U21630 (N_21630,N_17750,N_15550);
and U21631 (N_21631,N_16320,N_17902);
or U21632 (N_21632,N_17626,N_15733);
and U21633 (N_21633,N_19556,N_19959);
nand U21634 (N_21634,N_17984,N_15877);
or U21635 (N_21635,N_17114,N_15381);
or U21636 (N_21636,N_17982,N_16879);
and U21637 (N_21637,N_19394,N_18435);
nand U21638 (N_21638,N_19583,N_16938);
nand U21639 (N_21639,N_19925,N_18187);
nand U21640 (N_21640,N_19677,N_19205);
and U21641 (N_21641,N_17103,N_16444);
or U21642 (N_21642,N_17255,N_19874);
nor U21643 (N_21643,N_15935,N_17704);
nand U21644 (N_21644,N_16163,N_19099);
or U21645 (N_21645,N_19721,N_19744);
xnor U21646 (N_21646,N_18546,N_18118);
and U21647 (N_21647,N_17024,N_16495);
or U21648 (N_21648,N_19951,N_15216);
and U21649 (N_21649,N_16016,N_19920);
xor U21650 (N_21650,N_18024,N_16359);
xor U21651 (N_21651,N_19927,N_17530);
nand U21652 (N_21652,N_16011,N_19093);
xnor U21653 (N_21653,N_15663,N_16354);
or U21654 (N_21654,N_19059,N_16817);
and U21655 (N_21655,N_17715,N_19828);
and U21656 (N_21656,N_16022,N_16846);
or U21657 (N_21657,N_15107,N_16253);
nand U21658 (N_21658,N_17181,N_18781);
nor U21659 (N_21659,N_19270,N_19979);
or U21660 (N_21660,N_16149,N_19832);
nor U21661 (N_21661,N_15345,N_17365);
and U21662 (N_21662,N_17149,N_19439);
nor U21663 (N_21663,N_16076,N_19108);
nand U21664 (N_21664,N_17017,N_16172);
nand U21665 (N_21665,N_16180,N_15764);
and U21666 (N_21666,N_18267,N_15253);
xor U21667 (N_21667,N_19356,N_17115);
nand U21668 (N_21668,N_17080,N_19192);
xnor U21669 (N_21669,N_15676,N_17186);
nor U21670 (N_21670,N_18179,N_18769);
or U21671 (N_21671,N_18660,N_15598);
nor U21672 (N_21672,N_15341,N_17254);
nand U21673 (N_21673,N_17965,N_16483);
or U21674 (N_21674,N_18283,N_19502);
xor U21675 (N_21675,N_18934,N_15662);
or U21676 (N_21676,N_19510,N_19690);
nor U21677 (N_21677,N_18678,N_15005);
nor U21678 (N_21678,N_16905,N_15565);
xor U21679 (N_21679,N_16088,N_15945);
and U21680 (N_21680,N_16537,N_16575);
and U21681 (N_21681,N_16436,N_16523);
and U21682 (N_21682,N_17742,N_15303);
or U21683 (N_21683,N_15710,N_17756);
nor U21684 (N_21684,N_19505,N_19523);
nand U21685 (N_21685,N_16985,N_15711);
and U21686 (N_21686,N_19950,N_15388);
xnor U21687 (N_21687,N_19124,N_16809);
nand U21688 (N_21688,N_18586,N_15912);
nor U21689 (N_21689,N_19009,N_18555);
nor U21690 (N_21690,N_17322,N_16765);
nor U21691 (N_21691,N_19342,N_18665);
or U21692 (N_21692,N_19960,N_16671);
nor U21693 (N_21693,N_18142,N_17660);
nand U21694 (N_21694,N_19934,N_18954);
nor U21695 (N_21695,N_15385,N_16110);
and U21696 (N_21696,N_16411,N_17027);
xor U21697 (N_21697,N_19153,N_16372);
nor U21698 (N_21698,N_19867,N_16854);
nor U21699 (N_21699,N_17744,N_17136);
nand U21700 (N_21700,N_16282,N_17596);
and U21701 (N_21701,N_17823,N_17624);
or U21702 (N_21702,N_16159,N_18029);
and U21703 (N_21703,N_18842,N_17820);
nor U21704 (N_21704,N_18376,N_19548);
xor U21705 (N_21705,N_17571,N_18949);
nand U21706 (N_21706,N_18706,N_18176);
nor U21707 (N_21707,N_16459,N_17848);
xor U21708 (N_21708,N_18630,N_19248);
nand U21709 (N_21709,N_18196,N_17105);
or U21710 (N_21710,N_15731,N_16348);
or U21711 (N_21711,N_15575,N_16960);
nand U21712 (N_21712,N_17675,N_17673);
or U21713 (N_21713,N_15149,N_15236);
and U21714 (N_21714,N_16923,N_19109);
or U21715 (N_21715,N_18309,N_16064);
and U21716 (N_21716,N_15229,N_16729);
or U21717 (N_21717,N_18069,N_19098);
or U21718 (N_21718,N_18872,N_18515);
nor U21719 (N_21719,N_17490,N_18675);
nand U21720 (N_21720,N_17416,N_17336);
xor U21721 (N_21721,N_16416,N_18714);
nor U21722 (N_21722,N_17002,N_17042);
xnor U21723 (N_21723,N_19826,N_18815);
nand U21724 (N_21724,N_17277,N_17745);
nor U21725 (N_21725,N_19648,N_16232);
nor U21726 (N_21726,N_15032,N_15995);
nand U21727 (N_21727,N_15084,N_17592);
nor U21728 (N_21728,N_18770,N_19569);
nand U21729 (N_21729,N_16328,N_15917);
xor U21730 (N_21730,N_17325,N_18937);
nor U21731 (N_21731,N_16790,N_19801);
nand U21732 (N_21732,N_17682,N_19724);
or U21733 (N_21733,N_19827,N_15719);
or U21734 (N_21734,N_19687,N_15412);
and U21735 (N_21735,N_16738,N_15615);
or U21736 (N_21736,N_15031,N_17515);
and U21737 (N_21737,N_17546,N_16989);
or U21738 (N_21738,N_19762,N_18598);
or U21739 (N_21739,N_17516,N_18926);
or U21740 (N_21740,N_17226,N_19482);
and U21741 (N_21741,N_19676,N_15845);
and U21742 (N_21742,N_15277,N_19806);
or U21743 (N_21743,N_19330,N_15337);
or U21744 (N_21744,N_16628,N_19396);
nor U21745 (N_21745,N_17562,N_17950);
and U21746 (N_21746,N_18635,N_16104);
nand U21747 (N_21747,N_16721,N_16655);
nor U21748 (N_21748,N_19426,N_15478);
nor U21749 (N_21749,N_16598,N_17366);
or U21750 (N_21750,N_19126,N_17069);
xnor U21751 (N_21751,N_18068,N_15362);
nor U21752 (N_21752,N_17239,N_18443);
nor U21753 (N_21753,N_16271,N_18611);
nor U21754 (N_21754,N_16066,N_15836);
nor U21755 (N_21755,N_16892,N_16934);
and U21756 (N_21756,N_18212,N_17276);
nand U21757 (N_21757,N_18305,N_15957);
or U21758 (N_21758,N_18111,N_19956);
or U21759 (N_21759,N_18696,N_16279);
nor U21760 (N_21760,N_19587,N_15124);
nor U21761 (N_21761,N_16337,N_17825);
nand U21762 (N_21762,N_16611,N_16505);
and U21763 (N_21763,N_17509,N_15843);
xnor U21764 (N_21764,N_15464,N_17710);
and U21765 (N_21765,N_15125,N_15871);
nor U21766 (N_21766,N_19857,N_16771);
nand U21767 (N_21767,N_17536,N_19557);
nand U21768 (N_21768,N_18701,N_18720);
or U21769 (N_21769,N_16169,N_15697);
or U21770 (N_21770,N_18092,N_16056);
or U21771 (N_21771,N_18386,N_17364);
or U21772 (N_21772,N_16793,N_19790);
nand U21773 (N_21773,N_18148,N_15169);
and U21774 (N_21774,N_18396,N_19412);
and U21775 (N_21775,N_17422,N_18837);
and U21776 (N_21776,N_18258,N_16231);
or U21777 (N_21777,N_15111,N_16440);
nand U21778 (N_21778,N_18533,N_18637);
or U21779 (N_21779,N_16034,N_17681);
and U21780 (N_21780,N_19851,N_16225);
nand U21781 (N_21781,N_15860,N_18314);
nor U21782 (N_21782,N_18255,N_16498);
nor U21783 (N_21783,N_18046,N_15904);
or U21784 (N_21784,N_16807,N_19480);
nor U21785 (N_21785,N_16235,N_15182);
nand U21786 (N_21786,N_15118,N_18641);
and U21787 (N_21787,N_17297,N_19037);
and U21788 (N_21788,N_16778,N_18367);
or U21789 (N_21789,N_19345,N_16797);
nand U21790 (N_21790,N_18311,N_19137);
and U21791 (N_21791,N_18152,N_19728);
and U21792 (N_21792,N_16710,N_18321);
and U21793 (N_21793,N_17958,N_18981);
nor U21794 (N_21794,N_16478,N_15950);
nor U21795 (N_21795,N_16160,N_19445);
nand U21796 (N_21796,N_16068,N_17369);
and U21797 (N_21797,N_15890,N_16465);
nand U21798 (N_21798,N_17781,N_15744);
nor U21799 (N_21799,N_16121,N_19221);
nor U21800 (N_21800,N_15212,N_15578);
and U21801 (N_21801,N_18967,N_19784);
nand U21802 (N_21802,N_18829,N_15556);
and U21803 (N_21803,N_15859,N_15217);
or U21804 (N_21804,N_16831,N_18150);
and U21805 (N_21805,N_17387,N_16332);
nor U21806 (N_21806,N_19206,N_15366);
nor U21807 (N_21807,N_15484,N_17492);
or U21808 (N_21808,N_17097,N_15878);
nand U21809 (N_21809,N_16761,N_16331);
or U21810 (N_21810,N_19619,N_17267);
nor U21811 (N_21811,N_15735,N_15417);
or U21812 (N_21812,N_15468,N_16596);
or U21813 (N_21813,N_15818,N_18836);
nor U21814 (N_21814,N_15926,N_19226);
nand U21815 (N_21815,N_19006,N_15187);
or U21816 (N_21816,N_17315,N_19405);
nor U21817 (N_21817,N_18909,N_18797);
and U21818 (N_21818,N_15130,N_15727);
nand U21819 (N_21819,N_15319,N_15056);
nor U21820 (N_21820,N_17137,N_19409);
nor U21821 (N_21821,N_18128,N_15373);
nor U21822 (N_21822,N_16285,N_17723);
nor U21823 (N_21823,N_15844,N_15333);
xnor U21824 (N_21824,N_15640,N_18248);
nor U21825 (N_21825,N_15421,N_15121);
nor U21826 (N_21826,N_19189,N_18618);
and U21827 (N_21827,N_19793,N_19669);
nand U21828 (N_21828,N_16130,N_15068);
or U21829 (N_21829,N_19481,N_15185);
nand U21830 (N_21830,N_16781,N_17401);
and U21831 (N_21831,N_18107,N_17925);
or U21832 (N_21832,N_16530,N_17317);
nor U21833 (N_21833,N_16908,N_19527);
or U21834 (N_21834,N_15400,N_18916);
and U21835 (N_21835,N_16647,N_19312);
and U21836 (N_21836,N_17373,N_19310);
or U21837 (N_21837,N_18677,N_17736);
and U21838 (N_21838,N_19633,N_17280);
nand U21839 (N_21839,N_17511,N_17694);
nor U21840 (N_21840,N_15268,N_19263);
nor U21841 (N_21841,N_16111,N_16882);
xor U21842 (N_21842,N_19764,N_16737);
xor U21843 (N_21843,N_15041,N_16224);
or U21844 (N_21844,N_16062,N_17645);
or U21845 (N_21845,N_17202,N_16442);
nor U21846 (N_21846,N_16423,N_16844);
or U21847 (N_21847,N_19068,N_15255);
xnor U21848 (N_21848,N_16573,N_17600);
nand U21849 (N_21849,N_16353,N_15766);
and U21850 (N_21850,N_16646,N_15195);
or U21851 (N_21851,N_15706,N_16398);
or U21852 (N_21852,N_16141,N_17059);
and U21853 (N_21853,N_17891,N_15944);
or U21854 (N_21854,N_19570,N_19796);
or U21855 (N_21855,N_16473,N_15503);
nand U21856 (N_21856,N_16803,N_17142);
and U21857 (N_21857,N_19082,N_19539);
xor U21858 (N_21858,N_19441,N_18219);
nand U21859 (N_21859,N_17104,N_17739);
or U21860 (N_21860,N_17627,N_16151);
and U21861 (N_21861,N_15491,N_17209);
nor U21862 (N_21862,N_16676,N_16693);
nand U21863 (N_21863,N_17860,N_16852);
nor U21864 (N_21864,N_18115,N_15043);
or U21865 (N_21865,N_15922,N_15955);
and U21866 (N_21866,N_15579,N_17120);
nor U21867 (N_21867,N_19623,N_18841);
nor U21868 (N_21868,N_16645,N_16198);
nor U21869 (N_21869,N_16181,N_17609);
and U21870 (N_21870,N_18932,N_18601);
nand U21871 (N_21871,N_17633,N_17344);
nor U21872 (N_21872,N_17778,N_16408);
xor U21873 (N_21873,N_18524,N_18602);
nor U21874 (N_21874,N_15644,N_17617);
nand U21875 (N_21875,N_18587,N_18168);
nand U21876 (N_21876,N_18273,N_15684);
nor U21877 (N_21877,N_16741,N_15203);
and U21878 (N_21878,N_18890,N_16963);
nor U21879 (N_21879,N_18917,N_17708);
nand U21880 (N_21880,N_15643,N_19467);
nand U21881 (N_21881,N_19324,N_16668);
xor U21882 (N_21882,N_15566,N_15064);
and U21883 (N_21883,N_17170,N_19885);
nand U21884 (N_21884,N_19781,N_16391);
nor U21885 (N_21885,N_18993,N_16664);
or U21886 (N_21886,N_18871,N_17729);
xor U21887 (N_21887,N_19457,N_18891);
xnor U21888 (N_21888,N_15375,N_16039);
nor U21889 (N_21889,N_15492,N_16040);
or U21890 (N_21890,N_19268,N_18138);
or U21891 (N_21891,N_15087,N_16695);
nor U21892 (N_21892,N_16255,N_15228);
nand U21893 (N_21893,N_16918,N_19708);
or U21894 (N_21894,N_17041,N_19710);
and U21895 (N_21895,N_17504,N_18944);
nor U21896 (N_21896,N_18288,N_15732);
and U21897 (N_21897,N_17486,N_19316);
nand U21898 (N_21898,N_16051,N_18778);
nor U21899 (N_21899,N_15050,N_17018);
or U21900 (N_21900,N_18591,N_15978);
and U21901 (N_21901,N_15269,N_18372);
or U21902 (N_21902,N_18431,N_17924);
and U21903 (N_21903,N_16496,N_16031);
nor U21904 (N_21904,N_18734,N_19999);
and U21905 (N_21905,N_17123,N_19652);
nand U21906 (N_21906,N_17119,N_17008);
nand U21907 (N_21907,N_15873,N_15568);
xnor U21908 (N_21908,N_15486,N_15712);
and U21909 (N_21909,N_15755,N_19733);
and U21910 (N_21910,N_17067,N_17191);
or U21911 (N_21911,N_19177,N_15749);
nand U21912 (N_21912,N_18748,N_15984);
xor U21913 (N_21913,N_16736,N_18102);
nand U21914 (N_21914,N_15499,N_18370);
nor U21915 (N_21915,N_19173,N_18726);
xnor U21916 (N_21916,N_16708,N_15862);
nor U21917 (N_21917,N_15052,N_19117);
or U21918 (N_21918,N_15820,N_19717);
nand U21919 (N_21919,N_15387,N_19018);
and U21920 (N_21920,N_16571,N_16926);
nor U21921 (N_21921,N_15703,N_15328);
nor U21922 (N_21922,N_17849,N_18412);
and U21923 (N_21923,N_19494,N_19931);
nand U21924 (N_21924,N_18382,N_19102);
or U21925 (N_21925,N_17423,N_18940);
nor U21926 (N_21926,N_19693,N_19080);
nor U21927 (N_21927,N_15266,N_18716);
nor U21928 (N_21928,N_17824,N_18804);
or U21929 (N_21929,N_17922,N_15677);
or U21930 (N_21930,N_19834,N_19606);
nand U21931 (N_21931,N_17651,N_18205);
xor U21932 (N_21932,N_16997,N_19306);
and U21933 (N_21933,N_19670,N_16648);
or U21934 (N_21934,N_16971,N_17629);
xor U21935 (N_21935,N_18574,N_18798);
nor U21936 (N_21936,N_18780,N_15833);
nand U21937 (N_21937,N_16435,N_17298);
and U21938 (N_21938,N_15367,N_18011);
nand U21939 (N_21939,N_19357,N_18072);
nor U21940 (N_21940,N_19145,N_19870);
nor U21941 (N_21941,N_17867,N_19702);
and U21942 (N_21942,N_19774,N_15938);
nand U21943 (N_21943,N_17890,N_19889);
nand U21944 (N_21944,N_16910,N_17889);
xnor U21945 (N_21945,N_16546,N_17985);
xnor U21946 (N_21946,N_16339,N_19629);
nand U21947 (N_21947,N_19657,N_15202);
nor U21948 (N_21948,N_19808,N_18374);
and U21949 (N_21949,N_19504,N_19036);
nor U21950 (N_21950,N_19869,N_18609);
nand U21951 (N_21951,N_19992,N_19191);
and U21952 (N_21952,N_17686,N_19681);
or U21953 (N_21953,N_19127,N_17074);
or U21954 (N_21954,N_19351,N_15789);
and U21955 (N_21955,N_17222,N_18659);
nor U21956 (N_21956,N_17455,N_18700);
and U21957 (N_21957,N_19765,N_17949);
nor U21958 (N_21958,N_16384,N_18833);
or U21959 (N_21959,N_15892,N_17050);
nor U21960 (N_21960,N_19530,N_15742);
nor U21961 (N_21961,N_19372,N_17585);
nor U21962 (N_21962,N_18846,N_19072);
nor U21963 (N_21963,N_18821,N_18339);
nor U21964 (N_21964,N_19071,N_17974);
and U21965 (N_21965,N_15004,N_17404);
and U21966 (N_21966,N_19247,N_16091);
nand U21967 (N_21967,N_15301,N_15399);
xnor U21968 (N_21968,N_15601,N_16032);
xor U21969 (N_21969,N_19898,N_18500);
and U21970 (N_21970,N_17434,N_15247);
and U21971 (N_21971,N_15940,N_15669);
nor U21972 (N_21972,N_19786,N_19825);
or U21973 (N_21973,N_16547,N_16851);
xnor U21974 (N_21974,N_15901,N_18033);
or U21975 (N_21975,N_15091,N_15872);
nand U21976 (N_21976,N_17969,N_17990);
or U21977 (N_21977,N_16903,N_15026);
and U21978 (N_21978,N_18048,N_17053);
and U21979 (N_21979,N_19712,N_15638);
and U21980 (N_21980,N_16924,N_15448);
xnor U21981 (N_21981,N_15148,N_17288);
or U21982 (N_21982,N_15475,N_19551);
or U21983 (N_21983,N_17238,N_19800);
nor U21984 (N_21984,N_16768,N_18233);
nand U21985 (N_21985,N_15540,N_17522);
nand U21986 (N_21986,N_18057,N_18496);
nand U21987 (N_21987,N_15280,N_17931);
nand U21988 (N_21988,N_18446,N_19789);
nand U21989 (N_21989,N_15179,N_15507);
or U21990 (N_21990,N_16643,N_16867);
nand U21991 (N_21991,N_16749,N_19360);
nand U21992 (N_21992,N_16396,N_19239);
or U21993 (N_21993,N_19637,N_17453);
nand U21994 (N_21994,N_17662,N_15778);
or U21995 (N_21995,N_19413,N_17553);
nand U21996 (N_21996,N_15039,N_16267);
nand U21997 (N_21997,N_16277,N_18817);
and U21998 (N_21998,N_19769,N_15784);
or U21999 (N_21999,N_17427,N_18619);
xnor U22000 (N_22000,N_19651,N_15044);
nor U22001 (N_22001,N_15411,N_19864);
and U22002 (N_22002,N_18845,N_16184);
or U22003 (N_22003,N_19561,N_16283);
and U22004 (N_22004,N_16783,N_19732);
nor U22005 (N_22005,N_17263,N_15014);
and U22006 (N_22006,N_15626,N_19662);
nor U22007 (N_22007,N_16452,N_15219);
and U22008 (N_22008,N_15451,N_17452);
nor U22009 (N_22009,N_19368,N_16543);
or U22010 (N_22010,N_17264,N_18625);
nand U22011 (N_22011,N_17019,N_17709);
or U22012 (N_22012,N_16357,N_15726);
nor U22013 (N_22013,N_19271,N_19215);
nor U22014 (N_22014,N_18667,N_16116);
or U22015 (N_22015,N_16367,N_17875);
and U22016 (N_22016,N_18870,N_18918);
nor U22017 (N_22017,N_19761,N_18519);
or U22018 (N_22018,N_16117,N_16972);
xor U22019 (N_22019,N_19705,N_18577);
nand U22020 (N_22020,N_15737,N_15610);
or U22021 (N_22021,N_19612,N_15306);
nand U22022 (N_22022,N_18760,N_19565);
and U22023 (N_22023,N_16047,N_19428);
and U22024 (N_22024,N_19540,N_18049);
and U22025 (N_22025,N_15815,N_16592);
nand U22026 (N_22026,N_17623,N_18942);
nand U22027 (N_22027,N_18054,N_18643);
nand U22028 (N_22028,N_17598,N_15884);
or U22029 (N_22029,N_16866,N_17488);
nor U22030 (N_22030,N_19969,N_17564);
or U22031 (N_22031,N_17078,N_18834);
nand U22032 (N_22032,N_18310,N_18575);
xor U22033 (N_22033,N_18375,N_19996);
and U22034 (N_22034,N_17044,N_16719);
nor U22035 (N_22035,N_19403,N_19275);
or U22036 (N_22036,N_17711,N_17429);
or U22037 (N_22037,N_16079,N_15355);
and U22038 (N_22038,N_15127,N_15386);
xor U22039 (N_22039,N_19649,N_18124);
nand U22040 (N_22040,N_18463,N_19197);
or U22041 (N_22041,N_16516,N_17563);
nand U22042 (N_22042,N_18089,N_19678);
nand U22043 (N_22043,N_16340,N_17952);
xor U22044 (N_22044,N_18553,N_15285);
nor U22045 (N_22045,N_17223,N_15335);
nor U22046 (N_22046,N_17869,N_17816);
nand U22047 (N_22047,N_15577,N_18203);
and U22048 (N_22048,N_18779,N_17072);
nor U22049 (N_22049,N_16245,N_17342);
nand U22050 (N_22050,N_17877,N_17150);
and U22051 (N_22051,N_16063,N_16463);
nand U22052 (N_22052,N_19593,N_17743);
nand U22053 (N_22053,N_19355,N_18985);
nand U22054 (N_22054,N_17199,N_18135);
and U22055 (N_22055,N_18805,N_18717);
nor U22056 (N_22056,N_17077,N_19435);
and U22057 (N_22057,N_16914,N_17208);
or U22058 (N_22058,N_17900,N_16156);
or U22059 (N_22059,N_15986,N_18514);
nor U22060 (N_22060,N_18277,N_19408);
nor U22061 (N_22061,N_18467,N_16680);
and U22062 (N_22062,N_18636,N_15057);
nor U22063 (N_22063,N_16162,N_18126);
and U22064 (N_22064,N_18289,N_17959);
nor U22065 (N_22065,N_16269,N_18349);
or U22066 (N_22066,N_15554,N_19986);
nand U22067 (N_22067,N_19768,N_17198);
and U22068 (N_22068,N_18269,N_18851);
and U22069 (N_22069,N_18260,N_15291);
nand U22070 (N_22070,N_17010,N_18035);
and U22071 (N_22071,N_17324,N_17581);
or U22072 (N_22072,N_18866,N_19667);
or U22073 (N_22073,N_15746,N_19010);
and U22074 (N_22074,N_18380,N_15997);
and U22075 (N_22075,N_16921,N_16237);
and U22076 (N_22076,N_17064,N_17013);
and U22077 (N_22077,N_15589,N_17671);
nor U22078 (N_22078,N_19167,N_16100);
or U22079 (N_22079,N_16002,N_15133);
or U22080 (N_22080,N_17559,N_18364);
nand U22081 (N_22081,N_17776,N_15304);
nand U22082 (N_22082,N_15141,N_17194);
and U22083 (N_22083,N_17471,N_16412);
nand U22084 (N_22084,N_16146,N_17561);
or U22085 (N_22085,N_15350,N_17054);
xnor U22086 (N_22086,N_15813,N_15351);
or U22087 (N_22087,N_15893,N_17063);
nor U22088 (N_22088,N_17474,N_19918);
or U22089 (N_22089,N_15788,N_18732);
xor U22090 (N_22090,N_17231,N_15911);
or U22091 (N_22091,N_16937,N_15019);
or U22092 (N_22092,N_17165,N_18291);
xnor U22093 (N_22093,N_17926,N_19486);
or U22094 (N_22094,N_18559,N_18513);
nor U22095 (N_22095,N_17936,N_17531);
nor U22096 (N_22096,N_15704,N_16000);
nand U22097 (N_22097,N_17665,N_17759);
nand U22098 (N_22098,N_17970,N_15240);
nor U22099 (N_22099,N_18642,N_17616);
nand U22100 (N_22100,N_16246,N_19600);
or U22101 (N_22101,N_16123,N_15769);
nand U22102 (N_22102,N_16143,N_18231);
xor U22103 (N_22103,N_16241,N_17107);
nor U22104 (N_22104,N_19361,N_16254);
nor U22105 (N_22105,N_18595,N_18028);
and U22106 (N_22106,N_17897,N_19092);
or U22107 (N_22107,N_18067,N_19779);
or U22108 (N_22108,N_17201,N_15377);
and U22109 (N_22109,N_16057,N_19465);
xor U22110 (N_22110,N_17537,N_19074);
or U22111 (N_22111,N_18488,N_15981);
and U22112 (N_22112,N_18850,N_15437);
or U22113 (N_22113,N_16800,N_15680);
or U22114 (N_22114,N_16548,N_17160);
nor U22115 (N_22115,N_18970,N_15175);
nand U22116 (N_22116,N_15326,N_17417);
nor U22117 (N_22117,N_17431,N_15509);
and U22118 (N_22118,N_18832,N_16681);
xnor U22119 (N_22119,N_16760,N_17145);
or U22120 (N_22120,N_15413,N_18286);
nand U22121 (N_22121,N_16711,N_16786);
nand U22122 (N_22122,N_15534,N_15180);
and U22123 (N_22123,N_17707,N_15759);
nand U22124 (N_22124,N_19056,N_16466);
nand U22125 (N_22125,N_19698,N_17595);
and U22126 (N_22126,N_16182,N_19123);
nor U22127 (N_22127,N_16657,N_19823);
nor U22128 (N_22128,N_15174,N_15508);
or U22129 (N_22129,N_16519,N_17693);
and U22130 (N_22130,N_16324,N_19729);
nand U22131 (N_22131,N_17821,N_19522);
and U22132 (N_22132,N_18787,N_16049);
nand U22133 (N_22133,N_17810,N_17408);
or U22134 (N_22134,N_15007,N_19161);
or U22135 (N_22135,N_16380,N_19314);
or U22136 (N_22136,N_19811,N_18041);
nand U22137 (N_22137,N_18143,N_17864);
or U22138 (N_22138,N_15028,N_15762);
or U22139 (N_22139,N_17076,N_18725);
xor U22140 (N_22140,N_18400,N_18910);
nor U22141 (N_22141,N_17001,N_19411);
nand U22142 (N_22142,N_18458,N_18958);
nor U22143 (N_22143,N_16197,N_16395);
nor U22144 (N_22144,N_18566,N_19739);
nand U22145 (N_22145,N_19382,N_18239);
or U22146 (N_22146,N_18405,N_17358);
nand U22147 (N_22147,N_15916,N_18474);
xnor U22148 (N_22148,N_16114,N_18572);
nand U22149 (N_22149,N_19973,N_15886);
nor U22150 (N_22150,N_19602,N_18959);
xnor U22151 (N_22151,N_19052,N_17611);
nor U22152 (N_22152,N_16188,N_18650);
or U22153 (N_22153,N_16689,N_15153);
nand U22154 (N_22154,N_15071,N_16700);
xnor U22155 (N_22155,N_18290,N_15714);
or U22156 (N_22156,N_19943,N_15942);
and U22157 (N_22157,N_15621,N_16675);
nor U22158 (N_22158,N_16631,N_17892);
nand U22159 (N_22159,N_17339,N_16004);
and U22160 (N_22160,N_17811,N_16821);
xor U22161 (N_22161,N_18263,N_17779);
nand U22162 (N_22162,N_19347,N_17215);
nor U22163 (N_22163,N_17642,N_15308);
nor U22164 (N_22164,N_18881,N_19492);
and U22165 (N_22165,N_16397,N_17786);
nand U22166 (N_22166,N_16779,N_19259);
nand U22167 (N_22167,N_16060,N_15548);
nand U22168 (N_22168,N_15259,N_15937);
and U22169 (N_22169,N_16122,N_19333);
or U22170 (N_22170,N_17903,N_19566);
nand U22171 (N_22171,N_16139,N_19103);
nand U22172 (N_22172,N_16873,N_19782);
nand U22173 (N_22173,N_15059,N_16427);
nor U22174 (N_22174,N_15654,N_17909);
and U22175 (N_22175,N_18931,N_15119);
nand U22176 (N_22176,N_18147,N_19442);
xnor U22177 (N_22177,N_16782,N_19856);
or U22178 (N_22178,N_19026,N_15629);
xor U22179 (N_22179,N_17797,N_15800);
and U22180 (N_22180,N_16912,N_19814);
nand U22181 (N_22181,N_16616,N_16687);
xor U22182 (N_22182,N_16770,N_16309);
nand U22183 (N_22183,N_17538,N_15101);
nor U22184 (N_22184,N_18543,N_17256);
and U22185 (N_22185,N_15538,N_17236);
nand U22186 (N_22186,N_17732,N_17780);
and U22187 (N_22187,N_17381,N_17666);
and U22188 (N_22188,N_17375,N_17332);
nand U22189 (N_22189,N_16089,N_15907);
nor U22190 (N_22190,N_16625,N_16185);
nand U22191 (N_22191,N_16304,N_16428);
and U22192 (N_22192,N_15757,N_15463);
and U22193 (N_22193,N_19621,N_19881);
nand U22194 (N_22194,N_16112,N_17986);
xnor U22195 (N_22195,N_15775,N_16717);
nand U22196 (N_22196,N_17062,N_17272);
and U22197 (N_22197,N_19751,N_16319);
and U22198 (N_22198,N_16641,N_19756);
xnor U22199 (N_22199,N_19804,N_17475);
nand U22200 (N_22200,N_16961,N_18141);
or U22201 (N_22201,N_17033,N_17953);
and U22202 (N_22202,N_19209,N_16095);
or U22203 (N_22203,N_15773,N_16366);
and U22204 (N_22204,N_17258,N_17140);
nor U22205 (N_22205,N_15628,N_17122);
nor U22206 (N_22206,N_15201,N_19097);
and U22207 (N_22207,N_17543,N_18765);
xor U22208 (N_22208,N_18681,N_16356);
xnor U22209 (N_22209,N_19459,N_16234);
nor U22210 (N_22210,N_15622,N_16842);
xor U22211 (N_22211,N_19341,N_16870);
nor U22212 (N_22212,N_15848,N_15519);
xnor U22213 (N_22213,N_16970,N_18294);
nor U22214 (N_22214,N_16953,N_19236);
and U22215 (N_22215,N_18186,N_15739);
and U22216 (N_22216,N_16977,N_19849);
xor U22217 (N_22217,N_16766,N_17383);
nor U22218 (N_22218,N_19399,N_16211);
or U22219 (N_22219,N_17755,N_19349);
or U22220 (N_22220,N_16297,N_18119);
nor U22221 (N_22221,N_18155,N_19666);
and U22222 (N_22222,N_15660,N_15701);
nand U22223 (N_22223,N_19616,N_18556);
and U22224 (N_22224,N_17650,N_18353);
or U22225 (N_22225,N_18006,N_15181);
nor U22226 (N_22226,N_17549,N_15998);
or U22227 (N_22227,N_15576,N_16904);
nor U22228 (N_22228,N_15258,N_16637);
or U22229 (N_22229,N_18130,N_15965);
nor U22230 (N_22230,N_15875,N_16658);
nand U22231 (N_22231,N_17430,N_16998);
nand U22232 (N_22232,N_15840,N_15173);
or U22233 (N_22233,N_18953,N_16128);
nor U22234 (N_22234,N_16607,N_16845);
nor U22235 (N_22235,N_17672,N_18893);
or U22236 (N_22236,N_17731,N_17697);
nand U22237 (N_22237,N_18816,N_16727);
and U22238 (N_22238,N_19576,N_16213);
nor U22239 (N_22239,N_18251,N_18322);
nand U22240 (N_22240,N_19422,N_18428);
xor U22241 (N_22241,N_15244,N_19410);
and U22242 (N_22242,N_18853,N_15256);
xnor U22243 (N_22243,N_17345,N_17748);
or U22244 (N_22244,N_17346,N_19024);
nor U22245 (N_22245,N_17132,N_16351);
nand U22246 (N_22246,N_16437,N_16580);
nand U22247 (N_22247,N_15382,N_18456);
nor U22248 (N_22248,N_19238,N_19216);
and U22249 (N_22249,N_18530,N_18903);
or U22250 (N_22250,N_18211,N_18783);
or U22251 (N_22251,N_18455,N_19741);
nor U22252 (N_22252,N_19343,N_17540);
nand U22253 (N_22253,N_19231,N_18266);
xnor U22254 (N_22254,N_15952,N_16362);
or U22255 (N_22255,N_17071,N_17977);
nand U22256 (N_22256,N_18688,N_16424);
nor U22257 (N_22257,N_16405,N_19454);
or U22258 (N_22258,N_18333,N_18707);
xnor U22259 (N_22259,N_17377,N_15754);
and U22260 (N_22260,N_19151,N_18042);
and U22261 (N_22261,N_16462,N_19105);
or U22262 (N_22262,N_17844,N_17569);
and U22263 (N_22263,N_18324,N_19185);
or U22264 (N_22264,N_19598,N_18101);
nor U22265 (N_22265,N_18499,N_16816);
and U22266 (N_22266,N_15470,N_15504);
nand U22267 (N_22267,N_19802,N_16078);
nor U22268 (N_22268,N_19747,N_16347);
nand U22269 (N_22269,N_19497,N_15526);
and U22270 (N_22270,N_16212,N_18568);
nand U22271 (N_22271,N_17917,N_18334);
nand U22272 (N_22272,N_17316,N_17565);
xnor U22273 (N_22273,N_18315,N_18924);
nand U22274 (N_22274,N_15434,N_19989);
or U22275 (N_22275,N_18014,N_15025);
and U22276 (N_22276,N_16099,N_15694);
nand U22277 (N_22277,N_17412,N_19579);
nand U22278 (N_22278,N_19178,N_17591);
or U22279 (N_22279,N_19942,N_17691);
or U22280 (N_22280,N_15641,N_17520);
nand U22281 (N_22281,N_17061,N_16090);
xor U22282 (N_22282,N_18237,N_19432);
or U22283 (N_22283,N_16893,N_17517);
and U22284 (N_22284,N_15632,N_16103);
and U22285 (N_22285,N_19266,N_15347);
nand U22286 (N_22286,N_18672,N_16855);
nor U22287 (N_22287,N_17735,N_17219);
xnor U22288 (N_22288,N_16291,N_19735);
or U22289 (N_22289,N_18825,N_19302);
nand U22290 (N_22290,N_16712,N_19574);
nor U22291 (N_22291,N_18199,N_18887);
nand U22292 (N_22292,N_18025,N_17220);
or U22293 (N_22293,N_18355,N_17966);
and U22294 (N_22294,N_18943,N_15476);
nand U22295 (N_22295,N_18536,N_17934);
nand U22296 (N_22296,N_18470,N_16906);
and U22297 (N_22297,N_16107,N_15549);
nor U22298 (N_22298,N_16012,N_18477);
nor U22299 (N_22299,N_16841,N_18045);
and U22300 (N_22300,N_15082,N_18806);
xnor U22301 (N_22301,N_15897,N_19868);
nor U22302 (N_22302,N_17512,N_17698);
or U22303 (N_22303,N_15561,N_15342);
or U22304 (N_22304,N_16859,N_15160);
nand U22305 (N_22305,N_19130,N_16230);
xnor U22306 (N_22306,N_19429,N_15237);
and U22307 (N_22307,N_18140,N_19427);
and U22308 (N_22308,N_18082,N_19013);
xor U22309 (N_22309,N_19878,N_18379);
and U22310 (N_22310,N_16531,N_15422);
nand U22311 (N_22311,N_17946,N_18005);
xnor U22312 (N_22312,N_15449,N_16720);
nand U22313 (N_22313,N_15390,N_15292);
nor U22314 (N_22314,N_19668,N_15473);
and U22315 (N_22315,N_19605,N_16310);
xnor U22316 (N_22316,N_19256,N_15505);
xnor U22317 (N_22317,N_18032,N_15322);
nand U22318 (N_22318,N_18064,N_17607);
and U22319 (N_22319,N_16265,N_19113);
nor U22320 (N_22320,N_15645,N_16986);
or U22321 (N_22321,N_16621,N_16135);
or U22322 (N_22322,N_19792,N_15930);
and U22323 (N_22323,N_17265,N_16382);
nor U22324 (N_22324,N_16417,N_15040);
nand U22325 (N_22325,N_19133,N_16257);
and U22326 (N_22326,N_17871,N_16243);
and U22327 (N_22327,N_18907,N_17360);
nor U22328 (N_22328,N_18282,N_16102);
xor U22329 (N_22329,N_16132,N_17976);
and U22330 (N_22330,N_16525,N_16312);
and U22331 (N_22331,N_19935,N_17046);
or U22332 (N_22332,N_15582,N_15770);
nor U22333 (N_22333,N_16176,N_19132);
or U22334 (N_22334,N_15810,N_19818);
or U22335 (N_22335,N_16560,N_17847);
nand U22336 (N_22336,N_19495,N_15874);
nand U22337 (N_22337,N_19012,N_16450);
and U22338 (N_22338,N_17290,N_15281);
and U22339 (N_22339,N_16557,N_17989);
or U22340 (N_22340,N_19290,N_17935);
nand U22341 (N_22341,N_18256,N_16223);
nand U22342 (N_22342,N_18824,N_17424);
nand U22343 (N_22343,N_16272,N_19008);
nor U22344 (N_22344,N_19400,N_18226);
nor U22345 (N_22345,N_17842,N_16383);
nand U22346 (N_22346,N_15218,N_19809);
xor U22347 (N_22347,N_18230,N_18232);
nor U22348 (N_22348,N_18091,N_16581);
xor U22349 (N_22349,N_15510,N_16205);
xnor U22350 (N_22350,N_16350,N_17070);
nor U22351 (N_22351,N_18433,N_19199);
nor U22352 (N_22352,N_19004,N_15140);
nor U22353 (N_22353,N_19118,N_19845);
nand U22354 (N_22354,N_17057,N_17809);
or U22355 (N_22355,N_16840,N_19136);
or U22356 (N_22356,N_16098,N_16701);
or U22357 (N_22357,N_19243,N_16978);
nand U22358 (N_22358,N_15116,N_18752);
and U22359 (N_22359,N_17961,N_18984);
and U22360 (N_22360,N_17301,N_19533);
or U22361 (N_22361,N_18627,N_16964);
or U22362 (N_22362,N_15105,N_19146);
nor U22363 (N_22363,N_19493,N_16639);
xnor U22364 (N_22364,N_19586,N_17242);
and U22365 (N_22365,N_18395,N_15616);
or U22366 (N_22366,N_18154,N_18332);
or U22367 (N_22367,N_15962,N_15048);
nand U22368 (N_22368,N_18451,N_15117);
nand U22369 (N_22369,N_17873,N_16227);
and U22370 (N_22370,N_19169,N_18099);
or U22371 (N_22371,N_19923,N_16679);
and U22372 (N_22372,N_17620,N_19365);
and U22373 (N_22373,N_16504,N_17438);
and U22374 (N_22374,N_19661,N_16959);
nor U22375 (N_22375,N_15674,N_18051);
or U22376 (N_22376,N_18703,N_16404);
nand U22377 (N_22377,N_18009,N_16652);
nand U22378 (N_22378,N_18502,N_19628);
or U22379 (N_22379,N_17135,N_18223);
xnor U22380 (N_22380,N_18620,N_18662);
xor U22381 (N_22381,N_18520,N_18646);
nand U22382 (N_22382,N_19001,N_18904);
or U22383 (N_22383,N_15324,N_18879);
and U22384 (N_22384,N_17659,N_19597);
and U22385 (N_22385,N_19871,N_19212);
nand U22386 (N_22386,N_16216,N_17167);
nor U22387 (N_22387,N_15595,N_15261);
nor U22388 (N_22388,N_17456,N_18737);
nor U22389 (N_22389,N_19620,N_15879);
nand U22390 (N_22390,N_17441,N_15441);
nand U22391 (N_22391,N_15881,N_15100);
nor U22392 (N_22392,N_15378,N_18132);
or U22393 (N_22393,N_16441,N_18090);
and U22394 (N_22394,N_18254,N_16732);
xor U22395 (N_22395,N_17021,N_18425);
or U22396 (N_22396,N_15442,N_18225);
or U22397 (N_22397,N_18070,N_18495);
and U22398 (N_22398,N_16696,N_16608);
nand U22399 (N_22399,N_19471,N_15569);
nand U22400 (N_22400,N_19201,N_19106);
nor U22401 (N_22401,N_19909,N_17087);
nand U22402 (N_22402,N_19591,N_18792);
nand U22403 (N_22403,N_19404,N_15969);
or U22404 (N_22404,N_17204,N_16043);
nor U22405 (N_22405,N_17541,N_18763);
nor U22406 (N_22406,N_19320,N_17898);
nor U22407 (N_22407,N_16941,N_18453);
and U22408 (N_22408,N_19407,N_15580);
nor U22409 (N_22409,N_17390,N_17338);
nor U22410 (N_22410,N_18162,N_17933);
nor U22411 (N_22411,N_18802,N_16662);
nand U22412 (N_22412,N_15906,N_17113);
nand U22413 (N_22413,N_17225,N_17722);
xor U22414 (N_22414,N_16485,N_16503);
nand U22415 (N_22415,N_19884,N_17521);
nor U22416 (N_22416,N_17355,N_18693);
and U22417 (N_22417,N_18750,N_18558);
or U22418 (N_22418,N_17765,N_19980);
nand U22419 (N_22419,N_16869,N_17260);
nor U22420 (N_22420,N_18666,N_19420);
or U22421 (N_22421,N_19077,N_19937);
and U22422 (N_22422,N_17166,N_16614);
nor U22423 (N_22423,N_15300,N_17035);
nor U22424 (N_22424,N_19214,N_15847);
and U22425 (N_22425,N_19737,N_16476);
or U22426 (N_22426,N_15729,N_19738);
xor U22427 (N_22427,N_19567,N_16533);
xnor U22428 (N_22428,N_16569,N_15129);
or U22429 (N_22429,N_16638,N_16922);
nand U22430 (N_22430,N_16931,N_17395);
or U22431 (N_22431,N_17758,N_16774);
and U22432 (N_22432,N_16420,N_16626);
or U22433 (N_22433,N_15110,N_18383);
nand U22434 (N_22434,N_15363,N_17567);
or U22435 (N_22435,N_18087,N_18847);
nor U22436 (N_22436,N_16545,N_17830);
or U22437 (N_22437,N_18019,N_16287);
and U22438 (N_22438,N_19924,N_15452);
nor U22439 (N_22439,N_19086,N_18652);
nor U22440 (N_22440,N_15284,N_15410);
nor U22441 (N_22441,N_17413,N_19844);
nand U22442 (N_22442,N_18983,N_16378);
xnor U22443 (N_22443,N_16594,N_19307);
nand U22444 (N_22444,N_18483,N_18705);
or U22445 (N_22445,N_16262,N_17907);
or U22446 (N_22446,N_15053,N_15910);
nor U22447 (N_22447,N_18812,N_17162);
or U22448 (N_22448,N_18579,N_15132);
and U22449 (N_22449,N_17716,N_15740);
nor U22450 (N_22450,N_17655,N_18583);
or U22451 (N_22451,N_15432,N_19203);
or U22452 (N_22452,N_15604,N_16179);
nor U22453 (N_22453,N_18923,N_18517);
and U22454 (N_22454,N_17396,N_15407);
nand U22455 (N_22455,N_16747,N_18831);
nor U22456 (N_22456,N_17172,N_17688);
nand U22457 (N_22457,N_17937,N_19833);
nor U22458 (N_22458,N_16755,N_19812);
or U22459 (N_22459,N_17468,N_15705);
nand U22460 (N_22460,N_17446,N_17147);
and U22461 (N_22461,N_19528,N_17532);
and U22462 (N_22462,N_16865,N_16858);
or U22463 (N_22463,N_15806,N_17161);
and U22464 (N_22464,N_19525,N_16486);
or U22465 (N_22465,N_18573,N_19340);
and U22466 (N_22466,N_18359,N_15817);
and U22467 (N_22467,N_19211,N_15230);
or U22468 (N_22468,N_16274,N_16916);
and U22469 (N_22469,N_18746,N_18534);
and U22470 (N_22470,N_16250,N_18055);
and U22471 (N_22471,N_16118,N_16306);
nor U22472 (N_22472,N_19139,N_18276);
or U22473 (N_22473,N_19982,N_19894);
nand U22474 (N_22474,N_16656,N_19558);
or U22475 (N_22475,N_16474,N_18439);
nand U22476 (N_22476,N_17411,N_17116);
or U22477 (N_22477,N_19264,N_16674);
nand U22478 (N_22478,N_18977,N_16798);
nand U22479 (N_22479,N_19083,N_15678);
or U22480 (N_22480,N_19122,N_17351);
and U22481 (N_22481,N_16373,N_18018);
nor U22482 (N_22482,N_19813,N_16752);
nor U22483 (N_22483,N_18358,N_15161);
or U22484 (N_22484,N_17835,N_16833);
nor U22485 (N_22485,N_15115,N_19965);
nor U22486 (N_22486,N_17228,N_19948);
nand U22487 (N_22487,N_19679,N_16748);
or U22488 (N_22488,N_17206,N_16555);
and U22489 (N_22489,N_19615,N_17128);
nand U22490 (N_22490,N_19142,N_16050);
or U22491 (N_22491,N_18287,N_15222);
nor U22492 (N_22492,N_19150,N_18131);
or U22493 (N_22493,N_19027,N_19699);
and U22494 (N_22494,N_17397,N_18476);
or U22495 (N_22495,N_18274,N_18228);
and U22496 (N_22496,N_17680,N_19622);
or U22497 (N_22497,N_16723,N_17178);
or U22498 (N_22498,N_19129,N_16698);
nor U22499 (N_22499,N_19902,N_17654);
nand U22500 (N_22500,N_16657,N_16421);
nand U22501 (N_22501,N_17017,N_16066);
or U22502 (N_22502,N_19465,N_16920);
xor U22503 (N_22503,N_18332,N_16259);
or U22504 (N_22504,N_16865,N_16860);
nor U22505 (N_22505,N_19960,N_18045);
nor U22506 (N_22506,N_16973,N_15628);
and U22507 (N_22507,N_15071,N_17637);
nand U22508 (N_22508,N_19425,N_19327);
or U22509 (N_22509,N_18397,N_18561);
xor U22510 (N_22510,N_18006,N_17911);
and U22511 (N_22511,N_18159,N_17012);
and U22512 (N_22512,N_16751,N_15964);
and U22513 (N_22513,N_18966,N_19138);
nor U22514 (N_22514,N_19222,N_17048);
or U22515 (N_22515,N_18446,N_17286);
or U22516 (N_22516,N_17395,N_15795);
and U22517 (N_22517,N_15316,N_18572);
and U22518 (N_22518,N_19418,N_17874);
nor U22519 (N_22519,N_18450,N_16068);
nand U22520 (N_22520,N_16383,N_15809);
or U22521 (N_22521,N_17068,N_18717);
xnor U22522 (N_22522,N_17870,N_18259);
xnor U22523 (N_22523,N_16351,N_18446);
nor U22524 (N_22524,N_16791,N_15441);
nand U22525 (N_22525,N_17053,N_18325);
nor U22526 (N_22526,N_15200,N_19694);
nand U22527 (N_22527,N_19556,N_18361);
xor U22528 (N_22528,N_17465,N_19905);
nand U22529 (N_22529,N_15851,N_19963);
or U22530 (N_22530,N_16961,N_18054);
nand U22531 (N_22531,N_18357,N_16481);
nand U22532 (N_22532,N_17637,N_19311);
xor U22533 (N_22533,N_17693,N_17876);
or U22534 (N_22534,N_17247,N_15406);
nand U22535 (N_22535,N_19607,N_15024);
or U22536 (N_22536,N_18058,N_18513);
and U22537 (N_22537,N_17082,N_15227);
nand U22538 (N_22538,N_18610,N_17336);
xor U22539 (N_22539,N_17923,N_18847);
nor U22540 (N_22540,N_19197,N_16167);
xnor U22541 (N_22541,N_17195,N_19149);
and U22542 (N_22542,N_15406,N_17773);
and U22543 (N_22543,N_19308,N_19440);
xor U22544 (N_22544,N_15738,N_17838);
xnor U22545 (N_22545,N_17590,N_15985);
nor U22546 (N_22546,N_18237,N_17311);
or U22547 (N_22547,N_18347,N_18933);
nor U22548 (N_22548,N_18787,N_18463);
nor U22549 (N_22549,N_16165,N_15380);
and U22550 (N_22550,N_17468,N_19813);
or U22551 (N_22551,N_18350,N_19281);
and U22552 (N_22552,N_15983,N_17367);
or U22553 (N_22553,N_18441,N_19176);
or U22554 (N_22554,N_15272,N_19264);
nand U22555 (N_22555,N_17149,N_17883);
or U22556 (N_22556,N_16104,N_19677);
and U22557 (N_22557,N_19596,N_17035);
nor U22558 (N_22558,N_18045,N_16090);
nor U22559 (N_22559,N_18226,N_18194);
and U22560 (N_22560,N_19294,N_19435);
nor U22561 (N_22561,N_15231,N_17702);
xnor U22562 (N_22562,N_18614,N_18828);
nand U22563 (N_22563,N_17000,N_16805);
nand U22564 (N_22564,N_15467,N_18085);
or U22565 (N_22565,N_18320,N_16008);
nand U22566 (N_22566,N_15801,N_16953);
or U22567 (N_22567,N_19959,N_19240);
nor U22568 (N_22568,N_19710,N_19774);
or U22569 (N_22569,N_18928,N_18288);
nand U22570 (N_22570,N_15182,N_17899);
nor U22571 (N_22571,N_17982,N_15468);
nor U22572 (N_22572,N_19952,N_18179);
and U22573 (N_22573,N_15617,N_16147);
nand U22574 (N_22574,N_15847,N_19400);
and U22575 (N_22575,N_19065,N_19140);
nor U22576 (N_22576,N_18879,N_16571);
and U22577 (N_22577,N_17514,N_19167);
nand U22578 (N_22578,N_18769,N_16576);
nand U22579 (N_22579,N_17292,N_17096);
xor U22580 (N_22580,N_16123,N_19134);
nand U22581 (N_22581,N_16536,N_18958);
xnor U22582 (N_22582,N_16184,N_18439);
nand U22583 (N_22583,N_19457,N_15424);
or U22584 (N_22584,N_16518,N_17209);
or U22585 (N_22585,N_16642,N_17813);
xor U22586 (N_22586,N_15111,N_17613);
and U22587 (N_22587,N_19747,N_17783);
nand U22588 (N_22588,N_16939,N_18624);
and U22589 (N_22589,N_15713,N_15430);
or U22590 (N_22590,N_17276,N_18803);
and U22591 (N_22591,N_19762,N_18151);
nand U22592 (N_22592,N_19600,N_16544);
xnor U22593 (N_22593,N_15330,N_17809);
nor U22594 (N_22594,N_17784,N_17190);
or U22595 (N_22595,N_16126,N_15277);
xnor U22596 (N_22596,N_16031,N_16032);
nor U22597 (N_22597,N_19199,N_18234);
nand U22598 (N_22598,N_19608,N_18060);
and U22599 (N_22599,N_18791,N_15806);
and U22600 (N_22600,N_16263,N_16654);
nand U22601 (N_22601,N_17653,N_18715);
and U22602 (N_22602,N_19664,N_15761);
nand U22603 (N_22603,N_19596,N_16399);
nor U22604 (N_22604,N_15021,N_19186);
nand U22605 (N_22605,N_18004,N_16500);
xnor U22606 (N_22606,N_15836,N_19885);
nand U22607 (N_22607,N_19705,N_17550);
or U22608 (N_22608,N_16788,N_16850);
and U22609 (N_22609,N_16124,N_15824);
nand U22610 (N_22610,N_16701,N_15244);
nor U22611 (N_22611,N_17972,N_16827);
nand U22612 (N_22612,N_17639,N_16831);
nand U22613 (N_22613,N_15469,N_19736);
nor U22614 (N_22614,N_16108,N_17048);
or U22615 (N_22615,N_18368,N_18902);
and U22616 (N_22616,N_19248,N_15097);
and U22617 (N_22617,N_16430,N_17012);
and U22618 (N_22618,N_16065,N_16883);
nand U22619 (N_22619,N_16665,N_15546);
or U22620 (N_22620,N_19382,N_17468);
and U22621 (N_22621,N_15671,N_17343);
and U22622 (N_22622,N_17842,N_17952);
xor U22623 (N_22623,N_17225,N_16673);
and U22624 (N_22624,N_19437,N_17793);
nand U22625 (N_22625,N_19504,N_18084);
nor U22626 (N_22626,N_16310,N_16413);
nand U22627 (N_22627,N_15132,N_16887);
or U22628 (N_22628,N_17914,N_17491);
or U22629 (N_22629,N_17188,N_16998);
xnor U22630 (N_22630,N_19361,N_16746);
nor U22631 (N_22631,N_18360,N_19871);
or U22632 (N_22632,N_17953,N_16554);
or U22633 (N_22633,N_18174,N_17515);
nand U22634 (N_22634,N_15424,N_15841);
and U22635 (N_22635,N_16220,N_16477);
nand U22636 (N_22636,N_19355,N_16118);
nand U22637 (N_22637,N_16334,N_18122);
nor U22638 (N_22638,N_17626,N_17027);
nand U22639 (N_22639,N_19547,N_16426);
nand U22640 (N_22640,N_15648,N_16096);
nor U22641 (N_22641,N_19142,N_19811);
and U22642 (N_22642,N_15590,N_15003);
and U22643 (N_22643,N_15432,N_19250);
xnor U22644 (N_22644,N_15676,N_17148);
or U22645 (N_22645,N_16076,N_18349);
nand U22646 (N_22646,N_18914,N_17795);
and U22647 (N_22647,N_15618,N_19584);
or U22648 (N_22648,N_16030,N_15892);
or U22649 (N_22649,N_18328,N_19760);
and U22650 (N_22650,N_15893,N_18478);
nor U22651 (N_22651,N_19389,N_17185);
nand U22652 (N_22652,N_16924,N_16420);
or U22653 (N_22653,N_19756,N_19809);
or U22654 (N_22654,N_15111,N_16111);
or U22655 (N_22655,N_19643,N_15842);
or U22656 (N_22656,N_18495,N_16882);
or U22657 (N_22657,N_18367,N_17977);
or U22658 (N_22658,N_17907,N_18788);
or U22659 (N_22659,N_16234,N_17950);
nand U22660 (N_22660,N_17168,N_15295);
and U22661 (N_22661,N_18598,N_18529);
or U22662 (N_22662,N_17808,N_15104);
and U22663 (N_22663,N_16082,N_19679);
nand U22664 (N_22664,N_15592,N_17103);
or U22665 (N_22665,N_17165,N_19997);
nand U22666 (N_22666,N_17217,N_16310);
or U22667 (N_22667,N_19492,N_16184);
xnor U22668 (N_22668,N_16780,N_18865);
and U22669 (N_22669,N_16152,N_18916);
nand U22670 (N_22670,N_16244,N_19778);
nor U22671 (N_22671,N_18154,N_19069);
and U22672 (N_22672,N_17013,N_15183);
and U22673 (N_22673,N_15913,N_18082);
nor U22674 (N_22674,N_16561,N_15249);
xnor U22675 (N_22675,N_18685,N_19465);
nor U22676 (N_22676,N_17113,N_16056);
xnor U22677 (N_22677,N_17383,N_19157);
nor U22678 (N_22678,N_16608,N_18450);
and U22679 (N_22679,N_18540,N_15892);
or U22680 (N_22680,N_15177,N_16453);
or U22681 (N_22681,N_19320,N_18389);
nor U22682 (N_22682,N_19275,N_19490);
nor U22683 (N_22683,N_17489,N_18792);
or U22684 (N_22684,N_16580,N_19134);
nor U22685 (N_22685,N_16519,N_17153);
nor U22686 (N_22686,N_19055,N_16251);
nand U22687 (N_22687,N_15676,N_17717);
nand U22688 (N_22688,N_18269,N_17818);
nand U22689 (N_22689,N_16011,N_19258);
nor U22690 (N_22690,N_17194,N_17032);
nand U22691 (N_22691,N_19753,N_18217);
nand U22692 (N_22692,N_15675,N_16919);
and U22693 (N_22693,N_17929,N_16378);
xnor U22694 (N_22694,N_19397,N_16430);
nor U22695 (N_22695,N_15891,N_15453);
and U22696 (N_22696,N_18802,N_15150);
nand U22697 (N_22697,N_16916,N_16299);
and U22698 (N_22698,N_15511,N_19332);
nand U22699 (N_22699,N_16932,N_17669);
nand U22700 (N_22700,N_16182,N_17548);
nor U22701 (N_22701,N_16537,N_16089);
or U22702 (N_22702,N_17708,N_17105);
nor U22703 (N_22703,N_18654,N_16820);
xnor U22704 (N_22704,N_19795,N_16060);
xnor U22705 (N_22705,N_18774,N_15057);
nand U22706 (N_22706,N_15083,N_18604);
nand U22707 (N_22707,N_19710,N_18339);
and U22708 (N_22708,N_16072,N_17514);
or U22709 (N_22709,N_16478,N_15783);
and U22710 (N_22710,N_16424,N_17455);
nand U22711 (N_22711,N_15509,N_18954);
and U22712 (N_22712,N_15509,N_18056);
nor U22713 (N_22713,N_19605,N_18491);
and U22714 (N_22714,N_15999,N_16525);
nand U22715 (N_22715,N_15501,N_18705);
nand U22716 (N_22716,N_17425,N_16965);
nor U22717 (N_22717,N_19387,N_19275);
nand U22718 (N_22718,N_15218,N_16428);
nand U22719 (N_22719,N_18348,N_16967);
or U22720 (N_22720,N_19821,N_19685);
xor U22721 (N_22721,N_17746,N_19412);
xnor U22722 (N_22722,N_15272,N_17526);
xor U22723 (N_22723,N_18014,N_17695);
and U22724 (N_22724,N_17482,N_19549);
nor U22725 (N_22725,N_19001,N_15518);
or U22726 (N_22726,N_16468,N_17041);
or U22727 (N_22727,N_18294,N_15655);
and U22728 (N_22728,N_19120,N_17640);
and U22729 (N_22729,N_15190,N_15887);
nor U22730 (N_22730,N_18360,N_16398);
nor U22731 (N_22731,N_19965,N_15706);
and U22732 (N_22732,N_17866,N_18059);
nor U22733 (N_22733,N_15811,N_16306);
nand U22734 (N_22734,N_19383,N_19072);
and U22735 (N_22735,N_18029,N_18459);
nand U22736 (N_22736,N_16924,N_16354);
or U22737 (N_22737,N_15091,N_18775);
xnor U22738 (N_22738,N_16719,N_16339);
nand U22739 (N_22739,N_16706,N_15773);
and U22740 (N_22740,N_16272,N_19561);
nor U22741 (N_22741,N_18186,N_16160);
nand U22742 (N_22742,N_15062,N_16706);
nand U22743 (N_22743,N_17333,N_15381);
nand U22744 (N_22744,N_17034,N_18729);
nand U22745 (N_22745,N_19290,N_16458);
or U22746 (N_22746,N_16574,N_15407);
or U22747 (N_22747,N_18580,N_18969);
nor U22748 (N_22748,N_16061,N_19873);
nor U22749 (N_22749,N_17802,N_17382);
nand U22750 (N_22750,N_16431,N_15485);
and U22751 (N_22751,N_15359,N_19192);
or U22752 (N_22752,N_16141,N_15557);
nand U22753 (N_22753,N_17645,N_18635);
nor U22754 (N_22754,N_17384,N_15749);
or U22755 (N_22755,N_18654,N_19520);
and U22756 (N_22756,N_19961,N_16823);
nand U22757 (N_22757,N_16829,N_17047);
nor U22758 (N_22758,N_17046,N_16802);
xor U22759 (N_22759,N_15096,N_17095);
and U22760 (N_22760,N_16235,N_17961);
and U22761 (N_22761,N_18227,N_18539);
nor U22762 (N_22762,N_18616,N_18293);
or U22763 (N_22763,N_18710,N_18214);
nand U22764 (N_22764,N_16414,N_17781);
or U22765 (N_22765,N_19369,N_18069);
xor U22766 (N_22766,N_17783,N_17806);
or U22767 (N_22767,N_18798,N_18029);
xor U22768 (N_22768,N_19208,N_19315);
and U22769 (N_22769,N_19693,N_15088);
and U22770 (N_22770,N_17822,N_15671);
or U22771 (N_22771,N_19281,N_19071);
or U22772 (N_22772,N_19892,N_17215);
and U22773 (N_22773,N_17867,N_16125);
xor U22774 (N_22774,N_18544,N_19949);
xor U22775 (N_22775,N_17424,N_15628);
or U22776 (N_22776,N_17901,N_15349);
and U22777 (N_22777,N_15823,N_17901);
xnor U22778 (N_22778,N_19396,N_17926);
and U22779 (N_22779,N_19388,N_15320);
and U22780 (N_22780,N_18772,N_19963);
nor U22781 (N_22781,N_16844,N_19797);
and U22782 (N_22782,N_15410,N_19525);
and U22783 (N_22783,N_17650,N_16925);
or U22784 (N_22784,N_15403,N_18865);
nand U22785 (N_22785,N_16617,N_15471);
and U22786 (N_22786,N_16965,N_17413);
and U22787 (N_22787,N_19245,N_19183);
or U22788 (N_22788,N_19485,N_17181);
or U22789 (N_22789,N_17831,N_16660);
nand U22790 (N_22790,N_15740,N_18153);
and U22791 (N_22791,N_18960,N_17691);
nor U22792 (N_22792,N_17773,N_15203);
nor U22793 (N_22793,N_17020,N_15412);
or U22794 (N_22794,N_15984,N_18882);
and U22795 (N_22795,N_17581,N_19694);
xnor U22796 (N_22796,N_15490,N_19936);
nor U22797 (N_22797,N_17390,N_19292);
or U22798 (N_22798,N_18719,N_19674);
xor U22799 (N_22799,N_17794,N_15754);
xnor U22800 (N_22800,N_19705,N_16593);
nor U22801 (N_22801,N_16184,N_17714);
nand U22802 (N_22802,N_19770,N_17177);
and U22803 (N_22803,N_19062,N_19699);
nor U22804 (N_22804,N_17811,N_18378);
nor U22805 (N_22805,N_17616,N_17478);
nand U22806 (N_22806,N_19093,N_18351);
nor U22807 (N_22807,N_16396,N_17568);
or U22808 (N_22808,N_16711,N_19829);
and U22809 (N_22809,N_19295,N_17092);
and U22810 (N_22810,N_18903,N_16199);
nor U22811 (N_22811,N_19850,N_19101);
and U22812 (N_22812,N_19364,N_16035);
nand U22813 (N_22813,N_19104,N_19637);
and U22814 (N_22814,N_15785,N_16088);
or U22815 (N_22815,N_19608,N_17236);
xor U22816 (N_22816,N_16356,N_16173);
or U22817 (N_22817,N_16028,N_17727);
nor U22818 (N_22818,N_19851,N_15593);
and U22819 (N_22819,N_17338,N_17090);
or U22820 (N_22820,N_16375,N_16766);
xnor U22821 (N_22821,N_18800,N_16186);
or U22822 (N_22822,N_16213,N_17580);
or U22823 (N_22823,N_17939,N_18610);
and U22824 (N_22824,N_19939,N_17105);
nor U22825 (N_22825,N_17664,N_17861);
and U22826 (N_22826,N_16076,N_15432);
or U22827 (N_22827,N_16258,N_17301);
and U22828 (N_22828,N_16234,N_17912);
nor U22829 (N_22829,N_18522,N_15577);
or U22830 (N_22830,N_15429,N_16245);
nand U22831 (N_22831,N_17438,N_16721);
xnor U22832 (N_22832,N_15237,N_15390);
or U22833 (N_22833,N_15507,N_15089);
and U22834 (N_22834,N_15255,N_16677);
or U22835 (N_22835,N_16563,N_17351);
and U22836 (N_22836,N_15087,N_18059);
nor U22837 (N_22837,N_18357,N_15872);
nand U22838 (N_22838,N_19531,N_19299);
or U22839 (N_22839,N_19234,N_17856);
nor U22840 (N_22840,N_16862,N_18694);
nand U22841 (N_22841,N_15165,N_19160);
nand U22842 (N_22842,N_18604,N_15802);
or U22843 (N_22843,N_16062,N_19453);
nand U22844 (N_22844,N_17422,N_16432);
or U22845 (N_22845,N_15989,N_16848);
xor U22846 (N_22846,N_17819,N_18332);
and U22847 (N_22847,N_17358,N_15552);
or U22848 (N_22848,N_16172,N_18934);
nor U22849 (N_22849,N_19002,N_15894);
xnor U22850 (N_22850,N_15528,N_15433);
or U22851 (N_22851,N_16808,N_18754);
nor U22852 (N_22852,N_17535,N_15039);
or U22853 (N_22853,N_17948,N_18708);
or U22854 (N_22854,N_18940,N_19572);
nand U22855 (N_22855,N_16471,N_17660);
and U22856 (N_22856,N_19682,N_15523);
nor U22857 (N_22857,N_17907,N_17677);
nor U22858 (N_22858,N_16786,N_17131);
nand U22859 (N_22859,N_15862,N_16868);
nand U22860 (N_22860,N_15396,N_15597);
or U22861 (N_22861,N_17087,N_16747);
or U22862 (N_22862,N_17226,N_18755);
nor U22863 (N_22863,N_15015,N_16643);
nor U22864 (N_22864,N_18210,N_18444);
nor U22865 (N_22865,N_18370,N_16004);
nor U22866 (N_22866,N_19012,N_17108);
nand U22867 (N_22867,N_19052,N_19127);
or U22868 (N_22868,N_15170,N_18104);
or U22869 (N_22869,N_17970,N_15501);
nor U22870 (N_22870,N_16805,N_19540);
and U22871 (N_22871,N_18444,N_15511);
nor U22872 (N_22872,N_18543,N_16401);
and U22873 (N_22873,N_18800,N_15991);
nor U22874 (N_22874,N_19137,N_19099);
or U22875 (N_22875,N_16386,N_16313);
or U22876 (N_22876,N_15188,N_17119);
nand U22877 (N_22877,N_19333,N_16023);
and U22878 (N_22878,N_15696,N_19953);
nand U22879 (N_22879,N_17291,N_17518);
xor U22880 (N_22880,N_15471,N_16339);
or U22881 (N_22881,N_16926,N_19953);
or U22882 (N_22882,N_19589,N_16141);
nor U22883 (N_22883,N_17159,N_17826);
nand U22884 (N_22884,N_15599,N_16153);
or U22885 (N_22885,N_15755,N_15851);
nor U22886 (N_22886,N_15825,N_19688);
nor U22887 (N_22887,N_19076,N_16648);
nor U22888 (N_22888,N_17691,N_16630);
nand U22889 (N_22889,N_19082,N_19421);
nand U22890 (N_22890,N_15846,N_17677);
nand U22891 (N_22891,N_18303,N_18144);
or U22892 (N_22892,N_19127,N_16983);
nor U22893 (N_22893,N_18600,N_18916);
nor U22894 (N_22894,N_19956,N_18436);
nor U22895 (N_22895,N_16424,N_16440);
xnor U22896 (N_22896,N_15395,N_19675);
nor U22897 (N_22897,N_15705,N_19733);
nand U22898 (N_22898,N_19475,N_18375);
nand U22899 (N_22899,N_19108,N_18422);
nand U22900 (N_22900,N_19680,N_19450);
nand U22901 (N_22901,N_19045,N_19292);
and U22902 (N_22902,N_15890,N_18996);
or U22903 (N_22903,N_16613,N_19481);
and U22904 (N_22904,N_17606,N_19255);
or U22905 (N_22905,N_18869,N_15875);
or U22906 (N_22906,N_16483,N_17137);
nand U22907 (N_22907,N_18494,N_17011);
nor U22908 (N_22908,N_16489,N_16749);
xnor U22909 (N_22909,N_19106,N_16945);
or U22910 (N_22910,N_15593,N_19823);
nor U22911 (N_22911,N_16672,N_16063);
nand U22912 (N_22912,N_18768,N_15885);
or U22913 (N_22913,N_16133,N_19653);
nand U22914 (N_22914,N_18939,N_17987);
and U22915 (N_22915,N_15989,N_19171);
nor U22916 (N_22916,N_15681,N_19225);
and U22917 (N_22917,N_16376,N_16268);
and U22918 (N_22918,N_17117,N_17992);
or U22919 (N_22919,N_15818,N_17958);
or U22920 (N_22920,N_19609,N_19749);
nor U22921 (N_22921,N_17974,N_19059);
nor U22922 (N_22922,N_19904,N_15488);
nand U22923 (N_22923,N_15416,N_17479);
nand U22924 (N_22924,N_18100,N_18270);
and U22925 (N_22925,N_16702,N_18659);
nand U22926 (N_22926,N_15087,N_19438);
nor U22927 (N_22927,N_16675,N_19695);
and U22928 (N_22928,N_18425,N_16680);
xor U22929 (N_22929,N_17275,N_16138);
or U22930 (N_22930,N_16819,N_18937);
nor U22931 (N_22931,N_17848,N_15996);
nand U22932 (N_22932,N_17097,N_17651);
or U22933 (N_22933,N_19670,N_17126);
and U22934 (N_22934,N_17272,N_18501);
or U22935 (N_22935,N_18668,N_16402);
or U22936 (N_22936,N_16765,N_18166);
or U22937 (N_22937,N_16225,N_19607);
nand U22938 (N_22938,N_17994,N_15679);
and U22939 (N_22939,N_19389,N_15768);
nor U22940 (N_22940,N_19074,N_18091);
xnor U22941 (N_22941,N_15452,N_18691);
and U22942 (N_22942,N_15646,N_18567);
nand U22943 (N_22943,N_15438,N_19037);
nor U22944 (N_22944,N_16361,N_19258);
or U22945 (N_22945,N_17121,N_16935);
xor U22946 (N_22946,N_15635,N_17754);
nor U22947 (N_22947,N_16998,N_19793);
xnor U22948 (N_22948,N_15528,N_18832);
or U22949 (N_22949,N_15569,N_15924);
and U22950 (N_22950,N_16309,N_17145);
and U22951 (N_22951,N_19456,N_15056);
xor U22952 (N_22952,N_18643,N_15262);
and U22953 (N_22953,N_16536,N_16951);
nand U22954 (N_22954,N_15525,N_17711);
or U22955 (N_22955,N_15662,N_18513);
or U22956 (N_22956,N_19356,N_15823);
or U22957 (N_22957,N_19966,N_17936);
nand U22958 (N_22958,N_18464,N_16793);
or U22959 (N_22959,N_18442,N_15543);
and U22960 (N_22960,N_15232,N_19558);
or U22961 (N_22961,N_16870,N_18295);
or U22962 (N_22962,N_16164,N_18295);
xor U22963 (N_22963,N_17937,N_18675);
and U22964 (N_22964,N_16593,N_16206);
nor U22965 (N_22965,N_17510,N_16602);
nand U22966 (N_22966,N_17206,N_18634);
and U22967 (N_22967,N_18305,N_15113);
or U22968 (N_22968,N_15491,N_16400);
or U22969 (N_22969,N_15488,N_19491);
or U22970 (N_22970,N_17391,N_15880);
or U22971 (N_22971,N_15863,N_17806);
nor U22972 (N_22972,N_15079,N_18798);
nor U22973 (N_22973,N_18848,N_16895);
xnor U22974 (N_22974,N_16791,N_18569);
nand U22975 (N_22975,N_15058,N_17087);
xnor U22976 (N_22976,N_16755,N_17706);
nor U22977 (N_22977,N_15419,N_17479);
and U22978 (N_22978,N_17439,N_18631);
and U22979 (N_22979,N_15203,N_15244);
xnor U22980 (N_22980,N_17379,N_19829);
and U22981 (N_22981,N_19548,N_19188);
nor U22982 (N_22982,N_18322,N_19813);
or U22983 (N_22983,N_16642,N_18378);
xor U22984 (N_22984,N_18248,N_15546);
nor U22985 (N_22985,N_18358,N_15214);
or U22986 (N_22986,N_19746,N_19170);
nor U22987 (N_22987,N_16940,N_19138);
nor U22988 (N_22988,N_19573,N_17866);
and U22989 (N_22989,N_16327,N_18288);
and U22990 (N_22990,N_19311,N_15300);
and U22991 (N_22991,N_17559,N_17806);
and U22992 (N_22992,N_15504,N_19598);
nor U22993 (N_22993,N_19263,N_18582);
and U22994 (N_22994,N_17578,N_18782);
nor U22995 (N_22995,N_15800,N_15253);
or U22996 (N_22996,N_18206,N_15113);
nand U22997 (N_22997,N_15086,N_19311);
nand U22998 (N_22998,N_17964,N_15333);
nand U22999 (N_22999,N_16832,N_15543);
nor U23000 (N_23000,N_15821,N_15959);
nand U23001 (N_23001,N_18426,N_18174);
or U23002 (N_23002,N_18354,N_19179);
nor U23003 (N_23003,N_17794,N_15544);
and U23004 (N_23004,N_17865,N_17546);
and U23005 (N_23005,N_15873,N_18625);
nand U23006 (N_23006,N_17767,N_17194);
nand U23007 (N_23007,N_18494,N_18485);
xor U23008 (N_23008,N_15258,N_17227);
nand U23009 (N_23009,N_19277,N_16963);
or U23010 (N_23010,N_16804,N_17642);
nor U23011 (N_23011,N_16757,N_19263);
nor U23012 (N_23012,N_18818,N_18250);
nand U23013 (N_23013,N_17418,N_15781);
or U23014 (N_23014,N_19803,N_17503);
or U23015 (N_23015,N_15070,N_18273);
and U23016 (N_23016,N_16729,N_16571);
nand U23017 (N_23017,N_18025,N_18079);
or U23018 (N_23018,N_18186,N_18855);
xor U23019 (N_23019,N_18999,N_16201);
nand U23020 (N_23020,N_15454,N_15260);
and U23021 (N_23021,N_16772,N_16349);
or U23022 (N_23022,N_17008,N_17498);
or U23023 (N_23023,N_16429,N_15986);
and U23024 (N_23024,N_17692,N_19883);
nand U23025 (N_23025,N_16949,N_17365);
xnor U23026 (N_23026,N_15302,N_18851);
or U23027 (N_23027,N_15233,N_15237);
and U23028 (N_23028,N_19958,N_19336);
xor U23029 (N_23029,N_16061,N_16864);
and U23030 (N_23030,N_15811,N_18589);
xnor U23031 (N_23031,N_17310,N_18242);
nor U23032 (N_23032,N_17263,N_17712);
nand U23033 (N_23033,N_17627,N_17266);
and U23034 (N_23034,N_15228,N_18256);
or U23035 (N_23035,N_16685,N_19430);
and U23036 (N_23036,N_16665,N_19888);
nor U23037 (N_23037,N_19500,N_16799);
or U23038 (N_23038,N_18106,N_18270);
nand U23039 (N_23039,N_19848,N_17473);
xor U23040 (N_23040,N_18166,N_19402);
nor U23041 (N_23041,N_16994,N_19756);
nor U23042 (N_23042,N_19616,N_19222);
nand U23043 (N_23043,N_16741,N_18711);
xnor U23044 (N_23044,N_19013,N_17162);
nand U23045 (N_23045,N_19667,N_18008);
and U23046 (N_23046,N_15308,N_15408);
or U23047 (N_23047,N_18014,N_19000);
xor U23048 (N_23048,N_15572,N_17278);
xor U23049 (N_23049,N_18602,N_19998);
or U23050 (N_23050,N_18662,N_18048);
and U23051 (N_23051,N_19422,N_15555);
or U23052 (N_23052,N_19731,N_16778);
and U23053 (N_23053,N_17482,N_18713);
or U23054 (N_23054,N_15491,N_19169);
or U23055 (N_23055,N_19053,N_18150);
or U23056 (N_23056,N_17534,N_17766);
nand U23057 (N_23057,N_17940,N_16029);
nand U23058 (N_23058,N_17597,N_15131);
and U23059 (N_23059,N_16140,N_19069);
nor U23060 (N_23060,N_16612,N_16468);
or U23061 (N_23061,N_15281,N_19976);
or U23062 (N_23062,N_16302,N_16608);
nor U23063 (N_23063,N_15711,N_15348);
nand U23064 (N_23064,N_15907,N_18554);
or U23065 (N_23065,N_17516,N_16223);
xor U23066 (N_23066,N_16140,N_17236);
nor U23067 (N_23067,N_17206,N_16813);
nor U23068 (N_23068,N_15304,N_16217);
or U23069 (N_23069,N_16038,N_16314);
or U23070 (N_23070,N_17850,N_16445);
xor U23071 (N_23071,N_15074,N_16691);
xor U23072 (N_23072,N_17230,N_17205);
xnor U23073 (N_23073,N_15210,N_16326);
and U23074 (N_23074,N_18644,N_18153);
nor U23075 (N_23075,N_19976,N_15981);
nand U23076 (N_23076,N_16966,N_17315);
nor U23077 (N_23077,N_15776,N_18016);
or U23078 (N_23078,N_17011,N_15270);
nand U23079 (N_23079,N_19539,N_19709);
nor U23080 (N_23080,N_15302,N_19383);
nand U23081 (N_23081,N_19623,N_19929);
nand U23082 (N_23082,N_15982,N_15025);
and U23083 (N_23083,N_16231,N_19446);
and U23084 (N_23084,N_18680,N_15262);
or U23085 (N_23085,N_16136,N_17642);
xnor U23086 (N_23086,N_15251,N_17412);
or U23087 (N_23087,N_18652,N_15417);
nand U23088 (N_23088,N_18771,N_19057);
nand U23089 (N_23089,N_19107,N_19514);
xnor U23090 (N_23090,N_18830,N_17392);
and U23091 (N_23091,N_17850,N_17913);
or U23092 (N_23092,N_19466,N_18858);
nand U23093 (N_23093,N_15204,N_16446);
nor U23094 (N_23094,N_18936,N_19742);
and U23095 (N_23095,N_17711,N_19488);
or U23096 (N_23096,N_19086,N_19975);
or U23097 (N_23097,N_15134,N_16330);
or U23098 (N_23098,N_15931,N_17259);
nor U23099 (N_23099,N_18233,N_16758);
and U23100 (N_23100,N_17027,N_15680);
or U23101 (N_23101,N_18944,N_16823);
xor U23102 (N_23102,N_16414,N_19975);
or U23103 (N_23103,N_16996,N_17598);
or U23104 (N_23104,N_16821,N_18681);
nand U23105 (N_23105,N_17644,N_15718);
nor U23106 (N_23106,N_17609,N_15167);
or U23107 (N_23107,N_16759,N_15630);
xnor U23108 (N_23108,N_15028,N_16687);
nor U23109 (N_23109,N_15262,N_19560);
nor U23110 (N_23110,N_17703,N_18405);
nand U23111 (N_23111,N_17095,N_19658);
and U23112 (N_23112,N_18420,N_18689);
nand U23113 (N_23113,N_18519,N_16238);
or U23114 (N_23114,N_17749,N_17080);
nand U23115 (N_23115,N_16923,N_15344);
nor U23116 (N_23116,N_19431,N_18988);
or U23117 (N_23117,N_15590,N_18814);
and U23118 (N_23118,N_19259,N_16970);
nand U23119 (N_23119,N_18567,N_16604);
or U23120 (N_23120,N_19141,N_15161);
or U23121 (N_23121,N_17472,N_17568);
or U23122 (N_23122,N_15368,N_19120);
and U23123 (N_23123,N_17045,N_15491);
and U23124 (N_23124,N_15491,N_19225);
xnor U23125 (N_23125,N_15334,N_15502);
nor U23126 (N_23126,N_15057,N_16345);
or U23127 (N_23127,N_16811,N_15916);
xnor U23128 (N_23128,N_17878,N_17927);
and U23129 (N_23129,N_15894,N_18264);
and U23130 (N_23130,N_16645,N_17792);
nor U23131 (N_23131,N_17539,N_17517);
nand U23132 (N_23132,N_18957,N_18704);
and U23133 (N_23133,N_19232,N_16827);
xor U23134 (N_23134,N_16213,N_16415);
or U23135 (N_23135,N_18976,N_18923);
nor U23136 (N_23136,N_16177,N_18751);
nand U23137 (N_23137,N_16247,N_18602);
nand U23138 (N_23138,N_15227,N_17110);
xor U23139 (N_23139,N_18251,N_18013);
nand U23140 (N_23140,N_19927,N_16047);
nor U23141 (N_23141,N_15063,N_15353);
or U23142 (N_23142,N_17837,N_17605);
or U23143 (N_23143,N_15982,N_18947);
or U23144 (N_23144,N_18203,N_16069);
or U23145 (N_23145,N_16585,N_19566);
or U23146 (N_23146,N_16430,N_19940);
nor U23147 (N_23147,N_17562,N_15480);
and U23148 (N_23148,N_15050,N_15569);
or U23149 (N_23149,N_18686,N_15135);
and U23150 (N_23150,N_18060,N_15046);
nor U23151 (N_23151,N_18675,N_15355);
and U23152 (N_23152,N_18523,N_17467);
and U23153 (N_23153,N_18837,N_19545);
and U23154 (N_23154,N_18210,N_17517);
or U23155 (N_23155,N_16765,N_19041);
nor U23156 (N_23156,N_17112,N_17337);
nand U23157 (N_23157,N_15053,N_17667);
nor U23158 (N_23158,N_18562,N_18185);
nand U23159 (N_23159,N_15832,N_19236);
and U23160 (N_23160,N_18267,N_16702);
and U23161 (N_23161,N_15263,N_15962);
and U23162 (N_23162,N_16506,N_15361);
and U23163 (N_23163,N_17297,N_16567);
and U23164 (N_23164,N_17856,N_15497);
or U23165 (N_23165,N_18296,N_16021);
or U23166 (N_23166,N_15121,N_16854);
or U23167 (N_23167,N_16411,N_16634);
or U23168 (N_23168,N_17747,N_18900);
or U23169 (N_23169,N_17372,N_18847);
and U23170 (N_23170,N_19908,N_18800);
and U23171 (N_23171,N_17033,N_15884);
nor U23172 (N_23172,N_17263,N_15280);
nor U23173 (N_23173,N_15564,N_16746);
nor U23174 (N_23174,N_19949,N_15493);
or U23175 (N_23175,N_15765,N_16808);
nand U23176 (N_23176,N_15565,N_19207);
nand U23177 (N_23177,N_18370,N_16436);
or U23178 (N_23178,N_18113,N_18337);
and U23179 (N_23179,N_19905,N_17840);
nor U23180 (N_23180,N_15113,N_18428);
nor U23181 (N_23181,N_18886,N_17885);
nand U23182 (N_23182,N_19767,N_18592);
nand U23183 (N_23183,N_18851,N_18724);
nor U23184 (N_23184,N_16341,N_19901);
or U23185 (N_23185,N_16355,N_17939);
nor U23186 (N_23186,N_16145,N_16307);
nor U23187 (N_23187,N_17593,N_15196);
nor U23188 (N_23188,N_16994,N_15396);
or U23189 (N_23189,N_15449,N_16209);
nor U23190 (N_23190,N_18148,N_19347);
nand U23191 (N_23191,N_19730,N_18691);
nand U23192 (N_23192,N_15318,N_19983);
and U23193 (N_23193,N_17019,N_17850);
nor U23194 (N_23194,N_17490,N_15825);
or U23195 (N_23195,N_17380,N_15435);
nand U23196 (N_23196,N_17185,N_15740);
and U23197 (N_23197,N_16943,N_16139);
nor U23198 (N_23198,N_16942,N_18514);
nand U23199 (N_23199,N_19290,N_16688);
xor U23200 (N_23200,N_16591,N_18982);
nand U23201 (N_23201,N_18868,N_19394);
nor U23202 (N_23202,N_17586,N_17542);
nand U23203 (N_23203,N_15876,N_18655);
xnor U23204 (N_23204,N_19583,N_16993);
nand U23205 (N_23205,N_18505,N_15968);
and U23206 (N_23206,N_18065,N_16452);
nand U23207 (N_23207,N_15940,N_15941);
or U23208 (N_23208,N_15172,N_17922);
nor U23209 (N_23209,N_19602,N_17815);
nor U23210 (N_23210,N_18792,N_17900);
and U23211 (N_23211,N_17972,N_19138);
or U23212 (N_23212,N_18751,N_17389);
and U23213 (N_23213,N_19730,N_16707);
and U23214 (N_23214,N_16344,N_15487);
nand U23215 (N_23215,N_19118,N_16652);
nor U23216 (N_23216,N_17225,N_17170);
nor U23217 (N_23217,N_16181,N_19212);
and U23218 (N_23218,N_15833,N_15552);
or U23219 (N_23219,N_19869,N_17010);
nor U23220 (N_23220,N_15263,N_16934);
nand U23221 (N_23221,N_16218,N_16054);
or U23222 (N_23222,N_18280,N_19156);
nand U23223 (N_23223,N_16565,N_17199);
nand U23224 (N_23224,N_17756,N_16914);
nand U23225 (N_23225,N_18009,N_15804);
nor U23226 (N_23226,N_19884,N_16187);
xor U23227 (N_23227,N_18912,N_16628);
and U23228 (N_23228,N_19792,N_17154);
nor U23229 (N_23229,N_19788,N_17951);
xor U23230 (N_23230,N_18767,N_17194);
nand U23231 (N_23231,N_19891,N_15948);
and U23232 (N_23232,N_15732,N_16127);
nand U23233 (N_23233,N_19684,N_18810);
xor U23234 (N_23234,N_17771,N_19657);
or U23235 (N_23235,N_17894,N_19619);
and U23236 (N_23236,N_19892,N_17960);
nand U23237 (N_23237,N_16921,N_17957);
nor U23238 (N_23238,N_17093,N_18429);
nand U23239 (N_23239,N_16117,N_18214);
nor U23240 (N_23240,N_19205,N_16967);
nand U23241 (N_23241,N_19333,N_19427);
or U23242 (N_23242,N_16747,N_19854);
nor U23243 (N_23243,N_17972,N_18000);
and U23244 (N_23244,N_17670,N_16618);
or U23245 (N_23245,N_19056,N_15333);
nor U23246 (N_23246,N_16168,N_16829);
or U23247 (N_23247,N_18706,N_15779);
nand U23248 (N_23248,N_19152,N_17110);
and U23249 (N_23249,N_19966,N_17346);
nor U23250 (N_23250,N_19674,N_19191);
or U23251 (N_23251,N_16443,N_18328);
or U23252 (N_23252,N_15772,N_16591);
xnor U23253 (N_23253,N_18754,N_15445);
and U23254 (N_23254,N_18921,N_19900);
nand U23255 (N_23255,N_15018,N_19235);
nor U23256 (N_23256,N_17431,N_19012);
nor U23257 (N_23257,N_18435,N_19676);
and U23258 (N_23258,N_17590,N_16940);
or U23259 (N_23259,N_16434,N_15921);
nand U23260 (N_23260,N_18574,N_16889);
nor U23261 (N_23261,N_18141,N_19900);
xor U23262 (N_23262,N_17177,N_16526);
nand U23263 (N_23263,N_18531,N_17670);
xnor U23264 (N_23264,N_15892,N_18435);
nor U23265 (N_23265,N_19276,N_16737);
nand U23266 (N_23266,N_16815,N_19601);
or U23267 (N_23267,N_19404,N_15477);
nor U23268 (N_23268,N_16485,N_15787);
or U23269 (N_23269,N_17667,N_17237);
and U23270 (N_23270,N_17837,N_15731);
or U23271 (N_23271,N_15890,N_18101);
and U23272 (N_23272,N_16311,N_19745);
nor U23273 (N_23273,N_19332,N_16628);
or U23274 (N_23274,N_16460,N_16610);
and U23275 (N_23275,N_16447,N_19343);
or U23276 (N_23276,N_16721,N_17945);
xnor U23277 (N_23277,N_15030,N_18677);
or U23278 (N_23278,N_18985,N_17167);
or U23279 (N_23279,N_19014,N_18475);
or U23280 (N_23280,N_15848,N_17282);
and U23281 (N_23281,N_18825,N_15049);
and U23282 (N_23282,N_15534,N_19542);
nor U23283 (N_23283,N_15808,N_18486);
or U23284 (N_23284,N_15891,N_18660);
and U23285 (N_23285,N_18095,N_19319);
nand U23286 (N_23286,N_16903,N_17083);
xnor U23287 (N_23287,N_17804,N_17712);
nor U23288 (N_23288,N_16925,N_15013);
or U23289 (N_23289,N_16669,N_17381);
xnor U23290 (N_23290,N_18946,N_18201);
and U23291 (N_23291,N_18644,N_15934);
and U23292 (N_23292,N_17416,N_15204);
and U23293 (N_23293,N_19609,N_19406);
xor U23294 (N_23294,N_15349,N_16961);
and U23295 (N_23295,N_15973,N_15601);
or U23296 (N_23296,N_16520,N_15331);
or U23297 (N_23297,N_17263,N_16355);
xor U23298 (N_23298,N_15282,N_19754);
nand U23299 (N_23299,N_15767,N_17204);
nand U23300 (N_23300,N_17986,N_19737);
and U23301 (N_23301,N_19726,N_18419);
or U23302 (N_23302,N_17887,N_15247);
and U23303 (N_23303,N_15877,N_16063);
nand U23304 (N_23304,N_19609,N_16834);
nor U23305 (N_23305,N_16282,N_18437);
and U23306 (N_23306,N_17575,N_16705);
nor U23307 (N_23307,N_15673,N_16813);
nor U23308 (N_23308,N_19110,N_17104);
nand U23309 (N_23309,N_18545,N_17614);
and U23310 (N_23310,N_17755,N_17094);
nor U23311 (N_23311,N_17575,N_18467);
nor U23312 (N_23312,N_15749,N_18186);
or U23313 (N_23313,N_16268,N_19552);
nand U23314 (N_23314,N_16553,N_19537);
and U23315 (N_23315,N_17392,N_18584);
nor U23316 (N_23316,N_16810,N_18457);
and U23317 (N_23317,N_15234,N_17613);
and U23318 (N_23318,N_19229,N_19928);
and U23319 (N_23319,N_16437,N_16098);
and U23320 (N_23320,N_19548,N_15628);
nor U23321 (N_23321,N_19559,N_17149);
xor U23322 (N_23322,N_18034,N_18677);
nand U23323 (N_23323,N_19974,N_16871);
nand U23324 (N_23324,N_18846,N_17136);
xor U23325 (N_23325,N_18126,N_19685);
or U23326 (N_23326,N_19495,N_19061);
or U23327 (N_23327,N_19831,N_15867);
nor U23328 (N_23328,N_18450,N_17938);
nor U23329 (N_23329,N_15916,N_16178);
and U23330 (N_23330,N_17901,N_17840);
xnor U23331 (N_23331,N_16173,N_17235);
and U23332 (N_23332,N_19792,N_15322);
nor U23333 (N_23333,N_16660,N_18574);
and U23334 (N_23334,N_15275,N_17865);
nor U23335 (N_23335,N_19645,N_18379);
and U23336 (N_23336,N_18233,N_15467);
and U23337 (N_23337,N_16760,N_15939);
or U23338 (N_23338,N_16963,N_19432);
and U23339 (N_23339,N_18360,N_17512);
xor U23340 (N_23340,N_15195,N_15185);
or U23341 (N_23341,N_15999,N_16819);
or U23342 (N_23342,N_19695,N_18566);
nor U23343 (N_23343,N_18668,N_15923);
nand U23344 (N_23344,N_19772,N_19900);
or U23345 (N_23345,N_17779,N_19620);
nand U23346 (N_23346,N_19965,N_15988);
and U23347 (N_23347,N_18620,N_19255);
or U23348 (N_23348,N_17895,N_18408);
xnor U23349 (N_23349,N_18064,N_17248);
nor U23350 (N_23350,N_17506,N_17408);
nand U23351 (N_23351,N_19225,N_18048);
nor U23352 (N_23352,N_17085,N_19856);
nand U23353 (N_23353,N_19465,N_17879);
and U23354 (N_23354,N_16315,N_19284);
nand U23355 (N_23355,N_18349,N_16963);
and U23356 (N_23356,N_19717,N_19665);
xnor U23357 (N_23357,N_16023,N_17714);
and U23358 (N_23358,N_17369,N_15257);
nand U23359 (N_23359,N_15722,N_17052);
nand U23360 (N_23360,N_15416,N_17665);
xnor U23361 (N_23361,N_19028,N_18552);
or U23362 (N_23362,N_18619,N_18730);
or U23363 (N_23363,N_18536,N_18177);
and U23364 (N_23364,N_18411,N_18937);
xnor U23365 (N_23365,N_19803,N_19682);
or U23366 (N_23366,N_18247,N_15049);
nand U23367 (N_23367,N_18350,N_19467);
xor U23368 (N_23368,N_17828,N_16116);
and U23369 (N_23369,N_17850,N_19213);
and U23370 (N_23370,N_18587,N_19274);
xnor U23371 (N_23371,N_18146,N_15090);
and U23372 (N_23372,N_19558,N_17360);
xnor U23373 (N_23373,N_16570,N_16572);
nor U23374 (N_23374,N_16868,N_18138);
or U23375 (N_23375,N_17562,N_18153);
nand U23376 (N_23376,N_17680,N_17461);
nand U23377 (N_23377,N_17793,N_19986);
or U23378 (N_23378,N_17646,N_16974);
nor U23379 (N_23379,N_16476,N_15165);
or U23380 (N_23380,N_16280,N_15967);
xnor U23381 (N_23381,N_15515,N_16650);
nand U23382 (N_23382,N_19720,N_18055);
nand U23383 (N_23383,N_18658,N_19844);
nand U23384 (N_23384,N_18936,N_17997);
or U23385 (N_23385,N_18871,N_16017);
nor U23386 (N_23386,N_16100,N_16027);
nor U23387 (N_23387,N_17137,N_15462);
or U23388 (N_23388,N_15998,N_16702);
and U23389 (N_23389,N_17871,N_16442);
and U23390 (N_23390,N_15350,N_15511);
nor U23391 (N_23391,N_19953,N_19226);
nand U23392 (N_23392,N_17094,N_17786);
xor U23393 (N_23393,N_18540,N_15142);
xnor U23394 (N_23394,N_18650,N_17447);
and U23395 (N_23395,N_15596,N_15665);
and U23396 (N_23396,N_19210,N_18095);
nor U23397 (N_23397,N_15296,N_18013);
xor U23398 (N_23398,N_18310,N_18745);
and U23399 (N_23399,N_19125,N_18867);
and U23400 (N_23400,N_18416,N_17636);
nor U23401 (N_23401,N_19967,N_18503);
nand U23402 (N_23402,N_18344,N_16792);
nor U23403 (N_23403,N_15099,N_19258);
nand U23404 (N_23404,N_19261,N_17086);
and U23405 (N_23405,N_15157,N_19554);
nand U23406 (N_23406,N_17541,N_18133);
nor U23407 (N_23407,N_18248,N_19357);
xnor U23408 (N_23408,N_18921,N_19523);
nand U23409 (N_23409,N_18591,N_18798);
xnor U23410 (N_23410,N_17035,N_19590);
xor U23411 (N_23411,N_16109,N_15683);
nand U23412 (N_23412,N_16619,N_18834);
nand U23413 (N_23413,N_17652,N_19150);
nand U23414 (N_23414,N_16346,N_18816);
or U23415 (N_23415,N_19153,N_16451);
nand U23416 (N_23416,N_16164,N_15547);
nand U23417 (N_23417,N_15602,N_16179);
and U23418 (N_23418,N_16259,N_18560);
nor U23419 (N_23419,N_18303,N_15242);
nand U23420 (N_23420,N_17628,N_17451);
nand U23421 (N_23421,N_15567,N_17185);
or U23422 (N_23422,N_17479,N_16162);
or U23423 (N_23423,N_17253,N_15274);
and U23424 (N_23424,N_19114,N_15419);
nand U23425 (N_23425,N_19643,N_16913);
nor U23426 (N_23426,N_18069,N_17918);
or U23427 (N_23427,N_19084,N_17549);
and U23428 (N_23428,N_18059,N_16634);
xnor U23429 (N_23429,N_15288,N_16039);
and U23430 (N_23430,N_19752,N_17907);
nand U23431 (N_23431,N_16909,N_15835);
nor U23432 (N_23432,N_18937,N_15465);
nor U23433 (N_23433,N_18496,N_17745);
nor U23434 (N_23434,N_19291,N_17983);
nor U23435 (N_23435,N_15805,N_16327);
or U23436 (N_23436,N_15329,N_16410);
nor U23437 (N_23437,N_18587,N_17572);
or U23438 (N_23438,N_16470,N_19464);
nor U23439 (N_23439,N_16049,N_16670);
nand U23440 (N_23440,N_15158,N_19116);
nand U23441 (N_23441,N_16546,N_17172);
or U23442 (N_23442,N_17352,N_16984);
xnor U23443 (N_23443,N_17353,N_17015);
or U23444 (N_23444,N_17859,N_19354);
and U23445 (N_23445,N_18163,N_19897);
nand U23446 (N_23446,N_16729,N_16795);
and U23447 (N_23447,N_19283,N_15267);
or U23448 (N_23448,N_19954,N_15382);
nand U23449 (N_23449,N_19264,N_17385);
xnor U23450 (N_23450,N_16735,N_16071);
xor U23451 (N_23451,N_16458,N_16431);
and U23452 (N_23452,N_19389,N_19854);
nor U23453 (N_23453,N_15551,N_17308);
and U23454 (N_23454,N_15044,N_18256);
or U23455 (N_23455,N_19066,N_15140);
nand U23456 (N_23456,N_19291,N_16936);
or U23457 (N_23457,N_18632,N_19533);
and U23458 (N_23458,N_15723,N_16316);
nor U23459 (N_23459,N_15666,N_17685);
nor U23460 (N_23460,N_15063,N_16313);
nand U23461 (N_23461,N_16841,N_15355);
or U23462 (N_23462,N_16210,N_17956);
nand U23463 (N_23463,N_16320,N_18188);
nand U23464 (N_23464,N_16434,N_17603);
nor U23465 (N_23465,N_17240,N_19824);
nand U23466 (N_23466,N_16224,N_16459);
nor U23467 (N_23467,N_15874,N_17985);
nand U23468 (N_23468,N_15865,N_18857);
nor U23469 (N_23469,N_19456,N_17451);
nor U23470 (N_23470,N_17247,N_17629);
nand U23471 (N_23471,N_17787,N_16062);
and U23472 (N_23472,N_17933,N_19011);
or U23473 (N_23473,N_17072,N_18956);
nand U23474 (N_23474,N_17673,N_16791);
nand U23475 (N_23475,N_16351,N_16898);
or U23476 (N_23476,N_15853,N_19882);
or U23477 (N_23477,N_16623,N_16649);
and U23478 (N_23478,N_16258,N_19902);
nand U23479 (N_23479,N_18661,N_17844);
nand U23480 (N_23480,N_17155,N_16490);
nand U23481 (N_23481,N_17661,N_18525);
or U23482 (N_23482,N_16993,N_17537);
nor U23483 (N_23483,N_18616,N_17064);
xor U23484 (N_23484,N_15600,N_16938);
nand U23485 (N_23485,N_16728,N_15659);
or U23486 (N_23486,N_15982,N_15218);
nor U23487 (N_23487,N_18454,N_19152);
or U23488 (N_23488,N_18215,N_18494);
or U23489 (N_23489,N_16942,N_19734);
nand U23490 (N_23490,N_15974,N_16382);
nor U23491 (N_23491,N_15255,N_18077);
nor U23492 (N_23492,N_16869,N_19867);
nand U23493 (N_23493,N_15238,N_18879);
nor U23494 (N_23494,N_18303,N_18891);
or U23495 (N_23495,N_18445,N_15195);
and U23496 (N_23496,N_16023,N_18290);
or U23497 (N_23497,N_19696,N_19732);
nand U23498 (N_23498,N_15297,N_16861);
and U23499 (N_23499,N_15903,N_15772);
or U23500 (N_23500,N_18579,N_19892);
nand U23501 (N_23501,N_15990,N_17153);
and U23502 (N_23502,N_18945,N_19154);
or U23503 (N_23503,N_17104,N_15134);
or U23504 (N_23504,N_17092,N_18128);
nand U23505 (N_23505,N_17338,N_19286);
or U23506 (N_23506,N_19783,N_15827);
and U23507 (N_23507,N_16477,N_19960);
nand U23508 (N_23508,N_17454,N_16643);
xor U23509 (N_23509,N_17849,N_19099);
and U23510 (N_23510,N_17413,N_16942);
and U23511 (N_23511,N_18585,N_19397);
nor U23512 (N_23512,N_19270,N_15059);
or U23513 (N_23513,N_18016,N_18832);
and U23514 (N_23514,N_15057,N_19874);
and U23515 (N_23515,N_15983,N_16599);
nor U23516 (N_23516,N_19133,N_15239);
nor U23517 (N_23517,N_16353,N_15265);
xnor U23518 (N_23518,N_16893,N_17646);
nand U23519 (N_23519,N_17323,N_15923);
xor U23520 (N_23520,N_15961,N_19111);
nand U23521 (N_23521,N_16343,N_19368);
xnor U23522 (N_23522,N_15528,N_18223);
and U23523 (N_23523,N_18674,N_17689);
and U23524 (N_23524,N_17101,N_19607);
and U23525 (N_23525,N_19878,N_15485);
or U23526 (N_23526,N_18187,N_18140);
and U23527 (N_23527,N_16233,N_17037);
nand U23528 (N_23528,N_19971,N_16094);
and U23529 (N_23529,N_17559,N_16807);
or U23530 (N_23530,N_18105,N_17967);
nor U23531 (N_23531,N_15851,N_16477);
xor U23532 (N_23532,N_19172,N_19244);
or U23533 (N_23533,N_16867,N_17706);
nand U23534 (N_23534,N_18453,N_17227);
nand U23535 (N_23535,N_18076,N_15814);
nand U23536 (N_23536,N_17104,N_15088);
and U23537 (N_23537,N_15917,N_16256);
or U23538 (N_23538,N_16205,N_15870);
or U23539 (N_23539,N_15865,N_18024);
or U23540 (N_23540,N_16680,N_19723);
nand U23541 (N_23541,N_17024,N_16288);
nor U23542 (N_23542,N_18609,N_16078);
and U23543 (N_23543,N_17551,N_19322);
or U23544 (N_23544,N_16148,N_16907);
nor U23545 (N_23545,N_19619,N_19774);
or U23546 (N_23546,N_16697,N_19886);
xnor U23547 (N_23547,N_18770,N_15544);
nand U23548 (N_23548,N_19341,N_18539);
xnor U23549 (N_23549,N_18068,N_19532);
nand U23550 (N_23550,N_19649,N_16172);
or U23551 (N_23551,N_16156,N_17405);
or U23552 (N_23552,N_18642,N_18976);
nor U23553 (N_23553,N_18746,N_15407);
nor U23554 (N_23554,N_15140,N_15514);
and U23555 (N_23555,N_18121,N_15656);
nand U23556 (N_23556,N_18621,N_17657);
nor U23557 (N_23557,N_19505,N_16051);
nand U23558 (N_23558,N_15940,N_16570);
or U23559 (N_23559,N_17316,N_15511);
nor U23560 (N_23560,N_16319,N_17875);
nand U23561 (N_23561,N_15151,N_19222);
and U23562 (N_23562,N_16800,N_19569);
nand U23563 (N_23563,N_19819,N_17524);
nor U23564 (N_23564,N_16870,N_16431);
xor U23565 (N_23565,N_18809,N_18020);
or U23566 (N_23566,N_19145,N_19441);
and U23567 (N_23567,N_16376,N_17214);
or U23568 (N_23568,N_19068,N_19165);
nand U23569 (N_23569,N_19974,N_19522);
and U23570 (N_23570,N_19513,N_18872);
nor U23571 (N_23571,N_15703,N_19722);
nor U23572 (N_23572,N_17875,N_15504);
or U23573 (N_23573,N_19744,N_15707);
nand U23574 (N_23574,N_18298,N_16628);
and U23575 (N_23575,N_15326,N_18306);
nor U23576 (N_23576,N_19182,N_17955);
nor U23577 (N_23577,N_17554,N_15902);
and U23578 (N_23578,N_16884,N_18879);
nand U23579 (N_23579,N_15883,N_17902);
or U23580 (N_23580,N_16942,N_19830);
nand U23581 (N_23581,N_18751,N_16892);
nor U23582 (N_23582,N_15052,N_15436);
or U23583 (N_23583,N_15235,N_17764);
nand U23584 (N_23584,N_18109,N_17537);
nor U23585 (N_23585,N_16537,N_17374);
and U23586 (N_23586,N_19021,N_18933);
nand U23587 (N_23587,N_18427,N_18889);
nand U23588 (N_23588,N_16781,N_19185);
or U23589 (N_23589,N_18191,N_15040);
nor U23590 (N_23590,N_18955,N_17535);
and U23591 (N_23591,N_18145,N_19079);
nor U23592 (N_23592,N_16120,N_19039);
nand U23593 (N_23593,N_16103,N_16951);
or U23594 (N_23594,N_19953,N_17014);
nor U23595 (N_23595,N_18586,N_15917);
xnor U23596 (N_23596,N_18289,N_18535);
or U23597 (N_23597,N_18791,N_16895);
and U23598 (N_23598,N_18939,N_19085);
xnor U23599 (N_23599,N_19283,N_17218);
and U23600 (N_23600,N_17199,N_17322);
nor U23601 (N_23601,N_17770,N_16402);
nand U23602 (N_23602,N_16499,N_15709);
nor U23603 (N_23603,N_17493,N_15552);
and U23604 (N_23604,N_18225,N_17893);
nor U23605 (N_23605,N_18569,N_15192);
or U23606 (N_23606,N_16133,N_19619);
nand U23607 (N_23607,N_17273,N_17155);
and U23608 (N_23608,N_15155,N_17082);
nand U23609 (N_23609,N_16986,N_19349);
and U23610 (N_23610,N_15946,N_16796);
or U23611 (N_23611,N_17540,N_18100);
nand U23612 (N_23612,N_15294,N_18452);
nand U23613 (N_23613,N_15243,N_19045);
or U23614 (N_23614,N_16892,N_18988);
nor U23615 (N_23615,N_18962,N_17110);
nor U23616 (N_23616,N_15109,N_18834);
or U23617 (N_23617,N_15877,N_19944);
or U23618 (N_23618,N_19005,N_18784);
nor U23619 (N_23619,N_17163,N_19624);
nor U23620 (N_23620,N_16003,N_19190);
nor U23621 (N_23621,N_17239,N_19701);
nor U23622 (N_23622,N_17709,N_17094);
or U23623 (N_23623,N_17823,N_16219);
and U23624 (N_23624,N_18723,N_17454);
nor U23625 (N_23625,N_19901,N_17318);
nand U23626 (N_23626,N_19325,N_15671);
and U23627 (N_23627,N_17684,N_17167);
and U23628 (N_23628,N_16011,N_19868);
and U23629 (N_23629,N_15649,N_19387);
xnor U23630 (N_23630,N_17663,N_18130);
and U23631 (N_23631,N_19417,N_15118);
nor U23632 (N_23632,N_16966,N_15839);
nor U23633 (N_23633,N_19714,N_18084);
xor U23634 (N_23634,N_17414,N_18300);
xor U23635 (N_23635,N_15881,N_17557);
and U23636 (N_23636,N_16071,N_16419);
nand U23637 (N_23637,N_18342,N_15538);
nor U23638 (N_23638,N_19078,N_17726);
and U23639 (N_23639,N_19270,N_18685);
nor U23640 (N_23640,N_15289,N_18247);
and U23641 (N_23641,N_19314,N_16124);
nor U23642 (N_23642,N_18248,N_16690);
and U23643 (N_23643,N_18036,N_17227);
or U23644 (N_23644,N_19821,N_17354);
nor U23645 (N_23645,N_15098,N_15353);
or U23646 (N_23646,N_18135,N_19890);
or U23647 (N_23647,N_15671,N_19507);
nand U23648 (N_23648,N_16814,N_16341);
and U23649 (N_23649,N_19893,N_19316);
nor U23650 (N_23650,N_16017,N_19236);
xor U23651 (N_23651,N_19523,N_19931);
or U23652 (N_23652,N_19919,N_17620);
and U23653 (N_23653,N_16931,N_19466);
nand U23654 (N_23654,N_15642,N_18308);
or U23655 (N_23655,N_16144,N_18693);
nor U23656 (N_23656,N_19553,N_17105);
and U23657 (N_23657,N_18757,N_18689);
nor U23658 (N_23658,N_17437,N_17573);
or U23659 (N_23659,N_15969,N_16851);
nor U23660 (N_23660,N_17732,N_18521);
or U23661 (N_23661,N_15722,N_17953);
nor U23662 (N_23662,N_19758,N_19128);
nor U23663 (N_23663,N_15693,N_16697);
nand U23664 (N_23664,N_17147,N_16279);
nand U23665 (N_23665,N_18943,N_17903);
and U23666 (N_23666,N_16387,N_19751);
or U23667 (N_23667,N_19822,N_19261);
xor U23668 (N_23668,N_18134,N_19098);
and U23669 (N_23669,N_17626,N_18777);
or U23670 (N_23670,N_17048,N_15245);
or U23671 (N_23671,N_15553,N_18427);
or U23672 (N_23672,N_15442,N_17614);
or U23673 (N_23673,N_16430,N_15375);
and U23674 (N_23674,N_19172,N_19519);
or U23675 (N_23675,N_19069,N_15073);
and U23676 (N_23676,N_16942,N_17892);
or U23677 (N_23677,N_19371,N_18746);
xnor U23678 (N_23678,N_17724,N_16138);
or U23679 (N_23679,N_16244,N_17574);
and U23680 (N_23680,N_17340,N_15308);
nor U23681 (N_23681,N_19355,N_17939);
and U23682 (N_23682,N_19269,N_18718);
nor U23683 (N_23683,N_17928,N_16570);
or U23684 (N_23684,N_15840,N_15142);
or U23685 (N_23685,N_16138,N_16129);
and U23686 (N_23686,N_18337,N_18208);
or U23687 (N_23687,N_18576,N_16891);
and U23688 (N_23688,N_17215,N_17763);
xor U23689 (N_23689,N_19997,N_18667);
and U23690 (N_23690,N_15161,N_15993);
xnor U23691 (N_23691,N_15219,N_16654);
nand U23692 (N_23692,N_15804,N_16297);
xnor U23693 (N_23693,N_16870,N_16038);
nor U23694 (N_23694,N_17430,N_16660);
and U23695 (N_23695,N_16228,N_19366);
and U23696 (N_23696,N_16949,N_15898);
or U23697 (N_23697,N_15490,N_18000);
nor U23698 (N_23698,N_16414,N_17068);
or U23699 (N_23699,N_15958,N_15107);
nand U23700 (N_23700,N_18854,N_16025);
and U23701 (N_23701,N_15628,N_16871);
nand U23702 (N_23702,N_15519,N_15786);
or U23703 (N_23703,N_17443,N_15745);
xor U23704 (N_23704,N_17558,N_19811);
nor U23705 (N_23705,N_15898,N_15655);
and U23706 (N_23706,N_18057,N_19962);
and U23707 (N_23707,N_19871,N_17003);
nor U23708 (N_23708,N_15341,N_15559);
and U23709 (N_23709,N_15278,N_16515);
nor U23710 (N_23710,N_15669,N_19143);
and U23711 (N_23711,N_19636,N_19218);
or U23712 (N_23712,N_17184,N_16891);
and U23713 (N_23713,N_19940,N_17169);
nor U23714 (N_23714,N_15507,N_15940);
or U23715 (N_23715,N_16580,N_15145);
nand U23716 (N_23716,N_17023,N_17974);
and U23717 (N_23717,N_15086,N_18922);
or U23718 (N_23718,N_16330,N_17326);
and U23719 (N_23719,N_16707,N_17233);
or U23720 (N_23720,N_15911,N_17398);
nor U23721 (N_23721,N_16175,N_19485);
or U23722 (N_23722,N_16508,N_19202);
nand U23723 (N_23723,N_18655,N_18185);
or U23724 (N_23724,N_15455,N_17725);
and U23725 (N_23725,N_17747,N_19736);
or U23726 (N_23726,N_16854,N_17652);
nand U23727 (N_23727,N_18905,N_18497);
nand U23728 (N_23728,N_19296,N_19374);
nor U23729 (N_23729,N_18506,N_16765);
xor U23730 (N_23730,N_17955,N_17176);
nor U23731 (N_23731,N_17991,N_16727);
nor U23732 (N_23732,N_15665,N_16873);
nor U23733 (N_23733,N_18102,N_17861);
or U23734 (N_23734,N_19934,N_16691);
or U23735 (N_23735,N_15249,N_15808);
or U23736 (N_23736,N_17893,N_19321);
nand U23737 (N_23737,N_18101,N_16834);
nor U23738 (N_23738,N_17756,N_19487);
nand U23739 (N_23739,N_15586,N_16181);
xor U23740 (N_23740,N_15677,N_19889);
nand U23741 (N_23741,N_19926,N_17158);
or U23742 (N_23742,N_18063,N_18326);
xor U23743 (N_23743,N_16238,N_15532);
nor U23744 (N_23744,N_18137,N_18279);
nor U23745 (N_23745,N_18110,N_19487);
nor U23746 (N_23746,N_17045,N_19509);
nand U23747 (N_23747,N_16991,N_16575);
and U23748 (N_23748,N_19106,N_15617);
or U23749 (N_23749,N_18047,N_15230);
and U23750 (N_23750,N_18372,N_16828);
nand U23751 (N_23751,N_19159,N_16187);
or U23752 (N_23752,N_16928,N_15368);
and U23753 (N_23753,N_16587,N_19021);
or U23754 (N_23754,N_15443,N_18952);
or U23755 (N_23755,N_17029,N_16288);
or U23756 (N_23756,N_16771,N_18895);
and U23757 (N_23757,N_15695,N_18786);
nand U23758 (N_23758,N_16134,N_17198);
and U23759 (N_23759,N_18148,N_19644);
nor U23760 (N_23760,N_16036,N_18175);
nand U23761 (N_23761,N_15527,N_16405);
xnor U23762 (N_23762,N_19641,N_15235);
nor U23763 (N_23763,N_17185,N_16341);
or U23764 (N_23764,N_16384,N_17931);
nand U23765 (N_23765,N_15353,N_18203);
nor U23766 (N_23766,N_16511,N_19562);
or U23767 (N_23767,N_16823,N_16888);
or U23768 (N_23768,N_17325,N_18115);
or U23769 (N_23769,N_19671,N_16713);
or U23770 (N_23770,N_16035,N_15732);
nor U23771 (N_23771,N_19905,N_17468);
or U23772 (N_23772,N_18457,N_16230);
or U23773 (N_23773,N_15270,N_18693);
xor U23774 (N_23774,N_15124,N_17109);
and U23775 (N_23775,N_18515,N_16478);
or U23776 (N_23776,N_17395,N_18425);
nand U23777 (N_23777,N_16081,N_16578);
and U23778 (N_23778,N_19686,N_19240);
nand U23779 (N_23779,N_15290,N_16797);
nor U23780 (N_23780,N_15157,N_16085);
or U23781 (N_23781,N_17969,N_19015);
nand U23782 (N_23782,N_18939,N_19632);
and U23783 (N_23783,N_15923,N_19588);
nand U23784 (N_23784,N_16019,N_15397);
and U23785 (N_23785,N_18102,N_15842);
nand U23786 (N_23786,N_15535,N_18294);
nand U23787 (N_23787,N_19476,N_16133);
nor U23788 (N_23788,N_15586,N_17979);
xnor U23789 (N_23789,N_19185,N_16513);
nor U23790 (N_23790,N_16229,N_15018);
or U23791 (N_23791,N_17036,N_17670);
or U23792 (N_23792,N_18447,N_18824);
nor U23793 (N_23793,N_19899,N_16749);
nor U23794 (N_23794,N_18692,N_16190);
nand U23795 (N_23795,N_17272,N_18189);
nor U23796 (N_23796,N_18333,N_17864);
and U23797 (N_23797,N_15641,N_15619);
nand U23798 (N_23798,N_17393,N_17002);
nand U23799 (N_23799,N_18426,N_16241);
xnor U23800 (N_23800,N_15571,N_19599);
or U23801 (N_23801,N_16289,N_15619);
nor U23802 (N_23802,N_15651,N_16575);
nand U23803 (N_23803,N_17848,N_15150);
nor U23804 (N_23804,N_19703,N_18607);
nor U23805 (N_23805,N_15672,N_19695);
or U23806 (N_23806,N_19257,N_16103);
or U23807 (N_23807,N_18361,N_18304);
xnor U23808 (N_23808,N_16635,N_19739);
or U23809 (N_23809,N_15108,N_15331);
nand U23810 (N_23810,N_18127,N_19373);
nor U23811 (N_23811,N_17900,N_18784);
nand U23812 (N_23812,N_19774,N_19782);
or U23813 (N_23813,N_19103,N_15966);
xor U23814 (N_23814,N_15376,N_18425);
nor U23815 (N_23815,N_18641,N_17769);
and U23816 (N_23816,N_19649,N_18273);
and U23817 (N_23817,N_18666,N_15197);
nor U23818 (N_23818,N_16392,N_15183);
xor U23819 (N_23819,N_18383,N_15976);
or U23820 (N_23820,N_17982,N_16204);
nor U23821 (N_23821,N_16351,N_16733);
and U23822 (N_23822,N_15999,N_15606);
nor U23823 (N_23823,N_19215,N_18198);
nand U23824 (N_23824,N_17790,N_19346);
or U23825 (N_23825,N_19411,N_16323);
nor U23826 (N_23826,N_15228,N_16220);
nor U23827 (N_23827,N_17248,N_16251);
nand U23828 (N_23828,N_19405,N_18968);
or U23829 (N_23829,N_15791,N_16507);
or U23830 (N_23830,N_18873,N_17245);
nand U23831 (N_23831,N_17170,N_15723);
nor U23832 (N_23832,N_19349,N_19906);
nand U23833 (N_23833,N_19246,N_16169);
nor U23834 (N_23834,N_18387,N_15388);
nand U23835 (N_23835,N_19865,N_18519);
nor U23836 (N_23836,N_16574,N_18494);
or U23837 (N_23837,N_18260,N_16015);
xnor U23838 (N_23838,N_18012,N_19372);
and U23839 (N_23839,N_17092,N_17511);
and U23840 (N_23840,N_19737,N_15189);
nor U23841 (N_23841,N_15156,N_17118);
nor U23842 (N_23842,N_15051,N_18376);
xor U23843 (N_23843,N_16896,N_17654);
and U23844 (N_23844,N_16020,N_16398);
or U23845 (N_23845,N_17818,N_16338);
nand U23846 (N_23846,N_18583,N_15931);
nand U23847 (N_23847,N_18260,N_17529);
and U23848 (N_23848,N_15190,N_19116);
and U23849 (N_23849,N_19301,N_17134);
or U23850 (N_23850,N_16633,N_16939);
nor U23851 (N_23851,N_16573,N_17678);
xnor U23852 (N_23852,N_16624,N_16579);
nor U23853 (N_23853,N_19340,N_16709);
and U23854 (N_23854,N_15828,N_16286);
and U23855 (N_23855,N_19949,N_16351);
nor U23856 (N_23856,N_15411,N_15982);
xor U23857 (N_23857,N_17029,N_17045);
nand U23858 (N_23858,N_17722,N_19445);
or U23859 (N_23859,N_15915,N_18668);
and U23860 (N_23860,N_17440,N_15925);
nor U23861 (N_23861,N_17284,N_16440);
or U23862 (N_23862,N_18849,N_17108);
and U23863 (N_23863,N_17741,N_17561);
and U23864 (N_23864,N_18819,N_15974);
nand U23865 (N_23865,N_17894,N_17531);
nor U23866 (N_23866,N_19299,N_16697);
or U23867 (N_23867,N_18088,N_17512);
nor U23868 (N_23868,N_15829,N_18759);
nor U23869 (N_23869,N_17959,N_17788);
nand U23870 (N_23870,N_16640,N_16716);
nand U23871 (N_23871,N_15734,N_15572);
or U23872 (N_23872,N_19753,N_15693);
and U23873 (N_23873,N_16346,N_15173);
or U23874 (N_23874,N_15587,N_18850);
xnor U23875 (N_23875,N_17490,N_15547);
or U23876 (N_23876,N_17565,N_19203);
nand U23877 (N_23877,N_18698,N_17863);
or U23878 (N_23878,N_16432,N_16135);
or U23879 (N_23879,N_19640,N_15239);
and U23880 (N_23880,N_19938,N_17303);
and U23881 (N_23881,N_17659,N_15862);
and U23882 (N_23882,N_18067,N_19062);
or U23883 (N_23883,N_19340,N_19859);
and U23884 (N_23884,N_17160,N_16053);
or U23885 (N_23885,N_16542,N_15013);
and U23886 (N_23886,N_18717,N_19463);
nor U23887 (N_23887,N_18650,N_17750);
xor U23888 (N_23888,N_17622,N_19077);
nor U23889 (N_23889,N_16868,N_17864);
nand U23890 (N_23890,N_18065,N_19795);
or U23891 (N_23891,N_16691,N_16660);
and U23892 (N_23892,N_15174,N_16375);
nor U23893 (N_23893,N_16331,N_19820);
or U23894 (N_23894,N_18126,N_16327);
and U23895 (N_23895,N_17818,N_15288);
nor U23896 (N_23896,N_15131,N_17119);
or U23897 (N_23897,N_17407,N_15035);
and U23898 (N_23898,N_15077,N_15006);
nor U23899 (N_23899,N_19674,N_17469);
nand U23900 (N_23900,N_18440,N_19224);
nand U23901 (N_23901,N_16024,N_18960);
nand U23902 (N_23902,N_15990,N_16512);
nor U23903 (N_23903,N_18641,N_18969);
nor U23904 (N_23904,N_15352,N_19675);
nand U23905 (N_23905,N_15825,N_17037);
nor U23906 (N_23906,N_17119,N_16912);
and U23907 (N_23907,N_19199,N_16346);
nor U23908 (N_23908,N_19408,N_18945);
nor U23909 (N_23909,N_19376,N_16885);
nor U23910 (N_23910,N_19170,N_17671);
nand U23911 (N_23911,N_17379,N_15008);
or U23912 (N_23912,N_18802,N_17806);
nand U23913 (N_23913,N_16308,N_16516);
nor U23914 (N_23914,N_16701,N_18185);
nor U23915 (N_23915,N_18750,N_19889);
nand U23916 (N_23916,N_18321,N_16970);
nor U23917 (N_23917,N_15476,N_16714);
and U23918 (N_23918,N_17306,N_19072);
or U23919 (N_23919,N_17570,N_15134);
and U23920 (N_23920,N_15956,N_16972);
and U23921 (N_23921,N_18760,N_16587);
xor U23922 (N_23922,N_16227,N_18481);
nor U23923 (N_23923,N_15319,N_16264);
xor U23924 (N_23924,N_18150,N_15430);
or U23925 (N_23925,N_19037,N_18113);
nand U23926 (N_23926,N_17237,N_18547);
and U23927 (N_23927,N_17052,N_18543);
nand U23928 (N_23928,N_15859,N_17966);
nand U23929 (N_23929,N_16965,N_16895);
nand U23930 (N_23930,N_15372,N_19820);
nand U23931 (N_23931,N_18352,N_15303);
or U23932 (N_23932,N_17616,N_18855);
xnor U23933 (N_23933,N_17676,N_15126);
or U23934 (N_23934,N_18274,N_18482);
nand U23935 (N_23935,N_17148,N_19902);
nand U23936 (N_23936,N_17315,N_18887);
or U23937 (N_23937,N_18103,N_15805);
or U23938 (N_23938,N_18978,N_19964);
nor U23939 (N_23939,N_16465,N_18435);
nor U23940 (N_23940,N_18409,N_19460);
and U23941 (N_23941,N_15737,N_19018);
or U23942 (N_23942,N_15030,N_17583);
or U23943 (N_23943,N_17302,N_16422);
nor U23944 (N_23944,N_18680,N_19681);
nor U23945 (N_23945,N_17650,N_18039);
and U23946 (N_23946,N_15622,N_18855);
and U23947 (N_23947,N_19719,N_18802);
and U23948 (N_23948,N_16079,N_17100);
nand U23949 (N_23949,N_16226,N_19389);
nor U23950 (N_23950,N_17863,N_18613);
xor U23951 (N_23951,N_15626,N_15977);
and U23952 (N_23952,N_15502,N_19721);
nor U23953 (N_23953,N_15075,N_17752);
and U23954 (N_23954,N_16622,N_18616);
nand U23955 (N_23955,N_18260,N_19435);
nand U23956 (N_23956,N_17704,N_18628);
nand U23957 (N_23957,N_15169,N_15638);
nor U23958 (N_23958,N_19168,N_15678);
nand U23959 (N_23959,N_18561,N_17054);
nand U23960 (N_23960,N_16837,N_18847);
nand U23961 (N_23961,N_17517,N_17276);
and U23962 (N_23962,N_18976,N_16277);
xnor U23963 (N_23963,N_18046,N_18346);
nor U23964 (N_23964,N_19185,N_17556);
and U23965 (N_23965,N_15943,N_16472);
nand U23966 (N_23966,N_16323,N_16114);
or U23967 (N_23967,N_15656,N_17438);
and U23968 (N_23968,N_17496,N_15291);
nor U23969 (N_23969,N_17728,N_19874);
nand U23970 (N_23970,N_15492,N_15008);
and U23971 (N_23971,N_17317,N_19720);
or U23972 (N_23972,N_19326,N_18886);
nand U23973 (N_23973,N_15153,N_19560);
nand U23974 (N_23974,N_17023,N_16018);
nand U23975 (N_23975,N_16401,N_15407);
and U23976 (N_23976,N_18587,N_15239);
nand U23977 (N_23977,N_19449,N_18930);
or U23978 (N_23978,N_19954,N_18092);
nand U23979 (N_23979,N_17060,N_17664);
or U23980 (N_23980,N_19545,N_18934);
nand U23981 (N_23981,N_18126,N_17418);
nand U23982 (N_23982,N_15586,N_15805);
and U23983 (N_23983,N_19891,N_17834);
nand U23984 (N_23984,N_18375,N_17340);
and U23985 (N_23985,N_19734,N_16938);
and U23986 (N_23986,N_15964,N_18392);
nand U23987 (N_23987,N_18333,N_16434);
and U23988 (N_23988,N_16168,N_16111);
and U23989 (N_23989,N_16461,N_18037);
nor U23990 (N_23990,N_17860,N_19358);
nand U23991 (N_23991,N_19836,N_15236);
or U23992 (N_23992,N_15914,N_18289);
nor U23993 (N_23993,N_16361,N_15691);
xnor U23994 (N_23994,N_15502,N_15923);
and U23995 (N_23995,N_15789,N_15595);
and U23996 (N_23996,N_18177,N_17611);
nand U23997 (N_23997,N_17875,N_17808);
nand U23998 (N_23998,N_16739,N_15080);
and U23999 (N_23999,N_16704,N_15590);
or U24000 (N_24000,N_18058,N_15051);
nor U24001 (N_24001,N_19060,N_19157);
nor U24002 (N_24002,N_18451,N_15953);
nor U24003 (N_24003,N_18678,N_16417);
xor U24004 (N_24004,N_15366,N_19591);
and U24005 (N_24005,N_15986,N_18577);
nor U24006 (N_24006,N_15921,N_15085);
nor U24007 (N_24007,N_17002,N_18577);
and U24008 (N_24008,N_17200,N_17664);
nand U24009 (N_24009,N_17511,N_17538);
nand U24010 (N_24010,N_17977,N_18542);
nor U24011 (N_24011,N_17253,N_18195);
or U24012 (N_24012,N_16005,N_15581);
and U24013 (N_24013,N_19294,N_18710);
and U24014 (N_24014,N_17098,N_15034);
nand U24015 (N_24015,N_15273,N_16673);
or U24016 (N_24016,N_16518,N_19577);
and U24017 (N_24017,N_18910,N_17790);
and U24018 (N_24018,N_15122,N_16382);
or U24019 (N_24019,N_17765,N_15601);
nand U24020 (N_24020,N_19655,N_15886);
and U24021 (N_24021,N_18993,N_18901);
nor U24022 (N_24022,N_18844,N_17738);
or U24023 (N_24023,N_19180,N_19098);
nand U24024 (N_24024,N_17979,N_18661);
and U24025 (N_24025,N_16065,N_16096);
and U24026 (N_24026,N_18853,N_18618);
or U24027 (N_24027,N_15109,N_16863);
nand U24028 (N_24028,N_16109,N_17188);
nand U24029 (N_24029,N_15532,N_15209);
nand U24030 (N_24030,N_15072,N_15775);
nand U24031 (N_24031,N_18897,N_16798);
nand U24032 (N_24032,N_15004,N_18976);
nand U24033 (N_24033,N_15663,N_16088);
nor U24034 (N_24034,N_17984,N_17934);
nand U24035 (N_24035,N_15322,N_17809);
and U24036 (N_24036,N_18764,N_17171);
nand U24037 (N_24037,N_16324,N_16678);
nand U24038 (N_24038,N_19274,N_16759);
and U24039 (N_24039,N_17900,N_16292);
nor U24040 (N_24040,N_15431,N_16863);
xnor U24041 (N_24041,N_16697,N_17811);
or U24042 (N_24042,N_17280,N_16181);
or U24043 (N_24043,N_19018,N_15447);
nor U24044 (N_24044,N_17671,N_15932);
xor U24045 (N_24045,N_19443,N_19467);
or U24046 (N_24046,N_15260,N_15205);
and U24047 (N_24047,N_19479,N_18294);
nor U24048 (N_24048,N_16093,N_18784);
xor U24049 (N_24049,N_19454,N_17989);
and U24050 (N_24050,N_17981,N_18478);
xnor U24051 (N_24051,N_16586,N_16044);
and U24052 (N_24052,N_17372,N_18975);
and U24053 (N_24053,N_15645,N_16528);
and U24054 (N_24054,N_18705,N_17508);
xnor U24055 (N_24055,N_15929,N_19400);
or U24056 (N_24056,N_16644,N_18725);
or U24057 (N_24057,N_15239,N_17405);
nand U24058 (N_24058,N_15176,N_15920);
nor U24059 (N_24059,N_19851,N_18694);
nand U24060 (N_24060,N_16277,N_16082);
and U24061 (N_24061,N_15308,N_15045);
xnor U24062 (N_24062,N_15117,N_19163);
or U24063 (N_24063,N_19612,N_15109);
or U24064 (N_24064,N_17257,N_18637);
and U24065 (N_24065,N_17060,N_16862);
and U24066 (N_24066,N_18905,N_18042);
nand U24067 (N_24067,N_18605,N_19696);
nand U24068 (N_24068,N_18253,N_16796);
and U24069 (N_24069,N_19828,N_15763);
or U24070 (N_24070,N_19829,N_15392);
nor U24071 (N_24071,N_16831,N_17451);
nor U24072 (N_24072,N_18642,N_19292);
nor U24073 (N_24073,N_17231,N_18847);
nand U24074 (N_24074,N_17661,N_16160);
nor U24075 (N_24075,N_19805,N_19780);
nor U24076 (N_24076,N_17057,N_15922);
and U24077 (N_24077,N_15193,N_16506);
xnor U24078 (N_24078,N_19334,N_15682);
and U24079 (N_24079,N_18222,N_19020);
nor U24080 (N_24080,N_16305,N_16087);
and U24081 (N_24081,N_17433,N_18914);
nor U24082 (N_24082,N_17987,N_18480);
nor U24083 (N_24083,N_17306,N_18740);
nand U24084 (N_24084,N_15063,N_16195);
or U24085 (N_24085,N_15466,N_15452);
and U24086 (N_24086,N_16619,N_19324);
or U24087 (N_24087,N_19378,N_18601);
nand U24088 (N_24088,N_18621,N_19691);
or U24089 (N_24089,N_19382,N_18958);
nand U24090 (N_24090,N_18165,N_18012);
nor U24091 (N_24091,N_18353,N_15837);
nand U24092 (N_24092,N_18028,N_15631);
nor U24093 (N_24093,N_16468,N_17583);
nand U24094 (N_24094,N_19887,N_16452);
nor U24095 (N_24095,N_19459,N_17404);
xnor U24096 (N_24096,N_15031,N_17782);
and U24097 (N_24097,N_15201,N_16161);
and U24098 (N_24098,N_16345,N_18800);
nand U24099 (N_24099,N_15732,N_17658);
and U24100 (N_24100,N_16533,N_15338);
nand U24101 (N_24101,N_15365,N_18822);
xnor U24102 (N_24102,N_15993,N_19716);
and U24103 (N_24103,N_16359,N_19095);
nand U24104 (N_24104,N_19649,N_18926);
nor U24105 (N_24105,N_15412,N_16676);
or U24106 (N_24106,N_17402,N_16880);
nand U24107 (N_24107,N_18502,N_19702);
xnor U24108 (N_24108,N_15382,N_17017);
and U24109 (N_24109,N_18235,N_18100);
or U24110 (N_24110,N_19311,N_16214);
nand U24111 (N_24111,N_15054,N_18679);
or U24112 (N_24112,N_17967,N_15239);
or U24113 (N_24113,N_19823,N_19316);
or U24114 (N_24114,N_16660,N_17410);
nor U24115 (N_24115,N_17756,N_19225);
nand U24116 (N_24116,N_18908,N_17515);
or U24117 (N_24117,N_15606,N_17443);
xnor U24118 (N_24118,N_17866,N_16122);
nand U24119 (N_24119,N_19797,N_16692);
or U24120 (N_24120,N_17925,N_15954);
or U24121 (N_24121,N_16003,N_17717);
or U24122 (N_24122,N_19665,N_18738);
nor U24123 (N_24123,N_16329,N_19346);
or U24124 (N_24124,N_17860,N_17256);
nand U24125 (N_24125,N_15229,N_18647);
nor U24126 (N_24126,N_15718,N_18700);
and U24127 (N_24127,N_19640,N_18614);
and U24128 (N_24128,N_16553,N_16971);
nand U24129 (N_24129,N_17352,N_16016);
and U24130 (N_24130,N_18694,N_19791);
nand U24131 (N_24131,N_15454,N_18782);
or U24132 (N_24132,N_17403,N_17327);
and U24133 (N_24133,N_15084,N_18898);
or U24134 (N_24134,N_18209,N_17434);
or U24135 (N_24135,N_17488,N_18249);
or U24136 (N_24136,N_17312,N_18067);
nor U24137 (N_24137,N_16271,N_17709);
nand U24138 (N_24138,N_17838,N_19784);
and U24139 (N_24139,N_18588,N_18165);
and U24140 (N_24140,N_17350,N_19419);
nor U24141 (N_24141,N_17085,N_16114);
xnor U24142 (N_24142,N_18470,N_16472);
or U24143 (N_24143,N_15781,N_17299);
or U24144 (N_24144,N_15521,N_19754);
nand U24145 (N_24145,N_19263,N_16587);
or U24146 (N_24146,N_17360,N_19172);
nand U24147 (N_24147,N_16607,N_19491);
nor U24148 (N_24148,N_15300,N_19362);
xor U24149 (N_24149,N_15183,N_17649);
nand U24150 (N_24150,N_17377,N_17402);
or U24151 (N_24151,N_19603,N_16957);
xnor U24152 (N_24152,N_18415,N_18942);
or U24153 (N_24153,N_17887,N_19321);
nand U24154 (N_24154,N_15253,N_15104);
and U24155 (N_24155,N_17693,N_19258);
or U24156 (N_24156,N_18288,N_18373);
and U24157 (N_24157,N_17578,N_17055);
nor U24158 (N_24158,N_16285,N_16357);
nor U24159 (N_24159,N_17652,N_15662);
and U24160 (N_24160,N_19673,N_16920);
nor U24161 (N_24161,N_15385,N_15511);
or U24162 (N_24162,N_16809,N_17253);
nand U24163 (N_24163,N_15713,N_15281);
nor U24164 (N_24164,N_19389,N_16851);
nand U24165 (N_24165,N_19806,N_19024);
or U24166 (N_24166,N_17820,N_15869);
nor U24167 (N_24167,N_19645,N_19529);
nand U24168 (N_24168,N_16940,N_18943);
and U24169 (N_24169,N_17314,N_15562);
nand U24170 (N_24170,N_18458,N_16757);
xor U24171 (N_24171,N_17329,N_15722);
and U24172 (N_24172,N_18434,N_17268);
nand U24173 (N_24173,N_18689,N_15787);
nor U24174 (N_24174,N_16000,N_15801);
and U24175 (N_24175,N_15823,N_18426);
and U24176 (N_24176,N_16690,N_15368);
nand U24177 (N_24177,N_15648,N_18308);
nor U24178 (N_24178,N_17217,N_15470);
and U24179 (N_24179,N_18521,N_15420);
nand U24180 (N_24180,N_16371,N_19829);
nand U24181 (N_24181,N_16073,N_17356);
nor U24182 (N_24182,N_15932,N_16253);
and U24183 (N_24183,N_19793,N_17213);
nor U24184 (N_24184,N_19884,N_16293);
or U24185 (N_24185,N_15072,N_18497);
or U24186 (N_24186,N_18693,N_16990);
nand U24187 (N_24187,N_19725,N_17946);
nor U24188 (N_24188,N_16913,N_16507);
or U24189 (N_24189,N_15300,N_19540);
or U24190 (N_24190,N_18636,N_19397);
nand U24191 (N_24191,N_17007,N_16854);
nor U24192 (N_24192,N_16569,N_19349);
nor U24193 (N_24193,N_17479,N_19571);
or U24194 (N_24194,N_16389,N_15604);
nand U24195 (N_24195,N_18526,N_18965);
nor U24196 (N_24196,N_15425,N_15206);
nor U24197 (N_24197,N_18756,N_18318);
nor U24198 (N_24198,N_17740,N_15515);
and U24199 (N_24199,N_15579,N_16550);
or U24200 (N_24200,N_16017,N_16927);
xnor U24201 (N_24201,N_16493,N_19821);
nor U24202 (N_24202,N_18228,N_17327);
and U24203 (N_24203,N_17105,N_19924);
or U24204 (N_24204,N_18082,N_15757);
or U24205 (N_24205,N_18949,N_15277);
nand U24206 (N_24206,N_17750,N_17045);
nand U24207 (N_24207,N_17878,N_18384);
nand U24208 (N_24208,N_16434,N_16894);
or U24209 (N_24209,N_17286,N_15123);
nor U24210 (N_24210,N_16808,N_19413);
nor U24211 (N_24211,N_15331,N_19157);
nand U24212 (N_24212,N_16583,N_16756);
nand U24213 (N_24213,N_17101,N_19328);
nor U24214 (N_24214,N_18337,N_15396);
nor U24215 (N_24215,N_17046,N_17921);
nor U24216 (N_24216,N_18779,N_16102);
nor U24217 (N_24217,N_15257,N_19724);
nor U24218 (N_24218,N_17686,N_17552);
nor U24219 (N_24219,N_17481,N_16710);
and U24220 (N_24220,N_15950,N_18959);
and U24221 (N_24221,N_17439,N_19861);
or U24222 (N_24222,N_15721,N_18480);
and U24223 (N_24223,N_16836,N_17795);
or U24224 (N_24224,N_18510,N_17532);
or U24225 (N_24225,N_15096,N_18026);
nand U24226 (N_24226,N_17892,N_19005);
nor U24227 (N_24227,N_19303,N_18364);
or U24228 (N_24228,N_15425,N_19524);
nand U24229 (N_24229,N_18663,N_19024);
nor U24230 (N_24230,N_18999,N_16560);
nand U24231 (N_24231,N_18676,N_15626);
or U24232 (N_24232,N_15050,N_19509);
xnor U24233 (N_24233,N_18813,N_17059);
nand U24234 (N_24234,N_19971,N_15404);
or U24235 (N_24235,N_16644,N_15395);
nand U24236 (N_24236,N_18807,N_16713);
nand U24237 (N_24237,N_18766,N_18322);
or U24238 (N_24238,N_16483,N_18793);
or U24239 (N_24239,N_19329,N_17183);
or U24240 (N_24240,N_17298,N_18686);
nand U24241 (N_24241,N_17847,N_19078);
nor U24242 (N_24242,N_16706,N_17280);
and U24243 (N_24243,N_18157,N_18921);
nand U24244 (N_24244,N_17798,N_16335);
xnor U24245 (N_24245,N_17365,N_17009);
and U24246 (N_24246,N_16545,N_18142);
nor U24247 (N_24247,N_16578,N_15211);
and U24248 (N_24248,N_17074,N_16197);
nand U24249 (N_24249,N_16028,N_18693);
and U24250 (N_24250,N_19315,N_19003);
nor U24251 (N_24251,N_16005,N_19057);
and U24252 (N_24252,N_19803,N_17394);
and U24253 (N_24253,N_17183,N_16568);
nor U24254 (N_24254,N_18071,N_16205);
nor U24255 (N_24255,N_17255,N_17825);
and U24256 (N_24256,N_19298,N_15877);
nand U24257 (N_24257,N_16676,N_18734);
nand U24258 (N_24258,N_15908,N_19067);
nor U24259 (N_24259,N_17106,N_16647);
and U24260 (N_24260,N_16199,N_19449);
nand U24261 (N_24261,N_17222,N_18535);
or U24262 (N_24262,N_19045,N_15068);
and U24263 (N_24263,N_15913,N_19914);
nand U24264 (N_24264,N_19111,N_16958);
and U24265 (N_24265,N_19295,N_15777);
nand U24266 (N_24266,N_16955,N_18910);
and U24267 (N_24267,N_15238,N_18765);
nor U24268 (N_24268,N_15987,N_19193);
and U24269 (N_24269,N_19864,N_16874);
or U24270 (N_24270,N_16361,N_16109);
nor U24271 (N_24271,N_18997,N_18880);
nand U24272 (N_24272,N_17980,N_18023);
xor U24273 (N_24273,N_16600,N_15941);
and U24274 (N_24274,N_16433,N_19293);
nor U24275 (N_24275,N_15024,N_19422);
nor U24276 (N_24276,N_18143,N_17378);
nor U24277 (N_24277,N_19673,N_17298);
nand U24278 (N_24278,N_18242,N_16636);
or U24279 (N_24279,N_15228,N_15046);
or U24280 (N_24280,N_19848,N_18157);
nand U24281 (N_24281,N_17454,N_17456);
or U24282 (N_24282,N_17236,N_16205);
or U24283 (N_24283,N_18053,N_17236);
or U24284 (N_24284,N_19778,N_19049);
and U24285 (N_24285,N_15377,N_15981);
nand U24286 (N_24286,N_17073,N_18502);
nor U24287 (N_24287,N_15430,N_15802);
xnor U24288 (N_24288,N_17390,N_15020);
nand U24289 (N_24289,N_15539,N_19181);
nor U24290 (N_24290,N_18165,N_16149);
and U24291 (N_24291,N_17572,N_16000);
or U24292 (N_24292,N_19652,N_16470);
nand U24293 (N_24293,N_16684,N_19537);
or U24294 (N_24294,N_19767,N_18774);
nand U24295 (N_24295,N_16312,N_18357);
nand U24296 (N_24296,N_17227,N_18391);
or U24297 (N_24297,N_15994,N_15168);
nand U24298 (N_24298,N_17040,N_15345);
nor U24299 (N_24299,N_15666,N_19795);
nand U24300 (N_24300,N_16228,N_18950);
and U24301 (N_24301,N_16361,N_15946);
nand U24302 (N_24302,N_15065,N_15594);
nand U24303 (N_24303,N_17027,N_16678);
and U24304 (N_24304,N_19278,N_15437);
or U24305 (N_24305,N_18948,N_18335);
nor U24306 (N_24306,N_16881,N_19114);
and U24307 (N_24307,N_18721,N_19359);
nand U24308 (N_24308,N_16212,N_16432);
xor U24309 (N_24309,N_17648,N_18255);
nand U24310 (N_24310,N_18730,N_17645);
nand U24311 (N_24311,N_16075,N_15474);
and U24312 (N_24312,N_17805,N_15030);
nand U24313 (N_24313,N_18703,N_18110);
nand U24314 (N_24314,N_19664,N_16938);
nand U24315 (N_24315,N_16967,N_17424);
or U24316 (N_24316,N_16778,N_16835);
nand U24317 (N_24317,N_18909,N_16966);
or U24318 (N_24318,N_17287,N_15877);
and U24319 (N_24319,N_17643,N_18731);
xnor U24320 (N_24320,N_18969,N_19606);
nor U24321 (N_24321,N_19447,N_18668);
nand U24322 (N_24322,N_18508,N_16969);
and U24323 (N_24323,N_16088,N_16434);
nand U24324 (N_24324,N_17097,N_18389);
and U24325 (N_24325,N_15720,N_19923);
nor U24326 (N_24326,N_17696,N_18218);
nor U24327 (N_24327,N_18105,N_16789);
and U24328 (N_24328,N_15171,N_19840);
and U24329 (N_24329,N_16113,N_17114);
and U24330 (N_24330,N_15268,N_15454);
or U24331 (N_24331,N_18307,N_15448);
and U24332 (N_24332,N_16565,N_16241);
and U24333 (N_24333,N_18484,N_15217);
nand U24334 (N_24334,N_16917,N_15896);
xnor U24335 (N_24335,N_16462,N_15289);
nand U24336 (N_24336,N_16690,N_17484);
nand U24337 (N_24337,N_15252,N_15640);
nor U24338 (N_24338,N_17703,N_19395);
or U24339 (N_24339,N_18545,N_16831);
and U24340 (N_24340,N_16552,N_19424);
and U24341 (N_24341,N_15887,N_16080);
xnor U24342 (N_24342,N_17503,N_17182);
or U24343 (N_24343,N_15862,N_17109);
or U24344 (N_24344,N_16753,N_17529);
and U24345 (N_24345,N_17295,N_15281);
and U24346 (N_24346,N_18548,N_16049);
and U24347 (N_24347,N_15490,N_17985);
nand U24348 (N_24348,N_19083,N_16170);
and U24349 (N_24349,N_16293,N_17031);
nand U24350 (N_24350,N_15200,N_17037);
or U24351 (N_24351,N_18802,N_17506);
nor U24352 (N_24352,N_18371,N_19990);
nand U24353 (N_24353,N_19668,N_16233);
nand U24354 (N_24354,N_16815,N_16939);
or U24355 (N_24355,N_18115,N_16862);
or U24356 (N_24356,N_15183,N_16099);
xnor U24357 (N_24357,N_16289,N_15557);
nor U24358 (N_24358,N_17558,N_15724);
or U24359 (N_24359,N_18260,N_15893);
or U24360 (N_24360,N_19626,N_19874);
and U24361 (N_24361,N_17847,N_15664);
xor U24362 (N_24362,N_17522,N_15230);
or U24363 (N_24363,N_18715,N_16578);
nor U24364 (N_24364,N_19005,N_15396);
nor U24365 (N_24365,N_17745,N_19615);
nand U24366 (N_24366,N_17138,N_15313);
xnor U24367 (N_24367,N_16560,N_16365);
nor U24368 (N_24368,N_16952,N_17199);
and U24369 (N_24369,N_18863,N_16650);
nor U24370 (N_24370,N_15905,N_18034);
or U24371 (N_24371,N_18945,N_15874);
nand U24372 (N_24372,N_18500,N_15059);
nor U24373 (N_24373,N_15286,N_15343);
or U24374 (N_24374,N_19186,N_15324);
or U24375 (N_24375,N_16500,N_16660);
and U24376 (N_24376,N_19588,N_15817);
or U24377 (N_24377,N_15728,N_15007);
and U24378 (N_24378,N_15137,N_17300);
nor U24379 (N_24379,N_19563,N_17239);
nand U24380 (N_24380,N_19123,N_16251);
or U24381 (N_24381,N_18505,N_19324);
nor U24382 (N_24382,N_15671,N_19065);
and U24383 (N_24383,N_15682,N_17529);
nor U24384 (N_24384,N_19007,N_15187);
or U24385 (N_24385,N_16871,N_17069);
or U24386 (N_24386,N_16750,N_15187);
xor U24387 (N_24387,N_16221,N_15356);
xnor U24388 (N_24388,N_17138,N_18971);
nand U24389 (N_24389,N_16767,N_18599);
nor U24390 (N_24390,N_17818,N_19972);
and U24391 (N_24391,N_17452,N_17876);
xor U24392 (N_24392,N_16837,N_18183);
or U24393 (N_24393,N_16310,N_16269);
and U24394 (N_24394,N_16706,N_17176);
and U24395 (N_24395,N_19365,N_19697);
xor U24396 (N_24396,N_16617,N_17532);
nand U24397 (N_24397,N_16247,N_19923);
nor U24398 (N_24398,N_18162,N_15499);
xor U24399 (N_24399,N_18171,N_18322);
or U24400 (N_24400,N_18492,N_17171);
or U24401 (N_24401,N_18375,N_18082);
or U24402 (N_24402,N_18725,N_18671);
nor U24403 (N_24403,N_19904,N_17292);
nor U24404 (N_24404,N_17252,N_15210);
nor U24405 (N_24405,N_18074,N_15840);
xnor U24406 (N_24406,N_17788,N_18062);
nand U24407 (N_24407,N_15328,N_17275);
nand U24408 (N_24408,N_16473,N_16521);
nand U24409 (N_24409,N_17298,N_18320);
nor U24410 (N_24410,N_19182,N_18587);
and U24411 (N_24411,N_17674,N_19482);
and U24412 (N_24412,N_17768,N_15404);
nand U24413 (N_24413,N_16989,N_17000);
nand U24414 (N_24414,N_18760,N_19161);
nor U24415 (N_24415,N_19516,N_16987);
and U24416 (N_24416,N_18565,N_18262);
and U24417 (N_24417,N_19649,N_16975);
or U24418 (N_24418,N_17444,N_16697);
nand U24419 (N_24419,N_18877,N_15818);
or U24420 (N_24420,N_19893,N_18443);
nor U24421 (N_24421,N_17948,N_17077);
or U24422 (N_24422,N_17063,N_16952);
and U24423 (N_24423,N_16865,N_17153);
or U24424 (N_24424,N_17647,N_17040);
nor U24425 (N_24425,N_15305,N_18909);
nor U24426 (N_24426,N_15894,N_16556);
or U24427 (N_24427,N_16933,N_19419);
nand U24428 (N_24428,N_19558,N_15087);
or U24429 (N_24429,N_16620,N_19422);
nor U24430 (N_24430,N_18884,N_17285);
and U24431 (N_24431,N_19765,N_15416);
nand U24432 (N_24432,N_18574,N_16309);
xor U24433 (N_24433,N_18692,N_16310);
or U24434 (N_24434,N_18516,N_19459);
or U24435 (N_24435,N_18031,N_18476);
nand U24436 (N_24436,N_19800,N_19181);
nor U24437 (N_24437,N_17716,N_16525);
or U24438 (N_24438,N_17507,N_15979);
nand U24439 (N_24439,N_19575,N_16887);
nor U24440 (N_24440,N_15208,N_17931);
or U24441 (N_24441,N_17954,N_15509);
or U24442 (N_24442,N_16852,N_16734);
or U24443 (N_24443,N_15694,N_15336);
or U24444 (N_24444,N_19182,N_15000);
or U24445 (N_24445,N_17449,N_17366);
or U24446 (N_24446,N_17669,N_17751);
nor U24447 (N_24447,N_16421,N_15781);
and U24448 (N_24448,N_16027,N_16613);
and U24449 (N_24449,N_15580,N_18223);
nor U24450 (N_24450,N_19821,N_17534);
and U24451 (N_24451,N_16473,N_15994);
nand U24452 (N_24452,N_15017,N_16540);
xor U24453 (N_24453,N_19558,N_15040);
or U24454 (N_24454,N_19805,N_18448);
nand U24455 (N_24455,N_19321,N_18113);
nor U24456 (N_24456,N_15451,N_17574);
or U24457 (N_24457,N_15680,N_15942);
and U24458 (N_24458,N_15714,N_16847);
or U24459 (N_24459,N_15537,N_19861);
or U24460 (N_24460,N_18820,N_16337);
or U24461 (N_24461,N_17267,N_17252);
nand U24462 (N_24462,N_19434,N_18208);
nor U24463 (N_24463,N_19054,N_18959);
and U24464 (N_24464,N_18266,N_19247);
or U24465 (N_24465,N_15700,N_19944);
nor U24466 (N_24466,N_16715,N_15649);
or U24467 (N_24467,N_17850,N_17343);
or U24468 (N_24468,N_15520,N_19489);
nor U24469 (N_24469,N_19743,N_18994);
or U24470 (N_24470,N_18505,N_17187);
or U24471 (N_24471,N_17241,N_17254);
and U24472 (N_24472,N_18031,N_19125);
and U24473 (N_24473,N_19230,N_16299);
nor U24474 (N_24474,N_15554,N_17230);
or U24475 (N_24475,N_15346,N_19615);
and U24476 (N_24476,N_18532,N_18373);
and U24477 (N_24477,N_17456,N_15898);
or U24478 (N_24478,N_17723,N_18507);
nor U24479 (N_24479,N_18462,N_18303);
nand U24480 (N_24480,N_17701,N_15681);
or U24481 (N_24481,N_19032,N_17404);
and U24482 (N_24482,N_15935,N_15287);
nand U24483 (N_24483,N_17671,N_17888);
or U24484 (N_24484,N_18606,N_19433);
or U24485 (N_24485,N_17802,N_18242);
and U24486 (N_24486,N_19990,N_19562);
nand U24487 (N_24487,N_18887,N_17008);
nand U24488 (N_24488,N_18065,N_19575);
nor U24489 (N_24489,N_19951,N_16624);
and U24490 (N_24490,N_18072,N_17806);
nor U24491 (N_24491,N_17573,N_17254);
or U24492 (N_24492,N_15120,N_19394);
and U24493 (N_24493,N_19292,N_16893);
xnor U24494 (N_24494,N_15833,N_17399);
or U24495 (N_24495,N_17869,N_19977);
and U24496 (N_24496,N_15639,N_18146);
xor U24497 (N_24497,N_17243,N_15466);
xnor U24498 (N_24498,N_15594,N_18995);
nand U24499 (N_24499,N_16624,N_17972);
and U24500 (N_24500,N_19223,N_19677);
or U24501 (N_24501,N_16676,N_17347);
nor U24502 (N_24502,N_17092,N_19063);
and U24503 (N_24503,N_17701,N_17353);
nor U24504 (N_24504,N_15464,N_19924);
nand U24505 (N_24505,N_17906,N_18496);
or U24506 (N_24506,N_17565,N_19404);
nor U24507 (N_24507,N_16637,N_19064);
xor U24508 (N_24508,N_19792,N_17598);
nor U24509 (N_24509,N_17149,N_18754);
nand U24510 (N_24510,N_19222,N_19276);
and U24511 (N_24511,N_17770,N_19246);
and U24512 (N_24512,N_15651,N_19158);
xnor U24513 (N_24513,N_16986,N_15566);
xnor U24514 (N_24514,N_17917,N_18640);
nor U24515 (N_24515,N_15314,N_15101);
nor U24516 (N_24516,N_17834,N_18589);
and U24517 (N_24517,N_15494,N_17858);
nand U24518 (N_24518,N_19802,N_16514);
nor U24519 (N_24519,N_17624,N_15274);
or U24520 (N_24520,N_16301,N_15055);
nor U24521 (N_24521,N_17725,N_15170);
or U24522 (N_24522,N_16197,N_17970);
nor U24523 (N_24523,N_16078,N_16845);
xor U24524 (N_24524,N_16530,N_19687);
and U24525 (N_24525,N_19732,N_16456);
nor U24526 (N_24526,N_15589,N_16639);
or U24527 (N_24527,N_16968,N_18681);
and U24528 (N_24528,N_18259,N_15188);
xor U24529 (N_24529,N_15477,N_15985);
and U24530 (N_24530,N_19409,N_17914);
xor U24531 (N_24531,N_16265,N_18574);
nor U24532 (N_24532,N_16050,N_17107);
and U24533 (N_24533,N_19468,N_15594);
nand U24534 (N_24534,N_18684,N_19852);
and U24535 (N_24535,N_15329,N_18075);
nor U24536 (N_24536,N_19979,N_17126);
nand U24537 (N_24537,N_17693,N_17308);
and U24538 (N_24538,N_16060,N_17378);
or U24539 (N_24539,N_15187,N_18883);
nand U24540 (N_24540,N_18182,N_16579);
nand U24541 (N_24541,N_19684,N_19157);
xor U24542 (N_24542,N_19360,N_17878);
or U24543 (N_24543,N_18320,N_17673);
nand U24544 (N_24544,N_17828,N_17618);
xor U24545 (N_24545,N_18546,N_17348);
and U24546 (N_24546,N_19040,N_16492);
nand U24547 (N_24547,N_18761,N_19823);
nand U24548 (N_24548,N_18754,N_15607);
and U24549 (N_24549,N_15104,N_17436);
nor U24550 (N_24550,N_19786,N_15883);
or U24551 (N_24551,N_15298,N_19019);
xnor U24552 (N_24552,N_15716,N_16429);
or U24553 (N_24553,N_16105,N_15147);
or U24554 (N_24554,N_19857,N_18725);
or U24555 (N_24555,N_17640,N_18171);
or U24556 (N_24556,N_17383,N_16824);
and U24557 (N_24557,N_16432,N_16783);
nor U24558 (N_24558,N_18941,N_18578);
or U24559 (N_24559,N_18430,N_19686);
xor U24560 (N_24560,N_19407,N_15322);
nor U24561 (N_24561,N_18853,N_17518);
or U24562 (N_24562,N_18847,N_15501);
and U24563 (N_24563,N_15078,N_18368);
nor U24564 (N_24564,N_18689,N_15140);
nor U24565 (N_24565,N_17970,N_18346);
and U24566 (N_24566,N_16732,N_19385);
and U24567 (N_24567,N_17900,N_16422);
or U24568 (N_24568,N_16395,N_17601);
or U24569 (N_24569,N_19502,N_15437);
nor U24570 (N_24570,N_19781,N_15467);
nand U24571 (N_24571,N_19681,N_17847);
nor U24572 (N_24572,N_18704,N_18880);
or U24573 (N_24573,N_18051,N_18813);
nand U24574 (N_24574,N_19329,N_17663);
nand U24575 (N_24575,N_18672,N_15718);
and U24576 (N_24576,N_17352,N_19884);
or U24577 (N_24577,N_17346,N_19591);
nor U24578 (N_24578,N_18434,N_19608);
xor U24579 (N_24579,N_15424,N_17942);
xnor U24580 (N_24580,N_19568,N_18079);
nand U24581 (N_24581,N_17678,N_15733);
nor U24582 (N_24582,N_16673,N_16944);
nand U24583 (N_24583,N_19666,N_15060);
and U24584 (N_24584,N_17884,N_16286);
nor U24585 (N_24585,N_15003,N_16663);
or U24586 (N_24586,N_19132,N_16946);
and U24587 (N_24587,N_19631,N_18929);
nand U24588 (N_24588,N_16402,N_15412);
or U24589 (N_24589,N_17493,N_17590);
and U24590 (N_24590,N_17254,N_15908);
nor U24591 (N_24591,N_16984,N_16859);
nor U24592 (N_24592,N_15010,N_19455);
nor U24593 (N_24593,N_17246,N_16034);
and U24594 (N_24594,N_19212,N_18290);
nand U24595 (N_24595,N_19282,N_18132);
nor U24596 (N_24596,N_17517,N_18687);
and U24597 (N_24597,N_16616,N_15963);
or U24598 (N_24598,N_18134,N_16924);
nor U24599 (N_24599,N_16715,N_16697);
nand U24600 (N_24600,N_16004,N_18695);
nor U24601 (N_24601,N_16290,N_15374);
xor U24602 (N_24602,N_18969,N_17219);
and U24603 (N_24603,N_16848,N_15569);
xor U24604 (N_24604,N_19753,N_18760);
and U24605 (N_24605,N_16135,N_15590);
or U24606 (N_24606,N_15130,N_16259);
and U24607 (N_24607,N_17095,N_19992);
nor U24608 (N_24608,N_16238,N_15820);
and U24609 (N_24609,N_18600,N_16128);
nor U24610 (N_24610,N_16039,N_18427);
nor U24611 (N_24611,N_16910,N_19499);
nor U24612 (N_24612,N_17234,N_16352);
nand U24613 (N_24613,N_19993,N_18604);
nand U24614 (N_24614,N_16721,N_19533);
nor U24615 (N_24615,N_19868,N_16600);
nand U24616 (N_24616,N_17839,N_15939);
and U24617 (N_24617,N_17749,N_18754);
nand U24618 (N_24618,N_17387,N_17685);
and U24619 (N_24619,N_19208,N_16200);
or U24620 (N_24620,N_18807,N_17679);
or U24621 (N_24621,N_19640,N_18709);
nor U24622 (N_24622,N_19468,N_15827);
and U24623 (N_24623,N_17599,N_17021);
nand U24624 (N_24624,N_18718,N_18325);
or U24625 (N_24625,N_18224,N_15386);
nand U24626 (N_24626,N_16492,N_18778);
or U24627 (N_24627,N_16968,N_15504);
nor U24628 (N_24628,N_18120,N_15163);
xnor U24629 (N_24629,N_18033,N_16975);
nand U24630 (N_24630,N_17461,N_17626);
nor U24631 (N_24631,N_18609,N_18693);
nand U24632 (N_24632,N_19719,N_19416);
or U24633 (N_24633,N_18699,N_19310);
nor U24634 (N_24634,N_19264,N_19950);
or U24635 (N_24635,N_15235,N_15923);
and U24636 (N_24636,N_16741,N_18863);
and U24637 (N_24637,N_19570,N_15786);
and U24638 (N_24638,N_16962,N_16813);
or U24639 (N_24639,N_15278,N_16051);
and U24640 (N_24640,N_15706,N_15306);
nand U24641 (N_24641,N_16916,N_15086);
or U24642 (N_24642,N_18161,N_18872);
xnor U24643 (N_24643,N_17550,N_16738);
nand U24644 (N_24644,N_17818,N_16441);
nand U24645 (N_24645,N_15396,N_18136);
nor U24646 (N_24646,N_19621,N_17813);
nor U24647 (N_24647,N_16824,N_16775);
and U24648 (N_24648,N_15915,N_18349);
xor U24649 (N_24649,N_16674,N_19387);
or U24650 (N_24650,N_17314,N_15415);
nor U24651 (N_24651,N_17243,N_15014);
or U24652 (N_24652,N_18198,N_17530);
nor U24653 (N_24653,N_17586,N_18805);
or U24654 (N_24654,N_16495,N_15411);
xor U24655 (N_24655,N_15056,N_18972);
or U24656 (N_24656,N_19935,N_18839);
or U24657 (N_24657,N_18648,N_15972);
nand U24658 (N_24658,N_18786,N_17521);
nand U24659 (N_24659,N_17550,N_19890);
xor U24660 (N_24660,N_17834,N_15046);
nor U24661 (N_24661,N_18850,N_18505);
nor U24662 (N_24662,N_18419,N_17280);
nor U24663 (N_24663,N_16902,N_18661);
nand U24664 (N_24664,N_16639,N_17315);
nor U24665 (N_24665,N_17549,N_17443);
and U24666 (N_24666,N_15672,N_15531);
nor U24667 (N_24667,N_15891,N_19274);
xnor U24668 (N_24668,N_19864,N_15388);
nor U24669 (N_24669,N_16252,N_16452);
and U24670 (N_24670,N_19342,N_19505);
nand U24671 (N_24671,N_19567,N_17399);
or U24672 (N_24672,N_17288,N_18785);
nand U24673 (N_24673,N_18645,N_15202);
and U24674 (N_24674,N_16937,N_19196);
or U24675 (N_24675,N_17877,N_18318);
nor U24676 (N_24676,N_16068,N_18467);
nand U24677 (N_24677,N_19290,N_15127);
xor U24678 (N_24678,N_15334,N_18990);
nor U24679 (N_24679,N_15180,N_15884);
or U24680 (N_24680,N_15151,N_19464);
nand U24681 (N_24681,N_15543,N_16269);
xnor U24682 (N_24682,N_16329,N_19015);
or U24683 (N_24683,N_15951,N_18584);
nor U24684 (N_24684,N_18587,N_17721);
nand U24685 (N_24685,N_18765,N_19536);
and U24686 (N_24686,N_16465,N_19201);
nand U24687 (N_24687,N_15182,N_17455);
nor U24688 (N_24688,N_17636,N_17615);
and U24689 (N_24689,N_16210,N_19932);
nand U24690 (N_24690,N_16020,N_16326);
nor U24691 (N_24691,N_19084,N_19290);
xnor U24692 (N_24692,N_15999,N_15551);
nand U24693 (N_24693,N_15876,N_17959);
or U24694 (N_24694,N_16616,N_18160);
or U24695 (N_24695,N_18197,N_18811);
nand U24696 (N_24696,N_19278,N_15879);
or U24697 (N_24697,N_17458,N_17182);
and U24698 (N_24698,N_17353,N_16734);
nor U24699 (N_24699,N_16364,N_16961);
nand U24700 (N_24700,N_19286,N_18441);
nor U24701 (N_24701,N_15849,N_17537);
or U24702 (N_24702,N_16084,N_18451);
nand U24703 (N_24703,N_16048,N_19945);
nor U24704 (N_24704,N_18772,N_17829);
or U24705 (N_24705,N_17127,N_18899);
nand U24706 (N_24706,N_18332,N_19365);
nor U24707 (N_24707,N_17728,N_19329);
or U24708 (N_24708,N_17709,N_19185);
nor U24709 (N_24709,N_15466,N_19396);
and U24710 (N_24710,N_15035,N_18672);
or U24711 (N_24711,N_19548,N_15100);
xnor U24712 (N_24712,N_17528,N_15834);
nand U24713 (N_24713,N_17513,N_16264);
nand U24714 (N_24714,N_15050,N_17047);
and U24715 (N_24715,N_19309,N_15416);
xor U24716 (N_24716,N_18224,N_15866);
nand U24717 (N_24717,N_15430,N_19301);
nand U24718 (N_24718,N_16087,N_17918);
xor U24719 (N_24719,N_17186,N_17165);
or U24720 (N_24720,N_17958,N_15286);
and U24721 (N_24721,N_17957,N_17772);
xnor U24722 (N_24722,N_19920,N_15154);
nor U24723 (N_24723,N_17442,N_16248);
and U24724 (N_24724,N_17687,N_18972);
nor U24725 (N_24725,N_18973,N_15199);
nand U24726 (N_24726,N_15794,N_19979);
or U24727 (N_24727,N_17524,N_16566);
xor U24728 (N_24728,N_17043,N_18607);
and U24729 (N_24729,N_15715,N_18132);
nand U24730 (N_24730,N_16937,N_19263);
or U24731 (N_24731,N_19389,N_16203);
and U24732 (N_24732,N_19265,N_15203);
nand U24733 (N_24733,N_18609,N_16983);
nand U24734 (N_24734,N_15775,N_16077);
and U24735 (N_24735,N_18913,N_19264);
nor U24736 (N_24736,N_17082,N_15871);
and U24737 (N_24737,N_15734,N_19845);
nor U24738 (N_24738,N_17418,N_17192);
nand U24739 (N_24739,N_17436,N_16016);
or U24740 (N_24740,N_15125,N_16859);
nand U24741 (N_24741,N_17235,N_17137);
or U24742 (N_24742,N_15531,N_19121);
or U24743 (N_24743,N_19857,N_19492);
and U24744 (N_24744,N_15008,N_16556);
or U24745 (N_24745,N_19194,N_18498);
or U24746 (N_24746,N_19432,N_19522);
and U24747 (N_24747,N_15956,N_15933);
nor U24748 (N_24748,N_19124,N_16425);
nand U24749 (N_24749,N_15555,N_15535);
xor U24750 (N_24750,N_17185,N_17541);
and U24751 (N_24751,N_16657,N_18517);
or U24752 (N_24752,N_16191,N_15109);
or U24753 (N_24753,N_17808,N_17382);
and U24754 (N_24754,N_17397,N_15282);
nand U24755 (N_24755,N_15976,N_15062);
or U24756 (N_24756,N_15899,N_19207);
and U24757 (N_24757,N_16668,N_18242);
nand U24758 (N_24758,N_16831,N_17806);
and U24759 (N_24759,N_18366,N_15080);
or U24760 (N_24760,N_16702,N_16277);
xor U24761 (N_24761,N_17812,N_18802);
and U24762 (N_24762,N_15027,N_17690);
nand U24763 (N_24763,N_15976,N_19057);
nor U24764 (N_24764,N_17983,N_16997);
and U24765 (N_24765,N_16502,N_15589);
nor U24766 (N_24766,N_18826,N_19211);
nand U24767 (N_24767,N_19688,N_17510);
and U24768 (N_24768,N_19523,N_15458);
xor U24769 (N_24769,N_16285,N_19680);
and U24770 (N_24770,N_18914,N_15340);
and U24771 (N_24771,N_16578,N_18150);
and U24772 (N_24772,N_15349,N_18371);
or U24773 (N_24773,N_18660,N_18723);
and U24774 (N_24774,N_19542,N_19356);
nand U24775 (N_24775,N_18197,N_18356);
nor U24776 (N_24776,N_15827,N_19508);
xnor U24777 (N_24777,N_19833,N_15466);
or U24778 (N_24778,N_16258,N_15389);
xor U24779 (N_24779,N_18624,N_16249);
or U24780 (N_24780,N_18761,N_18580);
or U24781 (N_24781,N_15582,N_18490);
xnor U24782 (N_24782,N_17526,N_16908);
or U24783 (N_24783,N_18506,N_17142);
nand U24784 (N_24784,N_19518,N_19424);
or U24785 (N_24785,N_18615,N_18077);
xnor U24786 (N_24786,N_18297,N_15629);
or U24787 (N_24787,N_19267,N_18466);
xnor U24788 (N_24788,N_19364,N_18005);
or U24789 (N_24789,N_15794,N_18692);
or U24790 (N_24790,N_15016,N_18012);
xnor U24791 (N_24791,N_18032,N_16490);
nor U24792 (N_24792,N_18364,N_17220);
and U24793 (N_24793,N_16001,N_17271);
nor U24794 (N_24794,N_18999,N_17861);
and U24795 (N_24795,N_18705,N_19204);
nand U24796 (N_24796,N_16027,N_17688);
nor U24797 (N_24797,N_19575,N_18764);
and U24798 (N_24798,N_16964,N_16720);
nand U24799 (N_24799,N_18368,N_16145);
xor U24800 (N_24800,N_16091,N_18321);
nor U24801 (N_24801,N_18872,N_16430);
or U24802 (N_24802,N_18744,N_15321);
nor U24803 (N_24803,N_16619,N_17960);
nand U24804 (N_24804,N_16462,N_16308);
or U24805 (N_24805,N_18703,N_17195);
nand U24806 (N_24806,N_17816,N_18486);
nor U24807 (N_24807,N_15166,N_15753);
and U24808 (N_24808,N_17567,N_15772);
nand U24809 (N_24809,N_16929,N_15673);
or U24810 (N_24810,N_19049,N_17047);
and U24811 (N_24811,N_15989,N_17797);
xnor U24812 (N_24812,N_17942,N_19903);
xor U24813 (N_24813,N_16566,N_15906);
or U24814 (N_24814,N_16560,N_18360);
xnor U24815 (N_24815,N_18113,N_17822);
nand U24816 (N_24816,N_18932,N_17698);
or U24817 (N_24817,N_18139,N_19042);
nand U24818 (N_24818,N_16640,N_17508);
xor U24819 (N_24819,N_17467,N_18172);
nand U24820 (N_24820,N_15696,N_17904);
and U24821 (N_24821,N_15675,N_15662);
and U24822 (N_24822,N_16401,N_15367);
or U24823 (N_24823,N_15392,N_18303);
nor U24824 (N_24824,N_15527,N_18148);
and U24825 (N_24825,N_18169,N_16330);
nor U24826 (N_24826,N_18146,N_19185);
nand U24827 (N_24827,N_15006,N_16266);
or U24828 (N_24828,N_18480,N_15946);
nand U24829 (N_24829,N_19241,N_17835);
and U24830 (N_24830,N_19336,N_16616);
nand U24831 (N_24831,N_15398,N_19340);
nor U24832 (N_24832,N_17685,N_18917);
or U24833 (N_24833,N_16656,N_16132);
xor U24834 (N_24834,N_17275,N_16333);
or U24835 (N_24835,N_16753,N_19114);
and U24836 (N_24836,N_18338,N_16366);
or U24837 (N_24837,N_17633,N_15410);
or U24838 (N_24838,N_16890,N_18472);
nand U24839 (N_24839,N_16920,N_16194);
and U24840 (N_24840,N_18597,N_19292);
or U24841 (N_24841,N_19777,N_17610);
nor U24842 (N_24842,N_17186,N_18001);
and U24843 (N_24843,N_19576,N_18279);
nor U24844 (N_24844,N_15246,N_17194);
nand U24845 (N_24845,N_17085,N_15289);
nor U24846 (N_24846,N_15967,N_15382);
nor U24847 (N_24847,N_18893,N_19900);
nor U24848 (N_24848,N_18748,N_16404);
nand U24849 (N_24849,N_19069,N_17144);
nor U24850 (N_24850,N_17821,N_18802);
nor U24851 (N_24851,N_16723,N_17888);
or U24852 (N_24852,N_15317,N_19512);
or U24853 (N_24853,N_19698,N_16772);
and U24854 (N_24854,N_15735,N_19468);
nor U24855 (N_24855,N_19229,N_15473);
or U24856 (N_24856,N_16503,N_16290);
and U24857 (N_24857,N_16778,N_18633);
or U24858 (N_24858,N_16954,N_15120);
nor U24859 (N_24859,N_15671,N_17065);
nor U24860 (N_24860,N_16648,N_15397);
and U24861 (N_24861,N_16812,N_18275);
xnor U24862 (N_24862,N_18057,N_18778);
xnor U24863 (N_24863,N_16991,N_16464);
and U24864 (N_24864,N_19512,N_17800);
and U24865 (N_24865,N_18449,N_17316);
or U24866 (N_24866,N_19065,N_19445);
and U24867 (N_24867,N_19219,N_15122);
or U24868 (N_24868,N_16321,N_18314);
nor U24869 (N_24869,N_17502,N_19882);
and U24870 (N_24870,N_18647,N_18193);
and U24871 (N_24871,N_19565,N_16171);
and U24872 (N_24872,N_16907,N_15737);
or U24873 (N_24873,N_15721,N_18929);
nor U24874 (N_24874,N_19390,N_16693);
nor U24875 (N_24875,N_17337,N_15041);
and U24876 (N_24876,N_15949,N_15027);
nand U24877 (N_24877,N_15121,N_18760);
and U24878 (N_24878,N_19396,N_18681);
or U24879 (N_24879,N_16056,N_16535);
and U24880 (N_24880,N_16119,N_17815);
nand U24881 (N_24881,N_18063,N_19594);
nand U24882 (N_24882,N_16882,N_17828);
and U24883 (N_24883,N_16989,N_18009);
nand U24884 (N_24884,N_15773,N_15743);
or U24885 (N_24885,N_17040,N_18807);
and U24886 (N_24886,N_16159,N_18666);
nor U24887 (N_24887,N_16117,N_17393);
and U24888 (N_24888,N_15488,N_19950);
nand U24889 (N_24889,N_15089,N_16904);
nand U24890 (N_24890,N_18968,N_16610);
nor U24891 (N_24891,N_16063,N_18634);
or U24892 (N_24892,N_15524,N_18856);
nand U24893 (N_24893,N_18924,N_17961);
nor U24894 (N_24894,N_15505,N_15418);
xor U24895 (N_24895,N_18367,N_17092);
nand U24896 (N_24896,N_16928,N_19387);
nand U24897 (N_24897,N_19082,N_16405);
or U24898 (N_24898,N_19120,N_19864);
xnor U24899 (N_24899,N_19795,N_18520);
or U24900 (N_24900,N_18237,N_16134);
and U24901 (N_24901,N_15052,N_17090);
nand U24902 (N_24902,N_16276,N_18321);
or U24903 (N_24903,N_15953,N_18061);
and U24904 (N_24904,N_18054,N_19727);
or U24905 (N_24905,N_18725,N_17390);
and U24906 (N_24906,N_16853,N_16798);
or U24907 (N_24907,N_17772,N_16264);
nor U24908 (N_24908,N_17681,N_15861);
nor U24909 (N_24909,N_16780,N_18821);
nor U24910 (N_24910,N_18531,N_17715);
nor U24911 (N_24911,N_18686,N_16541);
or U24912 (N_24912,N_19487,N_19402);
nand U24913 (N_24913,N_15111,N_18045);
nor U24914 (N_24914,N_15044,N_18668);
and U24915 (N_24915,N_19299,N_17075);
or U24916 (N_24916,N_19982,N_15891);
nand U24917 (N_24917,N_18602,N_15692);
or U24918 (N_24918,N_15498,N_19817);
xnor U24919 (N_24919,N_18286,N_17496);
or U24920 (N_24920,N_18752,N_16166);
nand U24921 (N_24921,N_15830,N_19653);
and U24922 (N_24922,N_19455,N_19609);
or U24923 (N_24923,N_19766,N_19916);
and U24924 (N_24924,N_19443,N_17329);
nor U24925 (N_24925,N_17412,N_15398);
nor U24926 (N_24926,N_15556,N_18409);
nand U24927 (N_24927,N_17340,N_18806);
nand U24928 (N_24928,N_18348,N_16553);
nand U24929 (N_24929,N_15945,N_16281);
nor U24930 (N_24930,N_19794,N_17953);
nand U24931 (N_24931,N_18797,N_16234);
or U24932 (N_24932,N_16035,N_16746);
or U24933 (N_24933,N_16322,N_15346);
or U24934 (N_24934,N_15617,N_18561);
and U24935 (N_24935,N_15911,N_19864);
nor U24936 (N_24936,N_19839,N_19220);
and U24937 (N_24937,N_18833,N_17671);
nor U24938 (N_24938,N_19763,N_15121);
or U24939 (N_24939,N_18670,N_17911);
nand U24940 (N_24940,N_19500,N_15417);
and U24941 (N_24941,N_19124,N_16050);
xnor U24942 (N_24942,N_18813,N_15307);
and U24943 (N_24943,N_17528,N_16501);
or U24944 (N_24944,N_18369,N_18866);
nand U24945 (N_24945,N_18518,N_15687);
nand U24946 (N_24946,N_16362,N_18147);
or U24947 (N_24947,N_16298,N_19058);
nor U24948 (N_24948,N_19278,N_16673);
or U24949 (N_24949,N_18805,N_16873);
or U24950 (N_24950,N_18950,N_19069);
and U24951 (N_24951,N_17053,N_17655);
and U24952 (N_24952,N_15398,N_19110);
nand U24953 (N_24953,N_15150,N_17105);
nand U24954 (N_24954,N_16773,N_17489);
nand U24955 (N_24955,N_19438,N_16857);
or U24956 (N_24956,N_17518,N_15568);
and U24957 (N_24957,N_15356,N_18360);
xor U24958 (N_24958,N_19140,N_19234);
nand U24959 (N_24959,N_18533,N_16231);
and U24960 (N_24960,N_15606,N_15491);
xor U24961 (N_24961,N_16250,N_18023);
or U24962 (N_24962,N_19996,N_15785);
nor U24963 (N_24963,N_17457,N_19924);
nor U24964 (N_24964,N_17197,N_17632);
nand U24965 (N_24965,N_18387,N_18393);
and U24966 (N_24966,N_18602,N_15645);
or U24967 (N_24967,N_15096,N_19186);
xor U24968 (N_24968,N_18154,N_15285);
or U24969 (N_24969,N_18718,N_16188);
xor U24970 (N_24970,N_17651,N_17364);
or U24971 (N_24971,N_15642,N_19265);
and U24972 (N_24972,N_18680,N_15052);
and U24973 (N_24973,N_16502,N_16504);
nand U24974 (N_24974,N_15127,N_15777);
nor U24975 (N_24975,N_19829,N_16855);
nand U24976 (N_24976,N_15292,N_18878);
or U24977 (N_24977,N_18134,N_16870);
nor U24978 (N_24978,N_18758,N_16570);
nand U24979 (N_24979,N_17066,N_17258);
and U24980 (N_24980,N_18146,N_17991);
nand U24981 (N_24981,N_19092,N_17337);
or U24982 (N_24982,N_17979,N_19940);
nand U24983 (N_24983,N_15620,N_18924);
and U24984 (N_24984,N_18608,N_15634);
nor U24985 (N_24985,N_18806,N_15244);
nand U24986 (N_24986,N_19520,N_17516);
or U24987 (N_24987,N_19130,N_19292);
nand U24988 (N_24988,N_19713,N_17930);
nand U24989 (N_24989,N_17247,N_19947);
or U24990 (N_24990,N_19839,N_18441);
or U24991 (N_24991,N_15978,N_17994);
xnor U24992 (N_24992,N_18059,N_15759);
nor U24993 (N_24993,N_15412,N_17217);
and U24994 (N_24994,N_17772,N_18350);
nor U24995 (N_24995,N_16052,N_19785);
xnor U24996 (N_24996,N_18384,N_17919);
nor U24997 (N_24997,N_17231,N_19983);
nor U24998 (N_24998,N_18436,N_17336);
or U24999 (N_24999,N_19570,N_15389);
xor U25000 (N_25000,N_23435,N_24234);
nand U25001 (N_25001,N_20970,N_20812);
xor U25002 (N_25002,N_24855,N_24504);
or U25003 (N_25003,N_24209,N_21546);
nor U25004 (N_25004,N_22835,N_23302);
nand U25005 (N_25005,N_22679,N_22307);
nor U25006 (N_25006,N_20412,N_22209);
and U25007 (N_25007,N_21870,N_20557);
nand U25008 (N_25008,N_24172,N_20836);
or U25009 (N_25009,N_24016,N_22255);
and U25010 (N_25010,N_21795,N_20338);
nor U25011 (N_25011,N_23393,N_21639);
nand U25012 (N_25012,N_21695,N_23361);
nand U25013 (N_25013,N_22365,N_21591);
or U25014 (N_25014,N_20990,N_22667);
and U25015 (N_25015,N_21682,N_20509);
nand U25016 (N_25016,N_24212,N_23181);
and U25017 (N_25017,N_22511,N_21997);
and U25018 (N_25018,N_24254,N_24207);
xnor U25019 (N_25019,N_20712,N_22238);
and U25020 (N_25020,N_20986,N_22986);
nand U25021 (N_25021,N_20906,N_23833);
nor U25022 (N_25022,N_24849,N_21509);
nor U25023 (N_25023,N_24693,N_20435);
nor U25024 (N_25024,N_24577,N_23224);
nand U25025 (N_25025,N_23561,N_22089);
and U25026 (N_25026,N_24665,N_23053);
or U25027 (N_25027,N_22176,N_22792);
nand U25028 (N_25028,N_22999,N_22827);
nand U25029 (N_25029,N_20735,N_20516);
and U25030 (N_25030,N_24673,N_21621);
or U25031 (N_25031,N_22322,N_21897);
nor U25032 (N_25032,N_21864,N_20955);
nor U25033 (N_25033,N_22861,N_21961);
or U25034 (N_25034,N_22126,N_22149);
and U25035 (N_25035,N_21972,N_22570);
or U25036 (N_25036,N_22973,N_22968);
and U25037 (N_25037,N_22914,N_21475);
xor U25038 (N_25038,N_21121,N_20785);
and U25039 (N_25039,N_20388,N_24318);
or U25040 (N_25040,N_20695,N_21882);
or U25041 (N_25041,N_24407,N_22682);
and U25042 (N_25042,N_24628,N_21089);
or U25043 (N_25043,N_20567,N_24345);
nor U25044 (N_25044,N_23108,N_20157);
or U25045 (N_25045,N_22744,N_22996);
nor U25046 (N_25046,N_21743,N_21545);
or U25047 (N_25047,N_22035,N_21287);
nor U25048 (N_25048,N_24513,N_20947);
and U25049 (N_25049,N_24439,N_22358);
nand U25050 (N_25050,N_24330,N_21854);
nand U25051 (N_25051,N_23754,N_22109);
and U25052 (N_25052,N_23848,N_21815);
xor U25053 (N_25053,N_23348,N_24590);
nor U25054 (N_25054,N_20225,N_22512);
or U25055 (N_25055,N_21304,N_21818);
or U25056 (N_25056,N_23425,N_24866);
nor U25057 (N_25057,N_20723,N_24206);
nand U25058 (N_25058,N_23459,N_21525);
nand U25059 (N_25059,N_21608,N_20458);
nand U25060 (N_25060,N_20896,N_24013);
nand U25061 (N_25061,N_22295,N_20886);
or U25062 (N_25062,N_24214,N_22446);
or U25063 (N_25063,N_22435,N_24377);
nand U25064 (N_25064,N_22854,N_24908);
xnor U25065 (N_25065,N_24552,N_24089);
nor U25066 (N_25066,N_20775,N_23633);
xnor U25067 (N_25067,N_22502,N_22677);
nand U25068 (N_25068,N_23956,N_20211);
or U25069 (N_25069,N_23385,N_23607);
nand U25070 (N_25070,N_21480,N_21582);
or U25071 (N_25071,N_23723,N_23146);
xnor U25072 (N_25072,N_22706,N_21804);
or U25073 (N_25073,N_23000,N_20314);
nor U25074 (N_25074,N_22586,N_21796);
nor U25075 (N_25075,N_23946,N_23211);
and U25076 (N_25076,N_23855,N_22545);
nand U25077 (N_25077,N_20964,N_21022);
or U25078 (N_25078,N_20422,N_21188);
nor U25079 (N_25079,N_22998,N_20400);
nor U25080 (N_25080,N_24793,N_22098);
nand U25081 (N_25081,N_24178,N_21152);
xor U25082 (N_25082,N_23358,N_20615);
or U25083 (N_25083,N_21573,N_23470);
and U25084 (N_25084,N_22666,N_22179);
or U25085 (N_25085,N_21189,N_20767);
nor U25086 (N_25086,N_20256,N_22641);
or U25087 (N_25087,N_23781,N_22216);
nand U25088 (N_25088,N_23680,N_23977);
or U25089 (N_25089,N_20020,N_23274);
nand U25090 (N_25090,N_22001,N_20163);
or U25091 (N_25091,N_23487,N_20654);
or U25092 (N_25092,N_21960,N_21452);
nand U25093 (N_25093,N_20015,N_23481);
and U25094 (N_25094,N_21229,N_23111);
and U25095 (N_25095,N_21737,N_21209);
or U25096 (N_25096,N_20579,N_24134);
or U25097 (N_25097,N_22463,N_20880);
or U25098 (N_25098,N_20559,N_24687);
nor U25099 (N_25099,N_21176,N_23960);
nand U25100 (N_25100,N_24691,N_24306);
and U25101 (N_25101,N_24356,N_21421);
and U25102 (N_25102,N_22655,N_22548);
nand U25103 (N_25103,N_21555,N_20278);
and U25104 (N_25104,N_21801,N_23290);
nand U25105 (N_25105,N_23472,N_23475);
nand U25106 (N_25106,N_23340,N_23789);
nor U25107 (N_25107,N_23372,N_20003);
or U25108 (N_25108,N_23457,N_21060);
and U25109 (N_25109,N_24718,N_21858);
nand U25110 (N_25110,N_23350,N_23996);
and U25111 (N_25111,N_22724,N_21023);
nand U25112 (N_25112,N_24763,N_22060);
xnor U25113 (N_25113,N_24004,N_23471);
nand U25114 (N_25114,N_20308,N_20645);
nor U25115 (N_25115,N_21810,N_23642);
nand U25116 (N_25116,N_20073,N_24889);
nand U25117 (N_25117,N_22870,N_22290);
and U25118 (N_25118,N_23606,N_20231);
and U25119 (N_25119,N_21698,N_23896);
and U25120 (N_25120,N_21167,N_21297);
or U25121 (N_25121,N_20737,N_20530);
xor U25122 (N_25122,N_21148,N_21539);
nand U25123 (N_25123,N_20887,N_22627);
nor U25124 (N_25124,N_23987,N_24405);
nor U25125 (N_25125,N_24309,N_22492);
or U25126 (N_25126,N_23814,N_23344);
nor U25127 (N_25127,N_21093,N_24143);
xnor U25128 (N_25128,N_22116,N_23582);
or U25129 (N_25129,N_23605,N_23635);
or U25130 (N_25130,N_23081,N_23534);
nand U25131 (N_25131,N_23811,N_21277);
and U25132 (N_25132,N_22993,N_24477);
xor U25133 (N_25133,N_22913,N_22066);
nand U25134 (N_25134,N_23812,N_21044);
nor U25135 (N_25135,N_23375,N_22036);
nor U25136 (N_25136,N_24743,N_20273);
xor U25137 (N_25137,N_21399,N_22782);
nand U25138 (N_25138,N_24991,N_22232);
xnor U25139 (N_25139,N_23755,N_23866);
nand U25140 (N_25140,N_24805,N_22153);
nand U25141 (N_25141,N_22762,N_20480);
nand U25142 (N_25142,N_20022,N_20001);
and U25143 (N_25143,N_20716,N_20543);
or U25144 (N_25144,N_20550,N_24277);
nor U25145 (N_25145,N_23636,N_20856);
or U25146 (N_25146,N_20203,N_20726);
or U25147 (N_25147,N_23863,N_20113);
xnor U25148 (N_25148,N_20407,N_24390);
nor U25149 (N_25149,N_22202,N_22242);
nand U25150 (N_25150,N_22620,N_24150);
or U25151 (N_25151,N_20552,N_23469);
or U25152 (N_25152,N_20968,N_21441);
and U25153 (N_25153,N_22268,N_23734);
and U25154 (N_25154,N_21569,N_21881);
xor U25155 (N_25155,N_24807,N_24457);
nand U25156 (N_25156,N_20434,N_20583);
nand U25157 (N_25157,N_22263,N_20133);
or U25158 (N_25158,N_22793,N_20883);
nand U25159 (N_25159,N_23911,N_24817);
nand U25160 (N_25160,N_24905,N_21606);
nor U25161 (N_25161,N_20063,N_22270);
nand U25162 (N_25162,N_21785,N_21657);
nor U25163 (N_25163,N_22194,N_23955);
or U25164 (N_25164,N_21109,N_24963);
and U25165 (N_25165,N_22693,N_23617);
nor U25166 (N_25166,N_23984,N_23058);
nand U25167 (N_25167,N_23632,N_24620);
and U25168 (N_25168,N_23659,N_21885);
and U25169 (N_25169,N_23029,N_24989);
and U25170 (N_25170,N_21631,N_21351);
or U25171 (N_25171,N_24595,N_22305);
nand U25172 (N_25172,N_20507,N_24675);
nor U25173 (N_25173,N_22475,N_21294);
xnor U25174 (N_25174,N_20491,N_23940);
nor U25175 (N_25175,N_23428,N_21928);
nand U25176 (N_25176,N_23882,N_23041);
or U25177 (N_25177,N_22201,N_21625);
and U25178 (N_25178,N_21068,N_22625);
nand U25179 (N_25179,N_23669,N_21630);
or U25180 (N_25180,N_20622,N_24154);
nor U25181 (N_25181,N_20111,N_20833);
nand U25182 (N_25182,N_20123,N_24401);
xor U25183 (N_25183,N_20217,N_21074);
or U25184 (N_25184,N_22525,N_22286);
or U25185 (N_25185,N_23787,N_22980);
xnor U25186 (N_25186,N_21713,N_22729);
or U25187 (N_25187,N_20710,N_24317);
nor U25188 (N_25188,N_23722,N_21381);
and U25189 (N_25189,N_23953,N_23176);
nand U25190 (N_25190,N_24796,N_22046);
and U25191 (N_25191,N_20998,N_21720);
and U25192 (N_25192,N_20066,N_20206);
or U25193 (N_25193,N_21149,N_21243);
and U25194 (N_25194,N_23159,N_21083);
and U25195 (N_25195,N_24970,N_20824);
or U25196 (N_25196,N_24662,N_23704);
and U25197 (N_25197,N_24219,N_21146);
and U25198 (N_25198,N_24153,N_20598);
nor U25199 (N_25199,N_20146,N_23851);
xnor U25200 (N_25200,N_24075,N_23979);
and U25201 (N_25201,N_23551,N_20055);
nand U25202 (N_25202,N_20379,N_23141);
xor U25203 (N_25203,N_20465,N_22317);
and U25204 (N_25204,N_23918,N_20238);
or U25205 (N_25205,N_22595,N_21444);
and U25206 (N_25206,N_20593,N_22758);
or U25207 (N_25207,N_22722,N_23758);
and U25208 (N_25208,N_24259,N_24081);
or U25209 (N_25209,N_20832,N_24860);
or U25210 (N_25210,N_21353,N_23529);
and U25211 (N_25211,N_23584,N_20074);
and U25212 (N_25212,N_24922,N_23210);
nor U25213 (N_25213,N_20352,N_24140);
or U25214 (N_25214,N_23281,N_21218);
nor U25215 (N_25215,N_23881,N_22629);
and U25216 (N_25216,N_23062,N_20941);
xnor U25217 (N_25217,N_22946,N_22774);
xnor U25218 (N_25218,N_22079,N_21678);
nand U25219 (N_25219,N_22369,N_20870);
nor U25220 (N_25220,N_22389,N_22632);
and U25221 (N_25221,N_21021,N_23388);
nand U25222 (N_25222,N_23868,N_23877);
nor U25223 (N_25223,N_23152,N_23986);
and U25224 (N_25224,N_23075,N_23328);
xnor U25225 (N_25225,N_21194,N_24139);
or U25226 (N_25226,N_20177,N_24814);
and U25227 (N_25227,N_23906,N_23491);
nand U25228 (N_25228,N_21503,N_22166);
nand U25229 (N_25229,N_23500,N_22649);
nand U25230 (N_25230,N_23107,N_23154);
nor U25231 (N_25231,N_24525,N_22838);
xor U25232 (N_25232,N_22982,N_24488);
and U25233 (N_25233,N_21724,N_22842);
nor U25234 (N_25234,N_21833,N_24830);
and U25235 (N_25235,N_23850,N_22325);
xor U25236 (N_25236,N_23715,N_21413);
xnor U25237 (N_25237,N_21586,N_21157);
and U25238 (N_25238,N_23043,N_20834);
nand U25239 (N_25239,N_23175,N_21267);
or U25240 (N_25240,N_23024,N_24419);
nor U25241 (N_25241,N_24574,N_24692);
or U25242 (N_25242,N_22534,N_23552);
nor U25243 (N_25243,N_23068,N_24142);
nor U25244 (N_25244,N_23884,N_21099);
nor U25245 (N_25245,N_23038,N_20302);
xor U25246 (N_25246,N_24274,N_23801);
nand U25247 (N_25247,N_21255,N_20118);
nand U25248 (N_25248,N_23228,N_24184);
and U25249 (N_25249,N_23046,N_21211);
and U25250 (N_25250,N_24618,N_22908);
nand U25251 (N_25251,N_20331,N_20991);
nor U25252 (N_25252,N_22233,N_20221);
and U25253 (N_25253,N_22972,N_23123);
and U25254 (N_25254,N_20769,N_22125);
nor U25255 (N_25255,N_22464,N_23902);
xor U25256 (N_25256,N_21493,N_23624);
nand U25257 (N_25257,N_20818,N_20130);
or U25258 (N_25258,N_24031,N_21759);
or U25259 (N_25259,N_23718,N_24449);
xor U25260 (N_25260,N_24284,N_23645);
nor U25261 (N_25261,N_23702,N_20104);
nand U25262 (N_25262,N_24302,N_24825);
nand U25263 (N_25263,N_24508,N_23941);
nand U25264 (N_25264,N_24812,N_22636);
and U25265 (N_25265,N_20428,N_21105);
nand U25266 (N_25266,N_20080,N_22364);
nor U25267 (N_25267,N_21504,N_20497);
and U25268 (N_25268,N_24934,N_22957);
xnor U25269 (N_25269,N_22752,N_21220);
nand U25270 (N_25270,N_23729,N_21607);
and U25271 (N_25271,N_24430,N_23920);
nor U25272 (N_25272,N_23962,N_20081);
and U25273 (N_25273,N_21755,N_21921);
nand U25274 (N_25274,N_24049,N_22420);
xnor U25275 (N_25275,N_24785,N_22207);
or U25276 (N_25276,N_21394,N_22720);
or U25277 (N_25277,N_23686,N_20738);
or U25278 (N_25278,N_20058,N_21617);
nand U25279 (N_25279,N_24223,N_22193);
nand U25280 (N_25280,N_23069,N_24775);
nand U25281 (N_25281,N_22716,N_24250);
nand U25282 (N_25282,N_22123,N_22877);
nor U25283 (N_25283,N_21174,N_21315);
nand U25284 (N_25284,N_22097,N_24500);
nand U25285 (N_25285,N_20444,N_24882);
and U25286 (N_25286,N_22719,N_20373);
or U25287 (N_25287,N_21623,N_24593);
and U25288 (N_25288,N_23478,N_24028);
or U25289 (N_25289,N_22203,N_20069);
nor U25290 (N_25290,N_20090,N_22592);
nor U25291 (N_25291,N_23001,N_23852);
or U25292 (N_25292,N_22298,N_23883);
xnor U25293 (N_25293,N_20072,N_21723);
or U25294 (N_25294,N_21239,N_20354);
nand U25295 (N_25295,N_23816,N_21027);
xnor U25296 (N_25296,N_21227,N_21846);
nand U25297 (N_25297,N_22612,N_21199);
nand U25298 (N_25298,N_24005,N_22817);
and U25299 (N_25299,N_23629,N_24845);
or U25300 (N_25300,N_21793,N_22165);
or U25301 (N_25301,N_23720,N_21827);
or U25302 (N_25302,N_23429,N_21797);
or U25303 (N_25303,N_21474,N_24398);
or U25304 (N_25304,N_22495,N_21551);
and U25305 (N_25305,N_23291,N_23278);
nor U25306 (N_25306,N_20031,N_24017);
xor U25307 (N_25307,N_24000,N_24964);
nand U25308 (N_25308,N_23072,N_24490);
nor U25309 (N_25309,N_23751,N_20250);
and U25310 (N_25310,N_23978,N_20089);
xnor U25311 (N_25311,N_24828,N_23761);
and U25312 (N_25312,N_22223,N_23580);
and U25313 (N_25313,N_22014,N_23540);
nor U25314 (N_25314,N_24364,N_21590);
nand U25315 (N_25315,N_24097,N_20076);
or U25316 (N_25316,N_22024,N_21633);
nand U25317 (N_25317,N_20156,N_20105);
xnor U25318 (N_25318,N_24975,N_23620);
or U25319 (N_25319,N_23737,N_22418);
or U25320 (N_25320,N_21522,N_24363);
nor U25321 (N_25321,N_21802,N_23351);
nand U25322 (N_25322,N_24819,N_23296);
or U25323 (N_25323,N_23499,N_20169);
nor U25324 (N_25324,N_21982,N_23251);
xor U25325 (N_25325,N_24900,N_22254);
nor U25326 (N_25326,N_20647,N_20688);
nor U25327 (N_25327,N_24119,N_22910);
or U25328 (N_25328,N_23837,N_21041);
nand U25329 (N_25329,N_24400,N_23065);
nor U25330 (N_25330,N_22481,N_23673);
or U25331 (N_25331,N_23386,N_20555);
nand U25332 (N_25332,N_20402,N_21537);
and U25333 (N_25333,N_23783,N_20666);
and U25334 (N_25334,N_24899,N_20188);
nor U25335 (N_25335,N_24251,N_21873);
and U25336 (N_25336,N_23546,N_22346);
nand U25337 (N_25337,N_20770,N_22170);
or U25338 (N_25338,N_24783,N_22673);
nor U25339 (N_25339,N_24193,N_20734);
nor U25340 (N_25340,N_24984,N_21547);
nand U25341 (N_25341,N_22276,N_21417);
nor U25342 (N_25342,N_23307,N_22830);
or U25343 (N_25343,N_22520,N_24327);
nand U25344 (N_25344,N_21282,N_21122);
nor U25345 (N_25345,N_22734,N_21283);
or U25346 (N_25346,N_22936,N_22969);
nand U25347 (N_25347,N_21223,N_24231);
nand U25348 (N_25348,N_21448,N_22763);
or U25349 (N_25349,N_21519,N_20096);
or U25350 (N_25350,N_22139,N_24024);
nor U25351 (N_25351,N_22015,N_22575);
nand U25352 (N_25352,N_21426,N_22384);
or U25353 (N_25353,N_22228,N_22181);
or U25354 (N_25354,N_21050,N_24926);
nand U25355 (N_25355,N_24957,N_22903);
nor U25356 (N_25356,N_20449,N_23971);
and U25357 (N_25357,N_23148,N_23219);
nand U25358 (N_25358,N_21242,N_24703);
nand U25359 (N_25359,N_21420,N_23262);
nand U25360 (N_25360,N_24344,N_23473);
xnor U25361 (N_25361,N_21436,N_22362);
or U25362 (N_25362,N_24579,N_20167);
or U25363 (N_25363,N_22219,N_24465);
nand U25364 (N_25364,N_24086,N_22497);
or U25365 (N_25365,N_24598,N_23409);
xor U25366 (N_25366,N_21530,N_20115);
nand U25367 (N_25367,N_24745,N_22319);
nand U25368 (N_25368,N_21548,N_21677);
nand U25369 (N_25369,N_23791,N_20235);
or U25370 (N_25370,N_20023,N_22544);
or U25371 (N_25371,N_22940,N_22010);
or U25372 (N_25372,N_21322,N_24832);
nand U25373 (N_25373,N_24539,N_24227);
nor U25374 (N_25374,N_23447,N_22188);
xor U25375 (N_25375,N_21645,N_22563);
or U25376 (N_25376,N_24535,N_23229);
or U25377 (N_25377,N_20823,N_21541);
xnor U25378 (N_25378,N_21675,N_24612);
nor U25379 (N_25379,N_23594,N_21328);
nor U25380 (N_25380,N_20774,N_21574);
nor U25381 (N_25381,N_23912,N_20587);
nor U25382 (N_25382,N_23450,N_20576);
nand U25383 (N_25383,N_24560,N_24591);
or U25384 (N_25384,N_23690,N_24945);
or U25385 (N_25385,N_23028,N_21129);
or U25386 (N_25386,N_24600,N_22656);
xnor U25387 (N_25387,N_21952,N_23609);
xnor U25388 (N_25388,N_21138,N_22312);
nor U25389 (N_25389,N_22959,N_21392);
or U25390 (N_25390,N_21604,N_22327);
and U25391 (N_25391,N_23039,N_21779);
and U25392 (N_25392,N_20474,N_20100);
nor U25393 (N_25393,N_20733,N_20298);
nor U25394 (N_25394,N_22761,N_24441);
nor U25395 (N_25395,N_20699,N_23543);
nor U25396 (N_25396,N_20320,N_20008);
xnor U25397 (N_25397,N_22448,N_20742);
nor U25398 (N_25398,N_21663,N_24810);
nand U25399 (N_25399,N_22076,N_21418);
or U25400 (N_25400,N_22439,N_20925);
xnor U25401 (N_25401,N_22155,N_24505);
nand U25402 (N_25402,N_24782,N_24839);
nand U25403 (N_25403,N_22626,N_21140);
nand U25404 (N_25404,N_24268,N_22743);
and U25405 (N_25405,N_20838,N_21279);
or U25406 (N_25406,N_23698,N_21831);
xnor U25407 (N_25407,N_21671,N_23799);
or U25408 (N_25408,N_22415,N_21688);
nand U25409 (N_25409,N_22905,N_20045);
nor U25410 (N_25410,N_21020,N_20237);
or U25411 (N_25411,N_22971,N_23179);
or U25412 (N_25412,N_24396,N_22469);
or U25413 (N_25413,N_22549,N_20881);
xor U25414 (N_25414,N_23516,N_20650);
nor U25415 (N_25415,N_23929,N_23989);
or U25416 (N_25416,N_23027,N_23272);
xor U25417 (N_25417,N_24052,N_24104);
nor U25418 (N_25418,N_22985,N_24655);
or U25419 (N_25419,N_21440,N_20591);
or U25420 (N_25420,N_20884,N_20164);
and U25421 (N_25421,N_23293,N_22360);
nand U25422 (N_25422,N_20663,N_22902);
nand U25423 (N_25423,N_22361,N_20272);
nor U25424 (N_25424,N_21934,N_23144);
nand U25425 (N_25425,N_24019,N_23103);
nand U25426 (N_25426,N_24597,N_23910);
and U25427 (N_25427,N_24079,N_21403);
and U25428 (N_25428,N_21108,N_22546);
and U25429 (N_25429,N_21288,N_21757);
nor U25430 (N_25430,N_24395,N_24462);
or U25431 (N_25431,N_22794,N_20929);
nand U25432 (N_25432,N_24823,N_22450);
nand U25433 (N_25433,N_22933,N_23846);
xnor U25434 (N_25434,N_24348,N_21124);
nor U25435 (N_25435,N_23903,N_24025);
xnor U25436 (N_25436,N_20623,N_24165);
nor U25437 (N_25437,N_24246,N_22206);
and U25438 (N_25438,N_20585,N_20805);
or U25439 (N_25439,N_23049,N_20995);
and U25440 (N_25440,N_20420,N_24599);
nor U25441 (N_25441,N_22948,N_21907);
nor U25442 (N_25442,N_23449,N_24791);
nand U25443 (N_25443,N_23364,N_24766);
xnor U25444 (N_25444,N_22859,N_23926);
nor U25445 (N_25445,N_24290,N_23667);
or U25446 (N_25446,N_24857,N_22218);
or U25447 (N_25447,N_22990,N_24841);
nor U25448 (N_25448,N_22726,N_23333);
nand U25449 (N_25449,N_20365,N_21372);
or U25450 (N_25450,N_24282,N_21766);
and U25451 (N_25451,N_20496,N_20141);
and U25452 (N_25452,N_21339,N_21332);
nor U25453 (N_25453,N_22490,N_20972);
nor U25454 (N_25454,N_21857,N_22302);
or U25455 (N_25455,N_23188,N_20924);
nand U25456 (N_25456,N_21772,N_23894);
or U25457 (N_25457,N_24846,N_21821);
and U25458 (N_25458,N_21366,N_24243);
nor U25459 (N_25459,N_21003,N_22467);
or U25460 (N_25460,N_24478,N_20762);
or U25461 (N_25461,N_20077,N_24608);
or U25462 (N_25462,N_21753,N_20321);
or U25463 (N_25463,N_23446,N_22260);
or U25464 (N_25464,N_21196,N_23611);
and U25465 (N_25465,N_20265,N_22006);
or U25466 (N_25466,N_23055,N_24994);
xnor U25467 (N_25467,N_20129,N_20503);
or U25468 (N_25468,N_22237,N_22961);
or U25469 (N_25469,N_22065,N_21517);
and U25470 (N_25470,N_21906,N_23453);
and U25471 (N_25471,N_24808,N_22550);
or U25472 (N_25472,N_24879,N_21313);
and U25473 (N_25473,N_20335,N_23138);
nor U25474 (N_25474,N_24448,N_21234);
xor U25475 (N_25475,N_23007,N_23724);
or U25476 (N_25476,N_20050,N_22584);
nand U25477 (N_25477,N_21959,N_20943);
or U25478 (N_25478,N_22494,N_20124);
and U25479 (N_25479,N_21690,N_21042);
nand U25480 (N_25480,N_22642,N_20212);
or U25481 (N_25481,N_20686,N_24602);
or U25482 (N_25482,N_20529,N_20556);
and U25483 (N_25483,N_21251,N_22825);
nor U25484 (N_25484,N_20918,N_21847);
nor U25485 (N_25485,N_21526,N_24541);
and U25486 (N_25486,N_22934,N_23283);
or U25487 (N_25487,N_23448,N_20535);
nand U25488 (N_25488,N_24756,N_20617);
and U25489 (N_25489,N_24792,N_23662);
xnor U25490 (N_25490,N_21762,N_24469);
or U25491 (N_25491,N_20161,N_24651);
nand U25492 (N_25492,N_24393,N_21273);
and U25493 (N_25493,N_21280,N_22354);
nand U25494 (N_25494,N_20382,N_21927);
nand U25495 (N_25495,N_23511,N_23285);
or U25496 (N_25496,N_23652,N_20706);
nand U25497 (N_25497,N_22199,N_24114);
nor U25498 (N_25498,N_20461,N_21727);
nor U25499 (N_25499,N_24068,N_22564);
nor U25500 (N_25500,N_21516,N_24434);
and U25501 (N_25501,N_23312,N_20674);
or U25502 (N_25502,N_20814,N_21697);
and U25503 (N_25503,N_24511,N_21076);
nor U25504 (N_25504,N_21655,N_22653);
or U25505 (N_25505,N_22652,N_20872);
nand U25506 (N_25506,N_24631,N_24789);
nor U25507 (N_25507,N_20983,N_23542);
or U25508 (N_25508,N_24901,N_21320);
or U25509 (N_25509,N_24360,N_22185);
nor U25510 (N_25510,N_22618,N_21518);
or U25511 (N_25511,N_23600,N_24942);
xnor U25512 (N_25512,N_22912,N_22177);
and U25513 (N_25513,N_21528,N_23074);
or U25514 (N_25514,N_22528,N_24906);
or U25515 (N_25515,N_23016,N_23433);
and U25516 (N_25516,N_22950,N_24834);
or U25517 (N_25517,N_21704,N_20323);
nor U25518 (N_25518,N_24294,N_24515);
nand U25519 (N_25519,N_21616,N_23401);
nor U25520 (N_25520,N_21919,N_22853);
or U25521 (N_25521,N_24533,N_24506);
nor U25522 (N_25522,N_22489,N_21396);
nand U25523 (N_25523,N_21808,N_20804);
or U25524 (N_25524,N_20675,N_20239);
or U25525 (N_25525,N_20334,N_24313);
nor U25526 (N_25526,N_24871,N_22243);
nor U25527 (N_25527,N_24528,N_23689);
and U25528 (N_25528,N_24741,N_22157);
xor U25529 (N_25529,N_23992,N_20811);
and U25530 (N_25530,N_23379,N_23657);
or U25531 (N_25531,N_21389,N_20882);
nand U25532 (N_25532,N_21184,N_21600);
and U25533 (N_25533,N_23128,N_20751);
xor U25534 (N_25534,N_20916,N_20952);
and U25535 (N_25535,N_23872,N_23663);
or U25536 (N_25536,N_22474,N_22868);
or U25537 (N_25537,N_22355,N_22906);
xnor U25538 (N_25538,N_20160,N_22701);
xor U25539 (N_25539,N_22651,N_22247);
nor U25540 (N_25540,N_24365,N_20378);
or U25541 (N_25541,N_22480,N_22577);
and U25542 (N_25542,N_21387,N_24040);
or U25543 (N_25543,N_23891,N_23384);
xor U25544 (N_25544,N_24605,N_21082);
and U25545 (N_25545,N_23909,N_24359);
nor U25546 (N_25546,N_22404,N_24753);
xor U25547 (N_25547,N_21741,N_24397);
nor U25548 (N_25548,N_21913,N_22379);
nand U25549 (N_25549,N_22120,N_24615);
xnor U25550 (N_25550,N_20739,N_23426);
xor U25551 (N_25551,N_23867,N_24180);
or U25552 (N_25552,N_23368,N_24854);
nand U25553 (N_25553,N_20510,N_23047);
and U25554 (N_25554,N_24437,N_21637);
or U25555 (N_25555,N_20898,N_20019);
or U25556 (N_25556,N_20387,N_24135);
or U25557 (N_25557,N_20180,N_21686);
xor U25558 (N_25558,N_23951,N_23820);
nand U25559 (N_25559,N_21114,N_24204);
nor U25560 (N_25560,N_24787,N_24670);
or U25561 (N_25561,N_20065,N_23392);
nand U25562 (N_25562,N_24194,N_20633);
or U25563 (N_25563,N_22039,N_24242);
nand U25564 (N_25564,N_24532,N_24873);
nand U25565 (N_25565,N_22433,N_23042);
or U25566 (N_25566,N_24530,N_22991);
or U25567 (N_25567,N_23022,N_23120);
and U25568 (N_25568,N_22624,N_22602);
xor U25569 (N_25569,N_20079,N_24717);
and U25570 (N_25570,N_24494,N_22566);
nand U25571 (N_25571,N_23494,N_20581);
nor U25572 (N_25572,N_22703,N_23949);
or U25573 (N_25573,N_21627,N_24995);
and U25574 (N_25574,N_20506,N_21559);
or U25575 (N_25575,N_20519,N_21987);
nor U25576 (N_25576,N_22321,N_24780);
and U25577 (N_25577,N_21107,N_23760);
xor U25578 (N_25578,N_23060,N_21078);
and U25579 (N_25579,N_24296,N_20042);
and U25580 (N_25580,N_22493,N_24529);
nand U25581 (N_25581,N_23225,N_22663);
nor U25582 (N_25582,N_22925,N_23936);
nor U25583 (N_25583,N_22114,N_21871);
nor U25584 (N_25584,N_22009,N_23098);
and U25585 (N_25585,N_23099,N_24071);
nand U25586 (N_25586,N_23279,N_21567);
or U25587 (N_25587,N_23236,N_20218);
nand U25588 (N_25588,N_23404,N_23961);
nor U25589 (N_25589,N_21067,N_21489);
nand U25590 (N_25590,N_23231,N_20722);
nor U25591 (N_25591,N_23017,N_21700);
nor U25592 (N_25592,N_21711,N_21164);
and U25593 (N_25593,N_22088,N_21859);
and U25594 (N_25594,N_22129,N_22809);
xnor U25595 (N_25595,N_22888,N_23116);
xnor U25596 (N_25596,N_21894,N_20960);
nand U25597 (N_25597,N_22606,N_20743);
or U25598 (N_25598,N_23521,N_23654);
nor U25599 (N_25599,N_20607,N_23467);
xnor U25600 (N_25600,N_23419,N_20415);
nand U25601 (N_25601,N_22110,N_24794);
and U25602 (N_25602,N_22727,N_20869);
and U25603 (N_25603,N_22274,N_23003);
or U25604 (N_25604,N_22572,N_21973);
or U25605 (N_25605,N_20974,N_21009);
and U25606 (N_25606,N_22824,N_23567);
xor U25607 (N_25607,N_20099,N_22638);
nor U25608 (N_25608,N_22881,N_20935);
nand U25609 (N_25609,N_20830,N_21974);
xor U25610 (N_25610,N_24411,N_22997);
nand U25611 (N_25611,N_24236,N_23145);
or U25612 (N_25612,N_21529,N_20172);
nor U25613 (N_25613,N_24305,N_20857);
nor U25614 (N_25614,N_21661,N_22135);
nand U25615 (N_25615,N_20083,N_23477);
or U25616 (N_25616,N_22623,N_24026);
nor U25617 (N_25617,N_24270,N_20197);
nor U25618 (N_25618,N_22140,N_20705);
nand U25619 (N_25619,N_20729,N_21842);
and U25620 (N_25620,N_23343,N_21935);
nand U25621 (N_25621,N_21984,N_24913);
nand U25622 (N_25622,N_24295,N_21648);
nor U25623 (N_25623,N_20915,N_22732);
nand U25624 (N_25624,N_22173,N_21342);
nand U25625 (N_25625,N_21014,N_23779);
or U25626 (N_25626,N_23463,N_20253);
xnor U25627 (N_25627,N_24454,N_21767);
nand U25628 (N_25628,N_23217,N_24788);
nor U25629 (N_25629,N_22004,N_24838);
or U25630 (N_25630,N_20657,N_23458);
and U25631 (N_25631,N_23907,N_23610);
nor U25632 (N_25632,N_22900,N_24376);
nor U25633 (N_25633,N_20441,N_21470);
or U25634 (N_25634,N_24724,N_24299);
nand U25635 (N_25635,N_23876,N_24580);
or U25636 (N_25636,N_22044,N_23443);
or U25637 (N_25637,N_20874,N_23164);
xnor U25638 (N_25638,N_22523,N_20759);
or U25639 (N_25639,N_20690,N_23432);
and U25640 (N_25640,N_20088,N_23740);
nand U25641 (N_25641,N_20993,N_24925);
nand U25642 (N_25642,N_20483,N_20311);
nor U25643 (N_25643,N_21253,N_21683);
nand U25644 (N_25644,N_21428,N_24217);
xnor U25645 (N_25645,N_21760,N_24061);
nand U25646 (N_25646,N_24550,N_22956);
and U25647 (N_25647,N_22021,N_21407);
nor U25648 (N_25648,N_20837,N_20578);
and U25649 (N_25649,N_21742,N_21340);
nand U25650 (N_25650,N_23900,N_24021);
nand U25651 (N_25651,N_21127,N_20229);
nor U25652 (N_25652,N_20185,N_22210);
and U25653 (N_25653,N_20835,N_23819);
or U25654 (N_25654,N_21162,N_22396);
nor U25655 (N_25655,N_22963,N_20424);
and U25656 (N_25656,N_21676,N_24537);
nand U25657 (N_25657,N_24661,N_22611);
nor U25658 (N_25658,N_21434,N_23454);
nand U25659 (N_25659,N_21781,N_20827);
nor U25660 (N_25660,N_23577,N_20264);
and U25661 (N_25661,N_22334,N_20630);
and U25662 (N_25662,N_21497,N_22685);
and U25663 (N_25663,N_23444,N_21261);
or U25664 (N_25664,N_22037,N_21788);
and U25665 (N_25665,N_20667,N_24341);
and U25666 (N_25666,N_23665,N_22952);
or U25667 (N_25667,N_21026,N_24795);
nand U25668 (N_25668,N_20306,N_20512);
or U25669 (N_25669,N_20809,N_20829);
or U25670 (N_25670,N_22645,N_24131);
and U25671 (N_25671,N_24240,N_21705);
nand U25672 (N_25672,N_22454,N_20110);
nor U25673 (N_25673,N_22075,N_24969);
and U25674 (N_25674,N_20603,N_22073);
and U25675 (N_25675,N_22514,N_21778);
nand U25676 (N_25676,N_21749,N_22485);
or U25677 (N_25677,N_20171,N_21286);
and U25678 (N_25678,N_20490,N_22191);
or U25679 (N_25679,N_20243,N_22231);
nand U25680 (N_25680,N_21929,N_23277);
nor U25681 (N_25681,N_20282,N_22215);
or U25682 (N_25682,N_20563,N_21837);
and U25683 (N_25683,N_23070,N_21197);
and U25684 (N_25684,N_23982,N_21568);
and U25685 (N_25685,N_22955,N_22146);
or U25686 (N_25686,N_23040,N_21807);
nand U25687 (N_25687,N_21978,N_24516);
nand U25688 (N_25688,N_20370,N_24898);
xnor U25689 (N_25689,N_24837,N_24098);
nand U25690 (N_25690,N_21673,N_24215);
and U25691 (N_25691,N_23400,N_21654);
and U25692 (N_25692,N_24610,N_22128);
nand U25693 (N_25693,N_23639,N_22372);
and U25694 (N_25694,N_20456,N_24954);
or U25695 (N_25695,N_20806,N_24229);
or U25696 (N_25696,N_22387,N_21071);
or U25697 (N_25697,N_21423,N_20801);
and U25698 (N_25698,N_21324,N_20891);
nor U25699 (N_25699,N_23717,N_21414);
or U25700 (N_25700,N_22407,N_22800);
nand U25701 (N_25701,N_24069,N_20126);
and U25702 (N_25702,N_24008,N_23503);
or U25703 (N_25703,N_24667,N_21106);
and U25704 (N_25704,N_20979,N_23126);
or U25705 (N_25705,N_24534,N_23998);
nand U25706 (N_25706,N_20875,N_23885);
xnor U25707 (N_25707,N_23315,N_22573);
and U25708 (N_25708,N_20589,N_23818);
and U25709 (N_25709,N_24197,N_20642);
and U25710 (N_25710,N_22954,N_24311);
nor U25711 (N_25711,N_24872,N_22635);
nor U25712 (N_25712,N_24230,N_20047);
nand U25713 (N_25713,N_23768,N_22524);
nor U25714 (N_25714,N_23966,N_21325);
nor U25715 (N_25715,N_21156,N_22863);
and U25716 (N_25716,N_21499,N_20524);
or U25717 (N_25717,N_22283,N_20939);
nand U25718 (N_25718,N_20057,N_21790);
nand U25719 (N_25719,N_20219,N_20620);
and U25720 (N_25720,N_21769,N_20268);
xnor U25721 (N_25721,N_23835,N_23365);
xnor U25722 (N_25722,N_23066,N_24144);
xnor U25723 (N_25723,N_23294,N_21036);
nand U25724 (N_25724,N_22917,N_20965);
and U25725 (N_25725,N_21643,N_24876);
and U25726 (N_25726,N_20553,N_24540);
or U25727 (N_25727,N_21744,N_22668);
or U25728 (N_25728,N_22002,N_20651);
nor U25729 (N_25729,N_20385,N_20190);
nand U25730 (N_25730,N_24672,N_21812);
nor U25731 (N_25731,N_21385,N_22221);
xor U25732 (N_25732,N_20849,N_20611);
nor U25733 (N_25733,N_20101,N_21835);
and U25734 (N_25734,N_21780,N_22617);
or U25735 (N_25735,N_24378,N_20901);
nand U25736 (N_25736,N_24475,N_23928);
nor U25737 (N_25737,N_22168,N_20950);
nand U25738 (N_25738,N_23905,N_21331);
or U25739 (N_25739,N_22144,N_21012);
and U25740 (N_25740,N_21893,N_20132);
or U25741 (N_25741,N_22300,N_20269);
nand U25742 (N_25742,N_22208,N_20725);
nand U25743 (N_25743,N_24386,N_20527);
or U25744 (N_25744,N_22000,N_22328);
and U25745 (N_25745,N_23020,N_22811);
nor U25746 (N_25746,N_22068,N_23504);
and U25747 (N_25747,N_22500,N_22513);
xnor U25748 (N_25748,N_24947,N_21464);
and U25749 (N_25749,N_24538,N_22425);
or U25750 (N_25750,N_24616,N_21587);
nand U25751 (N_25751,N_21030,N_24634);
nor U25752 (N_25752,N_20877,N_23773);
or U25753 (N_25753,N_20395,N_24056);
nand U25754 (N_25754,N_21991,N_24806);
xnor U25755 (N_25755,N_23745,N_24289);
nand U25756 (N_25756,N_24228,N_20908);
nor U25757 (N_25757,N_22051,N_23149);
or U25758 (N_25758,N_21902,N_22603);
nor U25759 (N_25759,N_22576,N_20011);
nor U25760 (N_25760,N_20152,N_21079);
or U25761 (N_25761,N_21910,N_24911);
and U25762 (N_25762,N_20468,N_24575);
or U25763 (N_25763,N_24815,N_24708);
nand U25764 (N_25764,N_22718,N_20602);
or U25765 (N_25765,N_23875,N_22865);
and U25766 (N_25766,N_23981,N_22261);
nor U25767 (N_25767,N_23390,N_22034);
or U25768 (N_25768,N_21667,N_24476);
nand U25769 (N_25769,N_24883,N_22751);
or U25770 (N_25770,N_22819,N_22022);
nor U25771 (N_25771,N_24728,N_21213);
nand U25772 (N_25772,N_23644,N_23420);
or U25773 (N_25773,N_24286,N_20210);
nand U25774 (N_25774,N_23096,N_20779);
and U25775 (N_25775,N_24063,N_24151);
nor U25776 (N_25776,N_24492,N_22347);
and U25777 (N_25777,N_22466,N_24875);
nand U25778 (N_25778,N_20694,N_20636);
and U25779 (N_25779,N_20430,N_24485);
nand U25780 (N_25780,N_24157,N_24573);
nand U25781 (N_25781,N_22483,N_23335);
and U25782 (N_25782,N_22688,N_22735);
and U25783 (N_25783,N_21185,N_21594);
or U25784 (N_25784,N_23451,N_24225);
xnor U25785 (N_25785,N_24076,N_24734);
or U25786 (N_25786,N_21694,N_21250);
or U25787 (N_25787,N_24859,N_20669);
and U25788 (N_25788,N_20085,N_22390);
or U25789 (N_25789,N_20333,N_24438);
nand U25790 (N_25790,N_20102,N_24321);
or U25791 (N_25791,N_22134,N_21245);
nand U25792 (N_25792,N_21965,N_23933);
nand U25793 (N_25793,N_24208,N_22598);
or U25794 (N_25794,N_20671,N_21986);
nor U25795 (N_25795,N_21999,N_23045);
xor U25796 (N_25796,N_22025,N_21747);
nand U25797 (N_25797,N_22802,N_23397);
nor U25798 (N_25798,N_22226,N_20892);
nor U25799 (N_25799,N_22029,N_21877);
or U25800 (N_25800,N_20061,N_21900);
and U25801 (N_25801,N_21449,N_23092);
or U25802 (N_25802,N_21577,N_23461);
nand U25803 (N_25803,N_24087,N_24442);
nand U25804 (N_25804,N_21636,N_22893);
nor U25805 (N_25805,N_23794,N_20016);
nor U25806 (N_25806,N_20844,N_21895);
nor U25807 (N_25807,N_21649,N_21160);
nand U25808 (N_25808,N_20494,N_24821);
nor U25809 (N_25809,N_21491,N_22296);
or U25810 (N_25810,N_20060,N_24951);
nor U25811 (N_25811,N_22262,N_21454);
or U25812 (N_25812,N_23889,N_20398);
nor U25813 (N_25813,N_24629,N_22768);
and U25814 (N_25814,N_22061,N_21299);
and U25815 (N_25815,N_20485,N_21154);
or U25816 (N_25816,N_24474,N_23051);
nand U25817 (N_25817,N_21040,N_21656);
xor U25818 (N_25818,N_20969,N_22979);
and U25819 (N_25819,N_22159,N_20517);
or U25820 (N_25820,N_23174,N_21576);
nor U25821 (N_25821,N_21585,N_21719);
xor U25822 (N_25822,N_21845,N_23847);
or U25823 (N_25823,N_22175,N_24779);
and U25824 (N_25824,N_21733,N_23362);
or U25825 (N_25825,N_20195,N_20934);
nor U25826 (N_25826,N_24366,N_22335);
nand U25827 (N_25827,N_23954,N_22700);
nor U25828 (N_25828,N_22411,N_22038);
nor U25829 (N_25829,N_24256,N_21102);
nor U25830 (N_25830,N_24948,N_24952);
nor U25831 (N_25831,N_20013,N_22301);
nor U25832 (N_25832,N_21212,N_20046);
and U25833 (N_25833,N_24632,N_24958);
or U25834 (N_25834,N_24353,N_23205);
or U25835 (N_25835,N_22852,N_22491);
or U25836 (N_25836,N_20295,N_24126);
nor U25837 (N_25837,N_22694,N_24443);
and U25838 (N_25838,N_23115,N_20764);
and U25839 (N_25839,N_20170,N_20052);
and U25840 (N_25840,N_22820,N_20928);
xor U25841 (N_25841,N_24035,N_24440);
nor U25842 (N_25842,N_21811,N_21552);
nor U25843 (N_25843,N_23287,N_20867);
xnor U25844 (N_25844,N_24658,N_20317);
or U25845 (N_25845,N_24863,N_20325);
nand U25846 (N_25846,N_22190,N_24827);
nor U25847 (N_25847,N_21247,N_22436);
nand U25848 (N_25848,N_23859,N_21143);
nor U25849 (N_25849,N_24965,N_20709);
xor U25850 (N_25850,N_24847,N_24128);
xor U25851 (N_25851,N_20502,N_22150);
nor U25852 (N_25852,N_24704,N_21084);
nor U25853 (N_25853,N_23013,N_23917);
xnor U25854 (N_25854,N_23777,N_23897);
nor U25855 (N_25855,N_21031,N_23380);
or U25856 (N_25856,N_22965,N_24174);
nand U25857 (N_25857,N_21205,N_23257);
nor U25858 (N_25858,N_20902,N_22775);
and U25859 (N_25859,N_21825,N_20966);
nor U25860 (N_25860,N_20692,N_24731);
and U25861 (N_25861,N_21970,N_22967);
or U25862 (N_25862,N_24109,N_22394);
nor U25863 (N_25863,N_20041,N_22594);
or U25864 (N_25864,N_24938,N_24623);
and U25865 (N_25865,N_21909,N_24116);
or U25866 (N_25866,N_20755,N_20910);
and U25867 (N_25867,N_20000,N_23100);
xnor U25868 (N_25868,N_22558,N_24503);
nand U25869 (N_25869,N_23950,N_22386);
and U25870 (N_25870,N_21777,N_22148);
nor U25871 (N_25871,N_21629,N_22351);
or U25872 (N_25872,N_21145,N_22182);
nor U25873 (N_25873,N_21096,N_23506);
or U25874 (N_25874,N_21257,N_23018);
or U25875 (N_25875,N_21356,N_23276);
xor U25876 (N_25876,N_24387,N_21611);
nor U25877 (N_25877,N_20713,N_21588);
or U25878 (N_25878,N_22018,N_20249);
nand U25879 (N_25879,N_21359,N_24099);
or U25880 (N_25880,N_21553,N_22745);
or U25881 (N_25881,N_24408,N_22427);
nor U25882 (N_25882,N_24727,N_23121);
nand U25883 (N_25883,N_23821,N_21217);
nor U25884 (N_25884,N_23813,N_22406);
nor U25885 (N_25885,N_22643,N_21373);
or U25886 (N_25886,N_23346,N_20927);
nand U25887 (N_25887,N_20006,N_21126);
nor U25888 (N_25888,N_24486,N_23815);
nor U25889 (N_25889,N_22264,N_21310);
or U25890 (N_25890,N_23681,N_21216);
xor U25891 (N_25891,N_20348,N_21832);
or U25892 (N_25892,N_21956,N_20746);
nor U25893 (N_25893,N_22329,N_20797);
or U25894 (N_25894,N_20418,N_23788);
nor U25895 (N_25895,N_21967,N_22970);
nand U25896 (N_25896,N_24709,N_21039);
nand U25897 (N_25897,N_24636,N_24674);
nor U25898 (N_25898,N_21560,N_20439);
xnor U25899 (N_25899,N_23721,N_24768);
and U25900 (N_25900,N_23887,N_20730);
and U25901 (N_25901,N_20279,N_21878);
or U25902 (N_25902,N_20410,N_24381);
or U25903 (N_25903,N_23649,N_21120);
nand U25904 (N_25904,N_22767,N_20005);
or U25905 (N_25905,N_23147,N_22552);
and U25906 (N_25906,N_21765,N_23133);
nand U25907 (N_25907,N_22753,N_23901);
and U25908 (N_25908,N_24446,N_21019);
and U25909 (N_25909,N_22622,N_20258);
nand U25910 (N_25910,N_23849,N_22806);
nand U25911 (N_25911,N_22516,N_21028);
and U25912 (N_25912,N_22899,N_20796);
nand U25913 (N_25913,N_24427,N_23869);
and U25914 (N_25914,N_20158,N_23084);
nand U25915 (N_25915,N_21348,N_23945);
nor U25916 (N_25916,N_23033,N_20597);
nor U25917 (N_25917,N_24856,N_23502);
or U25918 (N_25918,N_20511,N_23305);
nor U25919 (N_25919,N_23189,N_21691);
or U25920 (N_25920,N_21401,N_22543);
nor U25921 (N_25921,N_24183,N_24426);
nor U25922 (N_25922,N_22941,N_23354);
or U25923 (N_25923,N_22251,N_24861);
nor U25924 (N_25924,N_23215,N_22341);
nor U25925 (N_25925,N_23169,N_20588);
or U25926 (N_25926,N_24987,N_22779);
and U25927 (N_25927,N_23304,N_23378);
nand U25928 (N_25928,N_24813,N_21693);
or U25929 (N_25929,N_21784,N_22339);
nor U25930 (N_25930,N_23766,N_22781);
nor U25931 (N_25931,N_23774,N_20703);
nand U25932 (N_25932,N_24809,N_24774);
and U25933 (N_25933,N_23268,N_20613);
or U25934 (N_25934,N_23925,N_22441);
nor U25935 (N_25935,N_20953,N_22094);
nor U25936 (N_25936,N_23999,N_21650);
nand U25937 (N_25937,N_20802,N_21971);
and U25938 (N_25938,N_21035,N_21302);
nand U25939 (N_25939,N_24041,N_23326);
nor U25940 (N_25940,N_24373,N_20541);
and U25941 (N_25941,N_23329,N_21751);
nand U25942 (N_25942,N_22275,N_20534);
or U25943 (N_25943,N_22689,N_24587);
nor U25944 (N_25944,N_23465,N_24985);
nor U25945 (N_25945,N_22918,N_24200);
or U25946 (N_25946,N_20084,N_23841);
nand U25947 (N_25947,N_23265,N_24149);
and U25948 (N_25948,N_23413,N_24974);
or U25949 (N_25949,N_20828,N_23212);
and U25950 (N_25950,N_21200,N_24100);
or U25951 (N_25951,N_20949,N_24735);
nand U25952 (N_25952,N_23248,N_23975);
nand U25953 (N_25953,N_21186,N_20135);
xnor U25954 (N_25954,N_24011,N_22043);
xnor U25955 (N_25955,N_22313,N_20336);
and U25956 (N_25956,N_22371,N_21175);
nor U25957 (N_25957,N_20499,N_22342);
or U25958 (N_25958,N_20192,N_21013);
nand U25959 (N_25959,N_24981,N_24685);
xnor U25960 (N_25960,N_21976,N_24695);
xor U25961 (N_25961,N_22599,N_24238);
or U25962 (N_25962,N_22100,N_21393);
nor U25963 (N_25963,N_20122,N_24978);
nand U25964 (N_25964,N_21383,N_22708);
nor U25965 (N_25965,N_24480,N_22198);
xnor U25966 (N_25966,N_22397,N_23186);
or U25967 (N_25967,N_23595,N_22147);
nor U25968 (N_25968,N_21901,N_24630);
or U25969 (N_25969,N_22770,N_24760);
or U25970 (N_25970,N_20148,N_24831);
nor U25971 (N_25971,N_23209,N_22256);
xor U25972 (N_25972,N_20493,N_20794);
and U25973 (N_25973,N_23763,N_23442);
nand U25974 (N_25974,N_21549,N_20909);
xnor U25975 (N_25975,N_24334,N_21670);
and U25976 (N_25976,N_22695,N_23888);
or U25977 (N_25977,N_22647,N_24639);
nor U25978 (N_25978,N_21791,N_23173);
xor U25979 (N_25979,N_23994,N_24931);
and U25980 (N_25980,N_23327,N_24325);
and U25981 (N_25981,N_22103,N_21712);
nand U25982 (N_25982,N_23009,N_22823);
or U25983 (N_25983,N_23844,N_22555);
or U25984 (N_25984,N_20655,N_20241);
and U25985 (N_25985,N_24066,N_21316);
nand U25986 (N_25986,N_24032,N_24258);
and U25987 (N_25987,N_21903,N_22234);
nor U25988 (N_25988,N_23353,N_22013);
or U25989 (N_25989,N_20391,N_24252);
nor U25990 (N_25990,N_21734,N_23958);
or U25991 (N_25991,N_24235,N_21301);
nor U25992 (N_25992,N_21679,N_23710);
nand U25993 (N_25993,N_21706,N_21319);
or U25994 (N_25994,N_23517,N_24464);
and U25995 (N_25995,N_22320,N_24239);
or U25996 (N_25996,N_24986,N_22669);
nor U25997 (N_25997,N_20071,N_21303);
xor U25998 (N_25998,N_20193,N_21666);
and U25999 (N_25999,N_21064,N_20183);
xnor U26000 (N_26000,N_21128,N_20029);
nor U26001 (N_26001,N_20372,N_23856);
and U26002 (N_26002,N_24713,N_23497);
or U26003 (N_26003,N_21263,N_22568);
nand U26004 (N_26004,N_23550,N_22330);
and U26005 (N_26005,N_24862,N_22904);
and U26006 (N_26006,N_22634,N_22821);
nand U26007 (N_26007,N_22087,N_21602);
nand U26008 (N_26008,N_23261,N_20393);
nor U26009 (N_26009,N_20839,N_24484);
and U26010 (N_26010,N_20932,N_20711);
or U26011 (N_26011,N_22417,N_20290);
or U26012 (N_26012,N_22591,N_23204);
or U26013 (N_26013,N_24420,N_23044);
nor U26014 (N_26014,N_20977,N_20668);
or U26015 (N_26015,N_22962,N_22983);
or U26016 (N_26016,N_20168,N_20570);
or U26017 (N_26017,N_20799,N_22860);
and U26018 (N_26018,N_24022,N_22578);
nand U26019 (N_26019,N_21215,N_20351);
or U26020 (N_26020,N_20201,N_21622);
nor U26021 (N_26021,N_22085,N_24992);
nand U26022 (N_26022,N_22174,N_24769);
nand U26023 (N_26023,N_21483,N_21944);
nor U26024 (N_26024,N_24932,N_22885);
nand U26025 (N_26025,N_21710,N_24497);
nor U26026 (N_26026,N_23916,N_22064);
nor U26027 (N_26027,N_21641,N_21181);
nor U26028 (N_26028,N_22604,N_22637);
or U26029 (N_26029,N_21357,N_22241);
and U26030 (N_26030,N_23807,N_20377);
and U26031 (N_26031,N_24581,N_20360);
and U26032 (N_26032,N_21799,N_22282);
nand U26033 (N_26033,N_20429,N_23725);
or U26034 (N_26034,N_20488,N_24055);
and U26035 (N_26035,N_20930,N_22471);
or U26036 (N_26036,N_21786,N_23832);
xnor U26037 (N_26037,N_22780,N_20004);
xnor U26038 (N_26038,N_23823,N_24388);
or U26039 (N_26039,N_23731,N_24425);
nand U26040 (N_26040,N_20166,N_23556);
or U26041 (N_26041,N_23555,N_22605);
and U26042 (N_26042,N_24354,N_20443);
nor U26043 (N_26043,N_23893,N_21988);
and U26044 (N_26044,N_22131,N_20287);
xor U26045 (N_26045,N_21379,N_20501);
or U26046 (N_26046,N_21498,N_24747);
nand U26047 (N_26047,N_21125,N_22984);
nor U26048 (N_26048,N_20889,N_24333);
nand U26049 (N_26049,N_23666,N_22187);
or U26050 (N_26050,N_24850,N_23317);
xor U26051 (N_26051,N_23638,N_22442);
nand U26052 (N_26052,N_22382,N_21327);
xnor U26053 (N_26053,N_23762,N_23790);
nand U26054 (N_26054,N_21544,N_20244);
nand U26055 (N_26055,N_22423,N_24122);
nor U26056 (N_26056,N_23330,N_23522);
nor U26057 (N_26057,N_22016,N_22003);
or U26058 (N_26058,N_21445,N_20687);
or U26059 (N_26059,N_24444,N_23817);
nor U26060 (N_26060,N_23661,N_24549);
and U26061 (N_26061,N_21595,N_20498);
xnor U26062 (N_26062,N_21570,N_20500);
nor U26063 (N_26063,N_24105,N_20266);
or U26064 (N_26064,N_24171,N_24342);
and U26065 (N_26065,N_23756,N_21222);
or U26066 (N_26066,N_23122,N_20114);
nor U26067 (N_26067,N_22897,N_21872);
nand U26068 (N_26068,N_24222,N_20840);
xnor U26069 (N_26069,N_20207,N_20215);
nand U26070 (N_26070,N_24869,N_20445);
or U26071 (N_26071,N_20843,N_23355);
xnor U26072 (N_26072,N_23012,N_23011);
xor U26073 (N_26073,N_21047,N_21850);
nand U26074 (N_26074,N_23309,N_20653);
nor U26075 (N_26075,N_23143,N_20448);
nand U26076 (N_26076,N_20182,N_20327);
nor U26077 (N_26077,N_23973,N_24750);
nand U26078 (N_26078,N_22801,N_24953);
xnor U26079 (N_26079,N_24090,N_22421);
nor U26080 (N_26080,N_22924,N_22938);
nor U26081 (N_26081,N_23671,N_23156);
and U26082 (N_26082,N_21374,N_24767);
nand U26083 (N_26083,N_23967,N_20270);
and U26084 (N_26084,N_22225,N_22023);
and U26085 (N_26085,N_24493,N_22053);
xor U26086 (N_26086,N_21368,N_20572);
nand U26087 (N_26087,N_22683,N_20394);
and U26088 (N_26088,N_20017,N_24800);
nor U26089 (N_26089,N_20937,N_23456);
nand U26090 (N_26090,N_22919,N_23980);
or U26091 (N_26091,N_24358,N_23119);
nand U26092 (N_26092,N_20191,N_21435);
or U26093 (N_26093,N_23699,N_24112);
xnor U26094 (N_26094,N_23622,N_23127);
nand U26095 (N_26095,N_21226,N_24389);
or U26096 (N_26096,N_20815,N_22027);
or U26097 (N_26097,N_21466,N_23234);
and U26098 (N_26098,N_22281,N_21386);
nand U26099 (N_26099,N_20789,N_23323);
or U26100 (N_26100,N_20715,N_20214);
and U26101 (N_26101,N_24919,N_20401);
and U26102 (N_26102,N_23389,N_23474);
nor U26103 (N_26103,N_20423,N_21450);
nor U26104 (N_26104,N_20254,N_24027);
nand U26105 (N_26105,N_23712,N_23310);
nor U26106 (N_26106,N_24761,N_24960);
and U26107 (N_26107,N_20677,N_24058);
and U26108 (N_26108,N_22717,N_24611);
or U26109 (N_26109,N_22156,N_22482);
nor U26110 (N_26110,N_24169,N_20560);
nor U26111 (N_26111,N_21564,N_23106);
nor U26112 (N_26112,N_23831,N_24677);
or U26113 (N_26113,N_21123,N_22533);
and U26114 (N_26114,N_22892,N_22443);
xor U26115 (N_26115,N_20554,N_23676);
or U26116 (N_26116,N_22621,N_23767);
nor U26117 (N_26117,N_22409,N_21318);
and U26118 (N_26118,N_22879,N_24759);
or U26119 (N_26119,N_20540,N_20292);
nand U26120 (N_26120,N_21892,N_20098);
nand U26121 (N_26121,N_23408,N_20807);
and U26122 (N_26122,N_20459,N_20693);
nor U26123 (N_26123,N_20637,N_23436);
nor U26124 (N_26124,N_20263,N_24053);
nand U26125 (N_26125,N_22019,N_21662);
and U26126 (N_26126,N_24141,N_21904);
nor U26127 (N_26127,N_20380,N_21259);
nor U26128 (N_26128,N_24576,N_21080);
nand U26129 (N_26129,N_23273,N_23037);
nor U26130 (N_26130,N_21896,N_22833);
and U26131 (N_26131,N_20413,N_23313);
nor U26132 (N_26132,N_20196,N_20032);
and U26133 (N_26133,N_23243,N_21456);
nand U26134 (N_26134,N_24412,N_20736);
xnor U26135 (N_26135,N_23759,N_21424);
nor U26136 (N_26136,N_22684,N_21187);
nand U26137 (N_26137,N_22648,N_24403);
or U26138 (N_26138,N_22163,N_23415);
and U26139 (N_26139,N_21070,N_22461);
or U26140 (N_26140,N_23244,N_22760);
or U26141 (N_26141,N_23412,N_24836);
and U26142 (N_26142,N_21207,N_24754);
xor U26143 (N_26143,N_23746,N_20917);
and U26144 (N_26144,N_23965,N_23201);
nor U26145 (N_26145,N_24495,N_21479);
xnor U26146 (N_26146,N_24357,N_22449);
or U26147 (N_26147,N_24941,N_24829);
or U26148 (N_26148,N_24265,N_23109);
or U26149 (N_26149,N_24527,N_21278);
xor U26150 (N_26150,N_23238,N_20154);
nor U26151 (N_26151,N_23230,N_22975);
nor U26152 (N_26152,N_20851,N_20731);
nor U26153 (N_26153,N_23804,N_24826);
and U26154 (N_26154,N_22915,N_21346);
nand U26155 (N_26155,N_22926,N_24088);
nand U26156 (N_26156,N_23250,N_23547);
or U26157 (N_26157,N_20853,N_24473);
nand U26158 (N_26158,N_21739,N_24697);
nand U26159 (N_26159,N_21350,N_22848);
nand U26160 (N_26160,N_20696,N_21463);
or U26161 (N_26161,N_22815,N_22289);
nand U26162 (N_26162,N_22338,N_23387);
nor U26163 (N_26163,N_24566,N_23300);
and U26164 (N_26164,N_21168,N_24679);
nand U26165 (N_26165,N_21890,N_22995);
nand U26166 (N_26166,N_20222,N_20389);
and U26167 (N_26167,N_24189,N_21938);
xor U26168 (N_26168,N_21151,N_20639);
xnor U26169 (N_26169,N_22772,N_20116);
nor U26170 (N_26170,N_21433,N_20894);
nor U26171 (N_26171,N_23656,N_20720);
or U26172 (N_26172,N_21367,N_20450);
or U26173 (N_26173,N_22239,N_24977);
nor U26174 (N_26174,N_24175,N_20956);
and U26175 (N_26175,N_23612,N_24959);
or U26176 (N_26176,N_23919,N_22987);
or U26177 (N_26177,N_24563,N_23240);
nand U26178 (N_26178,N_20704,N_21674);
and U26179 (N_26179,N_20260,N_23548);
nand U26180 (N_26180,N_23683,N_21352);
or U26181 (N_26181,N_21964,N_24177);
or U26182 (N_26182,N_23713,N_22143);
nand U26183 (N_26183,N_22571,N_21874);
nor U26184 (N_26184,N_24554,N_24993);
and U26185 (N_26185,N_22786,N_22333);
or U26186 (N_26186,N_24578,N_23086);
nor U26187 (N_26187,N_20109,N_24544);
nor U26188 (N_26188,N_21510,N_20863);
nand U26189 (N_26189,N_21843,N_24647);
nor U26190 (N_26190,N_23678,N_22348);
or U26191 (N_26191,N_23997,N_20719);
xor U26192 (N_26192,N_22294,N_24002);
or U26193 (N_26193,N_23545,N_23255);
nand U26194 (N_26194,N_24567,N_20324);
and U26195 (N_26195,N_23167,N_21681);
or U26196 (N_26196,N_23947,N_20223);
nor U26197 (N_26197,N_20304,N_24073);
nand U26198 (N_26198,N_20186,N_24106);
nor U26199 (N_26199,N_20198,N_24472);
or U26200 (N_26200,N_20594,N_20879);
nor U26201 (N_26201,N_24878,N_20533);
nand U26202 (N_26202,N_22452,N_21937);
nand U26203 (N_26203,N_21899,N_24641);
and U26204 (N_26204,N_24037,N_21502);
or U26205 (N_26205,N_24886,N_20251);
nor U26206 (N_26206,N_23083,N_20165);
nand U26207 (N_26207,N_24609,N_24683);
or U26208 (N_26208,N_21848,N_21391);
and U26209 (N_26209,N_20532,N_22740);
or U26210 (N_26210,N_24949,N_23843);
and U26211 (N_26211,N_22867,N_21535);
nor U26212 (N_26212,N_22506,N_24918);
nand U26213 (N_26213,N_21268,N_23360);
and U26214 (N_26214,N_22180,N_23034);
or U26215 (N_26215,N_20432,N_22880);
xnor U26216 (N_26216,N_22011,N_23752);
or U26217 (N_26217,N_22921,N_22696);
nand U26218 (N_26218,N_23489,N_21806);
nand U26219 (N_26219,N_22138,N_24936);
or U26220 (N_26220,N_20194,N_20271);
nor U26221 (N_26221,N_22367,N_21912);
nor U26222 (N_26222,N_20907,N_20513);
nor U26223 (N_26223,N_20549,N_20470);
xnor U26224 (N_26224,N_20426,N_24650);
nand U26225 (N_26225,N_20048,N_23396);
nand U26226 (N_26226,N_22395,N_23157);
or U26227 (N_26227,N_23549,N_22878);
xnor U26228 (N_26228,N_22287,N_24127);
nand U26229 (N_26229,N_22799,N_24297);
and U26230 (N_26230,N_20757,N_24203);
nand U26231 (N_26231,N_23537,N_23565);
xor U26232 (N_26232,N_20153,N_23407);
nor U26233 (N_26233,N_23026,N_24548);
nor U26234 (N_26234,N_22426,N_22844);
and U26235 (N_26235,N_21975,N_21378);
nand U26236 (N_26236,N_24891,N_22989);
nand U26237 (N_26237,N_21680,N_23603);
or U26238 (N_26238,N_23539,N_23422);
nand U26239 (N_26239,N_23241,N_20093);
or U26240 (N_26240,N_24148,N_21538);
nor U26241 (N_26241,N_24298,N_23311);
nor U26242 (N_26242,N_24152,N_22405);
nor U26243 (N_26243,N_23198,N_21771);
and U26244 (N_26244,N_23935,N_21718);
xor U26245 (N_26245,N_24367,N_20728);
nor U26246 (N_26246,N_22686,N_20707);
or U26247 (N_26247,N_21191,N_24285);
nand U26248 (N_26248,N_21888,N_20531);
xnor U26249 (N_26249,N_23728,N_21476);
and U26250 (N_26250,N_20994,N_22167);
nand U26251 (N_26251,N_24107,N_23780);
and U26252 (N_26252,N_22220,N_22186);
nor U26253 (N_26253,N_21492,N_20945);
nor U26254 (N_26254,N_24777,N_20396);
nand U26255 (N_26255,N_21018,N_21052);
or U26256 (N_26256,N_24361,N_24436);
nor U26257 (N_26257,N_24453,N_21344);
xor U26258 (N_26258,N_21272,N_22841);
nand U26259 (N_26259,N_21550,N_20149);
nand U26260 (N_26260,N_23709,N_21354);
nand U26261 (N_26261,N_24101,N_24262);
nor U26262 (N_26262,N_24887,N_24291);
nor U26263 (N_26263,N_20772,N_22613);
nand U26264 (N_26264,N_20472,N_24211);
xor U26265 (N_26265,N_22607,N_22070);
xnor U26266 (N_26266,N_24196,N_22690);
and U26267 (N_26267,N_24312,N_20504);
nor U26268 (N_26268,N_21447,N_20284);
nor U26269 (N_26269,N_22291,N_23357);
xor U26270 (N_26270,N_22284,N_22864);
nor U26271 (N_26271,N_20200,N_23112);
nor U26272 (N_26272,N_22095,N_20786);
and U26273 (N_26273,N_20357,N_21905);
or U26274 (N_26274,N_23076,N_23237);
nor U26275 (N_26275,N_24572,N_21763);
nor U26276 (N_26276,N_21924,N_23208);
nand U26277 (N_26277,N_21053,N_20850);
nand U26278 (N_26278,N_21130,N_23411);
nor U26279 (N_26279,N_23110,N_24370);
or U26280 (N_26280,N_24943,N_21664);
and U26281 (N_26281,N_24716,N_20761);
and U26282 (N_26282,N_20978,N_21689);
or U26283 (N_26283,N_20753,N_20520);
and U26284 (N_26284,N_20313,N_20569);
xor U26285 (N_26285,N_22154,N_24249);
nand U26286 (N_26286,N_20660,N_20368);
or U26287 (N_26287,N_24545,N_21104);
nand U26288 (N_26288,N_22639,N_23336);
or U26289 (N_26289,N_21887,N_21774);
or U26290 (N_26290,N_21314,N_23974);
and U26291 (N_26291,N_21775,N_24562);
nor U26292 (N_26292,N_24110,N_22944);
or U26293 (N_26293,N_24350,N_20322);
and U26294 (N_26294,N_24496,N_22032);
nand U26295 (N_26295,N_24331,N_20297);
or U26296 (N_26296,N_21275,N_21202);
xnor U26297 (N_26297,N_20859,N_21110);
nor U26298 (N_26298,N_20680,N_23879);
nor U26299 (N_26299,N_20717,N_21968);
nand U26300 (N_26300,N_23089,N_22542);
nor U26301 (N_26301,N_21057,N_21111);
xnor U26302 (N_26302,N_23747,N_23834);
and U26303 (N_26303,N_20803,N_23269);
nor U26304 (N_26304,N_23604,N_23934);
and U26305 (N_26305,N_24536,N_20575);
or U26306 (N_26306,N_21144,N_21046);
or U26307 (N_26307,N_21343,N_23221);
or U26308 (N_26308,N_23711,N_23703);
and U26309 (N_26309,N_22810,N_21860);
nor U26310 (N_26310,N_21119,N_23324);
or U26311 (N_26311,N_24523,N_24195);
xnor U26312 (N_26312,N_21941,N_24921);
or U26313 (N_26313,N_21063,N_21254);
or U26314 (N_26314,N_22040,N_21575);
xor U26315 (N_26315,N_21262,N_22200);
xor U26316 (N_26316,N_24895,N_24124);
or U26317 (N_26317,N_22804,N_21580);
or U26318 (N_26318,N_21088,N_24521);
nand U26319 (N_26319,N_24637,N_20776);
nor U26320 (N_26320,N_22790,N_20684);
and U26321 (N_26321,N_21038,N_20679);
nand U26322 (N_26322,N_22172,N_24912);
and U26323 (N_26323,N_22316,N_21930);
nor U26324 (N_26324,N_22152,N_21073);
or U26325 (N_26325,N_22428,N_23078);
nand U26326 (N_26326,N_22496,N_23964);
and U26327 (N_26327,N_20638,N_21155);
nand U26328 (N_26328,N_24799,N_23438);
nand U26329 (N_26329,N_22412,N_24546);
or U26330 (N_26330,N_20574,N_24406);
nor U26331 (N_26331,N_23239,N_20790);
nand U26332 (N_26332,N_20363,N_22547);
nand U26333 (N_26333,N_24280,N_24339);
nor U26334 (N_26334,N_20933,N_20817);
nor U26335 (N_26335,N_20876,N_20064);
or U26336 (N_26336,N_20299,N_23944);
xor U26337 (N_26337,N_23564,N_24308);
and U26338 (N_26338,N_24146,N_22822);
nor U26339 (N_26339,N_20242,N_20438);
or U26340 (N_26340,N_22318,N_22357);
nand U26341 (N_26341,N_20708,N_22857);
xnor U26342 (N_26342,N_20330,N_21347);
or U26343 (N_26343,N_23371,N_21849);
and U26344 (N_26344,N_23770,N_21614);
nand U26345 (N_26345,N_23207,N_21955);
or U26346 (N_26346,N_21507,N_21117);
and U26347 (N_26347,N_21773,N_21323);
nand U26348 (N_26348,N_23748,N_20010);
and U26349 (N_26349,N_22832,N_24786);
or U26350 (N_26350,N_23249,N_20628);
and U26351 (N_26351,N_22736,N_21048);
xnor U26352 (N_26352,N_24979,N_20778);
nor U26353 (N_26353,N_23739,N_20240);
or U26354 (N_26354,N_20714,N_23382);
or U26355 (N_26355,N_23347,N_22311);
or U26356 (N_26356,N_20565,N_22445);
and U26357 (N_26357,N_21007,N_23626);
and U26358 (N_26358,N_21284,N_22373);
and U26359 (N_26359,N_24399,N_21512);
and U26360 (N_26360,N_24619,N_23514);
or U26361 (N_26361,N_21236,N_23258);
and U26362 (N_26362,N_23402,N_22249);
and U26363 (N_26363,N_22416,N_24233);
and U26364 (N_26364,N_24310,N_23525);
and U26365 (N_26365,N_23507,N_23860);
nand U26366 (N_26366,N_23095,N_22030);
nor U26367 (N_26367,N_20175,N_24314);
nor U26368 (N_26368,N_24569,N_20605);
or U26369 (N_26369,N_24678,N_24980);
or U26370 (N_26370,N_20566,N_22890);
xor U26371 (N_26371,N_22681,N_23643);
nand U26372 (N_26372,N_22424,N_24748);
nor U26373 (N_26373,N_20283,N_20750);
nor U26374 (N_26374,N_24983,N_22583);
nand U26375 (N_26375,N_23130,N_20232);
nor U26376 (N_26376,N_22093,N_21954);
nor U26377 (N_26377,N_23245,N_22224);
or U26378 (N_26378,N_20230,N_21942);
and U26379 (N_26379,N_20792,N_21410);
nor U26380 (N_26380,N_21274,N_21950);
and U26381 (N_26381,N_21171,N_21001);
and U26382 (N_26382,N_22931,N_21309);
nand U26383 (N_26383,N_22553,N_24657);
xor U26384 (N_26384,N_21725,N_22303);
or U26385 (N_26385,N_23316,N_22324);
or U26386 (N_26386,N_20462,N_21840);
nand U26387 (N_26387,N_21886,N_24186);
nor U26388 (N_26388,N_24617,N_22398);
nand U26389 (N_26389,N_21844,N_22650);
or U26390 (N_26390,N_21244,N_24034);
or U26391 (N_26391,N_21615,N_23839);
nor U26392 (N_26392,N_24160,N_22658);
or U26393 (N_26393,N_21729,N_20040);
nor U26394 (N_26394,N_23688,N_23568);
nor U26395 (N_26395,N_24710,N_20868);
nor U26396 (N_26396,N_20855,N_21321);
nand U26397 (N_26397,N_21817,N_20199);
nor U26398 (N_26398,N_21298,N_21334);
nor U26399 (N_26399,N_20359,N_23631);
or U26400 (N_26400,N_20205,N_22646);
and U26401 (N_26401,N_22889,N_23025);
or U26402 (N_26402,N_23796,N_23321);
and U26403 (N_26403,N_21008,N_21005);
nor U26404 (N_26404,N_23492,N_23857);
nand U26405 (N_26405,N_22090,N_22212);
or U26406 (N_26406,N_21365,N_22071);
and U26407 (N_26407,N_21438,N_23213);
or U26408 (N_26408,N_23322,N_20159);
and U26409 (N_26409,N_23318,N_21265);
xor U26410 (N_26410,N_23963,N_22055);
and U26411 (N_26411,N_21947,N_23035);
or U26412 (N_26412,N_24450,N_24048);
and U26413 (N_26413,N_22532,N_24271);
and U26414 (N_26414,N_21233,N_24797);
and U26415 (N_26415,N_23870,N_24781);
nor U26416 (N_26416,N_21583,N_22608);
or U26417 (N_26417,N_24688,N_22675);
xnor U26418 (N_26418,N_23405,N_23246);
nand U26419 (N_26419,N_21484,N_20518);
nand U26420 (N_26420,N_21736,N_22929);
nor U26421 (N_26421,N_23730,N_20948);
nand U26422 (N_26422,N_24084,N_23452);
or U26423 (N_26423,N_24842,N_20255);
nand U26424 (N_26424,N_24822,N_24043);
or U26425 (N_26425,N_24108,N_21416);
nand U26426 (N_26426,N_23803,N_23184);
or U26427 (N_26427,N_21642,N_21473);
nand U26428 (N_26428,N_22710,N_23840);
or U26429 (N_26429,N_21462,N_23943);
or U26430 (N_26430,N_21782,N_20926);
nor U26431 (N_26431,N_23284,N_23496);
and U26432 (N_26432,N_23809,N_20936);
xor U26433 (N_26433,N_22213,N_20386);
nor U26434 (N_26434,N_22887,N_22759);
nor U26435 (N_26435,N_22137,N_24355);
nand U26436 (N_26436,N_22704,N_21103);
nand U26437 (N_26437,N_20577,N_21405);
nand U26438 (N_26438,N_22557,N_20619);
nor U26439 (N_26439,N_22551,N_23005);
nor U26440 (N_26440,N_20234,N_20397);
nor U26441 (N_26441,N_24896,N_24394);
or U26442 (N_26442,N_22473,N_21330);
and U26443 (N_26443,N_23684,N_23558);
nor U26444 (N_26444,N_22245,N_23827);
or U26445 (N_26445,N_22054,N_20136);
nand U26446 (N_26446,N_23418,N_21169);
nor U26447 (N_26447,N_21136,N_23695);
nor U26448 (N_26448,N_24253,N_22831);
xnor U26449 (N_26449,N_24968,N_23719);
and U26450 (N_26450,N_21783,N_20551);
nand U26451 (N_26451,N_24163,N_24374);
nor U26452 (N_26452,N_20685,N_21443);
and U26453 (N_26453,N_20044,N_24892);
and U26454 (N_26454,N_23014,N_20142);
or U26455 (N_26455,N_24451,N_20900);
xor U26456 (N_26456,N_22855,N_24145);
and U26457 (N_26457,N_23057,N_23178);
and U26458 (N_26458,N_24064,N_23226);
and U26459 (N_26459,N_20012,N_22419);
and U26460 (N_26460,N_22705,N_20732);
or U26461 (N_26461,N_21296,N_22847);
and U26462 (N_26462,N_22507,N_24470);
and U26463 (N_26463,N_23200,N_23180);
and U26464 (N_26464,N_20033,N_23129);
and U26465 (N_26465,N_22049,N_24586);
or U26466 (N_26466,N_23431,N_21115);
nor U26467 (N_26467,N_21722,N_22127);
nor U26468 (N_26468,N_20139,N_20366);
nand U26469 (N_26469,N_20646,N_21364);
nand U26470 (N_26470,N_23810,N_23338);
nand U26471 (N_26471,N_20793,N_22829);
or U26472 (N_26472,N_22240,N_20070);
nor U26473 (N_26473,N_22375,N_22048);
nand U26474 (N_26474,N_20681,N_22184);
or U26475 (N_26475,N_20043,N_21494);
and U26476 (N_26476,N_21646,N_20931);
or U26477 (N_26477,N_22399,N_20782);
xnor U26478 (N_26478,N_21652,N_22873);
nor U26479 (N_26479,N_22408,N_24129);
or U26480 (N_26480,N_22227,N_21599);
xor U26481 (N_26481,N_21010,N_24705);
or U26482 (N_26482,N_21684,N_23289);
nand U26483 (N_26483,N_23254,N_22935);
or U26484 (N_26484,N_21794,N_22805);
and U26485 (N_26485,N_24682,N_20455);
or U26486 (N_26486,N_21159,N_20131);
xor U26487 (N_26487,N_24915,N_24380);
nand U26488 (N_26488,N_23485,N_24601);
and U26489 (N_26489,N_20224,N_24046);
or U26490 (N_26490,N_21523,N_24332);
nand U26491 (N_26491,N_22765,N_21610);
and U26492 (N_26492,N_23733,N_20691);
or U26493 (N_26493,N_20453,N_21836);
or U26494 (N_26494,N_22750,N_21651);
nand U26495 (N_26495,N_24125,N_23805);
nand U26496 (N_26496,N_22059,N_22730);
nand U26497 (N_26497,N_22102,N_24455);
and U26498 (N_26498,N_23769,N_22587);
or U26499 (N_26499,N_21338,N_24561);
or U26500 (N_26500,N_22456,N_24382);
and U26501 (N_26501,N_20035,N_23242);
nor U26502 (N_26502,N_22122,N_21015);
and U26503 (N_26503,N_21880,N_22403);
nand U26504 (N_26504,N_20262,N_20414);
nor U26505 (N_26505,N_23952,N_23535);
xor U26506 (N_26506,N_20981,N_21536);
nand U26507 (N_26507,N_20871,N_23486);
nand U26508 (N_26508,N_21307,N_23714);
nand U26509 (N_26509,N_21916,N_21085);
nand U26510 (N_26510,N_24933,N_22422);
or U26511 (N_26511,N_21069,N_24564);
nor U26512 (N_26512,N_22713,N_20808);
nand U26513 (N_26513,N_21228,N_21029);
xor U26514 (N_26514,N_21822,N_23376);
or U26515 (N_26515,N_22503,N_21051);
or U26516 (N_26516,N_23927,N_24263);
nor U26517 (N_26517,N_20957,N_20562);
and U26518 (N_26518,N_23094,N_21116);
or U26519 (N_26519,N_24870,N_22345);
or U26520 (N_26520,N_22600,N_20227);
xnor U26521 (N_26521,N_24749,N_24201);
or U26522 (N_26522,N_23314,N_22808);
nor U26523 (N_26523,N_22273,N_23286);
and U26524 (N_26524,N_23233,N_23693);
or U26525 (N_26525,N_23576,N_22943);
or U26526 (N_26526,N_22196,N_20798);
or U26527 (N_26527,N_23679,N_21011);
nor U26528 (N_26528,N_23969,N_21514);
nand U26529 (N_26529,N_22366,N_21482);
xnor U26530 (N_26530,N_21496,N_24764);
nand U26531 (N_26531,N_23223,N_21669);
and U26532 (N_26532,N_23776,N_22788);
nand U26533 (N_26533,N_23168,N_22092);
nand U26534 (N_26534,N_23510,N_20463);
or U26535 (N_26535,N_23369,N_20920);
nor U26536 (N_26536,N_20447,N_21866);
nor U26537 (N_26537,N_23579,N_20189);
or U26538 (N_26538,N_23898,N_20409);
nor U26539 (N_26539,N_24432,N_24843);
and U26540 (N_26540,N_24322,N_21628);
nand U26541 (N_26541,N_22279,N_21113);
xnor U26542 (N_26542,N_23757,N_21025);
and U26543 (N_26543,N_21311,N_21994);
xnor U26544 (N_26544,N_24720,N_20296);
or U26545 (N_26545,N_20813,N_22189);
xor U26546 (N_26546,N_24429,N_24347);
nand U26547 (N_26547,N_22766,N_21601);
nand U26548 (N_26548,N_20431,N_24966);
xor U26549 (N_26549,N_23059,N_23394);
or U26550 (N_26550,N_20525,N_23532);
or U26551 (N_26551,N_20652,N_20962);
xnor U26552 (N_26552,N_20905,N_22541);
or U26553 (N_26553,N_23363,N_23495);
and U26554 (N_26554,N_22081,N_20885);
nand U26555 (N_26555,N_22843,N_22771);
nand U26556 (N_26556,N_23921,N_24020);
and U26557 (N_26557,N_20457,N_20341);
nand U26558 (N_26558,N_22529,N_21603);
xnor U26559 (N_26559,N_21558,N_20312);
nand U26560 (N_26560,N_22976,N_22460);
and U26561 (N_26561,N_23476,N_20545);
and U26562 (N_26562,N_23743,N_24740);
or U26563 (N_26563,N_23566,N_20586);
or U26564 (N_26564,N_24962,N_24300);
nand U26565 (N_26565,N_23166,N_23523);
nor U26566 (N_26566,N_20454,N_20810);
or U26567 (N_26567,N_22561,N_20293);
and U26568 (N_26568,N_24770,N_24998);
or U26569 (N_26569,N_23124,N_21208);
nor U26570 (N_26570,N_21841,N_22299);
nand U26571 (N_26571,N_23183,N_23513);
nand U26572 (N_26572,N_21406,N_21983);
and U26573 (N_26573,N_24404,N_21898);
nand U26574 (N_26574,N_22304,N_24621);
or U26575 (N_26575,N_23836,N_22697);
and U26576 (N_26576,N_23301,N_20795);
nand U26577 (N_26577,N_24224,N_24656);
and U26578 (N_26578,N_23806,N_21908);
nor U26579 (N_26579,N_22737,N_22540);
xor U26580 (N_26580,N_21852,N_21658);
nor U26581 (N_26581,N_20475,N_22522);
and U26582 (N_26582,N_21884,N_23391);
xnor U26583 (N_26583,N_20701,N_24130);
xor U26584 (N_26584,N_23253,N_24972);
nand U26585 (N_26585,N_23480,N_22660);
or U26586 (N_26586,N_21419,N_24512);
or U26587 (N_26587,N_20339,N_24955);
and U26588 (N_26588,N_24391,N_22657);
nor U26589 (N_26589,N_20117,N_20756);
xnor U26590 (N_26590,N_22739,N_21183);
xnor U26591 (N_26591,N_23150,N_22994);
xnor U26592 (N_26592,N_22531,N_22045);
and U26593 (N_26593,N_21062,N_21206);
nor U26594 (N_26594,N_21190,N_24868);
or U26595 (N_26595,N_24603,N_23483);
xnor U26596 (N_26596,N_20997,N_23334);
and U26597 (N_26597,N_20315,N_22376);
and U26598 (N_26598,N_22749,N_22937);
or U26599 (N_26599,N_21177,N_20009);
nor U26600 (N_26600,N_23488,N_21397);
or U26601 (N_26601,N_22818,N_23512);
or U26602 (N_26602,N_24479,N_20209);
or U26603 (N_26603,N_20523,N_22204);
nand U26604 (N_26604,N_22951,N_22539);
nand U26605 (N_26605,N_20376,N_20702);
or U26606 (N_26606,N_21161,N_23434);
or U26607 (N_26607,N_20134,N_20526);
and U26608 (N_26608,N_24681,N_22112);
xor U26609 (N_26609,N_20460,N_24626);
nor U26610 (N_26610,N_21638,N_20187);
nand U26611 (N_26611,N_24320,N_21260);
nand U26612 (N_26612,N_22026,N_22964);
and U26613 (N_26613,N_24659,N_20748);
nand U26614 (N_26614,N_22579,N_23097);
nand U26615 (N_26615,N_24547,N_22400);
nand U26616 (N_26616,N_24607,N_21112);
nand U26617 (N_26617,N_21469,N_20075);
nand U26618 (N_26618,N_23370,N_20547);
and U26619 (N_26619,N_23858,N_21533);
nand U26620 (N_26620,N_20784,N_22922);
nand U26621 (N_26621,N_20220,N_21605);
nand U26622 (N_26622,N_20476,N_22927);
nand U26623 (N_26623,N_22725,N_24592);
or U26624 (N_26624,N_24594,N_22438);
nand U26625 (N_26625,N_22084,N_20584);
and U26626 (N_26626,N_24267,N_21032);
or U26627 (N_26627,N_21056,N_23052);
nand U26628 (N_26628,N_21701,N_23125);
nand U26629 (N_26629,N_20328,N_22077);
nand U26630 (N_26630,N_21920,N_22106);
nor U26631 (N_26631,N_23036,N_21527);
nand U26632 (N_26632,N_21963,N_23972);
nor U26633 (N_26633,N_23306,N_24247);
nor U26634 (N_26634,N_20573,N_21467);
nor U26635 (N_26635,N_22151,N_23574);
nand U26636 (N_26636,N_22378,N_20208);
nand U26637 (N_26637,N_21761,N_21943);
nand U26638 (N_26638,N_23586,N_20002);
nand U26639 (N_26639,N_21856,N_24187);
nand U26640 (N_26640,N_21153,N_23990);
and U26641 (N_26641,N_21077,N_24798);
nor U26642 (N_26642,N_20673,N_21940);
or U26643 (N_26643,N_20247,N_23319);
xnor U26644 (N_26644,N_20353,N_20921);
nand U26645 (N_26645,N_23930,N_20747);
and U26646 (N_26646,N_20958,N_20473);
or U26647 (N_26647,N_21501,N_24542);
or U26648 (N_26648,N_23585,N_21933);
nand U26649 (N_26649,N_24288,N_20989);
nor U26650 (N_26650,N_22017,N_22118);
or U26651 (N_26651,N_22280,N_23056);
and U26652 (N_26652,N_21002,N_23942);
xor U26653 (N_26653,N_22458,N_20895);
or U26654 (N_26654,N_22977,N_20288);
nand U26655 (N_26655,N_24221,N_24852);
nor U26656 (N_26656,N_20825,N_22171);
or U26657 (N_26657,N_21726,N_21853);
or U26658 (N_26658,N_20309,N_20121);
and U26659 (N_26659,N_24526,N_23959);
nand U26660 (N_26660,N_24093,N_23938);
xor U26661 (N_26661,N_22711,N_23464);
and U26662 (N_26662,N_24491,N_22465);
or U26663 (N_26663,N_22217,N_24047);
and U26664 (N_26664,N_23741,N_22310);
xnor U26665 (N_26665,N_24324,N_20614);
and U26666 (N_26666,N_22615,N_21951);
nor U26667 (N_26667,N_22430,N_23628);
nor U26668 (N_26668,N_21862,N_24383);
nor U26669 (N_26669,N_23646,N_24517);
and U26670 (N_26670,N_20992,N_20151);
or U26671 (N_26671,N_21770,N_24458);
nand U26672 (N_26672,N_20471,N_22082);
nand U26673 (N_26673,N_20744,N_22527);
nor U26674 (N_26674,N_20248,N_22945);
or U26675 (N_26675,N_21855,N_23218);
nor U26676 (N_26676,N_24614,N_24990);
and U26677 (N_26677,N_24468,N_23599);
nor U26678 (N_26678,N_24001,N_22559);
or U26679 (N_26679,N_24182,N_23171);
xor U26680 (N_26680,N_24220,N_23508);
and U26681 (N_26681,N_20635,N_20913);
nand U26682 (N_26682,N_20173,N_21400);
nand U26683 (N_26683,N_21714,N_22178);
or U26684 (N_26684,N_24773,N_24241);
nand U26685 (N_26685,N_21561,N_22197);
nand U26686 (N_26686,N_22041,N_20984);
nor U26687 (N_26687,N_24018,N_24287);
or U26688 (N_26688,N_20281,N_23800);
nor U26689 (N_26689,N_23554,N_24702);
nor U26690 (N_26690,N_21926,N_23750);
and U26691 (N_26691,N_24967,N_24920);
nor U26692 (N_26692,N_23165,N_24435);
nand U26693 (N_26693,N_22791,N_24613);
xnor U26694 (N_26694,N_21619,N_22949);
nand U26695 (N_26695,N_24997,N_23440);
nor U26696 (N_26696,N_22108,N_21521);
nor U26697 (N_26697,N_23280,N_20343);
and U26698 (N_26698,N_20865,N_21065);
and U26699 (N_26699,N_24498,N_21597);
nor U26700 (N_26700,N_24746,N_24337);
and U26701 (N_26701,N_24392,N_20127);
nor U26702 (N_26702,N_20847,N_20971);
nor U26703 (N_26703,N_24433,N_24029);
or U26704 (N_26704,N_24074,N_24711);
and U26705 (N_26705,N_21415,N_20362);
and U26706 (N_26706,N_21292,N_21221);
xnor U26707 (N_26707,N_22519,N_24784);
and U26708 (N_26708,N_21439,N_24164);
nor U26709 (N_26709,N_22866,N_24897);
and U26710 (N_26710,N_20788,N_21565);
nand U26711 (N_26711,N_24937,N_21179);
nand U26712 (N_26712,N_24907,N_22340);
xnor U26713 (N_26713,N_21990,N_21409);
and U26714 (N_26714,N_21745,N_24326);
xnor U26715 (N_26715,N_22562,N_21946);
nor U26716 (N_26716,N_22271,N_22252);
xnor U26717 (N_26717,N_24642,N_22777);
xor U26718 (N_26718,N_20745,N_21204);
nand U26719 (N_26719,N_24045,N_23177);
nand U26720 (N_26720,N_20275,N_20539);
nand U26721 (N_26721,N_23597,N_23260);
and U26722 (N_26722,N_23352,N_22343);
nand U26723 (N_26723,N_21306,N_21752);
nor U26724 (N_26724,N_20095,N_21524);
nor U26725 (N_26725,N_24645,N_23623);
nand U26726 (N_26726,N_21329,N_20985);
or U26727 (N_26727,N_24909,N_23793);
or U26728 (N_26728,N_23765,N_23573);
nand U26729 (N_26729,N_24864,N_20783);
nand U26730 (N_26730,N_20542,N_21515);
and U26731 (N_26731,N_21460,N_20466);
nand U26732 (N_26732,N_22738,N_24033);
xnor U26733 (N_26733,N_22589,N_21376);
or U26734 (N_26734,N_23685,N_22258);
xor U26735 (N_26735,N_24635,N_23325);
nor U26736 (N_26736,N_20963,N_22269);
xnor U26737 (N_26737,N_21581,N_23531);
nor U26738 (N_26738,N_21335,N_21731);
and U26739 (N_26739,N_24509,N_23970);
nor U26740 (N_26740,N_22007,N_20301);
nand U26741 (N_26741,N_24733,N_24078);
nand U26742 (N_26742,N_21458,N_21634);
nand U26743 (N_26743,N_20291,N_22554);
nor U26744 (N_26744,N_23421,N_24640);
nor U26745 (N_26745,N_21672,N_24556);
and U26746 (N_26746,N_24232,N_22047);
and U26747 (N_26747,N_21300,N_24166);
and U26748 (N_26748,N_24279,N_22535);
or U26749 (N_26749,N_21055,N_22687);
nor U26750 (N_26750,N_22850,N_22654);
nand U26751 (N_26751,N_21178,N_23785);
or U26752 (N_26752,N_22067,N_20027);
nand U26753 (N_26753,N_24689,N_20982);
and U26754 (N_26754,N_20781,N_21488);
or U26755 (N_26755,N_24070,N_22920);
xor U26756 (N_26756,N_20406,N_22383);
and U26757 (N_26757,N_20346,N_24445);
or U26758 (N_26758,N_20592,N_24136);
and U26759 (N_26759,N_22083,N_21293);
or U26760 (N_26760,N_24038,N_21059);
or U26761 (N_26761,N_21101,N_23085);
and U26762 (N_26762,N_22356,N_21097);
nor U26763 (N_26763,N_21948,N_21660);
nand U26764 (N_26764,N_20144,N_20018);
nor U26765 (N_26765,N_21738,N_20846);
or U26766 (N_26766,N_22676,N_23079);
nand U26767 (N_26767,N_22884,N_21098);
nor U26768 (N_26768,N_24091,N_21592);
xnor U26769 (N_26769,N_21922,N_23742);
or U26770 (N_26770,N_23187,N_22816);
xnor U26771 (N_26771,N_21086,N_20596);
nand U26772 (N_26772,N_24858,N_23701);
and U26773 (N_26773,N_22104,N_20820);
xnor U26774 (N_26774,N_22691,N_23191);
or U26775 (N_26775,N_24928,N_23104);
nand U26776 (N_26776,N_24865,N_21258);
xnor U26777 (N_26777,N_21740,N_23593);
nand U26778 (N_26778,N_22911,N_21256);
nor U26779 (N_26779,N_21563,N_24668);
and U26780 (N_26780,N_23275,N_20440);
nor U26781 (N_26781,N_20609,N_22715);
or U26782 (N_26782,N_23010,N_22285);
nor U26783 (N_26783,N_21809,N_20923);
and U26784 (N_26784,N_20419,N_24418);
and U26785 (N_26785,N_24123,N_22380);
and U26786 (N_26786,N_20861,N_22741);
or U26787 (N_26787,N_23572,N_20959);
nor U26788 (N_26788,N_21556,N_20780);
nor U26789 (N_26789,N_20682,N_24190);
nor U26790 (N_26790,N_24273,N_20318);
nand U26791 (N_26791,N_24255,N_21081);
and U26792 (N_26792,N_23826,N_22909);
nor U26793 (N_26793,N_23414,N_23995);
nor U26794 (N_26794,N_24816,N_23672);
and U26795 (N_26795,N_21459,N_24776);
nand U26796 (N_26796,N_20184,N_23383);
nor U26797 (N_26797,N_23527,N_23155);
or U26798 (N_26798,N_20659,N_22856);
nand U26799 (N_26799,N_21506,N_23142);
nand U26800 (N_26800,N_24633,N_22031);
nand U26801 (N_26801,N_20632,N_23267);
or U26802 (N_26802,N_24137,N_24596);
xor U26803 (N_26803,N_20537,N_22350);
nor U26804 (N_26804,N_22099,N_23736);
nand U26805 (N_26805,N_24185,N_24006);
or U26806 (N_26806,N_22883,N_23441);
nor U26807 (N_26807,N_22974,N_24543);
nor U26808 (N_26808,N_22871,N_23923);
nor U26809 (N_26809,N_22582,N_22947);
nor U26810 (N_26810,N_24877,N_22141);
nor U26811 (N_26811,N_20155,N_23403);
or U26812 (N_26812,N_20062,N_22451);
and U26813 (N_26813,N_20107,N_20355);
nor U26814 (N_26814,N_22413,N_21004);
or U26815 (N_26815,N_23798,N_21090);
and U26816 (N_26816,N_23559,N_21219);
nand U26817 (N_26817,N_21384,N_22755);
and U26818 (N_26818,N_21135,N_22692);
or U26819 (N_26819,N_21923,N_22052);
nand U26820 (N_26820,N_20492,N_21863);
or U26821 (N_26821,N_23073,N_20860);
xor U26822 (N_26822,N_20903,N_23158);
and U26823 (N_26823,N_24102,N_21091);
and U26824 (N_26824,N_22429,N_20897);
nand U26825 (N_26825,N_24340,N_23874);
or U26826 (N_26826,N_24010,N_24757);
or U26827 (N_26827,N_21453,N_21708);
nand U26828 (N_26828,N_24410,N_24042);
or U26829 (N_26829,N_21173,N_22778);
nand U26830 (N_26830,N_23557,N_23067);
nor U26831 (N_26831,N_22309,N_23468);
or U26832 (N_26832,N_20252,N_22898);
or U26833 (N_26833,N_21412,N_20034);
nor U26834 (N_26834,N_20174,N_22923);
or U26835 (N_26835,N_22115,N_22742);
or U26836 (N_26836,N_22244,N_20561);
nor U26837 (N_26837,N_24362,N_21252);
or U26838 (N_26838,N_20626,N_21166);
nor U26839 (N_26839,N_24009,N_24893);
nor U26840 (N_26840,N_22757,N_24916);
xnor U26841 (N_26841,N_20021,N_22444);
or U26842 (N_26842,N_22896,N_24062);
nand U26843 (N_26843,N_24328,N_21380);
and U26844 (N_26844,N_23417,N_21375);
nand U26845 (N_26845,N_20261,N_20741);
and U26846 (N_26846,N_20078,N_20150);
or U26847 (N_26847,N_21024,N_20178);
nor U26848 (N_26848,N_20086,N_24304);
xor U26849 (N_26849,N_20616,N_20108);
nand U26850 (N_26850,N_20112,N_22353);
or U26851 (N_26851,N_23061,N_21058);
nor U26852 (N_26852,N_21349,N_22183);
nor U26853 (N_26853,N_22731,N_21408);
nand U26854 (N_26854,N_20664,N_23589);
nand U26855 (N_26855,N_23132,N_20740);
or U26856 (N_26856,N_21620,N_20007);
and U26857 (N_26857,N_20054,N_21993);
xnor U26858 (N_26858,N_22331,N_22756);
and U26859 (N_26859,N_22501,N_20951);
or U26860 (N_26860,N_21016,N_22826);
nand U26861 (N_26861,N_23553,N_24346);
and U26862 (N_26862,N_23256,N_22437);
nor U26863 (N_26863,N_22161,N_23802);
nor U26864 (N_26864,N_20621,N_21006);
or U26865 (N_26865,N_21478,N_23749);
and U26866 (N_26866,N_22593,N_23484);
nand U26867 (N_26867,N_24721,N_23778);
xor U26868 (N_26868,N_22785,N_23416);
and U26869 (N_26869,N_21702,N_20437);
nand U26870 (N_26870,N_22136,N_20912);
xnor U26871 (N_26871,N_21532,N_20873);
nand U26872 (N_26872,N_24402,N_23015);
and U26873 (N_26873,N_20922,N_23445);
xnor U26874 (N_26874,N_20538,N_21180);
and U26875 (N_26875,N_21049,N_22988);
or U26876 (N_26876,N_20495,N_21290);
or U26877 (N_26877,N_20179,N_21249);
and U26878 (N_26878,N_21490,N_24676);
and U26879 (N_26879,N_22628,N_22257);
nand U26880 (N_26880,N_22062,N_24551);
nand U26881 (N_26881,N_22248,N_23538);
nand U26882 (N_26882,N_24198,N_24319);
or U26883 (N_26883,N_24758,N_24384);
xnor U26884 (N_26884,N_24686,N_24973);
and U26885 (N_26885,N_20858,N_21432);
nor U26886 (N_26886,N_21072,N_21246);
or U26887 (N_26887,N_20878,N_21721);
nor U26888 (N_26888,N_21317,N_24167);
or U26889 (N_26889,N_24159,N_21276);
nor U26890 (N_26890,N_21596,N_20904);
nor U26891 (N_26891,N_24571,N_23830);
and U26892 (N_26892,N_22796,N_20467);
nor U26893 (N_26893,N_20940,N_24851);
nand U26894 (N_26894,N_22479,N_20405);
nand U26895 (N_26895,N_24557,N_24818);
and U26896 (N_26896,N_24368,N_24722);
or U26897 (N_26897,N_21214,N_24999);
nand U26898 (N_26898,N_23292,N_23904);
and U26899 (N_26899,N_23374,N_22063);
or U26900 (N_26900,N_24218,N_23162);
nor U26901 (N_26901,N_21578,N_21609);
nor U26902 (N_26902,N_20289,N_24820);
xor U26903 (N_26903,N_23588,N_23808);
nor U26904 (N_26904,N_21883,N_22932);
and U26905 (N_26905,N_24459,N_21838);
and U26906 (N_26906,N_22876,N_22812);
nand U26907 (N_26907,N_21248,N_23932);
nand U26908 (N_26908,N_21411,N_23782);
and U26909 (N_26909,N_23653,N_22133);
nor U26910 (N_26910,N_24690,N_24719);
nor U26911 (N_26911,N_22377,N_23682);
nand U26912 (N_26912,N_22728,N_23792);
or U26913 (N_26913,N_20049,N_23575);
or U26914 (N_26914,N_21977,N_23349);
nand U26915 (N_26915,N_20329,N_24336);
and U26916 (N_26916,N_23694,N_22851);
nand U26917 (N_26917,N_20024,N_22837);
nand U26918 (N_26918,N_24371,N_24096);
and U26919 (N_26919,N_20143,N_24646);
xnor U26920 (N_26920,N_24910,N_21668);
or U26921 (N_26921,N_20610,N_20631);
and U26922 (N_26922,N_21355,N_21163);
and U26923 (N_26923,N_23341,N_22930);
or U26924 (N_26924,N_24706,N_24481);
nor U26925 (N_26925,N_20056,N_23571);
or U26926 (N_26926,N_22505,N_20942);
nor U26927 (N_26927,N_23915,N_20067);
and U26928 (N_26928,N_22078,N_22537);
and U26929 (N_26929,N_24456,N_24739);
xor U26930 (N_26930,N_22158,N_23528);
nand U26931 (N_26931,N_20618,N_23006);
nor U26932 (N_26932,N_23509,N_20257);
nor U26933 (N_26933,N_24044,N_22538);
xor U26934 (N_26934,N_23214,N_22769);
or U26935 (N_26935,N_24216,N_22160);
nor U26936 (N_26936,N_21095,N_21455);
and U26937 (N_26937,N_21017,N_22459);
or U26938 (N_26938,N_22521,N_21911);
nand U26939 (N_26939,N_22614,N_24315);
and U26940 (N_26940,N_22928,N_20721);
nand U26941 (N_26941,N_24293,N_22714);
nor U26942 (N_26942,N_22509,N_22370);
nand U26943 (N_26943,N_22698,N_24057);
xnor U26944 (N_26944,N_21427,N_24039);
and U26945 (N_26945,N_21061,N_23063);
or U26946 (N_26946,N_22567,N_21326);
or U26947 (N_26947,N_21210,N_23482);
nand U26948 (N_26948,N_22058,N_24589);
xor U26949 (N_26949,N_22230,N_22834);
or U26950 (N_26950,N_23625,N_20162);
xor U26951 (N_26951,N_22721,N_22132);
nand U26952 (N_26952,N_23948,N_23117);
nand U26953 (N_26953,N_20522,N_24085);
nor U26954 (N_26954,N_24030,N_20300);
or U26955 (N_26955,N_22250,N_23861);
nand U26956 (N_26956,N_20484,N_22992);
or U26957 (N_26957,N_20612,N_21264);
nand U26958 (N_26958,N_23873,N_23139);
and U26959 (N_26959,N_21195,N_23295);
and U26960 (N_26960,N_23113,N_23105);
nor U26961 (N_26961,N_21803,N_23991);
nor U26962 (N_26962,N_22363,N_23501);
nand U26963 (N_26963,N_22266,N_20946);
or U26964 (N_26964,N_23716,N_20442);
nor U26965 (N_26965,N_24588,N_23786);
xor U26966 (N_26966,N_22164,N_21653);
xor U26967 (N_26967,N_21291,N_22246);
and U26968 (N_26968,N_21295,N_23194);
and U26969 (N_26969,N_20629,N_21754);
or U26970 (N_26970,N_24133,N_21225);
nor U26971 (N_26971,N_23299,N_23048);
nor U26972 (N_26972,N_20436,N_24023);
nor U26973 (N_26973,N_20303,N_20718);
and U26974 (N_26974,N_20599,N_23615);
and U26975 (N_26975,N_22402,N_22631);
and U26976 (N_26976,N_20274,N_23195);
nand U26977 (N_26977,N_21172,N_22874);
nor U26978 (N_26978,N_23398,N_20773);
nor U26979 (N_26979,N_24237,N_24452);
nor U26980 (N_26980,N_22773,N_20976);
nor U26981 (N_26981,N_23019,N_22468);
or U26982 (N_26982,N_22845,N_23976);
and U26983 (N_26983,N_24161,N_23331);
and U26984 (N_26984,N_22124,N_23266);
or U26985 (N_26985,N_23674,N_23031);
nor U26986 (N_26986,N_21717,N_23519);
and U26987 (N_26987,N_21949,N_21889);
nand U26988 (N_26988,N_23091,N_20307);
nor U26989 (N_26989,N_20399,N_21165);
and U26990 (N_26990,N_20727,N_24414);
nor U26991 (N_26991,N_21969,N_20749);
or U26992 (N_26992,N_24155,N_23530);
xor U26993 (N_26993,N_21998,N_21875);
nor U26994 (N_26994,N_24666,N_23196);
nor U26995 (N_26995,N_20698,N_24835);
nand U26996 (N_26996,N_22958,N_20358);
nor U26997 (N_26997,N_20528,N_23308);
or U26998 (N_26998,N_21237,N_20890);
xor U26999 (N_26999,N_23895,N_23619);
nand U27000 (N_27000,N_20213,N_21034);
or U27001 (N_27001,N_23140,N_23988);
and U27002 (N_27002,N_23203,N_23232);
and U27003 (N_27003,N_23071,N_24080);
nand U27004 (N_27004,N_24671,N_23131);
xnor U27005 (N_27005,N_24007,N_20831);
nand U27006 (N_27006,N_24874,N_22162);
or U27007 (N_27007,N_24103,N_22836);
and U27008 (N_27008,N_22169,N_23939);
nor U27009 (N_27009,N_24790,N_21861);
and U27010 (N_27010,N_20176,N_22086);
nor U27011 (N_27011,N_23297,N_22121);
or U27012 (N_27012,N_20337,N_22455);
or U27013 (N_27013,N_22297,N_23367);
and U27014 (N_27014,N_20356,N_24083);
and U27015 (N_27015,N_24844,N_22385);
nor U27016 (N_27016,N_21500,N_20852);
and U27017 (N_27017,N_22733,N_20119);
nor U27018 (N_27018,N_21572,N_20147);
and U27019 (N_27019,N_23583,N_21513);
nand U27020 (N_27020,N_24522,N_20087);
and U27021 (N_27021,N_21829,N_21687);
or U27022 (N_27022,N_20014,N_22862);
nor U27023 (N_27023,N_20624,N_21624);
or U27024 (N_27024,N_21868,N_20854);
and U27025 (N_27025,N_21511,N_22916);
and U27026 (N_27026,N_24885,N_24372);
nand U27027 (N_27027,N_23824,N_22640);
nand U27028 (N_27028,N_20670,N_21371);
or U27029 (N_27029,N_23163,N_23822);
xor U27030 (N_27030,N_23570,N_20482);
and U27031 (N_27031,N_24730,N_24060);
xor U27032 (N_27032,N_24755,N_22265);
nor U27033 (N_27033,N_24751,N_20752);
xor U27034 (N_27034,N_20536,N_23298);
or U27035 (N_27035,N_20961,N_22414);
and U27036 (N_27036,N_22374,N_21134);
nor U27037 (N_27037,N_24226,N_22478);
or U27038 (N_27038,N_22323,N_23899);
nand U27039 (N_27039,N_22470,N_22707);
nand U27040 (N_27040,N_21865,N_23023);
and U27041 (N_27041,N_24385,N_23772);
xor U27042 (N_27042,N_23004,N_21644);
or U27043 (N_27043,N_20285,N_23602);
or U27044 (N_27044,N_23664,N_22272);
xor U27045 (N_27045,N_21461,N_24555);
nor U27046 (N_27046,N_22410,N_21437);
nor U27047 (N_27047,N_23775,N_20938);
nor U27048 (N_27048,N_23088,N_23641);
or U27049 (N_27049,N_20106,N_24111);
or U27050 (N_27050,N_20648,N_23735);
nand U27051 (N_27051,N_24416,N_24520);
or U27052 (N_27052,N_21758,N_24696);
or U27053 (N_27053,N_24266,N_21345);
and U27054 (N_27054,N_21834,N_20091);
xor U27055 (N_27055,N_22619,N_24191);
nor U27056 (N_27056,N_23687,N_22486);
nand U27057 (N_27057,N_20037,N_20371);
nand U27058 (N_27058,N_21732,N_23185);
and U27059 (N_27059,N_24264,N_24950);
or U27060 (N_27060,N_20478,N_22336);
and U27061 (N_27061,N_23220,N_23697);
or U27062 (N_27062,N_21388,N_22462);
nand U27063 (N_27063,N_22432,N_22288);
or U27064 (N_27064,N_24210,N_22192);
or U27065 (N_27065,N_24275,N_23264);
nor U27066 (N_27066,N_20125,N_21647);
or U27067 (N_27067,N_24976,N_24065);
or U27068 (N_27068,N_22028,N_24281);
nor U27069 (N_27069,N_24507,N_23235);
and U27070 (N_27070,N_24424,N_21289);
and U27071 (N_27071,N_23581,N_23437);
nor U27072 (N_27072,N_21094,N_24524);
and U27073 (N_27073,N_22117,N_24272);
nand U27074 (N_27074,N_21823,N_21789);
xnor U27075 (N_27075,N_23601,N_22776);
nor U27076 (N_27076,N_21395,N_21728);
nand U27077 (N_27077,N_22315,N_21468);
and U27078 (N_27078,N_21270,N_22145);
nor U27079 (N_27079,N_24147,N_21989);
nand U27080 (N_27080,N_21931,N_23064);
or U27081 (N_27081,N_22828,N_20608);
xor U27082 (N_27082,N_21879,N_23505);
or U27083 (N_27083,N_24729,N_23908);
or U27084 (N_27084,N_20595,N_22259);
nor U27085 (N_27085,N_22680,N_23640);
and U27086 (N_27086,N_22314,N_24487);
nand U27087 (N_27087,N_23691,N_24301);
xnor U27088 (N_27088,N_21281,N_24946);
nor U27089 (N_27089,N_21776,N_24248);
nand U27090 (N_27090,N_23199,N_21442);
nand U27091 (N_27091,N_23738,N_23560);
nand U27092 (N_27092,N_23878,N_21404);
or U27093 (N_27093,N_20975,N_22797);
nand U27094 (N_27094,N_21612,N_21945);
or U27095 (N_27095,N_24269,N_20246);
and U27096 (N_27096,N_20787,N_20305);
or U27097 (N_27097,N_23647,N_24565);
and U27098 (N_27098,N_24742,N_20558);
xnor U27099 (N_27099,N_23339,N_24423);
xnor U27100 (N_27100,N_23634,N_23303);
xnor U27101 (N_27101,N_24351,N_20987);
nor U27102 (N_27102,N_22747,N_21562);
and U27103 (N_27103,N_24712,N_21936);
and U27104 (N_27104,N_24568,N_20204);
and U27105 (N_27105,N_23270,N_21485);
nor U27106 (N_27106,N_24192,N_23838);
nand U27107 (N_27107,N_23050,N_23077);
and U27108 (N_27108,N_22515,N_20590);
or U27109 (N_27109,N_20202,N_20914);
and U27110 (N_27110,N_21542,N_24935);
and U27111 (N_27111,N_22787,N_23608);
xor U27112 (N_27112,N_23651,N_20259);
nor U27113 (N_27113,N_23137,N_20128);
or U27114 (N_27114,N_22764,N_21735);
nand U27115 (N_27115,N_20375,N_23032);
or U27116 (N_27116,N_23460,N_22308);
nor U27117 (N_27117,N_24260,N_23771);
nand U27118 (N_27118,N_24162,N_22453);
nor U27119 (N_27119,N_23937,N_20826);
xor U27120 (N_27120,N_21066,N_23590);
nand U27121 (N_27121,N_21203,N_24553);
and U27122 (N_27122,N_21830,N_21716);
and U27123 (N_27123,N_20137,N_22211);
nand U27124 (N_27124,N_21333,N_24736);
nand U27125 (N_27125,N_22293,N_20845);
nand U27126 (N_27126,N_23259,N_20546);
and U27127 (N_27127,N_22978,N_24482);
or U27128 (N_27128,N_24924,N_20138);
and U27129 (N_27129,N_24570,N_23222);
or U27130 (N_27130,N_23288,N_24257);
or U27131 (N_27131,N_22581,N_23216);
xnor U27132 (N_27132,N_24701,N_22610);
or U27133 (N_27133,N_23924,N_20777);
xor U27134 (N_27134,N_21240,N_24082);
and U27135 (N_27135,N_24698,N_23271);
nor U27136 (N_27136,N_21826,N_22882);
or U27137 (N_27137,N_22205,N_20374);
nand U27138 (N_27138,N_23692,N_21787);
or U27139 (N_27139,N_20345,N_24323);
or U27140 (N_27140,N_24583,N_20689);
nand U27141 (N_27141,N_24335,N_20332);
or U27142 (N_27142,N_22849,N_20310);
or U27143 (N_27143,N_22510,N_23892);
nor U27144 (N_27144,N_23356,N_24417);
or U27145 (N_27145,N_24811,N_20350);
nor U27146 (N_27146,N_20226,N_24737);
xnor U27147 (N_27147,N_23616,N_24649);
and U27148 (N_27148,N_22508,N_23160);
nand U27149 (N_27149,N_20700,N_21534);
or U27150 (N_27150,N_22101,N_24752);
and U27151 (N_27151,N_20319,N_23621);
and U27152 (N_27152,N_24118,N_20544);
nor U27153 (N_27153,N_21531,N_23395);
nand U27154 (N_27154,N_22953,N_22447);
xor U27155 (N_27155,N_20600,N_23890);
and U27156 (N_27156,N_24431,N_24489);
nand U27157 (N_27157,N_21992,N_21363);
nor U27158 (N_27158,N_24930,N_21425);
xnor U27159 (N_27159,N_20381,N_21361);
xor U27160 (N_27160,N_24744,N_24421);
nand U27161 (N_27161,N_21037,N_22477);
nor U27162 (N_27162,N_22942,N_21158);
nor U27163 (N_27163,N_20754,N_24292);
nand U27164 (N_27164,N_24329,N_23744);
or U27165 (N_27165,N_20625,N_20411);
or U27166 (N_27166,N_20661,N_23410);
nand U27167 (N_27167,N_22074,N_20390);
or U27168 (N_27168,N_23732,N_22278);
nand U27169 (N_27169,N_23853,N_21962);
nand U27170 (N_27170,N_20548,N_20604);
nand U27171 (N_27171,N_23423,N_20489);
and U27172 (N_27172,N_21224,N_22672);
or U27173 (N_27173,N_24606,N_21756);
nand U27174 (N_27174,N_22748,N_20316);
nand U27175 (N_27175,N_21045,N_24276);
or U27176 (N_27176,N_23533,N_24095);
nor U27177 (N_27177,N_22536,N_22590);
nor U27178 (N_27178,N_21422,N_24460);
nor U27179 (N_27179,N_22401,N_20768);
xnor U27180 (N_27180,N_24982,N_22702);
and U27181 (N_27181,N_22005,N_21985);
or U27182 (N_27182,N_20433,N_21917);
and U27183 (N_27183,N_22381,N_21486);
and U27184 (N_27184,N_23795,N_20697);
nor U27185 (N_27185,N_20403,N_24669);
nor U27186 (N_27186,N_23706,N_22107);
nand U27187 (N_27187,N_22907,N_23377);
nand U27188 (N_27188,N_23263,N_22960);
and U27189 (N_27189,N_21730,N_21635);
nand U27190 (N_27190,N_20280,N_23524);
nor U27191 (N_27191,N_20340,N_20899);
or U27192 (N_27192,N_22875,N_21891);
xnor U27193 (N_27193,N_20367,N_21966);
nor U27194 (N_27194,N_20421,N_24939);
and U27195 (N_27195,N_21813,N_24558);
and U27196 (N_27196,N_22670,N_20676);
nand U27197 (N_27197,N_22472,N_24307);
nand U27198 (N_27198,N_22487,N_23591);
nor U27199 (N_27199,N_24648,N_23498);
nand U27200 (N_27200,N_22326,N_20644);
nor U27201 (N_27201,N_20582,N_20988);
nand U27202 (N_27202,N_20568,N_20038);
nand U27203 (N_27203,N_24663,N_24050);
nand U27204 (N_27204,N_20277,N_21285);
nor U27205 (N_27205,N_22795,N_21520);
and U27206 (N_27206,N_22368,N_21271);
or U27207 (N_27207,N_22644,N_23983);
and U27208 (N_27208,N_21798,N_24158);
nor U27209 (N_27209,N_20026,N_22746);
nand U27210 (N_27210,N_24014,N_24707);
or U27211 (N_27211,N_22130,N_21540);
nor U27212 (N_27212,N_23406,N_20888);
nand U27213 (N_27213,N_21495,N_24067);
nand U27214 (N_27214,N_23439,N_22222);
and U27215 (N_27215,N_23596,N_22042);
or U27216 (N_27216,N_21824,N_24684);
or U27217 (N_27217,N_20758,N_21692);
nand U27218 (N_27218,N_21699,N_22080);
xor U27219 (N_27219,N_23871,N_22662);
nand U27220 (N_27220,N_20973,N_21820);
or U27221 (N_27221,N_21370,N_24121);
nand U27222 (N_27222,N_21231,N_20097);
and U27223 (N_27223,N_20841,N_24738);
xnor U27224 (N_27224,N_21980,N_20092);
nand U27225 (N_27225,N_20361,N_24961);
nor U27226 (N_27226,N_24283,N_22530);
nand U27227 (N_27227,N_24880,N_24138);
or U27228 (N_27228,N_22111,N_20683);
or U27229 (N_27229,N_24170,N_22012);
nand U27230 (N_27230,N_20791,N_22277);
or U27231 (N_27231,N_24051,N_21764);
or U27232 (N_27232,N_23520,N_22498);
or U27233 (N_27233,N_21819,N_24772);
nand U27234 (N_27234,N_21092,N_24940);
or U27235 (N_27235,N_22807,N_23135);
nor U27236 (N_27236,N_20640,N_24501);
or U27237 (N_27237,N_22872,N_21033);
nand U27238 (N_27238,N_23430,N_20954);
xnor U27239 (N_27239,N_24036,N_24559);
and U27240 (N_27240,N_23784,N_22253);
xor U27241 (N_27241,N_20369,N_22886);
nand U27242 (N_27242,N_23182,N_20760);
or U27243 (N_27243,N_21876,N_23455);
and U27244 (N_27244,N_23541,N_22723);
nor U27245 (N_27245,N_24113,N_23914);
nand U27246 (N_27246,N_21571,N_24213);
and U27247 (N_27247,N_20326,N_24188);
nor U27248 (N_27248,N_22091,N_23282);
and U27249 (N_27249,N_22008,N_20656);
nand U27250 (N_27250,N_20068,N_21000);
or U27251 (N_27251,N_24115,N_20036);
nor U27252 (N_27252,N_24903,N_23886);
or U27253 (N_27253,N_24483,N_20464);
or U27254 (N_27254,N_21554,N_23345);
nand U27255 (N_27255,N_23854,N_23865);
or U27256 (N_27256,N_20627,N_22235);
and U27257 (N_27257,N_21816,N_22891);
nor U27258 (N_27258,N_20487,N_23707);
and U27259 (N_27259,N_23087,N_24694);
xor U27260 (N_27260,N_21709,N_24168);
nor U27261 (N_27261,N_23845,N_24117);
nor U27262 (N_27262,N_24622,N_22616);
and U27263 (N_27263,N_21201,N_24801);
or U27264 (N_27264,N_22056,N_24853);
and U27265 (N_27265,N_21133,N_23479);
and U27266 (N_27266,N_21851,N_21360);
nor U27267 (N_27267,N_24833,N_21839);
nor U27268 (N_27268,N_22560,N_23592);
and U27269 (N_27269,N_22359,N_21266);
nor U27270 (N_27270,N_24463,N_21137);
and U27271 (N_27271,N_23829,N_23544);
xnor U27272 (N_27272,N_24499,N_22665);
or U27273 (N_27273,N_21750,N_20481);
xor U27274 (N_27274,N_22783,N_24627);
nor U27275 (N_27275,N_22569,N_22236);
and U27276 (N_27276,N_23828,N_22661);
and U27277 (N_27277,N_21805,N_23660);
nor U27278 (N_27278,N_21193,N_24003);
and U27279 (N_27279,N_24415,N_24176);
or U27280 (N_27280,N_20822,N_24072);
or U27281 (N_27281,N_23466,N_22020);
and U27282 (N_27282,N_20967,N_21566);
nand U27283 (N_27283,N_23587,N_20816);
nor U27284 (N_27284,N_20427,N_23399);
nor U27285 (N_27285,N_22674,N_21768);
nand U27286 (N_27286,N_23161,N_24840);
nand U27287 (N_27287,N_21170,N_21800);
nand U27288 (N_27288,N_21139,N_21192);
nor U27289 (N_27289,N_21746,N_20181);
or U27290 (N_27290,N_23320,N_24461);
and U27291 (N_27291,N_22846,N_23627);
or U27292 (N_27292,N_23101,N_23090);
or U27293 (N_27293,N_23332,N_23490);
nand U27294 (N_27294,N_21431,N_24409);
nand U27295 (N_27295,N_22214,N_24120);
and U27296 (N_27296,N_20294,N_21132);
and U27297 (N_27297,N_21487,N_22633);
and U27298 (N_27298,N_23700,N_24902);
xor U27299 (N_27299,N_21996,N_20364);
or U27300 (N_27300,N_22858,N_23880);
or U27301 (N_27301,N_23726,N_21932);
or U27302 (N_27302,N_23842,N_22105);
nand U27303 (N_27303,N_23424,N_21557);
and U27304 (N_27304,N_20606,N_23002);
and U27305 (N_27305,N_20508,N_23613);
and U27306 (N_27306,N_21337,N_22434);
nor U27307 (N_27307,N_24644,N_24202);
xor U27308 (N_27308,N_23093,N_24059);
or U27309 (N_27309,N_21589,N_23668);
nand U27310 (N_27310,N_20103,N_21958);
nor U27311 (N_27311,N_21981,N_20521);
nand U27312 (N_27312,N_21584,N_23862);
or U27313 (N_27313,N_23247,N_21792);
nor U27314 (N_27314,N_23102,N_21703);
nor U27315 (N_27315,N_20819,N_24012);
or U27316 (N_27316,N_22814,N_23753);
or U27317 (N_27317,N_24349,N_24471);
nor U27318 (N_27318,N_24824,N_20842);
or U27319 (N_27319,N_21598,N_23864);
nor U27320 (N_27320,N_21618,N_20505);
and U27321 (N_27321,N_20120,N_21054);
and U27322 (N_27322,N_22671,N_24803);
and U27323 (N_27323,N_24604,N_24904);
nor U27324 (N_27324,N_24077,N_24971);
nor U27325 (N_27325,N_21995,N_21312);
nor U27326 (N_27326,N_24352,N_24519);
nand U27327 (N_27327,N_21100,N_21915);
nor U27328 (N_27328,N_20641,N_23797);
nand U27329 (N_27329,N_22585,N_22267);
xnor U27330 (N_27330,N_23614,N_22388);
and U27331 (N_27331,N_22664,N_20800);
nand U27332 (N_27332,N_22556,N_23206);
nor U27333 (N_27333,N_20864,N_22517);
and U27334 (N_27334,N_22344,N_24664);
nand U27335 (N_27335,N_22195,N_20658);
or U27336 (N_27336,N_20025,N_22119);
xnor U27337 (N_27337,N_21626,N_23825);
nor U27338 (N_27338,N_21471,N_22895);
and U27339 (N_27339,N_21451,N_21593);
and U27340 (N_27340,N_24660,N_21087);
nand U27341 (N_27341,N_20140,N_24638);
nand U27342 (N_27342,N_24582,N_24245);
nand U27343 (N_27343,N_22484,N_23008);
xnor U27344 (N_27344,N_21075,N_22609);
nor U27345 (N_27345,N_22840,N_22803);
and U27346 (N_27346,N_23366,N_20051);
and U27347 (N_27347,N_24944,N_23708);
nand U27348 (N_27348,N_20665,N_21659);
nand U27349 (N_27349,N_24643,N_23957);
and U27350 (N_27350,N_20765,N_21685);
xnor U27351 (N_27351,N_20672,N_22391);
nand U27352 (N_27352,N_24996,N_23227);
nor U27353 (N_27353,N_24927,N_23197);
and U27354 (N_27354,N_22292,N_23080);
nor U27355 (N_27355,N_24802,N_21341);
xnor U27356 (N_27356,N_22678,N_20662);
nor U27357 (N_27357,N_21235,N_23618);
xnor U27358 (N_27358,N_20425,N_20643);
nand U27359 (N_27359,N_24654,N_24771);
or U27360 (N_27360,N_23193,N_24584);
and U27361 (N_27361,N_22392,N_20866);
nand U27362 (N_27362,N_23968,N_20771);
nor U27363 (N_27363,N_21979,N_24867);
nand U27364 (N_27364,N_20821,N_20919);
nor U27365 (N_27365,N_21358,N_23696);
and U27366 (N_27366,N_23170,N_23342);
nand U27367 (N_27367,N_23578,N_24890);
and U27368 (N_27368,N_21182,N_22488);
and U27369 (N_27369,N_22789,N_20408);
nor U27370 (N_27370,N_24881,N_23563);
nand U27371 (N_27371,N_21632,N_22565);
nor U27372 (N_27372,N_22393,N_21308);
or U27373 (N_27373,N_20286,N_23598);
nand U27374 (N_27374,N_24653,N_22601);
or U27375 (N_27375,N_24804,N_23136);
nor U27376 (N_27376,N_23190,N_24199);
or U27377 (N_27377,N_22142,N_21505);
and U27378 (N_27378,N_23153,N_22229);
xnor U27379 (N_27379,N_21481,N_20848);
and U27380 (N_27380,N_23373,N_21305);
or U27381 (N_27381,N_23054,N_20030);
or U27382 (N_27382,N_20342,N_21696);
or U27383 (N_27383,N_21382,N_24181);
nand U27384 (N_27384,N_20245,N_20862);
or U27385 (N_27385,N_21141,N_24762);
and U27386 (N_27386,N_23655,N_23677);
nand U27387 (N_27387,N_24699,N_21579);
nor U27388 (N_27388,N_21477,N_22518);
and U27389 (N_27389,N_23202,N_21925);
or U27390 (N_27390,N_23637,N_23913);
nor U27391 (N_27391,N_20634,N_20059);
or U27392 (N_27392,N_20911,N_24732);
nand U27393 (N_27393,N_23536,N_24467);
nand U27394 (N_27394,N_23114,N_21402);
nand U27395 (N_27395,N_21230,N_20724);
and U27396 (N_27396,N_21508,N_23985);
and U27397 (N_27397,N_23922,N_23192);
nand U27398 (N_27398,N_22440,N_22057);
nor U27399 (N_27399,N_23493,N_24884);
nor U27400 (N_27400,N_22526,N_21198);
nor U27401 (N_27401,N_20486,N_20053);
and U27402 (N_27402,N_20384,N_24917);
and U27403 (N_27403,N_20145,N_24156);
nand U27404 (N_27404,N_22050,N_23151);
or U27405 (N_27405,N_21238,N_21043);
or U27406 (N_27406,N_23030,N_24585);
nand U27407 (N_27407,N_24714,N_22901);
or U27408 (N_27408,N_24988,N_23648);
nand U27409 (N_27409,N_20564,N_24725);
and U27410 (N_27410,N_21336,N_23252);
nand U27411 (N_27411,N_22798,N_23670);
nor U27412 (N_27412,N_24132,N_22712);
and U27413 (N_27413,N_22332,N_20392);
nand U27414 (N_27414,N_20451,N_24054);
or U27415 (N_27415,N_23727,N_21957);
and U27416 (N_27416,N_24715,N_21918);
nand U27417 (N_27417,N_23381,N_24369);
or U27418 (N_27418,N_24428,N_21446);
nand U27419 (N_27419,N_20216,N_23359);
nor U27420 (N_27420,N_22813,N_23658);
nor U27421 (N_27421,N_21147,N_20349);
nor U27422 (N_27422,N_20763,N_21613);
nor U27423 (N_27423,N_21640,N_24343);
xor U27424 (N_27424,N_24652,N_22574);
nor U27425 (N_27425,N_22476,N_20944);
or U27426 (N_27426,N_21377,N_24888);
and U27427 (N_27427,N_21241,N_23569);
nand U27428 (N_27428,N_24518,N_21131);
nand U27429 (N_27429,N_23764,N_20276);
or U27430 (N_27430,N_24303,N_24015);
nand U27431 (N_27431,N_20601,N_24502);
nand U27432 (N_27432,N_22709,N_21828);
and U27433 (N_27433,N_21867,N_21869);
nor U27434 (N_27434,N_21362,N_21232);
nand U27435 (N_27435,N_20094,N_22306);
xor U27436 (N_27436,N_22069,N_21543);
nor U27437 (N_27437,N_21472,N_24778);
nand U27438 (N_27438,N_20514,N_24765);
nand U27439 (N_27439,N_20039,N_22966);
and U27440 (N_27440,N_24956,N_22754);
and U27441 (N_27441,N_22580,N_20996);
or U27442 (N_27442,N_24179,N_22659);
nor U27443 (N_27443,N_20028,N_20228);
or U27444 (N_27444,N_23562,N_20236);
nor U27445 (N_27445,N_24316,N_24923);
nor U27446 (N_27446,N_24726,N_23650);
xnor U27447 (N_27447,N_20383,N_20344);
nor U27448 (N_27448,N_24338,N_21369);
or U27449 (N_27449,N_23462,N_23518);
and U27450 (N_27450,N_20446,N_23526);
nand U27451 (N_27451,N_20649,N_24092);
xor U27452 (N_27452,N_22596,N_21118);
or U27453 (N_27453,N_23134,N_24514);
nand U27454 (N_27454,N_21429,N_24375);
or U27455 (N_27455,N_20980,N_23630);
nor U27456 (N_27456,N_24261,N_22096);
or U27457 (N_27457,N_20416,N_23931);
or U27458 (N_27458,N_24278,N_20452);
and U27459 (N_27459,N_24848,N_20571);
nand U27460 (N_27460,N_21390,N_20347);
or U27461 (N_27461,N_24094,N_24625);
nor U27462 (N_27462,N_21814,N_22699);
and U27463 (N_27463,N_24723,N_23118);
and U27464 (N_27464,N_21939,N_24929);
nor U27465 (N_27465,N_24379,N_22431);
nor U27466 (N_27466,N_20766,N_24510);
or U27467 (N_27467,N_21269,N_24894);
nor U27468 (N_27468,N_22784,N_22504);
xnor U27469 (N_27469,N_20417,N_24173);
nor U27470 (N_27470,N_23515,N_20404);
nor U27471 (N_27471,N_21914,N_24244);
nand U27472 (N_27472,N_22869,N_20082);
nor U27473 (N_27473,N_21748,N_21430);
nor U27474 (N_27474,N_24531,N_21142);
or U27475 (N_27475,N_22630,N_24422);
nor U27476 (N_27476,N_24624,N_21150);
and U27477 (N_27477,N_21953,N_20678);
and U27478 (N_27478,N_24466,N_24914);
and U27479 (N_27479,N_23172,N_21465);
nor U27480 (N_27480,N_22033,N_21457);
nor U27481 (N_27481,N_21665,N_20479);
or U27482 (N_27482,N_22349,N_22352);
nor U27483 (N_27483,N_24447,N_20515);
nor U27484 (N_27484,N_24413,N_22981);
or U27485 (N_27485,N_22597,N_20477);
xor U27486 (N_27486,N_21715,N_23675);
nor U27487 (N_27487,N_22939,N_23427);
and U27488 (N_27488,N_22588,N_22894);
and U27489 (N_27489,N_20893,N_22113);
nor U27490 (N_27490,N_20580,N_23021);
nand U27491 (N_27491,N_23337,N_23993);
nor U27492 (N_27492,N_23082,N_21707);
and U27493 (N_27493,N_21398,N_22337);
nand U27494 (N_27494,N_20469,N_22499);
or U27495 (N_27495,N_22457,N_24680);
and U27496 (N_27496,N_23705,N_22072);
or U27497 (N_27497,N_20267,N_20999);
nor U27498 (N_27498,N_20233,N_22839);
nand U27499 (N_27499,N_24205,N_24700);
nor U27500 (N_27500,N_22930,N_22079);
and U27501 (N_27501,N_24620,N_24049);
and U27502 (N_27502,N_24428,N_23375);
nand U27503 (N_27503,N_24097,N_23799);
or U27504 (N_27504,N_23662,N_24687);
nand U27505 (N_27505,N_23616,N_20480);
and U27506 (N_27506,N_24627,N_24854);
and U27507 (N_27507,N_20904,N_23981);
nand U27508 (N_27508,N_20497,N_24939);
or U27509 (N_27509,N_22436,N_23358);
nand U27510 (N_27510,N_21526,N_21269);
or U27511 (N_27511,N_21690,N_24400);
xor U27512 (N_27512,N_22653,N_23456);
and U27513 (N_27513,N_21008,N_24199);
and U27514 (N_27514,N_20606,N_24488);
and U27515 (N_27515,N_21214,N_23635);
xnor U27516 (N_27516,N_22926,N_24095);
nand U27517 (N_27517,N_23877,N_20606);
nor U27518 (N_27518,N_23669,N_21372);
nor U27519 (N_27519,N_20817,N_23868);
nand U27520 (N_27520,N_21107,N_23912);
nor U27521 (N_27521,N_23510,N_20004);
nand U27522 (N_27522,N_22534,N_20044);
or U27523 (N_27523,N_21893,N_20428);
nand U27524 (N_27524,N_21244,N_21216);
nand U27525 (N_27525,N_20910,N_23311);
and U27526 (N_27526,N_20489,N_20047);
or U27527 (N_27527,N_22021,N_22198);
nand U27528 (N_27528,N_20942,N_24742);
nor U27529 (N_27529,N_20587,N_23741);
or U27530 (N_27530,N_20753,N_21362);
nor U27531 (N_27531,N_20160,N_24062);
and U27532 (N_27532,N_20199,N_23102);
nand U27533 (N_27533,N_21230,N_21446);
and U27534 (N_27534,N_23407,N_20331);
nor U27535 (N_27535,N_20103,N_22729);
or U27536 (N_27536,N_21180,N_21241);
nor U27537 (N_27537,N_21602,N_20016);
nand U27538 (N_27538,N_20750,N_20775);
nor U27539 (N_27539,N_24252,N_24307);
nor U27540 (N_27540,N_20970,N_21109);
nand U27541 (N_27541,N_22608,N_21616);
and U27542 (N_27542,N_21690,N_21078);
nand U27543 (N_27543,N_24302,N_21800);
nor U27544 (N_27544,N_20580,N_24873);
nand U27545 (N_27545,N_24683,N_23874);
xnor U27546 (N_27546,N_23403,N_20531);
or U27547 (N_27547,N_21820,N_23441);
nor U27548 (N_27548,N_20651,N_22441);
nand U27549 (N_27549,N_20688,N_23310);
or U27550 (N_27550,N_21697,N_22074);
nand U27551 (N_27551,N_20858,N_21337);
nand U27552 (N_27552,N_24378,N_22687);
and U27553 (N_27553,N_22230,N_24139);
and U27554 (N_27554,N_23448,N_23236);
nand U27555 (N_27555,N_24010,N_22404);
xnor U27556 (N_27556,N_22278,N_23826);
nor U27557 (N_27557,N_22249,N_23284);
or U27558 (N_27558,N_20654,N_23008);
or U27559 (N_27559,N_24489,N_24145);
nand U27560 (N_27560,N_24632,N_22883);
nor U27561 (N_27561,N_24663,N_22421);
nor U27562 (N_27562,N_22633,N_21563);
nand U27563 (N_27563,N_22272,N_20498);
nand U27564 (N_27564,N_24471,N_21103);
and U27565 (N_27565,N_21900,N_21302);
nand U27566 (N_27566,N_24575,N_21835);
nand U27567 (N_27567,N_21771,N_20067);
nor U27568 (N_27568,N_23224,N_20311);
nand U27569 (N_27569,N_24367,N_21458);
and U27570 (N_27570,N_22625,N_21335);
nand U27571 (N_27571,N_22069,N_21628);
and U27572 (N_27572,N_20402,N_23262);
nand U27573 (N_27573,N_22190,N_23027);
nand U27574 (N_27574,N_21791,N_24943);
and U27575 (N_27575,N_21370,N_21896);
and U27576 (N_27576,N_21963,N_21570);
or U27577 (N_27577,N_21545,N_20838);
xnor U27578 (N_27578,N_23359,N_23324);
or U27579 (N_27579,N_22775,N_23596);
nor U27580 (N_27580,N_24180,N_24253);
or U27581 (N_27581,N_20662,N_21045);
or U27582 (N_27582,N_21786,N_21725);
or U27583 (N_27583,N_24442,N_21401);
and U27584 (N_27584,N_20610,N_21423);
nand U27585 (N_27585,N_21137,N_24836);
nor U27586 (N_27586,N_24866,N_24501);
nor U27587 (N_27587,N_20107,N_20368);
nor U27588 (N_27588,N_20345,N_23507);
nor U27589 (N_27589,N_23171,N_23739);
nor U27590 (N_27590,N_21220,N_24919);
and U27591 (N_27591,N_23199,N_24995);
xnor U27592 (N_27592,N_23901,N_21091);
and U27593 (N_27593,N_24146,N_21654);
nand U27594 (N_27594,N_22644,N_20728);
nand U27595 (N_27595,N_23725,N_23904);
nand U27596 (N_27596,N_24429,N_21595);
and U27597 (N_27597,N_23709,N_20042);
or U27598 (N_27598,N_21055,N_23067);
nor U27599 (N_27599,N_23925,N_20188);
and U27600 (N_27600,N_22742,N_22695);
nor U27601 (N_27601,N_21743,N_22655);
or U27602 (N_27602,N_20229,N_23428);
nor U27603 (N_27603,N_23215,N_24726);
and U27604 (N_27604,N_21529,N_24042);
or U27605 (N_27605,N_21069,N_22922);
and U27606 (N_27606,N_21937,N_22240);
nor U27607 (N_27607,N_22701,N_23348);
and U27608 (N_27608,N_21526,N_20200);
nor U27609 (N_27609,N_22783,N_22501);
or U27610 (N_27610,N_20258,N_20850);
nand U27611 (N_27611,N_22363,N_21347);
and U27612 (N_27612,N_20814,N_21014);
nand U27613 (N_27613,N_21136,N_21235);
nand U27614 (N_27614,N_22819,N_21661);
nand U27615 (N_27615,N_23554,N_20600);
nor U27616 (N_27616,N_22495,N_20850);
nand U27617 (N_27617,N_22482,N_20583);
nand U27618 (N_27618,N_21486,N_20190);
nand U27619 (N_27619,N_22107,N_24983);
xnor U27620 (N_27620,N_22827,N_21662);
and U27621 (N_27621,N_23669,N_22068);
or U27622 (N_27622,N_23245,N_20575);
nand U27623 (N_27623,N_23924,N_21459);
nand U27624 (N_27624,N_21544,N_21395);
nor U27625 (N_27625,N_21614,N_24141);
or U27626 (N_27626,N_22697,N_23169);
or U27627 (N_27627,N_24753,N_24132);
nand U27628 (N_27628,N_24830,N_23290);
or U27629 (N_27629,N_22787,N_23814);
and U27630 (N_27630,N_21511,N_23987);
and U27631 (N_27631,N_20804,N_20429);
xnor U27632 (N_27632,N_23975,N_24538);
and U27633 (N_27633,N_22124,N_24936);
or U27634 (N_27634,N_22067,N_20516);
and U27635 (N_27635,N_23963,N_24693);
and U27636 (N_27636,N_20797,N_23611);
nor U27637 (N_27637,N_22577,N_22525);
nor U27638 (N_27638,N_20408,N_24687);
and U27639 (N_27639,N_21234,N_24675);
and U27640 (N_27640,N_21310,N_21362);
nor U27641 (N_27641,N_21430,N_24568);
xor U27642 (N_27642,N_21209,N_24915);
xor U27643 (N_27643,N_22623,N_24779);
or U27644 (N_27644,N_21831,N_21984);
nor U27645 (N_27645,N_20388,N_24830);
nand U27646 (N_27646,N_20052,N_24299);
nand U27647 (N_27647,N_24979,N_24322);
or U27648 (N_27648,N_24992,N_20797);
nor U27649 (N_27649,N_22213,N_21539);
nor U27650 (N_27650,N_22892,N_23065);
and U27651 (N_27651,N_24650,N_21658);
and U27652 (N_27652,N_21226,N_23947);
nand U27653 (N_27653,N_20915,N_23131);
or U27654 (N_27654,N_22719,N_20763);
xnor U27655 (N_27655,N_22308,N_21568);
or U27656 (N_27656,N_23306,N_23983);
and U27657 (N_27657,N_22661,N_24851);
or U27658 (N_27658,N_23759,N_24373);
or U27659 (N_27659,N_21826,N_24927);
and U27660 (N_27660,N_23284,N_24431);
nor U27661 (N_27661,N_24164,N_20909);
or U27662 (N_27662,N_22234,N_20404);
xnor U27663 (N_27663,N_23679,N_24056);
nor U27664 (N_27664,N_22560,N_22015);
nand U27665 (N_27665,N_22590,N_23116);
nand U27666 (N_27666,N_20342,N_23090);
and U27667 (N_27667,N_21745,N_23167);
nor U27668 (N_27668,N_24579,N_22876);
or U27669 (N_27669,N_23641,N_22468);
or U27670 (N_27670,N_22894,N_23070);
nor U27671 (N_27671,N_23181,N_22680);
nand U27672 (N_27672,N_21975,N_24163);
nand U27673 (N_27673,N_22558,N_24942);
xor U27674 (N_27674,N_22785,N_23685);
and U27675 (N_27675,N_20217,N_23105);
and U27676 (N_27676,N_24327,N_24338);
or U27677 (N_27677,N_22382,N_23028);
or U27678 (N_27678,N_22182,N_24673);
or U27679 (N_27679,N_22636,N_24747);
nand U27680 (N_27680,N_22283,N_22092);
xor U27681 (N_27681,N_22117,N_22453);
xor U27682 (N_27682,N_24052,N_23977);
nand U27683 (N_27683,N_24918,N_22597);
nand U27684 (N_27684,N_20299,N_23029);
nand U27685 (N_27685,N_22393,N_21016);
nor U27686 (N_27686,N_23650,N_20486);
or U27687 (N_27687,N_21729,N_23717);
nand U27688 (N_27688,N_20985,N_23693);
and U27689 (N_27689,N_24545,N_20813);
nand U27690 (N_27690,N_20185,N_23378);
nor U27691 (N_27691,N_20280,N_21135);
xor U27692 (N_27692,N_22122,N_21825);
xor U27693 (N_27693,N_22689,N_22575);
nand U27694 (N_27694,N_20852,N_21160);
or U27695 (N_27695,N_22671,N_23421);
or U27696 (N_27696,N_21909,N_22791);
nor U27697 (N_27697,N_24542,N_21894);
nor U27698 (N_27698,N_20712,N_21201);
nand U27699 (N_27699,N_20358,N_24057);
nand U27700 (N_27700,N_24035,N_22891);
nand U27701 (N_27701,N_21493,N_21258);
or U27702 (N_27702,N_21912,N_21506);
xnor U27703 (N_27703,N_23460,N_20639);
or U27704 (N_27704,N_20136,N_24134);
nand U27705 (N_27705,N_24347,N_23107);
and U27706 (N_27706,N_23237,N_20702);
or U27707 (N_27707,N_21224,N_22018);
nor U27708 (N_27708,N_23546,N_21701);
and U27709 (N_27709,N_22249,N_22769);
or U27710 (N_27710,N_21455,N_22974);
nand U27711 (N_27711,N_24030,N_21896);
and U27712 (N_27712,N_21260,N_20780);
or U27713 (N_27713,N_23898,N_24212);
nor U27714 (N_27714,N_24539,N_23281);
nor U27715 (N_27715,N_24245,N_23105);
xor U27716 (N_27716,N_21207,N_21288);
and U27717 (N_27717,N_20348,N_21512);
and U27718 (N_27718,N_22956,N_24544);
nand U27719 (N_27719,N_20709,N_21237);
xor U27720 (N_27720,N_20647,N_24421);
nand U27721 (N_27721,N_20382,N_23132);
nand U27722 (N_27722,N_24798,N_22933);
nor U27723 (N_27723,N_20387,N_23804);
and U27724 (N_27724,N_20503,N_20386);
and U27725 (N_27725,N_22541,N_24164);
nor U27726 (N_27726,N_22771,N_24925);
nand U27727 (N_27727,N_20087,N_22648);
and U27728 (N_27728,N_24326,N_21706);
or U27729 (N_27729,N_20519,N_24746);
xnor U27730 (N_27730,N_20307,N_24195);
and U27731 (N_27731,N_24964,N_22651);
or U27732 (N_27732,N_20751,N_22655);
and U27733 (N_27733,N_22775,N_24927);
nor U27734 (N_27734,N_20719,N_23999);
nand U27735 (N_27735,N_20888,N_20528);
nand U27736 (N_27736,N_22172,N_20585);
nor U27737 (N_27737,N_21460,N_24921);
nand U27738 (N_27738,N_23810,N_21744);
and U27739 (N_27739,N_20583,N_24539);
or U27740 (N_27740,N_24905,N_22876);
nor U27741 (N_27741,N_20222,N_20792);
nand U27742 (N_27742,N_21799,N_20632);
nand U27743 (N_27743,N_20661,N_24724);
and U27744 (N_27744,N_22196,N_20886);
nand U27745 (N_27745,N_20929,N_22564);
nand U27746 (N_27746,N_24182,N_22758);
or U27747 (N_27747,N_20464,N_24126);
or U27748 (N_27748,N_23376,N_20904);
and U27749 (N_27749,N_20912,N_20134);
or U27750 (N_27750,N_20253,N_23095);
nor U27751 (N_27751,N_22029,N_20787);
and U27752 (N_27752,N_24675,N_22969);
or U27753 (N_27753,N_21667,N_21351);
and U27754 (N_27754,N_21944,N_23599);
nand U27755 (N_27755,N_21430,N_23311);
nor U27756 (N_27756,N_24068,N_22073);
and U27757 (N_27757,N_22392,N_24008);
or U27758 (N_27758,N_20342,N_22899);
or U27759 (N_27759,N_21278,N_24296);
or U27760 (N_27760,N_21840,N_22757);
or U27761 (N_27761,N_20096,N_24789);
nand U27762 (N_27762,N_20245,N_21124);
nand U27763 (N_27763,N_23899,N_24998);
nand U27764 (N_27764,N_21012,N_22287);
nor U27765 (N_27765,N_22801,N_21939);
nand U27766 (N_27766,N_20993,N_24576);
nand U27767 (N_27767,N_20555,N_24608);
xor U27768 (N_27768,N_20731,N_21650);
and U27769 (N_27769,N_20648,N_23714);
xnor U27770 (N_27770,N_22209,N_23593);
nor U27771 (N_27771,N_24502,N_21217);
xor U27772 (N_27772,N_22426,N_20860);
and U27773 (N_27773,N_24074,N_21364);
nand U27774 (N_27774,N_20422,N_23638);
nand U27775 (N_27775,N_24067,N_22676);
or U27776 (N_27776,N_24771,N_22712);
nand U27777 (N_27777,N_20177,N_20543);
nor U27778 (N_27778,N_20923,N_20832);
or U27779 (N_27779,N_20271,N_22944);
nor U27780 (N_27780,N_22583,N_24257);
nand U27781 (N_27781,N_24204,N_23218);
xor U27782 (N_27782,N_23817,N_21027);
or U27783 (N_27783,N_21174,N_24937);
nand U27784 (N_27784,N_24685,N_20274);
nor U27785 (N_27785,N_23421,N_24556);
or U27786 (N_27786,N_22438,N_22411);
or U27787 (N_27787,N_20687,N_21337);
xnor U27788 (N_27788,N_21342,N_20589);
and U27789 (N_27789,N_22905,N_22920);
and U27790 (N_27790,N_24842,N_21030);
xnor U27791 (N_27791,N_21073,N_21067);
or U27792 (N_27792,N_23531,N_23059);
and U27793 (N_27793,N_20715,N_23909);
or U27794 (N_27794,N_23432,N_22946);
and U27795 (N_27795,N_24214,N_23134);
and U27796 (N_27796,N_22651,N_23327);
nand U27797 (N_27797,N_20252,N_20289);
or U27798 (N_27798,N_23818,N_20837);
nand U27799 (N_27799,N_21624,N_23894);
and U27800 (N_27800,N_21660,N_20978);
xnor U27801 (N_27801,N_20097,N_22876);
or U27802 (N_27802,N_24256,N_23483);
or U27803 (N_27803,N_22814,N_20197);
xnor U27804 (N_27804,N_20389,N_24542);
nand U27805 (N_27805,N_23195,N_22557);
nor U27806 (N_27806,N_22343,N_21331);
and U27807 (N_27807,N_22576,N_24543);
and U27808 (N_27808,N_23425,N_21613);
nand U27809 (N_27809,N_22801,N_20277);
nand U27810 (N_27810,N_20437,N_24238);
nor U27811 (N_27811,N_20940,N_21009);
nor U27812 (N_27812,N_21842,N_21253);
or U27813 (N_27813,N_22732,N_23521);
nand U27814 (N_27814,N_21236,N_20250);
or U27815 (N_27815,N_20834,N_22985);
and U27816 (N_27816,N_23324,N_20758);
or U27817 (N_27817,N_21211,N_24995);
nand U27818 (N_27818,N_22023,N_21961);
nand U27819 (N_27819,N_21497,N_24984);
nand U27820 (N_27820,N_21430,N_22325);
nand U27821 (N_27821,N_24974,N_21098);
and U27822 (N_27822,N_22921,N_22979);
nor U27823 (N_27823,N_21253,N_20935);
nor U27824 (N_27824,N_23422,N_21487);
nand U27825 (N_27825,N_23829,N_24615);
and U27826 (N_27826,N_21119,N_20327);
and U27827 (N_27827,N_20094,N_20615);
nand U27828 (N_27828,N_24379,N_20061);
xnor U27829 (N_27829,N_23478,N_21679);
xor U27830 (N_27830,N_20023,N_23829);
or U27831 (N_27831,N_24169,N_20980);
nand U27832 (N_27832,N_24806,N_20885);
nor U27833 (N_27833,N_22728,N_20325);
nor U27834 (N_27834,N_22008,N_23755);
and U27835 (N_27835,N_22995,N_24540);
nor U27836 (N_27836,N_20384,N_23092);
or U27837 (N_27837,N_21189,N_22557);
nand U27838 (N_27838,N_24860,N_24838);
xor U27839 (N_27839,N_20871,N_21481);
nor U27840 (N_27840,N_21728,N_24124);
and U27841 (N_27841,N_24669,N_21781);
or U27842 (N_27842,N_24008,N_20477);
nand U27843 (N_27843,N_24177,N_22326);
xor U27844 (N_27844,N_24893,N_22553);
and U27845 (N_27845,N_20232,N_20765);
and U27846 (N_27846,N_22160,N_20556);
nand U27847 (N_27847,N_23923,N_22915);
or U27848 (N_27848,N_21401,N_21332);
nor U27849 (N_27849,N_20755,N_21124);
nor U27850 (N_27850,N_23556,N_23675);
nand U27851 (N_27851,N_20139,N_21367);
nand U27852 (N_27852,N_23338,N_21172);
and U27853 (N_27853,N_23587,N_20331);
nor U27854 (N_27854,N_24455,N_22940);
nand U27855 (N_27855,N_22379,N_24936);
nand U27856 (N_27856,N_21541,N_21655);
or U27857 (N_27857,N_22027,N_21333);
nor U27858 (N_27858,N_20985,N_24697);
and U27859 (N_27859,N_20370,N_20588);
or U27860 (N_27860,N_22741,N_23718);
xor U27861 (N_27861,N_22129,N_24639);
xor U27862 (N_27862,N_21300,N_23261);
and U27863 (N_27863,N_23410,N_20063);
and U27864 (N_27864,N_22386,N_23706);
nor U27865 (N_27865,N_24667,N_20410);
nor U27866 (N_27866,N_21050,N_20764);
xor U27867 (N_27867,N_20550,N_22074);
nor U27868 (N_27868,N_20021,N_23278);
or U27869 (N_27869,N_20860,N_24418);
nand U27870 (N_27870,N_22366,N_24961);
xnor U27871 (N_27871,N_22840,N_20050);
nand U27872 (N_27872,N_24595,N_20041);
nand U27873 (N_27873,N_22737,N_22055);
nand U27874 (N_27874,N_23947,N_24384);
nand U27875 (N_27875,N_23456,N_20524);
xor U27876 (N_27876,N_22147,N_21511);
and U27877 (N_27877,N_24536,N_21498);
or U27878 (N_27878,N_22410,N_21691);
nor U27879 (N_27879,N_22771,N_22044);
or U27880 (N_27880,N_23421,N_22527);
or U27881 (N_27881,N_20979,N_21721);
or U27882 (N_27882,N_23337,N_21220);
xnor U27883 (N_27883,N_21179,N_20414);
nor U27884 (N_27884,N_23705,N_24467);
nor U27885 (N_27885,N_20790,N_21035);
or U27886 (N_27886,N_20195,N_20382);
nor U27887 (N_27887,N_21829,N_23674);
xnor U27888 (N_27888,N_24108,N_22214);
or U27889 (N_27889,N_22091,N_20757);
and U27890 (N_27890,N_22449,N_23021);
and U27891 (N_27891,N_23973,N_21017);
nand U27892 (N_27892,N_24647,N_21190);
or U27893 (N_27893,N_24532,N_21670);
nor U27894 (N_27894,N_23532,N_24779);
nand U27895 (N_27895,N_22204,N_23430);
nor U27896 (N_27896,N_24393,N_23305);
and U27897 (N_27897,N_22222,N_21822);
and U27898 (N_27898,N_23414,N_23236);
nor U27899 (N_27899,N_21296,N_22753);
nand U27900 (N_27900,N_24838,N_22634);
or U27901 (N_27901,N_21355,N_22401);
or U27902 (N_27902,N_23044,N_22225);
nand U27903 (N_27903,N_22938,N_20335);
and U27904 (N_27904,N_20820,N_22059);
or U27905 (N_27905,N_23409,N_24551);
nand U27906 (N_27906,N_23009,N_23145);
and U27907 (N_27907,N_24907,N_24040);
nor U27908 (N_27908,N_23962,N_20828);
nand U27909 (N_27909,N_20673,N_21959);
nand U27910 (N_27910,N_24153,N_22771);
or U27911 (N_27911,N_23213,N_24168);
and U27912 (N_27912,N_22657,N_22024);
or U27913 (N_27913,N_23961,N_21754);
or U27914 (N_27914,N_23057,N_21183);
and U27915 (N_27915,N_23359,N_22848);
or U27916 (N_27916,N_21802,N_23976);
nor U27917 (N_27917,N_20930,N_24182);
and U27918 (N_27918,N_20104,N_24866);
nand U27919 (N_27919,N_21793,N_24927);
nor U27920 (N_27920,N_24640,N_24230);
or U27921 (N_27921,N_20156,N_24292);
or U27922 (N_27922,N_23803,N_20339);
nand U27923 (N_27923,N_21685,N_24191);
or U27924 (N_27924,N_22620,N_21276);
and U27925 (N_27925,N_21755,N_23513);
nor U27926 (N_27926,N_22535,N_24677);
or U27927 (N_27927,N_23929,N_22510);
and U27928 (N_27928,N_24621,N_21457);
nor U27929 (N_27929,N_24314,N_23450);
nor U27930 (N_27930,N_23919,N_22304);
nor U27931 (N_27931,N_22269,N_23037);
and U27932 (N_27932,N_23532,N_20438);
nor U27933 (N_27933,N_24326,N_21674);
nor U27934 (N_27934,N_20704,N_21965);
or U27935 (N_27935,N_21985,N_22176);
nor U27936 (N_27936,N_23705,N_22234);
or U27937 (N_27937,N_20155,N_24686);
or U27938 (N_27938,N_23142,N_24320);
nor U27939 (N_27939,N_22657,N_20301);
and U27940 (N_27940,N_22018,N_23021);
or U27941 (N_27941,N_23800,N_20847);
and U27942 (N_27942,N_21539,N_22598);
nor U27943 (N_27943,N_21393,N_24760);
nand U27944 (N_27944,N_22114,N_20747);
nand U27945 (N_27945,N_22081,N_21439);
and U27946 (N_27946,N_20080,N_23596);
nand U27947 (N_27947,N_23796,N_23530);
nand U27948 (N_27948,N_21695,N_21346);
or U27949 (N_27949,N_23358,N_21230);
or U27950 (N_27950,N_24193,N_21260);
and U27951 (N_27951,N_21680,N_23043);
nor U27952 (N_27952,N_20208,N_21602);
and U27953 (N_27953,N_22041,N_23633);
nor U27954 (N_27954,N_24056,N_20068);
xnor U27955 (N_27955,N_22236,N_24702);
nand U27956 (N_27956,N_20804,N_20352);
nor U27957 (N_27957,N_24347,N_20475);
nand U27958 (N_27958,N_20949,N_24756);
nor U27959 (N_27959,N_22869,N_21129);
or U27960 (N_27960,N_23879,N_21890);
and U27961 (N_27961,N_23625,N_22347);
xnor U27962 (N_27962,N_22003,N_20712);
nand U27963 (N_27963,N_22836,N_22496);
xor U27964 (N_27964,N_24760,N_24748);
nand U27965 (N_27965,N_24174,N_21693);
nor U27966 (N_27966,N_23915,N_21296);
and U27967 (N_27967,N_21359,N_24850);
nand U27968 (N_27968,N_24107,N_24008);
and U27969 (N_27969,N_22841,N_23645);
xnor U27970 (N_27970,N_20531,N_20897);
and U27971 (N_27971,N_20960,N_23254);
nand U27972 (N_27972,N_20913,N_24806);
nand U27973 (N_27973,N_20627,N_24955);
nand U27974 (N_27974,N_22432,N_24377);
and U27975 (N_27975,N_24271,N_23177);
and U27976 (N_27976,N_22409,N_20599);
nand U27977 (N_27977,N_21176,N_21377);
and U27978 (N_27978,N_23261,N_20551);
and U27979 (N_27979,N_22538,N_20862);
and U27980 (N_27980,N_23719,N_21449);
or U27981 (N_27981,N_24553,N_23008);
and U27982 (N_27982,N_23526,N_20084);
and U27983 (N_27983,N_20111,N_22699);
nor U27984 (N_27984,N_23808,N_23252);
nor U27985 (N_27985,N_21353,N_22969);
or U27986 (N_27986,N_22442,N_21087);
nand U27987 (N_27987,N_24908,N_24583);
xor U27988 (N_27988,N_21361,N_20437);
nand U27989 (N_27989,N_23416,N_22920);
nand U27990 (N_27990,N_21695,N_24452);
nor U27991 (N_27991,N_21479,N_22182);
xnor U27992 (N_27992,N_23175,N_21607);
or U27993 (N_27993,N_22287,N_23765);
or U27994 (N_27994,N_22658,N_24253);
nand U27995 (N_27995,N_20247,N_21071);
nand U27996 (N_27996,N_23092,N_20248);
nand U27997 (N_27997,N_24291,N_24992);
nand U27998 (N_27998,N_21743,N_22469);
or U27999 (N_27999,N_24396,N_20276);
nand U28000 (N_28000,N_24092,N_21609);
or U28001 (N_28001,N_22643,N_23155);
nand U28002 (N_28002,N_23019,N_22675);
or U28003 (N_28003,N_20629,N_21044);
nand U28004 (N_28004,N_21929,N_20175);
and U28005 (N_28005,N_24022,N_20763);
nand U28006 (N_28006,N_24532,N_20259);
nand U28007 (N_28007,N_20736,N_22445);
nand U28008 (N_28008,N_20535,N_20016);
or U28009 (N_28009,N_21532,N_23617);
nor U28010 (N_28010,N_20557,N_22286);
and U28011 (N_28011,N_20582,N_24834);
nand U28012 (N_28012,N_24559,N_20869);
xor U28013 (N_28013,N_22837,N_20488);
and U28014 (N_28014,N_20032,N_21431);
xnor U28015 (N_28015,N_20244,N_20762);
or U28016 (N_28016,N_24307,N_21851);
and U28017 (N_28017,N_20945,N_23996);
nand U28018 (N_28018,N_20860,N_22996);
nor U28019 (N_28019,N_20754,N_23857);
or U28020 (N_28020,N_20485,N_24915);
nor U28021 (N_28021,N_21697,N_20365);
nor U28022 (N_28022,N_23064,N_22047);
and U28023 (N_28023,N_23284,N_21953);
nand U28024 (N_28024,N_20993,N_22842);
nor U28025 (N_28025,N_20623,N_21624);
or U28026 (N_28026,N_21254,N_23595);
or U28027 (N_28027,N_21554,N_21788);
or U28028 (N_28028,N_20204,N_24386);
nand U28029 (N_28029,N_24021,N_21019);
or U28030 (N_28030,N_22173,N_21164);
xor U28031 (N_28031,N_20709,N_24392);
or U28032 (N_28032,N_23293,N_23252);
and U28033 (N_28033,N_23772,N_21485);
and U28034 (N_28034,N_22859,N_24002);
nand U28035 (N_28035,N_21903,N_23973);
xnor U28036 (N_28036,N_22525,N_23504);
or U28037 (N_28037,N_23384,N_22494);
xnor U28038 (N_28038,N_24788,N_23917);
or U28039 (N_28039,N_23582,N_23852);
nand U28040 (N_28040,N_24647,N_22426);
or U28041 (N_28041,N_23456,N_22432);
nor U28042 (N_28042,N_20843,N_24225);
nor U28043 (N_28043,N_24083,N_24704);
or U28044 (N_28044,N_21604,N_21943);
nor U28045 (N_28045,N_23235,N_24039);
or U28046 (N_28046,N_21286,N_24375);
nand U28047 (N_28047,N_22587,N_24163);
and U28048 (N_28048,N_23462,N_20487);
and U28049 (N_28049,N_22940,N_24834);
or U28050 (N_28050,N_21546,N_22991);
nand U28051 (N_28051,N_20955,N_23406);
or U28052 (N_28052,N_21358,N_21479);
and U28053 (N_28053,N_21229,N_24226);
and U28054 (N_28054,N_22423,N_20811);
and U28055 (N_28055,N_21311,N_22407);
and U28056 (N_28056,N_23321,N_23582);
xnor U28057 (N_28057,N_20724,N_20738);
or U28058 (N_28058,N_22789,N_24000);
nor U28059 (N_28059,N_23604,N_22572);
or U28060 (N_28060,N_23366,N_20662);
or U28061 (N_28061,N_21970,N_22656);
xnor U28062 (N_28062,N_24687,N_23289);
nor U28063 (N_28063,N_22831,N_20556);
or U28064 (N_28064,N_24574,N_23932);
or U28065 (N_28065,N_22544,N_23801);
nor U28066 (N_28066,N_22661,N_23077);
nor U28067 (N_28067,N_21360,N_23990);
or U28068 (N_28068,N_24275,N_24717);
nand U28069 (N_28069,N_24126,N_23490);
nand U28070 (N_28070,N_22970,N_21257);
and U28071 (N_28071,N_22017,N_23527);
and U28072 (N_28072,N_22217,N_23422);
and U28073 (N_28073,N_21981,N_23207);
nor U28074 (N_28074,N_24023,N_20553);
and U28075 (N_28075,N_24264,N_20386);
nand U28076 (N_28076,N_24984,N_22897);
or U28077 (N_28077,N_21952,N_20732);
xor U28078 (N_28078,N_23605,N_20469);
and U28079 (N_28079,N_24070,N_23487);
xnor U28080 (N_28080,N_24472,N_24273);
nor U28081 (N_28081,N_22673,N_22105);
xnor U28082 (N_28082,N_20423,N_21124);
or U28083 (N_28083,N_21043,N_22838);
nor U28084 (N_28084,N_21257,N_22991);
nor U28085 (N_28085,N_22404,N_20508);
nand U28086 (N_28086,N_24092,N_24030);
and U28087 (N_28087,N_24855,N_23018);
nand U28088 (N_28088,N_24838,N_23381);
xor U28089 (N_28089,N_23037,N_23997);
and U28090 (N_28090,N_21456,N_21056);
xnor U28091 (N_28091,N_21425,N_23761);
or U28092 (N_28092,N_21595,N_22011);
and U28093 (N_28093,N_20703,N_20068);
nand U28094 (N_28094,N_23938,N_24143);
or U28095 (N_28095,N_20824,N_22265);
xor U28096 (N_28096,N_24174,N_23508);
or U28097 (N_28097,N_24718,N_22767);
xor U28098 (N_28098,N_24533,N_23045);
xor U28099 (N_28099,N_22661,N_24156);
or U28100 (N_28100,N_24141,N_23092);
and U28101 (N_28101,N_20302,N_22120);
and U28102 (N_28102,N_21053,N_21347);
and U28103 (N_28103,N_21445,N_24376);
or U28104 (N_28104,N_20396,N_23366);
nand U28105 (N_28105,N_24672,N_22433);
nand U28106 (N_28106,N_21968,N_21772);
or U28107 (N_28107,N_20719,N_22020);
and U28108 (N_28108,N_24399,N_20378);
nand U28109 (N_28109,N_23194,N_24805);
nand U28110 (N_28110,N_21673,N_23710);
or U28111 (N_28111,N_24670,N_24890);
nor U28112 (N_28112,N_21066,N_22390);
nand U28113 (N_28113,N_24716,N_20555);
nand U28114 (N_28114,N_24841,N_22206);
nor U28115 (N_28115,N_21458,N_22714);
nand U28116 (N_28116,N_20081,N_23937);
xor U28117 (N_28117,N_23077,N_20329);
nor U28118 (N_28118,N_23162,N_21182);
nor U28119 (N_28119,N_22263,N_22667);
and U28120 (N_28120,N_21264,N_23122);
nand U28121 (N_28121,N_23080,N_23492);
nor U28122 (N_28122,N_24358,N_24738);
or U28123 (N_28123,N_22488,N_21124);
xor U28124 (N_28124,N_23223,N_24775);
nand U28125 (N_28125,N_21209,N_21190);
or U28126 (N_28126,N_24071,N_20217);
nand U28127 (N_28127,N_22010,N_21076);
and U28128 (N_28128,N_23910,N_23682);
nor U28129 (N_28129,N_21199,N_23075);
and U28130 (N_28130,N_24569,N_21684);
xor U28131 (N_28131,N_20402,N_21226);
and U28132 (N_28132,N_23314,N_23062);
and U28133 (N_28133,N_23174,N_24981);
or U28134 (N_28134,N_23725,N_22404);
or U28135 (N_28135,N_23233,N_23595);
nor U28136 (N_28136,N_24256,N_22971);
nand U28137 (N_28137,N_21560,N_23933);
nor U28138 (N_28138,N_24894,N_21416);
and U28139 (N_28139,N_22423,N_24698);
and U28140 (N_28140,N_20634,N_21814);
or U28141 (N_28141,N_20278,N_24512);
nand U28142 (N_28142,N_21620,N_24503);
or U28143 (N_28143,N_23267,N_21790);
xnor U28144 (N_28144,N_23700,N_24140);
xnor U28145 (N_28145,N_24874,N_23893);
or U28146 (N_28146,N_22386,N_20848);
and U28147 (N_28147,N_20543,N_20938);
nand U28148 (N_28148,N_22168,N_22669);
and U28149 (N_28149,N_22217,N_24803);
or U28150 (N_28150,N_23529,N_21839);
nand U28151 (N_28151,N_24598,N_23329);
or U28152 (N_28152,N_21006,N_21976);
nor U28153 (N_28153,N_21673,N_20115);
or U28154 (N_28154,N_20734,N_20562);
nand U28155 (N_28155,N_23624,N_21631);
and U28156 (N_28156,N_21413,N_23250);
nand U28157 (N_28157,N_22756,N_22275);
nand U28158 (N_28158,N_24516,N_22510);
nor U28159 (N_28159,N_24577,N_22456);
and U28160 (N_28160,N_23939,N_20132);
nor U28161 (N_28161,N_23146,N_20053);
or U28162 (N_28162,N_20271,N_21362);
and U28163 (N_28163,N_24955,N_24774);
and U28164 (N_28164,N_22622,N_23056);
and U28165 (N_28165,N_22422,N_23610);
nor U28166 (N_28166,N_21026,N_23118);
or U28167 (N_28167,N_24783,N_23629);
nand U28168 (N_28168,N_23450,N_24162);
and U28169 (N_28169,N_22514,N_24987);
nand U28170 (N_28170,N_22070,N_21366);
nand U28171 (N_28171,N_23225,N_24930);
or U28172 (N_28172,N_21790,N_21989);
or U28173 (N_28173,N_21280,N_21092);
nor U28174 (N_28174,N_24647,N_24050);
nand U28175 (N_28175,N_22512,N_20942);
or U28176 (N_28176,N_24173,N_22797);
nand U28177 (N_28177,N_23673,N_23970);
xnor U28178 (N_28178,N_22912,N_22457);
nand U28179 (N_28179,N_22221,N_24580);
nand U28180 (N_28180,N_20329,N_20469);
or U28181 (N_28181,N_24200,N_21437);
nor U28182 (N_28182,N_20837,N_23647);
nor U28183 (N_28183,N_20422,N_22368);
and U28184 (N_28184,N_21906,N_20049);
or U28185 (N_28185,N_24979,N_23242);
nand U28186 (N_28186,N_22335,N_20612);
or U28187 (N_28187,N_22304,N_20624);
xor U28188 (N_28188,N_23326,N_24379);
nand U28189 (N_28189,N_24068,N_20104);
and U28190 (N_28190,N_23858,N_24067);
and U28191 (N_28191,N_20505,N_20096);
nor U28192 (N_28192,N_24178,N_24277);
nor U28193 (N_28193,N_20898,N_21477);
xor U28194 (N_28194,N_22247,N_22510);
or U28195 (N_28195,N_23463,N_22926);
nor U28196 (N_28196,N_21209,N_24843);
nor U28197 (N_28197,N_22663,N_21478);
and U28198 (N_28198,N_20258,N_22059);
nor U28199 (N_28199,N_24094,N_23487);
or U28200 (N_28200,N_20540,N_22710);
nand U28201 (N_28201,N_23366,N_24821);
xnor U28202 (N_28202,N_20463,N_21905);
or U28203 (N_28203,N_24628,N_24140);
nor U28204 (N_28204,N_20323,N_23391);
or U28205 (N_28205,N_23583,N_24530);
nor U28206 (N_28206,N_21524,N_21705);
and U28207 (N_28207,N_21999,N_21267);
nor U28208 (N_28208,N_20133,N_21364);
and U28209 (N_28209,N_20178,N_23605);
or U28210 (N_28210,N_20586,N_23628);
nor U28211 (N_28211,N_21086,N_21408);
nor U28212 (N_28212,N_22001,N_22078);
or U28213 (N_28213,N_22549,N_21969);
nor U28214 (N_28214,N_24558,N_21827);
nand U28215 (N_28215,N_23533,N_24397);
and U28216 (N_28216,N_21052,N_21484);
nor U28217 (N_28217,N_20616,N_24516);
or U28218 (N_28218,N_22834,N_23404);
nand U28219 (N_28219,N_23850,N_20851);
xor U28220 (N_28220,N_21115,N_24200);
xnor U28221 (N_28221,N_21499,N_21600);
nand U28222 (N_28222,N_23222,N_20912);
or U28223 (N_28223,N_21692,N_22306);
or U28224 (N_28224,N_22427,N_21472);
xor U28225 (N_28225,N_21930,N_21143);
or U28226 (N_28226,N_23310,N_22677);
nor U28227 (N_28227,N_24235,N_21920);
or U28228 (N_28228,N_24525,N_23361);
and U28229 (N_28229,N_24431,N_23409);
or U28230 (N_28230,N_22816,N_24697);
nor U28231 (N_28231,N_20187,N_21780);
or U28232 (N_28232,N_22131,N_22775);
nor U28233 (N_28233,N_21924,N_23512);
nand U28234 (N_28234,N_23681,N_24734);
and U28235 (N_28235,N_22895,N_24745);
nor U28236 (N_28236,N_24927,N_22264);
nand U28237 (N_28237,N_20154,N_23060);
or U28238 (N_28238,N_20928,N_23657);
or U28239 (N_28239,N_22881,N_22849);
nor U28240 (N_28240,N_23810,N_23203);
nand U28241 (N_28241,N_23988,N_23181);
nand U28242 (N_28242,N_20178,N_20236);
nand U28243 (N_28243,N_22067,N_22877);
and U28244 (N_28244,N_22524,N_24115);
and U28245 (N_28245,N_23271,N_24735);
nand U28246 (N_28246,N_24771,N_22507);
xnor U28247 (N_28247,N_22049,N_21008);
and U28248 (N_28248,N_24871,N_21141);
and U28249 (N_28249,N_20185,N_21100);
nand U28250 (N_28250,N_21140,N_24971);
and U28251 (N_28251,N_20091,N_20842);
xnor U28252 (N_28252,N_23493,N_21446);
nand U28253 (N_28253,N_21863,N_21053);
and U28254 (N_28254,N_21248,N_20593);
and U28255 (N_28255,N_22974,N_22654);
and U28256 (N_28256,N_22842,N_20697);
or U28257 (N_28257,N_20422,N_22384);
nand U28258 (N_28258,N_21267,N_21079);
and U28259 (N_28259,N_21895,N_24667);
nor U28260 (N_28260,N_20941,N_24154);
and U28261 (N_28261,N_20331,N_20422);
nor U28262 (N_28262,N_20299,N_20226);
nor U28263 (N_28263,N_24037,N_21374);
nand U28264 (N_28264,N_23787,N_24452);
nand U28265 (N_28265,N_20128,N_20029);
or U28266 (N_28266,N_23579,N_22961);
and U28267 (N_28267,N_23943,N_21318);
nand U28268 (N_28268,N_20596,N_20853);
nand U28269 (N_28269,N_22369,N_24503);
or U28270 (N_28270,N_20316,N_20761);
nand U28271 (N_28271,N_23654,N_21552);
nand U28272 (N_28272,N_22163,N_23396);
xnor U28273 (N_28273,N_21316,N_21630);
or U28274 (N_28274,N_20092,N_23891);
nand U28275 (N_28275,N_21387,N_22210);
and U28276 (N_28276,N_20741,N_23856);
or U28277 (N_28277,N_23542,N_24699);
nor U28278 (N_28278,N_22295,N_23533);
and U28279 (N_28279,N_21585,N_21420);
and U28280 (N_28280,N_21978,N_24252);
or U28281 (N_28281,N_21093,N_24547);
nand U28282 (N_28282,N_20657,N_24872);
or U28283 (N_28283,N_23628,N_21098);
and U28284 (N_28284,N_21457,N_20986);
nor U28285 (N_28285,N_22843,N_23833);
nor U28286 (N_28286,N_23730,N_21267);
or U28287 (N_28287,N_23160,N_23294);
nand U28288 (N_28288,N_23316,N_24087);
nand U28289 (N_28289,N_23010,N_22422);
and U28290 (N_28290,N_20927,N_24045);
and U28291 (N_28291,N_23221,N_22770);
or U28292 (N_28292,N_22954,N_24920);
nor U28293 (N_28293,N_24830,N_23430);
xnor U28294 (N_28294,N_22757,N_22269);
xor U28295 (N_28295,N_23998,N_22904);
nand U28296 (N_28296,N_24674,N_21346);
nand U28297 (N_28297,N_20192,N_24615);
and U28298 (N_28298,N_21915,N_24835);
or U28299 (N_28299,N_23672,N_24139);
or U28300 (N_28300,N_23419,N_23053);
xnor U28301 (N_28301,N_20783,N_24732);
nand U28302 (N_28302,N_22854,N_24325);
and U28303 (N_28303,N_21139,N_23964);
or U28304 (N_28304,N_22829,N_20292);
nand U28305 (N_28305,N_23992,N_24762);
nor U28306 (N_28306,N_23834,N_20798);
xnor U28307 (N_28307,N_23109,N_21991);
nand U28308 (N_28308,N_20063,N_24036);
and U28309 (N_28309,N_22135,N_21821);
xnor U28310 (N_28310,N_24340,N_20123);
and U28311 (N_28311,N_21106,N_23466);
nor U28312 (N_28312,N_23021,N_24613);
and U28313 (N_28313,N_21187,N_21322);
and U28314 (N_28314,N_23052,N_23552);
or U28315 (N_28315,N_24209,N_23157);
or U28316 (N_28316,N_21588,N_20667);
nor U28317 (N_28317,N_21647,N_20857);
or U28318 (N_28318,N_22422,N_23521);
nand U28319 (N_28319,N_21203,N_24938);
nor U28320 (N_28320,N_20899,N_22630);
nand U28321 (N_28321,N_23443,N_23888);
xor U28322 (N_28322,N_20153,N_24986);
nor U28323 (N_28323,N_21145,N_24628);
nor U28324 (N_28324,N_20277,N_20774);
or U28325 (N_28325,N_24596,N_23108);
and U28326 (N_28326,N_24244,N_24148);
nor U28327 (N_28327,N_23825,N_20615);
xor U28328 (N_28328,N_21980,N_22664);
nand U28329 (N_28329,N_23840,N_24359);
xnor U28330 (N_28330,N_24960,N_23623);
nor U28331 (N_28331,N_20844,N_20412);
nand U28332 (N_28332,N_20024,N_22992);
or U28333 (N_28333,N_22859,N_24547);
nand U28334 (N_28334,N_23785,N_21970);
nor U28335 (N_28335,N_21998,N_24945);
nand U28336 (N_28336,N_20851,N_20347);
and U28337 (N_28337,N_20510,N_24597);
nand U28338 (N_28338,N_22975,N_24879);
nor U28339 (N_28339,N_20833,N_22138);
and U28340 (N_28340,N_22904,N_21166);
or U28341 (N_28341,N_20088,N_20854);
or U28342 (N_28342,N_21344,N_24978);
and U28343 (N_28343,N_24371,N_20378);
nand U28344 (N_28344,N_23926,N_22556);
nand U28345 (N_28345,N_24219,N_21719);
nand U28346 (N_28346,N_23355,N_23815);
and U28347 (N_28347,N_20284,N_24948);
nor U28348 (N_28348,N_20240,N_24424);
xnor U28349 (N_28349,N_21247,N_23525);
or U28350 (N_28350,N_22550,N_22119);
nand U28351 (N_28351,N_22334,N_24739);
and U28352 (N_28352,N_20812,N_23733);
or U28353 (N_28353,N_24051,N_24267);
and U28354 (N_28354,N_24104,N_24688);
nor U28355 (N_28355,N_20972,N_23190);
nor U28356 (N_28356,N_22781,N_21131);
nor U28357 (N_28357,N_24661,N_20105);
and U28358 (N_28358,N_23895,N_22654);
or U28359 (N_28359,N_24164,N_22444);
and U28360 (N_28360,N_21145,N_21021);
or U28361 (N_28361,N_20480,N_21686);
or U28362 (N_28362,N_23155,N_24953);
nand U28363 (N_28363,N_24055,N_24384);
nand U28364 (N_28364,N_22931,N_21086);
nand U28365 (N_28365,N_20062,N_22766);
and U28366 (N_28366,N_20551,N_21198);
nor U28367 (N_28367,N_24427,N_23579);
nor U28368 (N_28368,N_21857,N_22295);
and U28369 (N_28369,N_22023,N_23996);
nor U28370 (N_28370,N_20901,N_20520);
and U28371 (N_28371,N_22419,N_21083);
nand U28372 (N_28372,N_20978,N_22764);
and U28373 (N_28373,N_23434,N_23958);
or U28374 (N_28374,N_20202,N_20739);
or U28375 (N_28375,N_23430,N_23221);
nor U28376 (N_28376,N_21849,N_24197);
xor U28377 (N_28377,N_20281,N_23216);
or U28378 (N_28378,N_20726,N_22611);
and U28379 (N_28379,N_20665,N_20668);
nor U28380 (N_28380,N_23577,N_24590);
and U28381 (N_28381,N_23878,N_24918);
nor U28382 (N_28382,N_23993,N_23571);
and U28383 (N_28383,N_22949,N_21559);
nor U28384 (N_28384,N_23584,N_20966);
nor U28385 (N_28385,N_20511,N_22436);
or U28386 (N_28386,N_24995,N_22190);
and U28387 (N_28387,N_22182,N_21528);
nor U28388 (N_28388,N_20196,N_20329);
nand U28389 (N_28389,N_20190,N_23746);
nor U28390 (N_28390,N_20182,N_20283);
nor U28391 (N_28391,N_22655,N_21681);
nor U28392 (N_28392,N_20456,N_24042);
nand U28393 (N_28393,N_21335,N_22796);
nand U28394 (N_28394,N_20615,N_22622);
and U28395 (N_28395,N_24395,N_20129);
xor U28396 (N_28396,N_20578,N_22975);
nor U28397 (N_28397,N_21813,N_20556);
and U28398 (N_28398,N_21003,N_22997);
and U28399 (N_28399,N_24133,N_20232);
nand U28400 (N_28400,N_22956,N_21595);
nand U28401 (N_28401,N_24711,N_20460);
nand U28402 (N_28402,N_21506,N_24973);
nand U28403 (N_28403,N_24004,N_22331);
nand U28404 (N_28404,N_20015,N_22221);
or U28405 (N_28405,N_24308,N_20553);
or U28406 (N_28406,N_24953,N_22288);
nand U28407 (N_28407,N_22198,N_22867);
nor U28408 (N_28408,N_23166,N_24553);
and U28409 (N_28409,N_24544,N_23595);
and U28410 (N_28410,N_22156,N_24048);
nor U28411 (N_28411,N_22270,N_21128);
or U28412 (N_28412,N_23281,N_23921);
nor U28413 (N_28413,N_22758,N_22727);
nand U28414 (N_28414,N_21670,N_21742);
xor U28415 (N_28415,N_24398,N_23753);
or U28416 (N_28416,N_24619,N_21557);
or U28417 (N_28417,N_24946,N_24256);
and U28418 (N_28418,N_22928,N_24290);
or U28419 (N_28419,N_21154,N_24003);
nor U28420 (N_28420,N_24496,N_20995);
and U28421 (N_28421,N_23983,N_23080);
or U28422 (N_28422,N_22901,N_20971);
nor U28423 (N_28423,N_22669,N_22475);
nand U28424 (N_28424,N_24092,N_22590);
nand U28425 (N_28425,N_20650,N_21007);
nor U28426 (N_28426,N_21443,N_24001);
xnor U28427 (N_28427,N_22568,N_22425);
nor U28428 (N_28428,N_21246,N_21434);
nand U28429 (N_28429,N_20838,N_22908);
nor U28430 (N_28430,N_23701,N_22910);
xor U28431 (N_28431,N_21234,N_23578);
or U28432 (N_28432,N_22469,N_23395);
or U28433 (N_28433,N_23852,N_24231);
nor U28434 (N_28434,N_22086,N_21399);
nor U28435 (N_28435,N_20855,N_22361);
nor U28436 (N_28436,N_22083,N_21752);
or U28437 (N_28437,N_20877,N_22639);
nor U28438 (N_28438,N_21900,N_24605);
nand U28439 (N_28439,N_23191,N_21645);
nor U28440 (N_28440,N_21656,N_24711);
and U28441 (N_28441,N_22624,N_21403);
nand U28442 (N_28442,N_20363,N_22662);
and U28443 (N_28443,N_21811,N_22262);
nand U28444 (N_28444,N_21572,N_24655);
or U28445 (N_28445,N_20144,N_22810);
nor U28446 (N_28446,N_21412,N_22196);
or U28447 (N_28447,N_23018,N_22156);
or U28448 (N_28448,N_22312,N_24268);
nand U28449 (N_28449,N_21569,N_22488);
and U28450 (N_28450,N_20718,N_23713);
or U28451 (N_28451,N_22794,N_21290);
and U28452 (N_28452,N_21659,N_21519);
nor U28453 (N_28453,N_24327,N_23477);
and U28454 (N_28454,N_20685,N_21191);
nor U28455 (N_28455,N_24778,N_20056);
nor U28456 (N_28456,N_23391,N_23273);
nand U28457 (N_28457,N_24207,N_22205);
or U28458 (N_28458,N_21923,N_21189);
and U28459 (N_28459,N_20630,N_24285);
and U28460 (N_28460,N_21145,N_21773);
and U28461 (N_28461,N_21768,N_22412);
xor U28462 (N_28462,N_24235,N_22810);
nor U28463 (N_28463,N_20637,N_24862);
nor U28464 (N_28464,N_24845,N_20064);
and U28465 (N_28465,N_22062,N_23575);
and U28466 (N_28466,N_21131,N_21494);
nand U28467 (N_28467,N_20302,N_23228);
nor U28468 (N_28468,N_21283,N_20380);
nor U28469 (N_28469,N_23121,N_24524);
nand U28470 (N_28470,N_23464,N_22694);
nor U28471 (N_28471,N_22429,N_23760);
nor U28472 (N_28472,N_22762,N_23577);
or U28473 (N_28473,N_22395,N_21763);
nor U28474 (N_28474,N_21470,N_24261);
nand U28475 (N_28475,N_22634,N_24156);
and U28476 (N_28476,N_21606,N_23605);
nor U28477 (N_28477,N_23368,N_22768);
nand U28478 (N_28478,N_22489,N_20466);
xor U28479 (N_28479,N_20300,N_24643);
nand U28480 (N_28480,N_24248,N_20559);
or U28481 (N_28481,N_23037,N_23308);
nor U28482 (N_28482,N_21491,N_24552);
and U28483 (N_28483,N_24420,N_20249);
or U28484 (N_28484,N_22828,N_21781);
and U28485 (N_28485,N_20927,N_21557);
or U28486 (N_28486,N_21193,N_21515);
nor U28487 (N_28487,N_21542,N_21646);
xnor U28488 (N_28488,N_24465,N_21272);
nand U28489 (N_28489,N_21094,N_24555);
and U28490 (N_28490,N_22134,N_20260);
nand U28491 (N_28491,N_22698,N_23872);
nand U28492 (N_28492,N_24900,N_22457);
nand U28493 (N_28493,N_23515,N_23017);
nand U28494 (N_28494,N_23288,N_20935);
and U28495 (N_28495,N_22446,N_20185);
nor U28496 (N_28496,N_24240,N_24162);
nor U28497 (N_28497,N_20627,N_22761);
and U28498 (N_28498,N_23856,N_23910);
and U28499 (N_28499,N_23704,N_22680);
nand U28500 (N_28500,N_20079,N_20537);
or U28501 (N_28501,N_24342,N_23836);
xnor U28502 (N_28502,N_21511,N_21103);
and U28503 (N_28503,N_20267,N_21311);
or U28504 (N_28504,N_22353,N_23815);
or U28505 (N_28505,N_20112,N_23865);
and U28506 (N_28506,N_23080,N_23058);
nand U28507 (N_28507,N_23774,N_22934);
nor U28508 (N_28508,N_22268,N_20541);
xnor U28509 (N_28509,N_23725,N_22712);
or U28510 (N_28510,N_22393,N_23065);
and U28511 (N_28511,N_20722,N_20146);
nor U28512 (N_28512,N_24925,N_23646);
nand U28513 (N_28513,N_20292,N_22073);
or U28514 (N_28514,N_23312,N_22681);
nor U28515 (N_28515,N_21635,N_23444);
or U28516 (N_28516,N_24183,N_24296);
nor U28517 (N_28517,N_23500,N_24316);
nand U28518 (N_28518,N_20722,N_20901);
xor U28519 (N_28519,N_22224,N_21694);
nand U28520 (N_28520,N_24940,N_23470);
nand U28521 (N_28521,N_24470,N_23274);
nand U28522 (N_28522,N_24225,N_20106);
and U28523 (N_28523,N_21399,N_24933);
and U28524 (N_28524,N_21644,N_24752);
and U28525 (N_28525,N_23589,N_20779);
nor U28526 (N_28526,N_22417,N_21495);
and U28527 (N_28527,N_22379,N_22633);
or U28528 (N_28528,N_23027,N_21088);
nor U28529 (N_28529,N_24934,N_23349);
xor U28530 (N_28530,N_21508,N_24172);
or U28531 (N_28531,N_20806,N_20879);
or U28532 (N_28532,N_22072,N_24273);
and U28533 (N_28533,N_20473,N_24908);
nand U28534 (N_28534,N_24228,N_20563);
nor U28535 (N_28535,N_24365,N_23539);
or U28536 (N_28536,N_21886,N_23594);
nor U28537 (N_28537,N_24458,N_22614);
or U28538 (N_28538,N_21862,N_23292);
nor U28539 (N_28539,N_20289,N_24369);
or U28540 (N_28540,N_21837,N_24342);
nor U28541 (N_28541,N_20164,N_23708);
or U28542 (N_28542,N_20641,N_20149);
and U28543 (N_28543,N_24977,N_21675);
xor U28544 (N_28544,N_22052,N_24117);
nand U28545 (N_28545,N_23249,N_21470);
and U28546 (N_28546,N_20079,N_20831);
xor U28547 (N_28547,N_21900,N_24343);
nor U28548 (N_28548,N_23146,N_22406);
nand U28549 (N_28549,N_20389,N_22311);
nor U28550 (N_28550,N_20436,N_24731);
or U28551 (N_28551,N_23344,N_23157);
nand U28552 (N_28552,N_21107,N_23976);
or U28553 (N_28553,N_24605,N_24571);
or U28554 (N_28554,N_20423,N_20870);
or U28555 (N_28555,N_23337,N_22485);
and U28556 (N_28556,N_22278,N_22642);
or U28557 (N_28557,N_24320,N_23036);
or U28558 (N_28558,N_23683,N_21590);
or U28559 (N_28559,N_23870,N_24062);
or U28560 (N_28560,N_23271,N_22584);
xnor U28561 (N_28561,N_21668,N_23893);
nand U28562 (N_28562,N_24293,N_21043);
nor U28563 (N_28563,N_23880,N_22058);
nor U28564 (N_28564,N_21973,N_23831);
nor U28565 (N_28565,N_20860,N_20541);
nand U28566 (N_28566,N_20743,N_22586);
or U28567 (N_28567,N_23423,N_20284);
or U28568 (N_28568,N_20597,N_22932);
nor U28569 (N_28569,N_23396,N_24881);
nand U28570 (N_28570,N_20638,N_21187);
nor U28571 (N_28571,N_22279,N_23852);
nand U28572 (N_28572,N_20283,N_23513);
and U28573 (N_28573,N_20766,N_24978);
nor U28574 (N_28574,N_24564,N_22554);
nor U28575 (N_28575,N_23337,N_23480);
and U28576 (N_28576,N_20545,N_20228);
nor U28577 (N_28577,N_24952,N_22514);
nand U28578 (N_28578,N_22450,N_23416);
or U28579 (N_28579,N_21254,N_22888);
and U28580 (N_28580,N_20805,N_21773);
nor U28581 (N_28581,N_20121,N_24885);
and U28582 (N_28582,N_21764,N_24530);
nand U28583 (N_28583,N_20728,N_21176);
nand U28584 (N_28584,N_22108,N_21849);
nand U28585 (N_28585,N_22435,N_24271);
nand U28586 (N_28586,N_24267,N_20217);
or U28587 (N_28587,N_24436,N_23506);
nand U28588 (N_28588,N_20156,N_24597);
and U28589 (N_28589,N_24243,N_23355);
nor U28590 (N_28590,N_22313,N_24680);
nand U28591 (N_28591,N_20681,N_21206);
nor U28592 (N_28592,N_20984,N_21282);
nand U28593 (N_28593,N_22333,N_24950);
nor U28594 (N_28594,N_23154,N_24579);
nor U28595 (N_28595,N_21976,N_22980);
or U28596 (N_28596,N_21085,N_21758);
nor U28597 (N_28597,N_23127,N_21620);
nor U28598 (N_28598,N_20592,N_20503);
and U28599 (N_28599,N_22005,N_23002);
xor U28600 (N_28600,N_24892,N_21539);
nand U28601 (N_28601,N_24789,N_22261);
nand U28602 (N_28602,N_22571,N_22527);
nand U28603 (N_28603,N_20119,N_20983);
or U28604 (N_28604,N_21723,N_21318);
nand U28605 (N_28605,N_23285,N_24869);
nor U28606 (N_28606,N_24954,N_24833);
and U28607 (N_28607,N_24937,N_21724);
nor U28608 (N_28608,N_23741,N_20349);
nor U28609 (N_28609,N_23467,N_20570);
or U28610 (N_28610,N_21830,N_23562);
xnor U28611 (N_28611,N_24138,N_24596);
nand U28612 (N_28612,N_23981,N_21114);
nand U28613 (N_28613,N_20501,N_24806);
nand U28614 (N_28614,N_24655,N_23064);
and U28615 (N_28615,N_21593,N_20822);
or U28616 (N_28616,N_21339,N_20221);
and U28617 (N_28617,N_22208,N_21359);
and U28618 (N_28618,N_20102,N_24028);
nor U28619 (N_28619,N_22425,N_22864);
and U28620 (N_28620,N_21968,N_24722);
or U28621 (N_28621,N_24921,N_23282);
or U28622 (N_28622,N_20713,N_23281);
nor U28623 (N_28623,N_24725,N_22464);
or U28624 (N_28624,N_20416,N_20117);
or U28625 (N_28625,N_22544,N_23067);
and U28626 (N_28626,N_23727,N_23902);
or U28627 (N_28627,N_22093,N_22762);
xor U28628 (N_28628,N_21617,N_20951);
nand U28629 (N_28629,N_24466,N_24289);
and U28630 (N_28630,N_21383,N_21887);
or U28631 (N_28631,N_20679,N_21149);
nor U28632 (N_28632,N_24733,N_24658);
nor U28633 (N_28633,N_20559,N_23801);
nand U28634 (N_28634,N_24456,N_24929);
nor U28635 (N_28635,N_23413,N_22187);
xnor U28636 (N_28636,N_22158,N_23701);
nor U28637 (N_28637,N_23312,N_21835);
or U28638 (N_28638,N_20971,N_21181);
and U28639 (N_28639,N_20863,N_21292);
nor U28640 (N_28640,N_22354,N_21500);
xnor U28641 (N_28641,N_21536,N_23554);
and U28642 (N_28642,N_20080,N_21117);
and U28643 (N_28643,N_24762,N_20777);
nor U28644 (N_28644,N_22308,N_23047);
or U28645 (N_28645,N_21626,N_20320);
or U28646 (N_28646,N_22444,N_22199);
and U28647 (N_28647,N_24661,N_23616);
nand U28648 (N_28648,N_24933,N_24666);
nand U28649 (N_28649,N_21156,N_22977);
or U28650 (N_28650,N_21237,N_24772);
xnor U28651 (N_28651,N_23799,N_21980);
xnor U28652 (N_28652,N_24204,N_21432);
nand U28653 (N_28653,N_21276,N_23470);
and U28654 (N_28654,N_21209,N_23228);
nand U28655 (N_28655,N_23112,N_20854);
nand U28656 (N_28656,N_23073,N_23992);
and U28657 (N_28657,N_20487,N_22201);
or U28658 (N_28658,N_22970,N_24810);
and U28659 (N_28659,N_20383,N_22572);
and U28660 (N_28660,N_23469,N_20562);
nand U28661 (N_28661,N_20132,N_22851);
or U28662 (N_28662,N_24974,N_21808);
xnor U28663 (N_28663,N_20517,N_21382);
nor U28664 (N_28664,N_22578,N_21580);
and U28665 (N_28665,N_21832,N_21343);
nand U28666 (N_28666,N_21599,N_21024);
nand U28667 (N_28667,N_22527,N_20616);
or U28668 (N_28668,N_20334,N_23860);
nor U28669 (N_28669,N_21519,N_21861);
or U28670 (N_28670,N_23576,N_21805);
or U28671 (N_28671,N_20695,N_20458);
nand U28672 (N_28672,N_20612,N_21496);
or U28673 (N_28673,N_20996,N_20961);
or U28674 (N_28674,N_22118,N_21882);
or U28675 (N_28675,N_23339,N_22059);
nor U28676 (N_28676,N_23280,N_23477);
or U28677 (N_28677,N_23669,N_24713);
xor U28678 (N_28678,N_23901,N_20123);
nand U28679 (N_28679,N_23237,N_23783);
and U28680 (N_28680,N_20444,N_22467);
or U28681 (N_28681,N_20770,N_23866);
or U28682 (N_28682,N_20204,N_21626);
and U28683 (N_28683,N_20570,N_21318);
xnor U28684 (N_28684,N_24575,N_21253);
and U28685 (N_28685,N_20738,N_23889);
nor U28686 (N_28686,N_21838,N_21040);
or U28687 (N_28687,N_24468,N_23961);
nand U28688 (N_28688,N_22985,N_22215);
and U28689 (N_28689,N_23837,N_21606);
or U28690 (N_28690,N_23420,N_24816);
xor U28691 (N_28691,N_20824,N_20501);
and U28692 (N_28692,N_22865,N_22449);
or U28693 (N_28693,N_22740,N_23399);
and U28694 (N_28694,N_23431,N_24706);
xor U28695 (N_28695,N_23861,N_24628);
or U28696 (N_28696,N_23929,N_22817);
or U28697 (N_28697,N_24616,N_20880);
nor U28698 (N_28698,N_22307,N_20737);
nand U28699 (N_28699,N_23007,N_24985);
nand U28700 (N_28700,N_21090,N_20846);
nand U28701 (N_28701,N_24880,N_20366);
or U28702 (N_28702,N_23965,N_22669);
and U28703 (N_28703,N_21152,N_20961);
nor U28704 (N_28704,N_21737,N_20917);
or U28705 (N_28705,N_21276,N_23845);
or U28706 (N_28706,N_24390,N_21605);
nand U28707 (N_28707,N_21075,N_23492);
xnor U28708 (N_28708,N_24348,N_20245);
or U28709 (N_28709,N_21631,N_21597);
or U28710 (N_28710,N_20261,N_24551);
or U28711 (N_28711,N_20847,N_22603);
nor U28712 (N_28712,N_23903,N_22416);
nand U28713 (N_28713,N_23852,N_21622);
nor U28714 (N_28714,N_21615,N_20219);
nand U28715 (N_28715,N_22570,N_21171);
nand U28716 (N_28716,N_20124,N_23592);
nand U28717 (N_28717,N_24595,N_24645);
nor U28718 (N_28718,N_20921,N_20881);
and U28719 (N_28719,N_22209,N_22644);
or U28720 (N_28720,N_22888,N_20696);
or U28721 (N_28721,N_22596,N_22773);
and U28722 (N_28722,N_20272,N_24031);
nor U28723 (N_28723,N_21611,N_22705);
xnor U28724 (N_28724,N_22994,N_23764);
nor U28725 (N_28725,N_22670,N_21554);
and U28726 (N_28726,N_20173,N_23978);
and U28727 (N_28727,N_20678,N_23518);
xnor U28728 (N_28728,N_20409,N_22287);
nor U28729 (N_28729,N_20901,N_22169);
and U28730 (N_28730,N_20090,N_23026);
or U28731 (N_28731,N_23137,N_21237);
or U28732 (N_28732,N_20349,N_20632);
nand U28733 (N_28733,N_23346,N_23516);
xor U28734 (N_28734,N_24048,N_21877);
or U28735 (N_28735,N_22123,N_23162);
nand U28736 (N_28736,N_21126,N_20972);
and U28737 (N_28737,N_21690,N_21470);
nand U28738 (N_28738,N_23574,N_21171);
and U28739 (N_28739,N_23815,N_22951);
nor U28740 (N_28740,N_21645,N_21027);
nand U28741 (N_28741,N_22191,N_22488);
nand U28742 (N_28742,N_23847,N_21219);
nand U28743 (N_28743,N_21962,N_22627);
and U28744 (N_28744,N_20152,N_23007);
or U28745 (N_28745,N_24459,N_20934);
and U28746 (N_28746,N_24277,N_22996);
or U28747 (N_28747,N_23534,N_23475);
or U28748 (N_28748,N_20534,N_23625);
and U28749 (N_28749,N_21358,N_24596);
and U28750 (N_28750,N_24340,N_24096);
nor U28751 (N_28751,N_20839,N_20298);
nor U28752 (N_28752,N_23517,N_21565);
or U28753 (N_28753,N_24180,N_23505);
nor U28754 (N_28754,N_22136,N_20738);
nand U28755 (N_28755,N_21125,N_20907);
nor U28756 (N_28756,N_21152,N_23245);
and U28757 (N_28757,N_21360,N_20402);
xnor U28758 (N_28758,N_21675,N_23524);
nor U28759 (N_28759,N_22441,N_24273);
and U28760 (N_28760,N_20965,N_21167);
nor U28761 (N_28761,N_21728,N_21371);
nor U28762 (N_28762,N_24494,N_21092);
nor U28763 (N_28763,N_20419,N_22632);
nor U28764 (N_28764,N_22924,N_23064);
or U28765 (N_28765,N_20845,N_24246);
and U28766 (N_28766,N_21949,N_24255);
nand U28767 (N_28767,N_20966,N_21727);
and U28768 (N_28768,N_24911,N_21745);
and U28769 (N_28769,N_24718,N_23098);
nand U28770 (N_28770,N_22960,N_23093);
nand U28771 (N_28771,N_24514,N_20391);
nand U28772 (N_28772,N_22475,N_20934);
nor U28773 (N_28773,N_22100,N_22633);
and U28774 (N_28774,N_24184,N_20248);
xor U28775 (N_28775,N_22386,N_22420);
or U28776 (N_28776,N_20257,N_22850);
nand U28777 (N_28777,N_24708,N_20630);
nand U28778 (N_28778,N_21290,N_22044);
nand U28779 (N_28779,N_21032,N_20688);
and U28780 (N_28780,N_23801,N_20317);
nor U28781 (N_28781,N_22423,N_20786);
or U28782 (N_28782,N_20720,N_22869);
or U28783 (N_28783,N_23413,N_24817);
or U28784 (N_28784,N_24309,N_21786);
or U28785 (N_28785,N_20279,N_23644);
nand U28786 (N_28786,N_23583,N_24187);
nand U28787 (N_28787,N_22173,N_20146);
xor U28788 (N_28788,N_24795,N_22777);
nor U28789 (N_28789,N_24473,N_23650);
nor U28790 (N_28790,N_24849,N_22147);
nand U28791 (N_28791,N_22803,N_21819);
nand U28792 (N_28792,N_21985,N_20452);
xnor U28793 (N_28793,N_21224,N_20420);
nand U28794 (N_28794,N_20699,N_21727);
nand U28795 (N_28795,N_24793,N_24051);
or U28796 (N_28796,N_22710,N_22695);
nor U28797 (N_28797,N_23887,N_22625);
xnor U28798 (N_28798,N_23258,N_22052);
or U28799 (N_28799,N_22614,N_24346);
and U28800 (N_28800,N_21428,N_20185);
nand U28801 (N_28801,N_22430,N_22464);
nor U28802 (N_28802,N_21120,N_23700);
nand U28803 (N_28803,N_23144,N_24572);
nor U28804 (N_28804,N_21891,N_24752);
or U28805 (N_28805,N_22310,N_22659);
nor U28806 (N_28806,N_20366,N_21685);
nor U28807 (N_28807,N_20438,N_24935);
nand U28808 (N_28808,N_21261,N_24220);
xor U28809 (N_28809,N_23889,N_21442);
nor U28810 (N_28810,N_21550,N_24876);
nor U28811 (N_28811,N_23105,N_24398);
nand U28812 (N_28812,N_21806,N_21253);
or U28813 (N_28813,N_24924,N_24055);
nor U28814 (N_28814,N_21447,N_20898);
and U28815 (N_28815,N_24587,N_23065);
nand U28816 (N_28816,N_20801,N_21976);
xor U28817 (N_28817,N_23570,N_21140);
and U28818 (N_28818,N_22563,N_22794);
or U28819 (N_28819,N_20558,N_22759);
and U28820 (N_28820,N_22859,N_20057);
nand U28821 (N_28821,N_23937,N_22560);
nand U28822 (N_28822,N_23658,N_21943);
nand U28823 (N_28823,N_21830,N_23800);
and U28824 (N_28824,N_24081,N_20408);
or U28825 (N_28825,N_21127,N_22794);
xor U28826 (N_28826,N_23836,N_20099);
xnor U28827 (N_28827,N_20290,N_20562);
nand U28828 (N_28828,N_23992,N_22610);
nor U28829 (N_28829,N_21713,N_20355);
nor U28830 (N_28830,N_24803,N_22813);
nor U28831 (N_28831,N_23904,N_22475);
nand U28832 (N_28832,N_22201,N_22360);
nand U28833 (N_28833,N_23666,N_21872);
nand U28834 (N_28834,N_21580,N_21924);
or U28835 (N_28835,N_20846,N_23899);
nand U28836 (N_28836,N_21200,N_23648);
and U28837 (N_28837,N_22365,N_22085);
nand U28838 (N_28838,N_23693,N_23615);
and U28839 (N_28839,N_20996,N_20516);
or U28840 (N_28840,N_24747,N_24319);
or U28841 (N_28841,N_24126,N_22646);
or U28842 (N_28842,N_20344,N_24391);
xnor U28843 (N_28843,N_22342,N_24440);
nand U28844 (N_28844,N_20803,N_22276);
and U28845 (N_28845,N_22112,N_23070);
and U28846 (N_28846,N_23923,N_21498);
nor U28847 (N_28847,N_23190,N_20857);
or U28848 (N_28848,N_23477,N_21792);
and U28849 (N_28849,N_23323,N_23297);
or U28850 (N_28850,N_22763,N_22086);
nand U28851 (N_28851,N_24387,N_20180);
nor U28852 (N_28852,N_21469,N_23519);
nor U28853 (N_28853,N_24927,N_23812);
nor U28854 (N_28854,N_22109,N_23140);
nand U28855 (N_28855,N_23294,N_22036);
and U28856 (N_28856,N_22105,N_23630);
nand U28857 (N_28857,N_24043,N_23303);
nor U28858 (N_28858,N_23368,N_23579);
nand U28859 (N_28859,N_24233,N_23268);
nand U28860 (N_28860,N_20685,N_21216);
nor U28861 (N_28861,N_23797,N_22719);
and U28862 (N_28862,N_21843,N_20591);
nor U28863 (N_28863,N_22818,N_23320);
nand U28864 (N_28864,N_23337,N_24927);
xnor U28865 (N_28865,N_20498,N_24536);
nor U28866 (N_28866,N_24653,N_21411);
and U28867 (N_28867,N_20540,N_21096);
or U28868 (N_28868,N_24409,N_21365);
and U28869 (N_28869,N_20995,N_22079);
xor U28870 (N_28870,N_20426,N_22302);
or U28871 (N_28871,N_20168,N_24031);
nor U28872 (N_28872,N_23124,N_22744);
and U28873 (N_28873,N_24380,N_24177);
and U28874 (N_28874,N_20240,N_21601);
nand U28875 (N_28875,N_23049,N_22917);
or U28876 (N_28876,N_24751,N_23608);
or U28877 (N_28877,N_23954,N_23896);
or U28878 (N_28878,N_22633,N_24895);
xnor U28879 (N_28879,N_20563,N_24893);
nand U28880 (N_28880,N_21497,N_23309);
nor U28881 (N_28881,N_21647,N_23030);
or U28882 (N_28882,N_20465,N_22582);
or U28883 (N_28883,N_22911,N_21790);
nor U28884 (N_28884,N_20425,N_24321);
nor U28885 (N_28885,N_23145,N_21097);
nand U28886 (N_28886,N_23465,N_20396);
nor U28887 (N_28887,N_20882,N_21216);
xor U28888 (N_28888,N_21890,N_24870);
nor U28889 (N_28889,N_21844,N_23635);
nand U28890 (N_28890,N_20503,N_24870);
and U28891 (N_28891,N_21275,N_23413);
nor U28892 (N_28892,N_22045,N_21561);
and U28893 (N_28893,N_20554,N_24002);
and U28894 (N_28894,N_22651,N_21755);
nor U28895 (N_28895,N_22652,N_21298);
or U28896 (N_28896,N_21549,N_20109);
nand U28897 (N_28897,N_22499,N_20083);
or U28898 (N_28898,N_24361,N_22441);
or U28899 (N_28899,N_22999,N_22875);
nor U28900 (N_28900,N_22452,N_20981);
or U28901 (N_28901,N_22304,N_24472);
xnor U28902 (N_28902,N_22385,N_20965);
nor U28903 (N_28903,N_20629,N_20347);
and U28904 (N_28904,N_24703,N_21975);
or U28905 (N_28905,N_20594,N_21876);
nor U28906 (N_28906,N_24240,N_23154);
or U28907 (N_28907,N_21924,N_24965);
and U28908 (N_28908,N_24700,N_22096);
and U28909 (N_28909,N_20166,N_23056);
nand U28910 (N_28910,N_20713,N_23473);
nand U28911 (N_28911,N_24428,N_24566);
nor U28912 (N_28912,N_21387,N_21755);
or U28913 (N_28913,N_23771,N_23231);
nand U28914 (N_28914,N_22019,N_22376);
and U28915 (N_28915,N_22845,N_24308);
or U28916 (N_28916,N_20462,N_22344);
nand U28917 (N_28917,N_20754,N_24023);
nand U28918 (N_28918,N_20962,N_23965);
nor U28919 (N_28919,N_20024,N_22496);
and U28920 (N_28920,N_20046,N_21002);
nor U28921 (N_28921,N_22856,N_21472);
and U28922 (N_28922,N_21908,N_22625);
nand U28923 (N_28923,N_20760,N_21589);
nor U28924 (N_28924,N_23168,N_24344);
xor U28925 (N_28925,N_20000,N_23787);
nor U28926 (N_28926,N_24499,N_21485);
nand U28927 (N_28927,N_20046,N_20297);
or U28928 (N_28928,N_22113,N_21102);
and U28929 (N_28929,N_24167,N_20196);
or U28930 (N_28930,N_22682,N_21441);
nor U28931 (N_28931,N_24596,N_20274);
or U28932 (N_28932,N_20846,N_23866);
xor U28933 (N_28933,N_20049,N_21873);
nand U28934 (N_28934,N_22339,N_23863);
or U28935 (N_28935,N_21763,N_24824);
or U28936 (N_28936,N_23744,N_22330);
or U28937 (N_28937,N_24200,N_24955);
nand U28938 (N_28938,N_22925,N_21785);
or U28939 (N_28939,N_21661,N_23000);
xor U28940 (N_28940,N_24164,N_22175);
and U28941 (N_28941,N_21947,N_20178);
nand U28942 (N_28942,N_20835,N_21912);
xor U28943 (N_28943,N_22061,N_22714);
or U28944 (N_28944,N_24704,N_20382);
xnor U28945 (N_28945,N_23847,N_20192);
xor U28946 (N_28946,N_20746,N_21995);
and U28947 (N_28947,N_24078,N_24138);
nand U28948 (N_28948,N_22047,N_23120);
and U28949 (N_28949,N_21245,N_24222);
xnor U28950 (N_28950,N_22122,N_21849);
or U28951 (N_28951,N_21528,N_23199);
nand U28952 (N_28952,N_24588,N_22245);
nand U28953 (N_28953,N_23697,N_24593);
and U28954 (N_28954,N_20812,N_21081);
xnor U28955 (N_28955,N_24727,N_20200);
nor U28956 (N_28956,N_20301,N_22504);
or U28957 (N_28957,N_21607,N_23434);
and U28958 (N_28958,N_24154,N_23852);
nor U28959 (N_28959,N_22710,N_21742);
and U28960 (N_28960,N_20401,N_20998);
nand U28961 (N_28961,N_21292,N_22874);
nand U28962 (N_28962,N_20834,N_23168);
nor U28963 (N_28963,N_22566,N_24229);
nand U28964 (N_28964,N_21547,N_24270);
nor U28965 (N_28965,N_20185,N_23450);
nor U28966 (N_28966,N_22672,N_22122);
xor U28967 (N_28967,N_23549,N_24162);
nor U28968 (N_28968,N_21252,N_22336);
nor U28969 (N_28969,N_24449,N_21258);
or U28970 (N_28970,N_24200,N_20190);
xnor U28971 (N_28971,N_23547,N_22925);
nand U28972 (N_28972,N_21302,N_21216);
and U28973 (N_28973,N_24534,N_20854);
and U28974 (N_28974,N_20775,N_23539);
and U28975 (N_28975,N_21145,N_21203);
and U28976 (N_28976,N_22136,N_24661);
and U28977 (N_28977,N_22104,N_21552);
xnor U28978 (N_28978,N_24048,N_21896);
xnor U28979 (N_28979,N_20116,N_23314);
nor U28980 (N_28980,N_20493,N_21675);
nand U28981 (N_28981,N_21554,N_21017);
nand U28982 (N_28982,N_21456,N_22346);
and U28983 (N_28983,N_21634,N_21779);
or U28984 (N_28984,N_24097,N_24555);
or U28985 (N_28985,N_23215,N_24435);
nand U28986 (N_28986,N_22181,N_24964);
nand U28987 (N_28987,N_23703,N_22075);
and U28988 (N_28988,N_23085,N_20842);
or U28989 (N_28989,N_22663,N_22858);
nand U28990 (N_28990,N_22055,N_24782);
and U28991 (N_28991,N_24248,N_23431);
and U28992 (N_28992,N_22601,N_23479);
nor U28993 (N_28993,N_22718,N_24878);
nand U28994 (N_28994,N_23569,N_21122);
and U28995 (N_28995,N_21211,N_21631);
nor U28996 (N_28996,N_21581,N_22756);
and U28997 (N_28997,N_24464,N_22668);
nor U28998 (N_28998,N_22171,N_20851);
and U28999 (N_28999,N_23499,N_20146);
nand U29000 (N_29000,N_23005,N_21767);
nor U29001 (N_29001,N_24061,N_22228);
nor U29002 (N_29002,N_21821,N_21479);
nand U29003 (N_29003,N_21723,N_24931);
or U29004 (N_29004,N_21222,N_22926);
and U29005 (N_29005,N_23300,N_21252);
nor U29006 (N_29006,N_22709,N_23558);
or U29007 (N_29007,N_20476,N_22307);
xnor U29008 (N_29008,N_21552,N_21017);
or U29009 (N_29009,N_22007,N_20167);
or U29010 (N_29010,N_21272,N_23553);
nand U29011 (N_29011,N_24329,N_20420);
and U29012 (N_29012,N_24005,N_23885);
nand U29013 (N_29013,N_23953,N_24700);
or U29014 (N_29014,N_23607,N_20736);
nand U29015 (N_29015,N_22271,N_22856);
nand U29016 (N_29016,N_21780,N_20967);
or U29017 (N_29017,N_20170,N_22684);
nand U29018 (N_29018,N_23146,N_23152);
and U29019 (N_29019,N_24820,N_23538);
or U29020 (N_29020,N_24815,N_23267);
nor U29021 (N_29021,N_21540,N_22017);
nand U29022 (N_29022,N_20800,N_23945);
nand U29023 (N_29023,N_23524,N_21070);
and U29024 (N_29024,N_20975,N_22219);
nand U29025 (N_29025,N_20307,N_20338);
and U29026 (N_29026,N_24816,N_22142);
nand U29027 (N_29027,N_24079,N_20727);
xor U29028 (N_29028,N_21308,N_21079);
nand U29029 (N_29029,N_20926,N_21871);
and U29030 (N_29030,N_24881,N_21020);
or U29031 (N_29031,N_20687,N_24679);
nor U29032 (N_29032,N_20666,N_23692);
nand U29033 (N_29033,N_22664,N_24748);
nor U29034 (N_29034,N_21219,N_24694);
and U29035 (N_29035,N_20041,N_21807);
and U29036 (N_29036,N_20740,N_22778);
xor U29037 (N_29037,N_20091,N_23843);
and U29038 (N_29038,N_22953,N_21742);
nor U29039 (N_29039,N_24859,N_20190);
nor U29040 (N_29040,N_22091,N_24208);
and U29041 (N_29041,N_23279,N_21406);
or U29042 (N_29042,N_23590,N_21522);
or U29043 (N_29043,N_21533,N_22036);
nor U29044 (N_29044,N_21062,N_24264);
or U29045 (N_29045,N_23405,N_21169);
xor U29046 (N_29046,N_20349,N_23148);
nand U29047 (N_29047,N_24272,N_24211);
nand U29048 (N_29048,N_23109,N_20058);
nor U29049 (N_29049,N_21551,N_22275);
nor U29050 (N_29050,N_21843,N_23951);
and U29051 (N_29051,N_22717,N_21064);
nand U29052 (N_29052,N_20011,N_20271);
nor U29053 (N_29053,N_23546,N_23619);
or U29054 (N_29054,N_22282,N_24014);
nor U29055 (N_29055,N_20628,N_21572);
nor U29056 (N_29056,N_24823,N_22185);
nand U29057 (N_29057,N_21824,N_20461);
and U29058 (N_29058,N_20393,N_20918);
xnor U29059 (N_29059,N_20099,N_24518);
and U29060 (N_29060,N_21570,N_21502);
and U29061 (N_29061,N_23719,N_20150);
xnor U29062 (N_29062,N_21492,N_21707);
xnor U29063 (N_29063,N_24927,N_24461);
xnor U29064 (N_29064,N_23284,N_24962);
and U29065 (N_29065,N_24731,N_20447);
nor U29066 (N_29066,N_20030,N_22596);
and U29067 (N_29067,N_22080,N_22913);
or U29068 (N_29068,N_23032,N_24307);
nand U29069 (N_29069,N_21452,N_23125);
nand U29070 (N_29070,N_22826,N_24455);
or U29071 (N_29071,N_22219,N_24213);
or U29072 (N_29072,N_20824,N_24942);
or U29073 (N_29073,N_20808,N_22501);
nand U29074 (N_29074,N_23081,N_20008);
nand U29075 (N_29075,N_20776,N_21207);
xor U29076 (N_29076,N_21596,N_22391);
and U29077 (N_29077,N_21996,N_24633);
nor U29078 (N_29078,N_22584,N_24356);
nand U29079 (N_29079,N_21926,N_24088);
and U29080 (N_29080,N_23624,N_23596);
xnor U29081 (N_29081,N_22694,N_24440);
nor U29082 (N_29082,N_21213,N_20556);
and U29083 (N_29083,N_20602,N_21652);
or U29084 (N_29084,N_23229,N_20430);
xnor U29085 (N_29085,N_22684,N_21551);
or U29086 (N_29086,N_23507,N_21577);
and U29087 (N_29087,N_21740,N_20339);
and U29088 (N_29088,N_24854,N_23691);
or U29089 (N_29089,N_24439,N_21093);
nor U29090 (N_29090,N_22207,N_20351);
or U29091 (N_29091,N_21431,N_20350);
nand U29092 (N_29092,N_21944,N_20551);
nand U29093 (N_29093,N_20367,N_20382);
nor U29094 (N_29094,N_21745,N_23857);
and U29095 (N_29095,N_22615,N_22637);
nand U29096 (N_29096,N_21409,N_24344);
or U29097 (N_29097,N_21310,N_23706);
or U29098 (N_29098,N_24198,N_20414);
and U29099 (N_29099,N_22771,N_22386);
or U29100 (N_29100,N_20490,N_21965);
nor U29101 (N_29101,N_23528,N_20336);
or U29102 (N_29102,N_20782,N_24225);
or U29103 (N_29103,N_24418,N_23089);
or U29104 (N_29104,N_23344,N_21272);
nor U29105 (N_29105,N_24478,N_23034);
xnor U29106 (N_29106,N_20917,N_21444);
or U29107 (N_29107,N_24423,N_22251);
and U29108 (N_29108,N_24764,N_21671);
and U29109 (N_29109,N_24926,N_24640);
nor U29110 (N_29110,N_22643,N_24251);
xor U29111 (N_29111,N_22848,N_22626);
and U29112 (N_29112,N_21052,N_24108);
or U29113 (N_29113,N_22598,N_20507);
nor U29114 (N_29114,N_20861,N_20129);
or U29115 (N_29115,N_21830,N_22144);
nand U29116 (N_29116,N_20491,N_21703);
or U29117 (N_29117,N_24649,N_21663);
nor U29118 (N_29118,N_22166,N_23092);
and U29119 (N_29119,N_22478,N_21433);
nand U29120 (N_29120,N_20424,N_23027);
or U29121 (N_29121,N_21108,N_23273);
nand U29122 (N_29122,N_24527,N_23233);
xor U29123 (N_29123,N_23454,N_21208);
nor U29124 (N_29124,N_24022,N_20881);
nor U29125 (N_29125,N_23414,N_21527);
nand U29126 (N_29126,N_21712,N_24601);
xnor U29127 (N_29127,N_20378,N_21185);
nand U29128 (N_29128,N_20617,N_21288);
nor U29129 (N_29129,N_23509,N_24340);
nand U29130 (N_29130,N_20850,N_23454);
nand U29131 (N_29131,N_22303,N_24112);
nand U29132 (N_29132,N_20207,N_21824);
or U29133 (N_29133,N_24819,N_22653);
nand U29134 (N_29134,N_24283,N_24666);
nand U29135 (N_29135,N_21275,N_24271);
nor U29136 (N_29136,N_20993,N_20630);
xnor U29137 (N_29137,N_23518,N_20334);
or U29138 (N_29138,N_21052,N_21604);
or U29139 (N_29139,N_21523,N_20823);
nor U29140 (N_29140,N_20478,N_22702);
and U29141 (N_29141,N_22752,N_21983);
nor U29142 (N_29142,N_22768,N_21176);
and U29143 (N_29143,N_21007,N_23865);
nor U29144 (N_29144,N_21601,N_24035);
or U29145 (N_29145,N_24757,N_24993);
or U29146 (N_29146,N_21454,N_20773);
nor U29147 (N_29147,N_21820,N_22259);
or U29148 (N_29148,N_24761,N_22975);
or U29149 (N_29149,N_21847,N_22041);
nand U29150 (N_29150,N_21299,N_21385);
nand U29151 (N_29151,N_24172,N_21341);
or U29152 (N_29152,N_21692,N_24528);
and U29153 (N_29153,N_20692,N_20607);
or U29154 (N_29154,N_22140,N_24173);
nor U29155 (N_29155,N_21602,N_24169);
nor U29156 (N_29156,N_20604,N_20325);
xor U29157 (N_29157,N_22570,N_21871);
and U29158 (N_29158,N_24334,N_20298);
or U29159 (N_29159,N_24348,N_22906);
nand U29160 (N_29160,N_22870,N_24256);
and U29161 (N_29161,N_20661,N_20292);
or U29162 (N_29162,N_24852,N_24853);
nand U29163 (N_29163,N_21457,N_21681);
nand U29164 (N_29164,N_24845,N_23249);
nand U29165 (N_29165,N_20736,N_21902);
nand U29166 (N_29166,N_24298,N_23929);
or U29167 (N_29167,N_20099,N_20132);
nor U29168 (N_29168,N_22728,N_21276);
nand U29169 (N_29169,N_20111,N_24720);
or U29170 (N_29170,N_20107,N_22019);
and U29171 (N_29171,N_20278,N_20938);
xor U29172 (N_29172,N_22503,N_23404);
or U29173 (N_29173,N_22154,N_23925);
nand U29174 (N_29174,N_22469,N_24628);
or U29175 (N_29175,N_22314,N_22519);
or U29176 (N_29176,N_23246,N_20431);
nor U29177 (N_29177,N_23942,N_20563);
and U29178 (N_29178,N_23297,N_24248);
xor U29179 (N_29179,N_22956,N_22703);
or U29180 (N_29180,N_24707,N_20635);
nor U29181 (N_29181,N_22838,N_21128);
nor U29182 (N_29182,N_24617,N_23349);
or U29183 (N_29183,N_21030,N_21651);
nand U29184 (N_29184,N_23237,N_23164);
nand U29185 (N_29185,N_22061,N_23274);
or U29186 (N_29186,N_24010,N_22277);
and U29187 (N_29187,N_24828,N_22177);
nand U29188 (N_29188,N_20623,N_23765);
and U29189 (N_29189,N_23240,N_21379);
nand U29190 (N_29190,N_21065,N_21553);
or U29191 (N_29191,N_21812,N_21635);
or U29192 (N_29192,N_22835,N_22431);
or U29193 (N_29193,N_23570,N_21061);
nand U29194 (N_29194,N_21004,N_20978);
and U29195 (N_29195,N_24484,N_22916);
and U29196 (N_29196,N_20847,N_20913);
nand U29197 (N_29197,N_21286,N_21714);
and U29198 (N_29198,N_22179,N_24815);
and U29199 (N_29199,N_24229,N_22762);
and U29200 (N_29200,N_21211,N_20667);
nand U29201 (N_29201,N_22647,N_22105);
xnor U29202 (N_29202,N_20753,N_22079);
nand U29203 (N_29203,N_21837,N_21032);
nand U29204 (N_29204,N_23723,N_21271);
nand U29205 (N_29205,N_24881,N_20016);
nand U29206 (N_29206,N_24372,N_22727);
nand U29207 (N_29207,N_24240,N_21100);
xnor U29208 (N_29208,N_23817,N_22198);
nand U29209 (N_29209,N_22271,N_23614);
and U29210 (N_29210,N_23784,N_21063);
nor U29211 (N_29211,N_24592,N_24472);
nor U29212 (N_29212,N_24259,N_24676);
nor U29213 (N_29213,N_24342,N_22527);
nor U29214 (N_29214,N_22161,N_20463);
nand U29215 (N_29215,N_23551,N_24011);
or U29216 (N_29216,N_23306,N_22712);
and U29217 (N_29217,N_24662,N_20110);
xnor U29218 (N_29218,N_20975,N_20675);
nand U29219 (N_29219,N_21096,N_21810);
xor U29220 (N_29220,N_24351,N_22639);
nand U29221 (N_29221,N_24165,N_24935);
nor U29222 (N_29222,N_22652,N_24782);
xor U29223 (N_29223,N_20102,N_23802);
xor U29224 (N_29224,N_21177,N_22960);
nand U29225 (N_29225,N_24763,N_20096);
nor U29226 (N_29226,N_23060,N_20341);
nand U29227 (N_29227,N_24075,N_20913);
or U29228 (N_29228,N_22842,N_21583);
nor U29229 (N_29229,N_21483,N_24648);
and U29230 (N_29230,N_21819,N_24914);
and U29231 (N_29231,N_23756,N_23134);
nand U29232 (N_29232,N_20488,N_24326);
and U29233 (N_29233,N_22401,N_20279);
and U29234 (N_29234,N_22976,N_23047);
and U29235 (N_29235,N_20551,N_24922);
xor U29236 (N_29236,N_23124,N_20074);
nand U29237 (N_29237,N_21629,N_23361);
nand U29238 (N_29238,N_20614,N_24436);
nand U29239 (N_29239,N_22268,N_21659);
nand U29240 (N_29240,N_20111,N_20376);
or U29241 (N_29241,N_20100,N_22046);
xnor U29242 (N_29242,N_23141,N_24711);
and U29243 (N_29243,N_22385,N_21615);
or U29244 (N_29244,N_21983,N_24243);
and U29245 (N_29245,N_21879,N_24236);
or U29246 (N_29246,N_22109,N_23120);
and U29247 (N_29247,N_23836,N_20858);
nor U29248 (N_29248,N_23511,N_22151);
nor U29249 (N_29249,N_24319,N_22945);
nand U29250 (N_29250,N_23041,N_20836);
xor U29251 (N_29251,N_22867,N_20172);
xor U29252 (N_29252,N_24024,N_22312);
nor U29253 (N_29253,N_22405,N_20256);
or U29254 (N_29254,N_23574,N_23045);
xor U29255 (N_29255,N_23560,N_23064);
nand U29256 (N_29256,N_22073,N_23836);
or U29257 (N_29257,N_24477,N_22512);
and U29258 (N_29258,N_22628,N_20452);
and U29259 (N_29259,N_24413,N_23611);
nor U29260 (N_29260,N_24582,N_21959);
nand U29261 (N_29261,N_21574,N_24752);
xnor U29262 (N_29262,N_22778,N_21084);
xor U29263 (N_29263,N_22701,N_23928);
and U29264 (N_29264,N_20964,N_21230);
or U29265 (N_29265,N_20869,N_20658);
nor U29266 (N_29266,N_22575,N_24187);
and U29267 (N_29267,N_21779,N_22827);
xnor U29268 (N_29268,N_21639,N_21425);
or U29269 (N_29269,N_20931,N_20581);
and U29270 (N_29270,N_22164,N_22122);
nand U29271 (N_29271,N_20716,N_22037);
xor U29272 (N_29272,N_20819,N_21717);
or U29273 (N_29273,N_20697,N_23213);
nand U29274 (N_29274,N_22376,N_20284);
or U29275 (N_29275,N_24507,N_22103);
nor U29276 (N_29276,N_24586,N_20337);
xnor U29277 (N_29277,N_20662,N_23215);
or U29278 (N_29278,N_20082,N_20996);
nor U29279 (N_29279,N_23130,N_23702);
xor U29280 (N_29280,N_20321,N_21451);
and U29281 (N_29281,N_22331,N_20444);
nand U29282 (N_29282,N_23178,N_22278);
nand U29283 (N_29283,N_23821,N_23513);
nor U29284 (N_29284,N_23516,N_21765);
nor U29285 (N_29285,N_24070,N_20488);
xnor U29286 (N_29286,N_22748,N_20184);
nand U29287 (N_29287,N_20448,N_24532);
nand U29288 (N_29288,N_23086,N_20796);
nor U29289 (N_29289,N_23622,N_24650);
nor U29290 (N_29290,N_23216,N_20334);
xnor U29291 (N_29291,N_24277,N_24660);
nor U29292 (N_29292,N_20418,N_24620);
nand U29293 (N_29293,N_22765,N_21794);
nand U29294 (N_29294,N_24840,N_21986);
or U29295 (N_29295,N_24075,N_24556);
nand U29296 (N_29296,N_22746,N_20729);
or U29297 (N_29297,N_21501,N_21984);
nor U29298 (N_29298,N_23470,N_20850);
and U29299 (N_29299,N_24358,N_23600);
or U29300 (N_29300,N_24953,N_22289);
xor U29301 (N_29301,N_22067,N_20174);
nand U29302 (N_29302,N_22284,N_22896);
nand U29303 (N_29303,N_24910,N_24058);
or U29304 (N_29304,N_20483,N_20050);
nand U29305 (N_29305,N_21927,N_23505);
nor U29306 (N_29306,N_24173,N_21584);
xor U29307 (N_29307,N_21448,N_23383);
and U29308 (N_29308,N_24455,N_23809);
nor U29309 (N_29309,N_24484,N_20805);
nor U29310 (N_29310,N_20856,N_21429);
nor U29311 (N_29311,N_23057,N_22233);
and U29312 (N_29312,N_22659,N_20353);
and U29313 (N_29313,N_22849,N_24093);
or U29314 (N_29314,N_22484,N_21048);
or U29315 (N_29315,N_23041,N_20022);
and U29316 (N_29316,N_21252,N_23798);
nand U29317 (N_29317,N_23505,N_24791);
and U29318 (N_29318,N_20832,N_21487);
or U29319 (N_29319,N_22187,N_20750);
nor U29320 (N_29320,N_20189,N_20610);
xor U29321 (N_29321,N_21750,N_24716);
or U29322 (N_29322,N_23949,N_22869);
nor U29323 (N_29323,N_24847,N_23626);
and U29324 (N_29324,N_23517,N_21591);
nor U29325 (N_29325,N_20661,N_21376);
or U29326 (N_29326,N_24454,N_20124);
nand U29327 (N_29327,N_22285,N_21303);
xor U29328 (N_29328,N_20674,N_21708);
or U29329 (N_29329,N_23169,N_21476);
or U29330 (N_29330,N_24700,N_20768);
and U29331 (N_29331,N_20702,N_23114);
or U29332 (N_29332,N_23230,N_22265);
and U29333 (N_29333,N_20854,N_24494);
nor U29334 (N_29334,N_23704,N_24508);
or U29335 (N_29335,N_23932,N_24811);
nand U29336 (N_29336,N_24860,N_20106);
nor U29337 (N_29337,N_21708,N_21885);
or U29338 (N_29338,N_20855,N_23734);
nor U29339 (N_29339,N_23177,N_23835);
nor U29340 (N_29340,N_24843,N_21114);
and U29341 (N_29341,N_22993,N_22651);
or U29342 (N_29342,N_20477,N_22309);
and U29343 (N_29343,N_22763,N_23491);
nand U29344 (N_29344,N_24832,N_24238);
xor U29345 (N_29345,N_24220,N_24842);
nand U29346 (N_29346,N_21938,N_20787);
xor U29347 (N_29347,N_23644,N_21992);
and U29348 (N_29348,N_24970,N_20257);
and U29349 (N_29349,N_23284,N_21980);
nor U29350 (N_29350,N_20401,N_21573);
nor U29351 (N_29351,N_20869,N_24590);
and U29352 (N_29352,N_24202,N_24578);
or U29353 (N_29353,N_24634,N_22416);
or U29354 (N_29354,N_20742,N_23235);
or U29355 (N_29355,N_24619,N_22246);
and U29356 (N_29356,N_22882,N_23877);
or U29357 (N_29357,N_23422,N_20186);
nand U29358 (N_29358,N_20415,N_24973);
xor U29359 (N_29359,N_22030,N_22956);
nor U29360 (N_29360,N_21867,N_20938);
and U29361 (N_29361,N_24827,N_23126);
or U29362 (N_29362,N_22924,N_22647);
and U29363 (N_29363,N_21874,N_24373);
nor U29364 (N_29364,N_20435,N_24441);
nor U29365 (N_29365,N_23583,N_21985);
xor U29366 (N_29366,N_20079,N_22957);
or U29367 (N_29367,N_21684,N_21134);
nand U29368 (N_29368,N_23047,N_24135);
and U29369 (N_29369,N_23694,N_21022);
nand U29370 (N_29370,N_24441,N_23232);
nand U29371 (N_29371,N_20845,N_21153);
or U29372 (N_29372,N_22607,N_20214);
xor U29373 (N_29373,N_24988,N_20441);
nand U29374 (N_29374,N_23377,N_24713);
and U29375 (N_29375,N_20630,N_22786);
xor U29376 (N_29376,N_20218,N_23468);
and U29377 (N_29377,N_22788,N_20177);
or U29378 (N_29378,N_24660,N_24557);
and U29379 (N_29379,N_21429,N_20782);
and U29380 (N_29380,N_24433,N_22075);
xnor U29381 (N_29381,N_22696,N_22638);
or U29382 (N_29382,N_20847,N_24454);
xnor U29383 (N_29383,N_22057,N_21681);
and U29384 (N_29384,N_20529,N_21886);
and U29385 (N_29385,N_23173,N_24168);
and U29386 (N_29386,N_22682,N_24044);
or U29387 (N_29387,N_22269,N_24470);
or U29388 (N_29388,N_24504,N_22662);
and U29389 (N_29389,N_23656,N_20910);
or U29390 (N_29390,N_24829,N_23701);
and U29391 (N_29391,N_22101,N_22765);
nand U29392 (N_29392,N_22485,N_24764);
nor U29393 (N_29393,N_22545,N_21988);
nand U29394 (N_29394,N_22552,N_21971);
and U29395 (N_29395,N_23867,N_21379);
and U29396 (N_29396,N_21919,N_22787);
or U29397 (N_29397,N_20285,N_20063);
xnor U29398 (N_29398,N_22378,N_20546);
and U29399 (N_29399,N_20853,N_20540);
or U29400 (N_29400,N_24394,N_22167);
nand U29401 (N_29401,N_24229,N_21942);
nor U29402 (N_29402,N_20813,N_22685);
nor U29403 (N_29403,N_20923,N_24530);
nand U29404 (N_29404,N_22987,N_23451);
and U29405 (N_29405,N_20324,N_22998);
and U29406 (N_29406,N_22586,N_24023);
and U29407 (N_29407,N_24097,N_22136);
and U29408 (N_29408,N_22112,N_23149);
or U29409 (N_29409,N_20175,N_22711);
or U29410 (N_29410,N_20838,N_20270);
and U29411 (N_29411,N_20084,N_20046);
or U29412 (N_29412,N_20522,N_21021);
and U29413 (N_29413,N_24931,N_23435);
nor U29414 (N_29414,N_24843,N_24280);
and U29415 (N_29415,N_20483,N_20295);
and U29416 (N_29416,N_22443,N_22201);
and U29417 (N_29417,N_21242,N_22562);
and U29418 (N_29418,N_24803,N_21822);
nand U29419 (N_29419,N_21205,N_22530);
nand U29420 (N_29420,N_20524,N_22866);
or U29421 (N_29421,N_24098,N_20023);
and U29422 (N_29422,N_24456,N_24443);
nand U29423 (N_29423,N_22591,N_22291);
and U29424 (N_29424,N_23231,N_23368);
and U29425 (N_29425,N_21844,N_23901);
nor U29426 (N_29426,N_24840,N_21312);
or U29427 (N_29427,N_24250,N_24306);
and U29428 (N_29428,N_23143,N_20028);
nand U29429 (N_29429,N_23046,N_24853);
nand U29430 (N_29430,N_24326,N_21757);
nor U29431 (N_29431,N_23723,N_20282);
xnor U29432 (N_29432,N_24250,N_20111);
nand U29433 (N_29433,N_21470,N_21213);
and U29434 (N_29434,N_20076,N_21435);
nand U29435 (N_29435,N_24603,N_23621);
nand U29436 (N_29436,N_24719,N_23735);
and U29437 (N_29437,N_22798,N_23306);
nor U29438 (N_29438,N_23329,N_21256);
nor U29439 (N_29439,N_21163,N_24004);
nor U29440 (N_29440,N_22921,N_20726);
or U29441 (N_29441,N_23991,N_21571);
nand U29442 (N_29442,N_21483,N_24221);
and U29443 (N_29443,N_21867,N_20022);
nor U29444 (N_29444,N_20972,N_22680);
nor U29445 (N_29445,N_24578,N_24204);
or U29446 (N_29446,N_23475,N_24867);
and U29447 (N_29447,N_23055,N_23956);
nor U29448 (N_29448,N_22782,N_21468);
or U29449 (N_29449,N_20843,N_23137);
and U29450 (N_29450,N_22988,N_22526);
and U29451 (N_29451,N_23392,N_20553);
and U29452 (N_29452,N_23237,N_20880);
nand U29453 (N_29453,N_22248,N_23779);
and U29454 (N_29454,N_24042,N_20742);
nand U29455 (N_29455,N_21393,N_21522);
and U29456 (N_29456,N_23763,N_20938);
nor U29457 (N_29457,N_22658,N_21874);
xor U29458 (N_29458,N_21640,N_22600);
or U29459 (N_29459,N_21258,N_20776);
nor U29460 (N_29460,N_20190,N_22523);
or U29461 (N_29461,N_23408,N_22511);
nand U29462 (N_29462,N_22928,N_21467);
and U29463 (N_29463,N_21154,N_24349);
and U29464 (N_29464,N_24165,N_21170);
or U29465 (N_29465,N_23335,N_21066);
nor U29466 (N_29466,N_21659,N_21490);
or U29467 (N_29467,N_20378,N_20285);
nand U29468 (N_29468,N_20616,N_22022);
and U29469 (N_29469,N_24911,N_21972);
and U29470 (N_29470,N_23559,N_24109);
and U29471 (N_29471,N_20137,N_21861);
or U29472 (N_29472,N_23601,N_20041);
xnor U29473 (N_29473,N_20358,N_24105);
or U29474 (N_29474,N_20501,N_24098);
and U29475 (N_29475,N_24276,N_22654);
nand U29476 (N_29476,N_24298,N_23805);
nand U29477 (N_29477,N_20678,N_23617);
and U29478 (N_29478,N_22369,N_20641);
nand U29479 (N_29479,N_20734,N_22925);
or U29480 (N_29480,N_20563,N_23668);
nand U29481 (N_29481,N_22444,N_21558);
and U29482 (N_29482,N_22330,N_22085);
and U29483 (N_29483,N_24196,N_21955);
and U29484 (N_29484,N_22285,N_20260);
nand U29485 (N_29485,N_22604,N_24292);
or U29486 (N_29486,N_23856,N_23513);
and U29487 (N_29487,N_20211,N_23634);
nand U29488 (N_29488,N_23251,N_22639);
nand U29489 (N_29489,N_20554,N_20340);
nor U29490 (N_29490,N_20884,N_21137);
nand U29491 (N_29491,N_20400,N_21978);
or U29492 (N_29492,N_24896,N_20874);
nor U29493 (N_29493,N_24226,N_20129);
and U29494 (N_29494,N_22214,N_20802);
and U29495 (N_29495,N_24319,N_20674);
nand U29496 (N_29496,N_24618,N_20138);
nand U29497 (N_29497,N_23555,N_23161);
xnor U29498 (N_29498,N_20196,N_20051);
or U29499 (N_29499,N_20239,N_22106);
nor U29500 (N_29500,N_21075,N_21079);
nand U29501 (N_29501,N_21485,N_23096);
nor U29502 (N_29502,N_23561,N_22559);
xnor U29503 (N_29503,N_21112,N_22760);
xnor U29504 (N_29504,N_22339,N_23901);
and U29505 (N_29505,N_24122,N_20211);
and U29506 (N_29506,N_24099,N_20507);
nand U29507 (N_29507,N_24105,N_23304);
and U29508 (N_29508,N_22511,N_21043);
and U29509 (N_29509,N_24225,N_22001);
nor U29510 (N_29510,N_24828,N_22692);
xnor U29511 (N_29511,N_20183,N_20837);
or U29512 (N_29512,N_22223,N_20814);
and U29513 (N_29513,N_21432,N_21951);
xor U29514 (N_29514,N_21370,N_24147);
nor U29515 (N_29515,N_21923,N_22654);
nor U29516 (N_29516,N_24375,N_22866);
nor U29517 (N_29517,N_20375,N_23472);
or U29518 (N_29518,N_24381,N_22760);
nor U29519 (N_29519,N_21432,N_23881);
or U29520 (N_29520,N_20178,N_22761);
nand U29521 (N_29521,N_22192,N_20328);
nor U29522 (N_29522,N_23995,N_21022);
and U29523 (N_29523,N_22277,N_20203);
nor U29524 (N_29524,N_22144,N_23888);
and U29525 (N_29525,N_22720,N_24158);
xnor U29526 (N_29526,N_23727,N_22155);
and U29527 (N_29527,N_22082,N_21636);
nor U29528 (N_29528,N_20845,N_21732);
or U29529 (N_29529,N_21583,N_22962);
and U29530 (N_29530,N_21247,N_21860);
xor U29531 (N_29531,N_22643,N_24683);
or U29532 (N_29532,N_22049,N_22847);
and U29533 (N_29533,N_24224,N_20718);
or U29534 (N_29534,N_20009,N_20559);
nor U29535 (N_29535,N_23512,N_24322);
nor U29536 (N_29536,N_21497,N_20959);
nor U29537 (N_29537,N_24120,N_21313);
and U29538 (N_29538,N_23875,N_21437);
nor U29539 (N_29539,N_20729,N_23161);
and U29540 (N_29540,N_20131,N_20231);
or U29541 (N_29541,N_24331,N_23431);
xnor U29542 (N_29542,N_22054,N_20507);
or U29543 (N_29543,N_23464,N_20765);
nor U29544 (N_29544,N_23847,N_23314);
and U29545 (N_29545,N_21751,N_24844);
nor U29546 (N_29546,N_20463,N_21238);
or U29547 (N_29547,N_24520,N_20003);
nand U29548 (N_29548,N_21013,N_23509);
or U29549 (N_29549,N_20591,N_21993);
nor U29550 (N_29550,N_20055,N_20076);
and U29551 (N_29551,N_22645,N_20756);
nor U29552 (N_29552,N_20203,N_23467);
nand U29553 (N_29553,N_22029,N_22687);
nand U29554 (N_29554,N_22716,N_20548);
or U29555 (N_29555,N_20298,N_22870);
nand U29556 (N_29556,N_24675,N_20872);
xnor U29557 (N_29557,N_23705,N_21120);
nand U29558 (N_29558,N_22319,N_22748);
nand U29559 (N_29559,N_24964,N_20220);
nand U29560 (N_29560,N_20007,N_24101);
and U29561 (N_29561,N_20568,N_21500);
or U29562 (N_29562,N_24274,N_21078);
nor U29563 (N_29563,N_21688,N_23069);
nand U29564 (N_29564,N_23922,N_21828);
xor U29565 (N_29565,N_20804,N_20313);
nor U29566 (N_29566,N_22286,N_23482);
or U29567 (N_29567,N_23847,N_21804);
nand U29568 (N_29568,N_21862,N_23526);
and U29569 (N_29569,N_20599,N_20845);
or U29570 (N_29570,N_22445,N_23000);
nor U29571 (N_29571,N_21972,N_21172);
and U29572 (N_29572,N_21371,N_22378);
and U29573 (N_29573,N_21777,N_21476);
nand U29574 (N_29574,N_23556,N_24974);
nand U29575 (N_29575,N_24726,N_21278);
nand U29576 (N_29576,N_24414,N_20493);
nor U29577 (N_29577,N_24859,N_20578);
xor U29578 (N_29578,N_22136,N_21969);
nor U29579 (N_29579,N_22109,N_21765);
or U29580 (N_29580,N_22215,N_21558);
xor U29581 (N_29581,N_20472,N_22119);
nor U29582 (N_29582,N_22306,N_20102);
xor U29583 (N_29583,N_21929,N_22865);
and U29584 (N_29584,N_21452,N_22473);
nand U29585 (N_29585,N_21179,N_22261);
nand U29586 (N_29586,N_22940,N_22525);
nor U29587 (N_29587,N_23153,N_22300);
nor U29588 (N_29588,N_21416,N_22564);
xnor U29589 (N_29589,N_22085,N_23434);
or U29590 (N_29590,N_20075,N_24737);
nand U29591 (N_29591,N_23283,N_20287);
or U29592 (N_29592,N_24720,N_22022);
xor U29593 (N_29593,N_24485,N_20753);
and U29594 (N_29594,N_23827,N_20623);
nor U29595 (N_29595,N_24758,N_24687);
nand U29596 (N_29596,N_20227,N_24977);
and U29597 (N_29597,N_21958,N_20593);
and U29598 (N_29598,N_23450,N_23449);
and U29599 (N_29599,N_23392,N_23281);
nand U29600 (N_29600,N_23773,N_21060);
nor U29601 (N_29601,N_21543,N_20614);
xnor U29602 (N_29602,N_23674,N_24258);
nor U29603 (N_29603,N_23365,N_22747);
xnor U29604 (N_29604,N_21672,N_22026);
nor U29605 (N_29605,N_21324,N_23034);
or U29606 (N_29606,N_23649,N_20148);
and U29607 (N_29607,N_20755,N_21878);
nand U29608 (N_29608,N_20877,N_22240);
nand U29609 (N_29609,N_24671,N_23970);
or U29610 (N_29610,N_24017,N_24197);
nor U29611 (N_29611,N_20318,N_20712);
nor U29612 (N_29612,N_21392,N_22175);
and U29613 (N_29613,N_20332,N_22669);
nand U29614 (N_29614,N_22428,N_20493);
or U29615 (N_29615,N_24886,N_22575);
nor U29616 (N_29616,N_20609,N_24309);
nor U29617 (N_29617,N_24895,N_21580);
nand U29618 (N_29618,N_23110,N_22304);
or U29619 (N_29619,N_23800,N_22135);
and U29620 (N_29620,N_22128,N_20611);
or U29621 (N_29621,N_22935,N_21937);
nand U29622 (N_29622,N_23983,N_23405);
or U29623 (N_29623,N_22057,N_20634);
nor U29624 (N_29624,N_23460,N_23501);
and U29625 (N_29625,N_23942,N_24385);
and U29626 (N_29626,N_22367,N_23462);
xor U29627 (N_29627,N_20926,N_24543);
or U29628 (N_29628,N_20306,N_24977);
nand U29629 (N_29629,N_21219,N_22746);
or U29630 (N_29630,N_21352,N_23188);
nor U29631 (N_29631,N_21254,N_20542);
nand U29632 (N_29632,N_21188,N_22377);
nand U29633 (N_29633,N_21709,N_23759);
or U29634 (N_29634,N_21993,N_21312);
nand U29635 (N_29635,N_23053,N_23628);
or U29636 (N_29636,N_20825,N_21973);
xor U29637 (N_29637,N_24951,N_23971);
nand U29638 (N_29638,N_20411,N_23887);
or U29639 (N_29639,N_22782,N_20705);
or U29640 (N_29640,N_20316,N_20341);
and U29641 (N_29641,N_24845,N_21367);
and U29642 (N_29642,N_23285,N_23113);
nand U29643 (N_29643,N_20961,N_22361);
and U29644 (N_29644,N_21948,N_23629);
or U29645 (N_29645,N_20873,N_22535);
and U29646 (N_29646,N_23423,N_21060);
nand U29647 (N_29647,N_20939,N_22881);
nor U29648 (N_29648,N_24355,N_24900);
nand U29649 (N_29649,N_22028,N_23388);
or U29650 (N_29650,N_20125,N_21210);
nor U29651 (N_29651,N_23966,N_23704);
nor U29652 (N_29652,N_23832,N_24982);
nor U29653 (N_29653,N_23515,N_21478);
or U29654 (N_29654,N_23126,N_20090);
or U29655 (N_29655,N_21395,N_24541);
xnor U29656 (N_29656,N_21489,N_22955);
or U29657 (N_29657,N_24177,N_23735);
nor U29658 (N_29658,N_20089,N_20439);
nor U29659 (N_29659,N_20996,N_24084);
nor U29660 (N_29660,N_24211,N_20813);
and U29661 (N_29661,N_21342,N_20803);
or U29662 (N_29662,N_24564,N_20450);
and U29663 (N_29663,N_22300,N_20392);
or U29664 (N_29664,N_22453,N_22561);
and U29665 (N_29665,N_24023,N_20640);
and U29666 (N_29666,N_23064,N_23093);
nor U29667 (N_29667,N_20825,N_20330);
nand U29668 (N_29668,N_23760,N_22644);
xor U29669 (N_29669,N_21436,N_23532);
nor U29670 (N_29670,N_21413,N_21703);
or U29671 (N_29671,N_21794,N_23567);
nand U29672 (N_29672,N_22321,N_24597);
nand U29673 (N_29673,N_22957,N_21341);
nor U29674 (N_29674,N_21542,N_22469);
nor U29675 (N_29675,N_23486,N_22820);
nor U29676 (N_29676,N_22305,N_23029);
or U29677 (N_29677,N_22658,N_21120);
or U29678 (N_29678,N_24187,N_23050);
nand U29679 (N_29679,N_24752,N_20383);
or U29680 (N_29680,N_20379,N_24744);
nor U29681 (N_29681,N_21568,N_21955);
nand U29682 (N_29682,N_24471,N_24384);
nor U29683 (N_29683,N_22580,N_24330);
nand U29684 (N_29684,N_22903,N_23493);
xor U29685 (N_29685,N_23628,N_21232);
and U29686 (N_29686,N_21995,N_23995);
xor U29687 (N_29687,N_23022,N_24508);
xor U29688 (N_29688,N_24283,N_24041);
and U29689 (N_29689,N_21866,N_23827);
nand U29690 (N_29690,N_23111,N_20309);
or U29691 (N_29691,N_21273,N_23137);
xor U29692 (N_29692,N_20612,N_21664);
and U29693 (N_29693,N_22309,N_20395);
or U29694 (N_29694,N_23712,N_22292);
nand U29695 (N_29695,N_23640,N_21841);
nor U29696 (N_29696,N_21573,N_21266);
nand U29697 (N_29697,N_23168,N_20245);
nor U29698 (N_29698,N_23952,N_24134);
and U29699 (N_29699,N_20220,N_21667);
nand U29700 (N_29700,N_24264,N_24668);
nor U29701 (N_29701,N_21750,N_20722);
and U29702 (N_29702,N_24177,N_21367);
or U29703 (N_29703,N_21481,N_20891);
nand U29704 (N_29704,N_20183,N_20705);
nand U29705 (N_29705,N_21379,N_23758);
nor U29706 (N_29706,N_20435,N_23078);
or U29707 (N_29707,N_24223,N_20518);
nor U29708 (N_29708,N_23569,N_21970);
nor U29709 (N_29709,N_20861,N_21525);
nor U29710 (N_29710,N_23910,N_22521);
and U29711 (N_29711,N_22633,N_22520);
and U29712 (N_29712,N_22057,N_24237);
nor U29713 (N_29713,N_24667,N_24669);
nor U29714 (N_29714,N_20989,N_23678);
nor U29715 (N_29715,N_23444,N_21949);
or U29716 (N_29716,N_20656,N_23521);
or U29717 (N_29717,N_20286,N_20068);
nor U29718 (N_29718,N_21965,N_22845);
nor U29719 (N_29719,N_22742,N_23791);
nand U29720 (N_29720,N_24360,N_22197);
xor U29721 (N_29721,N_20923,N_20943);
nor U29722 (N_29722,N_21484,N_23647);
nor U29723 (N_29723,N_23994,N_24540);
nor U29724 (N_29724,N_24987,N_20878);
nand U29725 (N_29725,N_20693,N_20837);
nor U29726 (N_29726,N_22792,N_23395);
nand U29727 (N_29727,N_24738,N_24249);
and U29728 (N_29728,N_21754,N_23484);
or U29729 (N_29729,N_20899,N_22806);
or U29730 (N_29730,N_21233,N_20788);
or U29731 (N_29731,N_20747,N_22363);
and U29732 (N_29732,N_24285,N_22858);
nor U29733 (N_29733,N_24815,N_24883);
and U29734 (N_29734,N_21459,N_20482);
or U29735 (N_29735,N_23051,N_24689);
nand U29736 (N_29736,N_24730,N_24719);
and U29737 (N_29737,N_23926,N_23668);
xor U29738 (N_29738,N_22796,N_22447);
or U29739 (N_29739,N_21292,N_23731);
nand U29740 (N_29740,N_23782,N_23605);
or U29741 (N_29741,N_20684,N_22013);
nor U29742 (N_29742,N_20052,N_22157);
nor U29743 (N_29743,N_21101,N_23383);
nand U29744 (N_29744,N_24845,N_23008);
nor U29745 (N_29745,N_21747,N_22064);
nor U29746 (N_29746,N_20558,N_23813);
or U29747 (N_29747,N_24013,N_20969);
and U29748 (N_29748,N_22709,N_22310);
nand U29749 (N_29749,N_20245,N_22787);
nand U29750 (N_29750,N_21706,N_23862);
or U29751 (N_29751,N_23752,N_21238);
nand U29752 (N_29752,N_23076,N_24953);
and U29753 (N_29753,N_20006,N_21726);
nor U29754 (N_29754,N_22174,N_21210);
or U29755 (N_29755,N_23314,N_21833);
or U29756 (N_29756,N_22814,N_23255);
nor U29757 (N_29757,N_24295,N_20205);
or U29758 (N_29758,N_23449,N_21962);
and U29759 (N_29759,N_22099,N_21271);
nor U29760 (N_29760,N_24113,N_20100);
and U29761 (N_29761,N_21256,N_22763);
xor U29762 (N_29762,N_24951,N_24767);
nand U29763 (N_29763,N_22898,N_23856);
nand U29764 (N_29764,N_23265,N_23957);
nand U29765 (N_29765,N_21445,N_23730);
xor U29766 (N_29766,N_20241,N_20700);
nand U29767 (N_29767,N_22751,N_21952);
nor U29768 (N_29768,N_21747,N_24483);
nand U29769 (N_29769,N_20037,N_21220);
nor U29770 (N_29770,N_24114,N_20132);
xnor U29771 (N_29771,N_20931,N_21453);
or U29772 (N_29772,N_24788,N_22901);
nor U29773 (N_29773,N_22970,N_24127);
and U29774 (N_29774,N_23854,N_21661);
nor U29775 (N_29775,N_21489,N_23988);
and U29776 (N_29776,N_24671,N_21426);
nand U29777 (N_29777,N_21328,N_22872);
nand U29778 (N_29778,N_20256,N_21971);
xnor U29779 (N_29779,N_24075,N_24379);
or U29780 (N_29780,N_21704,N_23835);
nor U29781 (N_29781,N_22166,N_24553);
and U29782 (N_29782,N_22219,N_22552);
or U29783 (N_29783,N_23748,N_20579);
nand U29784 (N_29784,N_21891,N_23486);
and U29785 (N_29785,N_20147,N_23529);
and U29786 (N_29786,N_24303,N_23179);
nor U29787 (N_29787,N_23054,N_24601);
and U29788 (N_29788,N_21496,N_22819);
and U29789 (N_29789,N_22858,N_20423);
nand U29790 (N_29790,N_21896,N_21238);
or U29791 (N_29791,N_24136,N_22372);
xor U29792 (N_29792,N_22128,N_24169);
or U29793 (N_29793,N_21067,N_20082);
xnor U29794 (N_29794,N_20721,N_24896);
nand U29795 (N_29795,N_23218,N_22369);
and U29796 (N_29796,N_22555,N_24052);
nand U29797 (N_29797,N_20625,N_24812);
nor U29798 (N_29798,N_23369,N_23463);
and U29799 (N_29799,N_21860,N_21669);
and U29800 (N_29800,N_24323,N_22995);
xnor U29801 (N_29801,N_21419,N_24728);
xnor U29802 (N_29802,N_23790,N_20336);
nand U29803 (N_29803,N_20544,N_24226);
and U29804 (N_29804,N_20655,N_20195);
xor U29805 (N_29805,N_20532,N_21521);
nor U29806 (N_29806,N_20239,N_23128);
and U29807 (N_29807,N_24100,N_22247);
or U29808 (N_29808,N_22274,N_23525);
nand U29809 (N_29809,N_23705,N_23902);
and U29810 (N_29810,N_21649,N_23255);
or U29811 (N_29811,N_22272,N_21382);
and U29812 (N_29812,N_21780,N_21103);
and U29813 (N_29813,N_21501,N_24302);
or U29814 (N_29814,N_23433,N_21053);
nor U29815 (N_29815,N_24166,N_24046);
and U29816 (N_29816,N_24254,N_21857);
and U29817 (N_29817,N_22892,N_21512);
and U29818 (N_29818,N_23241,N_23606);
and U29819 (N_29819,N_21353,N_24909);
nor U29820 (N_29820,N_23979,N_21334);
and U29821 (N_29821,N_24782,N_22965);
nand U29822 (N_29822,N_21675,N_20955);
nand U29823 (N_29823,N_24302,N_24616);
nand U29824 (N_29824,N_24102,N_24670);
or U29825 (N_29825,N_22644,N_21229);
or U29826 (N_29826,N_22334,N_21942);
or U29827 (N_29827,N_22135,N_23003);
xnor U29828 (N_29828,N_23746,N_22166);
nor U29829 (N_29829,N_23686,N_21698);
and U29830 (N_29830,N_23871,N_20833);
or U29831 (N_29831,N_21127,N_23137);
nor U29832 (N_29832,N_23438,N_21185);
and U29833 (N_29833,N_24725,N_24727);
nor U29834 (N_29834,N_24551,N_20792);
nor U29835 (N_29835,N_24345,N_23715);
and U29836 (N_29836,N_23721,N_20626);
nor U29837 (N_29837,N_22895,N_24097);
xor U29838 (N_29838,N_21780,N_20392);
nand U29839 (N_29839,N_22008,N_21135);
xnor U29840 (N_29840,N_22583,N_20026);
or U29841 (N_29841,N_23864,N_21455);
nand U29842 (N_29842,N_22569,N_24191);
xnor U29843 (N_29843,N_24746,N_21379);
or U29844 (N_29844,N_24158,N_21570);
xnor U29845 (N_29845,N_24747,N_21721);
nor U29846 (N_29846,N_24130,N_23393);
and U29847 (N_29847,N_23148,N_21333);
and U29848 (N_29848,N_23359,N_22624);
nand U29849 (N_29849,N_20748,N_23027);
and U29850 (N_29850,N_21695,N_21269);
xor U29851 (N_29851,N_21249,N_20909);
xor U29852 (N_29852,N_21231,N_20122);
xor U29853 (N_29853,N_23626,N_24854);
and U29854 (N_29854,N_22062,N_21700);
and U29855 (N_29855,N_22460,N_23669);
nor U29856 (N_29856,N_24842,N_24073);
or U29857 (N_29857,N_24309,N_24199);
or U29858 (N_29858,N_21774,N_23377);
nor U29859 (N_29859,N_24052,N_20641);
nand U29860 (N_29860,N_24958,N_21185);
nand U29861 (N_29861,N_21041,N_22382);
and U29862 (N_29862,N_21205,N_23239);
and U29863 (N_29863,N_21644,N_21042);
nor U29864 (N_29864,N_23323,N_24597);
nand U29865 (N_29865,N_20665,N_20453);
or U29866 (N_29866,N_23533,N_23797);
nand U29867 (N_29867,N_22581,N_24590);
and U29868 (N_29868,N_21833,N_21841);
xnor U29869 (N_29869,N_22450,N_20386);
nand U29870 (N_29870,N_22195,N_20201);
and U29871 (N_29871,N_24861,N_20207);
or U29872 (N_29872,N_20459,N_20061);
nand U29873 (N_29873,N_20486,N_21972);
xor U29874 (N_29874,N_22621,N_22723);
and U29875 (N_29875,N_20557,N_21421);
and U29876 (N_29876,N_20146,N_22902);
or U29877 (N_29877,N_21320,N_24409);
nor U29878 (N_29878,N_22975,N_20719);
or U29879 (N_29879,N_22609,N_22817);
and U29880 (N_29880,N_23963,N_24154);
nand U29881 (N_29881,N_24117,N_24907);
and U29882 (N_29882,N_20593,N_21557);
and U29883 (N_29883,N_22659,N_23000);
nor U29884 (N_29884,N_22969,N_22613);
nand U29885 (N_29885,N_24897,N_24136);
or U29886 (N_29886,N_24274,N_24615);
nand U29887 (N_29887,N_20780,N_23929);
and U29888 (N_29888,N_23828,N_24724);
xor U29889 (N_29889,N_20812,N_20122);
nand U29890 (N_29890,N_20150,N_22848);
nand U29891 (N_29891,N_22575,N_22781);
nor U29892 (N_29892,N_20549,N_20238);
nand U29893 (N_29893,N_24690,N_21119);
nor U29894 (N_29894,N_24448,N_22605);
nor U29895 (N_29895,N_23415,N_20701);
nand U29896 (N_29896,N_22406,N_22442);
or U29897 (N_29897,N_22497,N_20479);
xnor U29898 (N_29898,N_24075,N_22215);
xnor U29899 (N_29899,N_20270,N_22234);
nor U29900 (N_29900,N_24062,N_20130);
and U29901 (N_29901,N_20646,N_23029);
nor U29902 (N_29902,N_24489,N_20167);
nor U29903 (N_29903,N_23393,N_21215);
xor U29904 (N_29904,N_24061,N_20753);
and U29905 (N_29905,N_23931,N_21300);
or U29906 (N_29906,N_23340,N_24411);
xnor U29907 (N_29907,N_23465,N_22139);
or U29908 (N_29908,N_23099,N_21932);
or U29909 (N_29909,N_21097,N_21840);
or U29910 (N_29910,N_21804,N_21984);
xor U29911 (N_29911,N_24399,N_24002);
and U29912 (N_29912,N_23464,N_22323);
and U29913 (N_29913,N_21051,N_20165);
and U29914 (N_29914,N_24985,N_23654);
nand U29915 (N_29915,N_21337,N_20661);
nor U29916 (N_29916,N_24691,N_21575);
or U29917 (N_29917,N_23630,N_24318);
nor U29918 (N_29918,N_22412,N_22340);
and U29919 (N_29919,N_23033,N_24305);
nand U29920 (N_29920,N_23110,N_22544);
nand U29921 (N_29921,N_20629,N_23190);
and U29922 (N_29922,N_23181,N_20938);
and U29923 (N_29923,N_22398,N_22870);
and U29924 (N_29924,N_24173,N_24976);
nor U29925 (N_29925,N_22205,N_23369);
nand U29926 (N_29926,N_24784,N_22922);
or U29927 (N_29927,N_21746,N_22693);
and U29928 (N_29928,N_24332,N_22107);
nor U29929 (N_29929,N_21981,N_24991);
nand U29930 (N_29930,N_24132,N_23101);
nand U29931 (N_29931,N_24514,N_23577);
nor U29932 (N_29932,N_23940,N_20494);
or U29933 (N_29933,N_21700,N_20146);
or U29934 (N_29934,N_22121,N_21552);
nand U29935 (N_29935,N_22594,N_20815);
and U29936 (N_29936,N_22912,N_23254);
or U29937 (N_29937,N_21727,N_20581);
nor U29938 (N_29938,N_22410,N_22626);
nand U29939 (N_29939,N_23468,N_20480);
and U29940 (N_29940,N_24794,N_21463);
nand U29941 (N_29941,N_20186,N_22150);
or U29942 (N_29942,N_21183,N_23308);
nor U29943 (N_29943,N_23876,N_24099);
or U29944 (N_29944,N_24928,N_20730);
nor U29945 (N_29945,N_24999,N_20180);
and U29946 (N_29946,N_20639,N_21470);
nor U29947 (N_29947,N_21966,N_21445);
nor U29948 (N_29948,N_24048,N_21693);
xor U29949 (N_29949,N_20015,N_21451);
nand U29950 (N_29950,N_21789,N_20140);
nand U29951 (N_29951,N_21268,N_24389);
nor U29952 (N_29952,N_20109,N_21258);
nand U29953 (N_29953,N_22400,N_23059);
nand U29954 (N_29954,N_22316,N_21754);
or U29955 (N_29955,N_21440,N_24144);
nor U29956 (N_29956,N_24898,N_20311);
nor U29957 (N_29957,N_20241,N_24366);
nor U29958 (N_29958,N_23335,N_22407);
nand U29959 (N_29959,N_22085,N_21071);
or U29960 (N_29960,N_20851,N_21740);
nor U29961 (N_29961,N_24064,N_23759);
nor U29962 (N_29962,N_20527,N_22526);
and U29963 (N_29963,N_23497,N_22065);
and U29964 (N_29964,N_21901,N_21974);
and U29965 (N_29965,N_21021,N_24196);
nor U29966 (N_29966,N_23639,N_24622);
nor U29967 (N_29967,N_20117,N_23397);
or U29968 (N_29968,N_20104,N_22341);
nand U29969 (N_29969,N_20996,N_24509);
or U29970 (N_29970,N_23541,N_24686);
or U29971 (N_29971,N_21613,N_21692);
nand U29972 (N_29972,N_20248,N_22571);
or U29973 (N_29973,N_24276,N_22073);
or U29974 (N_29974,N_24424,N_23427);
nor U29975 (N_29975,N_22131,N_21093);
or U29976 (N_29976,N_22357,N_20783);
and U29977 (N_29977,N_23366,N_22508);
or U29978 (N_29978,N_22223,N_24832);
xnor U29979 (N_29979,N_24976,N_22925);
and U29980 (N_29980,N_20539,N_22205);
nor U29981 (N_29981,N_20454,N_20576);
xor U29982 (N_29982,N_24110,N_23584);
and U29983 (N_29983,N_23994,N_22805);
nor U29984 (N_29984,N_21211,N_21360);
or U29985 (N_29985,N_20616,N_24384);
and U29986 (N_29986,N_22778,N_24741);
or U29987 (N_29987,N_24530,N_22112);
xnor U29988 (N_29988,N_20393,N_22662);
and U29989 (N_29989,N_24051,N_24233);
nor U29990 (N_29990,N_22389,N_22799);
nor U29991 (N_29991,N_24638,N_21047);
or U29992 (N_29992,N_20166,N_23396);
nand U29993 (N_29993,N_24902,N_20936);
or U29994 (N_29994,N_21246,N_20048);
nand U29995 (N_29995,N_21235,N_22551);
nand U29996 (N_29996,N_24112,N_21382);
or U29997 (N_29997,N_23250,N_20500);
and U29998 (N_29998,N_20443,N_23498);
xnor U29999 (N_29999,N_20839,N_21986);
and UO_0 (O_0,N_26201,N_26163);
nor UO_1 (O_1,N_29921,N_29655);
nor UO_2 (O_2,N_26513,N_27667);
nor UO_3 (O_3,N_29057,N_26859);
nand UO_4 (O_4,N_26339,N_25692);
or UO_5 (O_5,N_26943,N_28604);
and UO_6 (O_6,N_29618,N_27137);
and UO_7 (O_7,N_28900,N_28983);
or UO_8 (O_8,N_26349,N_25171);
nor UO_9 (O_9,N_28741,N_28307);
and UO_10 (O_10,N_25518,N_29547);
nor UO_11 (O_11,N_29546,N_25765);
nor UO_12 (O_12,N_28205,N_26614);
nand UO_13 (O_13,N_26505,N_28776);
xor UO_14 (O_14,N_25013,N_26952);
or UO_15 (O_15,N_25343,N_25564);
and UO_16 (O_16,N_27682,N_28171);
or UO_17 (O_17,N_26200,N_27767);
or UO_18 (O_18,N_29550,N_29661);
and UO_19 (O_19,N_27449,N_28317);
nor UO_20 (O_20,N_25122,N_25687);
or UO_21 (O_21,N_27694,N_25834);
or UO_22 (O_22,N_27648,N_27198);
or UO_23 (O_23,N_25408,N_25238);
nand UO_24 (O_24,N_29089,N_25295);
and UO_25 (O_25,N_27446,N_29024);
xor UO_26 (O_26,N_27023,N_28860);
nor UO_27 (O_27,N_28611,N_27974);
xnor UO_28 (O_28,N_25086,N_27164);
or UO_29 (O_29,N_26500,N_25534);
nand UO_30 (O_30,N_26192,N_27812);
nor UO_31 (O_31,N_26093,N_26292);
nand UO_32 (O_32,N_27459,N_27235);
nor UO_33 (O_33,N_29568,N_27064);
or UO_34 (O_34,N_28754,N_27129);
nand UO_35 (O_35,N_27157,N_26341);
nand UO_36 (O_36,N_28898,N_27580);
and UO_37 (O_37,N_26627,N_26363);
xnor UO_38 (O_38,N_27708,N_27621);
and UO_39 (O_39,N_27674,N_29253);
nor UO_40 (O_40,N_25414,N_25293);
nand UO_41 (O_41,N_26127,N_25395);
and UO_42 (O_42,N_25315,N_28400);
xnor UO_43 (O_43,N_25341,N_25451);
nor UO_44 (O_44,N_29318,N_25832);
and UO_45 (O_45,N_27758,N_26951);
nand UO_46 (O_46,N_29572,N_25389);
nand UO_47 (O_47,N_26174,N_26609);
and UO_48 (O_48,N_26631,N_28661);
xor UO_49 (O_49,N_27300,N_25225);
nand UO_50 (O_50,N_26262,N_29076);
nor UO_51 (O_51,N_25527,N_28113);
nand UO_52 (O_52,N_27709,N_29218);
xnor UO_53 (O_53,N_25557,N_28727);
nand UO_54 (O_54,N_29874,N_27835);
or UO_55 (O_55,N_27640,N_28214);
nor UO_56 (O_56,N_27221,N_29890);
and UO_57 (O_57,N_29879,N_25284);
nor UO_58 (O_58,N_25397,N_26249);
nand UO_59 (O_59,N_29946,N_25049);
xor UO_60 (O_60,N_25226,N_28642);
or UO_61 (O_61,N_25491,N_26670);
nand UO_62 (O_62,N_29490,N_27509);
xnor UO_63 (O_63,N_26877,N_26465);
nand UO_64 (O_64,N_28079,N_25673);
or UO_65 (O_65,N_25465,N_29381);
or UO_66 (O_66,N_25381,N_26424);
or UO_67 (O_67,N_26265,N_26849);
and UO_68 (O_68,N_29138,N_29088);
nand UO_69 (O_69,N_28685,N_29978);
and UO_70 (O_70,N_27199,N_27266);
and UO_71 (O_71,N_25066,N_27833);
and UO_72 (O_72,N_27942,N_26980);
or UO_73 (O_73,N_27894,N_28034);
and UO_74 (O_74,N_25883,N_27042);
nand UO_75 (O_75,N_27697,N_26421);
nor UO_76 (O_76,N_27093,N_27739);
and UO_77 (O_77,N_28092,N_25936);
and UO_78 (O_78,N_27555,N_28529);
xor UO_79 (O_79,N_27900,N_25870);
nand UO_80 (O_80,N_26153,N_28259);
nor UO_81 (O_81,N_27774,N_28279);
nand UO_82 (O_82,N_29472,N_29231);
or UO_83 (O_83,N_26824,N_27190);
or UO_84 (O_84,N_28890,N_27022);
or UO_85 (O_85,N_27991,N_28610);
and UO_86 (O_86,N_26625,N_25143);
or UO_87 (O_87,N_26018,N_28624);
or UO_88 (O_88,N_26662,N_27314);
and UO_89 (O_89,N_28510,N_26460);
and UO_90 (O_90,N_29329,N_27663);
and UO_91 (O_91,N_28668,N_25023);
or UO_92 (O_92,N_27250,N_26255);
nor UO_93 (O_93,N_28028,N_29344);
and UO_94 (O_94,N_29308,N_25710);
or UO_95 (O_95,N_27360,N_26385);
nand UO_96 (O_96,N_27258,N_28915);
xor UO_97 (O_97,N_28519,N_28176);
and UO_98 (O_98,N_28740,N_29540);
nor UO_99 (O_99,N_25046,N_25730);
and UO_100 (O_100,N_28858,N_26468);
nor UO_101 (O_101,N_28375,N_25747);
nor UO_102 (O_102,N_25633,N_29241);
nor UO_103 (O_103,N_27996,N_26253);
and UO_104 (O_104,N_25379,N_29722);
and UO_105 (O_105,N_25098,N_28138);
xnor UO_106 (O_106,N_26914,N_29098);
nand UO_107 (O_107,N_25110,N_25075);
nand UO_108 (O_108,N_25691,N_26629);
nand UO_109 (O_109,N_25327,N_25124);
nand UO_110 (O_110,N_25555,N_27229);
and UO_111 (O_111,N_28587,N_25458);
nand UO_112 (O_112,N_25189,N_28350);
nand UO_113 (O_113,N_27576,N_28304);
nor UO_114 (O_114,N_29534,N_28326);
and UO_115 (O_115,N_29450,N_26739);
or UO_116 (O_116,N_27055,N_25173);
xnor UO_117 (O_117,N_28190,N_25240);
nor UO_118 (O_118,N_29934,N_27245);
and UO_119 (O_119,N_29559,N_26068);
or UO_120 (O_120,N_25971,N_28826);
nor UO_121 (O_121,N_27813,N_27294);
and UO_122 (O_122,N_25647,N_27471);
or UO_123 (O_123,N_26263,N_29852);
and UO_124 (O_124,N_29336,N_27223);
and UO_125 (O_125,N_26960,N_26526);
or UO_126 (O_126,N_27210,N_29999);
nand UO_127 (O_127,N_29525,N_25019);
or UO_128 (O_128,N_25498,N_29268);
nor UO_129 (O_129,N_25210,N_25749);
nor UO_130 (O_130,N_27106,N_28179);
and UO_131 (O_131,N_28870,N_29826);
nand UO_132 (O_132,N_26872,N_27751);
or UO_133 (O_133,N_28369,N_25289);
nand UO_134 (O_134,N_25776,N_29147);
nand UO_135 (O_135,N_26359,N_28756);
and UO_136 (O_136,N_29654,N_26748);
nor UO_137 (O_137,N_29959,N_25619);
nor UO_138 (O_138,N_29407,N_25551);
nor UO_139 (O_139,N_25968,N_29338);
nand UO_140 (O_140,N_26125,N_29632);
and UO_141 (O_141,N_27066,N_29944);
xor UO_142 (O_142,N_26126,N_26475);
nand UO_143 (O_143,N_26308,N_29576);
nor UO_144 (O_144,N_29793,N_27565);
nand UO_145 (O_145,N_29090,N_28647);
or UO_146 (O_146,N_28622,N_29666);
or UO_147 (O_147,N_27853,N_28000);
nor UO_148 (O_148,N_29393,N_29447);
or UO_149 (O_149,N_27881,N_29755);
and UO_150 (O_150,N_25490,N_29504);
or UO_151 (O_151,N_29283,N_26531);
or UO_152 (O_152,N_29264,N_25431);
xnor UO_153 (O_153,N_29179,N_29692);
nand UO_154 (O_154,N_27582,N_27799);
xnor UO_155 (O_155,N_26556,N_25304);
nor UO_156 (O_156,N_25552,N_28427);
nor UO_157 (O_157,N_25157,N_26242);
nor UO_158 (O_158,N_28527,N_25184);
nand UO_159 (O_159,N_29561,N_25073);
nor UO_160 (O_160,N_26793,N_25665);
nor UO_161 (O_161,N_27347,N_29465);
or UO_162 (O_162,N_28110,N_28973);
nand UO_163 (O_163,N_29911,N_27743);
and UO_164 (O_164,N_28100,N_27716);
xnor UO_165 (O_165,N_26254,N_26621);
nand UO_166 (O_166,N_27242,N_25837);
and UO_167 (O_167,N_28729,N_27930);
and UO_168 (O_168,N_29462,N_25982);
xnor UO_169 (O_169,N_28571,N_28008);
or UO_170 (O_170,N_26876,N_26347);
or UO_171 (O_171,N_29769,N_28193);
and UO_172 (O_172,N_28447,N_25858);
xor UO_173 (O_173,N_27656,N_25700);
nand UO_174 (O_174,N_27399,N_28812);
and UO_175 (O_175,N_29323,N_29097);
nor UO_176 (O_176,N_26733,N_29920);
nor UO_177 (O_177,N_26170,N_27626);
or UO_178 (O_178,N_27348,N_26903);
and UO_179 (O_179,N_25215,N_26796);
and UO_180 (O_180,N_27172,N_28974);
and UO_181 (O_181,N_27989,N_28507);
and UO_182 (O_182,N_29259,N_28908);
and UO_183 (O_183,N_27069,N_26161);
nand UO_184 (O_184,N_27939,N_26769);
xnor UO_185 (O_185,N_28015,N_29758);
or UO_186 (O_186,N_27834,N_26854);
nor UO_187 (O_187,N_26141,N_25689);
and UO_188 (O_188,N_25648,N_25152);
or UO_189 (O_189,N_27549,N_26470);
and UO_190 (O_190,N_26867,N_26709);
nand UO_191 (O_191,N_26934,N_29896);
nand UO_192 (O_192,N_25093,N_29485);
and UO_193 (O_193,N_26528,N_26319);
nand UO_194 (O_194,N_26365,N_29935);
nor UO_195 (O_195,N_29172,N_26384);
and UO_196 (O_196,N_26821,N_29951);
or UO_197 (O_197,N_27283,N_27091);
and UO_198 (O_198,N_29481,N_29244);
nand UO_199 (O_199,N_26819,N_26996);
or UO_200 (O_200,N_29892,N_26097);
or UO_201 (O_201,N_27062,N_29137);
xor UO_202 (O_202,N_26399,N_28448);
xor UO_203 (O_203,N_25282,N_28545);
and UO_204 (O_204,N_28584,N_29840);
nor UO_205 (O_205,N_28497,N_25961);
nor UO_206 (O_206,N_28819,N_27869);
or UO_207 (O_207,N_29558,N_25867);
xor UO_208 (O_208,N_29022,N_29217);
and UO_209 (O_209,N_26922,N_26166);
or UO_210 (O_210,N_26033,N_27008);
nor UO_211 (O_211,N_27529,N_29782);
or UO_212 (O_212,N_26437,N_26218);
nor UO_213 (O_213,N_25434,N_29280);
and UO_214 (O_214,N_29120,N_29523);
nand UO_215 (O_215,N_29206,N_25108);
nand UO_216 (O_216,N_25768,N_27722);
nand UO_217 (O_217,N_25789,N_29304);
nand UO_218 (O_218,N_27264,N_26527);
nand UO_219 (O_219,N_26239,N_29479);
nor UO_220 (O_220,N_25997,N_27720);
nand UO_221 (O_221,N_28710,N_25892);
nand UO_222 (O_222,N_27601,N_26603);
nand UO_223 (O_223,N_25781,N_27849);
xor UO_224 (O_224,N_25898,N_29423);
xor UO_225 (O_225,N_25622,N_28280);
or UO_226 (O_226,N_27354,N_28737);
nand UO_227 (O_227,N_27249,N_25056);
and UO_228 (O_228,N_28335,N_27121);
or UO_229 (O_229,N_28802,N_27019);
and UO_230 (O_230,N_26155,N_29190);
nor UO_231 (O_231,N_29684,N_26016);
or UO_232 (O_232,N_26521,N_27005);
xnor UO_233 (O_233,N_28431,N_28846);
and UO_234 (O_234,N_26969,N_26569);
nor UO_235 (O_235,N_26507,N_26970);
and UO_236 (O_236,N_25271,N_28018);
and UO_237 (O_237,N_29464,N_27263);
nor UO_238 (O_238,N_28355,N_27158);
nor UO_239 (O_239,N_29819,N_25478);
and UO_240 (O_240,N_26535,N_28155);
xor UO_241 (O_241,N_28924,N_28440);
and UO_242 (O_242,N_27434,N_25055);
xnor UO_243 (O_243,N_26401,N_26508);
nor UO_244 (O_244,N_28765,N_26790);
xor UO_245 (O_245,N_29274,N_27961);
nor UO_246 (O_246,N_29605,N_28650);
xor UO_247 (O_247,N_27362,N_25720);
nand UO_248 (O_248,N_28017,N_26599);
or UO_249 (O_249,N_27032,N_29453);
nor UO_250 (O_250,N_28251,N_27034);
nand UO_251 (O_251,N_25370,N_26655);
or UO_252 (O_252,N_26873,N_28743);
nor UO_253 (O_253,N_29792,N_25766);
nor UO_254 (O_254,N_25894,N_25112);
or UO_255 (O_255,N_25872,N_27824);
nand UO_256 (O_256,N_28823,N_27843);
nand UO_257 (O_257,N_29480,N_25485);
nand UO_258 (O_258,N_29201,N_25664);
and UO_259 (O_259,N_25609,N_25231);
nand UO_260 (O_260,N_29502,N_26457);
and UO_261 (O_261,N_27937,N_29562);
or UO_262 (O_262,N_27504,N_29298);
and UO_263 (O_263,N_26855,N_27292);
or UO_264 (O_264,N_27233,N_28559);
and UO_265 (O_265,N_26687,N_27220);
nor UO_266 (O_266,N_26910,N_29067);
nor UO_267 (O_267,N_25167,N_25348);
and UO_268 (O_268,N_27015,N_25909);
nand UO_269 (O_269,N_25076,N_29560);
nor UO_270 (O_270,N_29055,N_25918);
or UO_271 (O_271,N_28137,N_28364);
nor UO_272 (O_272,N_25421,N_26813);
or UO_273 (O_273,N_26717,N_27173);
or UO_274 (O_274,N_25649,N_26644);
or UO_275 (O_275,N_26443,N_28365);
nor UO_276 (O_276,N_27252,N_25260);
and UO_277 (O_277,N_28594,N_27257);
or UO_278 (O_278,N_25702,N_25081);
nand UO_279 (O_279,N_26622,N_26946);
nor UO_280 (O_280,N_27593,N_27317);
nand UO_281 (O_281,N_26888,N_27809);
and UO_282 (O_282,N_28945,N_25705);
or UO_283 (O_283,N_28867,N_27128);
and UO_284 (O_284,N_26327,N_28778);
nor UO_285 (O_285,N_28630,N_29730);
and UO_286 (O_286,N_25965,N_26520);
or UO_287 (O_287,N_28827,N_27451);
xor UO_288 (O_288,N_29918,N_29455);
nor UO_289 (O_289,N_29282,N_27867);
xnor UO_290 (O_290,N_28725,N_28485);
nor UO_291 (O_291,N_27478,N_26752);
and UO_292 (O_292,N_28608,N_26967);
and UO_293 (O_293,N_27563,N_27759);
or UO_294 (O_294,N_28912,N_27038);
or UO_295 (O_295,N_26591,N_29810);
nand UO_296 (O_296,N_26912,N_29907);
or UO_297 (O_297,N_27613,N_29733);
and UO_298 (O_298,N_29419,N_27048);
nand UO_299 (O_299,N_28123,N_25694);
nand UO_300 (O_300,N_25668,N_29924);
or UO_301 (O_301,N_28881,N_28060);
nand UO_302 (O_302,N_29037,N_29783);
nand UO_303 (O_303,N_25636,N_25342);
nor UO_304 (O_304,N_28136,N_28578);
nor UO_305 (O_305,N_25109,N_28759);
and UO_306 (O_306,N_27929,N_28050);
or UO_307 (O_307,N_25088,N_28486);
xor UO_308 (O_308,N_28324,N_26495);
and UO_309 (O_309,N_27778,N_29477);
or UO_310 (O_310,N_28960,N_29746);
and UO_311 (O_311,N_29590,N_27234);
nand UO_312 (O_312,N_25077,N_29357);
nand UO_313 (O_313,N_26745,N_25548);
nor UO_314 (O_314,N_26302,N_27384);
nor UO_315 (O_315,N_25751,N_27714);
xnor UO_316 (O_316,N_25712,N_29588);
xor UO_317 (O_317,N_26073,N_27395);
nor UO_318 (O_318,N_25933,N_26881);
nand UO_319 (O_319,N_27819,N_28520);
nor UO_320 (O_320,N_27790,N_28139);
nor UO_321 (O_321,N_27311,N_28201);
xor UO_322 (O_322,N_28583,N_25848);
nor UO_323 (O_323,N_27369,N_27203);
xnor UO_324 (O_324,N_25535,N_29048);
and UO_325 (O_325,N_28892,N_29273);
and UO_326 (O_326,N_29953,N_27830);
nor UO_327 (O_327,N_27113,N_28690);
nor UO_328 (O_328,N_29327,N_25369);
and UO_329 (O_329,N_27423,N_27359);
nor UO_330 (O_330,N_26393,N_27897);
and UO_331 (O_331,N_28184,N_29994);
or UO_332 (O_332,N_28374,N_29262);
nor UO_333 (O_333,N_26856,N_25446);
and UO_334 (O_334,N_28683,N_29272);
nor UO_335 (O_335,N_29131,N_27782);
nand UO_336 (O_336,N_25537,N_29254);
nor UO_337 (O_337,N_25409,N_26270);
nand UO_338 (O_338,N_25262,N_29598);
xnor UO_339 (O_339,N_26012,N_25158);
xor UO_340 (O_340,N_27548,N_28321);
xor UO_341 (O_341,N_27006,N_27046);
xnor UO_342 (O_342,N_28805,N_29569);
nor UO_343 (O_343,N_26235,N_26410);
xor UO_344 (O_344,N_27176,N_29404);
nor UO_345 (O_345,N_25992,N_29230);
and UO_346 (O_346,N_27126,N_27461);
xor UO_347 (O_347,N_25041,N_26886);
and UO_348 (O_348,N_29864,N_29827);
and UO_349 (O_349,N_25213,N_25674);
and UO_350 (O_350,N_25233,N_26378);
or UO_351 (O_351,N_28186,N_29341);
xnor UO_352 (O_352,N_26459,N_29250);
xnor UO_353 (O_353,N_27142,N_25764);
xor UO_354 (O_354,N_25711,N_29965);
and UO_355 (O_355,N_27707,N_28884);
nand UO_356 (O_356,N_27094,N_25516);
xor UO_357 (O_357,N_29938,N_25686);
xnor UO_358 (O_358,N_28733,N_26369);
and UO_359 (O_359,N_25021,N_28435);
nand UO_360 (O_360,N_26822,N_25254);
and UO_361 (O_361,N_28874,N_26286);
xor UO_362 (O_362,N_29467,N_27202);
and UO_363 (O_363,N_27842,N_25525);
nor UO_364 (O_364,N_29612,N_28401);
or UO_365 (O_365,N_26909,N_25347);
nor UO_366 (O_366,N_28348,N_28336);
and UO_367 (O_367,N_26798,N_26023);
and UO_368 (O_368,N_25107,N_29331);
nand UO_369 (O_369,N_26742,N_27789);
or UO_370 (O_370,N_28426,N_29156);
nor UO_371 (O_371,N_27584,N_29884);
or UO_372 (O_372,N_25773,N_25955);
or UO_373 (O_373,N_26534,N_26466);
and UO_374 (O_374,N_25199,N_27765);
xor UO_375 (O_375,N_28966,N_29609);
and UO_376 (O_376,N_27412,N_27999);
nand UO_377 (O_377,N_27905,N_25371);
and UO_378 (O_378,N_25921,N_27185);
nor UO_379 (O_379,N_27306,N_28885);
or UO_380 (O_380,N_27702,N_27779);
nand UO_381 (O_381,N_26323,N_25573);
nor UO_382 (O_382,N_27717,N_28523);
or UO_383 (O_383,N_27839,N_25726);
nand UO_384 (O_384,N_27891,N_26635);
nand UO_385 (O_385,N_26522,N_28086);
nor UO_386 (O_386,N_27057,N_28202);
nor UO_387 (O_387,N_28031,N_28552);
nor UO_388 (O_388,N_28981,N_26005);
or UO_389 (O_389,N_27297,N_26212);
nor UO_390 (O_390,N_28976,N_29159);
nor UO_391 (O_391,N_28509,N_25453);
and UO_392 (O_392,N_26791,N_29977);
nor UO_393 (O_393,N_25817,N_29683);
or UO_394 (O_394,N_29996,N_26060);
and UO_395 (O_395,N_28859,N_27002);
or UO_396 (O_396,N_29084,N_25117);
or UO_397 (O_397,N_27180,N_29132);
nor UO_398 (O_398,N_25136,N_29092);
or UO_399 (O_399,N_25078,N_28875);
or UO_400 (O_400,N_25303,N_26202);
or UO_401 (O_401,N_27770,N_25952);
or UO_402 (O_402,N_28029,N_27868);
nor UO_403 (O_403,N_28800,N_27856);
nor UO_404 (O_404,N_25162,N_29705);
nor UO_405 (O_405,N_27545,N_28775);
xnor UO_406 (O_406,N_28325,N_26087);
and UO_407 (O_407,N_29050,N_27847);
nand UO_408 (O_408,N_25266,N_29768);
and UO_409 (O_409,N_28215,N_29489);
or UO_410 (O_410,N_28476,N_28586);
or UO_411 (O_411,N_28402,N_25441);
and UO_412 (O_412,N_27322,N_25068);
nor UO_413 (O_413,N_28234,N_26990);
xor UO_414 (O_414,N_29675,N_29780);
nor UO_415 (O_415,N_27017,N_29038);
or UO_416 (O_416,N_28806,N_27662);
or UO_417 (O_417,N_28418,N_28063);
and UO_418 (O_418,N_29202,N_27916);
and UO_419 (O_419,N_27159,N_28542);
or UO_420 (O_420,N_28699,N_25051);
and UO_421 (O_421,N_29509,N_27453);
or UO_422 (O_422,N_28061,N_29858);
nand UO_423 (O_423,N_27913,N_28739);
nor UO_424 (O_424,N_26774,N_29957);
or UO_425 (O_425,N_27726,N_27806);
xor UO_426 (O_426,N_29972,N_26780);
nor UO_427 (O_427,N_29971,N_27296);
and UO_428 (O_428,N_25950,N_28393);
nor UO_429 (O_429,N_26035,N_26289);
or UO_430 (O_430,N_29514,N_27704);
and UO_431 (O_431,N_28276,N_26560);
or UO_432 (O_432,N_29401,N_29856);
xnor UO_433 (O_433,N_29051,N_27538);
nand UO_434 (O_434,N_26448,N_25227);
xor UO_435 (O_435,N_26371,N_28302);
or UO_436 (O_436,N_26808,N_28799);
nor UO_437 (O_437,N_27882,N_26593);
nand UO_438 (O_438,N_27239,N_28300);
nor UO_439 (O_439,N_28457,N_28169);
nand UO_440 (O_440,N_28016,N_27950);
nand UO_441 (O_441,N_29045,N_25026);
or UO_442 (O_442,N_29281,N_27775);
and UO_443 (O_443,N_25835,N_28045);
nand UO_444 (O_444,N_29784,N_25194);
nand UO_445 (O_445,N_25376,N_26129);
and UO_446 (O_446,N_26493,N_25926);
nand UO_447 (O_447,N_25312,N_29163);
nor UO_448 (O_448,N_26483,N_26340);
or UO_449 (O_449,N_27418,N_28600);
or UO_450 (O_450,N_27401,N_27166);
or UO_451 (O_451,N_29518,N_29503);
xnor UO_452 (O_452,N_28346,N_28597);
nor UO_453 (O_453,N_28682,N_25324);
nor UO_454 (O_454,N_25630,N_26017);
nor UO_455 (O_455,N_25216,N_26149);
and UO_456 (O_456,N_25533,N_27293);
and UO_457 (O_457,N_25917,N_25799);
and UO_458 (O_458,N_25111,N_28617);
nor UO_459 (O_459,N_25187,N_29725);
and UO_460 (O_460,N_28894,N_28697);
xor UO_461 (O_461,N_26831,N_26285);
xnor UO_462 (O_462,N_28226,N_27192);
or UO_463 (O_463,N_25221,N_28387);
or UO_464 (O_464,N_25559,N_29321);
nor UO_465 (O_465,N_28704,N_29302);
or UO_466 (O_466,N_25940,N_28413);
nor UO_467 (O_467,N_25344,N_25599);
nand UO_468 (O_468,N_26740,N_25653);
nand UO_469 (O_469,N_28004,N_28992);
or UO_470 (O_470,N_29984,N_26266);
and UO_471 (O_471,N_28388,N_29804);
nand UO_472 (O_472,N_28453,N_27865);
and UO_473 (O_473,N_25724,N_29717);
or UO_474 (O_474,N_27797,N_29277);
nand UO_475 (O_475,N_28764,N_26386);
and UO_476 (O_476,N_28428,N_28511);
xnor UO_477 (O_477,N_26875,N_25214);
and UO_478 (O_478,N_27490,N_27328);
nor UO_479 (O_479,N_26545,N_25200);
or UO_480 (O_480,N_25806,N_28582);
xor UO_481 (O_481,N_27163,N_26217);
xnor UO_482 (O_482,N_28189,N_29410);
nand UO_483 (O_483,N_29071,N_26968);
nor UO_484 (O_484,N_26864,N_26203);
nand UO_485 (O_485,N_29350,N_25703);
or UO_486 (O_486,N_26431,N_25605);
nand UO_487 (O_487,N_28373,N_26427);
xnor UO_488 (O_488,N_26688,N_26778);
nor UO_489 (O_489,N_27928,N_28020);
nand UO_490 (O_490,N_28910,N_29563);
nor UO_491 (O_491,N_28021,N_29983);
nand UO_492 (O_492,N_26305,N_27200);
or UO_493 (O_493,N_26057,N_29434);
and UO_494 (O_494,N_29516,N_29492);
and UO_495 (O_495,N_25241,N_26866);
or UO_496 (O_496,N_29413,N_27193);
xnor UO_497 (O_497,N_26324,N_25887);
xor UO_498 (O_498,N_26123,N_25246);
and UO_499 (O_499,N_27056,N_28546);
and UO_500 (O_500,N_27893,N_25586);
or UO_501 (O_501,N_28012,N_27725);
nand UO_502 (O_502,N_28558,N_29813);
nand UO_503 (O_503,N_27895,N_29375);
nand UO_504 (O_504,N_28356,N_26337);
nand UO_505 (O_505,N_28999,N_26314);
and UO_506 (O_506,N_25652,N_25641);
and UO_507 (O_507,N_29814,N_26026);
nand UO_508 (O_508,N_27195,N_25774);
and UO_509 (O_509,N_25357,N_26729);
or UO_510 (O_510,N_28352,N_28262);
and UO_511 (O_511,N_26134,N_29161);
nor UO_512 (O_512,N_25025,N_28475);
nor UO_513 (O_513,N_29881,N_25886);
or UO_514 (O_514,N_27781,N_29351);
nand UO_515 (O_515,N_27124,N_26422);
nand UO_516 (O_516,N_26247,N_26165);
or UO_517 (O_517,N_25772,N_27493);
or UO_518 (O_518,N_25864,N_28389);
or UO_519 (O_519,N_27814,N_25283);
nor UO_520 (O_520,N_27552,N_25280);
nor UO_521 (O_521,N_27099,N_29243);
nand UO_522 (O_522,N_29236,N_25275);
nor UO_523 (O_523,N_29880,N_25778);
nand UO_524 (O_524,N_25583,N_26027);
or UO_525 (O_525,N_26426,N_25882);
and UO_526 (O_526,N_26160,N_27816);
nand UO_527 (O_527,N_27026,N_28577);
or UO_528 (O_528,N_27037,N_29680);
or UO_529 (O_529,N_29859,N_26634);
or UO_530 (O_530,N_25662,N_29976);
nand UO_531 (O_531,N_25356,N_26021);
and UO_532 (O_532,N_29371,N_26956);
nand UO_533 (O_533,N_27922,N_27303);
and UO_534 (O_534,N_26312,N_27456);
nand UO_535 (O_535,N_28358,N_28105);
or UO_536 (O_536,N_26084,N_26974);
xnor UO_537 (O_537,N_25368,N_27411);
nand UO_538 (O_538,N_26015,N_25511);
and UO_539 (O_539,N_29279,N_29893);
nand UO_540 (O_540,N_25337,N_28657);
and UO_541 (O_541,N_27599,N_26279);
nor UO_542 (O_542,N_26233,N_28522);
and UO_543 (O_543,N_27579,N_27815);
nor UO_544 (O_544,N_25713,N_25290);
and UO_545 (O_545,N_25203,N_28643);
or UO_546 (O_546,N_29541,N_26984);
and UO_547 (O_547,N_29069,N_27416);
nor UO_548 (O_548,N_27277,N_26678);
nand UO_549 (O_549,N_25980,N_26906);
and UO_550 (O_550,N_29903,N_25219);
and UO_551 (O_551,N_28614,N_29638);
nor UO_552 (O_552,N_29713,N_29760);
or UO_553 (O_553,N_27209,N_27109);
and UO_554 (O_554,N_25330,N_25580);
nor UO_555 (O_555,N_26751,N_28667);
nand UO_556 (O_556,N_25180,N_27885);
and UO_557 (O_557,N_25310,N_29335);
xnor UO_558 (O_558,N_27736,N_26804);
nand UO_559 (O_559,N_28926,N_29307);
nand UO_560 (O_560,N_26848,N_26389);
and UO_561 (O_561,N_28244,N_25292);
and UO_562 (O_562,N_28718,N_28693);
xor UO_563 (O_563,N_29672,N_29724);
and UO_564 (O_564,N_28196,N_28026);
nor UO_565 (O_565,N_29975,N_28728);
nor UO_566 (O_566,N_26382,N_27054);
nor UO_567 (O_567,N_26897,N_29296);
xor UO_568 (O_568,N_29685,N_29807);
nor UO_569 (O_569,N_29284,N_29016);
nor UO_570 (O_570,N_27361,N_27608);
and UO_571 (O_571,N_25927,N_25838);
or UO_572 (O_572,N_27492,N_29747);
and UO_573 (O_573,N_25553,N_29942);
or UO_574 (O_574,N_25951,N_28853);
or UO_575 (O_575,N_28556,N_26691);
or UO_576 (O_576,N_28856,N_26425);
nor UO_577 (O_577,N_27612,N_28591);
and UO_578 (O_578,N_25496,N_29260);
nand UO_579 (O_579,N_29630,N_26182);
nand UO_580 (O_580,N_28731,N_25727);
nand UO_581 (O_581,N_28318,N_29449);
xor UO_582 (O_582,N_29029,N_29991);
nor UO_583 (O_583,N_27838,N_28386);
nor UO_584 (O_584,N_25069,N_26904);
or UO_585 (O_585,N_28633,N_27946);
or UO_586 (O_586,N_29442,N_27721);
nor UO_587 (O_587,N_25494,N_27216);
and UO_588 (O_588,N_29738,N_27562);
nand UO_589 (O_589,N_25132,N_29396);
and UO_590 (O_590,N_26588,N_28461);
nand UO_591 (O_591,N_26638,N_29266);
nand UO_592 (O_592,N_25582,N_28815);
xnor UO_593 (O_593,N_25539,N_29099);
or UO_594 (O_594,N_29548,N_27116);
or UO_595 (O_595,N_28277,N_27494);
nor UO_596 (O_596,N_26089,N_28851);
or UO_597 (O_597,N_27696,N_25515);
or UO_598 (O_598,N_27706,N_27050);
or UO_599 (O_599,N_25159,N_27899);
and UO_600 (O_600,N_27324,N_27547);
nor UO_601 (O_601,N_28069,N_25018);
xnor UO_602 (O_602,N_25106,N_28157);
xor UO_603 (O_603,N_26771,N_25182);
or UO_604 (O_604,N_27407,N_29036);
xor UO_605 (O_605,N_28688,N_27191);
and UO_606 (O_606,N_26447,N_25758);
or UO_607 (O_607,N_29967,N_29712);
and UO_608 (O_608,N_29860,N_27327);
or UO_609 (O_609,N_29299,N_27826);
nand UO_610 (O_610,N_29468,N_25212);
and UO_611 (O_611,N_28705,N_25074);
or UO_612 (O_612,N_29042,N_25201);
or UO_613 (O_613,N_28811,N_28637);
xnor UO_614 (O_614,N_28271,N_28786);
nor UO_615 (O_615,N_28084,N_28390);
xnor UO_616 (O_616,N_28872,N_29301);
and UO_617 (O_617,N_29194,N_25393);
and UO_618 (O_618,N_25061,N_26541);
and UO_619 (O_619,N_26490,N_26602);
and UO_620 (O_620,N_27020,N_27858);
xnor UO_621 (O_621,N_29107,N_28439);
and UO_622 (O_622,N_27052,N_27860);
xnor UO_623 (O_623,N_29604,N_28167);
xnor UO_624 (O_624,N_28782,N_25188);
or UO_625 (O_625,N_25775,N_25745);
nor UO_626 (O_626,N_27321,N_28087);
nand UO_627 (O_627,N_28404,N_28187);
nand UO_628 (O_628,N_28175,N_29948);
nand UO_629 (O_629,N_27307,N_29316);
or UO_630 (O_630,N_29932,N_25874);
nand UO_631 (O_631,N_28726,N_29429);
nor UO_632 (O_632,N_29762,N_28033);
and UO_633 (O_633,N_28297,N_29033);
nand UO_634 (O_634,N_25660,N_29227);
and UO_635 (O_635,N_25737,N_28014);
or UO_636 (O_636,N_27043,N_27151);
or UO_637 (O_637,N_29438,N_28059);
nor UO_638 (O_638,N_25697,N_29828);
nor UO_639 (O_639,N_28396,N_25611);
and UO_640 (O_640,N_28677,N_27155);
and UO_641 (O_641,N_26845,N_27941);
nand UO_642 (O_642,N_28467,N_26164);
xnor UO_643 (O_643,N_27330,N_29440);
xor UO_644 (O_644,N_28022,N_29674);
and UO_645 (O_645,N_29818,N_29352);
and UO_646 (O_646,N_26226,N_29652);
nand UO_647 (O_647,N_28531,N_28755);
xnor UO_648 (O_648,N_26862,N_28770);
or UO_649 (O_649,N_28882,N_26954);
or UO_650 (O_650,N_29524,N_25354);
nand UO_651 (O_651,N_25466,N_28935);
and UO_652 (O_652,N_25486,N_28504);
nor UO_653 (O_653,N_25090,N_27733);
nand UO_654 (O_654,N_26981,N_25116);
and UO_655 (O_655,N_25010,N_29265);
nor UO_656 (O_656,N_29641,N_26908);
and UO_657 (O_657,N_29809,N_25708);
nor UO_658 (O_658,N_29745,N_29741);
nor UO_659 (O_659,N_27440,N_27425);
nand UO_660 (O_660,N_26797,N_26962);
nor UO_661 (O_661,N_27866,N_27926);
and UO_662 (O_662,N_29169,N_25916);
xnor UO_663 (O_663,N_26045,N_26643);
or UO_664 (O_664,N_28342,N_26991);
nand UO_665 (O_665,N_25364,N_29646);
nand UO_666 (O_666,N_25941,N_25272);
or UO_667 (O_667,N_27127,N_27345);
and UO_668 (O_668,N_29153,N_29181);
nor UO_669 (O_669,N_28085,N_26111);
and UO_670 (O_670,N_26171,N_25362);
and UO_671 (O_671,N_28385,N_25318);
and UO_672 (O_672,N_27460,N_29643);
and UO_673 (O_673,N_26313,N_25914);
nand UO_674 (O_674,N_26293,N_27089);
nor UO_675 (O_675,N_27165,N_29074);
nor UO_676 (O_676,N_29586,N_28267);
nor UO_677 (O_677,N_25651,N_28818);
nand UO_678 (O_678,N_29034,N_27730);
xnor UO_679 (O_679,N_26597,N_29322);
nand UO_680 (O_680,N_25547,N_26451);
nor UO_681 (O_681,N_28188,N_25541);
and UO_682 (O_682,N_26509,N_26479);
nand UO_683 (O_683,N_29451,N_25334);
nor UO_684 (O_684,N_29386,N_28744);
or UO_685 (O_685,N_28181,N_27956);
nor UO_686 (O_686,N_29732,N_28229);
nor UO_687 (O_687,N_25889,N_28292);
and UO_688 (O_688,N_25170,N_26842);
or UO_689 (O_689,N_28857,N_26186);
and UO_690 (O_690,N_28148,N_29862);
or UO_691 (O_691,N_27935,N_25001);
nor UO_692 (O_692,N_27875,N_26277);
nand UO_693 (O_693,N_26557,N_27540);
nand UO_694 (O_694,N_29075,N_27243);
or UO_695 (O_695,N_28395,N_25263);
or UO_696 (O_696,N_27740,N_26179);
nor UO_697 (O_697,N_28248,N_27325);
nand UO_698 (O_698,N_27161,N_27557);
nand UO_699 (O_699,N_29119,N_29941);
nor UO_700 (O_700,N_28253,N_25037);
nand UO_701 (O_701,N_28944,N_27138);
nand UO_702 (O_702,N_25234,N_26002);
and UO_703 (O_703,N_27665,N_29554);
or UO_704 (O_704,N_27188,N_26777);
nor UO_705 (O_705,N_29461,N_26231);
and UO_706 (O_706,N_27993,N_27658);
nand UO_707 (O_707,N_29936,N_26439);
nand UO_708 (O_708,N_26190,N_29000);
nor UO_709 (O_709,N_25612,N_25603);
or UO_710 (O_710,N_29209,N_26983);
nor UO_711 (O_711,N_29167,N_27452);
and UO_712 (O_712,N_26659,N_25197);
nor UO_713 (O_713,N_26899,N_26360);
nand UO_714 (O_714,N_29821,N_29662);
nand UO_715 (O_715,N_28824,N_27445);
nor UO_716 (O_716,N_28601,N_26350);
or UO_717 (O_717,N_29542,N_29584);
nor UO_718 (O_718,N_28686,N_29059);
nand UO_719 (O_719,N_26563,N_29671);
and UO_720 (O_720,N_27871,N_28096);
nand UO_721 (O_721,N_25976,N_29297);
xor UO_722 (O_722,N_26196,N_26374);
nor UO_723 (O_723,N_29011,N_25558);
and UO_724 (O_724,N_25281,N_26379);
or UO_725 (O_725,N_29791,N_25487);
nand UO_726 (O_726,N_26768,N_27598);
and UO_727 (O_727,N_27021,N_29126);
or UO_728 (O_728,N_26574,N_29046);
or UO_729 (O_729,N_27238,N_25340);
nor UO_730 (O_730,N_29372,N_29535);
and UO_731 (O_731,N_27585,N_29992);
or UO_732 (O_732,N_29007,N_25699);
or UO_733 (O_733,N_29943,N_25499);
or UO_734 (O_734,N_28141,N_27473);
nand UO_735 (O_735,N_28788,N_29019);
or UO_736 (O_736,N_26444,N_29904);
nor UO_737 (O_737,N_29114,N_25034);
and UO_738 (O_738,N_25524,N_25877);
and UO_739 (O_739,N_28019,N_29578);
and UO_740 (O_740,N_27502,N_26518);
nand UO_741 (O_741,N_26616,N_26434);
or UO_742 (O_742,N_26388,N_29412);
xor UO_743 (O_743,N_27821,N_29645);
nand UO_744 (O_744,N_28410,N_28191);
or UO_745 (O_745,N_27684,N_26803);
xor UO_746 (O_746,N_28261,N_26608);
nor UO_747 (O_747,N_29956,N_25995);
nor UO_748 (O_748,N_26400,N_25947);
or UO_749 (O_749,N_28047,N_26536);
or UO_750 (O_750,N_26753,N_26334);
or UO_751 (O_751,N_29557,N_26920);
or UO_752 (O_752,N_25690,N_25420);
and UO_753 (O_753,N_28866,N_26637);
nand UO_754 (O_754,N_29543,N_27918);
or UO_755 (O_755,N_27532,N_29647);
nand UO_756 (O_756,N_28422,N_28801);
nand UO_757 (O_757,N_26006,N_28088);
and UO_758 (O_758,N_29734,N_28282);
or UO_759 (O_759,N_29580,N_27679);
nor UO_760 (O_760,N_29473,N_28498);
nor UO_761 (O_761,N_27332,N_29778);
xor UO_762 (O_762,N_26636,N_27783);
nor UO_763 (O_763,N_27764,N_29018);
nor UO_764 (O_764,N_28508,N_28967);
and UO_765 (O_765,N_25601,N_28821);
and UO_766 (O_766,N_29032,N_26979);
nor UO_767 (O_767,N_25148,N_28549);
and UO_768 (O_768,N_26940,N_26222);
or UO_769 (O_769,N_25814,N_27344);
and UO_770 (O_770,N_29233,N_27448);
and UO_771 (O_771,N_28102,N_27854);
nand UO_772 (O_772,N_29798,N_25160);
nand UO_773 (O_773,N_26352,N_25503);
and UO_774 (O_774,N_29197,N_28257);
nand UO_775 (O_775,N_29628,N_26724);
nor UO_776 (O_776,N_29512,N_27168);
nor UO_777 (O_777,N_29141,N_29927);
nor UO_778 (O_778,N_26046,N_27086);
nor UO_779 (O_779,N_26686,N_27108);
nand UO_780 (O_780,N_25053,N_28090);
xor UO_781 (O_781,N_26834,N_25970);
and UO_782 (O_782,N_28715,N_29855);
nand UO_783 (O_783,N_28753,N_25418);
xor UO_784 (O_784,N_26972,N_28499);
or UO_785 (O_785,N_25352,N_28108);
and UO_786 (O_786,N_29597,N_29182);
or UO_787 (O_787,N_25492,N_26482);
and UO_788 (O_788,N_28991,N_29753);
and UO_789 (O_789,N_29801,N_28200);
and UO_790 (O_790,N_26442,N_29969);
or UO_791 (O_791,N_26646,N_28289);
and UO_792 (O_792,N_29116,N_25363);
nor UO_793 (O_793,N_27212,N_27983);
and UO_794 (O_794,N_26999,N_27503);
xnor UO_795 (O_795,N_27267,N_27525);
nand UO_796 (O_796,N_29754,N_28627);
and UO_797 (O_797,N_27218,N_29409);
nor UO_798 (O_798,N_25593,N_26604);
and UO_799 (O_799,N_25050,N_27995);
or UO_800 (O_800,N_28524,N_27031);
nand UO_801 (O_801,N_26278,N_25688);
or UO_802 (O_802,N_28848,N_26098);
xnor UO_803 (O_803,N_28816,N_27417);
nand UO_804 (O_804,N_28091,N_26478);
nor UO_805 (O_805,N_27256,N_29135);
nor UO_806 (O_806,N_29010,N_25884);
nand UO_807 (O_807,N_29506,N_29234);
nand UO_808 (O_808,N_26446,N_25899);
nor UO_809 (O_809,N_28918,N_29706);
nand UO_810 (O_810,N_28331,N_28834);
nor UO_811 (O_811,N_29817,N_26645);
and UO_812 (O_812,N_29292,N_27510);
or UO_813 (O_813,N_26503,N_29415);
nand UO_814 (O_814,N_26827,N_26596);
or UO_815 (O_815,N_29545,N_29749);
nand UO_816 (O_816,N_28540,N_27769);
nand UO_817 (O_817,N_25323,N_29897);
nor UO_818 (O_818,N_27947,N_29475);
nand UO_819 (O_819,N_28180,N_28252);
and UO_820 (O_820,N_29627,N_26851);
nand UO_821 (O_821,N_26491,N_26765);
xor UO_822 (O_822,N_26533,N_26680);
xnor UO_823 (O_823,N_29248,N_25788);
nand UO_824 (O_824,N_29536,N_28536);
xor UO_825 (O_825,N_28897,N_27701);
or UO_826 (O_826,N_26607,N_26932);
nand UO_827 (O_827,N_26215,N_28496);
nand UO_828 (O_828,N_25752,N_25991);
xor UO_829 (O_829,N_25901,N_27206);
and UO_830 (O_830,N_29278,N_28409);
nand UO_831 (O_831,N_28011,N_26871);
nand UO_832 (O_832,N_25928,N_28576);
or UO_833 (O_833,N_27495,N_26061);
nand UO_834 (O_834,N_27241,N_26759);
and UO_835 (O_835,N_28362,N_26880);
nand UO_836 (O_836,N_29223,N_26373);
nand UO_837 (O_837,N_28825,N_28424);
xor UO_838 (O_838,N_25896,N_28417);
and UO_839 (O_839,N_29017,N_25291);
or UO_840 (O_840,N_27972,N_26965);
xnor UO_841 (O_841,N_29624,N_28695);
nand UO_842 (O_842,N_28236,N_26586);
or UO_843 (O_843,N_25484,N_29993);
and UO_844 (O_844,N_26896,N_25591);
xnor UO_845 (O_845,N_29295,N_27025);
and UO_846 (O_846,N_28414,N_27068);
nor UO_847 (O_847,N_25632,N_25429);
or UO_848 (O_848,N_26036,N_28165);
xor UO_849 (O_849,N_27376,N_27352);
nand UO_850 (O_850,N_27776,N_26072);
and UO_851 (O_851,N_28493,N_27215);
nand UO_852 (O_852,N_25588,N_28354);
xnor UO_853 (O_853,N_28140,N_26100);
or UO_854 (O_854,N_29751,N_26076);
or UO_855 (O_855,N_28379,N_27786);
and UO_856 (O_856,N_28284,N_27831);
xnor UO_857 (O_857,N_29796,N_28246);
and UO_858 (O_858,N_25404,N_26624);
nand UO_859 (O_859,N_27275,N_29836);
and UO_860 (O_860,N_27825,N_25607);
nor UO_861 (O_861,N_25501,N_26694);
nor UO_862 (O_862,N_29251,N_29395);
xnor UO_863 (O_863,N_27840,N_27270);
xor UO_864 (O_864,N_25011,N_29072);
nand UO_865 (O_865,N_28796,N_27623);
nor UO_866 (O_866,N_29602,N_26939);
or UO_867 (O_867,N_25461,N_25335);
nand UO_868 (O_868,N_28748,N_28199);
nor UO_869 (O_869,N_27810,N_26814);
xor UO_870 (O_870,N_29533,N_29521);
nor UO_871 (O_871,N_29103,N_27546);
nand UO_872 (O_872,N_29637,N_28076);
nor UO_873 (O_873,N_28405,N_28423);
nor UO_874 (O_874,N_27260,N_26601);
nor UO_875 (O_875,N_29228,N_27225);
and UO_876 (O_876,N_25036,N_29361);
and UO_877 (O_877,N_26014,N_28221);
xnor UO_878 (O_878,N_29701,N_28674);
xor UO_879 (O_879,N_25089,N_25902);
nor UO_880 (O_880,N_28436,N_29484);
nand UO_881 (O_881,N_26720,N_26390);
nor UO_882 (O_882,N_27368,N_28330);
xor UO_883 (O_883,N_28114,N_28691);
or UO_884 (O_884,N_28049,N_28367);
nor UO_885 (O_885,N_29154,N_26976);
and UO_886 (O_886,N_29592,N_29513);
nand UO_887 (O_887,N_29648,N_25684);
or UO_888 (O_888,N_27591,N_27182);
xnor UO_889 (O_889,N_25276,N_26453);
or UO_890 (O_890,N_26836,N_28025);
nand UO_891 (O_891,N_27001,N_29191);
or UO_892 (O_892,N_26056,N_28903);
xor UO_893 (O_893,N_27365,N_27876);
nand UO_894 (O_894,N_25017,N_27791);
xor UO_895 (O_895,N_26887,N_27827);
nor UO_896 (O_896,N_26584,N_25823);
or UO_897 (O_897,N_25422,N_27635);
and UO_898 (O_898,N_29869,N_25326);
and UO_899 (O_899,N_25530,N_29898);
nor UO_900 (O_900,N_27883,N_27226);
nand UO_901 (O_901,N_26812,N_25790);
and UO_902 (O_902,N_25030,N_25058);
nand UO_903 (O_903,N_25964,N_28081);
or UO_904 (O_904,N_27463,N_29109);
and UO_905 (O_905,N_29004,N_26354);
or UO_906 (O_906,N_25657,N_29062);
and UO_907 (O_907,N_29607,N_28316);
nand UO_908 (O_908,N_26498,N_29865);
nor UO_909 (O_909,N_25578,N_28065);
nand UO_910 (O_910,N_26613,N_25721);
nand UO_911 (O_911,N_25209,N_28581);
or UO_912 (O_912,N_29866,N_25000);
xor UO_913 (O_913,N_26863,N_25994);
nand UO_914 (O_914,N_28035,N_27174);
nor UO_915 (O_915,N_28969,N_28146);
or UO_916 (O_916,N_27917,N_28183);
and UO_917 (O_917,N_28098,N_26997);
or UO_918 (O_918,N_25103,N_27377);
or UO_919 (O_919,N_29369,N_28798);
nand UO_920 (O_920,N_25818,N_29526);
and UO_921 (O_921,N_28692,N_27214);
nor UO_922 (O_922,N_28847,N_26931);
or UO_923 (O_923,N_28072,N_26449);
or UO_924 (O_924,N_29177,N_25731);
or UO_925 (O_925,N_29130,N_29428);
nor UO_926 (O_926,N_25885,N_26716);
and UO_927 (O_927,N_25678,N_28416);
or UO_928 (O_928,N_28515,N_25707);
or UO_929 (O_929,N_26993,N_28380);
or UO_930 (O_930,N_29324,N_27527);
xnor UO_931 (O_931,N_29950,N_27286);
nand UO_932 (O_932,N_29347,N_25975);
and UO_933 (O_933,N_27908,N_27695);
nand UO_934 (O_934,N_28605,N_26847);
and UO_935 (O_935,N_27370,N_28980);
and UO_936 (O_936,N_27271,N_29670);
xnor UO_937 (O_937,N_29857,N_26456);
nand UO_938 (O_938,N_28249,N_26818);
and UO_939 (O_939,N_28420,N_29765);
and UO_940 (O_940,N_28077,N_27102);
nor UO_941 (O_941,N_29611,N_26025);
nand UO_942 (O_942,N_25786,N_26580);
nand UO_943 (O_943,N_27934,N_27131);
nand UO_944 (O_944,N_27095,N_27571);
nand UO_945 (O_945,N_29998,N_25401);
and UO_946 (O_946,N_26510,N_29709);
nor UO_947 (O_947,N_25852,N_25753);
nor UO_948 (O_948,N_27627,N_29719);
xor UO_949 (O_949,N_27431,N_26898);
or UO_950 (O_950,N_27530,N_25631);
nand UO_951 (O_951,N_27047,N_29315);
and UO_952 (O_952,N_25579,N_28946);
and UO_953 (O_953,N_28895,N_27703);
and UO_954 (O_954,N_28896,N_26559);
nand UO_955 (O_955,N_25373,N_29064);
xor UO_956 (O_956,N_28565,N_25130);
or UO_957 (O_957,N_28194,N_28250);
or UO_958 (O_958,N_25843,N_27975);
and UO_959 (O_959,N_29726,N_26001);
xor UO_960 (O_960,N_28937,N_26549);
nor UO_961 (O_961,N_25146,N_28239);
nor UO_962 (O_962,N_26712,N_29878);
and UO_963 (O_963,N_27213,N_28574);
nor UO_964 (O_964,N_25377,N_27718);
and UO_965 (O_965,N_26758,N_28281);
or UO_966 (O_966,N_26252,N_28570);
xnor UO_967 (O_967,N_27634,N_29414);
or UO_968 (O_968,N_26564,N_25045);
nand UO_969 (O_969,N_25836,N_27358);
or UO_970 (O_970,N_28299,N_26648);
or UO_971 (O_971,N_25382,N_28174);
nand UO_972 (O_972,N_25175,N_28285);
and UO_973 (O_973,N_28979,N_25308);
or UO_974 (O_974,N_29027,N_27666);
or UO_975 (O_975,N_28807,N_27750);
or UO_976 (O_976,N_29235,N_28106);
or UO_977 (O_977,N_25827,N_29127);
nand UO_978 (O_978,N_27534,N_29343);
or UO_979 (O_979,N_26978,N_29133);
nand UO_980 (O_980,N_26971,N_26746);
or UO_981 (O_981,N_25444,N_25070);
nor UO_982 (O_982,N_27715,N_25338);
and UO_983 (O_983,N_29208,N_26376);
and UO_984 (O_984,N_27171,N_29691);
xnor UO_985 (O_985,N_29929,N_27573);
and UO_986 (O_986,N_26394,N_25044);
and UO_987 (O_987,N_26237,N_28233);
nand UO_988 (O_988,N_29448,N_29229);
or UO_989 (O_989,N_27011,N_26059);
and UO_990 (O_990,N_25717,N_29567);
nor UO_991 (O_991,N_28977,N_26829);
and UO_992 (O_992,N_29173,N_29873);
and UO_993 (O_993,N_27528,N_29742);
or UO_994 (O_994,N_26852,N_27156);
and UO_995 (O_995,N_26761,N_26392);
nor UO_996 (O_996,N_28648,N_25155);
nand UO_997 (O_997,N_25079,N_29785);
or UO_998 (O_998,N_25456,N_29794);
nor UO_999 (O_999,N_28948,N_27925);
nand UO_1000 (O_1000,N_28408,N_25207);
and UO_1001 (O_1001,N_29061,N_28323);
nand UO_1002 (O_1002,N_29682,N_26860);
xnor UO_1003 (O_1003,N_28766,N_26280);
and UO_1004 (O_1004,N_29600,N_28972);
or UO_1005 (O_1005,N_25767,N_25113);
nand UO_1006 (O_1006,N_26933,N_28024);
nand UO_1007 (O_1007,N_25750,N_27911);
xnor UO_1008 (O_1008,N_26704,N_26409);
nand UO_1009 (O_1009,N_25270,N_28917);
nand UO_1010 (O_1010,N_27803,N_25473);
and UO_1011 (O_1011,N_25411,N_28689);
nor UO_1012 (O_1012,N_27927,N_25628);
and UO_1013 (O_1013,N_25626,N_27424);
or UO_1014 (O_1014,N_28238,N_27073);
nor UO_1015 (O_1015,N_25346,N_27279);
nor UO_1016 (O_1016,N_26137,N_26543);
or UO_1017 (O_1017,N_26172,N_26044);
nand UO_1018 (O_1018,N_26082,N_28833);
nand UO_1019 (O_1019,N_25502,N_27984);
and UO_1020 (O_1020,N_27619,N_25645);
nand UO_1021 (O_1021,N_26874,N_28671);
or UO_1022 (O_1022,N_26248,N_26357);
nand UO_1023 (O_1023,N_27641,N_26671);
or UO_1024 (O_1024,N_28793,N_29527);
or UO_1025 (O_1025,N_26290,N_25598);
nand UO_1026 (O_1026,N_27862,N_29319);
or UO_1027 (O_1027,N_27181,N_29861);
and UO_1028 (O_1028,N_25732,N_29669);
nand UO_1029 (O_1029,N_27101,N_26789);
nand UO_1030 (O_1030,N_26395,N_29808);
xor UO_1031 (O_1031,N_26486,N_28097);
nor UO_1032 (O_1032,N_29922,N_26406);
xor UO_1033 (O_1033,N_26885,N_29220);
nand UO_1034 (O_1034,N_25634,N_29779);
and UO_1035 (O_1035,N_25104,N_28327);
nor UO_1036 (O_1036,N_29966,N_26606);
or UO_1037 (O_1037,N_25388,N_28009);
nor UO_1038 (O_1038,N_26869,N_29081);
nor UO_1039 (O_1039,N_25450,N_26295);
nor UO_1040 (O_1040,N_28294,N_26542);
nor UO_1041 (O_1041,N_28283,N_25808);
nor UO_1042 (O_1042,N_26207,N_26322);
and UO_1043 (O_1043,N_25477,N_26346);
nand UO_1044 (O_1044,N_29593,N_26122);
and UO_1045 (O_1045,N_26474,N_29520);
and UO_1046 (O_1046,N_25423,N_27189);
and UO_1047 (O_1047,N_26702,N_28933);
nor UO_1048 (O_1048,N_28517,N_26611);
and UO_1049 (O_1049,N_29690,N_26722);
or UO_1050 (O_1050,N_26553,N_28589);
and UO_1051 (O_1051,N_27144,N_28142);
xor UO_1052 (O_1052,N_28984,N_27817);
or UO_1053 (O_1053,N_27699,N_28771);
xnor UO_1054 (O_1054,N_26146,N_28644);
nor UO_1055 (O_1055,N_27114,N_29332);
and UO_1056 (O_1056,N_28790,N_25906);
nand UO_1057 (O_1057,N_26229,N_29112);
and UO_1058 (O_1058,N_28635,N_25597);
nand UO_1059 (O_1059,N_29009,N_26467);
xor UO_1060 (O_1060,N_29041,N_25529);
or UO_1061 (O_1061,N_27643,N_27964);
nand UO_1062 (O_1062,N_29456,N_26891);
nor UO_1063 (O_1063,N_27382,N_26995);
nor UO_1064 (O_1064,N_28242,N_25576);
and UO_1065 (O_1065,N_25002,N_29906);
and UO_1066 (O_1066,N_25174,N_28521);
nor UO_1067 (O_1067,N_27522,N_25442);
and UO_1068 (O_1068,N_28932,N_26718);
nor UO_1069 (O_1069,N_29964,N_25129);
xor UO_1070 (O_1070,N_29761,N_29320);
and UO_1071 (O_1071,N_25550,N_26110);
or UO_1072 (O_1072,N_26085,N_26246);
nand UO_1073 (O_1073,N_29973,N_27805);
xor UO_1074 (O_1074,N_27428,N_26139);
or UO_1075 (O_1075,N_28996,N_26492);
nor UO_1076 (O_1076,N_25169,N_27357);
nor UO_1077 (O_1077,N_27500,N_25121);
and UO_1078 (O_1078,N_25881,N_28429);
and UO_1079 (O_1079,N_27651,N_28143);
xor UO_1080 (O_1080,N_28838,N_26318);
or UO_1081 (O_1081,N_29249,N_27464);
and UO_1082 (O_1082,N_29656,N_25287);
or UO_1083 (O_1083,N_28306,N_28567);
nand UO_1084 (O_1084,N_25138,N_27632);
or UO_1085 (O_1085,N_26868,N_25661);
or UO_1086 (O_1086,N_28734,N_26558);
nand UO_1087 (O_1087,N_26911,N_27763);
nand UO_1088 (O_1088,N_25922,N_29142);
and UO_1089 (O_1089,N_25331,N_25519);
nor UO_1090 (O_1090,N_29620,N_29095);
nor UO_1091 (O_1091,N_27350,N_28899);
nand UO_1092 (O_1092,N_28438,N_29342);
and UO_1093 (O_1093,N_28534,N_28154);
and UO_1094 (O_1094,N_25072,N_25211);
or UO_1095 (O_1095,N_29196,N_27175);
or UO_1096 (O_1096,N_26128,N_29517);
and UO_1097 (O_1097,N_26119,N_28237);
nor UO_1098 (O_1098,N_27071,N_27570);
nand UO_1099 (O_1099,N_25128,N_27337);
nor UO_1100 (O_1100,N_25869,N_25683);
and UO_1101 (O_1101,N_29774,N_26180);
nor UO_1102 (O_1102,N_29537,N_27637);
and UO_1103 (O_1103,N_25147,N_28590);
and UO_1104 (O_1104,N_26404,N_26271);
and UO_1105 (O_1105,N_28883,N_29636);
and UO_1106 (O_1106,N_29986,N_28471);
nor UO_1107 (O_1107,N_28368,N_26103);
nor UO_1108 (O_1108,N_29155,N_28149);
and UO_1109 (O_1109,N_25755,N_28732);
and UO_1110 (O_1110,N_26661,N_27581);
nor UO_1111 (O_1111,N_26890,N_28563);
and UO_1112 (O_1112,N_25780,N_28495);
xor UO_1113 (O_1113,N_29891,N_29073);
and UO_1114 (O_1114,N_28785,N_28357);
nor UO_1115 (O_1115,N_25756,N_29711);
nand UO_1116 (O_1116,N_25004,N_27615);
or UO_1117 (O_1117,N_28506,N_27752);
nand UO_1118 (O_1118,N_25840,N_28125);
or UO_1119 (O_1119,N_28957,N_25394);
nand UO_1120 (O_1120,N_25457,N_29788);
nor UO_1121 (O_1121,N_25365,N_29145);
nor UO_1122 (O_1122,N_27829,N_26701);
nor UO_1123 (O_1123,N_29420,N_25998);
nand UO_1124 (O_1124,N_25589,N_26832);
xor UO_1125 (O_1125,N_27153,N_29005);
and UO_1126 (O_1126,N_28411,N_27801);
nor UO_1127 (O_1127,N_27920,N_29370);
and UO_1128 (O_1128,N_25345,N_27923);
or UO_1129 (O_1129,N_26304,N_29846);
nand UO_1130 (O_1130,N_25459,N_29470);
and UO_1131 (O_1131,N_27556,N_26776);
nand UO_1132 (O_1132,N_26685,N_26489);
nand UO_1133 (O_1133,N_27919,N_26353);
nor UO_1134 (O_1134,N_27288,N_26665);
or UO_1135 (O_1135,N_25729,N_25822);
and UO_1136 (O_1136,N_28678,N_28445);
or UO_1137 (O_1137,N_28158,N_27110);
xnor UO_1138 (O_1138,N_27049,N_25329);
and UO_1139 (O_1139,N_29240,N_26598);
or UO_1140 (O_1140,N_26223,N_25430);
or UO_1141 (O_1141,N_29406,N_29469);
or UO_1142 (O_1142,N_25911,N_25454);
nor UO_1143 (O_1143,N_25784,N_26408);
nand UO_1144 (O_1144,N_29348,N_26177);
and UO_1145 (O_1145,N_29445,N_26770);
or UO_1146 (O_1146,N_27485,N_28665);
xnor UO_1147 (O_1147,N_25372,N_26261);
nor UO_1148 (O_1148,N_25856,N_29144);
nor UO_1149 (O_1149,N_27692,N_29122);
nor UO_1150 (O_1150,N_29180,N_28768);
or UO_1151 (O_1151,N_25488,N_25412);
and UO_1152 (O_1152,N_28227,N_28487);
nand UO_1153 (O_1153,N_25301,N_27886);
nor UO_1154 (O_1154,N_27207,N_28646);
nor UO_1155 (O_1155,N_28609,N_28382);
nor UO_1156 (O_1156,N_26582,N_26697);
nor UO_1157 (O_1157,N_26878,N_26578);
nand UO_1158 (O_1158,N_28832,N_25987);
nand UO_1159 (O_1159,N_27572,N_26566);
nor UO_1160 (O_1160,N_27065,N_29544);
xnor UO_1161 (O_1161,N_28621,N_26698);
nand UO_1162 (O_1162,N_29200,N_26245);
nand UO_1163 (O_1163,N_26516,N_27987);
nand UO_1164 (O_1164,N_26679,N_26438);
xor UO_1165 (O_1165,N_27310,N_25261);
nand UO_1166 (O_1166,N_26366,N_25149);
and UO_1167 (O_1167,N_29083,N_26345);
nor UO_1168 (O_1168,N_28488,N_25913);
nor UO_1169 (O_1169,N_26907,N_27650);
nor UO_1170 (O_1170,N_25613,N_26047);
nand UO_1171 (O_1171,N_28794,N_25709);
nor UO_1172 (O_1172,N_25141,N_26669);
nor UO_1173 (O_1173,N_28041,N_27949);
nand UO_1174 (O_1174,N_25624,N_27442);
nor UO_1175 (O_1175,N_29519,N_26031);
or UO_1176 (O_1176,N_26116,N_25989);
nor UO_1177 (O_1177,N_26835,N_27484);
and UO_1178 (O_1178,N_28746,N_28968);
and UO_1179 (O_1179,N_25196,N_28455);
nor UO_1180 (O_1180,N_28670,N_28927);
and UO_1181 (O_1181,N_29198,N_27364);
nand UO_1182 (O_1182,N_27518,N_28070);
nor UO_1183 (O_1183,N_28164,N_28275);
and UO_1184 (O_1184,N_27298,N_27848);
nor UO_1185 (O_1185,N_28986,N_25449);
nand UO_1186 (O_1186,N_28465,N_29845);
nand UO_1187 (O_1187,N_27724,N_27470);
nor UO_1188 (O_1188,N_27804,N_27375);
and UO_1189 (O_1189,N_26298,N_29028);
nand UO_1190 (O_1190,N_25646,N_28109);
or UO_1191 (O_1191,N_26274,N_28073);
or UO_1192 (O_1192,N_27644,N_29698);
xor UO_1193 (O_1193,N_27302,N_28735);
or UO_1194 (O_1194,N_28636,N_29763);
or UO_1195 (O_1195,N_26081,N_27432);
nor UO_1196 (O_1196,N_25236,N_29405);
nand UO_1197 (O_1197,N_28943,N_28207);
or UO_1198 (O_1198,N_26469,N_27403);
and UO_1199 (O_1199,N_29735,N_27852);
nor UO_1200 (O_1200,N_28886,N_29979);
nand UO_1201 (O_1201,N_27654,N_27472);
nor UO_1202 (O_1202,N_28568,N_25042);
or UO_1203 (O_1203,N_25566,N_29478);
and UO_1204 (O_1204,N_25220,N_27481);
nor UO_1205 (O_1205,N_28462,N_27921);
or UO_1206 (O_1206,N_29432,N_28557);
nor UO_1207 (O_1207,N_25925,N_28863);
and UO_1208 (O_1208,N_28104,N_26654);
or UO_1209 (O_1209,N_27607,N_29192);
or UO_1210 (O_1210,N_29889,N_28606);
or UO_1211 (O_1211,N_29777,N_26929);
and UO_1212 (O_1212,N_27994,N_29631);
or UO_1213 (O_1213,N_27785,N_25253);
and UO_1214 (O_1214,N_29660,N_29949);
or UO_1215 (O_1215,N_25572,N_29824);
or UO_1216 (O_1216,N_29888,N_26273);
or UO_1217 (O_1217,N_28502,N_29930);
nor UO_1218 (O_1218,N_27569,N_28955);
and UO_1219 (O_1219,N_27820,N_25249);
and UO_1220 (O_1220,N_28269,N_28220);
nand UO_1221 (O_1221,N_27625,N_26723);
nor UO_1222 (O_1222,N_29575,N_29261);
xnor UO_1223 (O_1223,N_25740,N_25027);
xor UO_1224 (O_1224,N_26895,N_26696);
nand UO_1225 (O_1225,N_27892,N_25243);
nor UO_1226 (O_1226,N_26356,N_29997);
and UO_1227 (O_1227,N_28579,N_27766);
nand UO_1228 (O_1228,N_28941,N_27061);
and UO_1229 (O_1229,N_29634,N_29431);
nand UO_1230 (O_1230,N_26383,N_29113);
nand UO_1231 (O_1231,N_28478,N_26152);
nand UO_1232 (O_1232,N_28115,N_28612);
nor UO_1233 (O_1233,N_28528,N_26183);
nor UO_1234 (O_1234,N_26454,N_25924);
xor UO_1235 (O_1235,N_26915,N_25349);
and UO_1236 (O_1236,N_29867,N_29391);
nand UO_1237 (O_1237,N_26754,N_27523);
nand UO_1238 (O_1238,N_27907,N_29816);
nand UO_1239 (O_1239,N_25127,N_26830);
nand UO_1240 (O_1240,N_29164,N_26787);
nand UO_1241 (O_1241,N_25177,N_29837);
and UO_1242 (O_1242,N_29610,N_28415);
xor UO_1243 (O_1243,N_25761,N_27618);
xnor UO_1244 (O_1244,N_25410,N_25910);
and UO_1245 (O_1245,N_25514,N_28654);
nand UO_1246 (O_1246,N_28172,N_29764);
nor UO_1247 (O_1247,N_26755,N_29500);
xnor UO_1248 (O_1248,N_29082,N_25040);
and UO_1249 (O_1249,N_28803,N_25033);
and UO_1250 (O_1250,N_28965,N_27870);
or UO_1251 (O_1251,N_27693,N_25819);
or UO_1252 (O_1252,N_28441,N_29207);
and UO_1253 (O_1253,N_29596,N_28618);
nor UO_1254 (O_1254,N_28451,N_25931);
or UO_1255 (O_1255,N_27592,N_25863);
or UO_1256 (O_1256,N_29759,N_27762);
nand UO_1257 (O_1257,N_27614,N_29786);
nand UO_1258 (O_1258,N_29582,N_26132);
or UO_1259 (O_1259,N_25556,N_26440);
and UO_1260 (O_1260,N_25096,N_25610);
or UO_1261 (O_1261,N_25695,N_28696);
and UO_1262 (O_1262,N_29499,N_28925);
or UO_1263 (O_1263,N_25038,N_25416);
xor UO_1264 (O_1264,N_29421,N_26311);
xor UO_1265 (O_1265,N_29086,N_27219);
nand UO_1266 (O_1266,N_25064,N_26042);
nand UO_1267 (O_1267,N_26154,N_26772);
nand UO_1268 (O_1268,N_28763,N_25392);
nor UO_1269 (O_1269,N_28719,N_27299);
nor UO_1270 (O_1270,N_25084,N_25091);
nand UO_1271 (O_1271,N_28135,N_27590);
xor UO_1272 (O_1272,N_26397,N_27777);
nand UO_1273 (O_1273,N_29564,N_25802);
nand UO_1274 (O_1274,N_29232,N_29771);
nand UO_1275 (O_1275,N_27281,N_25071);
nor UO_1276 (O_1276,N_29056,N_25351);
and UO_1277 (O_1277,N_25915,N_29383);
xor UO_1278 (O_1278,N_25981,N_27072);
and UO_1279 (O_1279,N_27617,N_25561);
or UO_1280 (O_1280,N_27646,N_26762);
xnor UO_1281 (O_1281,N_26961,N_25279);
nand UO_1282 (O_1282,N_28293,N_27409);
or UO_1283 (O_1283,N_28784,N_27788);
nand UO_1284 (O_1284,N_29151,N_26064);
nor UO_1285 (O_1285,N_28588,N_26104);
xnor UO_1286 (O_1286,N_28513,N_25163);
and UO_1287 (O_1287,N_28032,N_27024);
and UO_1288 (O_1288,N_25974,N_27992);
or UO_1289 (O_1289,N_28641,N_29739);
nor UO_1290 (O_1290,N_28071,N_26168);
nand UO_1291 (O_1291,N_28038,N_26744);
nand UO_1292 (O_1292,N_28613,N_26977);
and UO_1293 (O_1293,N_27045,N_28353);
nor UO_1294 (O_1294,N_27237,N_28152);
and UO_1295 (O_1295,N_26547,N_26142);
and UO_1296 (O_1296,N_29213,N_29257);
or UO_1297 (O_1297,N_26861,N_29382);
nor UO_1298 (O_1298,N_27906,N_28052);
and UO_1299 (O_1299,N_27794,N_28708);
nor UO_1300 (O_1300,N_29531,N_29471);
and UO_1301 (O_1301,N_25154,N_27577);
nor UO_1302 (O_1302,N_26004,N_29805);
nor UO_1303 (O_1303,N_26944,N_26090);
xor UO_1304 (O_1304,N_29134,N_25540);
or UO_1305 (O_1305,N_29825,N_27597);
or UO_1306 (O_1306,N_25235,N_25771);
or UO_1307 (O_1307,N_25587,N_25417);
xnor UO_1308 (O_1308,N_25083,N_26568);
nand UO_1309 (O_1309,N_28773,N_26660);
nor UO_1310 (O_1310,N_26573,N_28151);
and UO_1311 (O_1311,N_27259,N_25512);
nor UO_1312 (O_1312,N_27313,N_25006);
nor UO_1313 (O_1313,N_29854,N_27690);
nand UO_1314 (O_1314,N_25860,N_29635);
nor UO_1315 (O_1315,N_27078,N_28232);
or UO_1316 (O_1316,N_28208,N_27167);
and UO_1317 (O_1317,N_28319,N_25604);
and UO_1318 (O_1318,N_29337,N_26264);
nand UO_1319 (O_1319,N_26032,N_26370);
nand UO_1320 (O_1320,N_27550,N_27139);
nor UO_1321 (O_1321,N_26653,N_29246);
or UO_1322 (O_1322,N_29963,N_25739);
or UO_1323 (O_1323,N_25248,N_28278);
nand UO_1324 (O_1324,N_28398,N_28861);
and UO_1325 (O_1325,N_26690,N_26632);
nor UO_1326 (O_1326,N_29902,N_28888);
or UO_1327 (O_1327,N_25722,N_25972);
nand UO_1328 (O_1328,N_28619,N_29174);
or UO_1329 (O_1329,N_27901,N_26656);
nand UO_1330 (O_1330,N_29040,N_29689);
and UO_1331 (O_1331,N_26107,N_27604);
or UO_1332 (O_1332,N_25567,N_28361);
and UO_1333 (O_1333,N_25195,N_27141);
or UO_1334 (O_1334,N_25297,N_26555);
nor UO_1335 (O_1335,N_26344,N_28985);
xor UO_1336 (O_1336,N_29658,N_25571);
nand UO_1337 (O_1337,N_28844,N_26581);
nor UO_1338 (O_1338,N_26785,N_25507);
and UO_1339 (O_1339,N_28730,N_27120);
xor UO_1340 (O_1340,N_25277,N_28687);
xnor UO_1341 (O_1341,N_27605,N_26839);
nor UO_1342 (O_1342,N_26550,N_29325);
xor UO_1343 (O_1343,N_29688,N_25741);
nand UO_1344 (O_1344,N_26462,N_27686);
nor UO_1345 (O_1345,N_27496,N_27823);
nor UO_1346 (O_1346,N_29100,N_26763);
nor UO_1347 (O_1347,N_29125,N_29263);
or UO_1348 (O_1348,N_25821,N_26473);
nand UO_1349 (O_1349,N_26148,N_26230);
xnor UO_1350 (O_1350,N_25890,N_26619);
xnor UO_1351 (O_1351,N_28575,N_25118);
nor UO_1352 (O_1352,N_26668,N_28698);
nand UO_1353 (O_1353,N_25333,N_28742);
nor UO_1354 (O_1354,N_27076,N_27560);
and UO_1355 (O_1355,N_27385,N_25545);
nor UO_1356 (O_1356,N_28906,N_28777);
and UO_1357 (O_1357,N_28792,N_29553);
and UO_1358 (O_1358,N_29364,N_26124);
xor UO_1359 (O_1359,N_25845,N_27035);
and UO_1360 (O_1360,N_29397,N_26377);
or UO_1361 (O_1361,N_27320,N_27474);
and UO_1362 (O_1362,N_28672,N_26708);
and UO_1363 (O_1363,N_25080,N_27793);
and UO_1364 (O_1364,N_28694,N_25542);
or UO_1365 (O_1365,N_29416,N_29917);
nand UO_1366 (O_1366,N_26713,N_27254);
xnor UO_1367 (O_1367,N_29841,N_26538);
xor UO_1368 (O_1368,N_29184,N_27564);
and UO_1369 (O_1369,N_25919,N_28950);
nor UO_1370 (O_1370,N_25228,N_29170);
nand UO_1371 (O_1371,N_28673,N_28301);
or UO_1372 (O_1372,N_27039,N_28942);
nor UO_1373 (O_1373,N_26795,N_28037);
or UO_1374 (O_1374,N_29367,N_28121);
or UO_1375 (O_1375,N_27515,N_25993);
and UO_1376 (O_1376,N_29511,N_25575);
nand UO_1377 (O_1377,N_26412,N_25862);
or UO_1378 (O_1378,N_26784,N_25543);
nor UO_1379 (O_1379,N_25126,N_25979);
nand UO_1380 (O_1380,N_29225,N_25258);
nand UO_1381 (O_1381,N_27940,N_25696);
or UO_1382 (O_1382,N_27184,N_27115);
nor UO_1383 (O_1383,N_25669,N_26011);
nor UO_1384 (O_1384,N_29118,N_25706);
nand UO_1385 (O_1385,N_26413,N_25339);
nand UO_1386 (O_1386,N_28828,N_28334);
nand UO_1387 (O_1387,N_26949,N_29882);
nand UO_1388 (O_1388,N_27355,N_26471);
xor UO_1389 (O_1389,N_26078,N_27196);
nand UO_1390 (O_1390,N_26532,N_29928);
or UO_1391 (O_1391,N_27308,N_29430);
nor UO_1392 (O_1392,N_26162,N_26048);
nand UO_1393 (O_1393,N_26109,N_25704);
nor UO_1394 (O_1394,N_27678,N_27535);
and UO_1395 (O_1395,N_26941,N_28126);
nand UO_1396 (O_1396,N_25544,N_26975);
or UO_1397 (O_1397,N_27426,N_26269);
or UO_1398 (O_1398,N_27010,N_28118);
nand UO_1399 (O_1399,N_27841,N_28835);
nand UO_1400 (O_1400,N_28631,N_29551);
or UO_1401 (O_1401,N_27962,N_27861);
nor UO_1402 (O_1402,N_26077,N_27075);
or UO_1403 (O_1403,N_28891,N_29483);
and UO_1404 (O_1404,N_29663,N_27624);
and UO_1405 (O_1405,N_27506,N_27400);
or UO_1406 (O_1406,N_25996,N_28433);
nor UO_1407 (O_1407,N_29910,N_29958);
nand UO_1408 (O_1408,N_27351,N_27976);
nor UO_1409 (O_1409,N_27438,N_27728);
nand UO_1410 (O_1410,N_29328,N_28841);
or UO_1411 (O_1411,N_25847,N_26623);
or UO_1412 (O_1412,N_28767,N_28209);
and UO_1413 (O_1413,N_26003,N_29399);
and UO_1414 (O_1414,N_28911,N_26823);
nor UO_1415 (O_1415,N_28255,N_29222);
and UO_1416 (O_1416,N_25144,N_25857);
or UO_1417 (O_1417,N_26336,N_28852);
nor UO_1418 (O_1418,N_28738,N_26130);
nand UO_1419 (O_1419,N_28308,N_26512);
nand UO_1420 (O_1420,N_27857,N_27660);
nor UO_1421 (O_1421,N_29716,N_27316);
and UO_1422 (O_1422,N_27284,N_29355);
nor UO_1423 (O_1423,N_28344,N_26066);
xnor UO_1424 (O_1424,N_26086,N_28543);
nor UO_1425 (O_1425,N_26998,N_29380);
nor UO_1426 (O_1426,N_26883,N_25305);
nor UO_1427 (O_1427,N_29528,N_28216);
nand UO_1428 (O_1428,N_28676,N_26537);
and UO_1429 (O_1429,N_29466,N_29385);
nor UO_1430 (O_1430,N_27872,N_26985);
nor UO_1431 (O_1431,N_25358,N_29340);
or UO_1432 (O_1432,N_29258,N_27466);
nand UO_1433 (O_1433,N_26865,N_29085);
nor UO_1434 (O_1434,N_27040,N_29068);
nand UO_1435 (O_1435,N_28470,N_28053);
nand UO_1436 (O_1436,N_28651,N_27586);
and UO_1437 (O_1437,N_29219,N_28434);
or UO_1438 (O_1438,N_26589,N_26730);
and UO_1439 (O_1439,N_28940,N_25986);
or UO_1440 (O_1440,N_28197,N_25035);
or UO_1441 (O_1441,N_29799,N_28758);
xor UO_1442 (O_1442,N_28469,N_25644);
and UO_1443 (O_1443,N_28333,N_27501);
nor UO_1444 (O_1444,N_26445,N_28658);
nand UO_1445 (O_1445,N_27544,N_26587);
and UO_1446 (O_1446,N_28512,N_27596);
or UO_1447 (O_1447,N_28706,N_27630);
and UO_1448 (O_1448,N_29583,N_27318);
nor UO_1449 (O_1449,N_26650,N_27458);
xnor UO_1450 (O_1450,N_28988,N_28211);
nand UO_1451 (O_1451,N_26571,N_26022);
or UO_1452 (O_1452,N_29150,N_28952);
nand UO_1453 (O_1453,N_25638,N_25244);
nor UO_1454 (O_1454,N_29832,N_26726);
xnor UO_1455 (O_1455,N_26955,N_29974);
xnor UO_1456 (O_1456,N_26657,N_28645);
nor UO_1457 (O_1457,N_26844,N_29293);
nor UO_1458 (O_1458,N_25467,N_27389);
or UO_1459 (O_1459,N_25517,N_27107);
nand UO_1460 (O_1460,N_26221,N_27672);
xor UO_1461 (O_1461,N_28377,N_28554);
and UO_1462 (O_1462,N_28399,N_27874);
nand UO_1463 (O_1463,N_28797,N_27273);
or UO_1464 (O_1464,N_25595,N_25367);
xnor UO_1465 (O_1465,N_27105,N_25432);
and UO_1466 (O_1466,N_26889,N_28264);
and UO_1467 (O_1467,N_26676,N_25462);
and UO_1468 (O_1468,N_27568,N_26488);
nand UO_1469 (O_1469,N_28585,N_28681);
or UO_1470 (O_1470,N_29988,N_29720);
nor UO_1471 (O_1471,N_26209,N_27539);
nor UO_1472 (O_1472,N_25880,N_26101);
and UO_1473 (O_1473,N_27945,N_27747);
nand UO_1474 (O_1474,N_29831,N_26240);
nand UO_1475 (O_1475,N_28849,N_27012);
and UO_1476 (O_1476,N_25521,N_25549);
and UO_1477 (O_1477,N_26405,N_28840);
or UO_1478 (O_1478,N_27575,N_27997);
nor UO_1479 (O_1479,N_26515,N_27936);
or UO_1480 (O_1480,N_29677,N_29425);
nor UO_1481 (O_1481,N_25546,N_27731);
xnor UO_1482 (O_1482,N_29291,N_29981);
nor UO_1483 (O_1483,N_25671,N_28503);
and UO_1484 (O_1484,N_27878,N_29157);
or UO_1485 (O_1485,N_28947,N_28287);
and UO_1486 (O_1486,N_29664,N_25302);
nand UO_1487 (O_1487,N_26841,N_29129);
nand UO_1488 (O_1488,N_28391,N_29104);
nand UO_1489 (O_1489,N_25407,N_26105);
and UO_1490 (O_1490,N_25675,N_27498);
or UO_1491 (O_1491,N_28551,N_28147);
and UO_1492 (O_1492,N_25059,N_26052);
or UO_1493 (O_1493,N_28939,N_25097);
and UO_1494 (O_1494,N_26737,N_27948);
xor UO_1495 (O_1495,N_25493,N_27183);
or UO_1496 (O_1496,N_26913,N_28931);
nand UO_1497 (O_1497,N_27081,N_29424);
or UO_1498 (O_1498,N_28185,N_29035);
nand UO_1499 (O_1499,N_27669,N_25937);
xnor UO_1500 (O_1500,N_27255,N_27413);
or UO_1501 (O_1501,N_25757,N_27077);
nor UO_1502 (O_1502,N_28170,N_25944);
or UO_1503 (O_1503,N_29822,N_29379);
and UO_1504 (O_1504,N_29096,N_28789);
or UO_1505 (O_1505,N_27441,N_26296);
nand UO_1506 (O_1506,N_29601,N_25804);
and UO_1507 (O_1507,N_29702,N_26198);
nor UO_1508 (O_1508,N_27675,N_25186);
nor UO_1509 (O_1509,N_29044,N_25082);
xnor UO_1510 (O_1510,N_28443,N_29330);
or UO_1511 (O_1511,N_29077,N_25796);
xnor UO_1512 (O_1512,N_27295,N_28760);
and UO_1513 (O_1513,N_25452,N_27074);
and UO_1514 (O_1514,N_25828,N_29740);
and UO_1515 (O_1515,N_28463,N_29123);
nor UO_1516 (O_1516,N_29012,N_25812);
or UO_1517 (O_1517,N_28640,N_26074);
nand UO_1518 (O_1518,N_29439,N_25067);
nor UO_1519 (O_1519,N_25028,N_27982);
or UO_1520 (O_1520,N_25007,N_29252);
or UO_1521 (O_1521,N_26213,N_25495);
or UO_1522 (O_1522,N_26040,N_27711);
or UO_1523 (O_1523,N_26757,N_28144);
and UO_1524 (O_1524,N_28412,N_27084);
nand UO_1525 (O_1525,N_29989,N_29776);
and UO_1526 (O_1526,N_29158,N_28376);
nand UO_1527 (O_1527,N_26806,N_29065);
and UO_1528 (O_1528,N_29171,N_29001);
nor UO_1529 (O_1529,N_28160,N_28580);
or UO_1530 (O_1530,N_28340,N_29345);
nand UO_1531 (O_1531,N_28959,N_25903);
and UO_1532 (O_1532,N_25384,N_25746);
or UO_1533 (O_1533,N_27710,N_25861);
nand UO_1534 (O_1534,N_27003,N_25504);
nor UO_1535 (O_1535,N_26181,N_26079);
and UO_1536 (O_1536,N_25139,N_25983);
or UO_1537 (O_1537,N_25193,N_26576);
or UO_1538 (O_1538,N_25801,N_26511);
nand UO_1539 (O_1539,N_25532,N_26315);
and UO_1540 (O_1540,N_28547,N_27746);
or UO_1541 (O_1541,N_27489,N_29555);
nor UO_1542 (O_1542,N_29708,N_28817);
nand UO_1543 (O_1543,N_26692,N_25267);
and UO_1544 (O_1544,N_29599,N_25500);
or UO_1545 (O_1545,N_25156,N_26435);
nand UO_1546 (O_1546,N_27224,N_27521);
nor UO_1547 (O_1547,N_29707,N_25202);
and UO_1548 (O_1548,N_26051,N_26297);
nor UO_1549 (O_1549,N_25949,N_27732);
or UO_1550 (O_1550,N_28532,N_25311);
nor UO_1551 (O_1551,N_25223,N_25536);
nor UO_1552 (O_1552,N_25574,N_25092);
nand UO_1553 (O_1553,N_28479,N_29868);
or UO_1554 (O_1554,N_26250,N_26317);
nand UO_1555 (O_1555,N_29614,N_29271);
nand UO_1556 (O_1556,N_29723,N_27744);
xor UO_1557 (O_1557,N_25655,N_28535);
and UO_1558 (O_1558,N_29356,N_27647);
and UO_1559 (O_1559,N_28680,N_25958);
nand UO_1560 (O_1560,N_26825,N_29049);
nor UO_1561 (O_1561,N_28781,N_25052);
nor UO_1562 (O_1562,N_27119,N_26476);
xnor UO_1563 (O_1563,N_26640,N_29495);
nor UO_1564 (O_1564,N_28452,N_29800);
and UO_1565 (O_1565,N_25176,N_28889);
nand UO_1566 (O_1566,N_29945,N_27603);
and UO_1567 (O_1567,N_29110,N_27098);
nor UO_1568 (O_1568,N_25398,N_29093);
nor UO_1569 (O_1569,N_25584,N_29699);
and UO_1570 (O_1570,N_26901,N_28772);
and UO_1571 (O_1571,N_27636,N_26595);
and UO_1572 (O_1572,N_27622,N_26414);
nor UO_1573 (O_1573,N_29314,N_25844);
nor UO_1574 (O_1574,N_28124,N_27609);
xor UO_1575 (O_1575,N_29895,N_25960);
nand UO_1576 (O_1576,N_28217,N_28921);
xor UO_1577 (O_1577,N_26224,N_27600);
nand UO_1578 (O_1578,N_29737,N_25400);
nand UO_1579 (O_1579,N_28783,N_28120);
and UO_1580 (O_1580,N_29497,N_25639);
or UO_1581 (O_1581,N_27796,N_26118);
or UO_1582 (O_1582,N_26007,N_27205);
or UO_1583 (O_1583,N_25654,N_25811);
xor UO_1584 (O_1584,N_25191,N_26539);
or UO_1585 (O_1585,N_25833,N_27282);
and UO_1586 (O_1586,N_25438,N_25563);
nor UO_1587 (O_1587,N_28561,N_26220);
nand UO_1588 (O_1588,N_27405,N_27990);
or UO_1589 (O_1589,N_28062,N_25798);
nor UO_1590 (O_1590,N_25900,N_25946);
or UO_1591 (O_1591,N_26710,N_26184);
and UO_1592 (O_1592,N_26672,N_25402);
and UO_1593 (O_1593,N_28273,N_29300);
or UO_1594 (O_1594,N_29721,N_26548);
nor UO_1595 (O_1595,N_29522,N_29374);
or UO_1596 (O_1596,N_26652,N_29285);
xor UO_1597 (O_1597,N_25435,N_26477);
nor UO_1598 (O_1598,N_29626,N_27507);
nor UO_1599 (O_1599,N_25483,N_29830);
xnor UO_1600 (O_1600,N_29290,N_26649);
nor UO_1601 (O_1601,N_28450,N_27661);
or UO_1602 (O_1602,N_29982,N_26523);
nor UO_1603 (O_1603,N_27381,N_27508);
nand UO_1604 (O_1604,N_26206,N_26884);
or UO_1605 (O_1605,N_25592,N_25859);
or UO_1606 (O_1606,N_28372,N_29030);
or UO_1607 (O_1607,N_28291,N_26281);
nor UO_1608 (O_1608,N_27559,N_28990);
nor UO_1609 (O_1609,N_26973,N_28747);
nor UO_1610 (O_1610,N_27393,N_25785);
nor UO_1611 (O_1611,N_29843,N_29309);
nor UO_1612 (O_1612,N_26936,N_29847);
or UO_1613 (O_1613,N_26131,N_26605);
nor UO_1614 (O_1614,N_25208,N_27685);
and UO_1615 (O_1615,N_29510,N_27343);
or UO_1616 (O_1616,N_27551,N_26734);
nor UO_1617 (O_1617,N_25875,N_28752);
or UO_1618 (O_1618,N_27988,N_29195);
nand UO_1619 (O_1619,N_25482,N_27691);
and UO_1620 (O_1620,N_25445,N_25316);
nor UO_1621 (O_1621,N_25562,N_25161);
nand UO_1622 (O_1622,N_25012,N_25447);
nand UO_1623 (O_1623,N_27537,N_28714);
and UO_1624 (O_1624,N_28240,N_26767);
or UO_1625 (O_1625,N_27450,N_28224);
xor UO_1626 (O_1626,N_26310,N_26925);
or UO_1627 (O_1627,N_28054,N_27268);
nand UO_1628 (O_1628,N_29968,N_29595);
and UO_1629 (O_1629,N_25904,N_28723);
nor UO_1630 (O_1630,N_28787,N_26853);
nor UO_1631 (O_1631,N_25424,N_28750);
or UO_1632 (O_1632,N_25274,N_29212);
nand UO_1633 (O_1633,N_26029,N_25437);
and UO_1634 (O_1634,N_26992,N_29772);
and UO_1635 (O_1635,N_25264,N_29757);
or UO_1636 (O_1636,N_27335,N_25094);
nand UO_1637 (O_1637,N_25742,N_26540);
nor UO_1638 (O_1638,N_29311,N_27027);
or UO_1639 (O_1639,N_29617,N_27953);
nand UO_1640 (O_1640,N_29186,N_29387);
or UO_1641 (O_1641,N_27079,N_25239);
nor UO_1642 (O_1642,N_29079,N_29623);
or UO_1643 (O_1643,N_26307,N_28964);
xor UO_1644 (O_1644,N_28639,N_26988);
nor UO_1645 (O_1645,N_29388,N_29353);
nand UO_1646 (O_1646,N_29426,N_25255);
xnor UO_1647 (O_1647,N_26300,N_25306);
and UO_1648 (O_1648,N_26058,N_27491);
or UO_1649 (O_1649,N_25614,N_26088);
nor UO_1650 (O_1650,N_25716,N_25328);
and UO_1651 (O_1651,N_29094,N_26054);
and UO_1652 (O_1652,N_28168,N_26028);
xnor UO_1653 (O_1653,N_26303,N_27468);
or UO_1654 (O_1654,N_28419,N_26157);
nand UO_1655 (O_1655,N_25554,N_26783);
or UO_1656 (O_1656,N_27933,N_26546);
xnor UO_1657 (O_1657,N_29883,N_29349);
and UO_1658 (O_1658,N_29909,N_26423);
nand UO_1659 (O_1659,N_29781,N_26403);
xor UO_1660 (O_1660,N_27567,N_26112);
and UO_1661 (O_1661,N_29245,N_29775);
nor UO_1662 (O_1662,N_25738,N_29962);
or UO_1663 (O_1663,N_29189,N_28156);
and UO_1664 (O_1664,N_27973,N_29216);
nand UO_1665 (O_1665,N_28311,N_25718);
nor UO_1666 (O_1666,N_27735,N_26986);
and UO_1667 (O_1667,N_29346,N_27859);
or UO_1668 (O_1668,N_25759,N_29452);
xnor UO_1669 (O_1669,N_28722,N_29790);
or UO_1670 (O_1670,N_28712,N_27688);
nand UO_1671 (O_1671,N_26579,N_26567);
or UO_1672 (O_1672,N_28780,N_25793);
and UO_1673 (O_1673,N_27007,N_28632);
nor UO_1674 (O_1674,N_26666,N_27457);
and UO_1675 (O_1675,N_29795,N_26441);
nand UO_1676 (O_1676,N_25286,N_28664);
nor UO_1677 (O_1677,N_29530,N_29043);
or UO_1678 (O_1678,N_27390,N_25268);
or UO_1679 (O_1679,N_27309,N_26485);
nand UO_1680 (O_1680,N_26947,N_26083);
nand UO_1681 (O_1681,N_26994,N_25637);
or UO_1682 (O_1682,N_26287,N_27639);
and UO_1683 (O_1683,N_28064,N_28103);
nand UO_1684 (O_1684,N_28804,N_26481);
nor UO_1685 (O_1685,N_27112,N_26826);
or UO_1686 (O_1686,N_28473,N_28916);
and UO_1687 (O_1687,N_29899,N_25192);
and UO_1688 (O_1688,N_28607,N_28560);
nand UO_1689 (O_1689,N_26544,N_29615);
nor UO_1690 (O_1690,N_29003,N_29842);
and UO_1691 (O_1691,N_25930,N_28182);
nor UO_1692 (O_1692,N_29589,N_29619);
xor UO_1693 (O_1693,N_27712,N_26227);
and UO_1694 (O_1694,N_26517,N_26463);
and UO_1695 (O_1695,N_28830,N_26309);
nor UO_1696 (O_1696,N_27051,N_26628);
or UO_1697 (O_1697,N_29581,N_27201);
nand UO_1698 (O_1698,N_29552,N_25265);
nor UO_1699 (O_1699,N_27378,N_26075);
or UO_1700 (O_1700,N_26683,N_25403);
or UO_1701 (O_1701,N_25719,N_25294);
and UO_1702 (O_1702,N_29608,N_25698);
nand UO_1703 (O_1703,N_25528,N_29806);
and UO_1704 (O_1704,N_29752,N_27483);
nor UO_1705 (O_1705,N_27136,N_27380);
nor UO_1706 (O_1706,N_28620,N_27924);
nor UO_1707 (O_1707,N_29269,N_28407);
nor UO_1708 (O_1708,N_28628,N_26728);
nor UO_1709 (O_1709,N_28929,N_27014);
nand UO_1710 (O_1710,N_28603,N_26775);
nand UO_1711 (O_1711,N_25256,N_26251);
nor UO_1712 (O_1712,N_25851,N_25396);
or UO_1713 (O_1713,N_28544,N_25463);
xnor UO_1714 (O_1714,N_28432,N_27553);
xor UO_1715 (O_1715,N_28961,N_25577);
and UO_1716 (O_1716,N_27422,N_27542);
or UO_1717 (O_1717,N_28310,N_26963);
or UO_1718 (O_1718,N_29894,N_26727);
nor UO_1719 (O_1719,N_28296,N_26138);
xnor UO_1720 (O_1720,N_28421,N_29242);
and UO_1721 (O_1721,N_29165,N_28494);
nor UO_1722 (O_1722,N_27088,N_26747);
or UO_1723 (O_1723,N_26282,N_25876);
and UO_1724 (O_1724,N_29947,N_25172);
or UO_1725 (O_1725,N_29487,N_26135);
nand UO_1726 (O_1726,N_28247,N_25967);
nand UO_1727 (O_1727,N_25807,N_29408);
or UO_1728 (O_1728,N_29613,N_26882);
nand UO_1729 (O_1729,N_28328,N_28975);
nand UO_1730 (O_1730,N_27649,N_27372);
nand UO_1731 (O_1731,N_25943,N_27240);
nand UO_1732 (O_1732,N_29021,N_28203);
xnor UO_1733 (O_1733,N_27896,N_25497);
nor UO_1734 (O_1734,N_27676,N_27889);
nand UO_1735 (O_1735,N_26257,N_26150);
nor UO_1736 (O_1736,N_29063,N_25667);
nor UO_1737 (O_1737,N_29579,N_27029);
or UO_1738 (O_1738,N_26288,N_25963);
nand UO_1739 (O_1739,N_25934,N_25969);
or UO_1740 (O_1740,N_28295,N_28713);
nand UO_1741 (O_1741,N_27063,N_26095);
or UO_1742 (O_1742,N_27957,N_25769);
nand UO_1743 (O_1743,N_28573,N_28466);
and UO_1744 (O_1744,N_25942,N_28371);
nor UO_1745 (O_1745,N_27754,N_29667);
xnor UO_1746 (O_1746,N_26700,N_26530);
nor UO_1747 (O_1747,N_27587,N_25945);
nand UO_1748 (O_1748,N_27488,N_29919);
nor UO_1749 (O_1749,N_25966,N_26069);
nand UO_1750 (O_1750,N_26858,N_29787);
or UO_1751 (O_1751,N_25164,N_27745);
nand UO_1752 (O_1752,N_27965,N_29900);
nor UO_1753 (O_1753,N_27543,N_27132);
nand UO_1754 (O_1754,N_25803,N_26173);
nand UO_1755 (O_1755,N_26120,N_25733);
nand UO_1756 (O_1756,N_26879,N_26918);
nand UO_1757 (O_1757,N_26658,N_27780);
and UO_1758 (O_1758,N_25715,N_29014);
nand UO_1759 (O_1759,N_25390,N_27887);
or UO_1760 (O_1760,N_29501,N_28288);
and UO_1761 (O_1761,N_26244,N_26301);
and UO_1762 (O_1762,N_29008,N_26731);
and UO_1763 (O_1763,N_27058,N_28616);
or UO_1764 (O_1764,N_28150,N_28930);
nand UO_1765 (O_1765,N_28006,N_28315);
and UO_1766 (O_1766,N_27392,N_26892);
nor UO_1767 (O_1767,N_27067,N_25309);
nor UO_1768 (O_1768,N_29333,N_25569);
and UO_1769 (O_1769,N_26430,N_27349);
and UO_1770 (O_1770,N_29872,N_27902);
nand UO_1771 (O_1771,N_28263,N_27959);
and UO_1772 (O_1772,N_25842,N_29491);
nand UO_1773 (O_1773,N_28514,N_26850);
or UO_1774 (O_1774,N_26682,N_26331);
xor UO_1775 (O_1775,N_28270,N_28397);
nand UO_1776 (O_1776,N_25150,N_26837);
or UO_1777 (O_1777,N_28669,N_28219);
nor UO_1778 (O_1778,N_28089,N_28241);
nor UO_1779 (O_1779,N_26398,N_25760);
nand UO_1780 (O_1780,N_29039,N_27979);
and UO_1781 (O_1781,N_28936,N_26415);
nor UO_1782 (O_1782,N_27904,N_28363);
nor UO_1783 (O_1783,N_26810,N_25538);
nor UO_1784 (O_1784,N_26684,N_27033);
or UO_1785 (O_1785,N_26807,N_29149);
and UO_1786 (O_1786,N_28305,N_28048);
xor UO_1787 (O_1787,N_29362,N_29176);
and UO_1788 (O_1788,N_29310,N_27787);
or UO_1789 (O_1789,N_29146,N_28655);
nand UO_1790 (O_1790,N_26923,N_29106);
and UO_1791 (O_1791,N_27873,N_25140);
or UO_1792 (O_1792,N_27231,N_26432);
or UO_1793 (O_1793,N_26358,N_26117);
and UO_1794 (O_1794,N_27657,N_26937);
nor UO_1795 (O_1795,N_26800,N_28978);
and UO_1796 (O_1796,N_26504,N_29389);
or UO_1797 (O_1797,N_27080,N_29686);
nand UO_1798 (O_1798,N_29715,N_26820);
or UO_1799 (O_1799,N_29488,N_29498);
or UO_1800 (O_1800,N_26067,N_27421);
xnor UO_1801 (O_1801,N_25218,N_26583);
and UO_1802 (O_1802,N_26050,N_25054);
nor UO_1803 (O_1803,N_29435,N_28095);
nor UO_1804 (O_1804,N_27505,N_25332);
and UO_1805 (O_1805,N_25990,N_29058);
and UO_1806 (O_1806,N_28010,N_27269);
or UO_1807 (O_1807,N_26019,N_28230);
and UO_1808 (O_1808,N_26953,N_25204);
nand UO_1809 (O_1809,N_26472,N_27749);
or UO_1810 (O_1810,N_27197,N_28245);
nand UO_1811 (O_1811,N_25907,N_28553);
nor UO_1812 (O_1812,N_28265,N_29247);
or UO_1813 (O_1813,N_26108,N_27683);
nor UO_1814 (O_1814,N_29640,N_29463);
or UO_1815 (O_1815,N_29326,N_28057);
nor UO_1816 (O_1816,N_27531,N_28913);
or UO_1817 (O_1817,N_25728,N_27807);
and UO_1818 (O_1818,N_29015,N_25782);
or UO_1819 (O_1819,N_26326,N_29354);
or UO_1820 (O_1820,N_26817,N_26989);
or UO_1821 (O_1821,N_26258,N_25336);
nand UO_1822 (O_1822,N_29496,N_28101);
nand UO_1823 (O_1823,N_26268,N_28225);
or UO_1824 (O_1824,N_26024,N_26749);
and UO_1825 (O_1825,N_29390,N_29215);
or UO_1826 (O_1826,N_28914,N_27958);
nor UO_1827 (O_1827,N_29436,N_26641);
and UO_1828 (O_1828,N_26416,N_25020);
nor UO_1829 (O_1829,N_28044,N_25062);
nor UO_1830 (O_1830,N_27097,N_29838);
xor UO_1831 (O_1831,N_26572,N_27230);
nor UO_1832 (O_1832,N_28007,N_26121);
or UO_1833 (O_1833,N_28195,N_27903);
nor UO_1834 (O_1834,N_28235,N_28757);
or UO_1835 (O_1835,N_27738,N_28040);
nand UO_1836 (O_1836,N_27388,N_27154);
nand UO_1837 (O_1837,N_27339,N_27475);
or UO_1838 (O_1838,N_28384,N_27134);
nor UO_1839 (O_1839,N_25658,N_27100);
nand UO_1840 (O_1840,N_28274,N_28480);
and UO_1841 (O_1841,N_25816,N_26094);
or UO_1842 (O_1842,N_25298,N_26284);
and UO_1843 (O_1843,N_25825,N_27628);
nand UO_1844 (O_1844,N_29870,N_27312);
and UO_1845 (O_1845,N_27954,N_25526);
and UO_1846 (O_1846,N_29876,N_29653);
or UO_1847 (O_1847,N_27602,N_27366);
nand UO_1848 (O_1848,N_28298,N_25022);
or UO_1849 (O_1849,N_26735,N_25470);
or UO_1850 (O_1850,N_25479,N_28518);
nor UO_1851 (O_1851,N_29539,N_29013);
nor UO_1852 (O_1852,N_29384,N_26037);
xnor UO_1853 (O_1853,N_27845,N_25285);
nand UO_1854 (O_1854,N_27391,N_29402);
and UO_1855 (O_1855,N_26020,N_25325);
and UO_1856 (O_1856,N_27652,N_27967);
and UO_1857 (O_1857,N_29160,N_25939);
and UO_1858 (O_1858,N_29678,N_28446);
or UO_1859 (O_1859,N_26703,N_26938);
nand UO_1860 (O_1860,N_27160,N_26816);
nand UO_1861 (O_1861,N_28920,N_25095);
xnor UO_1862 (O_1862,N_29606,N_26348);
nand UO_1863 (O_1863,N_27943,N_27558);
and UO_1864 (O_1864,N_25355,N_26178);
or UO_1865 (O_1865,N_29728,N_28002);
nor UO_1866 (O_1866,N_26930,N_25014);
nand UO_1867 (O_1867,N_29444,N_28068);
and UO_1868 (O_1868,N_25085,N_29875);
and UO_1869 (O_1869,N_29166,N_26562);
nand UO_1870 (O_1870,N_25743,N_29459);
nor UO_1871 (O_1871,N_27931,N_28598);
xor UO_1872 (O_1872,N_26063,N_26519);
nand UO_1873 (O_1873,N_29591,N_27864);
nand UO_1874 (O_1874,N_28809,N_28958);
nand UO_1875 (O_1875,N_29002,N_26633);
and UO_1876 (O_1876,N_27092,N_28490);
nor UO_1877 (O_1877,N_25829,N_25672);
nor UO_1878 (O_1878,N_29394,N_25375);
nand UO_1879 (O_1879,N_25888,N_28159);
and UO_1880 (O_1880,N_27620,N_27668);
nand UO_1881 (O_1881,N_28845,N_28345);
and UO_1882 (O_1882,N_29108,N_27334);
and UO_1883 (O_1883,N_25666,N_27520);
nor UO_1884 (O_1884,N_27117,N_29373);
and UO_1885 (O_1885,N_29078,N_26514);
nor UO_1886 (O_1886,N_28956,N_26674);
nand UO_1887 (O_1887,N_27280,N_29849);
and UO_1888 (O_1888,N_27476,N_25959);
and UO_1889 (O_1889,N_27909,N_25866);
xnor UO_1890 (O_1890,N_28736,N_29313);
nand UO_1891 (O_1891,N_27837,N_27383);
or UO_1892 (O_1892,N_27135,N_29255);
and UO_1893 (O_1893,N_27227,N_28854);
xor UO_1894 (O_1894,N_27512,N_26617);
and UO_1895 (O_1895,N_29023,N_27748);
nor UO_1896 (O_1896,N_27524,N_25307);
nor UO_1897 (O_1897,N_27723,N_28562);
nor UO_1898 (O_1898,N_28231,N_26216);
or UO_1899 (O_1899,N_29990,N_26585);
or UO_1900 (O_1900,N_28820,N_26794);
or UO_1901 (O_1901,N_28998,N_29748);
nand UO_1902 (O_1902,N_28078,N_28459);
or UO_1903 (O_1903,N_28721,N_26411);
nor UO_1904 (O_1904,N_27305,N_27863);
nand UO_1905 (O_1905,N_25137,N_28516);
or UO_1906 (O_1906,N_25413,N_28001);
and UO_1907 (O_1907,N_28505,N_26924);
nor UO_1908 (O_1908,N_26332,N_26199);
xor UO_1909 (O_1909,N_26647,N_26291);
nand UO_1910 (O_1910,N_28320,N_27122);
or UO_1911 (O_1911,N_27589,N_28564);
nor UO_1912 (O_1912,N_29267,N_26494);
or UO_1913 (O_1913,N_25360,N_29649);
nor UO_1914 (O_1914,N_29851,N_26099);
nand UO_1915 (O_1915,N_25003,N_26681);
xor UO_1916 (O_1916,N_26236,N_27336);
and UO_1917 (O_1917,N_26948,N_26846);
and UO_1918 (O_1918,N_25043,N_26306);
xnor UO_1919 (O_1919,N_29136,N_26506);
nand UO_1920 (O_1920,N_29931,N_25047);
xor UO_1921 (O_1921,N_26159,N_29570);
and UO_1922 (O_1922,N_28360,N_26065);
or UO_1923 (O_1923,N_25476,N_26639);
nor UO_1924 (O_1924,N_28500,N_25643);
and UO_1925 (O_1925,N_29152,N_29066);
or UO_1926 (O_1926,N_25617,N_27677);
xnor UO_1927 (O_1927,N_26764,N_29700);
and UO_1928 (O_1928,N_25153,N_28456);
and UO_1929 (O_1929,N_28492,N_28537);
nor UO_1930 (O_1930,N_26480,N_26902);
nand UO_1931 (O_1931,N_25602,N_26840);
nor UO_1932 (O_1932,N_26328,N_28258);
xor UO_1933 (O_1933,N_25744,N_29916);
xnor UO_1934 (O_1934,N_27960,N_26667);
and UO_1935 (O_1935,N_29443,N_27574);
and UO_1936 (O_1936,N_29556,N_25353);
nor UO_1937 (O_1937,N_26009,N_29128);
and UO_1938 (O_1938,N_26802,N_29696);
nor UO_1939 (O_1939,N_26738,N_28663);
xnor UO_1940 (O_1940,N_25676,N_25391);
xnor UO_1941 (O_1941,N_27680,N_25320);
nor UO_1942 (O_1942,N_27850,N_28003);
xnor UO_1943 (O_1943,N_26333,N_28653);
nand UO_1944 (O_1944,N_26958,N_28703);
and UO_1945 (O_1945,N_28058,N_27606);
and UO_1946 (O_1946,N_25237,N_29060);
nor UO_1947 (O_1947,N_25962,N_25060);
nand UO_1948 (O_1948,N_25251,N_25475);
and UO_1949 (O_1949,N_26316,N_26987);
and UO_1950 (O_1950,N_25809,N_28970);
nor UO_1951 (O_1951,N_26195,N_27386);
or UO_1952 (O_1952,N_28762,N_27828);
nor UO_1953 (O_1953,N_26525,N_29571);
or UO_1954 (O_1954,N_26458,N_29210);
nor UO_1955 (O_1955,N_28904,N_25005);
and UO_1956 (O_1956,N_25865,N_27727);
or UO_1957 (O_1957,N_28887,N_29549);
and UO_1958 (O_1958,N_26677,N_25278);
nor UO_1959 (O_1959,N_29850,N_26342);
or UO_1960 (O_1960,N_26870,N_29694);
nor UO_1961 (O_1961,N_25350,N_28153);
or UO_1962 (O_1962,N_28953,N_25642);
or UO_1963 (O_1963,N_25824,N_26499);
nand UO_1964 (O_1964,N_27795,N_29070);
or UO_1965 (O_1965,N_26325,N_27013);
and UO_1966 (O_1966,N_29577,N_25427);
or UO_1967 (O_1967,N_28286,N_25008);
or UO_1968 (O_1968,N_29305,N_26554);
and UO_1969 (O_1969,N_25794,N_26241);
and UO_1970 (O_1970,N_29143,N_25024);
and UO_1971 (O_1971,N_25415,N_27427);
or UO_1972 (O_1972,N_28198,N_26381);
xor UO_1973 (O_1973,N_29054,N_29294);
xor UO_1974 (O_1974,N_28313,N_27437);
nand UO_1975 (O_1975,N_29211,N_27756);
and UO_1976 (O_1976,N_27111,N_29925);
or UO_1977 (O_1977,N_29031,N_28212);
or UO_1978 (O_1978,N_29587,N_29403);
nand UO_1979 (O_1979,N_28107,N_29704);
xnor UO_1980 (O_1980,N_26642,N_25016);
xor UO_1981 (O_1981,N_29378,N_29886);
or UO_1982 (O_1982,N_28652,N_25954);
xor UO_1983 (O_1983,N_27566,N_28526);
xnor UO_1984 (O_1984,N_26689,N_27499);
nor UO_1985 (O_1985,N_27415,N_25321);
or UO_1986 (O_1986,N_25440,N_28539);
and UO_1987 (O_1987,N_25736,N_25190);
and UO_1988 (O_1988,N_27768,N_25820);
or UO_1989 (O_1989,N_28177,N_25057);
or UO_1990 (O_1990,N_28043,N_26049);
and UO_1991 (O_1991,N_26368,N_28707);
or UO_1992 (O_1992,N_29418,N_28814);
xor UO_1993 (O_1993,N_29811,N_27469);
or UO_1994 (O_1994,N_29937,N_29358);
or UO_1995 (O_1995,N_26788,N_27642);
xor UO_1996 (O_1996,N_27404,N_28879);
and UO_1997 (O_1997,N_29633,N_27742);
and UO_1998 (O_1998,N_25797,N_26053);
nor UO_1999 (O_1999,N_29940,N_26715);
nand UO_2000 (O_2000,N_26335,N_29770);
nor UO_2001 (O_2001,N_28684,N_27482);
and UO_2002 (O_2002,N_29980,N_26496);
nor UO_2003 (O_2003,N_29494,N_26197);
nor UO_2004 (O_2004,N_27291,N_25259);
nor UO_2005 (O_2005,N_27784,N_27374);
or UO_2006 (O_2006,N_27951,N_28533);
nand UO_2007 (O_2007,N_27030,N_28995);
nor UO_2008 (O_2008,N_29529,N_29914);
nor UO_2009 (O_2009,N_27760,N_27583);
nand UO_2010 (O_2010,N_27487,N_29629);
xor UO_2011 (O_2011,N_29736,N_28928);
nor UO_2012 (O_2012,N_25679,N_26905);
or UO_2013 (O_2013,N_29970,N_29433);
nand UO_2014 (O_2014,N_27236,N_28902);
nand UO_2015 (O_2015,N_25938,N_27244);
and UO_2016 (O_2016,N_25178,N_25471);
and UO_2017 (O_2017,N_27143,N_25853);
nand UO_2018 (O_2018,N_26805,N_29644);
and UO_2019 (O_2019,N_25725,N_26551);
or UO_2020 (O_2020,N_27968,N_26809);
nor UO_2021 (O_2021,N_28795,N_26030);
and UO_2022 (O_2022,N_27420,N_27179);
and UO_2023 (O_2023,N_25953,N_25439);
and UO_2024 (O_2024,N_27060,N_25878);
and UO_2025 (O_2025,N_27338,N_25230);
nor UO_2026 (O_2026,N_26484,N_28555);
nor UO_2027 (O_2027,N_26919,N_29188);
or UO_2028 (O_2028,N_25831,N_28213);
or UO_2029 (O_2029,N_29006,N_28880);
and UO_2030 (O_2030,N_27397,N_29224);
nor UO_2031 (O_2031,N_29312,N_26664);
nor UO_2032 (O_2032,N_26144,N_26452);
nand UO_2033 (O_2033,N_28702,N_29657);
nand UO_2034 (O_2034,N_27004,N_29087);
nor UO_2035 (O_2035,N_29650,N_29668);
and UO_2036 (O_2036,N_28862,N_28094);
nand UO_2037 (O_2037,N_28837,N_27455);
xor UO_2038 (O_2038,N_29474,N_29710);
or UO_2039 (O_2039,N_27855,N_25978);
nand UO_2040 (O_2040,N_28067,N_29823);
xnor UO_2041 (O_2041,N_28660,N_25923);
nor UO_2042 (O_2042,N_28437,N_25247);
or UO_2043 (O_2043,N_28868,N_28351);
nand UO_2044 (O_2044,N_27018,N_28876);
and UO_2045 (O_2045,N_26043,N_27379);
xnor UO_2046 (O_2046,N_28711,N_25105);
nand UO_2047 (O_2047,N_27981,N_25625);
xor UO_2048 (O_2048,N_29026,N_28893);
xor UO_2049 (O_2049,N_28615,N_26096);
nor UO_2050 (O_2050,N_28133,N_27342);
or UO_2051 (O_2051,N_28869,N_29053);
nor UO_2052 (O_2052,N_29505,N_29288);
or UO_2053 (O_2053,N_25754,N_26259);
and UO_2054 (O_2054,N_28989,N_27083);
or UO_2055 (O_2055,N_27980,N_28392);
nand UO_2056 (O_2056,N_27513,N_27802);
or UO_2057 (O_2057,N_29417,N_29183);
and UO_2058 (O_2058,N_27514,N_25300);
nand UO_2059 (O_2059,N_29101,N_25977);
or UO_2060 (O_2060,N_29727,N_27808);
or UO_2061 (O_2061,N_27561,N_28454);
or UO_2062 (O_2062,N_26187,N_29833);
nand UO_2063 (O_2063,N_29744,N_25115);
nand UO_2064 (O_2064,N_29987,N_25594);
or UO_2065 (O_2065,N_27319,N_25640);
nand UO_2066 (O_2066,N_26175,N_29185);
nor UO_2067 (O_2067,N_27133,N_29080);
nand UO_2068 (O_2068,N_29908,N_29933);
xnor UO_2069 (O_2069,N_26957,N_27170);
and UO_2070 (O_2070,N_26592,N_25871);
and UO_2071 (O_2071,N_27687,N_26102);
nor UO_2072 (O_2072,N_28339,N_25855);
nand UO_2073 (O_2073,N_27966,N_28268);
and UO_2074 (O_2074,N_26038,N_28134);
or UO_2075 (O_2075,N_25905,N_29651);
or UO_2076 (O_2076,N_25378,N_25763);
xor UO_2077 (O_2077,N_29306,N_27554);
nor UO_2078 (O_2078,N_25565,N_26501);
and UO_2079 (O_2079,N_25406,N_25123);
nand UO_2080 (O_2080,N_27289,N_29905);
and UO_2081 (O_2081,N_27729,N_27186);
or UO_2082 (O_2082,N_25101,N_29885);
and UO_2083 (O_2083,N_26921,N_26436);
and UO_2084 (O_2084,N_28662,N_27222);
and UO_2085 (O_2085,N_29365,N_28129);
nor UO_2086 (O_2086,N_26917,N_26719);
nor UO_2087 (O_2087,N_26055,N_27836);
and UO_2088 (O_2088,N_29574,N_26529);
and UO_2089 (O_2089,N_28349,N_29714);
xor UO_2090 (O_2090,N_25791,N_26575);
and UO_2091 (O_2091,N_28934,N_27734);
and UO_2092 (O_2092,N_27447,N_25448);
and UO_2093 (O_2093,N_28460,N_26211);
or UO_2094 (O_2094,N_28839,N_28425);
and UO_2095 (O_2095,N_25374,N_28791);
nand UO_2096 (O_2096,N_25425,N_27519);
nand UO_2097 (O_2097,N_26594,N_25426);
and UO_2098 (O_2098,N_25469,N_26367);
and UO_2099 (O_2099,N_27443,N_25087);
and UO_2100 (O_2100,N_26136,N_29437);
nor UO_2101 (O_2101,N_29091,N_28982);
nand UO_2102 (O_2102,N_29214,N_28666);
and UO_2103 (O_2103,N_28855,N_29913);
or UO_2104 (O_2104,N_29829,N_25387);
xnor UO_2105 (O_2105,N_28599,N_28005);
or UO_2106 (O_2106,N_25531,N_25912);
nand UO_2107 (O_2107,N_28343,N_28082);
and UO_2108 (O_2108,N_25618,N_25714);
nand UO_2109 (O_2109,N_28042,N_29400);
nor UO_2110 (O_2110,N_25957,N_25985);
or UO_2111 (O_2111,N_27915,N_25100);
nand UO_2112 (O_2112,N_25659,N_27363);
nor UO_2113 (O_2113,N_26225,N_29954);
and UO_2114 (O_2114,N_29457,N_28922);
nand UO_2115 (O_2115,N_25031,N_27998);
nand UO_2116 (O_2116,N_27594,N_27985);
nand UO_2117 (O_2117,N_28905,N_29622);
or UO_2118 (O_2118,N_26243,N_28629);
and UO_2119 (O_2119,N_28842,N_29767);
nor UO_2120 (O_2120,N_29955,N_27169);
or UO_2121 (O_2121,N_26966,N_26210);
nand UO_2122 (O_2122,N_25810,N_25873);
and UO_2123 (O_2123,N_27541,N_28720);
nand UO_2124 (O_2124,N_26610,N_28173);
nor UO_2125 (O_2125,N_28997,N_28836);
xor UO_2126 (O_2126,N_28332,N_25198);
nor UO_2127 (O_2127,N_27123,N_29923);
nand UO_2128 (O_2128,N_25168,N_25779);
or UO_2129 (O_2129,N_28949,N_26276);
or UO_2130 (O_2130,N_29995,N_27070);
nor UO_2131 (O_2131,N_26364,N_29486);
nand UO_2132 (O_2132,N_28444,N_28701);
nand UO_2133 (O_2133,N_28530,N_26320);
nor UO_2134 (O_2134,N_29901,N_26502);
and UO_2135 (O_2135,N_26034,N_25474);
xor UO_2136 (O_2136,N_26811,N_29187);
or UO_2137 (O_2137,N_26450,N_25680);
nand UO_2138 (O_2138,N_28749,N_27588);
nor UO_2139 (O_2139,N_25048,N_29853);
nand UO_2140 (O_2140,N_27719,N_29926);
nor UO_2141 (O_2141,N_27480,N_25800);
or UO_2142 (O_2142,N_26372,N_25948);
nor UO_2143 (O_2143,N_25846,N_27082);
or UO_2144 (O_2144,N_27394,N_27194);
or UO_2145 (O_2145,N_28569,N_25317);
xnor UO_2146 (O_2146,N_25506,N_25245);
and UO_2147 (O_2147,N_26433,N_29366);
and UO_2148 (O_2148,N_25891,N_25560);
nor UO_2149 (O_2149,N_28161,N_28865);
or UO_2150 (O_2150,N_27832,N_26428);
nor UO_2151 (O_2151,N_28843,N_27851);
or UO_2152 (O_2152,N_29226,N_29877);
nor UO_2153 (O_2153,N_29168,N_25841);
or UO_2154 (O_2154,N_27304,N_27914);
or UO_2155 (O_2155,N_29334,N_25596);
nand UO_2156 (O_2156,N_25895,N_25399);
nor UO_2157 (O_2157,N_26232,N_26561);
nand UO_2158 (O_2158,N_26982,N_26927);
or UO_2159 (O_2159,N_28477,N_29673);
or UO_2160 (O_2160,N_27880,N_26950);
nor UO_2161 (O_2161,N_25879,N_27955);
nand UO_2162 (O_2162,N_28538,N_28210);
nor UO_2163 (O_2163,N_26362,N_25296);
and UO_2164 (O_2164,N_27028,N_28206);
or UO_2165 (O_2165,N_28623,N_27969);
nand UO_2166 (O_2166,N_27439,N_27932);
or UO_2167 (O_2167,N_27757,N_26272);
and UO_2168 (O_2168,N_25568,N_28075);
xnor UO_2169 (O_2169,N_25777,N_27798);
and UO_2170 (O_2170,N_27096,N_26080);
and UO_2171 (O_2171,N_25102,N_29703);
or UO_2172 (O_2172,N_26756,N_29105);
or UO_2173 (O_2173,N_26464,N_29276);
and UO_2174 (O_2174,N_27454,N_26773);
nor UO_2175 (O_2175,N_27877,N_27329);
or UO_2176 (O_2176,N_28649,N_27846);
or UO_2177 (O_2177,N_26321,N_26630);
xnor UO_2178 (O_2178,N_27152,N_27659);
or UO_2179 (O_2179,N_27944,N_25232);
xnor UO_2180 (O_2180,N_26497,N_29047);
or UO_2181 (O_2181,N_29912,N_26461);
nand UO_2182 (O_2182,N_27090,N_25380);
and UO_2183 (O_2183,N_29743,N_27371);
and UO_2184 (O_2184,N_28595,N_25723);
nor UO_2185 (O_2185,N_27978,N_26705);
or UO_2186 (O_2186,N_25956,N_27130);
or UO_2187 (O_2187,N_28878,N_27616);
nand UO_2188 (O_2188,N_29115,N_29835);
and UO_2189 (O_2189,N_28329,N_25257);
nand UO_2190 (O_2190,N_27367,N_28808);
nand UO_2191 (O_2191,N_27655,N_29239);
nand UO_2192 (O_2192,N_28338,N_28131);
xnor UO_2193 (O_2193,N_25508,N_27145);
nand UO_2194 (O_2194,N_28769,N_29803);
and UO_2195 (O_2195,N_29193,N_26194);
nand UO_2196 (O_2196,N_27204,N_25929);
and UO_2197 (O_2197,N_28951,N_29625);
and UO_2198 (O_2198,N_25385,N_29532);
nand UO_2199 (O_2199,N_25455,N_25682);
and UO_2200 (O_2200,N_28919,N_25510);
or UO_2201 (O_2201,N_28112,N_27800);
nor UO_2202 (O_2202,N_29422,N_25813);
and UO_2203 (O_2203,N_27387,N_27671);
nor UO_2204 (O_2204,N_28027,N_27419);
nand UO_2205 (O_2205,N_27085,N_26396);
and UO_2206 (O_2206,N_27595,N_28341);
or UO_2207 (O_2207,N_26343,N_28083);
xor UO_2208 (O_2208,N_25428,N_25677);
and UO_2209 (O_2209,N_28675,N_29368);
and UO_2210 (O_2210,N_28592,N_26612);
nand UO_2211 (O_2211,N_25009,N_26707);
nor UO_2212 (O_2212,N_28489,N_26900);
xor UO_2213 (O_2213,N_28013,N_27278);
or UO_2214 (O_2214,N_28954,N_26828);
nor UO_2215 (O_2215,N_26651,N_26380);
nor UO_2216 (O_2216,N_26214,N_28659);
xor UO_2217 (O_2217,N_26391,N_28030);
xor UO_2218 (O_2218,N_27162,N_26706);
nand UO_2219 (O_2219,N_25313,N_25133);
nand UO_2220 (O_2220,N_28080,N_25685);
nor UO_2221 (O_2221,N_28716,N_27465);
nor UO_2222 (O_2222,N_28907,N_27228);
or UO_2223 (O_2223,N_25383,N_26407);
nor UO_2224 (O_2224,N_29665,N_25120);
xor UO_2225 (O_2225,N_27888,N_25224);
nor UO_2226 (O_2226,N_29848,N_25273);
or UO_2227 (O_2227,N_29117,N_25513);
or UO_2228 (O_2228,N_29454,N_29538);
or UO_2229 (O_2229,N_26721,N_25151);
nor UO_2230 (O_2230,N_26935,N_25629);
nor UO_2231 (O_2231,N_28626,N_28116);
nor UO_2232 (O_2232,N_29121,N_25242);
nor UO_2233 (O_2233,N_27761,N_27148);
or UO_2234 (O_2234,N_26590,N_25849);
or UO_2235 (O_2235,N_29961,N_27631);
xnor UO_2236 (O_2236,N_25932,N_27664);
xnor UO_2237 (O_2237,N_29052,N_28266);
nand UO_2238 (O_2238,N_27287,N_26626);
nand UO_2239 (O_2239,N_25119,N_28366);
nor UO_2240 (O_2240,N_29139,N_26524);
nor UO_2241 (O_2241,N_28051,N_27373);
and UO_2242 (O_2242,N_25868,N_26256);
nand UO_2243 (O_2243,N_27036,N_25142);
nand UO_2244 (O_2244,N_27670,N_29140);
nor UO_2245 (O_2245,N_27755,N_28036);
nor UO_2246 (O_2246,N_26219,N_28055);
or UO_2247 (O_2247,N_29815,N_29237);
nand UO_2248 (O_2248,N_27208,N_27253);
nand UO_2249 (O_2249,N_27436,N_28347);
nand UO_2250 (O_2250,N_29642,N_28223);
nand UO_2251 (O_2251,N_27822,N_25205);
xnor UO_2252 (O_2252,N_26618,N_28482);
and UO_2253 (O_2253,N_25250,N_28602);
nor UO_2254 (O_2254,N_29359,N_25181);
nor UO_2255 (O_2255,N_29148,N_29565);
nor UO_2256 (O_2256,N_28309,N_25405);
and UO_2257 (O_2257,N_28491,N_25166);
or UO_2258 (O_2258,N_26673,N_28831);
xnor UO_2259 (O_2259,N_29812,N_25635);
or UO_2260 (O_2260,N_27689,N_29175);
and UO_2261 (O_2261,N_25826,N_27698);
nor UO_2262 (O_2262,N_28909,N_27408);
nor UO_2263 (O_2263,N_29773,N_29221);
nand UO_2264 (O_2264,N_25319,N_26402);
nor UO_2265 (O_2265,N_28709,N_26158);
or UO_2266 (O_2266,N_26736,N_26114);
and UO_2267 (O_2267,N_26429,N_25608);
xnor UO_2268 (O_2268,N_29802,N_28963);
or UO_2269 (O_2269,N_27331,N_25522);
nor UO_2270 (O_2270,N_27248,N_28700);
and UO_2271 (O_2271,N_27753,N_28099);
or UO_2272 (O_2272,N_29871,N_27435);
and UO_2273 (O_2273,N_25481,N_26815);
xnor UO_2274 (O_2274,N_25299,N_28864);
and UO_2275 (O_2275,N_29317,N_25670);
or UO_2276 (O_2276,N_27276,N_25920);
nor UO_2277 (O_2277,N_29960,N_26176);
and UO_2278 (O_2278,N_27952,N_26714);
nor UO_2279 (O_2279,N_25854,N_29756);
or UO_2280 (O_2280,N_28162,N_26570);
nor UO_2281 (O_2281,N_26238,N_27700);
nand UO_2282 (O_2282,N_29679,N_25433);
nor UO_2283 (O_2283,N_25770,N_25436);
nand UO_2284 (O_2284,N_28066,N_28656);
or UO_2285 (O_2285,N_27251,N_25590);
or UO_2286 (O_2286,N_25145,N_25114);
xor UO_2287 (O_2287,N_25663,N_29303);
or UO_2288 (O_2288,N_28871,N_28370);
nor UO_2289 (O_2289,N_25480,N_28468);
nand UO_2290 (O_2290,N_26760,N_26552);
nor UO_2291 (O_2291,N_25523,N_29766);
or UO_2292 (O_2292,N_25029,N_26008);
nor UO_2293 (O_2293,N_29603,N_29460);
xnor UO_2294 (O_2294,N_25839,N_25908);
nand UO_2295 (O_2295,N_29985,N_26732);
and UO_2296 (O_2296,N_29441,N_28243);
nor UO_2297 (O_2297,N_25065,N_25681);
or UO_2298 (O_2298,N_29482,N_25570);
nand UO_2299 (O_2299,N_26260,N_27261);
nor UO_2300 (O_2300,N_25217,N_26156);
and UO_2301 (O_2301,N_28119,N_29203);
xor UO_2302 (O_2302,N_27346,N_27653);
and UO_2303 (O_2303,N_28272,N_25460);
or UO_2304 (O_2304,N_26620,N_27150);
nand UO_2305 (O_2305,N_28359,N_25131);
xnor UO_2306 (O_2306,N_26964,N_28130);
or UO_2307 (O_2307,N_29507,N_29515);
nand UO_2308 (O_2308,N_26799,N_27247);
or UO_2309 (O_2309,N_26926,N_27629);
xnor UO_2310 (O_2310,N_27971,N_27140);
nand UO_2311 (O_2311,N_29939,N_28383);
nand UO_2312 (O_2312,N_28074,N_27486);
nor UO_2313 (O_2313,N_29729,N_25792);
nand UO_2314 (O_2314,N_28596,N_26894);
nor UO_2315 (O_2315,N_25185,N_28046);
nor UO_2316 (O_2316,N_28717,N_26741);
nor UO_2317 (O_2317,N_28829,N_25361);
and UO_2318 (O_2318,N_27497,N_27610);
nor UO_2319 (O_2319,N_25229,N_25039);
nor UO_2320 (O_2320,N_25935,N_26208);
and UO_2321 (O_2321,N_29594,N_26600);
or UO_2322 (O_2322,N_26228,N_26071);
nand UO_2323 (O_2323,N_25650,N_25489);
and UO_2324 (O_2324,N_27323,N_29621);
nor UO_2325 (O_2325,N_28474,N_25222);
or UO_2326 (O_2326,N_27772,N_26779);
nand UO_2327 (O_2327,N_27713,N_27232);
nand UO_2328 (O_2328,N_29025,N_26418);
nand UO_2329 (O_2329,N_29287,N_27041);
or UO_2330 (O_2330,N_26711,N_27638);
and UO_2331 (O_2331,N_25783,N_29493);
xor UO_2332 (O_2332,N_29124,N_28056);
nor UO_2333 (O_2333,N_28093,N_28962);
or UO_2334 (O_2334,N_28166,N_28260);
xnor UO_2335 (O_2335,N_29566,N_28128);
and UO_2336 (O_2336,N_27149,N_27578);
xor UO_2337 (O_2337,N_28254,N_29731);
nor UO_2338 (O_2338,N_25135,N_26013);
nor UO_2339 (O_2339,N_28850,N_27970);
nand UO_2340 (O_2340,N_29687,N_27178);
nand UO_2341 (O_2341,N_28322,N_26188);
xor UO_2342 (O_2342,N_27301,N_28634);
nor UO_2343 (O_2343,N_26766,N_26234);
or UO_2344 (O_2344,N_29693,N_26092);
nor UO_2345 (O_2345,N_25581,N_29839);
nand UO_2346 (O_2346,N_28877,N_26743);
nand UO_2347 (O_2347,N_28774,N_29887);
or UO_2348 (O_2348,N_26387,N_29573);
and UO_2349 (O_2349,N_29286,N_29102);
and UO_2350 (O_2350,N_28312,N_28822);
nor UO_2351 (O_2351,N_27611,N_28256);
or UO_2352 (O_2352,N_25359,N_25179);
or UO_2353 (O_2353,N_27910,N_25606);
or UO_2354 (O_2354,N_26615,N_25623);
or UO_2355 (O_2355,N_28873,N_26133);
or UO_2356 (O_2356,N_26675,N_26833);
nor UO_2357 (O_2357,N_26283,N_26792);
or UO_2358 (O_2358,N_27516,N_27009);
nand UO_2359 (O_2359,N_26147,N_28430);
nand UO_2360 (O_2360,N_26351,N_29797);
or UO_2361 (O_2361,N_26577,N_28192);
or UO_2362 (O_2362,N_28901,N_26928);
nor UO_2363 (O_2363,N_27444,N_26375);
nor UO_2364 (O_2364,N_26361,N_25973);
xnor UO_2365 (O_2365,N_27526,N_29508);
nor UO_2366 (O_2366,N_26693,N_28449);
xor UO_2367 (O_2367,N_28303,N_28938);
and UO_2368 (O_2368,N_26663,N_29458);
and UO_2369 (O_2369,N_27844,N_26838);
nand UO_2370 (O_2370,N_28403,N_27771);
nor UO_2371 (O_2371,N_26275,N_27429);
nor UO_2372 (O_2372,N_28039,N_29376);
xnor UO_2373 (O_2373,N_28122,N_27177);
nand UO_2374 (O_2374,N_29695,N_26959);
and UO_2375 (O_2375,N_26916,N_27879);
and UO_2376 (O_2376,N_28679,N_25288);
nor UO_2377 (O_2377,N_25627,N_25620);
nor UO_2378 (O_2378,N_25735,N_25165);
or UO_2379 (O_2379,N_29270,N_27792);
or UO_2380 (O_2380,N_27479,N_29339);
or UO_2381 (O_2381,N_27104,N_28813);
and UO_2382 (O_2382,N_26189,N_29915);
nor UO_2383 (O_2383,N_25509,N_28406);
and UO_2384 (O_2384,N_25815,N_26942);
xnor UO_2385 (O_2385,N_25015,N_26420);
or UO_2386 (O_2386,N_26010,N_27118);
xnor UO_2387 (O_2387,N_29204,N_25762);
or UO_2388 (O_2388,N_27053,N_26294);
or UO_2389 (O_2389,N_29585,N_28394);
or UO_2390 (O_2390,N_26695,N_28163);
and UO_2391 (O_2391,N_25134,N_27811);
or UO_2392 (O_2392,N_26750,N_28550);
or UO_2393 (O_2393,N_29952,N_26338);
nand UO_2394 (O_2394,N_25616,N_28023);
and UO_2395 (O_2395,N_27633,N_25468);
nand UO_2396 (O_2396,N_28923,N_29162);
nand UO_2397 (O_2397,N_28593,N_27818);
nand UO_2398 (O_2398,N_26417,N_25419);
or UO_2399 (O_2399,N_26299,N_28127);
nor UO_2400 (O_2400,N_25269,N_26487);
or UO_2401 (O_2401,N_25505,N_29256);
nor UO_2402 (O_2402,N_26193,N_27265);
and UO_2403 (O_2403,N_27741,N_26786);
nor UO_2404 (O_2404,N_29363,N_28442);
nand UO_2405 (O_2405,N_28481,N_28761);
and UO_2406 (O_2406,N_29820,N_26801);
nand UO_2407 (O_2407,N_27737,N_29659);
nand UO_2408 (O_2408,N_26893,N_26191);
or UO_2409 (O_2409,N_25443,N_26857);
nand UO_2410 (O_2410,N_27146,N_28525);
nand UO_2411 (O_2411,N_27773,N_28971);
nor UO_2412 (O_2412,N_27963,N_28994);
nand UO_2413 (O_2413,N_25621,N_29697);
xnor UO_2414 (O_2414,N_27402,N_27433);
or UO_2415 (O_2415,N_26725,N_26039);
and UO_2416 (O_2416,N_27087,N_29476);
xnor UO_2417 (O_2417,N_27884,N_25787);
nor UO_2418 (O_2418,N_28145,N_28222);
nand UO_2419 (O_2419,N_29639,N_28111);
and UO_2420 (O_2420,N_29377,N_25988);
or UO_2421 (O_2421,N_28378,N_27044);
xnor UO_2422 (O_2422,N_25893,N_28472);
nor UO_2423 (O_2423,N_25125,N_27705);
nor UO_2424 (O_2424,N_25897,N_25830);
or UO_2425 (O_2425,N_25999,N_26945);
and UO_2426 (O_2426,N_25386,N_25206);
nand UO_2427 (O_2427,N_27340,N_28314);
and UO_2428 (O_2428,N_28625,N_29446);
or UO_2429 (O_2429,N_27517,N_28724);
nor UO_2430 (O_2430,N_27262,N_28638);
nor UO_2431 (O_2431,N_25656,N_27246);
nand UO_2432 (O_2432,N_28501,N_29289);
and UO_2433 (O_2433,N_27326,N_27898);
xor UO_2434 (O_2434,N_28228,N_28566);
nor UO_2435 (O_2435,N_28572,N_27059);
or UO_2436 (O_2436,N_26185,N_29844);
and UO_2437 (O_2437,N_27912,N_28484);
or UO_2438 (O_2438,N_27533,N_25322);
nor UO_2439 (O_2439,N_27673,N_26113);
nand UO_2440 (O_2440,N_26205,N_25520);
and UO_2441 (O_2441,N_27285,N_27986);
and UO_2442 (O_2442,N_25032,N_27333);
or UO_2443 (O_2443,N_25850,N_26329);
or UO_2444 (O_2444,N_26455,N_27211);
and UO_2445 (O_2445,N_29398,N_26167);
or UO_2446 (O_2446,N_26267,N_28810);
or UO_2447 (O_2447,N_29616,N_27396);
nand UO_2448 (O_2448,N_25748,N_27016);
xnor UO_2449 (O_2449,N_29238,N_29111);
or UO_2450 (O_2450,N_27315,N_27681);
and UO_2451 (O_2451,N_28548,N_27430);
or UO_2452 (O_2452,N_28464,N_28745);
and UO_2453 (O_2453,N_29834,N_27938);
or UO_2454 (O_2454,N_25984,N_27406);
nand UO_2455 (O_2455,N_25252,N_28204);
nor UO_2456 (O_2456,N_26843,N_26204);
or UO_2457 (O_2457,N_27341,N_25795);
and UO_2458 (O_2458,N_25805,N_29789);
and UO_2459 (O_2459,N_26151,N_25701);
or UO_2460 (O_2460,N_29392,N_25585);
or UO_2461 (O_2461,N_29427,N_26115);
and UO_2462 (O_2462,N_25183,N_27977);
nand UO_2463 (O_2463,N_25734,N_28987);
or UO_2464 (O_2464,N_25099,N_27290);
or UO_2465 (O_2465,N_25464,N_26355);
or UO_2466 (O_2466,N_29676,N_25314);
nor UO_2467 (O_2467,N_26140,N_26782);
nor UO_2468 (O_2468,N_26000,N_29199);
nor UO_2469 (O_2469,N_26419,N_29020);
xor UO_2470 (O_2470,N_26062,N_27477);
and UO_2471 (O_2471,N_26106,N_27467);
nor UO_2472 (O_2472,N_28483,N_27103);
xor UO_2473 (O_2473,N_27414,N_28290);
and UO_2474 (O_2474,N_27356,N_28541);
and UO_2475 (O_2475,N_28132,N_26091);
nand UO_2476 (O_2476,N_29863,N_28751);
or UO_2477 (O_2477,N_27890,N_29750);
nand UO_2478 (O_2478,N_25600,N_28779);
or UO_2479 (O_2479,N_29275,N_27217);
xnor UO_2480 (O_2480,N_28458,N_26145);
nand UO_2481 (O_2481,N_26330,N_27125);
or UO_2482 (O_2482,N_27462,N_27410);
nor UO_2483 (O_2483,N_29178,N_25693);
and UO_2484 (O_2484,N_27353,N_29681);
nand UO_2485 (O_2485,N_25615,N_27274);
xnor UO_2486 (O_2486,N_27511,N_29718);
nor UO_2487 (O_2487,N_27000,N_29205);
nor UO_2488 (O_2488,N_29360,N_27272);
nand UO_2489 (O_2489,N_29411,N_28337);
nor UO_2490 (O_2490,N_28218,N_27187);
and UO_2491 (O_2491,N_25366,N_27645);
or UO_2492 (O_2492,N_27398,N_27536);
or UO_2493 (O_2493,N_27147,N_28993);
nand UO_2494 (O_2494,N_26143,N_26169);
and UO_2495 (O_2495,N_26041,N_26565);
and UO_2496 (O_2496,N_28178,N_26699);
xor UO_2497 (O_2497,N_28117,N_28381);
nor UO_2498 (O_2498,N_25063,N_26781);
xnor UO_2499 (O_2499,N_25472,N_26070);
xor UO_2500 (O_2500,N_25005,N_29312);
xnor UO_2501 (O_2501,N_25928,N_28535);
or UO_2502 (O_2502,N_25251,N_26188);
or UO_2503 (O_2503,N_29509,N_28485);
or UO_2504 (O_2504,N_27955,N_27159);
nor UO_2505 (O_2505,N_26118,N_25927);
or UO_2506 (O_2506,N_27005,N_25360);
and UO_2507 (O_2507,N_28282,N_27002);
nand UO_2508 (O_2508,N_27892,N_28335);
and UO_2509 (O_2509,N_28526,N_26925);
nand UO_2510 (O_2510,N_28345,N_29418);
nand UO_2511 (O_2511,N_28888,N_29072);
and UO_2512 (O_2512,N_26402,N_25973);
nor UO_2513 (O_2513,N_26342,N_29511);
nand UO_2514 (O_2514,N_25348,N_25095);
and UO_2515 (O_2515,N_25881,N_25580);
xor UO_2516 (O_2516,N_28199,N_27173);
nand UO_2517 (O_2517,N_27016,N_25548);
nor UO_2518 (O_2518,N_25318,N_26684);
and UO_2519 (O_2519,N_27791,N_26754);
nand UO_2520 (O_2520,N_29718,N_27946);
and UO_2521 (O_2521,N_29798,N_27864);
nor UO_2522 (O_2522,N_28218,N_25625);
nand UO_2523 (O_2523,N_29805,N_26738);
or UO_2524 (O_2524,N_25387,N_26541);
nor UO_2525 (O_2525,N_27163,N_28514);
xor UO_2526 (O_2526,N_29348,N_25756);
or UO_2527 (O_2527,N_25919,N_28334);
nand UO_2528 (O_2528,N_28069,N_29398);
nor UO_2529 (O_2529,N_27754,N_27253);
nand UO_2530 (O_2530,N_29888,N_28524);
and UO_2531 (O_2531,N_25346,N_27261);
xor UO_2532 (O_2532,N_28165,N_26918);
and UO_2533 (O_2533,N_27851,N_28324);
or UO_2534 (O_2534,N_28402,N_29267);
xnor UO_2535 (O_2535,N_28377,N_28140);
and UO_2536 (O_2536,N_25918,N_28922);
or UO_2537 (O_2537,N_25266,N_28313);
and UO_2538 (O_2538,N_26951,N_28472);
or UO_2539 (O_2539,N_27066,N_27610);
nand UO_2540 (O_2540,N_27019,N_26437);
nor UO_2541 (O_2541,N_28688,N_26801);
nand UO_2542 (O_2542,N_29001,N_29880);
or UO_2543 (O_2543,N_29159,N_27840);
nor UO_2544 (O_2544,N_29902,N_26086);
nor UO_2545 (O_2545,N_29343,N_25384);
and UO_2546 (O_2546,N_29249,N_29294);
or UO_2547 (O_2547,N_26878,N_25716);
and UO_2548 (O_2548,N_27046,N_27346);
nand UO_2549 (O_2549,N_26481,N_26690);
and UO_2550 (O_2550,N_29332,N_26671);
nand UO_2551 (O_2551,N_25338,N_29746);
xnor UO_2552 (O_2552,N_25303,N_28593);
nor UO_2553 (O_2553,N_25377,N_26167);
xnor UO_2554 (O_2554,N_29793,N_25039);
or UO_2555 (O_2555,N_28523,N_28854);
or UO_2556 (O_2556,N_27673,N_27012);
and UO_2557 (O_2557,N_29708,N_26495);
xor UO_2558 (O_2558,N_26554,N_27931);
nand UO_2559 (O_2559,N_25285,N_29794);
or UO_2560 (O_2560,N_26893,N_29895);
nand UO_2561 (O_2561,N_29857,N_27626);
or UO_2562 (O_2562,N_25984,N_26921);
or UO_2563 (O_2563,N_28592,N_28605);
or UO_2564 (O_2564,N_29341,N_28827);
or UO_2565 (O_2565,N_25203,N_28055);
or UO_2566 (O_2566,N_29578,N_27876);
or UO_2567 (O_2567,N_27047,N_27584);
and UO_2568 (O_2568,N_25004,N_29806);
nand UO_2569 (O_2569,N_26234,N_29220);
nor UO_2570 (O_2570,N_28207,N_25910);
and UO_2571 (O_2571,N_29471,N_26273);
xor UO_2572 (O_2572,N_27395,N_28881);
nand UO_2573 (O_2573,N_25511,N_25463);
nor UO_2574 (O_2574,N_27369,N_28678);
xor UO_2575 (O_2575,N_27263,N_29068);
nand UO_2576 (O_2576,N_27322,N_26240);
and UO_2577 (O_2577,N_25924,N_27637);
and UO_2578 (O_2578,N_28016,N_27956);
nand UO_2579 (O_2579,N_27695,N_27157);
nor UO_2580 (O_2580,N_26782,N_25956);
and UO_2581 (O_2581,N_26290,N_25273);
xor UO_2582 (O_2582,N_26973,N_25638);
and UO_2583 (O_2583,N_27831,N_26810);
and UO_2584 (O_2584,N_29947,N_29762);
xnor UO_2585 (O_2585,N_28434,N_26923);
and UO_2586 (O_2586,N_26906,N_27042);
nor UO_2587 (O_2587,N_26147,N_28672);
or UO_2588 (O_2588,N_26878,N_25509);
and UO_2589 (O_2589,N_27593,N_29464);
nor UO_2590 (O_2590,N_25538,N_26046);
nor UO_2591 (O_2591,N_28972,N_28958);
and UO_2592 (O_2592,N_28797,N_28308);
nor UO_2593 (O_2593,N_29828,N_25399);
nor UO_2594 (O_2594,N_29584,N_26853);
nand UO_2595 (O_2595,N_29174,N_25874);
nor UO_2596 (O_2596,N_25381,N_29855);
and UO_2597 (O_2597,N_28861,N_29617);
nand UO_2598 (O_2598,N_28568,N_28953);
nor UO_2599 (O_2599,N_27202,N_26279);
or UO_2600 (O_2600,N_29462,N_26591);
or UO_2601 (O_2601,N_28627,N_27294);
or UO_2602 (O_2602,N_28466,N_27880);
and UO_2603 (O_2603,N_27995,N_28026);
nor UO_2604 (O_2604,N_28272,N_28431);
nand UO_2605 (O_2605,N_29740,N_27782);
and UO_2606 (O_2606,N_27351,N_25795);
nand UO_2607 (O_2607,N_28458,N_25503);
or UO_2608 (O_2608,N_27911,N_26243);
or UO_2609 (O_2609,N_28950,N_29046);
nand UO_2610 (O_2610,N_26424,N_29545);
or UO_2611 (O_2611,N_28278,N_27815);
or UO_2612 (O_2612,N_27469,N_29637);
or UO_2613 (O_2613,N_27811,N_27426);
nor UO_2614 (O_2614,N_28757,N_29159);
or UO_2615 (O_2615,N_28283,N_27881);
and UO_2616 (O_2616,N_29986,N_25448);
nor UO_2617 (O_2617,N_29411,N_26254);
nor UO_2618 (O_2618,N_25039,N_25778);
nor UO_2619 (O_2619,N_26760,N_26565);
or UO_2620 (O_2620,N_27727,N_27163);
nor UO_2621 (O_2621,N_29404,N_29856);
or UO_2622 (O_2622,N_25922,N_27303);
and UO_2623 (O_2623,N_29141,N_29035);
nor UO_2624 (O_2624,N_25861,N_29761);
or UO_2625 (O_2625,N_25088,N_27649);
nand UO_2626 (O_2626,N_29339,N_26270);
nor UO_2627 (O_2627,N_29885,N_29662);
nor UO_2628 (O_2628,N_27529,N_27073);
xnor UO_2629 (O_2629,N_27734,N_29105);
nand UO_2630 (O_2630,N_27342,N_28676);
and UO_2631 (O_2631,N_27184,N_29771);
and UO_2632 (O_2632,N_26188,N_29946);
nand UO_2633 (O_2633,N_26633,N_27722);
or UO_2634 (O_2634,N_28067,N_25621);
nor UO_2635 (O_2635,N_28063,N_25675);
nand UO_2636 (O_2636,N_25618,N_25105);
xnor UO_2637 (O_2637,N_25383,N_28677);
and UO_2638 (O_2638,N_28218,N_27132);
nor UO_2639 (O_2639,N_27383,N_29546);
and UO_2640 (O_2640,N_28557,N_26427);
and UO_2641 (O_2641,N_29813,N_28506);
nand UO_2642 (O_2642,N_28363,N_29968);
nand UO_2643 (O_2643,N_26739,N_29144);
nor UO_2644 (O_2644,N_29689,N_29504);
and UO_2645 (O_2645,N_28144,N_27209);
nor UO_2646 (O_2646,N_29323,N_26419);
and UO_2647 (O_2647,N_25422,N_25354);
nand UO_2648 (O_2648,N_29266,N_27030);
or UO_2649 (O_2649,N_26987,N_29745);
and UO_2650 (O_2650,N_25405,N_28192);
or UO_2651 (O_2651,N_29259,N_28823);
nor UO_2652 (O_2652,N_27006,N_29701);
and UO_2653 (O_2653,N_26834,N_26516);
or UO_2654 (O_2654,N_26361,N_29980);
or UO_2655 (O_2655,N_26572,N_27306);
or UO_2656 (O_2656,N_29975,N_28219);
and UO_2657 (O_2657,N_29004,N_26493);
or UO_2658 (O_2658,N_25688,N_28698);
nor UO_2659 (O_2659,N_25929,N_28268);
and UO_2660 (O_2660,N_28163,N_26119);
nand UO_2661 (O_2661,N_26425,N_25168);
nand UO_2662 (O_2662,N_27437,N_25045);
or UO_2663 (O_2663,N_25719,N_26277);
xnor UO_2664 (O_2664,N_28535,N_26141);
xor UO_2665 (O_2665,N_26395,N_27673);
nand UO_2666 (O_2666,N_25660,N_29629);
and UO_2667 (O_2667,N_29152,N_25075);
nand UO_2668 (O_2668,N_28932,N_27760);
nor UO_2669 (O_2669,N_25046,N_27774);
and UO_2670 (O_2670,N_26688,N_26307);
nand UO_2671 (O_2671,N_26802,N_26268);
xor UO_2672 (O_2672,N_28451,N_26644);
nor UO_2673 (O_2673,N_28503,N_29170);
nand UO_2674 (O_2674,N_28686,N_28224);
nand UO_2675 (O_2675,N_25177,N_25969);
xnor UO_2676 (O_2676,N_29703,N_27819);
nor UO_2677 (O_2677,N_26292,N_25350);
nand UO_2678 (O_2678,N_26744,N_26367);
nor UO_2679 (O_2679,N_29702,N_27179);
nor UO_2680 (O_2680,N_28179,N_29142);
nand UO_2681 (O_2681,N_25442,N_25884);
and UO_2682 (O_2682,N_29352,N_28652);
or UO_2683 (O_2683,N_27472,N_27760);
nor UO_2684 (O_2684,N_28000,N_29305);
nand UO_2685 (O_2685,N_26198,N_29512);
nand UO_2686 (O_2686,N_29331,N_25918);
nor UO_2687 (O_2687,N_27167,N_29890);
and UO_2688 (O_2688,N_28397,N_27838);
and UO_2689 (O_2689,N_26321,N_26348);
or UO_2690 (O_2690,N_29432,N_29722);
nand UO_2691 (O_2691,N_29560,N_27487);
nor UO_2692 (O_2692,N_27254,N_28500);
and UO_2693 (O_2693,N_29918,N_28168);
and UO_2694 (O_2694,N_26404,N_27115);
nor UO_2695 (O_2695,N_29506,N_28311);
and UO_2696 (O_2696,N_27654,N_26072);
nor UO_2697 (O_2697,N_28318,N_27110);
nor UO_2698 (O_2698,N_27175,N_25823);
nor UO_2699 (O_2699,N_26840,N_29852);
or UO_2700 (O_2700,N_25588,N_26784);
and UO_2701 (O_2701,N_25011,N_26439);
nand UO_2702 (O_2702,N_27866,N_29294);
nor UO_2703 (O_2703,N_28889,N_29953);
or UO_2704 (O_2704,N_29093,N_28386);
or UO_2705 (O_2705,N_29532,N_26789);
nand UO_2706 (O_2706,N_29670,N_29868);
xnor UO_2707 (O_2707,N_28564,N_25254);
nor UO_2708 (O_2708,N_26166,N_28073);
or UO_2709 (O_2709,N_26591,N_26361);
and UO_2710 (O_2710,N_27340,N_28251);
or UO_2711 (O_2711,N_26944,N_25519);
xnor UO_2712 (O_2712,N_28357,N_28668);
xnor UO_2713 (O_2713,N_26928,N_28170);
nor UO_2714 (O_2714,N_27435,N_29215);
or UO_2715 (O_2715,N_27869,N_28389);
nor UO_2716 (O_2716,N_25888,N_26156);
or UO_2717 (O_2717,N_28026,N_26053);
nand UO_2718 (O_2718,N_26611,N_25507);
nor UO_2719 (O_2719,N_29196,N_28638);
nor UO_2720 (O_2720,N_25718,N_26710);
and UO_2721 (O_2721,N_25764,N_29678);
nor UO_2722 (O_2722,N_26407,N_26056);
or UO_2723 (O_2723,N_27082,N_25780);
nor UO_2724 (O_2724,N_27873,N_25646);
or UO_2725 (O_2725,N_25763,N_28657);
or UO_2726 (O_2726,N_25075,N_27103);
and UO_2727 (O_2727,N_26186,N_29548);
or UO_2728 (O_2728,N_26894,N_25578);
or UO_2729 (O_2729,N_25979,N_28709);
or UO_2730 (O_2730,N_26794,N_29203);
or UO_2731 (O_2731,N_26013,N_29169);
nand UO_2732 (O_2732,N_25753,N_25817);
nor UO_2733 (O_2733,N_29822,N_29659);
and UO_2734 (O_2734,N_28768,N_27357);
nor UO_2735 (O_2735,N_28303,N_26198);
or UO_2736 (O_2736,N_28867,N_27642);
or UO_2737 (O_2737,N_25565,N_28676);
and UO_2738 (O_2738,N_27479,N_26764);
nor UO_2739 (O_2739,N_26637,N_29748);
nor UO_2740 (O_2740,N_25401,N_27324);
nand UO_2741 (O_2741,N_28237,N_26720);
nand UO_2742 (O_2742,N_29188,N_28415);
and UO_2743 (O_2743,N_28974,N_28704);
xnor UO_2744 (O_2744,N_26290,N_25794);
or UO_2745 (O_2745,N_25803,N_25015);
or UO_2746 (O_2746,N_25606,N_28754);
nor UO_2747 (O_2747,N_27784,N_25392);
or UO_2748 (O_2748,N_27186,N_26807);
nor UO_2749 (O_2749,N_25960,N_26532);
nand UO_2750 (O_2750,N_25748,N_27356);
xnor UO_2751 (O_2751,N_25278,N_25846);
and UO_2752 (O_2752,N_28098,N_29516);
nor UO_2753 (O_2753,N_27439,N_27014);
and UO_2754 (O_2754,N_26463,N_26756);
nor UO_2755 (O_2755,N_28708,N_27969);
nand UO_2756 (O_2756,N_27603,N_29972);
or UO_2757 (O_2757,N_28619,N_25072);
nor UO_2758 (O_2758,N_26114,N_26699);
or UO_2759 (O_2759,N_25243,N_26403);
and UO_2760 (O_2760,N_29095,N_29475);
nor UO_2761 (O_2761,N_28649,N_29228);
and UO_2762 (O_2762,N_26511,N_28740);
or UO_2763 (O_2763,N_25111,N_25799);
nand UO_2764 (O_2764,N_26162,N_25537);
nand UO_2765 (O_2765,N_27824,N_25794);
or UO_2766 (O_2766,N_26733,N_28660);
xor UO_2767 (O_2767,N_27794,N_28200);
or UO_2768 (O_2768,N_28808,N_28559);
and UO_2769 (O_2769,N_26472,N_26020);
or UO_2770 (O_2770,N_28227,N_28284);
or UO_2771 (O_2771,N_26126,N_25211);
or UO_2772 (O_2772,N_27677,N_26227);
or UO_2773 (O_2773,N_25125,N_28936);
or UO_2774 (O_2774,N_26679,N_28571);
and UO_2775 (O_2775,N_28634,N_28648);
and UO_2776 (O_2776,N_29956,N_29744);
nand UO_2777 (O_2777,N_28073,N_26592);
nand UO_2778 (O_2778,N_26329,N_26912);
nand UO_2779 (O_2779,N_26243,N_26033);
nand UO_2780 (O_2780,N_28687,N_26119);
nor UO_2781 (O_2781,N_26760,N_26075);
nand UO_2782 (O_2782,N_26776,N_27832);
or UO_2783 (O_2783,N_29491,N_27940);
and UO_2784 (O_2784,N_26922,N_26937);
or UO_2785 (O_2785,N_27040,N_28750);
nor UO_2786 (O_2786,N_25341,N_28509);
or UO_2787 (O_2787,N_25324,N_25686);
nand UO_2788 (O_2788,N_27317,N_29380);
or UO_2789 (O_2789,N_29353,N_27526);
or UO_2790 (O_2790,N_25822,N_26069);
nor UO_2791 (O_2791,N_29003,N_26220);
nor UO_2792 (O_2792,N_29092,N_25317);
or UO_2793 (O_2793,N_29862,N_25392);
and UO_2794 (O_2794,N_25157,N_25498);
xnor UO_2795 (O_2795,N_29674,N_29624);
nand UO_2796 (O_2796,N_25936,N_27249);
xnor UO_2797 (O_2797,N_29674,N_29052);
nand UO_2798 (O_2798,N_28521,N_28384);
xnor UO_2799 (O_2799,N_29651,N_26919);
nand UO_2800 (O_2800,N_27916,N_26481);
and UO_2801 (O_2801,N_25138,N_28854);
nor UO_2802 (O_2802,N_29406,N_29117);
or UO_2803 (O_2803,N_25680,N_26134);
nand UO_2804 (O_2804,N_28441,N_29936);
and UO_2805 (O_2805,N_27409,N_26808);
nand UO_2806 (O_2806,N_29537,N_26909);
xor UO_2807 (O_2807,N_25121,N_25213);
nand UO_2808 (O_2808,N_27953,N_25645);
or UO_2809 (O_2809,N_26313,N_28514);
or UO_2810 (O_2810,N_29009,N_29029);
nand UO_2811 (O_2811,N_27314,N_28288);
or UO_2812 (O_2812,N_29568,N_26073);
nand UO_2813 (O_2813,N_26511,N_25123);
and UO_2814 (O_2814,N_26281,N_28872);
or UO_2815 (O_2815,N_26895,N_25667);
nand UO_2816 (O_2816,N_27215,N_27646);
nor UO_2817 (O_2817,N_25896,N_25368);
xor UO_2818 (O_2818,N_28231,N_27793);
nor UO_2819 (O_2819,N_25615,N_29752);
nand UO_2820 (O_2820,N_28692,N_26218);
nor UO_2821 (O_2821,N_29684,N_25101);
or UO_2822 (O_2822,N_29246,N_25725);
nor UO_2823 (O_2823,N_25888,N_25421);
nand UO_2824 (O_2824,N_27188,N_26672);
or UO_2825 (O_2825,N_26057,N_26657);
nor UO_2826 (O_2826,N_25489,N_27384);
nand UO_2827 (O_2827,N_28038,N_25202);
and UO_2828 (O_2828,N_26694,N_26029);
nor UO_2829 (O_2829,N_27192,N_26077);
nor UO_2830 (O_2830,N_28880,N_27283);
xor UO_2831 (O_2831,N_25722,N_25020);
nor UO_2832 (O_2832,N_26597,N_29047);
nor UO_2833 (O_2833,N_26363,N_27502);
and UO_2834 (O_2834,N_25677,N_28475);
or UO_2835 (O_2835,N_28342,N_27467);
and UO_2836 (O_2836,N_29993,N_29920);
nand UO_2837 (O_2837,N_25078,N_26370);
nand UO_2838 (O_2838,N_26798,N_26105);
or UO_2839 (O_2839,N_28536,N_26933);
and UO_2840 (O_2840,N_27801,N_27890);
or UO_2841 (O_2841,N_29170,N_27928);
xor UO_2842 (O_2842,N_29459,N_27251);
xnor UO_2843 (O_2843,N_29444,N_29189);
nand UO_2844 (O_2844,N_26544,N_28080);
nand UO_2845 (O_2845,N_28940,N_29007);
or UO_2846 (O_2846,N_28819,N_25188);
or UO_2847 (O_2847,N_29061,N_26704);
xnor UO_2848 (O_2848,N_26146,N_25895);
nor UO_2849 (O_2849,N_26792,N_29828);
and UO_2850 (O_2850,N_25036,N_25090);
or UO_2851 (O_2851,N_25292,N_27308);
and UO_2852 (O_2852,N_25849,N_26899);
and UO_2853 (O_2853,N_26155,N_27308);
nand UO_2854 (O_2854,N_27911,N_28482);
and UO_2855 (O_2855,N_26696,N_28569);
or UO_2856 (O_2856,N_25542,N_25142);
and UO_2857 (O_2857,N_27073,N_29641);
or UO_2858 (O_2858,N_27860,N_25213);
xnor UO_2859 (O_2859,N_28320,N_29979);
and UO_2860 (O_2860,N_25642,N_27542);
nand UO_2861 (O_2861,N_25208,N_27397);
nand UO_2862 (O_2862,N_27678,N_25807);
or UO_2863 (O_2863,N_28300,N_29323);
nor UO_2864 (O_2864,N_26609,N_29811);
or UO_2865 (O_2865,N_28308,N_25234);
and UO_2866 (O_2866,N_26924,N_28809);
nand UO_2867 (O_2867,N_26987,N_27084);
xnor UO_2868 (O_2868,N_28634,N_26287);
and UO_2869 (O_2869,N_25164,N_29604);
nand UO_2870 (O_2870,N_27177,N_26092);
nand UO_2871 (O_2871,N_26554,N_29683);
and UO_2872 (O_2872,N_27255,N_27907);
nor UO_2873 (O_2873,N_27998,N_25385);
nand UO_2874 (O_2874,N_27302,N_29161);
or UO_2875 (O_2875,N_27322,N_28626);
or UO_2876 (O_2876,N_26008,N_25026);
nand UO_2877 (O_2877,N_26301,N_28236);
nor UO_2878 (O_2878,N_28547,N_27228);
xnor UO_2879 (O_2879,N_29505,N_29313);
and UO_2880 (O_2880,N_25470,N_28704);
or UO_2881 (O_2881,N_29195,N_28875);
nor UO_2882 (O_2882,N_25257,N_29658);
xnor UO_2883 (O_2883,N_26687,N_28482);
nand UO_2884 (O_2884,N_28691,N_25382);
nor UO_2885 (O_2885,N_29017,N_28742);
nand UO_2886 (O_2886,N_28803,N_28369);
xor UO_2887 (O_2887,N_25031,N_27982);
and UO_2888 (O_2888,N_28216,N_29789);
and UO_2889 (O_2889,N_25922,N_28298);
nor UO_2890 (O_2890,N_26781,N_27372);
nor UO_2891 (O_2891,N_26666,N_27723);
nor UO_2892 (O_2892,N_28097,N_26189);
and UO_2893 (O_2893,N_26190,N_27918);
and UO_2894 (O_2894,N_27986,N_25019);
or UO_2895 (O_2895,N_27984,N_29240);
and UO_2896 (O_2896,N_26979,N_25681);
and UO_2897 (O_2897,N_26775,N_29087);
nand UO_2898 (O_2898,N_27868,N_29841);
nand UO_2899 (O_2899,N_25421,N_25059);
xnor UO_2900 (O_2900,N_25015,N_27830);
or UO_2901 (O_2901,N_25305,N_25873);
nor UO_2902 (O_2902,N_28985,N_28444);
or UO_2903 (O_2903,N_29733,N_26038);
nor UO_2904 (O_2904,N_25663,N_29565);
nand UO_2905 (O_2905,N_26418,N_26088);
or UO_2906 (O_2906,N_29416,N_25408);
and UO_2907 (O_2907,N_25999,N_25408);
nand UO_2908 (O_2908,N_27886,N_27358);
or UO_2909 (O_2909,N_25715,N_28099);
nand UO_2910 (O_2910,N_25799,N_26263);
xnor UO_2911 (O_2911,N_25417,N_26947);
nand UO_2912 (O_2912,N_26444,N_29510);
or UO_2913 (O_2913,N_27005,N_25814);
nand UO_2914 (O_2914,N_25866,N_29067);
nor UO_2915 (O_2915,N_28189,N_29599);
nor UO_2916 (O_2916,N_26533,N_28661);
nor UO_2917 (O_2917,N_29366,N_29809);
or UO_2918 (O_2918,N_25792,N_25129);
nand UO_2919 (O_2919,N_25418,N_26671);
and UO_2920 (O_2920,N_28532,N_29229);
nor UO_2921 (O_2921,N_29233,N_25084);
nand UO_2922 (O_2922,N_29616,N_28050);
nor UO_2923 (O_2923,N_28280,N_28865);
or UO_2924 (O_2924,N_29533,N_29219);
nor UO_2925 (O_2925,N_27269,N_29184);
and UO_2926 (O_2926,N_26591,N_25521);
nand UO_2927 (O_2927,N_29157,N_25164);
or UO_2928 (O_2928,N_27275,N_28105);
nor UO_2929 (O_2929,N_27210,N_28501);
nor UO_2930 (O_2930,N_25092,N_25082);
nand UO_2931 (O_2931,N_26789,N_27151);
or UO_2932 (O_2932,N_25673,N_25273);
and UO_2933 (O_2933,N_25081,N_25076);
nor UO_2934 (O_2934,N_28825,N_27583);
or UO_2935 (O_2935,N_27250,N_27397);
nor UO_2936 (O_2936,N_26056,N_26718);
and UO_2937 (O_2937,N_25081,N_29859);
nand UO_2938 (O_2938,N_27319,N_27261);
nor UO_2939 (O_2939,N_25008,N_26542);
nor UO_2940 (O_2940,N_28919,N_27398);
nand UO_2941 (O_2941,N_25754,N_27292);
and UO_2942 (O_2942,N_28455,N_28635);
or UO_2943 (O_2943,N_28663,N_28879);
nand UO_2944 (O_2944,N_28763,N_25532);
xor UO_2945 (O_2945,N_25525,N_29720);
nor UO_2946 (O_2946,N_28846,N_29536);
or UO_2947 (O_2947,N_29739,N_27195);
or UO_2948 (O_2948,N_29358,N_26324);
and UO_2949 (O_2949,N_25903,N_26467);
nand UO_2950 (O_2950,N_26222,N_27893);
and UO_2951 (O_2951,N_25280,N_25453);
and UO_2952 (O_2952,N_27072,N_26346);
xor UO_2953 (O_2953,N_26382,N_25005);
nand UO_2954 (O_2954,N_29771,N_28929);
nand UO_2955 (O_2955,N_28288,N_25170);
nand UO_2956 (O_2956,N_29427,N_29614);
or UO_2957 (O_2957,N_28340,N_27915);
or UO_2958 (O_2958,N_27566,N_28990);
or UO_2959 (O_2959,N_27837,N_25832);
nor UO_2960 (O_2960,N_28737,N_26482);
or UO_2961 (O_2961,N_27889,N_25867);
or UO_2962 (O_2962,N_26994,N_29123);
nor UO_2963 (O_2963,N_29907,N_27807);
or UO_2964 (O_2964,N_28040,N_25917);
and UO_2965 (O_2965,N_27791,N_29419);
and UO_2966 (O_2966,N_28487,N_28163);
or UO_2967 (O_2967,N_27073,N_29873);
or UO_2968 (O_2968,N_26683,N_29739);
nand UO_2969 (O_2969,N_29377,N_25128);
nor UO_2970 (O_2970,N_29537,N_29359);
nand UO_2971 (O_2971,N_28220,N_28744);
xnor UO_2972 (O_2972,N_27364,N_28861);
nand UO_2973 (O_2973,N_25787,N_29358);
nand UO_2974 (O_2974,N_29199,N_25118);
xnor UO_2975 (O_2975,N_26862,N_25371);
or UO_2976 (O_2976,N_25089,N_28848);
nor UO_2977 (O_2977,N_28969,N_29503);
xor UO_2978 (O_2978,N_27675,N_28979);
nand UO_2979 (O_2979,N_27327,N_26124);
and UO_2980 (O_2980,N_27610,N_25614);
or UO_2981 (O_2981,N_25492,N_27542);
or UO_2982 (O_2982,N_26294,N_26801);
and UO_2983 (O_2983,N_27809,N_28684);
and UO_2984 (O_2984,N_29013,N_25434);
and UO_2985 (O_2985,N_27328,N_25817);
nor UO_2986 (O_2986,N_25480,N_25012);
nor UO_2987 (O_2987,N_26113,N_27458);
or UO_2988 (O_2988,N_28042,N_28370);
and UO_2989 (O_2989,N_27157,N_26185);
and UO_2990 (O_2990,N_25871,N_29170);
nor UO_2991 (O_2991,N_27620,N_25569);
nor UO_2992 (O_2992,N_26652,N_29321);
and UO_2993 (O_2993,N_28677,N_27844);
nand UO_2994 (O_2994,N_29372,N_27959);
xor UO_2995 (O_2995,N_27823,N_29077);
and UO_2996 (O_2996,N_25344,N_28996);
or UO_2997 (O_2997,N_25747,N_27110);
nor UO_2998 (O_2998,N_29908,N_29821);
and UO_2999 (O_2999,N_28084,N_29606);
nor UO_3000 (O_3000,N_27702,N_28939);
or UO_3001 (O_3001,N_27859,N_26170);
and UO_3002 (O_3002,N_29630,N_25292);
nand UO_3003 (O_3003,N_29173,N_26405);
nor UO_3004 (O_3004,N_27415,N_29407);
nor UO_3005 (O_3005,N_25496,N_28807);
xnor UO_3006 (O_3006,N_27775,N_25264);
and UO_3007 (O_3007,N_25123,N_28553);
or UO_3008 (O_3008,N_25032,N_27845);
nand UO_3009 (O_3009,N_26704,N_28302);
or UO_3010 (O_3010,N_28216,N_25682);
and UO_3011 (O_3011,N_26908,N_29116);
or UO_3012 (O_3012,N_27206,N_27309);
nor UO_3013 (O_3013,N_29333,N_28211);
or UO_3014 (O_3014,N_25781,N_28136);
nor UO_3015 (O_3015,N_29762,N_26480);
or UO_3016 (O_3016,N_28133,N_29763);
nor UO_3017 (O_3017,N_27024,N_29545);
or UO_3018 (O_3018,N_29155,N_29464);
and UO_3019 (O_3019,N_29433,N_25137);
and UO_3020 (O_3020,N_26646,N_25657);
or UO_3021 (O_3021,N_25059,N_28797);
nand UO_3022 (O_3022,N_28090,N_25016);
nor UO_3023 (O_3023,N_27046,N_25121);
xnor UO_3024 (O_3024,N_28717,N_28627);
nand UO_3025 (O_3025,N_28705,N_29756);
or UO_3026 (O_3026,N_25012,N_26654);
nand UO_3027 (O_3027,N_26323,N_27415);
nand UO_3028 (O_3028,N_26120,N_27640);
nand UO_3029 (O_3029,N_26647,N_28168);
nor UO_3030 (O_3030,N_26641,N_26296);
nand UO_3031 (O_3031,N_29347,N_29860);
nor UO_3032 (O_3032,N_25152,N_27369);
nor UO_3033 (O_3033,N_27450,N_29966);
or UO_3034 (O_3034,N_28688,N_25175);
or UO_3035 (O_3035,N_27350,N_28727);
or UO_3036 (O_3036,N_28693,N_28412);
nand UO_3037 (O_3037,N_29159,N_26808);
nor UO_3038 (O_3038,N_28484,N_26392);
and UO_3039 (O_3039,N_29812,N_27123);
nor UO_3040 (O_3040,N_26966,N_28240);
nor UO_3041 (O_3041,N_26838,N_28571);
or UO_3042 (O_3042,N_29056,N_25234);
and UO_3043 (O_3043,N_26778,N_29252);
and UO_3044 (O_3044,N_25432,N_26865);
and UO_3045 (O_3045,N_26006,N_29647);
or UO_3046 (O_3046,N_25310,N_28204);
or UO_3047 (O_3047,N_28431,N_27478);
nor UO_3048 (O_3048,N_26473,N_28726);
or UO_3049 (O_3049,N_27574,N_26417);
nor UO_3050 (O_3050,N_25593,N_29333);
or UO_3051 (O_3051,N_28716,N_27455);
nor UO_3052 (O_3052,N_25164,N_26108);
or UO_3053 (O_3053,N_29257,N_29128);
nor UO_3054 (O_3054,N_27588,N_26190);
and UO_3055 (O_3055,N_28577,N_27368);
or UO_3056 (O_3056,N_26919,N_26176);
or UO_3057 (O_3057,N_27279,N_25617);
nor UO_3058 (O_3058,N_26988,N_29297);
nand UO_3059 (O_3059,N_28712,N_28670);
and UO_3060 (O_3060,N_27185,N_26233);
or UO_3061 (O_3061,N_27898,N_29020);
or UO_3062 (O_3062,N_27126,N_28193);
xor UO_3063 (O_3063,N_25995,N_28530);
or UO_3064 (O_3064,N_25297,N_27046);
or UO_3065 (O_3065,N_29015,N_26522);
nor UO_3066 (O_3066,N_29473,N_26860);
and UO_3067 (O_3067,N_25132,N_28632);
nor UO_3068 (O_3068,N_29038,N_25415);
and UO_3069 (O_3069,N_25137,N_26445);
or UO_3070 (O_3070,N_28906,N_27858);
nand UO_3071 (O_3071,N_28334,N_28214);
or UO_3072 (O_3072,N_28660,N_26455);
xnor UO_3073 (O_3073,N_25693,N_28102);
or UO_3074 (O_3074,N_27989,N_26828);
or UO_3075 (O_3075,N_26488,N_28855);
nand UO_3076 (O_3076,N_27589,N_29096);
and UO_3077 (O_3077,N_29895,N_26522);
nor UO_3078 (O_3078,N_28570,N_27875);
nand UO_3079 (O_3079,N_25009,N_25529);
nor UO_3080 (O_3080,N_29795,N_25460);
and UO_3081 (O_3081,N_29855,N_28724);
xnor UO_3082 (O_3082,N_29653,N_27712);
nand UO_3083 (O_3083,N_27450,N_28805);
or UO_3084 (O_3084,N_27656,N_29311);
nor UO_3085 (O_3085,N_28170,N_26768);
and UO_3086 (O_3086,N_25568,N_28060);
xor UO_3087 (O_3087,N_26968,N_29806);
xnor UO_3088 (O_3088,N_29816,N_27553);
nor UO_3089 (O_3089,N_26641,N_27810);
nor UO_3090 (O_3090,N_26141,N_28478);
nand UO_3091 (O_3091,N_29075,N_28181);
or UO_3092 (O_3092,N_28600,N_25074);
nor UO_3093 (O_3093,N_25751,N_27629);
nand UO_3094 (O_3094,N_28407,N_26187);
xnor UO_3095 (O_3095,N_29950,N_28403);
or UO_3096 (O_3096,N_28000,N_25135);
nor UO_3097 (O_3097,N_28234,N_29155);
nor UO_3098 (O_3098,N_25610,N_29371);
nor UO_3099 (O_3099,N_25579,N_26652);
nand UO_3100 (O_3100,N_28365,N_29297);
nand UO_3101 (O_3101,N_29469,N_27188);
nand UO_3102 (O_3102,N_26014,N_27889);
and UO_3103 (O_3103,N_26006,N_27584);
nand UO_3104 (O_3104,N_28602,N_28379);
nand UO_3105 (O_3105,N_25975,N_26305);
and UO_3106 (O_3106,N_27189,N_26532);
nand UO_3107 (O_3107,N_28689,N_29447);
and UO_3108 (O_3108,N_25134,N_27324);
nor UO_3109 (O_3109,N_26747,N_28151);
nor UO_3110 (O_3110,N_28923,N_26945);
nand UO_3111 (O_3111,N_29151,N_26002);
and UO_3112 (O_3112,N_28338,N_25187);
or UO_3113 (O_3113,N_27064,N_29601);
or UO_3114 (O_3114,N_27211,N_26407);
xor UO_3115 (O_3115,N_27614,N_29536);
or UO_3116 (O_3116,N_27242,N_25118);
and UO_3117 (O_3117,N_25429,N_26601);
nand UO_3118 (O_3118,N_26659,N_25246);
nor UO_3119 (O_3119,N_27856,N_29382);
or UO_3120 (O_3120,N_29062,N_28298);
or UO_3121 (O_3121,N_25738,N_27510);
and UO_3122 (O_3122,N_26643,N_29483);
nand UO_3123 (O_3123,N_25599,N_28662);
xor UO_3124 (O_3124,N_27667,N_29413);
nand UO_3125 (O_3125,N_25309,N_27979);
nor UO_3126 (O_3126,N_28273,N_27521);
nor UO_3127 (O_3127,N_26121,N_29412);
nor UO_3128 (O_3128,N_29675,N_25876);
nor UO_3129 (O_3129,N_25186,N_27528);
and UO_3130 (O_3130,N_28431,N_27979);
and UO_3131 (O_3131,N_25185,N_29866);
nand UO_3132 (O_3132,N_27811,N_26368);
nor UO_3133 (O_3133,N_26496,N_27165);
nor UO_3134 (O_3134,N_25930,N_29939);
nand UO_3135 (O_3135,N_27892,N_27093);
and UO_3136 (O_3136,N_25116,N_28983);
or UO_3137 (O_3137,N_27502,N_29350);
and UO_3138 (O_3138,N_26587,N_27237);
or UO_3139 (O_3139,N_29304,N_26932);
nand UO_3140 (O_3140,N_27935,N_27205);
nor UO_3141 (O_3141,N_26590,N_27583);
or UO_3142 (O_3142,N_29529,N_27777);
nand UO_3143 (O_3143,N_25141,N_28427);
xor UO_3144 (O_3144,N_25001,N_29175);
nand UO_3145 (O_3145,N_28877,N_26453);
nand UO_3146 (O_3146,N_28240,N_25557);
nor UO_3147 (O_3147,N_27949,N_25702);
and UO_3148 (O_3148,N_28459,N_29424);
nand UO_3149 (O_3149,N_25319,N_25214);
nand UO_3150 (O_3150,N_29573,N_26062);
and UO_3151 (O_3151,N_26870,N_28442);
nor UO_3152 (O_3152,N_28538,N_27641);
nor UO_3153 (O_3153,N_27345,N_29125);
nor UO_3154 (O_3154,N_25266,N_27964);
nand UO_3155 (O_3155,N_26490,N_29387);
nand UO_3156 (O_3156,N_26995,N_25130);
and UO_3157 (O_3157,N_26047,N_28426);
nand UO_3158 (O_3158,N_28645,N_28687);
or UO_3159 (O_3159,N_28015,N_27888);
nand UO_3160 (O_3160,N_26747,N_26256);
or UO_3161 (O_3161,N_25359,N_29845);
xnor UO_3162 (O_3162,N_27321,N_29294);
nand UO_3163 (O_3163,N_26120,N_29145);
nor UO_3164 (O_3164,N_25408,N_29383);
or UO_3165 (O_3165,N_25431,N_26383);
or UO_3166 (O_3166,N_26545,N_26651);
or UO_3167 (O_3167,N_29869,N_29530);
nand UO_3168 (O_3168,N_27248,N_25661);
or UO_3169 (O_3169,N_27690,N_26149);
nor UO_3170 (O_3170,N_27147,N_25093);
nand UO_3171 (O_3171,N_28119,N_26636);
and UO_3172 (O_3172,N_28064,N_28586);
and UO_3173 (O_3173,N_29623,N_29878);
nand UO_3174 (O_3174,N_28242,N_25741);
and UO_3175 (O_3175,N_25772,N_26673);
nor UO_3176 (O_3176,N_29163,N_26437);
nand UO_3177 (O_3177,N_29429,N_28456);
nor UO_3178 (O_3178,N_26541,N_25362);
nand UO_3179 (O_3179,N_29176,N_29323);
and UO_3180 (O_3180,N_26564,N_27854);
and UO_3181 (O_3181,N_25960,N_27692);
or UO_3182 (O_3182,N_26264,N_29247);
xor UO_3183 (O_3183,N_27252,N_27649);
or UO_3184 (O_3184,N_26179,N_26076);
or UO_3185 (O_3185,N_29010,N_28125);
nor UO_3186 (O_3186,N_28136,N_29951);
nand UO_3187 (O_3187,N_26687,N_29311);
and UO_3188 (O_3188,N_25359,N_29335);
xnor UO_3189 (O_3189,N_29292,N_27987);
xor UO_3190 (O_3190,N_28307,N_29928);
and UO_3191 (O_3191,N_27165,N_29503);
or UO_3192 (O_3192,N_28193,N_25786);
nand UO_3193 (O_3193,N_26026,N_26314);
nor UO_3194 (O_3194,N_27292,N_29350);
nand UO_3195 (O_3195,N_28391,N_27886);
and UO_3196 (O_3196,N_28214,N_25100);
nand UO_3197 (O_3197,N_28993,N_27180);
nor UO_3198 (O_3198,N_29838,N_29630);
nor UO_3199 (O_3199,N_27941,N_29064);
and UO_3200 (O_3200,N_29955,N_25886);
nand UO_3201 (O_3201,N_27542,N_25886);
nor UO_3202 (O_3202,N_27344,N_27573);
nand UO_3203 (O_3203,N_27582,N_25253);
and UO_3204 (O_3204,N_28577,N_25283);
xnor UO_3205 (O_3205,N_26728,N_29858);
and UO_3206 (O_3206,N_25511,N_29231);
nand UO_3207 (O_3207,N_27426,N_27943);
and UO_3208 (O_3208,N_29054,N_25309);
nand UO_3209 (O_3209,N_28521,N_28632);
nor UO_3210 (O_3210,N_27497,N_28340);
nand UO_3211 (O_3211,N_29918,N_26508);
or UO_3212 (O_3212,N_27555,N_29108);
and UO_3213 (O_3213,N_25305,N_25945);
nor UO_3214 (O_3214,N_29608,N_29100);
xnor UO_3215 (O_3215,N_26656,N_27251);
nor UO_3216 (O_3216,N_28982,N_25151);
or UO_3217 (O_3217,N_26235,N_25077);
nor UO_3218 (O_3218,N_28625,N_25511);
nand UO_3219 (O_3219,N_27464,N_29885);
or UO_3220 (O_3220,N_27668,N_27625);
xor UO_3221 (O_3221,N_25933,N_26156);
xor UO_3222 (O_3222,N_28403,N_26163);
nand UO_3223 (O_3223,N_26700,N_27290);
and UO_3224 (O_3224,N_28190,N_28076);
nand UO_3225 (O_3225,N_28131,N_25224);
or UO_3226 (O_3226,N_26174,N_29496);
nor UO_3227 (O_3227,N_27941,N_27744);
or UO_3228 (O_3228,N_29530,N_25327);
and UO_3229 (O_3229,N_28043,N_28181);
nor UO_3230 (O_3230,N_27080,N_27025);
xor UO_3231 (O_3231,N_25378,N_27857);
nand UO_3232 (O_3232,N_27616,N_25837);
and UO_3233 (O_3233,N_25664,N_25971);
nor UO_3234 (O_3234,N_26013,N_27611);
xor UO_3235 (O_3235,N_29200,N_28649);
nor UO_3236 (O_3236,N_26739,N_29999);
nand UO_3237 (O_3237,N_26265,N_26618);
and UO_3238 (O_3238,N_26877,N_26750);
nor UO_3239 (O_3239,N_26447,N_28417);
nand UO_3240 (O_3240,N_26743,N_29146);
nor UO_3241 (O_3241,N_27431,N_28704);
nand UO_3242 (O_3242,N_27248,N_26344);
nand UO_3243 (O_3243,N_26253,N_25973);
nor UO_3244 (O_3244,N_25825,N_25892);
nor UO_3245 (O_3245,N_26529,N_28255);
nor UO_3246 (O_3246,N_26706,N_29262);
nand UO_3247 (O_3247,N_29278,N_27339);
xor UO_3248 (O_3248,N_29752,N_28885);
and UO_3249 (O_3249,N_26268,N_27629);
nand UO_3250 (O_3250,N_27380,N_29017);
nand UO_3251 (O_3251,N_29059,N_28755);
and UO_3252 (O_3252,N_28542,N_29966);
xor UO_3253 (O_3253,N_29118,N_25549);
xor UO_3254 (O_3254,N_26049,N_25163);
and UO_3255 (O_3255,N_27856,N_28828);
or UO_3256 (O_3256,N_28450,N_26770);
or UO_3257 (O_3257,N_26202,N_28968);
xor UO_3258 (O_3258,N_26108,N_26291);
nor UO_3259 (O_3259,N_29552,N_25277);
nand UO_3260 (O_3260,N_28636,N_25025);
or UO_3261 (O_3261,N_27853,N_25480);
and UO_3262 (O_3262,N_29931,N_28333);
and UO_3263 (O_3263,N_29690,N_28727);
nor UO_3264 (O_3264,N_26955,N_29447);
and UO_3265 (O_3265,N_29817,N_27958);
nor UO_3266 (O_3266,N_27103,N_28345);
and UO_3267 (O_3267,N_29803,N_26232);
nand UO_3268 (O_3268,N_25222,N_25414);
nand UO_3269 (O_3269,N_29284,N_28937);
nor UO_3270 (O_3270,N_29443,N_28028);
nor UO_3271 (O_3271,N_29016,N_28067);
nand UO_3272 (O_3272,N_27849,N_25393);
nand UO_3273 (O_3273,N_29969,N_25011);
and UO_3274 (O_3274,N_25528,N_25091);
nand UO_3275 (O_3275,N_26894,N_29828);
or UO_3276 (O_3276,N_25632,N_26905);
nor UO_3277 (O_3277,N_28931,N_28733);
nor UO_3278 (O_3278,N_27601,N_26474);
nand UO_3279 (O_3279,N_26303,N_25553);
nand UO_3280 (O_3280,N_26930,N_29284);
nor UO_3281 (O_3281,N_25752,N_28340);
nand UO_3282 (O_3282,N_26710,N_27377);
or UO_3283 (O_3283,N_27393,N_29226);
nor UO_3284 (O_3284,N_27176,N_27194);
nor UO_3285 (O_3285,N_25427,N_26750);
and UO_3286 (O_3286,N_25565,N_28927);
nor UO_3287 (O_3287,N_28746,N_25920);
nor UO_3288 (O_3288,N_29673,N_25187);
nor UO_3289 (O_3289,N_29081,N_28089);
nor UO_3290 (O_3290,N_25593,N_29101);
nor UO_3291 (O_3291,N_26023,N_26799);
and UO_3292 (O_3292,N_27534,N_25944);
and UO_3293 (O_3293,N_29635,N_29371);
nor UO_3294 (O_3294,N_29374,N_29627);
nand UO_3295 (O_3295,N_27216,N_26710);
nor UO_3296 (O_3296,N_27978,N_26916);
and UO_3297 (O_3297,N_27688,N_29703);
nand UO_3298 (O_3298,N_25860,N_26535);
and UO_3299 (O_3299,N_26438,N_26967);
and UO_3300 (O_3300,N_29690,N_25054);
and UO_3301 (O_3301,N_26097,N_29518);
and UO_3302 (O_3302,N_26308,N_29363);
or UO_3303 (O_3303,N_25305,N_25263);
and UO_3304 (O_3304,N_27527,N_28867);
nor UO_3305 (O_3305,N_28303,N_27115);
and UO_3306 (O_3306,N_26116,N_26109);
nand UO_3307 (O_3307,N_28627,N_28547);
nand UO_3308 (O_3308,N_28099,N_26829);
and UO_3309 (O_3309,N_26753,N_26682);
nor UO_3310 (O_3310,N_28723,N_28445);
or UO_3311 (O_3311,N_28346,N_26381);
or UO_3312 (O_3312,N_29271,N_28515);
and UO_3313 (O_3313,N_29057,N_25571);
nor UO_3314 (O_3314,N_25009,N_26769);
nand UO_3315 (O_3315,N_29263,N_28688);
and UO_3316 (O_3316,N_27314,N_28935);
nand UO_3317 (O_3317,N_25563,N_29564);
and UO_3318 (O_3318,N_25738,N_28554);
nand UO_3319 (O_3319,N_26229,N_27259);
or UO_3320 (O_3320,N_27407,N_29741);
nand UO_3321 (O_3321,N_25982,N_28810);
or UO_3322 (O_3322,N_29051,N_27143);
nor UO_3323 (O_3323,N_27329,N_26777);
nor UO_3324 (O_3324,N_26102,N_28930);
nor UO_3325 (O_3325,N_26078,N_28271);
or UO_3326 (O_3326,N_25095,N_28958);
and UO_3327 (O_3327,N_27841,N_26201);
or UO_3328 (O_3328,N_27757,N_27634);
nand UO_3329 (O_3329,N_26473,N_25738);
nor UO_3330 (O_3330,N_29229,N_27228);
nor UO_3331 (O_3331,N_28035,N_28283);
nand UO_3332 (O_3332,N_28928,N_27619);
nor UO_3333 (O_3333,N_26930,N_26935);
nor UO_3334 (O_3334,N_29286,N_25905);
nor UO_3335 (O_3335,N_29559,N_26144);
nor UO_3336 (O_3336,N_26650,N_29060);
nor UO_3337 (O_3337,N_28129,N_26628);
xnor UO_3338 (O_3338,N_28983,N_29733);
nand UO_3339 (O_3339,N_28276,N_28849);
and UO_3340 (O_3340,N_28657,N_28807);
or UO_3341 (O_3341,N_29950,N_29335);
nand UO_3342 (O_3342,N_28279,N_26308);
nand UO_3343 (O_3343,N_28846,N_27880);
or UO_3344 (O_3344,N_26714,N_28747);
and UO_3345 (O_3345,N_28992,N_29092);
nor UO_3346 (O_3346,N_29770,N_29978);
nand UO_3347 (O_3347,N_29124,N_28525);
nor UO_3348 (O_3348,N_28836,N_29419);
nor UO_3349 (O_3349,N_28280,N_25088);
or UO_3350 (O_3350,N_27881,N_25026);
nor UO_3351 (O_3351,N_29847,N_29260);
nand UO_3352 (O_3352,N_27321,N_25791);
or UO_3353 (O_3353,N_26051,N_25760);
and UO_3354 (O_3354,N_25439,N_25810);
nand UO_3355 (O_3355,N_28288,N_27883);
and UO_3356 (O_3356,N_29355,N_28015);
nor UO_3357 (O_3357,N_29575,N_25945);
nor UO_3358 (O_3358,N_29153,N_25170);
nand UO_3359 (O_3359,N_26618,N_25752);
nand UO_3360 (O_3360,N_29960,N_29671);
and UO_3361 (O_3361,N_29463,N_28730);
or UO_3362 (O_3362,N_28773,N_27573);
or UO_3363 (O_3363,N_26898,N_27338);
nand UO_3364 (O_3364,N_26302,N_25772);
nand UO_3365 (O_3365,N_29882,N_25200);
nor UO_3366 (O_3366,N_29763,N_26462);
nand UO_3367 (O_3367,N_28442,N_28631);
or UO_3368 (O_3368,N_29746,N_29111);
or UO_3369 (O_3369,N_25492,N_25232);
or UO_3370 (O_3370,N_26799,N_26854);
and UO_3371 (O_3371,N_26884,N_27130);
and UO_3372 (O_3372,N_28285,N_29065);
and UO_3373 (O_3373,N_25294,N_27188);
xnor UO_3374 (O_3374,N_28679,N_26871);
nand UO_3375 (O_3375,N_26564,N_28964);
nand UO_3376 (O_3376,N_28136,N_28333);
and UO_3377 (O_3377,N_29475,N_28585);
nand UO_3378 (O_3378,N_29844,N_28072);
or UO_3379 (O_3379,N_29493,N_27312);
or UO_3380 (O_3380,N_29401,N_29314);
and UO_3381 (O_3381,N_25912,N_25390);
or UO_3382 (O_3382,N_27260,N_25104);
nand UO_3383 (O_3383,N_27755,N_28406);
and UO_3384 (O_3384,N_25580,N_29596);
or UO_3385 (O_3385,N_29429,N_27574);
nor UO_3386 (O_3386,N_26200,N_26717);
or UO_3387 (O_3387,N_27412,N_25210);
nand UO_3388 (O_3388,N_25734,N_27368);
or UO_3389 (O_3389,N_25185,N_28839);
nand UO_3390 (O_3390,N_25801,N_26594);
or UO_3391 (O_3391,N_28900,N_27128);
or UO_3392 (O_3392,N_29188,N_29339);
and UO_3393 (O_3393,N_29351,N_27029);
nand UO_3394 (O_3394,N_26589,N_25104);
or UO_3395 (O_3395,N_27945,N_29809);
or UO_3396 (O_3396,N_28297,N_26016);
nor UO_3397 (O_3397,N_28428,N_29875);
nor UO_3398 (O_3398,N_29450,N_29723);
and UO_3399 (O_3399,N_25022,N_26380);
and UO_3400 (O_3400,N_29192,N_28153);
and UO_3401 (O_3401,N_26612,N_28986);
and UO_3402 (O_3402,N_28098,N_26502);
xor UO_3403 (O_3403,N_29576,N_26657);
nor UO_3404 (O_3404,N_27553,N_25775);
and UO_3405 (O_3405,N_29133,N_25745);
xor UO_3406 (O_3406,N_25056,N_29159);
nand UO_3407 (O_3407,N_25625,N_25504);
nor UO_3408 (O_3408,N_28593,N_28048);
nand UO_3409 (O_3409,N_25314,N_28073);
nor UO_3410 (O_3410,N_29868,N_26308);
nor UO_3411 (O_3411,N_28197,N_28052);
and UO_3412 (O_3412,N_28898,N_28841);
nand UO_3413 (O_3413,N_28664,N_25738);
or UO_3414 (O_3414,N_25194,N_28593);
and UO_3415 (O_3415,N_29665,N_28761);
xor UO_3416 (O_3416,N_26732,N_27558);
or UO_3417 (O_3417,N_26336,N_25503);
nor UO_3418 (O_3418,N_28960,N_29926);
or UO_3419 (O_3419,N_26916,N_26876);
and UO_3420 (O_3420,N_28363,N_26544);
or UO_3421 (O_3421,N_26853,N_28065);
and UO_3422 (O_3422,N_27727,N_27986);
nand UO_3423 (O_3423,N_25915,N_28731);
or UO_3424 (O_3424,N_26342,N_28834);
nand UO_3425 (O_3425,N_25478,N_25745);
nor UO_3426 (O_3426,N_25608,N_27576);
and UO_3427 (O_3427,N_28092,N_27302);
nor UO_3428 (O_3428,N_26648,N_28503);
and UO_3429 (O_3429,N_28315,N_29539);
xor UO_3430 (O_3430,N_26765,N_28678);
or UO_3431 (O_3431,N_28379,N_25261);
nor UO_3432 (O_3432,N_26395,N_26202);
nor UO_3433 (O_3433,N_27615,N_26552);
nand UO_3434 (O_3434,N_29675,N_27239);
and UO_3435 (O_3435,N_27761,N_25623);
and UO_3436 (O_3436,N_28738,N_29663);
nand UO_3437 (O_3437,N_27803,N_25394);
nand UO_3438 (O_3438,N_29930,N_27144);
nor UO_3439 (O_3439,N_28776,N_27639);
xnor UO_3440 (O_3440,N_26742,N_26554);
nor UO_3441 (O_3441,N_29139,N_27215);
xor UO_3442 (O_3442,N_29165,N_28631);
nand UO_3443 (O_3443,N_25443,N_27676);
or UO_3444 (O_3444,N_26332,N_26398);
nor UO_3445 (O_3445,N_27403,N_25505);
and UO_3446 (O_3446,N_28050,N_26126);
or UO_3447 (O_3447,N_25553,N_25507);
nor UO_3448 (O_3448,N_25970,N_28969);
or UO_3449 (O_3449,N_29722,N_29932);
and UO_3450 (O_3450,N_26323,N_26469);
nor UO_3451 (O_3451,N_25187,N_27493);
nand UO_3452 (O_3452,N_29124,N_29031);
and UO_3453 (O_3453,N_25026,N_26889);
or UO_3454 (O_3454,N_27696,N_28043);
and UO_3455 (O_3455,N_29130,N_29831);
and UO_3456 (O_3456,N_29880,N_27291);
or UO_3457 (O_3457,N_29019,N_29007);
nor UO_3458 (O_3458,N_28568,N_29299);
nor UO_3459 (O_3459,N_28391,N_26891);
xnor UO_3460 (O_3460,N_26503,N_26147);
nor UO_3461 (O_3461,N_29468,N_29995);
and UO_3462 (O_3462,N_29026,N_25928);
nand UO_3463 (O_3463,N_27602,N_26051);
and UO_3464 (O_3464,N_26814,N_29290);
and UO_3465 (O_3465,N_26761,N_28060);
and UO_3466 (O_3466,N_26671,N_27267);
nor UO_3467 (O_3467,N_28333,N_28669);
nand UO_3468 (O_3468,N_29905,N_28132);
or UO_3469 (O_3469,N_26154,N_26611);
nor UO_3470 (O_3470,N_29131,N_25605);
and UO_3471 (O_3471,N_27537,N_25062);
or UO_3472 (O_3472,N_28164,N_26155);
and UO_3473 (O_3473,N_25067,N_28195);
or UO_3474 (O_3474,N_29848,N_26039);
nor UO_3475 (O_3475,N_25372,N_26737);
nand UO_3476 (O_3476,N_28323,N_27028);
nor UO_3477 (O_3477,N_27296,N_26124);
and UO_3478 (O_3478,N_27372,N_25770);
nor UO_3479 (O_3479,N_26767,N_25882);
xnor UO_3480 (O_3480,N_27473,N_28267);
nand UO_3481 (O_3481,N_27808,N_27058);
and UO_3482 (O_3482,N_27909,N_27581);
nor UO_3483 (O_3483,N_26974,N_25463);
or UO_3484 (O_3484,N_28364,N_29456);
nor UO_3485 (O_3485,N_28699,N_26814);
nand UO_3486 (O_3486,N_29820,N_29079);
nand UO_3487 (O_3487,N_26253,N_29379);
nand UO_3488 (O_3488,N_29562,N_28564);
nand UO_3489 (O_3489,N_29820,N_27117);
or UO_3490 (O_3490,N_25930,N_25485);
nor UO_3491 (O_3491,N_25610,N_27811);
or UO_3492 (O_3492,N_29842,N_29122);
and UO_3493 (O_3493,N_27529,N_28974);
or UO_3494 (O_3494,N_29275,N_25884);
or UO_3495 (O_3495,N_26085,N_26840);
nand UO_3496 (O_3496,N_27800,N_27112);
or UO_3497 (O_3497,N_28718,N_28202);
and UO_3498 (O_3498,N_26269,N_27790);
and UO_3499 (O_3499,N_25637,N_25337);
endmodule