module basic_2500_25000_3000_8_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_1530,In_719);
nor U1 (N_1,In_952,In_349);
xor U2 (N_2,In_432,In_1600);
and U3 (N_3,In_1969,In_2304);
nand U4 (N_4,In_1382,In_350);
or U5 (N_5,In_1380,In_1781);
nand U6 (N_6,In_390,In_553);
nor U7 (N_7,In_448,In_478);
nor U8 (N_8,In_578,In_1129);
nor U9 (N_9,In_1044,In_1877);
xnor U10 (N_10,In_768,In_209);
nand U11 (N_11,In_2376,In_424);
or U12 (N_12,In_2494,In_2085);
or U13 (N_13,In_772,In_1880);
xnor U14 (N_14,In_391,In_1852);
and U15 (N_15,In_1424,In_375);
xnor U16 (N_16,In_2390,In_2311);
xor U17 (N_17,In_1422,In_155);
or U18 (N_18,In_866,In_2440);
xnor U19 (N_19,In_2087,In_2415);
nor U20 (N_20,In_2281,In_2312);
xnor U21 (N_21,In_1690,In_175);
or U22 (N_22,In_1923,In_1723);
nor U23 (N_23,In_118,In_454);
xnor U24 (N_24,In_214,In_2242);
xor U25 (N_25,In_912,In_1376);
xor U26 (N_26,In_184,In_1570);
nand U27 (N_27,In_1778,In_1579);
xnor U28 (N_28,In_557,In_867);
xnor U29 (N_29,In_1192,In_346);
nor U30 (N_30,In_584,In_527);
or U31 (N_31,In_1055,In_192);
nor U32 (N_32,In_825,In_2245);
or U33 (N_33,In_67,In_105);
nor U34 (N_34,In_2407,In_1047);
and U35 (N_35,In_2172,In_1910);
nand U36 (N_36,In_1872,In_1130);
nor U37 (N_37,In_2075,In_909);
or U38 (N_38,In_2306,In_1624);
or U39 (N_39,In_2350,In_2069);
or U40 (N_40,In_1306,In_571);
nand U41 (N_41,In_1832,In_2026);
xnor U42 (N_42,In_1788,In_61);
xnor U43 (N_43,In_1598,In_2447);
nor U44 (N_44,In_2394,In_2092);
xnor U45 (N_45,In_1360,In_2122);
nor U46 (N_46,In_750,In_1618);
nor U47 (N_47,In_1451,In_1891);
xor U48 (N_48,In_1709,In_1042);
nor U49 (N_49,In_1198,In_1409);
nor U50 (N_50,In_332,In_1372);
and U51 (N_51,In_1580,In_30);
nor U52 (N_52,In_2015,In_1289);
and U53 (N_53,In_1492,In_296);
xor U54 (N_54,In_1842,In_2315);
xor U55 (N_55,In_2317,In_309);
nand U56 (N_56,In_2046,In_1317);
nand U57 (N_57,In_2247,In_1020);
or U58 (N_58,In_1605,In_551);
and U59 (N_59,In_926,In_1185);
nand U60 (N_60,In_1241,In_872);
nand U61 (N_61,In_1377,In_306);
or U62 (N_62,In_953,In_2479);
nand U63 (N_63,In_1194,In_2208);
xnor U64 (N_64,In_762,In_2114);
or U65 (N_65,In_1909,In_335);
nor U66 (N_66,In_860,In_2078);
and U67 (N_67,In_530,In_876);
nor U68 (N_68,In_776,In_746);
nor U69 (N_69,In_1193,In_751);
nor U70 (N_70,In_1966,In_1133);
xor U71 (N_71,In_2464,In_2442);
xor U72 (N_72,In_1448,In_660);
nand U73 (N_73,In_2370,In_1225);
and U74 (N_74,In_2364,In_15);
xnor U75 (N_75,In_1186,In_2039);
nand U76 (N_76,In_841,In_1721);
nand U77 (N_77,In_2262,In_646);
and U78 (N_78,In_2051,In_1964);
xnor U79 (N_79,In_745,In_2427);
xnor U80 (N_80,In_112,In_1074);
xnor U81 (N_81,In_502,In_904);
xnor U82 (N_82,In_1714,In_2420);
and U83 (N_83,In_778,In_368);
xnor U84 (N_84,In_1655,In_504);
and U85 (N_85,In_986,In_2455);
xor U86 (N_86,In_1716,In_2024);
and U87 (N_87,In_1199,In_2068);
or U88 (N_88,In_738,In_987);
or U89 (N_89,In_942,In_2027);
nand U90 (N_90,In_1879,In_1371);
and U91 (N_91,In_1255,In_2182);
xnor U92 (N_92,In_483,In_2056);
nand U93 (N_93,In_948,In_1223);
nor U94 (N_94,In_1974,In_1062);
nor U95 (N_95,In_1623,In_1314);
nor U96 (N_96,In_1989,In_2426);
or U97 (N_97,In_2117,In_321);
and U98 (N_98,In_205,In_2058);
or U99 (N_99,In_1531,In_1678);
nor U100 (N_100,In_2012,In_2296);
or U101 (N_101,In_2169,In_617);
or U102 (N_102,In_2480,In_635);
nand U103 (N_103,In_2324,In_190);
and U104 (N_104,In_1119,In_605);
nand U105 (N_105,In_2082,In_1075);
and U106 (N_106,In_1845,In_556);
and U107 (N_107,In_2072,In_2166);
or U108 (N_108,In_2441,In_2177);
and U109 (N_109,In_903,In_1218);
nor U110 (N_110,In_651,In_1246);
nor U111 (N_111,In_1337,In_1549);
nor U112 (N_112,In_2237,In_918);
nor U113 (N_113,In_1578,In_1860);
xnor U114 (N_114,In_131,In_954);
or U115 (N_115,In_2196,In_1008);
or U116 (N_116,In_677,In_1819);
xor U117 (N_117,In_1743,In_1853);
and U118 (N_118,In_2385,In_207);
xnor U119 (N_119,In_717,In_995);
nand U120 (N_120,In_2071,In_2103);
or U121 (N_121,In_577,In_1379);
nand U122 (N_122,In_2498,In_1768);
nor U123 (N_123,In_927,In_1428);
or U124 (N_124,In_2272,In_1071);
or U125 (N_125,In_8,In_1958);
and U126 (N_126,In_307,In_1741);
and U127 (N_127,In_1975,In_1333);
and U128 (N_128,In_638,In_404);
or U129 (N_129,In_117,In_1340);
xnor U130 (N_130,In_1355,In_869);
nor U131 (N_131,In_1828,In_1951);
and U132 (N_132,In_1560,In_1747);
or U133 (N_133,In_1445,In_2485);
xor U134 (N_134,In_1058,In_1405);
and U135 (N_135,In_1722,In_832);
nor U136 (N_136,In_1341,In_1127);
nor U137 (N_137,In_965,In_905);
xor U138 (N_138,In_2421,In_411);
or U139 (N_139,In_264,In_27);
nand U140 (N_140,In_1458,In_2112);
nand U141 (N_141,In_758,In_2193);
nand U142 (N_142,In_2448,In_1940);
and U143 (N_143,In_1354,In_724);
and U144 (N_144,In_1191,In_1864);
xnor U145 (N_145,In_49,In_742);
and U146 (N_146,In_1801,In_1034);
xnor U147 (N_147,In_1095,In_1336);
nor U148 (N_148,In_1991,In_2481);
and U149 (N_149,In_1449,In_2150);
nor U150 (N_150,In_2229,In_539);
and U151 (N_151,In_453,In_100);
or U152 (N_152,In_1608,In_602);
and U153 (N_153,In_1569,In_524);
nor U154 (N_154,In_1988,In_973);
and U155 (N_155,In_450,In_883);
nor U156 (N_156,In_21,In_37);
nand U157 (N_157,In_993,In_2226);
or U158 (N_158,In_1196,In_135);
nand U159 (N_159,In_203,In_749);
and U160 (N_160,In_1719,In_398);
xnor U161 (N_161,In_179,In_1563);
nor U162 (N_162,In_2343,In_1415);
nand U163 (N_163,In_1472,In_354);
or U164 (N_164,In_1046,In_251);
nand U165 (N_165,In_2257,In_2469);
nand U166 (N_166,In_1524,In_1285);
and U167 (N_167,In_229,In_649);
xnor U168 (N_168,In_1259,In_2021);
nor U169 (N_169,In_366,In_1911);
nor U170 (N_170,In_1824,In_937);
nand U171 (N_171,In_809,In_480);
or U172 (N_172,In_1184,In_958);
and U173 (N_173,In_1815,In_753);
nand U174 (N_174,In_1443,In_115);
or U175 (N_175,In_1724,In_2280);
nand U176 (N_176,In_1307,In_1757);
or U177 (N_177,In_598,In_1630);
nand U178 (N_178,In_397,In_360);
and U179 (N_179,In_80,In_1452);
and U180 (N_180,In_122,In_1232);
and U181 (N_181,In_102,In_940);
or U182 (N_182,In_1632,In_1423);
xnor U183 (N_183,In_886,In_508);
and U184 (N_184,In_1677,In_1599);
nand U185 (N_185,In_1012,In_96);
or U186 (N_186,In_1992,In_2111);
nand U187 (N_187,In_689,In_1890);
and U188 (N_188,In_1142,In_1201);
or U189 (N_189,In_31,In_1827);
and U190 (N_190,In_1970,In_1150);
or U191 (N_191,In_2206,In_2236);
and U192 (N_192,In_2335,In_811);
nor U193 (N_193,In_2482,In_1844);
nand U194 (N_194,In_1594,In_380);
or U195 (N_195,In_2299,In_26);
nand U196 (N_196,In_523,In_951);
nand U197 (N_197,In_715,In_345);
nor U198 (N_198,In_600,In_1647);
and U199 (N_199,In_138,In_1750);
nand U200 (N_200,In_1421,In_1997);
or U201 (N_201,In_1636,In_2290);
nor U202 (N_202,In_7,In_648);
nor U203 (N_203,In_739,In_1111);
or U204 (N_204,In_1631,In_505);
nor U205 (N_205,In_407,In_1084);
and U206 (N_206,In_270,In_1851);
or U207 (N_207,In_1748,In_2393);
and U208 (N_208,In_1473,In_1670);
and U209 (N_209,In_1485,In_732);
nand U210 (N_210,In_1859,In_1215);
nand U211 (N_211,In_34,In_1510);
nand U212 (N_212,In_1038,In_1369);
and U213 (N_213,In_124,In_1892);
xor U214 (N_214,In_1526,In_1606);
nor U215 (N_215,In_1830,In_2466);
nor U216 (N_216,In_389,In_978);
or U217 (N_217,In_2002,In_2138);
xor U218 (N_218,In_1590,In_662);
nand U219 (N_219,In_2174,In_1260);
xor U220 (N_220,In_850,In_1782);
xor U221 (N_221,In_456,In_95);
or U222 (N_222,In_606,In_1871);
and U223 (N_223,In_2221,In_1460);
or U224 (N_224,In_1641,In_2282);
and U225 (N_225,In_1078,In_984);
and U226 (N_226,In_298,In_356);
or U227 (N_227,In_2373,In_889);
or U228 (N_228,In_844,In_466);
nor U229 (N_229,In_106,In_1274);
nand U230 (N_230,In_1921,In_1013);
nor U231 (N_231,In_1527,In_2310);
xnor U232 (N_232,In_2325,In_2278);
nand U233 (N_233,In_1658,In_84);
nor U234 (N_234,In_1922,In_2048);
and U235 (N_235,In_1941,In_1420);
or U236 (N_236,In_842,In_775);
or U237 (N_237,In_1917,In_1281);
or U238 (N_238,In_1407,In_2368);
and U239 (N_239,In_1004,In_1916);
xnor U240 (N_240,In_1258,In_1935);
xnor U241 (N_241,In_2366,In_2074);
or U242 (N_242,In_1764,In_1049);
xor U243 (N_243,In_2030,In_394);
or U244 (N_244,In_1731,In_1637);
and U245 (N_245,In_1302,In_202);
and U246 (N_246,In_70,In_812);
xnor U247 (N_247,In_2109,In_913);
nand U248 (N_248,In_656,In_1200);
and U249 (N_249,In_1567,In_2486);
or U250 (N_250,In_1924,In_1454);
nor U251 (N_251,In_1616,In_1108);
and U252 (N_252,In_788,In_562);
and U253 (N_253,In_2330,In_1848);
nor U254 (N_254,In_2007,In_1996);
nand U255 (N_255,In_547,In_2429);
and U256 (N_256,In_741,In_2472);
and U257 (N_257,In_2113,In_2277);
and U258 (N_258,In_1070,In_177);
xor U259 (N_259,In_2380,In_697);
nand U260 (N_260,In_2396,In_792);
xnor U261 (N_261,In_1659,In_898);
and U262 (N_262,In_761,In_1931);
xor U263 (N_263,In_1766,In_2107);
xor U264 (N_264,In_1539,In_414);
nand U265 (N_265,In_2295,In_2476);
and U266 (N_266,In_935,In_1332);
nor U267 (N_267,In_1434,In_125);
and U268 (N_268,In_2191,In_248);
xor U269 (N_269,In_2345,In_1168);
and U270 (N_270,In_558,In_782);
or U271 (N_271,In_2301,In_1520);
xnor U272 (N_272,In_862,In_1474);
and U273 (N_273,In_759,In_977);
nand U274 (N_274,In_1090,In_1684);
and U275 (N_275,In_1479,In_716);
or U276 (N_276,In_252,In_2126);
and U277 (N_277,In_2096,In_1106);
nand U278 (N_278,In_960,In_1865);
nor U279 (N_279,In_2367,In_111);
nand U280 (N_280,In_1235,In_2130);
xnor U281 (N_281,In_897,In_971);
nor U282 (N_282,In_259,In_733);
nand U283 (N_283,In_290,In_2129);
xnor U284 (N_284,In_2383,In_1236);
or U285 (N_285,In_1017,In_1884);
and U286 (N_286,In_2100,In_1553);
and U287 (N_287,In_386,In_1282);
and U288 (N_288,In_899,In_644);
or U289 (N_289,In_1505,In_1284);
xor U290 (N_290,In_2134,In_400);
xnor U291 (N_291,In_694,In_2384);
nor U292 (N_292,In_1596,In_2149);
xnor U293 (N_293,In_1547,In_2187);
and U294 (N_294,In_939,In_2408);
xnor U295 (N_295,In_710,In_2400);
and U296 (N_296,In_181,In_514);
nand U297 (N_297,In_1098,In_1103);
and U298 (N_298,In_1813,In_87);
and U299 (N_299,In_1759,In_443);
xor U300 (N_300,In_1809,In_2016);
nor U301 (N_301,In_462,In_1016);
nand U302 (N_302,In_591,In_2120);
nor U303 (N_303,In_126,In_534);
or U304 (N_304,In_678,In_76);
and U305 (N_305,In_342,In_1169);
nand U306 (N_306,In_1981,In_283);
xnor U307 (N_307,In_784,In_150);
and U308 (N_308,In_799,In_133);
xnor U309 (N_309,In_2035,In_1650);
and U310 (N_310,In_29,In_374);
xnor U311 (N_311,In_1643,In_2409);
and U312 (N_312,In_2207,In_1418);
nor U313 (N_313,In_1740,In_1475);
nor U314 (N_314,In_2478,In_1182);
nand U315 (N_315,In_2332,In_1595);
xnor U316 (N_316,In_1404,In_1378);
nand U317 (N_317,In_2417,In_982);
and U318 (N_318,In_1694,In_979);
and U319 (N_319,In_2352,In_1021);
and U320 (N_320,In_1551,In_1088);
and U321 (N_321,In_1022,In_2080);
and U322 (N_322,In_1311,In_1811);
nand U323 (N_323,In_281,In_774);
nand U324 (N_324,In_1575,In_1107);
nand U325 (N_325,In_323,In_121);
nand U326 (N_326,In_1870,In_2294);
and U327 (N_327,In_243,In_1277);
xor U328 (N_328,In_2451,In_1490);
xnor U329 (N_329,In_654,In_616);
or U330 (N_330,In_471,In_1908);
nand U331 (N_331,In_1459,In_1649);
xor U332 (N_332,In_408,In_172);
xnor U333 (N_333,In_526,In_1050);
and U334 (N_334,In_233,In_1948);
and U335 (N_335,In_1268,In_331);
xor U336 (N_336,In_1971,In_586);
nor U337 (N_337,In_1188,In_1706);
or U338 (N_338,In_1564,In_1519);
xor U339 (N_339,In_619,In_2270);
or U340 (N_340,In_763,In_1535);
and U341 (N_341,In_12,In_1993);
nand U342 (N_342,In_279,In_614);
nand U343 (N_343,In_2218,In_88);
and U344 (N_344,In_1814,In_1280);
nand U345 (N_345,In_1469,In_1622);
or U346 (N_346,In_914,In_1388);
xnor U347 (N_347,In_1346,In_896);
nand U348 (N_348,In_1698,In_707);
nor U349 (N_349,In_1794,In_2308);
or U350 (N_350,In_17,In_1689);
nand U351 (N_351,In_2318,In_583);
nand U352 (N_352,In_2488,In_569);
and U353 (N_353,In_71,In_1484);
nand U354 (N_354,In_1561,In_2121);
nor U355 (N_355,In_246,In_364);
nor U356 (N_356,In_302,In_293);
nor U357 (N_357,In_2135,In_920);
or U358 (N_358,In_2108,In_297);
xor U359 (N_359,In_1779,In_693);
and U360 (N_360,In_864,In_2001);
nand U361 (N_361,In_838,In_82);
nor U362 (N_362,In_263,In_396);
or U363 (N_363,In_1385,In_1166);
and U364 (N_364,In_1437,In_2209);
or U365 (N_365,In_1977,In_92);
and U366 (N_366,In_672,In_592);
nor U367 (N_367,In_743,In_928);
xor U368 (N_368,In_2362,In_997);
nor U369 (N_369,In_1653,In_2055);
xor U370 (N_370,In_344,In_119);
nor U371 (N_371,In_1523,In_856);
nand U372 (N_372,In_1628,In_1514);
or U373 (N_373,In_1701,In_2289);
nand U374 (N_374,In_618,In_791);
nand U375 (N_375,In_1293,In_1440);
or U376 (N_376,In_440,In_2406);
nand U377 (N_377,In_2379,In_62);
or U378 (N_378,In_1343,In_1629);
nand U379 (N_379,In_2241,In_13);
xnor U380 (N_380,In_1231,In_1439);
and U381 (N_381,In_857,In_1238);
and U382 (N_382,In_1374,In_2217);
and U383 (N_383,In_333,In_1160);
and U384 (N_384,In_572,In_1227);
nor U385 (N_385,In_2457,In_1733);
and U386 (N_386,In_464,In_824);
and U387 (N_387,In_831,In_521);
or U388 (N_388,In_1131,In_744);
xor U389 (N_389,In_24,In_511);
xnor U390 (N_390,In_66,In_74);
xor U391 (N_391,In_2361,In_2495);
and U392 (N_392,In_459,In_355);
or U393 (N_393,In_2381,In_1959);
xnor U394 (N_394,In_2168,In_1143);
nor U395 (N_395,In_510,In_2154);
nor U396 (N_396,In_416,In_727);
or U397 (N_397,In_1164,In_1967);
xnor U398 (N_398,In_20,In_300);
xnor U399 (N_399,In_1321,In_475);
and U400 (N_400,In_1398,In_839);
or U401 (N_401,In_288,In_1868);
nor U402 (N_402,In_1065,In_1541);
nand U403 (N_403,In_1893,In_2025);
nand U404 (N_404,In_371,In_1481);
xnor U405 (N_405,In_1059,In_0);
and U406 (N_406,In_1244,In_1758);
nand U407 (N_407,In_1081,In_1810);
and U408 (N_408,In_1888,In_103);
nand U409 (N_409,In_2298,In_2171);
nand U410 (N_410,In_1416,In_1825);
and U411 (N_411,In_561,In_156);
nand U412 (N_412,In_770,In_129);
nor U413 (N_413,In_240,In_988);
or U414 (N_414,In_2110,In_1401);
nor U415 (N_415,In_875,In_1117);
xor U416 (N_416,In_1645,In_216);
xor U417 (N_417,In_1537,In_1639);
xnor U418 (N_418,In_241,In_2157);
nand U419 (N_419,In_930,In_1943);
xor U420 (N_420,In_2065,In_433);
nand U421 (N_421,In_176,In_517);
xor U422 (N_422,In_2033,In_786);
and U423 (N_423,In_2003,In_2232);
xor U424 (N_424,In_921,In_2060);
nor U425 (N_425,In_2231,In_487);
xor U426 (N_426,In_1362,In_1760);
and U427 (N_427,In_789,In_163);
xor U428 (N_428,In_1461,In_1183);
and U429 (N_429,In_461,In_1203);
nand U430 (N_430,In_1543,In_823);
and U431 (N_431,In_1339,In_793);
and U432 (N_432,In_501,In_637);
and U433 (N_433,In_2084,In_902);
xor U434 (N_434,In_829,In_943);
and U435 (N_435,In_187,In_265);
and U436 (N_436,In_399,In_1904);
nor U437 (N_437,In_1532,In_1821);
nand U438 (N_438,In_885,In_1676);
nor U439 (N_439,In_89,In_2269);
xor U440 (N_440,In_1375,In_2450);
xnor U441 (N_441,In_2314,In_2165);
xnor U442 (N_442,In_2090,In_1926);
or U443 (N_443,In_1955,In_1945);
and U444 (N_444,In_1226,In_2418);
and U445 (N_445,In_859,In_99);
nor U446 (N_446,In_992,In_1761);
nand U447 (N_447,In_2369,In_589);
or U448 (N_448,In_310,In_908);
and U449 (N_449,In_75,In_33);
nor U450 (N_450,In_1635,In_169);
or U451 (N_451,In_1190,In_878);
and U452 (N_452,In_1515,In_166);
and U453 (N_453,In_140,In_2273);
or U454 (N_454,In_236,In_1667);
or U455 (N_455,In_1051,In_1179);
nor U456 (N_456,In_218,In_2313);
xor U457 (N_457,In_2249,In_2340);
or U458 (N_458,In_431,In_1897);
nor U459 (N_459,In_661,In_1242);
nand U460 (N_460,In_704,In_1446);
or U461 (N_461,In_702,In_785);
and U462 (N_462,In_1681,In_800);
or U463 (N_463,In_2458,In_2351);
nor U464 (N_464,In_2323,In_983);
or U465 (N_465,In_1121,In_1287);
nor U466 (N_466,In_130,In_1080);
xnor U467 (N_467,In_185,In_1973);
or U468 (N_468,In_830,In_2377);
and U469 (N_469,In_2211,In_764);
nor U470 (N_470,In_484,In_966);
or U471 (N_471,In_1116,In_540);
nand U472 (N_472,In_446,In_1576);
or U473 (N_473,In_341,In_1300);
xor U474 (N_474,In_804,In_1091);
and U475 (N_475,In_412,In_923);
xor U476 (N_476,In_78,In_363);
or U477 (N_477,In_247,In_1920);
nor U478 (N_478,In_1640,In_726);
nand U479 (N_479,In_1838,In_1901);
and U480 (N_480,In_2156,In_1367);
or U481 (N_481,In_806,In_1096);
xnor U482 (N_482,In_2142,In_2238);
or U483 (N_483,In_73,In_1807);
or U484 (N_484,In_1933,In_373);
nor U485 (N_485,In_1006,In_1041);
nand U486 (N_486,In_1358,In_1874);
xnor U487 (N_487,In_2354,In_748);
nand U488 (N_488,In_1400,In_113);
and U489 (N_489,In_2201,In_597);
or U490 (N_490,In_777,In_1999);
nor U491 (N_491,In_173,In_1585);
nor U492 (N_492,In_1795,In_322);
and U493 (N_493,In_1542,In_1470);
or U494 (N_494,In_2053,In_2437);
nand U495 (N_495,In_69,In_228);
or U496 (N_496,In_2292,In_1239);
nor U497 (N_497,In_2192,In_141);
or U498 (N_498,In_2372,In_1251);
xnor U499 (N_499,In_2052,In_1003);
or U500 (N_500,In_901,In_191);
nor U501 (N_501,In_1675,In_2022);
xor U502 (N_502,In_1278,In_642);
nor U503 (N_503,In_90,In_2047);
or U504 (N_504,In_709,In_1552);
nand U505 (N_505,In_2339,In_503);
and U506 (N_506,In_1387,In_104);
or U507 (N_507,In_924,In_1325);
nand U508 (N_508,In_2176,In_658);
nand U509 (N_509,In_1504,In_1019);
or U510 (N_510,In_1784,In_2255);
or U511 (N_511,In_1386,In_1397);
and U512 (N_512,In_362,In_1344);
and U513 (N_513,In_245,In_1330);
nor U514 (N_514,In_329,In_1097);
nor U515 (N_515,In_822,In_858);
nand U516 (N_516,In_1749,In_1033);
xnor U517 (N_517,In_2006,In_2240);
and U518 (N_518,In_1323,In_1513);
and U519 (N_519,In_1742,In_1949);
xor U520 (N_520,In_2336,In_932);
nor U521 (N_521,In_2202,In_2063);
and U522 (N_522,In_2199,In_168);
nor U523 (N_523,In_2293,In_895);
and U524 (N_524,In_706,In_1983);
and U525 (N_525,In_552,In_1037);
nand U526 (N_526,In_194,In_1835);
xor U527 (N_527,In_1392,In_1101);
and U528 (N_528,In_485,In_1480);
nor U529 (N_529,In_625,In_1985);
xor U530 (N_530,In_2214,In_964);
and U531 (N_531,In_2261,In_1335);
xnor U532 (N_532,In_154,In_65);
xor U533 (N_533,In_515,In_1666);
or U534 (N_534,In_611,In_1248);
and U535 (N_535,In_23,In_258);
and U536 (N_536,In_695,In_200);
nor U537 (N_537,In_1279,In_1654);
and U538 (N_538,In_1373,In_1348);
nor U539 (N_539,In_2032,In_2454);
xor U540 (N_540,In_2460,In_1927);
and U541 (N_541,In_146,In_1790);
and U542 (N_542,In_2449,In_2076);
xnor U543 (N_543,In_213,In_83);
xnor U544 (N_544,In_766,In_238);
nand U545 (N_545,In_1913,In_2334);
nand U546 (N_546,In_193,In_1438);
and U547 (N_547,In_1297,In_1023);
or U548 (N_548,In_1086,In_1288);
nor U549 (N_549,In_32,In_226);
or U550 (N_550,In_1855,In_347);
and U551 (N_551,In_1705,In_2416);
or U552 (N_552,In_50,In_1247);
nand U553 (N_553,In_2433,In_2307);
or U554 (N_554,In_2422,In_225);
and U555 (N_555,In_242,In_615);
xnor U556 (N_556,In_2194,In_1414);
nand U557 (N_557,In_1725,In_1726);
nor U558 (N_558,In_1299,In_231);
nor U559 (N_559,In_1237,In_1533);
nor U560 (N_560,In_328,In_132);
nand U561 (N_561,In_2179,In_735);
and U562 (N_562,In_1357,In_2101);
nand U563 (N_563,In_415,In_969);
and U564 (N_564,In_36,In_2467);
nand U565 (N_565,In_2094,In_813);
nand U566 (N_566,In_946,In_473);
nand U567 (N_567,In_1728,In_627);
and U568 (N_568,In_1114,In_1005);
or U569 (N_569,In_1732,In_711);
nand U570 (N_570,In_564,In_2497);
xor U571 (N_571,In_1291,In_165);
nor U572 (N_572,In_593,In_861);
xnor U573 (N_573,In_585,In_1092);
nor U574 (N_574,In_1984,In_1327);
nor U575 (N_575,In_1846,In_609);
nor U576 (N_576,In_1136,In_1456);
nand U577 (N_577,In_1412,In_1516);
or U578 (N_578,In_941,In_301);
or U579 (N_579,In_1644,In_666);
or U580 (N_580,In_1266,In_546);
or U581 (N_581,In_64,In_2216);
xor U582 (N_582,In_1109,In_1696);
or U583 (N_583,In_136,In_1755);
or U584 (N_584,In_538,In_910);
or U585 (N_585,In_2254,In_392);
nor U586 (N_586,In_684,In_212);
and U587 (N_587,In_1648,In_669);
xnor U588 (N_588,In_1320,In_933);
or U589 (N_589,In_421,In_1885);
xor U590 (N_590,In_377,In_1507);
nand U591 (N_591,In_2382,In_378);
or U592 (N_592,In_1433,In_1350);
nor U593 (N_593,In_1593,In_1110);
nand U594 (N_594,In_1660,In_97);
and U595 (N_595,In_1427,In_1816);
or U596 (N_596,In_1313,In_922);
or U597 (N_597,In_417,In_1269);
nor U598 (N_598,In_116,In_1365);
or U599 (N_599,In_499,In_54);
nor U600 (N_600,In_681,In_2239);
nor U601 (N_601,In_1918,In_311);
xor U602 (N_602,In_916,In_1271);
or U603 (N_603,In_2153,In_2017);
nor U604 (N_604,In_1256,In_2271);
nor U605 (N_605,In_1497,In_428);
and U606 (N_606,In_679,In_1273);
nand U607 (N_607,In_2088,In_2161);
nor U608 (N_608,In_1077,In_1115);
nor U609 (N_609,In_2327,In_2321);
xor U610 (N_610,In_320,In_419);
nor U611 (N_611,In_1869,In_1907);
xnor U612 (N_612,In_1318,In_269);
and U613 (N_613,In_1031,In_161);
xnor U614 (N_614,In_305,In_647);
nor U615 (N_615,In_1947,In_613);
xor U616 (N_616,In_1370,In_1803);
and U617 (N_617,In_2256,In_506);
and U618 (N_618,In_1230,In_234);
and U619 (N_619,In_1463,In_2331);
nand U620 (N_620,In_840,In_818);
and U621 (N_621,In_369,In_833);
xor U622 (N_622,In_1769,In_1583);
xnor U623 (N_623,In_686,In_795);
nor U624 (N_624,In_1048,In_874);
or U625 (N_625,In_2124,In_1173);
or U626 (N_626,In_1026,In_1994);
and U627 (N_627,In_1841,In_2115);
and U628 (N_628,In_1146,In_268);
nor U629 (N_629,In_1,In_152);
or U630 (N_630,In_1536,In_2093);
and U631 (N_631,In_1140,In_2474);
and U632 (N_632,In_2446,In_2287);
or U633 (N_633,In_2152,In_160);
xor U634 (N_634,In_528,In_1180);
or U635 (N_635,In_1032,In_603);
or U636 (N_636,In_847,In_1319);
xor U637 (N_637,In_1529,In_1496);
xor U638 (N_638,In_1035,In_1303);
nor U639 (N_639,In_976,In_1739);
nand U640 (N_640,In_773,In_722);
nand U641 (N_641,In_2356,In_513);
nand U642 (N_642,In_436,In_2081);
or U643 (N_643,In_575,In_255);
and U644 (N_644,In_814,In_1522);
nor U645 (N_645,In_2322,In_834);
nor U646 (N_646,In_197,In_1351);
nor U647 (N_647,In_1076,In_25);
nand U648 (N_648,In_1122,In_2233);
xor U649 (N_649,In_2357,In_1214);
nand U650 (N_650,In_2014,In_474);
xnor U651 (N_651,In_2000,In_1752);
xnor U652 (N_652,In_1316,In_756);
nand U653 (N_653,In_1968,In_2205);
and U654 (N_654,In_1573,In_352);
nor U655 (N_655,In_974,In_962);
and U656 (N_656,In_1734,In_2167);
xnor U657 (N_657,In_2215,In_1559);
or U658 (N_658,In_1442,In_9);
and U659 (N_659,In_1785,In_1953);
or U660 (N_660,In_1326,In_670);
nand U661 (N_661,In_148,In_2300);
nor U662 (N_662,In_2316,In_46);
xnor U663 (N_663,In_249,In_787);
xor U664 (N_664,In_1441,In_2244);
and U665 (N_665,In_760,In_2070);
nand U666 (N_666,In_2250,In_2264);
and U667 (N_667,In_1754,In_2395);
and U668 (N_668,In_1342,In_1207);
nor U669 (N_669,In_1987,In_2338);
or U670 (N_670,In_519,In_2346);
or U671 (N_671,In_486,In_608);
nand U672 (N_672,In_57,In_700);
or U673 (N_673,In_2309,In_730);
or U674 (N_674,In_1406,In_1134);
or U675 (N_675,In_845,In_1213);
nor U676 (N_676,In_2228,In_2089);
and U677 (N_677,In_554,In_2276);
nand U678 (N_678,In_755,In_1836);
nand U679 (N_679,In_1148,In_1053);
nor U680 (N_680,In_1688,In_2431);
nor U681 (N_681,In_1209,In_1224);
nand U682 (N_682,In_1123,In_2397);
nor U683 (N_683,In_1240,In_182);
and U684 (N_684,In_1562,In_2432);
or U685 (N_685,In_39,In_1499);
nand U686 (N_686,In_1359,In_79);
or U687 (N_687,In_1765,In_879);
nand U688 (N_688,In_1312,In_1153);
and U689 (N_689,In_1356,In_2151);
or U690 (N_690,In_1154,In_1787);
nand U691 (N_691,In_1691,In_1069);
xor U692 (N_692,In_1876,In_852);
nor U693 (N_693,In_139,In_612);
and U694 (N_694,In_601,In_219);
and U695 (N_695,In_388,In_308);
nand U696 (N_696,In_1652,In_1137);
nand U697 (N_697,In_384,In_1797);
nor U698 (N_698,In_2341,In_51);
or U699 (N_699,In_426,In_1408);
and U700 (N_700,In_1264,In_1982);
xor U701 (N_701,In_1417,In_595);
nand U702 (N_702,In_365,In_158);
or U703 (N_703,In_2342,In_289);
xor U704 (N_704,In_1471,In_162);
and U705 (N_705,In_2388,In_2183);
nor U706 (N_706,In_1338,In_137);
or U707 (N_707,In_1986,In_393);
nand U708 (N_708,In_1310,In_14);
nand U709 (N_709,In_1638,In_253);
nand U710 (N_710,In_1783,In_1212);
nor U711 (N_711,In_2144,In_576);
nand U712 (N_712,In_287,In_757);
nand U713 (N_713,In_1518,In_186);
or U714 (N_714,In_1491,In_1883);
or U715 (N_715,In_1763,In_1254);
and U716 (N_716,In_2062,In_671);
nand U717 (N_717,In_550,In_1894);
nor U718 (N_718,In_2031,In_470);
nand U719 (N_719,In_2411,In_479);
nor U720 (N_720,In_1952,In_1712);
xor U721 (N_721,In_2414,In_1837);
xor U722 (N_722,In_1620,In_420);
nand U723 (N_723,In_127,In_1886);
nor U724 (N_724,In_423,In_1729);
or U725 (N_725,In_1770,In_2164);
xor U726 (N_726,In_2391,In_1619);
xnor U727 (N_727,In_2008,In_1025);
nand U728 (N_728,In_1413,In_2077);
nand U729 (N_729,In_701,In_998);
nor U730 (N_730,In_1464,In_171);
xor U731 (N_731,In_1444,In_1538);
nor U732 (N_732,In_441,In_1615);
xor U733 (N_733,In_1938,In_1609);
or U734 (N_734,In_1646,In_919);
or U735 (N_735,In_1793,In_1211);
and U736 (N_736,In_1389,In_1294);
nand U737 (N_737,In_2359,In_972);
xor U738 (N_738,In_1208,In_1161);
nor U739 (N_739,In_713,In_599);
xnor U740 (N_740,In_1394,In_1856);
nand U741 (N_741,In_2487,In_2483);
nor U742 (N_742,In_81,In_956);
and U743 (N_743,In_1702,In_2365);
or U744 (N_744,In_680,In_149);
nor U745 (N_745,In_1436,In_1588);
nor U746 (N_746,In_114,In_1572);
nor U747 (N_747,In_1822,In_1128);
or U748 (N_748,In_1024,In_201);
nand U749 (N_749,In_2136,In_244);
nor U750 (N_750,In_1840,In_482);
or U751 (N_751,In_2018,In_1906);
xor U752 (N_752,In_1862,In_1403);
nor U753 (N_753,In_2145,In_2190);
nor U754 (N_754,In_667,In_535);
or U755 (N_755,In_1296,In_170);
nor U756 (N_756,In_2073,In_1455);
nand U757 (N_757,In_545,In_2410);
xor U758 (N_758,In_1699,In_955);
nor U759 (N_759,In_1205,In_1857);
and U760 (N_760,In_1447,In_1171);
nor U761 (N_761,In_338,In_548);
or U762 (N_762,In_2170,In_2484);
and U763 (N_763,In_1104,In_1780);
and U764 (N_764,In_223,In_493);
and U765 (N_765,In_1511,In_1545);
and U766 (N_766,In_1687,In_1685);
or U767 (N_767,In_685,In_1683);
xor U768 (N_768,In_1498,In_1250);
and U769 (N_769,In_541,In_1789);
xnor U770 (N_770,In_1322,In_1843);
nand U771 (N_771,In_215,In_1361);
nand U772 (N_772,In_2029,In_204);
or U773 (N_773,In_639,In_2274);
nand U774 (N_774,In_327,In_2105);
or U775 (N_775,In_383,In_110);
xor U776 (N_776,In_144,In_659);
or U777 (N_777,In_1990,In_2061);
or U778 (N_778,In_142,In_108);
xnor U779 (N_779,In_434,In_1159);
nor U780 (N_780,In_624,In_652);
nand U781 (N_781,In_1384,In_430);
nand U782 (N_782,In_1521,In_2425);
xor U783 (N_783,In_1756,In_2333);
xor U784 (N_784,In_1219,In_1089);
or U785 (N_785,In_1633,In_580);
and U786 (N_786,In_957,In_1798);
or U787 (N_787,In_1612,In_385);
nor U788 (N_788,In_1366,In_1867);
or U789 (N_789,In_1604,In_22);
xor U790 (N_790,In_1899,In_542);
or U791 (N_791,In_367,In_299);
or U792 (N_792,In_2128,In_911);
or U793 (N_793,In_1328,In_1976);
or U794 (N_794,In_1267,In_1902);
or U795 (N_795,In_846,In_2419);
or U796 (N_796,In_381,In_636);
and U797 (N_797,In_1738,In_153);
nand U798 (N_798,In_1762,In_1158);
or U799 (N_799,In_2413,In_1502);
or U800 (N_800,In_1257,In_1792);
or U801 (N_801,In_2155,In_1057);
or U802 (N_802,In_1261,In_747);
nand U803 (N_803,In_2227,In_673);
or U804 (N_804,In_1292,In_1878);
nand U805 (N_805,In_1673,In_1565);
xnor U806 (N_806,In_1138,In_2141);
xnor U807 (N_807,In_1896,In_1574);
or U808 (N_808,In_676,In_808);
nand U809 (N_809,In_1286,In_395);
nor U810 (N_810,In_275,In_358);
nor U811 (N_811,In_1220,In_1668);
and U812 (N_812,In_1528,In_1656);
or U813 (N_813,In_1954,In_1802);
or U814 (N_814,In_714,In_174);
xor U815 (N_815,In_1170,In_1775);
nor U816 (N_816,In_1555,In_1002);
nor U817 (N_817,In_488,In_1155);
or U818 (N_818,In_312,In_1093);
or U819 (N_819,In_2222,In_881);
and U820 (N_820,In_1072,In_1301);
or U821 (N_821,In_664,In_2091);
nand U822 (N_822,In_1275,In_1187);
or U823 (N_823,In_1568,In_2471);
nand U824 (N_824,In_10,In_848);
nand U825 (N_825,In_574,In_1800);
or U826 (N_826,In_590,In_55);
nor U827 (N_827,In_444,In_85);
and U828 (N_828,In_1493,In_1905);
xnor U829 (N_829,In_1946,In_1589);
and U830 (N_830,In_445,In_2);
nor U831 (N_831,In_1587,In_1483);
nor U832 (N_832,In_1249,In_2258);
or U833 (N_833,In_1625,In_961);
xnor U834 (N_834,In_991,In_2286);
and U835 (N_835,In_1937,In_1329);
xor U836 (N_836,In_422,In_357);
and U837 (N_837,In_1430,In_1998);
or U838 (N_838,In_409,In_437);
xor U839 (N_839,In_1029,In_2493);
and U840 (N_840,In_1141,In_888);
or U841 (N_841,In_1634,In_2219);
nor U842 (N_842,In_1253,In_180);
nand U843 (N_843,In_272,In_2013);
and U844 (N_844,In_720,In_284);
and U845 (N_845,In_868,In_665);
nor U846 (N_846,In_1820,In_1206);
and U847 (N_847,In_44,In_1826);
nand U848 (N_848,In_1204,In_2445);
xnor U849 (N_849,In_1833,In_224);
and U850 (N_850,In_2235,In_2200);
or U851 (N_851,In_1431,In_318);
xor U852 (N_852,In_1995,In_2020);
xor U853 (N_853,In_1847,In_566);
or U854 (N_854,In_2328,In_1679);
nand U855 (N_855,In_4,In_853);
and U856 (N_856,In_1895,In_1252);
xor U857 (N_857,In_1113,In_990);
and U858 (N_858,In_2326,In_2288);
and U859 (N_859,In_1544,In_2079);
xnor U860 (N_860,In_1557,In_900);
and U861 (N_861,In_1965,In_2050);
or U862 (N_862,In_2263,In_723);
and U863 (N_863,In_1028,In_2259);
nand U864 (N_864,In_72,In_779);
or U865 (N_865,In_2095,In_1601);
xor U866 (N_866,In_1602,In_570);
nand U867 (N_867,In_1478,In_1737);
and U868 (N_868,In_1746,In_1334);
nand U869 (N_869,In_18,In_2252);
or U870 (N_870,In_273,In_2019);
nor U871 (N_871,In_622,In_1290);
xor U872 (N_872,In_740,In_1085);
or U873 (N_873,In_1324,In_2010);
xor U874 (N_874,In_206,In_481);
or U875 (N_875,In_1295,In_1839);
and U876 (N_876,In_1174,In_520);
nand U877 (N_877,In_931,In_1079);
xor U878 (N_878,In_28,In_891);
nor U879 (N_879,In_2353,In_2163);
nor U880 (N_880,In_1468,In_361);
nand U881 (N_881,In_208,In_1001);
xor U882 (N_882,In_2005,In_490);
or U883 (N_883,In_1308,In_2443);
nand U884 (N_884,In_1162,In_1489);
nand U885 (N_885,In_1854,In_2392);
or U886 (N_886,In_1465,In_596);
nand U887 (N_887,In_1960,In_641);
xor U888 (N_888,In_1850,In_604);
and U889 (N_889,In_1736,In_565);
nand U890 (N_890,In_1125,In_1771);
or U891 (N_891,In_2195,In_1711);
xnor U892 (N_892,In_1197,In_145);
nand U893 (N_893,In_1087,In_5);
and U894 (N_894,In_1944,In_1508);
and U895 (N_895,In_2147,In_582);
xnor U896 (N_896,In_271,In_1626);
nor U897 (N_897,In_781,In_425);
nor U898 (N_898,In_980,In_2158);
nor U899 (N_899,In_1939,In_579);
or U900 (N_900,In_1304,In_560);
nor U901 (N_901,In_2402,In_492);
and U902 (N_902,In_465,In_157);
and U903 (N_903,In_1118,In_2143);
or U904 (N_904,In_1000,In_2401);
or U905 (N_905,In_42,In_351);
and U906 (N_906,In_737,In_682);
and U907 (N_907,In_516,In_1571);
xnor U908 (N_908,In_1165,In_250);
nand U909 (N_909,In_2198,In_1466);
nor U910 (N_910,In_43,In_178);
and U911 (N_911,In_405,In_628);
nor U912 (N_912,In_1915,In_2159);
and U913 (N_913,In_2224,In_797);
xnor U914 (N_914,In_1703,In_1082);
and U915 (N_915,In_2246,In_1546);
nor U916 (N_916,In_449,In_2435);
or U917 (N_917,In_1831,In_855);
nand U918 (N_918,In_1777,In_1692);
nand U919 (N_919,In_1695,In_783);
and U920 (N_920,In_1776,In_581);
and U921 (N_921,In_559,In_254);
and U922 (N_922,In_2499,In_587);
nand U923 (N_923,In_691,In_1582);
and U924 (N_924,In_2011,In_563);
nand U925 (N_925,In_2140,In_438);
or U926 (N_926,In_837,In_1402);
nand U927 (N_927,In_1858,In_690);
and U928 (N_928,In_2489,In_1503);
or U929 (N_929,In_1925,In_2320);
nand U930 (N_930,In_457,In_936);
nor U931 (N_931,In_968,In_1064);
nand U932 (N_932,In_198,In_429);
nor U933 (N_933,In_2490,In_819);
nor U934 (N_934,In_549,In_418);
and U935 (N_935,In_1067,In_2023);
or U936 (N_936,In_2098,In_1929);
and U937 (N_937,In_640,In_1581);
nand U938 (N_938,In_1730,In_1517);
nor U939 (N_939,In_1972,In_512);
or U940 (N_940,In_2127,In_1135);
or U941 (N_941,In_674,In_2119);
nor U942 (N_942,In_2468,In_675);
nor U943 (N_943,In_765,In_1928);
xor U944 (N_944,In_1477,In_261);
xor U945 (N_945,In_379,In_944);
xnor U946 (N_946,In_1061,In_221);
or U947 (N_947,In_2375,In_2374);
nand U948 (N_948,In_469,In_1584);
or U949 (N_949,In_2459,In_2456);
nand U950 (N_950,In_413,In_463);
or U951 (N_951,In_796,In_2404);
nor U952 (N_952,In_2213,In_543);
and U953 (N_953,In_1482,In_1054);
nor U954 (N_954,In_1345,In_2146);
nor U955 (N_955,In_2329,In_164);
xor U956 (N_956,In_1950,In_1147);
xor U957 (N_957,In_893,In_1980);
nand U958 (N_958,In_705,In_1715);
nor U959 (N_959,In_877,In_949);
nand U960 (N_960,In_607,In_1796);
or U961 (N_961,In_1124,In_2034);
nor U962 (N_962,In_1586,In_703);
or U963 (N_963,In_854,In_1665);
xor U964 (N_964,In_533,In_1349);
nor U965 (N_965,In_1611,In_94);
nand U966 (N_966,In_712,In_120);
and U967 (N_967,In_1512,In_235);
or U968 (N_968,In_536,In_1751);
nor U969 (N_969,In_2148,In_280);
nor U970 (N_970,In_2399,In_1352);
xor U971 (N_971,In_1425,In_1007);
nand U972 (N_972,In_810,In_2197);
and U973 (N_973,In_68,In_2028);
nor U974 (N_974,In_1799,In_494);
or U975 (N_975,In_1210,In_2189);
xor U976 (N_976,In_1773,In_1347);
and U977 (N_977,In_1534,In_1978);
or U978 (N_978,In_650,In_1315);
and U979 (N_979,In_568,In_295);
nand U980 (N_980,In_1607,In_1152);
or U981 (N_981,In_870,In_2378);
or U982 (N_982,In_2371,In_771);
and U983 (N_983,In_2291,In_2044);
nor U984 (N_984,In_497,In_1873);
nand U985 (N_985,In_2132,In_1713);
or U986 (N_986,In_274,In_1144);
xor U987 (N_987,In_668,In_500);
xor U988 (N_988,In_1621,In_1368);
or U989 (N_989,In_1120,In_907);
or U990 (N_990,In_239,In_708);
nand U991 (N_991,In_1613,In_1661);
xnor U992 (N_992,In_2248,In_1015);
xor U993 (N_993,In_663,In_655);
nand U994 (N_994,In_227,In_1399);
xor U995 (N_995,In_77,In_835);
xnor U996 (N_996,In_2461,In_1381);
nor U997 (N_997,In_337,In_2285);
and U998 (N_998,In_256,In_873);
nand U999 (N_999,In_1010,In_1066);
nand U1000 (N_1000,In_892,In_45);
xor U1001 (N_1001,In_52,In_836);
or U1002 (N_1002,In_1979,In_975);
or U1003 (N_1003,In_277,In_698);
or U1004 (N_1004,In_1556,In_2160);
and U1005 (N_1005,In_2186,In_2462);
and U1006 (N_1006,In_683,In_1298);
xor U1007 (N_1007,In_1942,In_1126);
xor U1008 (N_1008,In_1963,In_2203);
and U1009 (N_1009,In_2403,In_107);
nand U1010 (N_1010,In_2004,In_2086);
nand U1011 (N_1011,In_410,In_2104);
nand U1012 (N_1012,In_1099,In_2475);
xor U1013 (N_1013,In_2253,In_1172);
xnor U1014 (N_1014,In_2054,In_1727);
xor U1015 (N_1015,In_220,In_40);
xnor U1016 (N_1016,In_938,In_985);
nor U1017 (N_1017,In_134,In_626);
nand U1018 (N_1018,In_525,In_2225);
and U1019 (N_1019,In_1149,In_2139);
nor U1020 (N_1020,In_1956,In_1393);
xnor U1021 (N_1021,In_1866,In_696);
and U1022 (N_1022,In_820,In_2439);
nor U1023 (N_1023,In_402,In_1525);
nor U1024 (N_1024,In_1812,In_183);
or U1025 (N_1025,In_1222,In_2302);
xnor U1026 (N_1026,In_1063,In_1817);
and U1027 (N_1027,In_817,In_544);
xor U1028 (N_1028,In_1139,In_1697);
nor U1029 (N_1029,In_718,In_1151);
xor U1030 (N_1030,In_1603,In_2009);
xnor U1031 (N_1031,In_2106,In_1263);
nand U1032 (N_1032,In_1597,In_2363);
nor U1033 (N_1033,In_1056,In_2178);
xnor U1034 (N_1034,In_1919,In_2123);
nand U1035 (N_1035,In_632,In_699);
xnor U1036 (N_1036,In_1178,In_442);
or U1037 (N_1037,In_1030,In_1834);
xnor U1038 (N_1038,In_188,In_286);
or U1039 (N_1039,In_687,In_348);
nor U1040 (N_1040,In_925,In_1467);
or U1041 (N_1041,In_531,In_621);
nor U1042 (N_1042,In_447,In_458);
and U1043 (N_1043,In_1642,In_2348);
nor U1044 (N_1044,In_1829,In_1704);
nor U1045 (N_1045,In_633,In_588);
or U1046 (N_1046,In_573,In_325);
and U1047 (N_1047,In_1540,In_816);
nor U1048 (N_1048,In_1419,In_1176);
nor U1049 (N_1049,In_1887,In_439);
nand U1050 (N_1050,In_1276,In_736);
nand U1051 (N_1051,In_917,In_2036);
nand U1052 (N_1052,In_1450,In_56);
xnor U1053 (N_1053,In_2064,In_353);
or U1054 (N_1054,In_58,In_2137);
and U1055 (N_1055,In_1710,In_2181);
or U1056 (N_1056,In_2265,In_945);
nand U1057 (N_1057,In_2344,In_1094);
xor U1058 (N_1058,In_821,In_2477);
or U1059 (N_1059,In_1027,In_1396);
and U1060 (N_1060,In_1157,In_98);
nor U1061 (N_1061,In_2347,In_2125);
nor U1062 (N_1062,In_2043,In_645);
and U1063 (N_1063,In_2355,In_35);
or U1064 (N_1064,In_798,In_2260);
or U1065 (N_1065,In_237,In_509);
nand U1066 (N_1066,In_2049,In_634);
and U1067 (N_1067,In_1163,In_2173);
and U1068 (N_1068,In_489,In_1262);
or U1069 (N_1069,In_805,In_1962);
nor U1070 (N_1070,In_959,In_314);
and U1071 (N_1071,In_1432,In_476);
nor U1072 (N_1072,In_801,In_989);
or U1073 (N_1073,In_843,In_406);
or U1074 (N_1074,In_370,In_1305);
and U1075 (N_1075,In_1073,In_2387);
or U1076 (N_1076,In_1457,In_934);
nand U1077 (N_1077,In_2358,In_495);
or U1078 (N_1078,In_643,In_2412);
nand U1079 (N_1079,In_167,In_1669);
nor U1080 (N_1080,In_211,In_2389);
nor U1081 (N_1081,In_189,In_109);
xnor U1082 (N_1082,In_1011,In_1849);
nor U1083 (N_1083,In_276,In_880);
and U1084 (N_1084,In_2337,In_315);
xor U1085 (N_1085,In_1234,In_359);
nand U1086 (N_1086,In_1614,In_871);
xnor U1087 (N_1087,In_1708,In_1488);
nand U1088 (N_1088,In_2496,In_790);
or U1089 (N_1089,In_1720,In_1558);
nand U1090 (N_1090,In_1863,In_1881);
nand U1091 (N_1091,In_317,In_1353);
and U1092 (N_1092,In_555,In_319);
nor U1093 (N_1093,In_48,In_1898);
and U1094 (N_1094,In_1167,In_1217);
and U1095 (N_1095,In_1566,In_2162);
or U1096 (N_1096,In_1272,In_2041);
nand U1097 (N_1097,In_2175,In_1509);
nand U1098 (N_1098,In_2040,In_2398);
nand U1099 (N_1099,In_2430,In_196);
and U1100 (N_1100,In_2492,In_1476);
xor U1101 (N_1101,In_507,In_1961);
nor U1102 (N_1102,In_2279,In_610);
nand U1103 (N_1103,In_594,In_16);
and U1104 (N_1104,In_6,In_260);
or U1105 (N_1105,In_1245,In_623);
and U1106 (N_1106,In_1043,In_195);
or U1107 (N_1107,In_1767,In_1487);
nor U1108 (N_1108,In_257,In_1068);
and U1109 (N_1109,In_303,In_947);
xnor U1110 (N_1110,In_884,In_232);
nand U1111 (N_1111,In_863,In_1936);
xor U1112 (N_1112,In_1718,In_151);
xor U1113 (N_1113,In_1889,In_1664);
nor U1114 (N_1114,In_1550,In_2319);
nand U1115 (N_1115,In_887,In_1610);
nor U1116 (N_1116,In_1774,In_1363);
and U1117 (N_1117,In_721,In_455);
or U1118 (N_1118,In_1331,In_2220);
and U1119 (N_1119,In_1228,In_1554);
and U1120 (N_1120,In_1410,In_1083);
or U1121 (N_1121,In_496,In_1577);
xor U1122 (N_1122,In_387,In_970);
xor U1123 (N_1123,In_537,In_1014);
nand U1124 (N_1124,In_1662,In_472);
nand U1125 (N_1125,In_1500,In_1506);
or U1126 (N_1126,In_1808,In_1202);
nand U1127 (N_1127,In_1875,In_38);
xnor U1128 (N_1128,In_1818,In_159);
xor U1129 (N_1129,In_1671,In_1426);
and U1130 (N_1130,In_827,In_93);
and U1131 (N_1131,In_63,In_1912);
nand U1132 (N_1132,In_929,In_304);
xnor U1133 (N_1133,In_11,In_688);
and U1134 (N_1134,In_1674,In_262);
and U1135 (N_1135,In_382,In_1309);
xor U1136 (N_1136,In_330,In_1052);
nand U1137 (N_1137,In_2424,In_147);
and U1138 (N_1138,In_2037,In_1900);
nor U1139 (N_1139,In_401,In_1045);
nand U1140 (N_1140,In_1429,In_754);
or U1141 (N_1141,In_2428,In_1934);
nand U1142 (N_1142,In_452,In_950);
nand U1143 (N_1143,In_2083,In_2470);
nand U1144 (N_1144,In_123,In_890);
nand U1145 (N_1145,In_2185,In_2099);
and U1146 (N_1146,In_882,In_451);
and U1147 (N_1147,In_1494,In_1390);
nand U1148 (N_1148,In_324,In_1700);
and U1149 (N_1149,In_1657,In_1903);
and U1150 (N_1150,In_2283,In_2188);
or U1151 (N_1151,In_1672,In_1930);
nand U1152 (N_1152,In_2057,In_1105);
or U1153 (N_1153,In_522,In_1717);
nand U1154 (N_1154,In_692,In_2045);
nor U1155 (N_1155,In_1823,In_199);
and U1156 (N_1156,In_828,In_217);
xor U1157 (N_1157,In_53,In_2452);
nor U1158 (N_1158,In_340,In_1100);
and U1159 (N_1159,In_2184,In_1156);
nor U1160 (N_1160,In_2349,In_1112);
nor U1161 (N_1161,In_1018,In_963);
xnor U1162 (N_1162,In_2102,In_294);
nand U1163 (N_1163,In_780,In_230);
or U1164 (N_1164,In_631,In_2297);
nand U1165 (N_1165,In_802,In_2284);
and U1166 (N_1166,In_729,In_313);
xor U1167 (N_1167,In_1806,In_1735);
and U1168 (N_1168,In_339,In_60);
nand U1169 (N_1169,In_2453,In_1036);
nand U1170 (N_1170,In_1753,In_403);
nor U1171 (N_1171,In_994,In_630);
or U1172 (N_1172,In_460,In_567);
xor U1173 (N_1173,In_2305,In_86);
xnor U1174 (N_1174,In_728,In_326);
nand U1175 (N_1175,In_2436,In_2066);
nand U1176 (N_1176,In_1932,In_1495);
nand U1177 (N_1177,In_1395,In_1707);
xor U1178 (N_1178,In_222,In_653);
or U1179 (N_1179,In_767,In_1229);
nand U1180 (N_1180,In_2268,In_2210);
or U1181 (N_1181,In_1145,In_1364);
or U1182 (N_1182,In_435,In_529);
xor U1183 (N_1183,In_2204,In_101);
xnor U1184 (N_1184,In_1627,In_967);
nor U1185 (N_1185,In_427,In_996);
and U1186 (N_1186,In_467,In_734);
nor U1187 (N_1187,In_1772,In_1462);
nor U1188 (N_1188,In_1914,In_1411);
or U1189 (N_1189,In_915,In_2438);
nand U1190 (N_1190,In_498,In_210);
xor U1191 (N_1191,In_376,In_3);
nor U1192 (N_1192,In_2116,In_1435);
nand U1193 (N_1193,In_1177,In_803);
xor U1194 (N_1194,In_1233,In_2230);
nand U1195 (N_1195,In_285,In_278);
nand U1196 (N_1196,In_491,In_2465);
or U1197 (N_1197,In_2303,In_999);
nand U1198 (N_1198,In_1486,In_731);
or U1199 (N_1199,In_19,In_2491);
and U1200 (N_1200,In_518,In_2267);
or U1201 (N_1201,In_2444,In_2251);
nor U1202 (N_1202,In_1804,In_1391);
nor U1203 (N_1203,In_2266,In_128);
nand U1204 (N_1204,In_143,In_1791);
and U1205 (N_1205,In_2097,In_725);
nand U1206 (N_1206,In_2434,In_807);
nor U1207 (N_1207,In_1680,In_1132);
xor U1208 (N_1208,In_291,In_826);
nor U1209 (N_1209,In_2423,In_1501);
nand U1210 (N_1210,In_2131,In_794);
and U1211 (N_1211,In_1693,In_851);
xnor U1212 (N_1212,In_1060,In_1040);
and U1213 (N_1213,In_2180,In_2118);
xor U1214 (N_1214,In_2234,In_981);
nor U1215 (N_1215,In_2212,In_292);
nor U1216 (N_1216,In_1189,In_1102);
nand U1217 (N_1217,In_316,In_372);
xnor U1218 (N_1218,In_2042,In_849);
or U1219 (N_1219,In_532,In_1592);
or U1220 (N_1220,In_1243,In_1682);
and U1221 (N_1221,In_769,In_1383);
nor U1222 (N_1222,In_1181,In_1175);
nand U1223 (N_1223,In_1805,In_1453);
or U1224 (N_1224,In_894,In_2243);
and U1225 (N_1225,In_1745,In_752);
nor U1226 (N_1226,In_47,In_620);
nand U1227 (N_1227,In_815,In_267);
nor U1228 (N_1228,In_266,In_2463);
xor U1229 (N_1229,In_906,In_2360);
or U1230 (N_1230,In_2386,In_1039);
xor U1231 (N_1231,In_1009,In_2275);
or U1232 (N_1232,In_2405,In_657);
xnor U1233 (N_1233,In_865,In_1651);
nor U1234 (N_1234,In_2473,In_1882);
nor U1235 (N_1235,In_1270,In_1861);
nand U1236 (N_1236,In_1663,In_343);
xnor U1237 (N_1237,In_2067,In_1744);
or U1238 (N_1238,In_1957,In_1786);
and U1239 (N_1239,In_2133,In_1221);
and U1240 (N_1240,In_629,In_2038);
xnor U1241 (N_1241,In_334,In_41);
nor U1242 (N_1242,In_477,In_468);
or U1243 (N_1243,In_1548,In_59);
nor U1244 (N_1244,In_336,In_282);
or U1245 (N_1245,In_1195,In_2223);
nor U1246 (N_1246,In_91,In_1591);
or U1247 (N_1247,In_1686,In_1265);
and U1248 (N_1248,In_2059,In_1617);
nor U1249 (N_1249,In_1216,In_1283);
and U1250 (N_1250,In_9,In_1917);
nand U1251 (N_1251,In_1444,In_953);
or U1252 (N_1252,In_611,In_992);
xor U1253 (N_1253,In_862,In_1938);
or U1254 (N_1254,In_337,In_2345);
xor U1255 (N_1255,In_709,In_2205);
xnor U1256 (N_1256,In_1628,In_1456);
and U1257 (N_1257,In_625,In_2083);
xor U1258 (N_1258,In_688,In_885);
nand U1259 (N_1259,In_911,In_1895);
nand U1260 (N_1260,In_2354,In_1161);
and U1261 (N_1261,In_1926,In_539);
nand U1262 (N_1262,In_395,In_2227);
nor U1263 (N_1263,In_247,In_2391);
xnor U1264 (N_1264,In_2119,In_265);
or U1265 (N_1265,In_215,In_2197);
xnor U1266 (N_1266,In_630,In_1055);
or U1267 (N_1267,In_675,In_808);
nor U1268 (N_1268,In_1675,In_1606);
and U1269 (N_1269,In_442,In_614);
xnor U1270 (N_1270,In_453,In_347);
xor U1271 (N_1271,In_1302,In_1949);
or U1272 (N_1272,In_2033,In_2068);
xor U1273 (N_1273,In_1647,In_1585);
nor U1274 (N_1274,In_1335,In_919);
nor U1275 (N_1275,In_2199,In_1417);
nor U1276 (N_1276,In_2450,In_281);
or U1277 (N_1277,In_1600,In_37);
xor U1278 (N_1278,In_244,In_1102);
nor U1279 (N_1279,In_1820,In_2239);
nor U1280 (N_1280,In_1290,In_506);
nand U1281 (N_1281,In_716,In_1073);
xor U1282 (N_1282,In_1534,In_2107);
xnor U1283 (N_1283,In_1403,In_1907);
or U1284 (N_1284,In_1661,In_1440);
nand U1285 (N_1285,In_351,In_1950);
nor U1286 (N_1286,In_451,In_158);
nand U1287 (N_1287,In_1544,In_1872);
and U1288 (N_1288,In_1171,In_2414);
and U1289 (N_1289,In_25,In_530);
nor U1290 (N_1290,In_1134,In_610);
or U1291 (N_1291,In_726,In_1001);
nor U1292 (N_1292,In_1229,In_1512);
nor U1293 (N_1293,In_871,In_1891);
or U1294 (N_1294,In_1672,In_1620);
or U1295 (N_1295,In_725,In_53);
or U1296 (N_1296,In_1582,In_1231);
xnor U1297 (N_1297,In_2479,In_998);
or U1298 (N_1298,In_1275,In_2414);
nor U1299 (N_1299,In_1697,In_1514);
nand U1300 (N_1300,In_1860,In_1531);
nor U1301 (N_1301,In_163,In_2465);
or U1302 (N_1302,In_2415,In_286);
nor U1303 (N_1303,In_428,In_2333);
and U1304 (N_1304,In_875,In_417);
nand U1305 (N_1305,In_286,In_1482);
nand U1306 (N_1306,In_2238,In_2007);
nand U1307 (N_1307,In_1955,In_972);
xnor U1308 (N_1308,In_481,In_1343);
nand U1309 (N_1309,In_2199,In_2180);
nor U1310 (N_1310,In_1537,In_1157);
nand U1311 (N_1311,In_948,In_343);
and U1312 (N_1312,In_71,In_1659);
and U1313 (N_1313,In_670,In_1892);
nand U1314 (N_1314,In_1004,In_626);
or U1315 (N_1315,In_1022,In_189);
and U1316 (N_1316,In_58,In_354);
or U1317 (N_1317,In_1930,In_633);
xor U1318 (N_1318,In_129,In_1);
nor U1319 (N_1319,In_792,In_2247);
xnor U1320 (N_1320,In_1839,In_1340);
nor U1321 (N_1321,In_707,In_942);
or U1322 (N_1322,In_964,In_2018);
or U1323 (N_1323,In_487,In_580);
nor U1324 (N_1324,In_412,In_503);
nand U1325 (N_1325,In_114,In_1709);
and U1326 (N_1326,In_268,In_631);
or U1327 (N_1327,In_301,In_2006);
nand U1328 (N_1328,In_2311,In_1216);
xor U1329 (N_1329,In_1409,In_2257);
xnor U1330 (N_1330,In_140,In_1252);
or U1331 (N_1331,In_2123,In_1550);
and U1332 (N_1332,In_1856,In_2229);
nor U1333 (N_1333,In_1982,In_2079);
or U1334 (N_1334,In_1136,In_1130);
nor U1335 (N_1335,In_1560,In_104);
nor U1336 (N_1336,In_22,In_2018);
nor U1337 (N_1337,In_2312,In_47);
or U1338 (N_1338,In_1093,In_1482);
xor U1339 (N_1339,In_647,In_929);
nand U1340 (N_1340,In_1307,In_331);
and U1341 (N_1341,In_1746,In_521);
and U1342 (N_1342,In_149,In_2065);
nor U1343 (N_1343,In_413,In_893);
nand U1344 (N_1344,In_1295,In_1993);
or U1345 (N_1345,In_1045,In_186);
or U1346 (N_1346,In_878,In_1592);
xnor U1347 (N_1347,In_615,In_1202);
nor U1348 (N_1348,In_259,In_1764);
xnor U1349 (N_1349,In_694,In_448);
nor U1350 (N_1350,In_1192,In_1655);
or U1351 (N_1351,In_422,In_382);
xnor U1352 (N_1352,In_1754,In_2225);
xnor U1353 (N_1353,In_845,In_529);
or U1354 (N_1354,In_2075,In_630);
and U1355 (N_1355,In_2346,In_2073);
nor U1356 (N_1356,In_1078,In_429);
nor U1357 (N_1357,In_1614,In_1826);
xnor U1358 (N_1358,In_270,In_974);
and U1359 (N_1359,In_602,In_863);
nor U1360 (N_1360,In_1990,In_2197);
nor U1361 (N_1361,In_1624,In_1392);
nand U1362 (N_1362,In_45,In_1668);
xnor U1363 (N_1363,In_1675,In_671);
or U1364 (N_1364,In_1742,In_1270);
nor U1365 (N_1365,In_1883,In_353);
and U1366 (N_1366,In_1328,In_935);
nor U1367 (N_1367,In_1558,In_106);
nor U1368 (N_1368,In_671,In_2489);
and U1369 (N_1369,In_963,In_1239);
xnor U1370 (N_1370,In_2451,In_424);
and U1371 (N_1371,In_1379,In_421);
xnor U1372 (N_1372,In_916,In_680);
xnor U1373 (N_1373,In_1551,In_1095);
nor U1374 (N_1374,In_2480,In_743);
nor U1375 (N_1375,In_1791,In_1595);
xnor U1376 (N_1376,In_2315,In_1903);
xnor U1377 (N_1377,In_940,In_1425);
nor U1378 (N_1378,In_1709,In_2281);
xor U1379 (N_1379,In_215,In_2208);
nand U1380 (N_1380,In_1844,In_2433);
nand U1381 (N_1381,In_1365,In_2079);
and U1382 (N_1382,In_947,In_1706);
xor U1383 (N_1383,In_2253,In_655);
xor U1384 (N_1384,In_423,In_1867);
nand U1385 (N_1385,In_184,In_1968);
nor U1386 (N_1386,In_56,In_283);
nand U1387 (N_1387,In_377,In_465);
or U1388 (N_1388,In_1075,In_2104);
nor U1389 (N_1389,In_2116,In_765);
xnor U1390 (N_1390,In_222,In_1733);
or U1391 (N_1391,In_774,In_2183);
nor U1392 (N_1392,In_556,In_1014);
and U1393 (N_1393,In_1742,In_2203);
and U1394 (N_1394,In_2047,In_2425);
nor U1395 (N_1395,In_1996,In_545);
nand U1396 (N_1396,In_685,In_1769);
nand U1397 (N_1397,In_1669,In_529);
or U1398 (N_1398,In_1556,In_799);
nor U1399 (N_1399,In_1142,In_1874);
nand U1400 (N_1400,In_1887,In_2300);
or U1401 (N_1401,In_4,In_1388);
xor U1402 (N_1402,In_520,In_428);
or U1403 (N_1403,In_1353,In_1720);
nand U1404 (N_1404,In_459,In_1246);
or U1405 (N_1405,In_1136,In_1863);
and U1406 (N_1406,In_2404,In_317);
nand U1407 (N_1407,In_2014,In_1842);
xnor U1408 (N_1408,In_680,In_1841);
xnor U1409 (N_1409,In_380,In_1491);
or U1410 (N_1410,In_588,In_2022);
or U1411 (N_1411,In_1150,In_765);
or U1412 (N_1412,In_1462,In_351);
xnor U1413 (N_1413,In_612,In_1147);
or U1414 (N_1414,In_883,In_1835);
xor U1415 (N_1415,In_4,In_1066);
nand U1416 (N_1416,In_1410,In_694);
and U1417 (N_1417,In_2250,In_1772);
nand U1418 (N_1418,In_595,In_2319);
nor U1419 (N_1419,In_379,In_205);
xor U1420 (N_1420,In_1624,In_1086);
nand U1421 (N_1421,In_2434,In_1077);
or U1422 (N_1422,In_181,In_1924);
xnor U1423 (N_1423,In_612,In_899);
or U1424 (N_1424,In_2014,In_1422);
nand U1425 (N_1425,In_1999,In_2333);
or U1426 (N_1426,In_1831,In_770);
nor U1427 (N_1427,In_1761,In_2011);
nand U1428 (N_1428,In_1021,In_810);
and U1429 (N_1429,In_626,In_1852);
or U1430 (N_1430,In_1857,In_685);
xor U1431 (N_1431,In_1430,In_1826);
and U1432 (N_1432,In_1913,In_1147);
xor U1433 (N_1433,In_2080,In_1597);
nand U1434 (N_1434,In_1841,In_1414);
and U1435 (N_1435,In_801,In_786);
xnor U1436 (N_1436,In_1164,In_1756);
nand U1437 (N_1437,In_843,In_2052);
nor U1438 (N_1438,In_1512,In_145);
nor U1439 (N_1439,In_2219,In_558);
xor U1440 (N_1440,In_277,In_2041);
or U1441 (N_1441,In_1194,In_445);
nor U1442 (N_1442,In_2081,In_916);
and U1443 (N_1443,In_2066,In_640);
xnor U1444 (N_1444,In_1072,In_1195);
xor U1445 (N_1445,In_1358,In_1130);
nor U1446 (N_1446,In_2087,In_315);
nor U1447 (N_1447,In_2181,In_2486);
xor U1448 (N_1448,In_1582,In_1687);
nor U1449 (N_1449,In_2059,In_1311);
and U1450 (N_1450,In_1042,In_857);
nor U1451 (N_1451,In_2037,In_281);
and U1452 (N_1452,In_2093,In_2150);
or U1453 (N_1453,In_1298,In_1808);
nor U1454 (N_1454,In_946,In_1849);
and U1455 (N_1455,In_360,In_405);
xor U1456 (N_1456,In_501,In_2319);
nor U1457 (N_1457,In_1652,In_440);
nand U1458 (N_1458,In_1979,In_792);
nand U1459 (N_1459,In_437,In_2357);
and U1460 (N_1460,In_1008,In_692);
nand U1461 (N_1461,In_1289,In_650);
or U1462 (N_1462,In_854,In_1949);
or U1463 (N_1463,In_36,In_651);
or U1464 (N_1464,In_219,In_892);
nand U1465 (N_1465,In_2341,In_1743);
nand U1466 (N_1466,In_664,In_1098);
nor U1467 (N_1467,In_2015,In_2313);
nor U1468 (N_1468,In_773,In_1654);
and U1469 (N_1469,In_53,In_1288);
and U1470 (N_1470,In_1560,In_918);
nor U1471 (N_1471,In_278,In_2282);
nand U1472 (N_1472,In_411,In_543);
or U1473 (N_1473,In_2471,In_526);
xnor U1474 (N_1474,In_2164,In_308);
nor U1475 (N_1475,In_499,In_2393);
or U1476 (N_1476,In_313,In_1095);
or U1477 (N_1477,In_1918,In_1938);
xor U1478 (N_1478,In_2489,In_2221);
and U1479 (N_1479,In_1217,In_1590);
or U1480 (N_1480,In_1738,In_765);
and U1481 (N_1481,In_334,In_885);
or U1482 (N_1482,In_279,In_463);
or U1483 (N_1483,In_2170,In_8);
or U1484 (N_1484,In_43,In_1417);
xor U1485 (N_1485,In_717,In_2109);
xor U1486 (N_1486,In_2437,In_2124);
nor U1487 (N_1487,In_2410,In_249);
and U1488 (N_1488,In_1363,In_1385);
and U1489 (N_1489,In_1155,In_2131);
and U1490 (N_1490,In_1365,In_996);
nor U1491 (N_1491,In_1939,In_1389);
nand U1492 (N_1492,In_1640,In_2202);
nand U1493 (N_1493,In_765,In_1809);
or U1494 (N_1494,In_2292,In_2199);
nor U1495 (N_1495,In_481,In_1532);
nand U1496 (N_1496,In_293,In_1414);
nand U1497 (N_1497,In_881,In_1648);
and U1498 (N_1498,In_2284,In_1647);
nand U1499 (N_1499,In_699,In_843);
or U1500 (N_1500,In_1658,In_1988);
nor U1501 (N_1501,In_883,In_1151);
and U1502 (N_1502,In_223,In_2060);
nor U1503 (N_1503,In_2269,In_369);
nor U1504 (N_1504,In_1139,In_1693);
xor U1505 (N_1505,In_1716,In_1058);
nand U1506 (N_1506,In_1967,In_904);
nand U1507 (N_1507,In_2490,In_7);
nand U1508 (N_1508,In_1685,In_184);
nand U1509 (N_1509,In_2139,In_1013);
nor U1510 (N_1510,In_264,In_2420);
nor U1511 (N_1511,In_1968,In_1860);
xor U1512 (N_1512,In_1014,In_238);
xnor U1513 (N_1513,In_1708,In_98);
nand U1514 (N_1514,In_2044,In_2050);
or U1515 (N_1515,In_1948,In_123);
xor U1516 (N_1516,In_211,In_95);
xnor U1517 (N_1517,In_1801,In_401);
xnor U1518 (N_1518,In_1229,In_2347);
and U1519 (N_1519,In_90,In_1231);
xnor U1520 (N_1520,In_1534,In_1974);
nand U1521 (N_1521,In_119,In_1231);
and U1522 (N_1522,In_1795,In_1518);
nand U1523 (N_1523,In_976,In_1009);
nand U1524 (N_1524,In_1495,In_1019);
nor U1525 (N_1525,In_673,In_2161);
and U1526 (N_1526,In_761,In_1358);
nor U1527 (N_1527,In_365,In_1662);
nand U1528 (N_1528,In_1490,In_1940);
and U1529 (N_1529,In_640,In_501);
and U1530 (N_1530,In_201,In_2212);
or U1531 (N_1531,In_2039,In_613);
and U1532 (N_1532,In_1184,In_1937);
xnor U1533 (N_1533,In_2083,In_1459);
and U1534 (N_1534,In_1029,In_1317);
nand U1535 (N_1535,In_2432,In_1110);
nor U1536 (N_1536,In_1912,In_181);
nor U1537 (N_1537,In_1159,In_1307);
or U1538 (N_1538,In_1684,In_1009);
or U1539 (N_1539,In_2244,In_2307);
xnor U1540 (N_1540,In_487,In_1634);
xnor U1541 (N_1541,In_2413,In_306);
nor U1542 (N_1542,In_391,In_1986);
nand U1543 (N_1543,In_1375,In_204);
and U1544 (N_1544,In_2248,In_572);
or U1545 (N_1545,In_1043,In_1861);
xnor U1546 (N_1546,In_774,In_2369);
xnor U1547 (N_1547,In_406,In_538);
nand U1548 (N_1548,In_451,In_1455);
xnor U1549 (N_1549,In_120,In_1213);
and U1550 (N_1550,In_532,In_379);
nand U1551 (N_1551,In_2073,In_5);
or U1552 (N_1552,In_1163,In_535);
and U1553 (N_1553,In_185,In_209);
nor U1554 (N_1554,In_626,In_180);
nor U1555 (N_1555,In_2236,In_2043);
or U1556 (N_1556,In_1202,In_1211);
xor U1557 (N_1557,In_227,In_2098);
nor U1558 (N_1558,In_1852,In_1194);
and U1559 (N_1559,In_1270,In_1466);
and U1560 (N_1560,In_1887,In_1354);
xnor U1561 (N_1561,In_363,In_1126);
and U1562 (N_1562,In_1433,In_1764);
and U1563 (N_1563,In_34,In_2302);
nand U1564 (N_1564,In_467,In_1627);
xor U1565 (N_1565,In_254,In_1875);
and U1566 (N_1566,In_570,In_533);
or U1567 (N_1567,In_1568,In_2023);
nand U1568 (N_1568,In_2240,In_372);
or U1569 (N_1569,In_1459,In_2191);
nand U1570 (N_1570,In_585,In_1760);
nand U1571 (N_1571,In_572,In_208);
and U1572 (N_1572,In_865,In_2400);
and U1573 (N_1573,In_278,In_1173);
xor U1574 (N_1574,In_630,In_2387);
and U1575 (N_1575,In_1621,In_901);
nor U1576 (N_1576,In_2453,In_1348);
and U1577 (N_1577,In_1528,In_2105);
or U1578 (N_1578,In_1387,In_1323);
and U1579 (N_1579,In_2195,In_719);
and U1580 (N_1580,In_865,In_1583);
and U1581 (N_1581,In_2282,In_68);
nor U1582 (N_1582,In_1630,In_1767);
nand U1583 (N_1583,In_1991,In_2319);
and U1584 (N_1584,In_442,In_1614);
xnor U1585 (N_1585,In_984,In_62);
or U1586 (N_1586,In_2459,In_1246);
nor U1587 (N_1587,In_2275,In_1779);
xor U1588 (N_1588,In_1575,In_825);
nor U1589 (N_1589,In_1235,In_1031);
xnor U1590 (N_1590,In_598,In_942);
or U1591 (N_1591,In_2017,In_166);
or U1592 (N_1592,In_613,In_229);
nor U1593 (N_1593,In_284,In_1710);
nor U1594 (N_1594,In_1538,In_1345);
and U1595 (N_1595,In_2209,In_1336);
and U1596 (N_1596,In_1499,In_187);
or U1597 (N_1597,In_117,In_1788);
nand U1598 (N_1598,In_227,In_1429);
nor U1599 (N_1599,In_1371,In_1167);
nor U1600 (N_1600,In_2241,In_1302);
nand U1601 (N_1601,In_2205,In_1757);
nand U1602 (N_1602,In_1512,In_502);
nand U1603 (N_1603,In_1051,In_665);
nor U1604 (N_1604,In_2420,In_1506);
nand U1605 (N_1605,In_840,In_297);
nor U1606 (N_1606,In_1134,In_1379);
nor U1607 (N_1607,In_613,In_2361);
or U1608 (N_1608,In_7,In_609);
or U1609 (N_1609,In_178,In_79);
and U1610 (N_1610,In_1272,In_487);
or U1611 (N_1611,In_1373,In_915);
nor U1612 (N_1612,In_542,In_652);
or U1613 (N_1613,In_2371,In_1995);
or U1614 (N_1614,In_2308,In_507);
xor U1615 (N_1615,In_629,In_2372);
and U1616 (N_1616,In_2340,In_2375);
nand U1617 (N_1617,In_1035,In_1773);
or U1618 (N_1618,In_458,In_783);
nor U1619 (N_1619,In_476,In_837);
and U1620 (N_1620,In_596,In_1965);
xor U1621 (N_1621,In_295,In_1545);
and U1622 (N_1622,In_272,In_2388);
or U1623 (N_1623,In_434,In_1265);
or U1624 (N_1624,In_1029,In_1305);
and U1625 (N_1625,In_323,In_631);
nor U1626 (N_1626,In_1485,In_1649);
or U1627 (N_1627,In_539,In_1060);
or U1628 (N_1628,In_1478,In_271);
and U1629 (N_1629,In_1105,In_1383);
nor U1630 (N_1630,In_482,In_327);
and U1631 (N_1631,In_565,In_1127);
or U1632 (N_1632,In_1351,In_1151);
and U1633 (N_1633,In_315,In_1411);
nand U1634 (N_1634,In_2379,In_604);
xor U1635 (N_1635,In_825,In_1515);
nand U1636 (N_1636,In_823,In_1116);
xor U1637 (N_1637,In_430,In_1371);
nand U1638 (N_1638,In_1979,In_87);
or U1639 (N_1639,In_234,In_890);
nor U1640 (N_1640,In_605,In_1070);
nand U1641 (N_1641,In_2151,In_1726);
nand U1642 (N_1642,In_872,In_1265);
nand U1643 (N_1643,In_2121,In_1477);
or U1644 (N_1644,In_1217,In_413);
or U1645 (N_1645,In_1923,In_336);
and U1646 (N_1646,In_899,In_1163);
nand U1647 (N_1647,In_240,In_1749);
or U1648 (N_1648,In_1075,In_929);
nand U1649 (N_1649,In_262,In_1699);
and U1650 (N_1650,In_749,In_532);
xnor U1651 (N_1651,In_1996,In_1746);
and U1652 (N_1652,In_516,In_1357);
nor U1653 (N_1653,In_1993,In_1691);
nand U1654 (N_1654,In_1698,In_2044);
nand U1655 (N_1655,In_266,In_2145);
or U1656 (N_1656,In_1844,In_805);
or U1657 (N_1657,In_2401,In_1473);
nor U1658 (N_1658,In_1754,In_1769);
xnor U1659 (N_1659,In_1357,In_1283);
nor U1660 (N_1660,In_887,In_1427);
or U1661 (N_1661,In_2051,In_730);
nor U1662 (N_1662,In_2383,In_651);
nand U1663 (N_1663,In_1318,In_2447);
and U1664 (N_1664,In_1501,In_167);
nor U1665 (N_1665,In_1531,In_818);
nand U1666 (N_1666,In_901,In_800);
or U1667 (N_1667,In_185,In_1370);
xnor U1668 (N_1668,In_2084,In_1726);
nand U1669 (N_1669,In_2111,In_1975);
nand U1670 (N_1670,In_1887,In_1611);
or U1671 (N_1671,In_343,In_962);
and U1672 (N_1672,In_2109,In_305);
or U1673 (N_1673,In_1206,In_1856);
nand U1674 (N_1674,In_2269,In_954);
nand U1675 (N_1675,In_2129,In_2004);
and U1676 (N_1676,In_1927,In_562);
nand U1677 (N_1677,In_2337,In_1962);
or U1678 (N_1678,In_2189,In_2415);
nand U1679 (N_1679,In_2027,In_135);
xnor U1680 (N_1680,In_1826,In_1823);
nand U1681 (N_1681,In_1816,In_1040);
and U1682 (N_1682,In_2249,In_219);
and U1683 (N_1683,In_147,In_1818);
and U1684 (N_1684,In_433,In_1498);
nand U1685 (N_1685,In_1685,In_417);
xor U1686 (N_1686,In_696,In_1800);
and U1687 (N_1687,In_1462,In_937);
nand U1688 (N_1688,In_70,In_1464);
or U1689 (N_1689,In_988,In_454);
nand U1690 (N_1690,In_527,In_810);
nor U1691 (N_1691,In_774,In_1815);
nor U1692 (N_1692,In_782,In_1414);
xor U1693 (N_1693,In_2309,In_2094);
or U1694 (N_1694,In_1210,In_1121);
and U1695 (N_1695,In_367,In_1665);
and U1696 (N_1696,In_2070,In_581);
and U1697 (N_1697,In_445,In_2233);
or U1698 (N_1698,In_1725,In_291);
xor U1699 (N_1699,In_163,In_953);
and U1700 (N_1700,In_1069,In_1065);
or U1701 (N_1701,In_1390,In_645);
or U1702 (N_1702,In_947,In_1160);
and U1703 (N_1703,In_1828,In_734);
and U1704 (N_1704,In_1945,In_2100);
nand U1705 (N_1705,In_819,In_471);
and U1706 (N_1706,In_322,In_901);
and U1707 (N_1707,In_1741,In_1207);
or U1708 (N_1708,In_9,In_717);
or U1709 (N_1709,In_166,In_745);
nor U1710 (N_1710,In_74,In_1138);
xor U1711 (N_1711,In_90,In_1690);
xor U1712 (N_1712,In_1077,In_2055);
and U1713 (N_1713,In_67,In_1486);
or U1714 (N_1714,In_2120,In_690);
xor U1715 (N_1715,In_2273,In_2375);
nand U1716 (N_1716,In_1580,In_1515);
and U1717 (N_1717,In_2007,In_1051);
nand U1718 (N_1718,In_1383,In_1682);
nor U1719 (N_1719,In_1006,In_1308);
or U1720 (N_1720,In_2473,In_1947);
or U1721 (N_1721,In_1774,In_1986);
and U1722 (N_1722,In_1769,In_991);
xor U1723 (N_1723,In_1047,In_1948);
xnor U1724 (N_1724,In_801,In_1812);
and U1725 (N_1725,In_2234,In_1164);
and U1726 (N_1726,In_2335,In_2052);
nand U1727 (N_1727,In_1738,In_1709);
nand U1728 (N_1728,In_1885,In_1231);
nand U1729 (N_1729,In_2477,In_0);
and U1730 (N_1730,In_947,In_1036);
or U1731 (N_1731,In_1694,In_104);
xnor U1732 (N_1732,In_1502,In_2211);
xnor U1733 (N_1733,In_289,In_126);
nand U1734 (N_1734,In_1679,In_1845);
nor U1735 (N_1735,In_2140,In_1699);
nor U1736 (N_1736,In_2447,In_1912);
and U1737 (N_1737,In_155,In_379);
and U1738 (N_1738,In_613,In_1243);
or U1739 (N_1739,In_1187,In_2253);
nor U1740 (N_1740,In_834,In_2229);
and U1741 (N_1741,In_281,In_287);
or U1742 (N_1742,In_95,In_1211);
or U1743 (N_1743,In_360,In_1646);
nor U1744 (N_1744,In_2394,In_2344);
and U1745 (N_1745,In_513,In_1776);
nor U1746 (N_1746,In_369,In_2234);
nand U1747 (N_1747,In_1806,In_487);
or U1748 (N_1748,In_1240,In_2358);
nand U1749 (N_1749,In_981,In_449);
and U1750 (N_1750,In_1469,In_1859);
nand U1751 (N_1751,In_886,In_2270);
and U1752 (N_1752,In_2048,In_721);
nor U1753 (N_1753,In_1365,In_733);
nor U1754 (N_1754,In_282,In_521);
or U1755 (N_1755,In_974,In_1200);
nand U1756 (N_1756,In_1766,In_468);
nor U1757 (N_1757,In_1993,In_2146);
nand U1758 (N_1758,In_772,In_691);
xor U1759 (N_1759,In_1772,In_812);
and U1760 (N_1760,In_92,In_696);
or U1761 (N_1761,In_1241,In_759);
xor U1762 (N_1762,In_1379,In_2452);
xor U1763 (N_1763,In_2139,In_1895);
nand U1764 (N_1764,In_1930,In_58);
xor U1765 (N_1765,In_662,In_1628);
nand U1766 (N_1766,In_1694,In_1440);
or U1767 (N_1767,In_1973,In_783);
and U1768 (N_1768,In_598,In_1211);
xnor U1769 (N_1769,In_2497,In_2377);
nor U1770 (N_1770,In_1292,In_338);
nand U1771 (N_1771,In_2162,In_896);
and U1772 (N_1772,In_1282,In_540);
or U1773 (N_1773,In_1821,In_802);
nor U1774 (N_1774,In_1381,In_1001);
or U1775 (N_1775,In_1941,In_2413);
nand U1776 (N_1776,In_901,In_1883);
nand U1777 (N_1777,In_2495,In_347);
nor U1778 (N_1778,In_177,In_2033);
or U1779 (N_1779,In_628,In_1365);
nand U1780 (N_1780,In_1476,In_2023);
xnor U1781 (N_1781,In_2480,In_1047);
or U1782 (N_1782,In_1868,In_1323);
and U1783 (N_1783,In_566,In_358);
or U1784 (N_1784,In_2297,In_314);
nand U1785 (N_1785,In_443,In_1895);
nand U1786 (N_1786,In_2481,In_929);
nand U1787 (N_1787,In_2091,In_135);
and U1788 (N_1788,In_2331,In_1186);
and U1789 (N_1789,In_2240,In_1011);
and U1790 (N_1790,In_1329,In_469);
and U1791 (N_1791,In_1915,In_967);
and U1792 (N_1792,In_274,In_581);
xnor U1793 (N_1793,In_2449,In_1918);
and U1794 (N_1794,In_1112,In_1784);
or U1795 (N_1795,In_851,In_2012);
nand U1796 (N_1796,In_1847,In_2250);
and U1797 (N_1797,In_135,In_1569);
or U1798 (N_1798,In_1004,In_2090);
nand U1799 (N_1799,In_862,In_284);
or U1800 (N_1800,In_550,In_761);
and U1801 (N_1801,In_2471,In_1423);
nand U1802 (N_1802,In_1927,In_1221);
nor U1803 (N_1803,In_2063,In_912);
and U1804 (N_1804,In_1473,In_2121);
nor U1805 (N_1805,In_2263,In_2353);
and U1806 (N_1806,In_1788,In_576);
xor U1807 (N_1807,In_2334,In_158);
nor U1808 (N_1808,In_88,In_1872);
nand U1809 (N_1809,In_448,In_1979);
or U1810 (N_1810,In_290,In_1683);
and U1811 (N_1811,In_1852,In_12);
xnor U1812 (N_1812,In_1809,In_2297);
nand U1813 (N_1813,In_642,In_1909);
nand U1814 (N_1814,In_2257,In_2258);
nor U1815 (N_1815,In_2220,In_1224);
nor U1816 (N_1816,In_456,In_2156);
nor U1817 (N_1817,In_1658,In_260);
xor U1818 (N_1818,In_1926,In_1991);
xor U1819 (N_1819,In_1784,In_1257);
xor U1820 (N_1820,In_641,In_472);
nand U1821 (N_1821,In_36,In_1467);
and U1822 (N_1822,In_1754,In_328);
nor U1823 (N_1823,In_359,In_1273);
xnor U1824 (N_1824,In_1545,In_307);
nor U1825 (N_1825,In_1067,In_2140);
or U1826 (N_1826,In_1554,In_1074);
nor U1827 (N_1827,In_331,In_1972);
and U1828 (N_1828,In_2381,In_877);
or U1829 (N_1829,In_269,In_1286);
xnor U1830 (N_1830,In_464,In_1638);
xnor U1831 (N_1831,In_194,In_2377);
or U1832 (N_1832,In_1986,In_2482);
and U1833 (N_1833,In_1410,In_866);
xor U1834 (N_1834,In_2002,In_155);
xor U1835 (N_1835,In_1598,In_841);
and U1836 (N_1836,In_325,In_1721);
and U1837 (N_1837,In_365,In_1804);
and U1838 (N_1838,In_470,In_501);
nand U1839 (N_1839,In_2055,In_1447);
xnor U1840 (N_1840,In_1647,In_1494);
and U1841 (N_1841,In_1194,In_1279);
or U1842 (N_1842,In_71,In_1125);
and U1843 (N_1843,In_1005,In_601);
xor U1844 (N_1844,In_2150,In_2066);
nand U1845 (N_1845,In_158,In_1818);
or U1846 (N_1846,In_2350,In_676);
or U1847 (N_1847,In_1799,In_1902);
nor U1848 (N_1848,In_184,In_1919);
and U1849 (N_1849,In_2061,In_2117);
or U1850 (N_1850,In_435,In_855);
and U1851 (N_1851,In_345,In_912);
nor U1852 (N_1852,In_578,In_551);
and U1853 (N_1853,In_656,In_285);
nand U1854 (N_1854,In_276,In_2223);
nand U1855 (N_1855,In_1154,In_1688);
or U1856 (N_1856,In_2047,In_2162);
nor U1857 (N_1857,In_782,In_1780);
or U1858 (N_1858,In_1352,In_1769);
xnor U1859 (N_1859,In_1966,In_1498);
and U1860 (N_1860,In_2296,In_1879);
and U1861 (N_1861,In_320,In_2315);
xor U1862 (N_1862,In_2079,In_41);
nand U1863 (N_1863,In_1891,In_1019);
and U1864 (N_1864,In_823,In_2063);
or U1865 (N_1865,In_313,In_1235);
nor U1866 (N_1866,In_1002,In_1062);
nor U1867 (N_1867,In_1958,In_767);
nand U1868 (N_1868,In_2215,In_676);
nor U1869 (N_1869,In_1665,In_1892);
and U1870 (N_1870,In_1800,In_738);
nor U1871 (N_1871,In_1158,In_1208);
nor U1872 (N_1872,In_1327,In_776);
nand U1873 (N_1873,In_2255,In_1659);
or U1874 (N_1874,In_791,In_1411);
xnor U1875 (N_1875,In_288,In_228);
nand U1876 (N_1876,In_2046,In_1443);
and U1877 (N_1877,In_2408,In_649);
nand U1878 (N_1878,In_416,In_2471);
xnor U1879 (N_1879,In_204,In_1865);
and U1880 (N_1880,In_2044,In_712);
nor U1881 (N_1881,In_237,In_946);
nand U1882 (N_1882,In_24,In_42);
and U1883 (N_1883,In_1858,In_2424);
or U1884 (N_1884,In_157,In_1371);
and U1885 (N_1885,In_121,In_1677);
and U1886 (N_1886,In_2453,In_1815);
nor U1887 (N_1887,In_2097,In_1205);
or U1888 (N_1888,In_1731,In_1469);
nand U1889 (N_1889,In_2171,In_804);
nand U1890 (N_1890,In_1282,In_360);
and U1891 (N_1891,In_1446,In_2041);
and U1892 (N_1892,In_676,In_1860);
or U1893 (N_1893,In_406,In_746);
and U1894 (N_1894,In_1038,In_1818);
and U1895 (N_1895,In_84,In_2494);
xnor U1896 (N_1896,In_149,In_1379);
xor U1897 (N_1897,In_1550,In_1709);
and U1898 (N_1898,In_748,In_1228);
nand U1899 (N_1899,In_211,In_1399);
nand U1900 (N_1900,In_133,In_1290);
nand U1901 (N_1901,In_1592,In_2239);
or U1902 (N_1902,In_372,In_1787);
nand U1903 (N_1903,In_298,In_705);
nor U1904 (N_1904,In_2474,In_1500);
nand U1905 (N_1905,In_1813,In_1523);
xor U1906 (N_1906,In_592,In_769);
xnor U1907 (N_1907,In_2292,In_622);
or U1908 (N_1908,In_1190,In_2370);
or U1909 (N_1909,In_2320,In_668);
nor U1910 (N_1910,In_1118,In_1316);
and U1911 (N_1911,In_2441,In_1206);
and U1912 (N_1912,In_299,In_2151);
or U1913 (N_1913,In_2404,In_971);
nand U1914 (N_1914,In_2490,In_871);
or U1915 (N_1915,In_1356,In_1531);
nand U1916 (N_1916,In_1452,In_2277);
nand U1917 (N_1917,In_192,In_1967);
or U1918 (N_1918,In_980,In_1777);
and U1919 (N_1919,In_1518,In_1529);
xor U1920 (N_1920,In_1675,In_906);
xnor U1921 (N_1921,In_1732,In_1180);
nand U1922 (N_1922,In_1456,In_441);
nand U1923 (N_1923,In_556,In_1167);
nand U1924 (N_1924,In_1034,In_635);
or U1925 (N_1925,In_1392,In_1528);
nor U1926 (N_1926,In_653,In_328);
nor U1927 (N_1927,In_2285,In_699);
or U1928 (N_1928,In_2382,In_1684);
nand U1929 (N_1929,In_574,In_1810);
and U1930 (N_1930,In_1670,In_2392);
xor U1931 (N_1931,In_921,In_2001);
nand U1932 (N_1932,In_674,In_2179);
xnor U1933 (N_1933,In_1752,In_1924);
and U1934 (N_1934,In_2168,In_2072);
nand U1935 (N_1935,In_1626,In_1532);
nor U1936 (N_1936,In_879,In_41);
nor U1937 (N_1937,In_2280,In_742);
nand U1938 (N_1938,In_673,In_2286);
nor U1939 (N_1939,In_2135,In_2106);
nand U1940 (N_1940,In_534,In_859);
nor U1941 (N_1941,In_439,In_981);
xnor U1942 (N_1942,In_309,In_1230);
xnor U1943 (N_1943,In_384,In_2456);
nor U1944 (N_1944,In_1513,In_1529);
or U1945 (N_1945,In_2110,In_56);
or U1946 (N_1946,In_1340,In_255);
and U1947 (N_1947,In_90,In_2316);
nor U1948 (N_1948,In_1055,In_1039);
nand U1949 (N_1949,In_1708,In_500);
xnor U1950 (N_1950,In_674,In_205);
and U1951 (N_1951,In_2212,In_2077);
xnor U1952 (N_1952,In_830,In_992);
xnor U1953 (N_1953,In_1180,In_1309);
and U1954 (N_1954,In_1882,In_2116);
xnor U1955 (N_1955,In_111,In_1147);
nand U1956 (N_1956,In_1942,In_342);
nor U1957 (N_1957,In_1560,In_2221);
nand U1958 (N_1958,In_635,In_971);
nand U1959 (N_1959,In_454,In_2133);
and U1960 (N_1960,In_267,In_2153);
nor U1961 (N_1961,In_1881,In_189);
nand U1962 (N_1962,In_1346,In_1497);
nor U1963 (N_1963,In_2407,In_1777);
nand U1964 (N_1964,In_1352,In_645);
xor U1965 (N_1965,In_251,In_2236);
or U1966 (N_1966,In_202,In_2380);
nand U1967 (N_1967,In_174,In_1569);
or U1968 (N_1968,In_567,In_261);
xnor U1969 (N_1969,In_234,In_262);
or U1970 (N_1970,In_1345,In_1340);
xnor U1971 (N_1971,In_1592,In_1069);
nand U1972 (N_1972,In_214,In_410);
or U1973 (N_1973,In_883,In_1606);
or U1974 (N_1974,In_1528,In_21);
or U1975 (N_1975,In_2260,In_1112);
xnor U1976 (N_1976,In_396,In_758);
or U1977 (N_1977,In_1926,In_1361);
and U1978 (N_1978,In_13,In_787);
or U1979 (N_1979,In_359,In_819);
nand U1980 (N_1980,In_1609,In_642);
nor U1981 (N_1981,In_1280,In_1462);
and U1982 (N_1982,In_1678,In_258);
and U1983 (N_1983,In_452,In_112);
and U1984 (N_1984,In_1346,In_63);
nand U1985 (N_1985,In_1880,In_2398);
and U1986 (N_1986,In_218,In_40);
and U1987 (N_1987,In_1305,In_811);
xor U1988 (N_1988,In_619,In_914);
nand U1989 (N_1989,In_1677,In_54);
nor U1990 (N_1990,In_250,In_510);
and U1991 (N_1991,In_919,In_452);
or U1992 (N_1992,In_568,In_2430);
nand U1993 (N_1993,In_296,In_690);
nor U1994 (N_1994,In_1515,In_637);
xnor U1995 (N_1995,In_1455,In_1906);
or U1996 (N_1996,In_1817,In_1448);
and U1997 (N_1997,In_883,In_2127);
and U1998 (N_1998,In_775,In_2146);
and U1999 (N_1999,In_988,In_1731);
nor U2000 (N_2000,In_1781,In_1393);
and U2001 (N_2001,In_599,In_784);
xor U2002 (N_2002,In_1718,In_2078);
and U2003 (N_2003,In_1623,In_1102);
xor U2004 (N_2004,In_901,In_2209);
and U2005 (N_2005,In_923,In_1083);
and U2006 (N_2006,In_1586,In_2245);
and U2007 (N_2007,In_1636,In_2292);
and U2008 (N_2008,In_281,In_177);
xor U2009 (N_2009,In_269,In_2194);
and U2010 (N_2010,In_1760,In_1594);
or U2011 (N_2011,In_825,In_151);
xor U2012 (N_2012,In_479,In_325);
and U2013 (N_2013,In_1384,In_1698);
and U2014 (N_2014,In_1428,In_2042);
or U2015 (N_2015,In_2235,In_741);
and U2016 (N_2016,In_913,In_5);
nor U2017 (N_2017,In_2494,In_1599);
nand U2018 (N_2018,In_1248,In_2128);
and U2019 (N_2019,In_1121,In_1814);
and U2020 (N_2020,In_2484,In_846);
xor U2021 (N_2021,In_1934,In_527);
and U2022 (N_2022,In_500,In_97);
nand U2023 (N_2023,In_672,In_335);
nand U2024 (N_2024,In_1703,In_2308);
nand U2025 (N_2025,In_454,In_1669);
or U2026 (N_2026,In_149,In_2312);
nor U2027 (N_2027,In_1402,In_87);
or U2028 (N_2028,In_899,In_1214);
nor U2029 (N_2029,In_1521,In_1558);
nand U2030 (N_2030,In_1896,In_2194);
nor U2031 (N_2031,In_1441,In_1968);
xor U2032 (N_2032,In_2432,In_42);
nor U2033 (N_2033,In_225,In_1586);
nor U2034 (N_2034,In_1694,In_1864);
nor U2035 (N_2035,In_1612,In_92);
or U2036 (N_2036,In_322,In_713);
xor U2037 (N_2037,In_47,In_25);
nand U2038 (N_2038,In_2467,In_693);
or U2039 (N_2039,In_850,In_738);
nor U2040 (N_2040,In_803,In_154);
or U2041 (N_2041,In_220,In_1987);
or U2042 (N_2042,In_1976,In_1578);
xor U2043 (N_2043,In_148,In_2443);
or U2044 (N_2044,In_1497,In_596);
and U2045 (N_2045,In_741,In_1005);
nand U2046 (N_2046,In_206,In_1477);
and U2047 (N_2047,In_397,In_410);
nor U2048 (N_2048,In_66,In_1685);
xnor U2049 (N_2049,In_1218,In_1202);
or U2050 (N_2050,In_1252,In_529);
nand U2051 (N_2051,In_1220,In_51);
nand U2052 (N_2052,In_1767,In_800);
nand U2053 (N_2053,In_2386,In_1898);
nor U2054 (N_2054,In_1106,In_1303);
nor U2055 (N_2055,In_1321,In_219);
xnor U2056 (N_2056,In_414,In_1723);
nor U2057 (N_2057,In_1661,In_2429);
nor U2058 (N_2058,In_262,In_1725);
xnor U2059 (N_2059,In_930,In_2392);
or U2060 (N_2060,In_88,In_1903);
or U2061 (N_2061,In_2120,In_782);
or U2062 (N_2062,In_605,In_2100);
xnor U2063 (N_2063,In_1282,In_2216);
nand U2064 (N_2064,In_1713,In_46);
xnor U2065 (N_2065,In_307,In_1061);
xnor U2066 (N_2066,In_545,In_1191);
nor U2067 (N_2067,In_568,In_277);
and U2068 (N_2068,In_1088,In_1545);
or U2069 (N_2069,In_1979,In_408);
and U2070 (N_2070,In_2012,In_658);
xnor U2071 (N_2071,In_1058,In_550);
xor U2072 (N_2072,In_376,In_661);
nand U2073 (N_2073,In_93,In_828);
xnor U2074 (N_2074,In_1453,In_883);
xnor U2075 (N_2075,In_1650,In_1267);
or U2076 (N_2076,In_1828,In_2048);
nand U2077 (N_2077,In_539,In_2095);
and U2078 (N_2078,In_1396,In_137);
or U2079 (N_2079,In_834,In_1243);
xor U2080 (N_2080,In_1307,In_1900);
xor U2081 (N_2081,In_1541,In_2417);
xor U2082 (N_2082,In_526,In_111);
nand U2083 (N_2083,In_2387,In_1712);
and U2084 (N_2084,In_755,In_2122);
and U2085 (N_2085,In_274,In_1368);
xnor U2086 (N_2086,In_2306,In_782);
xnor U2087 (N_2087,In_2255,In_1909);
xnor U2088 (N_2088,In_77,In_1381);
nor U2089 (N_2089,In_2115,In_1499);
xor U2090 (N_2090,In_460,In_649);
xnor U2091 (N_2091,In_1091,In_1679);
and U2092 (N_2092,In_1905,In_1260);
or U2093 (N_2093,In_1321,In_838);
xnor U2094 (N_2094,In_1853,In_1155);
nor U2095 (N_2095,In_662,In_2101);
or U2096 (N_2096,In_1050,In_1450);
or U2097 (N_2097,In_1716,In_397);
nand U2098 (N_2098,In_1407,In_1549);
nor U2099 (N_2099,In_1759,In_1826);
nor U2100 (N_2100,In_2126,In_2450);
or U2101 (N_2101,In_1946,In_891);
xor U2102 (N_2102,In_1545,In_2175);
or U2103 (N_2103,In_2040,In_1285);
or U2104 (N_2104,In_324,In_1672);
nand U2105 (N_2105,In_74,In_2486);
nand U2106 (N_2106,In_715,In_1457);
or U2107 (N_2107,In_387,In_1434);
nor U2108 (N_2108,In_1122,In_229);
and U2109 (N_2109,In_1629,In_2494);
nand U2110 (N_2110,In_930,In_854);
and U2111 (N_2111,In_976,In_2288);
and U2112 (N_2112,In_1736,In_2308);
nor U2113 (N_2113,In_242,In_1685);
and U2114 (N_2114,In_900,In_1785);
nand U2115 (N_2115,In_222,In_1200);
xnor U2116 (N_2116,In_87,In_2343);
nor U2117 (N_2117,In_1908,In_1299);
nand U2118 (N_2118,In_574,In_1232);
nand U2119 (N_2119,In_2485,In_818);
or U2120 (N_2120,In_2305,In_1156);
or U2121 (N_2121,In_569,In_971);
nand U2122 (N_2122,In_2066,In_947);
nand U2123 (N_2123,In_1537,In_2057);
nor U2124 (N_2124,In_837,In_702);
and U2125 (N_2125,In_1389,In_1364);
xnor U2126 (N_2126,In_1715,In_866);
and U2127 (N_2127,In_370,In_1143);
nand U2128 (N_2128,In_2170,In_19);
or U2129 (N_2129,In_235,In_319);
nand U2130 (N_2130,In_1527,In_1189);
nand U2131 (N_2131,In_1278,In_1985);
or U2132 (N_2132,In_897,In_2243);
nor U2133 (N_2133,In_962,In_1492);
nor U2134 (N_2134,In_381,In_1628);
nand U2135 (N_2135,In_1845,In_2476);
nor U2136 (N_2136,In_851,In_153);
and U2137 (N_2137,In_2235,In_789);
nor U2138 (N_2138,In_2483,In_1621);
nand U2139 (N_2139,In_626,In_1393);
and U2140 (N_2140,In_144,In_1743);
or U2141 (N_2141,In_1149,In_911);
or U2142 (N_2142,In_1036,In_286);
nand U2143 (N_2143,In_313,In_2133);
nand U2144 (N_2144,In_671,In_662);
nor U2145 (N_2145,In_2476,In_1710);
nor U2146 (N_2146,In_90,In_2472);
or U2147 (N_2147,In_1052,In_1179);
nand U2148 (N_2148,In_1713,In_2239);
xor U2149 (N_2149,In_2375,In_1838);
xnor U2150 (N_2150,In_857,In_1363);
or U2151 (N_2151,In_1360,In_1370);
nor U2152 (N_2152,In_1314,In_893);
nand U2153 (N_2153,In_2253,In_1118);
or U2154 (N_2154,In_2141,In_488);
or U2155 (N_2155,In_1406,In_7);
xor U2156 (N_2156,In_1460,In_2337);
or U2157 (N_2157,In_1994,In_1179);
and U2158 (N_2158,In_727,In_374);
nand U2159 (N_2159,In_765,In_835);
or U2160 (N_2160,In_1803,In_767);
xnor U2161 (N_2161,In_547,In_429);
nand U2162 (N_2162,In_2152,In_134);
or U2163 (N_2163,In_609,In_1763);
or U2164 (N_2164,In_355,In_1296);
and U2165 (N_2165,In_860,In_1907);
and U2166 (N_2166,In_307,In_464);
xnor U2167 (N_2167,In_2156,In_644);
xor U2168 (N_2168,In_113,In_1547);
or U2169 (N_2169,In_1033,In_92);
nor U2170 (N_2170,In_446,In_1426);
or U2171 (N_2171,In_244,In_1602);
nor U2172 (N_2172,In_217,In_1048);
or U2173 (N_2173,In_352,In_2408);
nor U2174 (N_2174,In_1358,In_2259);
or U2175 (N_2175,In_1426,In_774);
and U2176 (N_2176,In_190,In_1101);
nand U2177 (N_2177,In_2484,In_866);
and U2178 (N_2178,In_2296,In_1042);
nand U2179 (N_2179,In_2309,In_636);
and U2180 (N_2180,In_21,In_1294);
xnor U2181 (N_2181,In_2305,In_2431);
xnor U2182 (N_2182,In_907,In_2214);
nor U2183 (N_2183,In_556,In_2271);
nor U2184 (N_2184,In_1843,In_1593);
or U2185 (N_2185,In_1999,In_610);
or U2186 (N_2186,In_399,In_518);
xor U2187 (N_2187,In_1932,In_692);
or U2188 (N_2188,In_1864,In_1042);
and U2189 (N_2189,In_1341,In_1018);
xor U2190 (N_2190,In_2440,In_590);
nor U2191 (N_2191,In_1997,In_1377);
nor U2192 (N_2192,In_376,In_365);
nand U2193 (N_2193,In_2039,In_958);
or U2194 (N_2194,In_1399,In_1836);
and U2195 (N_2195,In_1939,In_617);
xnor U2196 (N_2196,In_688,In_1189);
and U2197 (N_2197,In_1741,In_155);
and U2198 (N_2198,In_1402,In_1126);
xor U2199 (N_2199,In_304,In_555);
or U2200 (N_2200,In_381,In_1445);
xnor U2201 (N_2201,In_1869,In_1069);
nand U2202 (N_2202,In_595,In_1107);
nor U2203 (N_2203,In_520,In_1244);
xnor U2204 (N_2204,In_1825,In_531);
nor U2205 (N_2205,In_1995,In_1957);
xnor U2206 (N_2206,In_1077,In_529);
nor U2207 (N_2207,In_170,In_1663);
nand U2208 (N_2208,In_268,In_161);
or U2209 (N_2209,In_1216,In_42);
and U2210 (N_2210,In_696,In_174);
xor U2211 (N_2211,In_72,In_1231);
and U2212 (N_2212,In_1230,In_1797);
xor U2213 (N_2213,In_477,In_396);
or U2214 (N_2214,In_239,In_2144);
and U2215 (N_2215,In_1500,In_213);
nor U2216 (N_2216,In_61,In_2392);
or U2217 (N_2217,In_1867,In_668);
and U2218 (N_2218,In_1228,In_2446);
or U2219 (N_2219,In_2109,In_329);
and U2220 (N_2220,In_155,In_2325);
nand U2221 (N_2221,In_2369,In_2170);
xor U2222 (N_2222,In_2017,In_916);
nor U2223 (N_2223,In_1708,In_1509);
and U2224 (N_2224,In_1759,In_117);
nand U2225 (N_2225,In_1893,In_1784);
nand U2226 (N_2226,In_1433,In_882);
nand U2227 (N_2227,In_379,In_566);
or U2228 (N_2228,In_1987,In_1930);
or U2229 (N_2229,In_87,In_629);
and U2230 (N_2230,In_926,In_2459);
nand U2231 (N_2231,In_1742,In_2354);
or U2232 (N_2232,In_1203,In_1477);
nor U2233 (N_2233,In_260,In_975);
and U2234 (N_2234,In_1952,In_2236);
and U2235 (N_2235,In_1493,In_2174);
xnor U2236 (N_2236,In_412,In_194);
nor U2237 (N_2237,In_2413,In_2195);
nor U2238 (N_2238,In_1554,In_209);
nor U2239 (N_2239,In_2111,In_2081);
nand U2240 (N_2240,In_1289,In_361);
and U2241 (N_2241,In_1818,In_1911);
or U2242 (N_2242,In_2149,In_2042);
xor U2243 (N_2243,In_1345,In_838);
xor U2244 (N_2244,In_1975,In_1198);
or U2245 (N_2245,In_106,In_1901);
nor U2246 (N_2246,In_674,In_63);
and U2247 (N_2247,In_2250,In_1693);
and U2248 (N_2248,In_1330,In_1314);
or U2249 (N_2249,In_1559,In_335);
and U2250 (N_2250,In_294,In_2352);
or U2251 (N_2251,In_2314,In_764);
nor U2252 (N_2252,In_1928,In_2236);
xnor U2253 (N_2253,In_1453,In_870);
nand U2254 (N_2254,In_807,In_528);
nor U2255 (N_2255,In_1748,In_1455);
or U2256 (N_2256,In_397,In_1844);
nor U2257 (N_2257,In_173,In_1206);
xnor U2258 (N_2258,In_1657,In_2118);
and U2259 (N_2259,In_226,In_1115);
and U2260 (N_2260,In_943,In_636);
and U2261 (N_2261,In_501,In_2065);
and U2262 (N_2262,In_1092,In_517);
nand U2263 (N_2263,In_1287,In_1587);
xnor U2264 (N_2264,In_1157,In_655);
xnor U2265 (N_2265,In_1821,In_553);
xnor U2266 (N_2266,In_374,In_1557);
and U2267 (N_2267,In_830,In_2188);
xnor U2268 (N_2268,In_48,In_345);
or U2269 (N_2269,In_110,In_2276);
xor U2270 (N_2270,In_1962,In_2106);
nand U2271 (N_2271,In_705,In_118);
and U2272 (N_2272,In_1306,In_1122);
nand U2273 (N_2273,In_1055,In_321);
xor U2274 (N_2274,In_1672,In_1068);
xor U2275 (N_2275,In_784,In_1226);
or U2276 (N_2276,In_2363,In_416);
nor U2277 (N_2277,In_1953,In_1587);
and U2278 (N_2278,In_2484,In_1362);
nand U2279 (N_2279,In_956,In_418);
nand U2280 (N_2280,In_1000,In_387);
nor U2281 (N_2281,In_1952,In_1471);
or U2282 (N_2282,In_1744,In_907);
xnor U2283 (N_2283,In_837,In_2131);
xor U2284 (N_2284,In_1078,In_28);
xnor U2285 (N_2285,In_1195,In_1421);
or U2286 (N_2286,In_1490,In_1480);
and U2287 (N_2287,In_1539,In_446);
nor U2288 (N_2288,In_597,In_959);
nor U2289 (N_2289,In_791,In_1331);
and U2290 (N_2290,In_625,In_2125);
or U2291 (N_2291,In_509,In_1782);
or U2292 (N_2292,In_592,In_1623);
or U2293 (N_2293,In_2461,In_118);
xnor U2294 (N_2294,In_2292,In_861);
or U2295 (N_2295,In_1498,In_1101);
xor U2296 (N_2296,In_876,In_1424);
and U2297 (N_2297,In_830,In_1511);
xor U2298 (N_2298,In_1290,In_36);
xor U2299 (N_2299,In_1312,In_2478);
nor U2300 (N_2300,In_407,In_1478);
xor U2301 (N_2301,In_1334,In_213);
nand U2302 (N_2302,In_1897,In_2468);
and U2303 (N_2303,In_861,In_1439);
and U2304 (N_2304,In_332,In_964);
nor U2305 (N_2305,In_1459,In_652);
and U2306 (N_2306,In_454,In_456);
xnor U2307 (N_2307,In_1876,In_91);
xor U2308 (N_2308,In_2095,In_1135);
and U2309 (N_2309,In_582,In_122);
nor U2310 (N_2310,In_1386,In_412);
or U2311 (N_2311,In_908,In_1493);
xor U2312 (N_2312,In_582,In_2245);
nor U2313 (N_2313,In_2019,In_2269);
nor U2314 (N_2314,In_233,In_413);
or U2315 (N_2315,In_608,In_1639);
nor U2316 (N_2316,In_1102,In_531);
or U2317 (N_2317,In_185,In_734);
nand U2318 (N_2318,In_956,In_1473);
and U2319 (N_2319,In_1179,In_558);
nand U2320 (N_2320,In_696,In_322);
nor U2321 (N_2321,In_1528,In_543);
and U2322 (N_2322,In_714,In_171);
and U2323 (N_2323,In_434,In_2341);
or U2324 (N_2324,In_2275,In_260);
nand U2325 (N_2325,In_142,In_1859);
nor U2326 (N_2326,In_274,In_1864);
nand U2327 (N_2327,In_2248,In_1342);
xor U2328 (N_2328,In_33,In_1726);
nor U2329 (N_2329,In_1952,In_191);
nand U2330 (N_2330,In_817,In_2269);
nor U2331 (N_2331,In_233,In_723);
xor U2332 (N_2332,In_2230,In_1918);
or U2333 (N_2333,In_1558,In_2184);
xnor U2334 (N_2334,In_25,In_2303);
and U2335 (N_2335,In_1577,In_2463);
nand U2336 (N_2336,In_1388,In_2055);
and U2337 (N_2337,In_2297,In_1037);
or U2338 (N_2338,In_1864,In_49);
nand U2339 (N_2339,In_751,In_19);
nor U2340 (N_2340,In_700,In_1619);
xor U2341 (N_2341,In_1399,In_2073);
and U2342 (N_2342,In_645,In_1361);
xor U2343 (N_2343,In_921,In_283);
nand U2344 (N_2344,In_1402,In_953);
and U2345 (N_2345,In_640,In_2441);
or U2346 (N_2346,In_792,In_1412);
nor U2347 (N_2347,In_2058,In_616);
xor U2348 (N_2348,In_1588,In_1615);
xor U2349 (N_2349,In_788,In_2377);
nor U2350 (N_2350,In_179,In_345);
and U2351 (N_2351,In_1792,In_379);
or U2352 (N_2352,In_1944,In_2350);
nor U2353 (N_2353,In_1322,In_1792);
nand U2354 (N_2354,In_2412,In_1247);
or U2355 (N_2355,In_2125,In_2373);
or U2356 (N_2356,In_2454,In_1002);
or U2357 (N_2357,In_2093,In_2084);
xnor U2358 (N_2358,In_219,In_1652);
nand U2359 (N_2359,In_951,In_1010);
xnor U2360 (N_2360,In_1224,In_771);
xnor U2361 (N_2361,In_2092,In_253);
nand U2362 (N_2362,In_2196,In_1378);
or U2363 (N_2363,In_1146,In_2090);
nor U2364 (N_2364,In_644,In_424);
nor U2365 (N_2365,In_2483,In_2044);
and U2366 (N_2366,In_145,In_64);
and U2367 (N_2367,In_550,In_2069);
xor U2368 (N_2368,In_2447,In_748);
or U2369 (N_2369,In_868,In_1795);
nand U2370 (N_2370,In_2061,In_2244);
nor U2371 (N_2371,In_1776,In_791);
xnor U2372 (N_2372,In_758,In_714);
and U2373 (N_2373,In_1061,In_74);
or U2374 (N_2374,In_680,In_2151);
or U2375 (N_2375,In_1192,In_1750);
nand U2376 (N_2376,In_1486,In_168);
nor U2377 (N_2377,In_1429,In_2196);
nor U2378 (N_2378,In_287,In_856);
nor U2379 (N_2379,In_928,In_2182);
nor U2380 (N_2380,In_551,In_718);
nand U2381 (N_2381,In_300,In_713);
xnor U2382 (N_2382,In_1763,In_1979);
or U2383 (N_2383,In_1513,In_2263);
and U2384 (N_2384,In_74,In_697);
and U2385 (N_2385,In_1558,In_883);
nor U2386 (N_2386,In_1404,In_375);
nand U2387 (N_2387,In_1885,In_2429);
and U2388 (N_2388,In_66,In_158);
and U2389 (N_2389,In_2189,In_1732);
and U2390 (N_2390,In_1316,In_1058);
nand U2391 (N_2391,In_1317,In_311);
and U2392 (N_2392,In_1990,In_1934);
nor U2393 (N_2393,In_2342,In_119);
nor U2394 (N_2394,In_680,In_1996);
or U2395 (N_2395,In_1479,In_2461);
xor U2396 (N_2396,In_1847,In_1071);
or U2397 (N_2397,In_2341,In_292);
nand U2398 (N_2398,In_370,In_87);
nand U2399 (N_2399,In_1928,In_1151);
and U2400 (N_2400,In_2352,In_217);
nand U2401 (N_2401,In_1840,In_2039);
or U2402 (N_2402,In_29,In_1967);
or U2403 (N_2403,In_135,In_1436);
nand U2404 (N_2404,In_1324,In_20);
and U2405 (N_2405,In_676,In_953);
nand U2406 (N_2406,In_2451,In_171);
nor U2407 (N_2407,In_1197,In_1351);
nor U2408 (N_2408,In_2498,In_2361);
xor U2409 (N_2409,In_981,In_1016);
or U2410 (N_2410,In_1200,In_2492);
xnor U2411 (N_2411,In_2438,In_2475);
nor U2412 (N_2412,In_1855,In_1937);
nor U2413 (N_2413,In_1713,In_2108);
and U2414 (N_2414,In_2056,In_1426);
and U2415 (N_2415,In_2202,In_2112);
nand U2416 (N_2416,In_1243,In_1070);
and U2417 (N_2417,In_1487,In_1070);
or U2418 (N_2418,In_1280,In_1863);
or U2419 (N_2419,In_899,In_232);
or U2420 (N_2420,In_1866,In_1964);
or U2421 (N_2421,In_1745,In_1961);
or U2422 (N_2422,In_55,In_402);
nor U2423 (N_2423,In_55,In_1661);
nor U2424 (N_2424,In_240,In_1433);
nor U2425 (N_2425,In_2124,In_1004);
or U2426 (N_2426,In_29,In_1736);
or U2427 (N_2427,In_1511,In_1835);
xnor U2428 (N_2428,In_2454,In_1917);
or U2429 (N_2429,In_2287,In_387);
xnor U2430 (N_2430,In_270,In_2325);
xnor U2431 (N_2431,In_770,In_1719);
nor U2432 (N_2432,In_1639,In_2198);
and U2433 (N_2433,In_287,In_2452);
or U2434 (N_2434,In_1109,In_1050);
xor U2435 (N_2435,In_1,In_1417);
nand U2436 (N_2436,In_1565,In_1043);
and U2437 (N_2437,In_2398,In_194);
or U2438 (N_2438,In_445,In_552);
xnor U2439 (N_2439,In_1949,In_2150);
and U2440 (N_2440,In_1714,In_1896);
nand U2441 (N_2441,In_2280,In_1067);
or U2442 (N_2442,In_1563,In_2322);
xnor U2443 (N_2443,In_2482,In_2413);
nand U2444 (N_2444,In_1242,In_413);
nand U2445 (N_2445,In_948,In_55);
nor U2446 (N_2446,In_2293,In_1419);
nand U2447 (N_2447,In_2089,In_1113);
nand U2448 (N_2448,In_2307,In_2497);
nand U2449 (N_2449,In_2489,In_1203);
or U2450 (N_2450,In_1288,In_1924);
and U2451 (N_2451,In_1026,In_27);
or U2452 (N_2452,In_704,In_1776);
or U2453 (N_2453,In_972,In_2358);
and U2454 (N_2454,In_1299,In_993);
nor U2455 (N_2455,In_586,In_646);
or U2456 (N_2456,In_1686,In_1387);
nor U2457 (N_2457,In_1965,In_765);
or U2458 (N_2458,In_2417,In_1093);
nand U2459 (N_2459,In_935,In_758);
and U2460 (N_2460,In_1170,In_1564);
nor U2461 (N_2461,In_1505,In_984);
nor U2462 (N_2462,In_1500,In_1317);
or U2463 (N_2463,In_1764,In_689);
or U2464 (N_2464,In_2404,In_1756);
nor U2465 (N_2465,In_797,In_1101);
xnor U2466 (N_2466,In_1525,In_1476);
or U2467 (N_2467,In_2040,In_531);
or U2468 (N_2468,In_1991,In_2444);
xnor U2469 (N_2469,In_896,In_479);
or U2470 (N_2470,In_1873,In_2492);
nand U2471 (N_2471,In_2364,In_1079);
and U2472 (N_2472,In_1895,In_2493);
nor U2473 (N_2473,In_1466,In_1485);
and U2474 (N_2474,In_500,In_1208);
nor U2475 (N_2475,In_2395,In_166);
xnor U2476 (N_2476,In_94,In_699);
nand U2477 (N_2477,In_1805,In_2368);
nor U2478 (N_2478,In_2436,In_988);
nor U2479 (N_2479,In_695,In_1377);
nand U2480 (N_2480,In_399,In_755);
nor U2481 (N_2481,In_1859,In_862);
or U2482 (N_2482,In_2426,In_1355);
or U2483 (N_2483,In_1997,In_1226);
nor U2484 (N_2484,In_920,In_1807);
and U2485 (N_2485,In_202,In_2115);
and U2486 (N_2486,In_1652,In_168);
nor U2487 (N_2487,In_1352,In_1906);
or U2488 (N_2488,In_1877,In_1115);
or U2489 (N_2489,In_2235,In_694);
nor U2490 (N_2490,In_576,In_2453);
nor U2491 (N_2491,In_1105,In_2128);
nand U2492 (N_2492,In_2105,In_496);
nand U2493 (N_2493,In_949,In_492);
or U2494 (N_2494,In_2119,In_1810);
xnor U2495 (N_2495,In_792,In_1060);
xnor U2496 (N_2496,In_668,In_183);
xor U2497 (N_2497,In_307,In_524);
nor U2498 (N_2498,In_2371,In_981);
nor U2499 (N_2499,In_177,In_2281);
or U2500 (N_2500,In_1152,In_289);
or U2501 (N_2501,In_1190,In_2412);
nand U2502 (N_2502,In_250,In_676);
or U2503 (N_2503,In_154,In_2190);
or U2504 (N_2504,In_1813,In_2307);
xor U2505 (N_2505,In_1049,In_2490);
nand U2506 (N_2506,In_1916,In_1153);
or U2507 (N_2507,In_1315,In_682);
or U2508 (N_2508,In_476,In_446);
or U2509 (N_2509,In_322,In_633);
nor U2510 (N_2510,In_1208,In_1177);
and U2511 (N_2511,In_1732,In_1963);
nand U2512 (N_2512,In_632,In_1090);
nor U2513 (N_2513,In_1543,In_1937);
nand U2514 (N_2514,In_1163,In_2367);
nand U2515 (N_2515,In_792,In_368);
or U2516 (N_2516,In_1312,In_812);
or U2517 (N_2517,In_2111,In_1285);
and U2518 (N_2518,In_84,In_2087);
or U2519 (N_2519,In_812,In_428);
or U2520 (N_2520,In_1487,In_1377);
xnor U2521 (N_2521,In_1694,In_525);
xnor U2522 (N_2522,In_1202,In_1681);
xor U2523 (N_2523,In_1532,In_1403);
or U2524 (N_2524,In_51,In_452);
nand U2525 (N_2525,In_1541,In_2022);
nor U2526 (N_2526,In_458,In_2457);
and U2527 (N_2527,In_2208,In_2062);
or U2528 (N_2528,In_669,In_2164);
nand U2529 (N_2529,In_1879,In_1191);
nand U2530 (N_2530,In_1762,In_1444);
or U2531 (N_2531,In_2223,In_1490);
and U2532 (N_2532,In_602,In_2204);
nor U2533 (N_2533,In_56,In_1779);
nand U2534 (N_2534,In_686,In_1116);
and U2535 (N_2535,In_2004,In_2350);
and U2536 (N_2536,In_504,In_1505);
xnor U2537 (N_2537,In_1936,In_2423);
or U2538 (N_2538,In_932,In_2264);
xor U2539 (N_2539,In_661,In_1769);
or U2540 (N_2540,In_661,In_12);
or U2541 (N_2541,In_124,In_1865);
xor U2542 (N_2542,In_1531,In_1993);
xor U2543 (N_2543,In_323,In_274);
or U2544 (N_2544,In_2430,In_1588);
nor U2545 (N_2545,In_1600,In_72);
and U2546 (N_2546,In_2237,In_2463);
nor U2547 (N_2547,In_985,In_2173);
and U2548 (N_2548,In_1781,In_1802);
xor U2549 (N_2549,In_1158,In_1305);
and U2550 (N_2550,In_2209,In_166);
xnor U2551 (N_2551,In_315,In_77);
xor U2552 (N_2552,In_555,In_1620);
and U2553 (N_2553,In_750,In_1382);
and U2554 (N_2554,In_2492,In_858);
xnor U2555 (N_2555,In_2303,In_668);
nor U2556 (N_2556,In_2382,In_1239);
nand U2557 (N_2557,In_1588,In_1814);
nor U2558 (N_2558,In_1228,In_1526);
or U2559 (N_2559,In_400,In_873);
and U2560 (N_2560,In_1498,In_1714);
or U2561 (N_2561,In_637,In_663);
and U2562 (N_2562,In_1564,In_404);
nor U2563 (N_2563,In_265,In_1348);
xnor U2564 (N_2564,In_1492,In_993);
xor U2565 (N_2565,In_1405,In_312);
or U2566 (N_2566,In_2369,In_2346);
nor U2567 (N_2567,In_699,In_1985);
xor U2568 (N_2568,In_617,In_1054);
xnor U2569 (N_2569,In_1308,In_1840);
and U2570 (N_2570,In_2231,In_1540);
nand U2571 (N_2571,In_2362,In_1002);
or U2572 (N_2572,In_2056,In_94);
nand U2573 (N_2573,In_1894,In_2414);
xor U2574 (N_2574,In_2134,In_1583);
and U2575 (N_2575,In_2006,In_1533);
or U2576 (N_2576,In_1868,In_1364);
nor U2577 (N_2577,In_1717,In_1556);
xnor U2578 (N_2578,In_1103,In_1456);
or U2579 (N_2579,In_407,In_1833);
nand U2580 (N_2580,In_35,In_1663);
xor U2581 (N_2581,In_1417,In_335);
nor U2582 (N_2582,In_1994,In_2190);
xnor U2583 (N_2583,In_1251,In_2397);
nor U2584 (N_2584,In_1050,In_854);
nand U2585 (N_2585,In_2297,In_775);
nand U2586 (N_2586,In_2319,In_1564);
nand U2587 (N_2587,In_1388,In_1077);
nor U2588 (N_2588,In_2290,In_838);
xor U2589 (N_2589,In_1793,In_360);
nand U2590 (N_2590,In_2192,In_2370);
and U2591 (N_2591,In_2397,In_28);
nand U2592 (N_2592,In_1568,In_2295);
and U2593 (N_2593,In_1647,In_80);
or U2594 (N_2594,In_1753,In_2306);
or U2595 (N_2595,In_759,In_969);
xor U2596 (N_2596,In_1175,In_2290);
or U2597 (N_2597,In_51,In_1731);
xnor U2598 (N_2598,In_1227,In_238);
xor U2599 (N_2599,In_1356,In_1248);
and U2600 (N_2600,In_728,In_474);
nor U2601 (N_2601,In_2362,In_385);
nor U2602 (N_2602,In_1270,In_717);
xor U2603 (N_2603,In_1752,In_1746);
or U2604 (N_2604,In_2031,In_2125);
xnor U2605 (N_2605,In_1229,In_624);
xor U2606 (N_2606,In_453,In_1730);
nand U2607 (N_2607,In_1490,In_1498);
xnor U2608 (N_2608,In_1099,In_2499);
xor U2609 (N_2609,In_498,In_1680);
xnor U2610 (N_2610,In_162,In_1676);
xnor U2611 (N_2611,In_1756,In_1013);
and U2612 (N_2612,In_1764,In_538);
or U2613 (N_2613,In_1358,In_426);
or U2614 (N_2614,In_1207,In_2307);
nand U2615 (N_2615,In_2264,In_440);
nor U2616 (N_2616,In_2451,In_1954);
or U2617 (N_2617,In_392,In_2292);
and U2618 (N_2618,In_458,In_437);
and U2619 (N_2619,In_601,In_1987);
nand U2620 (N_2620,In_1328,In_963);
xor U2621 (N_2621,In_1013,In_1221);
nor U2622 (N_2622,In_2237,In_1402);
nand U2623 (N_2623,In_1857,In_318);
nor U2624 (N_2624,In_144,In_833);
and U2625 (N_2625,In_1373,In_2225);
nand U2626 (N_2626,In_1077,In_1879);
nand U2627 (N_2627,In_418,In_550);
nor U2628 (N_2628,In_1307,In_1380);
nor U2629 (N_2629,In_1760,In_258);
nand U2630 (N_2630,In_879,In_663);
nor U2631 (N_2631,In_1261,In_284);
or U2632 (N_2632,In_1844,In_106);
nor U2633 (N_2633,In_2256,In_1354);
nand U2634 (N_2634,In_510,In_795);
xnor U2635 (N_2635,In_267,In_769);
xnor U2636 (N_2636,In_1493,In_1430);
and U2637 (N_2637,In_2039,In_2015);
xnor U2638 (N_2638,In_1279,In_182);
or U2639 (N_2639,In_1670,In_207);
nand U2640 (N_2640,In_2242,In_1448);
nand U2641 (N_2641,In_2028,In_221);
and U2642 (N_2642,In_1503,In_906);
or U2643 (N_2643,In_718,In_2116);
or U2644 (N_2644,In_340,In_386);
and U2645 (N_2645,In_146,In_348);
nor U2646 (N_2646,In_1771,In_1504);
xnor U2647 (N_2647,In_975,In_1932);
and U2648 (N_2648,In_1229,In_742);
nand U2649 (N_2649,In_1215,In_1989);
xnor U2650 (N_2650,In_1231,In_1751);
xnor U2651 (N_2651,In_1994,In_2335);
xnor U2652 (N_2652,In_438,In_2011);
and U2653 (N_2653,In_679,In_587);
and U2654 (N_2654,In_1134,In_1722);
and U2655 (N_2655,In_318,In_818);
nand U2656 (N_2656,In_1138,In_1535);
and U2657 (N_2657,In_2359,In_1249);
and U2658 (N_2658,In_632,In_964);
and U2659 (N_2659,In_559,In_763);
xor U2660 (N_2660,In_1845,In_785);
and U2661 (N_2661,In_1295,In_2417);
and U2662 (N_2662,In_1258,In_641);
and U2663 (N_2663,In_419,In_176);
or U2664 (N_2664,In_710,In_311);
nand U2665 (N_2665,In_563,In_2387);
nand U2666 (N_2666,In_1102,In_205);
nand U2667 (N_2667,In_2418,In_1035);
xnor U2668 (N_2668,In_1017,In_2221);
nor U2669 (N_2669,In_54,In_644);
or U2670 (N_2670,In_599,In_1996);
nor U2671 (N_2671,In_7,In_1538);
nor U2672 (N_2672,In_1292,In_1045);
xnor U2673 (N_2673,In_71,In_1834);
nor U2674 (N_2674,In_2067,In_2150);
nor U2675 (N_2675,In_1663,In_1366);
or U2676 (N_2676,In_1063,In_1332);
or U2677 (N_2677,In_1788,In_1906);
nand U2678 (N_2678,In_1327,In_967);
and U2679 (N_2679,In_464,In_2264);
and U2680 (N_2680,In_2223,In_34);
nand U2681 (N_2681,In_482,In_1946);
nand U2682 (N_2682,In_2097,In_2358);
nor U2683 (N_2683,In_1072,In_2166);
or U2684 (N_2684,In_1545,In_1366);
nor U2685 (N_2685,In_821,In_1302);
and U2686 (N_2686,In_243,In_1972);
nand U2687 (N_2687,In_2067,In_1669);
nand U2688 (N_2688,In_1584,In_928);
nor U2689 (N_2689,In_1539,In_1432);
nand U2690 (N_2690,In_330,In_1252);
or U2691 (N_2691,In_255,In_1826);
xnor U2692 (N_2692,In_1057,In_997);
xnor U2693 (N_2693,In_378,In_78);
xnor U2694 (N_2694,In_1646,In_2338);
xor U2695 (N_2695,In_1242,In_1628);
or U2696 (N_2696,In_2241,In_1615);
xor U2697 (N_2697,In_141,In_1756);
nor U2698 (N_2698,In_727,In_2373);
nor U2699 (N_2699,In_1928,In_1488);
or U2700 (N_2700,In_1225,In_920);
or U2701 (N_2701,In_2080,In_1949);
nor U2702 (N_2702,In_832,In_794);
nand U2703 (N_2703,In_1531,In_1732);
xnor U2704 (N_2704,In_140,In_2405);
nor U2705 (N_2705,In_161,In_1040);
nor U2706 (N_2706,In_1253,In_260);
xor U2707 (N_2707,In_11,In_1262);
xor U2708 (N_2708,In_1848,In_117);
and U2709 (N_2709,In_420,In_908);
and U2710 (N_2710,In_115,In_437);
nor U2711 (N_2711,In_106,In_1941);
and U2712 (N_2712,In_2199,In_2193);
or U2713 (N_2713,In_1047,In_84);
nor U2714 (N_2714,In_1164,In_743);
or U2715 (N_2715,In_1083,In_1376);
nand U2716 (N_2716,In_1841,In_2278);
nor U2717 (N_2717,In_1629,In_1109);
xnor U2718 (N_2718,In_1291,In_2300);
nand U2719 (N_2719,In_178,In_298);
and U2720 (N_2720,In_277,In_1317);
and U2721 (N_2721,In_1016,In_1832);
and U2722 (N_2722,In_2417,In_1140);
nand U2723 (N_2723,In_1168,In_971);
nor U2724 (N_2724,In_1222,In_1134);
or U2725 (N_2725,In_911,In_1121);
xor U2726 (N_2726,In_1983,In_1886);
xnor U2727 (N_2727,In_2091,In_753);
nor U2728 (N_2728,In_65,In_359);
nor U2729 (N_2729,In_826,In_1500);
nor U2730 (N_2730,In_266,In_2415);
xor U2731 (N_2731,In_1877,In_1947);
nor U2732 (N_2732,In_1061,In_2454);
xor U2733 (N_2733,In_2254,In_711);
nor U2734 (N_2734,In_1204,In_2374);
nand U2735 (N_2735,In_1049,In_154);
nor U2736 (N_2736,In_734,In_2131);
nand U2737 (N_2737,In_2074,In_170);
xnor U2738 (N_2738,In_433,In_2066);
xor U2739 (N_2739,In_1397,In_30);
or U2740 (N_2740,In_2006,In_1020);
nor U2741 (N_2741,In_2256,In_79);
nand U2742 (N_2742,In_629,In_2039);
nand U2743 (N_2743,In_559,In_1356);
and U2744 (N_2744,In_1171,In_883);
nor U2745 (N_2745,In_1876,In_1256);
xnor U2746 (N_2746,In_567,In_463);
xor U2747 (N_2747,In_301,In_1384);
or U2748 (N_2748,In_197,In_906);
nand U2749 (N_2749,In_1441,In_2314);
and U2750 (N_2750,In_2418,In_1003);
xor U2751 (N_2751,In_232,In_932);
nand U2752 (N_2752,In_1129,In_750);
or U2753 (N_2753,In_2337,In_239);
nand U2754 (N_2754,In_1931,In_2251);
nor U2755 (N_2755,In_2379,In_261);
nor U2756 (N_2756,In_1268,In_1870);
nor U2757 (N_2757,In_1326,In_242);
or U2758 (N_2758,In_2456,In_1215);
nand U2759 (N_2759,In_1065,In_538);
and U2760 (N_2760,In_1134,In_2189);
xnor U2761 (N_2761,In_188,In_1767);
nand U2762 (N_2762,In_1573,In_868);
and U2763 (N_2763,In_1848,In_1684);
or U2764 (N_2764,In_1204,In_1242);
or U2765 (N_2765,In_1454,In_298);
or U2766 (N_2766,In_281,In_881);
xnor U2767 (N_2767,In_1964,In_2258);
or U2768 (N_2768,In_2110,In_1987);
or U2769 (N_2769,In_285,In_330);
nand U2770 (N_2770,In_1946,In_2313);
nand U2771 (N_2771,In_1805,In_2487);
or U2772 (N_2772,In_1111,In_1621);
nor U2773 (N_2773,In_2416,In_342);
nor U2774 (N_2774,In_650,In_181);
nand U2775 (N_2775,In_96,In_1242);
nor U2776 (N_2776,In_1737,In_348);
nor U2777 (N_2777,In_1917,In_2402);
nor U2778 (N_2778,In_819,In_1434);
or U2779 (N_2779,In_1228,In_953);
nor U2780 (N_2780,In_719,In_95);
xnor U2781 (N_2781,In_2088,In_783);
nor U2782 (N_2782,In_995,In_2277);
nor U2783 (N_2783,In_2391,In_71);
xnor U2784 (N_2784,In_443,In_1584);
nand U2785 (N_2785,In_748,In_2223);
or U2786 (N_2786,In_398,In_1832);
xnor U2787 (N_2787,In_2214,In_564);
xor U2788 (N_2788,In_837,In_2312);
nor U2789 (N_2789,In_2445,In_1071);
or U2790 (N_2790,In_176,In_339);
nor U2791 (N_2791,In_965,In_1902);
nand U2792 (N_2792,In_2485,In_1493);
nor U2793 (N_2793,In_1459,In_641);
nand U2794 (N_2794,In_561,In_1943);
and U2795 (N_2795,In_234,In_1996);
xnor U2796 (N_2796,In_1284,In_1013);
xor U2797 (N_2797,In_1594,In_325);
or U2798 (N_2798,In_850,In_2430);
nor U2799 (N_2799,In_286,In_2256);
and U2800 (N_2800,In_545,In_1659);
nand U2801 (N_2801,In_1609,In_2197);
and U2802 (N_2802,In_2455,In_1257);
nor U2803 (N_2803,In_2077,In_1513);
or U2804 (N_2804,In_2474,In_985);
nor U2805 (N_2805,In_1513,In_33);
or U2806 (N_2806,In_991,In_873);
and U2807 (N_2807,In_1636,In_988);
or U2808 (N_2808,In_1255,In_180);
nand U2809 (N_2809,In_161,In_1503);
and U2810 (N_2810,In_1103,In_1243);
and U2811 (N_2811,In_160,In_1091);
nand U2812 (N_2812,In_1683,In_376);
and U2813 (N_2813,In_2442,In_1810);
or U2814 (N_2814,In_1555,In_10);
nor U2815 (N_2815,In_1907,In_176);
nor U2816 (N_2816,In_2047,In_69);
nor U2817 (N_2817,In_795,In_2486);
or U2818 (N_2818,In_900,In_421);
and U2819 (N_2819,In_2048,In_1187);
and U2820 (N_2820,In_1850,In_841);
and U2821 (N_2821,In_2130,In_1786);
xor U2822 (N_2822,In_1737,In_2338);
or U2823 (N_2823,In_1258,In_876);
xor U2824 (N_2824,In_899,In_2133);
nand U2825 (N_2825,In_1221,In_1570);
or U2826 (N_2826,In_2473,In_2467);
and U2827 (N_2827,In_115,In_177);
xnor U2828 (N_2828,In_2178,In_2191);
nor U2829 (N_2829,In_1857,In_350);
xnor U2830 (N_2830,In_2091,In_1152);
xnor U2831 (N_2831,In_1854,In_1024);
xor U2832 (N_2832,In_1249,In_534);
xnor U2833 (N_2833,In_1352,In_2267);
nor U2834 (N_2834,In_1775,In_689);
and U2835 (N_2835,In_637,In_839);
or U2836 (N_2836,In_1928,In_1046);
nor U2837 (N_2837,In_1274,In_17);
or U2838 (N_2838,In_1935,In_160);
nand U2839 (N_2839,In_613,In_1823);
or U2840 (N_2840,In_1277,In_484);
or U2841 (N_2841,In_2299,In_1519);
or U2842 (N_2842,In_1245,In_602);
nor U2843 (N_2843,In_955,In_638);
and U2844 (N_2844,In_902,In_825);
nand U2845 (N_2845,In_688,In_25);
or U2846 (N_2846,In_1695,In_2384);
nand U2847 (N_2847,In_155,In_1791);
nand U2848 (N_2848,In_646,In_1268);
and U2849 (N_2849,In_683,In_2363);
nor U2850 (N_2850,In_998,In_117);
or U2851 (N_2851,In_1780,In_1960);
and U2852 (N_2852,In_83,In_199);
and U2853 (N_2853,In_1057,In_1123);
nand U2854 (N_2854,In_107,In_1303);
and U2855 (N_2855,In_721,In_565);
xnor U2856 (N_2856,In_1805,In_2141);
or U2857 (N_2857,In_1988,In_708);
or U2858 (N_2858,In_532,In_141);
nand U2859 (N_2859,In_836,In_369);
or U2860 (N_2860,In_1825,In_743);
and U2861 (N_2861,In_523,In_1684);
nor U2862 (N_2862,In_2006,In_309);
xor U2863 (N_2863,In_580,In_1037);
xnor U2864 (N_2864,In_1875,In_2275);
xnor U2865 (N_2865,In_1720,In_1897);
and U2866 (N_2866,In_281,In_2272);
or U2867 (N_2867,In_2441,In_746);
xnor U2868 (N_2868,In_628,In_1340);
nand U2869 (N_2869,In_2301,In_1127);
or U2870 (N_2870,In_216,In_1468);
nor U2871 (N_2871,In_352,In_870);
nor U2872 (N_2872,In_1700,In_1194);
nand U2873 (N_2873,In_2461,In_1803);
nor U2874 (N_2874,In_1550,In_1134);
and U2875 (N_2875,In_1388,In_550);
nand U2876 (N_2876,In_765,In_1604);
nor U2877 (N_2877,In_1772,In_1374);
and U2878 (N_2878,In_1015,In_1749);
or U2879 (N_2879,In_474,In_2204);
or U2880 (N_2880,In_1402,In_2209);
or U2881 (N_2881,In_844,In_9);
nor U2882 (N_2882,In_1732,In_914);
or U2883 (N_2883,In_400,In_1770);
or U2884 (N_2884,In_2237,In_1235);
nand U2885 (N_2885,In_1718,In_673);
and U2886 (N_2886,In_1339,In_2292);
nand U2887 (N_2887,In_1884,In_2259);
nand U2888 (N_2888,In_704,In_1301);
xor U2889 (N_2889,In_1103,In_577);
nand U2890 (N_2890,In_412,In_164);
nor U2891 (N_2891,In_635,In_278);
or U2892 (N_2892,In_601,In_645);
nand U2893 (N_2893,In_1980,In_373);
and U2894 (N_2894,In_1494,In_1839);
xnor U2895 (N_2895,In_1244,In_26);
xor U2896 (N_2896,In_1317,In_259);
nand U2897 (N_2897,In_2480,In_2275);
nor U2898 (N_2898,In_125,In_1307);
xor U2899 (N_2899,In_116,In_428);
nor U2900 (N_2900,In_1608,In_1440);
nor U2901 (N_2901,In_2271,In_1344);
and U2902 (N_2902,In_1380,In_736);
and U2903 (N_2903,In_1732,In_2164);
nand U2904 (N_2904,In_2232,In_45);
or U2905 (N_2905,In_2311,In_1554);
xor U2906 (N_2906,In_2104,In_1292);
xnor U2907 (N_2907,In_2351,In_501);
or U2908 (N_2908,In_1174,In_1305);
xnor U2909 (N_2909,In_2019,In_1515);
nand U2910 (N_2910,In_583,In_1113);
nand U2911 (N_2911,In_955,In_1890);
and U2912 (N_2912,In_2219,In_887);
nor U2913 (N_2913,In_45,In_1068);
or U2914 (N_2914,In_911,In_2049);
or U2915 (N_2915,In_933,In_1120);
and U2916 (N_2916,In_1202,In_90);
or U2917 (N_2917,In_1040,In_699);
nor U2918 (N_2918,In_2396,In_1723);
and U2919 (N_2919,In_403,In_1204);
nor U2920 (N_2920,In_732,In_869);
and U2921 (N_2921,In_2209,In_2411);
nand U2922 (N_2922,In_1001,In_1880);
nor U2923 (N_2923,In_2261,In_2250);
and U2924 (N_2924,In_2288,In_2328);
or U2925 (N_2925,In_2116,In_1982);
nand U2926 (N_2926,In_290,In_360);
xnor U2927 (N_2927,In_1502,In_2237);
nor U2928 (N_2928,In_2412,In_655);
and U2929 (N_2929,In_851,In_1806);
and U2930 (N_2930,In_2197,In_1686);
nand U2931 (N_2931,In_353,In_1952);
and U2932 (N_2932,In_613,In_1146);
nor U2933 (N_2933,In_604,In_1571);
nor U2934 (N_2934,In_624,In_879);
or U2935 (N_2935,In_783,In_1293);
nand U2936 (N_2936,In_1606,In_818);
nand U2937 (N_2937,In_2248,In_1051);
and U2938 (N_2938,In_1450,In_583);
and U2939 (N_2939,In_880,In_1254);
and U2940 (N_2940,In_1286,In_727);
nand U2941 (N_2941,In_1926,In_1637);
nand U2942 (N_2942,In_2438,In_38);
and U2943 (N_2943,In_1899,In_1929);
xnor U2944 (N_2944,In_1740,In_436);
nor U2945 (N_2945,In_207,In_182);
or U2946 (N_2946,In_1853,In_2082);
xnor U2947 (N_2947,In_235,In_1929);
or U2948 (N_2948,In_295,In_2206);
xnor U2949 (N_2949,In_1160,In_2094);
nand U2950 (N_2950,In_250,In_1716);
and U2951 (N_2951,In_271,In_1527);
and U2952 (N_2952,In_365,In_1281);
nand U2953 (N_2953,In_2197,In_617);
and U2954 (N_2954,In_272,In_765);
nor U2955 (N_2955,In_2372,In_306);
or U2956 (N_2956,In_1557,In_1677);
nand U2957 (N_2957,In_1787,In_1423);
xnor U2958 (N_2958,In_981,In_649);
or U2959 (N_2959,In_1355,In_2381);
xnor U2960 (N_2960,In_1865,In_1342);
and U2961 (N_2961,In_567,In_220);
nor U2962 (N_2962,In_2431,In_302);
nor U2963 (N_2963,In_749,In_1021);
nand U2964 (N_2964,In_1156,In_92);
nor U2965 (N_2965,In_2335,In_259);
and U2966 (N_2966,In_1006,In_545);
and U2967 (N_2967,In_673,In_1754);
xnor U2968 (N_2968,In_1228,In_1139);
nor U2969 (N_2969,In_1849,In_1756);
nor U2970 (N_2970,In_2396,In_1334);
and U2971 (N_2971,In_645,In_2414);
xnor U2972 (N_2972,In_134,In_1504);
xor U2973 (N_2973,In_144,In_1622);
nand U2974 (N_2974,In_540,In_2091);
nor U2975 (N_2975,In_566,In_1995);
nor U2976 (N_2976,In_1797,In_1944);
xnor U2977 (N_2977,In_1880,In_2458);
and U2978 (N_2978,In_859,In_2219);
nor U2979 (N_2979,In_1247,In_1605);
xor U2980 (N_2980,In_2119,In_1527);
nand U2981 (N_2981,In_1623,In_238);
or U2982 (N_2982,In_799,In_35);
or U2983 (N_2983,In_785,In_515);
and U2984 (N_2984,In_2043,In_2195);
nor U2985 (N_2985,In_710,In_1791);
nor U2986 (N_2986,In_261,In_929);
nor U2987 (N_2987,In_1447,In_545);
and U2988 (N_2988,In_591,In_99);
nand U2989 (N_2989,In_2497,In_495);
nand U2990 (N_2990,In_1407,In_1405);
and U2991 (N_2991,In_536,In_2120);
nand U2992 (N_2992,In_1882,In_323);
xor U2993 (N_2993,In_1939,In_1204);
or U2994 (N_2994,In_583,In_2174);
or U2995 (N_2995,In_545,In_1358);
xnor U2996 (N_2996,In_1977,In_1074);
xnor U2997 (N_2997,In_1709,In_2495);
nand U2998 (N_2998,In_2494,In_719);
nor U2999 (N_2999,In_1729,In_2385);
xor U3000 (N_3000,In_1321,In_285);
and U3001 (N_3001,In_974,In_2403);
nand U3002 (N_3002,In_1538,In_415);
and U3003 (N_3003,In_698,In_1829);
and U3004 (N_3004,In_1454,In_2357);
and U3005 (N_3005,In_598,In_1084);
or U3006 (N_3006,In_454,In_553);
nand U3007 (N_3007,In_1611,In_2341);
and U3008 (N_3008,In_1652,In_2381);
xnor U3009 (N_3009,In_296,In_935);
or U3010 (N_3010,In_10,In_2315);
xnor U3011 (N_3011,In_2326,In_297);
or U3012 (N_3012,In_2446,In_1103);
xnor U3013 (N_3013,In_2433,In_693);
and U3014 (N_3014,In_1704,In_27);
and U3015 (N_3015,In_2194,In_4);
and U3016 (N_3016,In_1054,In_1711);
and U3017 (N_3017,In_815,In_1913);
nor U3018 (N_3018,In_324,In_661);
nor U3019 (N_3019,In_2047,In_456);
xnor U3020 (N_3020,In_1852,In_591);
nor U3021 (N_3021,In_1327,In_1662);
and U3022 (N_3022,In_589,In_725);
nand U3023 (N_3023,In_1915,In_1679);
and U3024 (N_3024,In_342,In_1598);
and U3025 (N_3025,In_2421,In_698);
and U3026 (N_3026,In_1879,In_943);
xor U3027 (N_3027,In_1031,In_1933);
nand U3028 (N_3028,In_974,In_1460);
or U3029 (N_3029,In_2345,In_1157);
and U3030 (N_3030,In_443,In_2355);
nor U3031 (N_3031,In_611,In_207);
nor U3032 (N_3032,In_1128,In_2342);
or U3033 (N_3033,In_1649,In_2386);
xor U3034 (N_3034,In_442,In_2219);
xor U3035 (N_3035,In_62,In_2499);
nor U3036 (N_3036,In_2248,In_2103);
and U3037 (N_3037,In_1540,In_1786);
and U3038 (N_3038,In_2016,In_1098);
nor U3039 (N_3039,In_1471,In_453);
xor U3040 (N_3040,In_435,In_2149);
or U3041 (N_3041,In_1638,In_2255);
or U3042 (N_3042,In_1847,In_296);
nand U3043 (N_3043,In_641,In_442);
and U3044 (N_3044,In_1485,In_872);
or U3045 (N_3045,In_2059,In_1099);
and U3046 (N_3046,In_1958,In_1318);
nand U3047 (N_3047,In_1835,In_1810);
nand U3048 (N_3048,In_1637,In_1809);
nor U3049 (N_3049,In_925,In_2105);
xnor U3050 (N_3050,In_1065,In_2000);
and U3051 (N_3051,In_158,In_2296);
xor U3052 (N_3052,In_1151,In_801);
xor U3053 (N_3053,In_2124,In_572);
nand U3054 (N_3054,In_2404,In_2059);
xor U3055 (N_3055,In_584,In_157);
xnor U3056 (N_3056,In_467,In_1407);
nor U3057 (N_3057,In_100,In_2374);
nor U3058 (N_3058,In_2008,In_2003);
or U3059 (N_3059,In_2240,In_2403);
xnor U3060 (N_3060,In_1431,In_2356);
nand U3061 (N_3061,In_1598,In_363);
or U3062 (N_3062,In_2414,In_3);
or U3063 (N_3063,In_1090,In_300);
xor U3064 (N_3064,In_784,In_128);
xnor U3065 (N_3065,In_874,In_1849);
nand U3066 (N_3066,In_1971,In_369);
and U3067 (N_3067,In_2410,In_1498);
or U3068 (N_3068,In_1622,In_1557);
nor U3069 (N_3069,In_297,In_2453);
nand U3070 (N_3070,In_1623,In_1637);
xnor U3071 (N_3071,In_2302,In_1591);
nor U3072 (N_3072,In_522,In_2484);
nor U3073 (N_3073,In_2367,In_2355);
and U3074 (N_3074,In_535,In_2264);
nand U3075 (N_3075,In_31,In_1259);
nor U3076 (N_3076,In_678,In_920);
or U3077 (N_3077,In_2302,In_1921);
and U3078 (N_3078,In_1043,In_1436);
xor U3079 (N_3079,In_671,In_1226);
nor U3080 (N_3080,In_1466,In_2231);
nor U3081 (N_3081,In_278,In_722);
and U3082 (N_3082,In_2168,In_1018);
and U3083 (N_3083,In_1153,In_1490);
or U3084 (N_3084,In_2306,In_2368);
xnor U3085 (N_3085,In_2139,In_2311);
nand U3086 (N_3086,In_1702,In_384);
or U3087 (N_3087,In_961,In_1279);
xnor U3088 (N_3088,In_509,In_1117);
and U3089 (N_3089,In_2362,In_204);
xnor U3090 (N_3090,In_129,In_71);
xor U3091 (N_3091,In_1228,In_201);
and U3092 (N_3092,In_94,In_1678);
or U3093 (N_3093,In_554,In_1596);
and U3094 (N_3094,In_7,In_352);
and U3095 (N_3095,In_929,In_729);
or U3096 (N_3096,In_370,In_531);
xnor U3097 (N_3097,In_579,In_653);
nand U3098 (N_3098,In_1344,In_573);
nor U3099 (N_3099,In_2249,In_1065);
nand U3100 (N_3100,In_433,In_1842);
nor U3101 (N_3101,In_97,In_2087);
nand U3102 (N_3102,In_2320,In_368);
or U3103 (N_3103,In_1796,In_2235);
nand U3104 (N_3104,In_1085,In_1058);
nor U3105 (N_3105,In_1034,In_1570);
nand U3106 (N_3106,In_1117,In_599);
and U3107 (N_3107,In_2426,In_1930);
xnor U3108 (N_3108,In_2306,In_1874);
and U3109 (N_3109,In_493,In_2161);
nor U3110 (N_3110,In_1517,In_2113);
xor U3111 (N_3111,In_64,In_2432);
nor U3112 (N_3112,In_1785,In_1337);
xnor U3113 (N_3113,In_775,In_556);
xnor U3114 (N_3114,In_139,In_189);
or U3115 (N_3115,In_1709,In_833);
xor U3116 (N_3116,In_2051,In_727);
xnor U3117 (N_3117,In_1578,In_814);
and U3118 (N_3118,In_1357,In_267);
nand U3119 (N_3119,In_258,In_109);
xor U3120 (N_3120,In_1509,In_1507);
or U3121 (N_3121,In_1421,In_599);
nor U3122 (N_3122,In_875,In_849);
and U3123 (N_3123,In_441,In_1574);
or U3124 (N_3124,In_568,In_692);
nor U3125 (N_3125,N_287,N_1338);
or U3126 (N_3126,N_640,N_1008);
nand U3127 (N_3127,N_1570,N_2674);
or U3128 (N_3128,N_30,N_1414);
nand U3129 (N_3129,N_2248,N_2390);
or U3130 (N_3130,N_803,N_1676);
or U3131 (N_3131,N_987,N_196);
nand U3132 (N_3132,N_608,N_2693);
and U3133 (N_3133,N_1751,N_2210);
and U3134 (N_3134,N_892,N_2446);
nand U3135 (N_3135,N_569,N_1803);
and U3136 (N_3136,N_1245,N_3055);
or U3137 (N_3137,N_2331,N_2477);
nor U3138 (N_3138,N_1019,N_3000);
and U3139 (N_3139,N_2858,N_2193);
nor U3140 (N_3140,N_2527,N_2841);
and U3141 (N_3141,N_687,N_2132);
or U3142 (N_3142,N_1731,N_2142);
and U3143 (N_3143,N_75,N_80);
and U3144 (N_3144,N_2174,N_2654);
or U3145 (N_3145,N_3114,N_1481);
nand U3146 (N_3146,N_877,N_1643);
and U3147 (N_3147,N_1475,N_837);
and U3148 (N_3148,N_2608,N_2526);
nor U3149 (N_3149,N_590,N_3015);
nand U3150 (N_3150,N_2750,N_951);
xnor U3151 (N_3151,N_1749,N_197);
and U3152 (N_3152,N_1756,N_1869);
or U3153 (N_3153,N_3072,N_1916);
nand U3154 (N_3154,N_983,N_1202);
or U3155 (N_3155,N_417,N_528);
or U3156 (N_3156,N_1529,N_2330);
xnor U3157 (N_3157,N_792,N_3095);
or U3158 (N_3158,N_2351,N_34);
nand U3159 (N_3159,N_923,N_2424);
nand U3160 (N_3160,N_1021,N_1705);
or U3161 (N_3161,N_299,N_806);
and U3162 (N_3162,N_2660,N_3044);
and U3163 (N_3163,N_1949,N_2679);
nor U3164 (N_3164,N_2206,N_1124);
xor U3165 (N_3165,N_1205,N_2107);
nor U3166 (N_3166,N_2126,N_356);
and U3167 (N_3167,N_1953,N_1759);
nor U3168 (N_3168,N_1097,N_3046);
and U3169 (N_3169,N_503,N_1308);
or U3170 (N_3170,N_2383,N_2117);
nand U3171 (N_3171,N_2493,N_244);
nand U3172 (N_3172,N_1977,N_1209);
or U3173 (N_3173,N_2406,N_2101);
xnor U3174 (N_3174,N_3052,N_782);
nand U3175 (N_3175,N_1426,N_28);
or U3176 (N_3176,N_2458,N_611);
nor U3177 (N_3177,N_910,N_727);
and U3178 (N_3178,N_2775,N_2063);
nand U3179 (N_3179,N_950,N_756);
or U3180 (N_3180,N_454,N_1249);
or U3181 (N_3181,N_2354,N_1416);
nor U3182 (N_3182,N_2721,N_2053);
nor U3183 (N_3183,N_3063,N_2389);
xor U3184 (N_3184,N_1626,N_483);
xor U3185 (N_3185,N_2680,N_1336);
xor U3186 (N_3186,N_95,N_3023);
and U3187 (N_3187,N_831,N_2964);
nor U3188 (N_3188,N_2990,N_1736);
xor U3189 (N_3189,N_2599,N_823);
or U3190 (N_3190,N_2257,N_388);
xnor U3191 (N_3191,N_330,N_896);
nor U3192 (N_3192,N_859,N_418);
nor U3193 (N_3193,N_1261,N_1991);
nor U3194 (N_3194,N_2636,N_1240);
or U3195 (N_3195,N_2306,N_1403);
xnor U3196 (N_3196,N_1398,N_2386);
xor U3197 (N_3197,N_661,N_2629);
nand U3198 (N_3198,N_2637,N_937);
or U3199 (N_3199,N_317,N_1604);
or U3200 (N_3200,N_2357,N_1753);
nand U3201 (N_3201,N_2859,N_434);
nor U3202 (N_3202,N_1879,N_1627);
nand U3203 (N_3203,N_628,N_305);
nand U3204 (N_3204,N_2429,N_1958);
nor U3205 (N_3205,N_1796,N_2145);
nor U3206 (N_3206,N_1046,N_599);
nor U3207 (N_3207,N_788,N_1052);
or U3208 (N_3208,N_326,N_1588);
or U3209 (N_3209,N_1065,N_3014);
nor U3210 (N_3210,N_790,N_2308);
or U3211 (N_3211,N_382,N_3069);
xnor U3212 (N_3212,N_2044,N_646);
xor U3213 (N_3213,N_1142,N_2326);
xnor U3214 (N_3214,N_193,N_1427);
xnor U3215 (N_3215,N_137,N_2006);
and U3216 (N_3216,N_1044,N_2192);
nor U3217 (N_3217,N_233,N_280);
nand U3218 (N_3218,N_1113,N_2555);
and U3219 (N_3219,N_966,N_3080);
or U3220 (N_3220,N_2209,N_1174);
xnor U3221 (N_3221,N_164,N_345);
and U3222 (N_3222,N_1488,N_1809);
nand U3223 (N_3223,N_999,N_996);
xnor U3224 (N_3224,N_2180,N_2774);
or U3225 (N_3225,N_2633,N_672);
or U3226 (N_3226,N_2800,N_1973);
and U3227 (N_3227,N_2029,N_439);
and U3228 (N_3228,N_436,N_2199);
xnor U3229 (N_3229,N_1368,N_2512);
or U3230 (N_3230,N_970,N_332);
or U3231 (N_3231,N_460,N_2319);
nor U3232 (N_3232,N_517,N_2723);
and U3233 (N_3233,N_1284,N_173);
and U3234 (N_3234,N_1467,N_2157);
nand U3235 (N_3235,N_798,N_726);
and U3236 (N_3236,N_1171,N_1275);
or U3237 (N_3237,N_1066,N_625);
nor U3238 (N_3238,N_1301,N_1771);
nand U3239 (N_3239,N_2503,N_1792);
nor U3240 (N_3240,N_1628,N_1540);
or U3241 (N_3241,N_2656,N_720);
xnor U3242 (N_3242,N_53,N_2001);
or U3243 (N_3243,N_922,N_2065);
xnor U3244 (N_3244,N_1312,N_1419);
xnor U3245 (N_3245,N_2384,N_1439);
and U3246 (N_3246,N_2097,N_1913);
and U3247 (N_3247,N_2294,N_1175);
or U3248 (N_3248,N_1876,N_2953);
or U3249 (N_3249,N_290,N_2348);
nor U3250 (N_3250,N_592,N_1645);
nand U3251 (N_3251,N_2355,N_493);
and U3252 (N_3252,N_1180,N_1712);
and U3253 (N_3253,N_2104,N_725);
nand U3254 (N_3254,N_819,N_139);
and U3255 (N_3255,N_50,N_100);
xnor U3256 (N_3256,N_1048,N_684);
xnor U3257 (N_3257,N_1373,N_2609);
nor U3258 (N_3258,N_550,N_72);
nand U3259 (N_3259,N_323,N_3031);
and U3260 (N_3260,N_698,N_2233);
or U3261 (N_3261,N_2332,N_1232);
xor U3262 (N_3262,N_1817,N_1423);
nor U3263 (N_3263,N_926,N_1435);
and U3264 (N_3264,N_2795,N_2034);
or U3265 (N_3265,N_2899,N_1482);
nor U3266 (N_3266,N_1463,N_1994);
nor U3267 (N_3267,N_1120,N_67);
nand U3268 (N_3268,N_424,N_1178);
nand U3269 (N_3269,N_433,N_1964);
nor U3270 (N_3270,N_1888,N_2431);
and U3271 (N_3271,N_351,N_3076);
and U3272 (N_3272,N_747,N_731);
nor U3273 (N_3273,N_2338,N_3100);
nor U3274 (N_3274,N_2780,N_1459);
nand U3275 (N_3275,N_3013,N_2604);
nand U3276 (N_3276,N_654,N_201);
or U3277 (N_3277,N_574,N_4);
nor U3278 (N_3278,N_1279,N_1877);
nor U3279 (N_3279,N_88,N_2122);
or U3280 (N_3280,N_845,N_3042);
nand U3281 (N_3281,N_1606,N_732);
nand U3282 (N_3282,N_1624,N_2709);
and U3283 (N_3283,N_2646,N_1354);
xor U3284 (N_3284,N_2946,N_2268);
nor U3285 (N_3285,N_1512,N_1170);
nor U3286 (N_3286,N_3005,N_2222);
and U3287 (N_3287,N_3039,N_1236);
or U3288 (N_3288,N_711,N_1609);
and U3289 (N_3289,N_2418,N_1874);
nor U3290 (N_3290,N_2048,N_652);
xnor U3291 (N_3291,N_1377,N_1560);
xnor U3292 (N_3292,N_615,N_2753);
nor U3293 (N_3293,N_513,N_1496);
xor U3294 (N_3294,N_568,N_512);
or U3295 (N_3295,N_2261,N_2339);
or U3296 (N_3296,N_254,N_1852);
nand U3297 (N_3297,N_2094,N_1479);
and U3298 (N_3298,N_2987,N_2533);
or U3299 (N_3299,N_3048,N_3006);
and U3300 (N_3300,N_2369,N_2520);
or U3301 (N_3301,N_96,N_659);
nor U3302 (N_3302,N_355,N_1686);
nor U3303 (N_3303,N_1598,N_631);
xnor U3304 (N_3304,N_1060,N_600);
xor U3305 (N_3305,N_587,N_214);
and U3306 (N_3306,N_1914,N_765);
and U3307 (N_3307,N_1032,N_1824);
nor U3308 (N_3308,N_269,N_357);
and U3309 (N_3309,N_364,N_2398);
and U3310 (N_3310,N_2405,N_1378);
xnor U3311 (N_3311,N_2361,N_2620);
and U3312 (N_3312,N_130,N_2475);
and U3313 (N_3313,N_3074,N_716);
or U3314 (N_3314,N_2616,N_256);
nor U3315 (N_3315,N_2289,N_441);
xnor U3316 (N_3316,N_1417,N_195);
and U3317 (N_3317,N_1214,N_1611);
xor U3318 (N_3318,N_2364,N_561);
nand U3319 (N_3319,N_2494,N_2876);
xor U3320 (N_3320,N_36,N_2744);
or U3321 (N_3321,N_2639,N_2208);
nor U3322 (N_3322,N_1745,N_110);
or U3323 (N_3323,N_533,N_1658);
nor U3324 (N_3324,N_1025,N_307);
xnor U3325 (N_3325,N_1960,N_127);
and U3326 (N_3326,N_48,N_1890);
nor U3327 (N_3327,N_2849,N_1873);
nor U3328 (N_3328,N_2021,N_1151);
nand U3329 (N_3329,N_147,N_1962);
or U3330 (N_3330,N_986,N_300);
xnor U3331 (N_3331,N_66,N_1451);
xor U3332 (N_3332,N_653,N_331);
and U3333 (N_3333,N_1704,N_2352);
and U3334 (N_3334,N_1726,N_2854);
and U3335 (N_3335,N_2070,N_2948);
or U3336 (N_3336,N_224,N_2223);
xnor U3337 (N_3337,N_1440,N_2396);
nor U3338 (N_3338,N_810,N_1592);
and U3339 (N_3339,N_1525,N_3117);
nand U3340 (N_3340,N_2393,N_2264);
xor U3341 (N_3341,N_3124,N_828);
xnor U3342 (N_3342,N_1149,N_1267);
nand U3343 (N_3343,N_1667,N_1896);
or U3344 (N_3344,N_1564,N_1096);
nand U3345 (N_3345,N_609,N_2360);
and U3346 (N_3346,N_912,N_1901);
nand U3347 (N_3347,N_1057,N_212);
nand U3348 (N_3348,N_1028,N_1589);
or U3349 (N_3349,N_2856,N_1402);
and U3350 (N_3350,N_745,N_880);
and U3351 (N_3351,N_2936,N_1179);
nor U3352 (N_3352,N_2747,N_2543);
xor U3353 (N_3353,N_722,N_643);
nor U3354 (N_3354,N_2671,N_1310);
nor U3355 (N_3355,N_2941,N_2920);
or U3356 (N_3356,N_1760,N_2853);
and U3357 (N_3357,N_1442,N_2079);
nand U3358 (N_3358,N_2500,N_316);
xor U3359 (N_3359,N_2698,N_302);
nor U3360 (N_3360,N_835,N_3079);
xnor U3361 (N_3361,N_1775,N_2413);
nor U3362 (N_3362,N_404,N_2219);
or U3363 (N_3363,N_2614,N_1989);
xnor U3364 (N_3364,N_1734,N_1872);
nand U3365 (N_3365,N_2293,N_2752);
or U3366 (N_3366,N_759,N_1296);
nor U3367 (N_3367,N_2672,N_1905);
xnor U3368 (N_3368,N_981,N_2562);
or U3369 (N_3369,N_1729,N_2505);
and U3370 (N_3370,N_2976,N_2090);
or U3371 (N_3371,N_1965,N_0);
nand U3372 (N_3372,N_1251,N_2630);
xor U3373 (N_3373,N_850,N_1250);
or U3374 (N_3374,N_113,N_2365);
nor U3375 (N_3375,N_1685,N_2687);
xnor U3376 (N_3376,N_2912,N_2557);
or U3377 (N_3377,N_2486,N_1383);
xor U3378 (N_3378,N_1811,N_635);
and U3379 (N_3379,N_1750,N_2613);
xnor U3380 (N_3380,N_7,N_967);
or U3381 (N_3381,N_1707,N_669);
nor U3382 (N_3382,N_236,N_642);
and U3383 (N_3383,N_2880,N_1432);
or U3384 (N_3384,N_2971,N_40);
nor U3385 (N_3385,N_2595,N_2915);
nand U3386 (N_3386,N_3121,N_1349);
and U3387 (N_3387,N_516,N_2404);
and U3388 (N_3388,N_2563,N_2855);
and U3389 (N_3389,N_1342,N_717);
nand U3390 (N_3390,N_2965,N_1531);
nor U3391 (N_3391,N_1182,N_1298);
xor U3392 (N_3392,N_1246,N_809);
nor U3393 (N_3393,N_1022,N_2080);
and U3394 (N_3394,N_1614,N_472);
or U3395 (N_3395,N_2316,N_686);
or U3396 (N_3396,N_2865,N_1480);
and U3397 (N_3397,N_774,N_2565);
xnor U3398 (N_3398,N_723,N_1992);
or U3399 (N_3399,N_1072,N_3065);
or U3400 (N_3400,N_1927,N_2213);
nor U3401 (N_3401,N_821,N_566);
or U3402 (N_3402,N_151,N_1744);
xnor U3403 (N_3403,N_1146,N_1562);
or U3404 (N_3404,N_3009,N_1735);
xnor U3405 (N_3405,N_2519,N_977);
and U3406 (N_3406,N_1505,N_1150);
nor U3407 (N_3407,N_1866,N_1754);
nor U3408 (N_3408,N_2216,N_279);
or U3409 (N_3409,N_415,N_3081);
or U3410 (N_3410,N_2110,N_183);
and U3411 (N_3411,N_2764,N_862);
xnor U3412 (N_3412,N_1630,N_2755);
and U3413 (N_3413,N_350,N_2066);
nand U3414 (N_3414,N_1469,N_797);
nand U3415 (N_3415,N_2881,N_2727);
or U3416 (N_3416,N_2975,N_873);
xnor U3417 (N_3417,N_2454,N_3024);
or U3418 (N_3418,N_1216,N_1619);
or U3419 (N_3419,N_25,N_1011);
nor U3420 (N_3420,N_1774,N_2939);
nand U3421 (N_3421,N_1217,N_2716);
nor U3422 (N_3422,N_243,N_2521);
nor U3423 (N_3423,N_584,N_2017);
xnor U3424 (N_3424,N_2334,N_2191);
or U3425 (N_3425,N_2682,N_1823);
and U3426 (N_3426,N_499,N_1311);
nand U3427 (N_3427,N_2333,N_1095);
or U3428 (N_3428,N_2183,N_239);
xor U3429 (N_3429,N_2835,N_249);
or U3430 (N_3430,N_2872,N_1652);
xnor U3431 (N_3431,N_2974,N_268);
xnor U3432 (N_3432,N_2906,N_2414);
or U3433 (N_3433,N_2367,N_1389);
nor U3434 (N_3434,N_480,N_2897);
xnor U3435 (N_3435,N_1790,N_2678);
and U3436 (N_3436,N_361,N_2564);
or U3437 (N_3437,N_31,N_2045);
and U3438 (N_3438,N_1574,N_1909);
and U3439 (N_3439,N_468,N_1381);
and U3440 (N_3440,N_706,N_275);
nand U3441 (N_3441,N_2449,N_1094);
xor U3442 (N_3442,N_1671,N_1137);
xnor U3443 (N_3443,N_1003,N_283);
or U3444 (N_3444,N_1701,N_902);
or U3445 (N_3445,N_210,N_2258);
and U3446 (N_3446,N_1330,N_2701);
xor U3447 (N_3447,N_2020,N_282);
xnor U3448 (N_3448,N_1986,N_2194);
xnor U3449 (N_3449,N_1408,N_3116);
nand U3450 (N_3450,N_2415,N_395);
or U3451 (N_3451,N_2697,N_1815);
and U3452 (N_3452,N_1600,N_389);
nand U3453 (N_3453,N_2155,N_734);
or U3454 (N_3454,N_1347,N_817);
nand U3455 (N_3455,N_1010,N_108);
nand U3456 (N_3456,N_106,N_198);
and U3457 (N_3457,N_2700,N_2088);
nand U3458 (N_3458,N_1444,N_2978);
and U3459 (N_3459,N_89,N_250);
nor U3460 (N_3460,N_1450,N_459);
nor U3461 (N_3461,N_980,N_527);
xnor U3462 (N_3462,N_231,N_1421);
nand U3463 (N_3463,N_907,N_2497);
nor U3464 (N_3464,N_636,N_504);
nand U3465 (N_3465,N_2551,N_2811);
or U3466 (N_3466,N_2438,N_2981);
nor U3467 (N_3467,N_2814,N_2287);
or U3468 (N_3468,N_2204,N_2824);
and U3469 (N_3469,N_1407,N_960);
nor U3470 (N_3470,N_227,N_1518);
or U3471 (N_3471,N_1218,N_2274);
xor U3472 (N_3472,N_963,N_2955);
and U3473 (N_3473,N_1101,N_547);
and U3474 (N_3474,N_1608,N_1737);
or U3475 (N_3475,N_2411,N_2507);
nor U3476 (N_3476,N_5,N_1264);
nor U3477 (N_3477,N_2304,N_1623);
nand U3478 (N_3478,N_733,N_1242);
or U3479 (N_3479,N_1002,N_1007);
and U3480 (N_3480,N_857,N_2498);
nor U3481 (N_3481,N_163,N_2461);
xor U3482 (N_3482,N_1037,N_973);
or U3483 (N_3483,N_1086,N_2492);
nand U3484 (N_3484,N_1761,N_453);
nand U3485 (N_3485,N_2282,N_1268);
or U3486 (N_3486,N_914,N_2628);
and U3487 (N_3487,N_3032,N_1920);
and U3488 (N_3488,N_1014,N_1537);
xnor U3489 (N_3489,N_2696,N_1243);
nand U3490 (N_3490,N_800,N_2980);
xor U3491 (N_3491,N_1689,N_1618);
nor U3492 (N_3492,N_2127,N_1228);
nand U3493 (N_3493,N_3112,N_23);
or U3494 (N_3494,N_602,N_948);
and U3495 (N_3495,N_832,N_1290);
or U3496 (N_3496,N_1078,N_2465);
or U3497 (N_3497,N_2158,N_1680);
nor U3498 (N_3498,N_868,N_779);
nand U3499 (N_3499,N_252,N_2035);
xor U3500 (N_3500,N_690,N_1231);
xnor U3501 (N_3501,N_577,N_1023);
nor U3502 (N_3502,N_1320,N_2342);
or U3503 (N_3503,N_730,N_2647);
or U3504 (N_3504,N_20,N_346);
nor U3505 (N_3505,N_1001,N_773);
or U3506 (N_3506,N_1184,N_487);
or U3507 (N_3507,N_715,N_2002);
nand U3508 (N_3508,N_1083,N_2436);
xnor U3509 (N_3509,N_1302,N_1271);
and U3510 (N_3510,N_1176,N_1546);
nand U3511 (N_3511,N_1341,N_2247);
nand U3512 (N_3512,N_2069,N_400);
and U3513 (N_3513,N_1514,N_709);
nor U3514 (N_3514,N_2713,N_2568);
and U3515 (N_3515,N_1081,N_338);
and U3516 (N_3516,N_1840,N_1816);
and U3517 (N_3517,N_1321,N_860);
nor U3518 (N_3518,N_429,N_419);
xor U3519 (N_3519,N_2082,N_372);
and U3520 (N_3520,N_2518,N_1845);
and U3521 (N_3521,N_2238,N_2171);
nor U3522 (N_3522,N_883,N_2772);
xor U3523 (N_3523,N_2392,N_1340);
xnor U3524 (N_3524,N_2745,N_2025);
nand U3525 (N_3525,N_2770,N_2068);
nand U3526 (N_3526,N_656,N_1979);
or U3527 (N_3527,N_2453,N_585);
and U3528 (N_3528,N_3059,N_2799);
or U3529 (N_3529,N_396,N_2490);
xor U3530 (N_3530,N_2092,N_2908);
nor U3531 (N_3531,N_3034,N_2786);
and U3532 (N_3532,N_2592,N_248);
xor U3533 (N_3533,N_1262,N_1702);
nand U3534 (N_3534,N_976,N_2560);
or U3535 (N_3535,N_2462,N_278);
and U3536 (N_3536,N_1187,N_1122);
and U3537 (N_3537,N_211,N_1798);
and U3538 (N_3538,N_1720,N_749);
xnor U3539 (N_3539,N_905,N_184);
and U3540 (N_3540,N_2150,N_2485);
nor U3541 (N_3541,N_766,N_81);
and U3542 (N_3542,N_1212,N_328);
or U3543 (N_3543,N_1413,N_3088);
nor U3544 (N_3544,N_2007,N_750);
nand U3545 (N_3545,N_3050,N_1303);
or U3546 (N_3546,N_1476,N_2504);
and U3547 (N_3547,N_703,N_1105);
and U3548 (N_3548,N_549,N_442);
xnor U3549 (N_3549,N_755,N_2726);
or U3550 (N_3550,N_257,N_1473);
nand U3551 (N_3551,N_2483,N_2181);
nand U3552 (N_3552,N_576,N_161);
xor U3553 (N_3553,N_1177,N_1506);
nand U3554 (N_3554,N_721,N_2154);
or U3555 (N_3555,N_911,N_2100);
nor U3556 (N_3556,N_2036,N_241);
xnor U3557 (N_3557,N_1152,N_370);
and U3558 (N_3558,N_1846,N_1682);
or U3559 (N_3559,N_1213,N_2010);
nor U3560 (N_3560,N_55,N_526);
and U3561 (N_3561,N_1523,N_1358);
nor U3562 (N_3562,N_2582,N_2930);
and U3563 (N_3563,N_2889,N_802);
xnor U3564 (N_3564,N_87,N_3030);
nor U3565 (N_3565,N_2000,N_990);
and U3566 (N_3566,N_553,N_928);
and U3567 (N_3567,N_2026,N_1791);
nor U3568 (N_3568,N_222,N_141);
and U3569 (N_3569,N_1038,N_1056);
and U3570 (N_3570,N_1332,N_1053);
nor U3571 (N_3571,N_1309,N_1715);
and U3572 (N_3572,N_1462,N_1887);
nand U3573 (N_3573,N_2846,N_2862);
nand U3574 (N_3574,N_482,N_1145);
nor U3575 (N_3575,N_2816,N_674);
xor U3576 (N_3576,N_1577,N_1392);
or U3577 (N_3577,N_1665,N_534);
nand U3578 (N_3578,N_2241,N_440);
or U3579 (N_3579,N_125,N_1996);
xor U3580 (N_3580,N_1533,N_1693);
and U3581 (N_3581,N_1632,N_1333);
nand U3582 (N_3582,N_123,N_3083);
nor U3583 (N_3583,N_1859,N_743);
or U3584 (N_3584,N_2200,N_2240);
and U3585 (N_3585,N_154,N_1895);
nor U3586 (N_3586,N_1721,N_607);
nand U3587 (N_3587,N_1254,N_724);
xnor U3588 (N_3588,N_3038,N_955);
nand U3589 (N_3589,N_2165,N_3007);
xnor U3590 (N_3590,N_942,N_1654);
xnor U3591 (N_3591,N_741,N_872);
nor U3592 (N_3592,N_3106,N_2923);
and U3593 (N_3593,N_3091,N_2969);
and U3594 (N_3594,N_995,N_645);
and U3595 (N_3595,N_461,N_2347);
xor U3596 (N_3596,N_1445,N_1538);
nor U3597 (N_3597,N_2642,N_2435);
xnor U3598 (N_3598,N_2535,N_109);
nand U3599 (N_3599,N_1,N_701);
nand U3600 (N_3600,N_890,N_488);
and U3601 (N_3601,N_748,N_801);
xor U3602 (N_3602,N_2731,N_2631);
xor U3603 (N_3603,N_551,N_1870);
nor U3604 (N_3604,N_152,N_1993);
xor U3605 (N_3605,N_1112,N_2708);
nor U3606 (N_3606,N_699,N_245);
and U3607 (N_3607,N_1329,N_1728);
nor U3608 (N_3608,N_918,N_443);
and U3609 (N_3609,N_770,N_298);
xor U3610 (N_3610,N_2138,N_2099);
and U3611 (N_3611,N_2464,N_247);
xor U3612 (N_3612,N_2916,N_1783);
nand U3613 (N_3613,N_2997,N_1765);
nand U3614 (N_3614,N_466,N_2922);
and U3615 (N_3615,N_920,N_2894);
or U3616 (N_3616,N_2186,N_2224);
or U3617 (N_3617,N_2087,N_1711);
nand U3618 (N_3618,N_1222,N_2221);
or U3619 (N_3619,N_1270,N_56);
nor U3620 (N_3620,N_2172,N_2940);
nor U3621 (N_3621,N_1675,N_47);
xnor U3622 (N_3622,N_3040,N_1568);
and U3623 (N_3623,N_2423,N_2265);
and U3624 (N_3624,N_2106,N_728);
or U3625 (N_3625,N_1834,N_1637);
nor U3626 (N_3626,N_781,N_2506);
nand U3627 (N_3627,N_2979,N_386);
and U3628 (N_3628,N_1567,N_3084);
nand U3629 (N_3629,N_662,N_402);
and U3630 (N_3630,N_511,N_1984);
xnor U3631 (N_3631,N_2491,N_2479);
xor U3632 (N_3632,N_1018,N_988);
and U3633 (N_3633,N_458,N_2720);
nor U3634 (N_3634,N_2902,N_2318);
or U3635 (N_3635,N_1773,N_1304);
xnor U3636 (N_3636,N_359,N_29);
nor U3637 (N_3637,N_1510,N_2376);
xor U3638 (N_3638,N_2668,N_3123);
and U3639 (N_3639,N_1288,N_2686);
nor U3640 (N_3640,N_105,N_2866);
and U3641 (N_3641,N_144,N_1638);
and U3642 (N_3642,N_559,N_446);
xnor U3643 (N_3643,N_1069,N_1944);
or U3644 (N_3644,N_1795,N_2302);
nor U3645 (N_3645,N_1902,N_2201);
or U3646 (N_3646,N_391,N_463);
and U3647 (N_3647,N_2481,N_1234);
xnor U3648 (N_3648,N_495,N_1364);
and U3649 (N_3649,N_3061,N_1945);
and U3650 (N_3650,N_2416,N_70);
and U3651 (N_3651,N_1943,N_1189);
xor U3652 (N_3652,N_1844,N_381);
or U3653 (N_3653,N_159,N_1324);
or U3654 (N_3654,N_589,N_2779);
nand U3655 (N_3655,N_41,N_1397);
xor U3656 (N_3656,N_579,N_921);
or U3657 (N_3657,N_1800,N_1013);
xnor U3658 (N_3658,N_2681,N_2561);
nor U3659 (N_3659,N_941,N_1253);
xnor U3660 (N_3660,N_1248,N_327);
nand U3661 (N_3661,N_1148,N_1485);
and U3662 (N_3662,N_2607,N_2252);
nand U3663 (N_3663,N_1135,N_761);
and U3664 (N_3664,N_1957,N_1858);
nor U3665 (N_3665,N_2315,N_1516);
nand U3666 (N_3666,N_2918,N_2422);
or U3667 (N_3667,N_836,N_2826);
or U3668 (N_3668,N_882,N_2470);
or U3669 (N_3669,N_2892,N_1700);
nor U3670 (N_3670,N_620,N_2243);
xor U3671 (N_3671,N_491,N_2903);
or U3672 (N_3672,N_1807,N_2050);
and U3673 (N_3673,N_1061,N_537);
xor U3674 (N_3674,N_2489,N_24);
and U3675 (N_3675,N_1836,N_901);
or U3676 (N_3676,N_2659,N_2133);
nand U3677 (N_3677,N_2790,N_1871);
and U3678 (N_3678,N_2711,N_1280);
or U3679 (N_3679,N_1495,N_2719);
or U3680 (N_3680,N_2657,N_444);
xnor U3681 (N_3681,N_405,N_1323);
nand U3682 (N_3682,N_2016,N_1117);
nand U3683 (N_3683,N_1139,N_2129);
or U3684 (N_3684,N_785,N_2689);
and U3685 (N_3685,N_2801,N_2959);
or U3686 (N_3686,N_94,N_1143);
or U3687 (N_3687,N_841,N_1613);
nand U3688 (N_3688,N_189,N_496);
or U3689 (N_3689,N_1183,N_1483);
nor U3690 (N_3690,N_2484,N_438);
xnor U3691 (N_3691,N_1710,N_854);
and U3692 (N_3692,N_3110,N_1880);
xnor U3693 (N_3693,N_2381,N_663);
nor U3694 (N_3694,N_2860,N_1797);
nor U3695 (N_3695,N_2949,N_2942);
xnor U3696 (N_3696,N_3033,N_2717);
xor U3697 (N_3697,N_2634,N_1239);
xor U3698 (N_3698,N_1504,N_267);
and U3699 (N_3699,N_1043,N_2928);
and U3700 (N_3700,N_2197,N_612);
or U3701 (N_3701,N_1857,N_2541);
or U3702 (N_3702,N_1351,N_895);
and U3703 (N_3703,N_1699,N_2291);
and U3704 (N_3704,N_2402,N_194);
nand U3705 (N_3705,N_1741,N_1899);
xor U3706 (N_3706,N_1952,N_919);
nor U3707 (N_3707,N_1757,N_18);
and U3708 (N_3708,N_2322,N_936);
or U3709 (N_3709,N_1636,N_2960);
or U3710 (N_3710,N_946,N_560);
nand U3711 (N_3711,N_502,N_1557);
nor U3712 (N_3712,N_3049,N_2580);
nand U3713 (N_3713,N_1125,N_1738);
and U3714 (N_3714,N_2421,N_170);
and U3715 (N_3715,N_1532,N_1946);
or U3716 (N_3716,N_1694,N_2808);
nand U3717 (N_3717,N_1515,N_1983);
nand U3718 (N_3718,N_2451,N_510);
and U3719 (N_3719,N_1379,N_2993);
or U3720 (N_3720,N_2870,N_2195);
nor U3721 (N_3721,N_2175,N_2182);
nor U3722 (N_3722,N_2589,N_1237);
or U3723 (N_3723,N_1580,N_1535);
and U3724 (N_3724,N_719,N_1851);
and U3725 (N_3725,N_2913,N_1141);
and U3726 (N_3726,N_215,N_1063);
xor U3727 (N_3727,N_2280,N_2733);
and U3728 (N_3728,N_695,N_1306);
and U3729 (N_3729,N_1612,N_2954);
and U3730 (N_3730,N_1255,N_522);
nand U3731 (N_3731,N_1036,N_2119);
nor U3732 (N_3732,N_1576,N_3075);
or U3733 (N_3733,N_2588,N_536);
and U3734 (N_3734,N_2227,N_2886);
nand U3735 (N_3735,N_1969,N_2995);
or U3736 (N_3736,N_1315,N_1362);
and U3737 (N_3737,N_2741,N_2729);
or U3738 (N_3738,N_1159,N_2809);
and U3739 (N_3739,N_1541,N_2810);
or U3740 (N_3740,N_1447,N_2730);
nor U3741 (N_3741,N_1555,N_1825);
or U3742 (N_3742,N_2651,N_1227);
nor U3743 (N_3743,N_2879,N_1892);
nor U3744 (N_3744,N_190,N_689);
and U3745 (N_3745,N_153,N_432);
nor U3746 (N_3746,N_641,N_1465);
nand U3747 (N_3747,N_3035,N_626);
nand U3748 (N_3748,N_44,N_1646);
or U3749 (N_3749,N_751,N_2513);
nand U3750 (N_3750,N_2300,N_232);
nor U3751 (N_3751,N_886,N_1855);
nor U3752 (N_3752,N_2362,N_2473);
and U3753 (N_3753,N_76,N_3068);
xor U3754 (N_3754,N_1291,N_1733);
or U3755 (N_3755,N_411,N_2917);
nor U3756 (N_3756,N_259,N_112);
xnor U3757 (N_3757,N_515,N_1590);
nand U3758 (N_3758,N_408,N_729);
or U3759 (N_3759,N_341,N_827);
and U3760 (N_3760,N_2275,N_486);
nor U3761 (N_3761,N_2650,N_220);
nor U3762 (N_3762,N_1883,N_897);
and U3763 (N_3763,N_1067,N_1106);
or U3764 (N_3764,N_2188,N_713);
and U3765 (N_3765,N_1679,N_145);
or U3766 (N_3766,N_804,N_898);
nor U3767 (N_3767,N_1719,N_1530);
or U3768 (N_3768,N_3018,N_971);
or U3769 (N_3769,N_2324,N_1752);
and U3770 (N_3770,N_2353,N_1104);
xnor U3771 (N_3771,N_1838,N_1644);
xor U3772 (N_3772,N_312,N_272);
or U3773 (N_3773,N_2911,N_258);
and U3774 (N_3774,N_3012,N_2426);
nand U3775 (N_3775,N_2067,N_1670);
or U3776 (N_3776,N_3017,N_1829);
and U3777 (N_3777,N_1875,N_583);
xor U3778 (N_3778,N_2356,N_565);
nor U3779 (N_3779,N_893,N_1691);
nor U3780 (N_3780,N_2228,N_3029);
or U3781 (N_3781,N_1668,N_2895);
xnor U3782 (N_3782,N_33,N_1625);
nand U3783 (N_3783,N_1115,N_867);
xnor U3784 (N_3784,N_2214,N_799);
or U3785 (N_3785,N_1956,N_778);
and U3786 (N_3786,N_712,N_1770);
and U3787 (N_3787,N_1307,N_465);
nor U3788 (N_3788,N_1410,N_2130);
nand U3789 (N_3789,N_2317,N_2662);
nor U3790 (N_3790,N_2480,N_1258);
nand U3791 (N_3791,N_2921,N_1110);
nand U3792 (N_3792,N_1746,N_2412);
nor U3793 (N_3793,N_398,N_2784);
nor U3794 (N_3794,N_879,N_1903);
and U3795 (N_3795,N_64,N_2705);
nand U3796 (N_3796,N_2788,N_696);
nand U3797 (N_3797,N_2297,N_876);
nand U3798 (N_3798,N_2239,N_532);
nand U3799 (N_3799,N_148,N_2245);
and U3800 (N_3800,N_915,N_610);
and U3801 (N_3801,N_2757,N_2743);
or U3802 (N_3802,N_399,N_1490);
nor U3803 (N_3803,N_1204,N_2255);
and U3804 (N_3804,N_451,N_1316);
nor U3805 (N_3805,N_586,N_1804);
or U3806 (N_3806,N_1343,N_758);
or U3807 (N_3807,N_26,N_264);
xnor U3808 (N_3808,N_614,N_234);
nor U3809 (N_3809,N_2648,N_2673);
or U3810 (N_3810,N_1015,N_2832);
nor U3811 (N_3811,N_3096,N_944);
xnor U3812 (N_3812,N_2852,N_938);
xor U3813 (N_3813,N_348,N_2537);
or U3814 (N_3814,N_899,N_3064);
and U3815 (N_3815,N_667,N_1446);
and U3816 (N_3816,N_2724,N_849);
nand U3817 (N_3817,N_114,N_3105);
or U3818 (N_3818,N_111,N_61);
xor U3819 (N_3819,N_2804,N_2009);
nor U3820 (N_3820,N_1367,N_2618);
xor U3821 (N_3821,N_2896,N_908);
nor U3822 (N_3822,N_3016,N_474);
nor U3823 (N_3823,N_2621,N_455);
xor U3824 (N_3824,N_851,N_2591);
xnor U3825 (N_3825,N_2166,N_2690);
nand U3826 (N_3826,N_2468,N_2083);
nor U3827 (N_3827,N_251,N_1454);
nor U3828 (N_3828,N_2692,N_1223);
nand U3829 (N_3829,N_737,N_1327);
nand U3830 (N_3830,N_767,N_925);
nand U3831 (N_3831,N_2973,N_2598);
nor U3832 (N_3832,N_1633,N_492);
nor U3833 (N_3833,N_2298,N_2212);
xor U3834 (N_3834,N_309,N_2843);
or U3835 (N_3835,N_714,N_1128);
or U3836 (N_3836,N_2556,N_2336);
nor U3837 (N_3837,N_2242,N_301);
nand U3838 (N_3838,N_2225,N_853);
nand U3839 (N_3839,N_2161,N_376);
and U3840 (N_3840,N_2057,N_1325);
xnor U3841 (N_3841,N_556,N_1764);
or U3842 (N_3842,N_51,N_1908);
xor U3843 (N_3843,N_368,N_1990);
xnor U3844 (N_3844,N_575,N_422);
nor U3845 (N_3845,N_1660,N_2536);
xnor U3846 (N_3846,N_2910,N_1513);
and U3847 (N_3847,N_606,N_2441);
nand U3848 (N_3848,N_818,N_1192);
xnor U3849 (N_3849,N_1556,N_1810);
nor U3850 (N_3850,N_1108,N_296);
nor U3851 (N_3851,N_322,N_2781);
or U3852 (N_3852,N_2602,N_2830);
and U3853 (N_3853,N_1157,N_1334);
or U3854 (N_3854,N_1027,N_2267);
nand U3855 (N_3855,N_1907,N_1587);
xnor U3856 (N_3856,N_3058,N_2198);
xor U3857 (N_3857,N_1528,N_2296);
or U3858 (N_3858,N_128,N_1486);
or U3859 (N_3859,N_1164,N_1639);
or U3860 (N_3860,N_1452,N_2901);
and U3861 (N_3861,N_762,N_627);
and U3862 (N_3862,N_3027,N_2447);
and U3863 (N_3863,N_1390,N_199);
or U3864 (N_3864,N_2273,N_538);
and U3865 (N_3865,N_1103,N_1864);
and U3866 (N_3866,N_2259,N_1801);
xnor U3867 (N_3867,N_702,N_739);
or U3868 (N_3868,N_2619,N_353);
and U3869 (N_3869,N_1987,N_1073);
or U3870 (N_3870,N_169,N_2164);
nor U3871 (N_3871,N_1029,N_3037);
nor U3872 (N_3872,N_1331,N_1437);
xor U3873 (N_3873,N_1400,N_1016);
and U3874 (N_3874,N_321,N_1405);
and U3875 (N_3875,N_2715,N_889);
nand U3876 (N_3876,N_863,N_855);
or U3877 (N_3877,N_2666,N_2571);
nor U3878 (N_3878,N_2340,N_2173);
or U3879 (N_3879,N_814,N_2823);
nand U3880 (N_3880,N_1534,N_593);
xor U3881 (N_3881,N_2084,N_2077);
xor U3882 (N_3882,N_1375,N_2958);
nor U3883 (N_3883,N_2478,N_1087);
xnor U3884 (N_3884,N_2900,N_2675);
xnor U3885 (N_3885,N_2807,N_2649);
and U3886 (N_3886,N_1224,N_1548);
xor U3887 (N_3887,N_52,N_1650);
nand U3888 (N_3888,N_2570,N_1140);
nor U3889 (N_3889,N_186,N_1472);
xor U3890 (N_3890,N_2395,N_2516);
xnor U3891 (N_3891,N_2754,N_2218);
nor U3892 (N_3892,N_2793,N_2115);
or U3893 (N_3893,N_1478,N_1494);
or U3894 (N_3894,N_639,N_1130);
or U3895 (N_3895,N_1585,N_473);
and U3896 (N_3896,N_213,N_2487);
or U3897 (N_3897,N_2256,N_1820);
and U3898 (N_3898,N_3001,N_752);
xor U3899 (N_3899,N_221,N_82);
xor U3900 (N_3900,N_1466,N_2550);
or U3901 (N_3901,N_43,N_2663);
or U3902 (N_3902,N_1197,N_1766);
nand U3903 (N_3903,N_693,N_1193);
and U3904 (N_3904,N_557,N_470);
or U3905 (N_3905,N_2929,N_2857);
and U3906 (N_3906,N_1780,N_660);
nand U3907 (N_3907,N_1544,N_2179);
nor U3908 (N_3908,N_134,N_428);
nand U3909 (N_3909,N_869,N_894);
and U3910 (N_3910,N_2545,N_1477);
and U3911 (N_3911,N_2888,N_2290);
and U3912 (N_3912,N_2762,N_1219);
or U3913 (N_3913,N_2135,N_1659);
or U3914 (N_3914,N_1277,N_2271);
nor U3915 (N_3915,N_2448,N_318);
nor U3916 (N_3916,N_1622,N_965);
or U3917 (N_3917,N_1226,N_423);
nand U3918 (N_3918,N_826,N_2530);
nor U3919 (N_3919,N_1155,N_1376);
xnor U3920 (N_3920,N_1318,N_464);
xnor U3921 (N_3921,N_1539,N_844);
or U3922 (N_3922,N_603,N_1191);
or U3923 (N_3923,N_2434,N_49);
nor U3924 (N_3924,N_2051,N_2796);
nand U3925 (N_3925,N_979,N_1933);
and U3926 (N_3926,N_175,N_539);
nand U3927 (N_3927,N_1006,N_578);
nand U3928 (N_3928,N_2203,N_2064);
nand U3929 (N_3929,N_2401,N_2961);
xor U3930 (N_3930,N_1841,N_17);
and U3931 (N_3931,N_3026,N_13);
xnor U3932 (N_3932,N_2907,N_847);
and U3933 (N_3933,N_2037,N_815);
nand U3934 (N_3934,N_3073,N_1569);
and U3935 (N_3935,N_288,N_2012);
or U3936 (N_3936,N_146,N_54);
nand U3937 (N_3937,N_1634,N_738);
nand U3938 (N_3938,N_379,N_1503);
or U3939 (N_3939,N_2778,N_2103);
nor U3940 (N_3940,N_1997,N_2968);
nor U3941 (N_3941,N_1319,N_45);
nand U3942 (N_3942,N_2956,N_2771);
or U3943 (N_3943,N_1930,N_840);
xnor U3944 (N_3944,N_1190,N_2061);
and U3945 (N_3945,N_3122,N_2096);
nand U3946 (N_3946,N_2457,N_1166);
xnor U3947 (N_3947,N_1456,N_742);
xnor U3948 (N_3948,N_2098,N_2163);
xnor U3949 (N_3949,N_1917,N_3019);
or U3950 (N_3950,N_2160,N_1420);
nor U3951 (N_3951,N_1910,N_2460);
nor U3952 (N_3952,N_621,N_167);
and U3953 (N_3953,N_2792,N_1365);
nor U3954 (N_3954,N_2877,N_1509);
nor U3955 (N_3955,N_1678,N_2510);
nor U3956 (N_3956,N_2883,N_2593);
or U3957 (N_3957,N_1276,N_129);
nand U3958 (N_3958,N_1511,N_2286);
and U3959 (N_3959,N_1867,N_324);
nand U3960 (N_3960,N_665,N_1578);
nor U3961 (N_3961,N_1361,N_1366);
nor U3962 (N_3962,N_1942,N_1350);
or U3963 (N_3963,N_3082,N_1273);
nor U3964 (N_3964,N_1068,N_2935);
or U3965 (N_3965,N_1664,N_1126);
nor U3966 (N_3966,N_805,N_1269);
nand U3967 (N_3967,N_1904,N_456);
nand U3968 (N_3968,N_1040,N_2307);
and U3969 (N_3969,N_12,N_1434);
or U3970 (N_3970,N_3036,N_1758);
xnor U3971 (N_3971,N_2838,N_2581);
nand U3972 (N_3972,N_1947,N_555);
and U3973 (N_3973,N_812,N_546);
or U3974 (N_3974,N_2023,N_19);
xnor U3975 (N_3975,N_462,N_2851);
nor U3976 (N_3976,N_1940,N_2499);
nand U3977 (N_3977,N_2372,N_2211);
nand U3978 (N_3978,N_1884,N_1138);
xnor U3979 (N_3979,N_1339,N_1722);
nand U3980 (N_3980,N_856,N_3078);
nor U3981 (N_3981,N_1968,N_2988);
nor U3982 (N_3982,N_3118,N_685);
or U3983 (N_3983,N_3002,N_1107);
or U3984 (N_3984,N_617,N_2529);
and U3985 (N_3985,N_1926,N_260);
nand U3986 (N_3986,N_852,N_1386);
xnor U3987 (N_3987,N_1508,N_374);
and U3988 (N_3988,N_3099,N_2176);
or U3989 (N_3989,N_1114,N_932);
or U3990 (N_3990,N_1601,N_481);
nand U3991 (N_3991,N_1821,N_412);
and U3992 (N_3992,N_972,N_1718);
or U3993 (N_3993,N_58,N_15);
or U3994 (N_3994,N_875,N_644);
and U3995 (N_3995,N_1545,N_2018);
and U3996 (N_3996,N_1163,N_1049);
nor U3997 (N_3997,N_3097,N_598);
nor U3998 (N_3998,N_242,N_2382);
or U3999 (N_3999,N_1412,N_1372);
xnor U4000 (N_4000,N_2983,N_846);
and U4001 (N_4001,N_1294,N_1071);
nor U4002 (N_4002,N_479,N_1345);
or U4003 (N_4003,N_943,N_261);
and U4004 (N_4004,N_1985,N_2403);
or U4005 (N_4005,N_187,N_315);
nor U4006 (N_4006,N_2153,N_1837);
xnor U4007 (N_4007,N_1085,N_1244);
and U4008 (N_4008,N_1136,N_757);
nand U4009 (N_4009,N_2583,N_1524);
and U4010 (N_4010,N_2237,N_2577);
and U4011 (N_4011,N_416,N_2246);
xor U4012 (N_4012,N_2718,N_1449);
or U4013 (N_4013,N_1235,N_2664);
nand U4014 (N_4014,N_935,N_1173);
xor U4015 (N_4015,N_1161,N_507);
or U4016 (N_4016,N_2278,N_2003);
and U4017 (N_4017,N_1755,N_704);
nand U4018 (N_4018,N_1596,N_2295);
or U4019 (N_4019,N_2525,N_1111);
xor U4020 (N_4020,N_2924,N_1848);
or U4021 (N_4021,N_2893,N_906);
nor U4022 (N_4022,N_2059,N_1683);
or U4023 (N_4023,N_2850,N_1769);
nand U4024 (N_4024,N_2590,N_509);
nor U4025 (N_4025,N_2982,N_178);
nor U4026 (N_4026,N_237,N_1207);
or U4027 (N_4027,N_115,N_848);
and U4028 (N_4028,N_1169,N_1129);
and U4029 (N_4029,N_2232,N_1974);
and U4030 (N_4030,N_375,N_1573);
nor U4031 (N_4031,N_3111,N_2594);
or U4032 (N_4032,N_311,N_2472);
or U4033 (N_4033,N_2054,N_2947);
xor U4034 (N_4034,N_2371,N_917);
and U4035 (N_4035,N_2626,N_142);
or U4036 (N_4036,N_2469,N_2276);
and U4037 (N_4037,N_680,N_501);
and U4038 (N_4038,N_116,N_162);
or U4039 (N_4039,N_1371,N_984);
nand U4040 (N_4040,N_447,N_1299);
nor U4041 (N_4041,N_1470,N_2124);
and U4042 (N_4042,N_1436,N_545);
and U4043 (N_4043,N_471,N_864);
nor U4044 (N_4044,N_2288,N_325);
or U4045 (N_4045,N_1831,N_354);
xor U4046 (N_4046,N_2427,N_2710);
nor U4047 (N_4047,N_1527,N_188);
nor U4048 (N_4048,N_2144,N_99);
xnor U4049 (N_4049,N_580,N_124);
and U4050 (N_4050,N_514,N_2839);
nand U4051 (N_4051,N_708,N_842);
or U4052 (N_4052,N_2013,N_101);
or U4053 (N_4053,N_1272,N_2279);
xor U4054 (N_4054,N_1674,N_1925);
xor U4055 (N_4055,N_2640,N_168);
nor U4056 (N_4056,N_1549,N_1441);
nor U4057 (N_4057,N_2610,N_1035);
nor U4058 (N_4058,N_494,N_2071);
nand U4059 (N_4059,N_1889,N_1865);
nor U4060 (N_4060,N_2742,N_90);
nand U4061 (N_4061,N_2685,N_2829);
and U4062 (N_4062,N_347,N_2235);
or U4063 (N_4063,N_3108,N_2584);
nand U4064 (N_4064,N_2539,N_235);
nand U4065 (N_4065,N_1042,N_1832);
nor U4066 (N_4066,N_956,N_102);
nor U4067 (N_4067,N_2387,N_2748);
xnor U4068 (N_4068,N_1651,N_1293);
or U4069 (N_4069,N_710,N_1118);
or U4070 (N_4070,N_1448,N_2128);
or U4071 (N_4071,N_959,N_207);
xor U4072 (N_4072,N_520,N_413);
nand U4073 (N_4073,N_21,N_2346);
nor U4074 (N_4074,N_2931,N_156);
and U4075 (N_4075,N_1024,N_85);
and U4076 (N_4076,N_3047,N_650);
xor U4077 (N_4077,N_1091,N_1401);
and U4078 (N_4078,N_2187,N_1692);
nand U4079 (N_4079,N_2345,N_2060);
xnor U4080 (N_4080,N_2652,N_705);
nor U4081 (N_4081,N_2011,N_1154);
xor U4082 (N_4082,N_2944,N_452);
nor U4083 (N_4083,N_435,N_1484);
nor U4084 (N_4084,N_1229,N_2136);
xnor U4085 (N_4085,N_885,N_2215);
nand U4086 (N_4086,N_740,N_735);
xnor U4087 (N_4087,N_1605,N_1988);
and U4088 (N_4088,N_2072,N_619);
or U4089 (N_4089,N_485,N_563);
or U4090 (N_4090,N_293,N_68);
or U4091 (N_4091,N_1430,N_1922);
xor U4092 (N_4092,N_262,N_1360);
nor U4093 (N_4093,N_2374,N_63);
nand U4094 (N_4094,N_2432,N_962);
nor U4095 (N_4095,N_490,N_2645);
or U4096 (N_4096,N_2989,N_2611);
xnor U4097 (N_4097,N_2927,N_1286);
nand U4098 (N_4098,N_816,N_813);
or U4099 (N_4099,N_1394,N_616);
nor U4100 (N_4100,N_2391,N_913);
nor U4101 (N_4101,N_1385,N_59);
and U4102 (N_4102,N_203,N_1387);
nor U4103 (N_4103,N_1891,N_1406);
and U4104 (N_4104,N_985,N_2040);
nor U4105 (N_4105,N_2574,N_3028);
nand U4106 (N_4106,N_406,N_1714);
nand U4107 (N_4107,N_2875,N_2343);
nor U4108 (N_4108,N_2558,N_3045);
or U4109 (N_4109,N_223,N_1597);
nand U4110 (N_4110,N_1677,N_1725);
and U4111 (N_4111,N_136,N_2202);
nor U4112 (N_4112,N_2863,N_2143);
nand U4113 (N_4113,N_2984,N_3004);
nand U4114 (N_4114,N_1724,N_2603);
xor U4115 (N_4115,N_407,N_2482);
and U4116 (N_4116,N_1116,N_834);
or U4117 (N_4117,N_2818,N_2864);
nand U4118 (N_4118,N_1186,N_771);
xnor U4119 (N_4119,N_180,N_1830);
and U4120 (N_4120,N_1395,N_2030);
xnor U4121 (N_4121,N_1583,N_2624);
xor U4122 (N_4122,N_2758,N_1690);
and U4123 (N_4123,N_155,N_2488);
or U4124 (N_4124,N_2996,N_1461);
and U4125 (N_4125,N_2266,N_2349);
or U4126 (N_4126,N_1863,N_982);
nand U4127 (N_4127,N_1297,N_2042);
nand U4128 (N_4128,N_1794,N_2430);
or U4129 (N_4129,N_784,N_2495);
xnor U4130 (N_4130,N_1553,N_519);
and U4131 (N_4131,N_171,N_657);
or U4132 (N_4132,N_1808,N_3107);
or U4133 (N_4133,N_2821,N_1172);
and U4134 (N_4134,N_866,N_1935);
or U4135 (N_4135,N_2706,N_2399);
nor U4136 (N_4136,N_953,N_2834);
xnor U4137 (N_4137,N_624,N_2766);
nand U4138 (N_4138,N_1767,N_2951);
or U4139 (N_4139,N_2627,N_2812);
and U4140 (N_4140,N_1256,N_2085);
or U4141 (N_4141,N_2586,N_1850);
and U4142 (N_4142,N_1265,N_78);
nand U4143 (N_4143,N_2134,N_2986);
nor U4144 (N_4144,N_2523,N_1929);
or U4145 (N_4145,N_764,N_380);
nand U4146 (N_4146,N_1131,N_1076);
nand U4147 (N_4147,N_1344,N_1077);
nand U4148 (N_4148,N_2229,N_426);
xor U4149 (N_4149,N_870,N_874);
or U4150 (N_4150,N_1201,N_1862);
nor U4151 (N_4151,N_1536,N_1489);
and U4152 (N_4152,N_1921,N_1287);
xor U4153 (N_4153,N_2335,N_276);
or U4154 (N_4154,N_1967,N_968);
nand U4155 (N_4155,N_77,N_2756);
and U4156 (N_4156,N_655,N_2366);
or U4157 (N_4157,N_891,N_2375);
xor U4158 (N_4158,N_1088,N_2428);
or U4159 (N_4159,N_1579,N_1200);
and U4160 (N_4160,N_2833,N_952);
or U4161 (N_4161,N_1363,N_329);
or U4162 (N_4162,N_2410,N_2644);
xnor U4163 (N_4163,N_1932,N_476);
nand U4164 (N_4164,N_1055,N_292);
or U4165 (N_4165,N_2605,N_2625);
nand U4166 (N_4166,N_2444,N_1050);
and U4167 (N_4167,N_2102,N_2385);
and U4168 (N_4168,N_2028,N_253);
or U4169 (N_4169,N_420,N_1199);
nand U4170 (N_4170,N_1599,N_1709);
or U4171 (N_4171,N_1031,N_120);
or U4172 (N_4172,N_1641,N_1471);
or U4173 (N_4173,N_1854,N_1655);
or U4174 (N_4174,N_484,N_2871);
nand U4175 (N_4175,N_1975,N_2508);
xor U4176 (N_4176,N_2442,N_3103);
and U4177 (N_4177,N_3010,N_2794);
or U4178 (N_4178,N_1153,N_916);
nor U4179 (N_4179,N_1425,N_143);
xor U4180 (N_4180,N_181,N_2363);
and U4181 (N_4181,N_2337,N_700);
and U4182 (N_4182,N_2167,N_362);
or U4183 (N_4183,N_1221,N_518);
xor U4184 (N_4184,N_2653,N_945);
and U4185 (N_4185,N_119,N_2109);
and U4186 (N_4186,N_2909,N_581);
nand U4187 (N_4187,N_3120,N_2437);
nor U4188 (N_4188,N_16,N_1847);
and U4189 (N_4189,N_2409,N_469);
nand U4190 (N_4190,N_2452,N_2456);
and U4191 (N_4191,N_2538,N_521);
nand U4192 (N_4192,N_1897,N_679);
xnor U4193 (N_4193,N_573,N_1647);
and U4194 (N_4194,N_2704,N_769);
nand U4195 (N_4195,N_3098,N_2116);
nor U4196 (N_4196,N_2749,N_384);
nor U4197 (N_4197,N_1526,N_216);
nor U4198 (N_4198,N_427,N_1572);
or U4199 (N_4199,N_1813,N_2785);
or U4200 (N_4200,N_2842,N_564);
and U4201 (N_4201,N_1346,N_2615);
nand U4202 (N_4202,N_1502,N_791);
and U4203 (N_4203,N_1937,N_138);
and U4204 (N_4204,N_1109,N_1708);
or U4205 (N_4205,N_1900,N_1822);
or U4206 (N_4206,N_228,N_340);
or U4207 (N_4207,N_2596,N_2740);
nor U4208 (N_4208,N_2062,N_303);
or U4209 (N_4209,N_2534,N_2891);
nor U4210 (N_4210,N_2925,N_397);
or U4211 (N_4211,N_2635,N_157);
and U4212 (N_4212,N_754,N_2159);
nand U4213 (N_4213,N_2576,N_2141);
and U4214 (N_4214,N_65,N_1487);
or U4215 (N_4215,N_931,N_371);
xnor U4216 (N_4216,N_2952,N_1915);
or U4217 (N_4217,N_1328,N_2190);
nand U4218 (N_4218,N_1631,N_1093);
nand U4219 (N_4219,N_430,N_2962);
or U4220 (N_4220,N_2819,N_833);
nor U4221 (N_4221,N_1629,N_385);
nand U4222 (N_4222,N_2089,N_793);
or U4223 (N_4223,N_2950,N_1498);
xnor U4224 (N_4224,N_2655,N_205);
nor U4225 (N_4225,N_2024,N_1713);
and U4226 (N_4226,N_2047,N_1054);
and U4227 (N_4227,N_1030,N_498);
or U4228 (N_4228,N_271,N_2683);
or U4229 (N_4229,N_3066,N_425);
nand U4230 (N_4230,N_1428,N_2998);
nor U4231 (N_4231,N_2926,N_523);
and U4232 (N_4232,N_3,N_2885);
and U4233 (N_4233,N_1898,N_2547);
xnor U4234 (N_4234,N_158,N_2579);
and U4235 (N_4235,N_246,N_947);
or U4236 (N_4236,N_1982,N_217);
nor U4237 (N_4237,N_2425,N_567);
xor U4238 (N_4238,N_149,N_2569);
nand U4239 (N_4239,N_2777,N_1615);
nor U4240 (N_4240,N_1411,N_1610);
nor U4241 (N_4241,N_73,N_682);
nand U4242 (N_4242,N_1550,N_994);
xor U4243 (N_4243,N_339,N_1584);
or U4244 (N_4244,N_240,N_2041);
or U4245 (N_4245,N_1520,N_1698);
nand U4246 (N_4246,N_1241,N_478);
and U4247 (N_4247,N_623,N_1747);
or U4248 (N_4248,N_2957,N_991);
xor U4249 (N_4249,N_2575,N_1415);
xnor U4250 (N_4250,N_591,N_3077);
and U4251 (N_4251,N_285,N_2739);
or U4252 (N_4252,N_3071,N_554);
and U4253 (N_4253,N_1669,N_208);
nand U4254 (N_4254,N_2420,N_1090);
nand U4255 (N_4255,N_2439,N_795);
nand U4256 (N_4256,N_39,N_2691);
nand U4257 (N_4257,N_675,N_3102);
and U4258 (N_4258,N_365,N_2236);
xnor U4259 (N_4259,N_410,N_1642);
nand U4260 (N_4260,N_2358,N_1210);
and U4261 (N_4261,N_1620,N_383);
and U4262 (N_4262,N_1144,N_878);
xnor U4263 (N_4263,N_1238,N_3089);
xor U4264 (N_4264,N_107,N_2967);
nor U4265 (N_4265,N_2540,N_694);
nand U4266 (N_4266,N_1393,N_71);
nand U4267 (N_4267,N_1220,N_1203);
xor U4268 (N_4268,N_2004,N_62);
and U4269 (N_4269,N_2985,N_1878);
or U4270 (N_4270,N_2767,N_1961);
nor U4271 (N_4271,N_1919,N_605);
xor U4272 (N_4272,N_1230,N_1594);
nor U4273 (N_4273,N_209,N_2904);
xor U4274 (N_4274,N_437,N_2303);
and U4275 (N_4275,N_1955,N_1551);
xnor U4276 (N_4276,N_126,N_637);
or U4277 (N_4277,N_949,N_2049);
or U4278 (N_4278,N_2301,N_1687);
xnor U4279 (N_4279,N_2231,N_2813);
nand U4280 (N_4280,N_1353,N_2323);
nor U4281 (N_4281,N_2702,N_121);
or U4282 (N_4282,N_1882,N_182);
and U4283 (N_4283,N_824,N_2509);
xor U4284 (N_4284,N_2632,N_2217);
xnor U4285 (N_4285,N_3092,N_104);
nor U4286 (N_4286,N_22,N_337);
nor U4287 (N_4287,N_2327,N_506);
and U4288 (N_4288,N_1009,N_794);
xor U4289 (N_4289,N_993,N_783);
nand U4290 (N_4290,N_1789,N_692);
or U4291 (N_4291,N_570,N_2884);
nor U4292 (N_4292,N_265,N_1059);
nand U4293 (N_4293,N_2205,N_903);
and U4294 (N_4294,N_467,N_3085);
or U4295 (N_4295,N_1673,N_122);
xor U4296 (N_4296,N_2105,N_2732);
xnor U4297 (N_4297,N_1012,N_2226);
xor U4298 (N_4298,N_1493,N_1778);
and U4299 (N_4299,N_1147,N_777);
nand U4300 (N_4300,N_2272,N_3113);
or U4301 (N_4301,N_1772,N_344);
and U4302 (N_4302,N_1762,N_390);
or U4303 (N_4303,N_1763,N_2270);
nand U4304 (N_4304,N_572,N_2517);
xnor U4305 (N_4305,N_2815,N_2445);
or U4306 (N_4306,N_1026,N_604);
nor U4307 (N_4307,N_1828,N_2695);
nand U4308 (N_4308,N_140,N_1591);
nor U4309 (N_4309,N_308,N_335);
nor U4310 (N_4310,N_1206,N_313);
xor U4311 (N_4311,N_2837,N_924);
xnor U4312 (N_4312,N_2890,N_2768);
and U4313 (N_4313,N_2994,N_1196);
nor U4314 (N_4314,N_2311,N_1912);
nand U4315 (N_4315,N_1849,N_1805);
nor U4316 (N_4316,N_1777,N_1519);
xnor U4317 (N_4317,N_2573,N_500);
nor U4318 (N_4318,N_1326,N_958);
nand U4319 (N_4319,N_3021,N_543);
xor U4320 (N_4320,N_1322,N_2725);
and U4321 (N_4321,N_2400,N_1211);
nand U4322 (N_4322,N_448,N_2734);
nand U4323 (N_4323,N_1657,N_2325);
xnor U4324 (N_4324,N_664,N_84);
or U4325 (N_4325,N_3104,N_445);
and U4326 (N_4326,N_2253,N_2112);
nor U4327 (N_4327,N_2076,N_1966);
and U4328 (N_4328,N_2751,N_613);
nor U4329 (N_4329,N_1727,N_92);
and U4330 (N_4330,N_204,N_1616);
nand U4331 (N_4331,N_2440,N_2761);
and U4332 (N_4332,N_670,N_2168);
xor U4333 (N_4333,N_3062,N_1998);
or U4334 (N_4334,N_449,N_2379);
nand U4335 (N_4335,N_2378,N_1868);
nand U4336 (N_4336,N_1070,N_1593);
xnor U4337 (N_4337,N_2914,N_1274);
nor U4338 (N_4338,N_2585,N_2031);
nor U4339 (N_4339,N_1041,N_957);
or U4340 (N_4340,N_1156,N_1861);
xnor U4341 (N_4341,N_1603,N_2600);
nor U4342 (N_4342,N_2027,N_1045);
nor U4343 (N_4343,N_2368,N_393);
nor U4344 (N_4344,N_3053,N_3025);
nand U4345 (N_4345,N_1233,N_2805);
nand U4346 (N_4346,N_2137,N_10);
xnor U4347 (N_4347,N_2736,N_1404);
or U4348 (N_4348,N_91,N_2714);
nand U4349 (N_4349,N_1662,N_2377);
xor U4350 (N_4350,N_2408,N_2528);
xor U4351 (N_4351,N_358,N_671);
nor U4352 (N_4352,N_274,N_2120);
and U4353 (N_4353,N_8,N_707);
xor U4354 (N_4354,N_2162,N_676);
nor U4355 (N_4355,N_2114,N_3094);
nand U4356 (N_4356,N_2015,N_2108);
nor U4357 (N_4357,N_531,N_1102);
or U4358 (N_4358,N_192,N_2156);
and U4359 (N_4359,N_1856,N_2305);
xor U4360 (N_4360,N_2938,N_2827);
or U4361 (N_4361,N_1313,N_1352);
and U4362 (N_4362,N_2999,N_202);
xor U4363 (N_4363,N_1259,N_760);
nand U4364 (N_4364,N_226,N_2310);
nor U4365 (N_4365,N_1281,N_497);
nand U4366 (N_4366,N_582,N_1793);
nor U4367 (N_4367,N_2836,N_964);
xor U4368 (N_4368,N_366,N_2474);
xnor U4369 (N_4369,N_3067,N_2397);
nor U4370 (N_4370,N_3020,N_2292);
nand U4371 (N_4371,N_1950,N_1788);
xor U4372 (N_4372,N_174,N_200);
xnor U4373 (N_4373,N_1283,N_421);
nor U4374 (N_4374,N_552,N_2443);
and U4375 (N_4375,N_2033,N_367);
nor U4376 (N_4376,N_934,N_2669);
nand U4377 (N_4377,N_319,N_1522);
nand U4378 (N_4378,N_673,N_320);
and U4379 (N_4379,N_373,N_352);
or U4380 (N_4380,N_2121,N_103);
or U4381 (N_4381,N_1954,N_1082);
xnor U4382 (N_4382,N_1706,N_634);
nor U4383 (N_4383,N_1396,N_2667);
or U4384 (N_4384,N_218,N_2151);
and U4385 (N_4385,N_2797,N_172);
nor U4386 (N_4386,N_772,N_1017);
nor U4387 (N_4387,N_2623,N_2467);
xor U4388 (N_4388,N_2262,N_2798);
nand U4389 (N_4389,N_1812,N_597);
and U4390 (N_4390,N_2665,N_2803);
nand U4391 (N_4391,N_3056,N_1263);
nor U4392 (N_4392,N_697,N_1181);
nand U4393 (N_4393,N_2898,N_1064);
and U4394 (N_4394,N_2825,N_1429);
nand U4395 (N_4395,N_744,N_2299);
nor U4396 (N_4396,N_2676,N_1748);
xor U4397 (N_4397,N_3011,N_206);
nor U4398 (N_4398,N_2081,N_1978);
nand U4399 (N_4399,N_2712,N_166);
xor U4400 (N_4400,N_2783,N_2544);
xor U4401 (N_4401,N_1004,N_69);
nand U4402 (N_4402,N_843,N_992);
nand U4403 (N_4403,N_2152,N_1782);
and U4404 (N_4404,N_2321,N_1285);
xor U4405 (N_4405,N_887,N_2522);
xnor U4406 (N_4406,N_185,N_1084);
nor U4407 (N_4407,N_2178,N_377);
or U4408 (N_4408,N_2254,N_2746);
xor U4409 (N_4409,N_2277,N_933);
or U4410 (N_4410,N_2848,N_1924);
or U4411 (N_4411,N_2471,N_1563);
and U4412 (N_4412,N_1121,N_969);
nor U4413 (N_4413,N_1586,N_508);
or U4414 (N_4414,N_98,N_1827);
and U4415 (N_4415,N_295,N_2463);
nor U4416 (N_4416,N_681,N_2022);
nor U4417 (N_4417,N_314,N_1768);
nor U4418 (N_4418,N_74,N_2515);
nor U4419 (N_4419,N_2553,N_633);
nand U4420 (N_4420,N_1716,N_1886);
xnor U4421 (N_4421,N_2249,N_2822);
xnor U4422 (N_4422,N_334,N_2005);
or U4423 (N_4423,N_1422,N_2567);
nand U4424 (N_4424,N_2419,N_2869);
nor U4425 (N_4425,N_2977,N_2643);
xor U4426 (N_4426,N_2285,N_2380);
xnor U4427 (N_4427,N_2867,N_1399);
and U4428 (N_4428,N_2549,N_2283);
and U4429 (N_4429,N_649,N_2111);
nand U4430 (N_4430,N_2251,N_2407);
or U4431 (N_4431,N_1507,N_2622);
or U4432 (N_4432,N_1931,N_1565);
and U4433 (N_4433,N_1881,N_978);
xor U4434 (N_4434,N_191,N_2670);
xor U4435 (N_4435,N_2350,N_1355);
nor U4436 (N_4436,N_2776,N_2844);
nand U4437 (N_4437,N_629,N_1369);
and U4438 (N_4438,N_997,N_2782);
xor U4439 (N_4439,N_1460,N_2459);
nor U4440 (N_4440,N_2905,N_2820);
xnor U4441 (N_4441,N_540,N_1194);
xor U4442 (N_4442,N_562,N_2093);
and U4443 (N_4443,N_294,N_1696);
or U4444 (N_4444,N_2919,N_2123);
and U4445 (N_4445,N_1431,N_97);
and U4446 (N_4446,N_2840,N_270);
nand U4447 (N_4447,N_2606,N_1252);
or U4448 (N_4448,N_1005,N_839);
xnor U4449 (N_4449,N_1335,N_3041);
nand U4450 (N_4450,N_1786,N_1779);
xnor U4451 (N_4451,N_2073,N_2828);
and U4452 (N_4452,N_2078,N_2455);
nand U4453 (N_4453,N_1785,N_881);
and U4454 (N_4454,N_3057,N_1388);
xor U4455 (N_4455,N_2250,N_2320);
and U4456 (N_4456,N_2861,N_2284);
xnor U4457 (N_4457,N_1062,N_2532);
and U4458 (N_4458,N_266,N_2043);
nand U4459 (N_4459,N_2019,N_2945);
nand U4460 (N_4460,N_1595,N_1257);
xnor U4461 (N_4461,N_618,N_1160);
nor U4462 (N_4462,N_3051,N_1561);
xnor U4463 (N_4463,N_2677,N_2263);
and U4464 (N_4464,N_2966,N_594);
or U4465 (N_4465,N_2970,N_343);
and U4466 (N_4466,N_1458,N_1934);
and U4467 (N_4467,N_1491,N_1359);
nand U4468 (N_4468,N_796,N_1127);
xor U4469 (N_4469,N_333,N_2638);
xnor U4470 (N_4470,N_284,N_2769);
and U4471 (N_4471,N_647,N_1100);
nor U4472 (N_4472,N_2760,N_1433);
or U4473 (N_4473,N_1906,N_2170);
xor U4474 (N_4474,N_1582,N_3093);
or U4475 (N_4475,N_1939,N_1617);
and U4476 (N_4476,N_117,N_3119);
nor U4477 (N_4477,N_2281,N_1571);
or U4478 (N_4478,N_1835,N_1781);
xor U4479 (N_4479,N_306,N_683);
nand U4480 (N_4480,N_1672,N_1020);
nor U4481 (N_4481,N_2146,N_2791);
nand U4482 (N_4482,N_2688,N_219);
and U4483 (N_4483,N_2992,N_763);
nand U4484 (N_4484,N_1282,N_651);
nor U4485 (N_4485,N_940,N_387);
nand U4486 (N_4486,N_1195,N_998);
nor U4487 (N_4487,N_1972,N_2542);
nand U4488 (N_4488,N_2874,N_1776);
nand U4489 (N_4489,N_1928,N_1653);
nor U4490 (N_4490,N_736,N_277);
nor U4491 (N_4491,N_450,N_2737);
nand U4492 (N_4492,N_2601,N_1337);
and U4493 (N_4493,N_2501,N_46);
nand U4494 (N_4494,N_2738,N_1918);
nor U4495 (N_4495,N_1455,N_2052);
or U4496 (N_4496,N_830,N_2095);
nand U4497 (N_4497,N_1474,N_1370);
nand U4498 (N_4498,N_2763,N_909);
or U4499 (N_4499,N_2091,N_1976);
xor U4500 (N_4500,N_401,N_2511);
or U4501 (N_4501,N_1981,N_666);
nor U4502 (N_4502,N_1730,N_2313);
and U4503 (N_4503,N_858,N_1971);
nand U4504 (N_4504,N_1799,N_1640);
xnor U4505 (N_4505,N_1740,N_1951);
or U4506 (N_4506,N_9,N_2039);
nor U4507 (N_4507,N_1424,N_1058);
xor U4508 (N_4508,N_677,N_1819);
xor U4509 (N_4509,N_86,N_2868);
nor U4510 (N_4510,N_409,N_83);
and U4511 (N_4511,N_2055,N_1464);
xor U4512 (N_4512,N_1305,N_1959);
and U4513 (N_4513,N_746,N_1225);
and U4514 (N_4514,N_1581,N_1188);
and U4515 (N_4515,N_954,N_2433);
nand U4516 (N_4516,N_1911,N_904);
nand U4517 (N_4517,N_1559,N_1133);
nor U4518 (N_4518,N_2359,N_2765);
or U4519 (N_4519,N_1039,N_1885);
or U4520 (N_4520,N_135,N_820);
nand U4521 (N_4521,N_1717,N_3008);
or U4522 (N_4522,N_601,N_1034);
nor U4523 (N_4523,N_630,N_1438);
xnor U4524 (N_4524,N_2773,N_403);
nor U4525 (N_4525,N_2370,N_475);
or U4526 (N_4526,N_1457,N_787);
nor U4527 (N_4527,N_2658,N_2759);
or U4528 (N_4528,N_1047,N_150);
nor U4529 (N_4529,N_1165,N_2722);
nand U4530 (N_4530,N_2476,N_961);
or U4531 (N_4531,N_2038,N_176);
nor U4532 (N_4532,N_310,N_2787);
nor U4533 (N_4533,N_2548,N_975);
nor U4534 (N_4534,N_2189,N_238);
and U4535 (N_4535,N_1621,N_930);
nor U4536 (N_4536,N_1607,N_658);
and U4537 (N_4537,N_1695,N_1661);
or U4538 (N_4538,N_1826,N_229);
and U4539 (N_4539,N_2074,N_1558);
nand U4540 (N_4540,N_2684,N_530);
and U4541 (N_4541,N_807,N_6);
nor U4542 (N_4542,N_1656,N_2329);
or U4543 (N_4543,N_2014,N_1409);
and U4544 (N_4544,N_2882,N_2578);
nor U4545 (N_4545,N_3022,N_133);
or U4546 (N_4546,N_871,N_1391);
or U4547 (N_4547,N_2546,N_1649);
nor U4548 (N_4548,N_1162,N_524);
xor U4549 (N_4549,N_1948,N_1648);
nor U4550 (N_4550,N_2972,N_1198);
nand U4551 (N_4551,N_2641,N_3086);
xnor U4552 (N_4552,N_780,N_1697);
nor U4553 (N_4553,N_558,N_775);
or U4554 (N_4554,N_541,N_2177);
and U4555 (N_4555,N_2341,N_1295);
nor U4556 (N_4556,N_1260,N_1517);
xor U4557 (N_4557,N_2617,N_1099);
xor U4558 (N_4558,N_291,N_1941);
xnor U4559 (N_4559,N_1893,N_1575);
nor U4560 (N_4560,N_1566,N_2878);
nor U4561 (N_4561,N_1418,N_2703);
and U4562 (N_4562,N_177,N_2502);
or U4563 (N_4563,N_1499,N_1787);
and U4564 (N_4564,N_1208,N_989);
xnor U4565 (N_4565,N_1185,N_2309);
nor U4566 (N_4566,N_1842,N_165);
or U4567 (N_4567,N_1132,N_588);
xnor U4568 (N_4568,N_753,N_1123);
xor U4569 (N_4569,N_2314,N_2802);
and U4570 (N_4570,N_369,N_1134);
xnor U4571 (N_4571,N_2118,N_1543);
xnor U4572 (N_4572,N_2344,N_1938);
nor U4573 (N_4573,N_838,N_2699);
and U4574 (N_4574,N_160,N_2394);
nand U4575 (N_4575,N_1497,N_1080);
nand U4576 (N_4576,N_2559,N_3101);
nand U4577 (N_4577,N_1970,N_132);
or U4578 (N_4578,N_1703,N_2113);
xnor U4579 (N_4579,N_786,N_457);
nor U4580 (N_4580,N_1739,N_2125);
nor U4581 (N_4581,N_363,N_2328);
nor U4582 (N_4582,N_2169,N_2075);
nand U4583 (N_4583,N_1357,N_3003);
xor U4584 (N_4584,N_3087,N_1963);
or U4585 (N_4585,N_118,N_2388);
or U4586 (N_4586,N_60,N_1289);
and U4587 (N_4587,N_525,N_1742);
nor U4588 (N_4588,N_1382,N_1635);
nor U4589 (N_4589,N_2735,N_2131);
nand U4590 (N_4590,N_414,N_2887);
nor U4591 (N_4591,N_789,N_27);
xnor U4592 (N_4592,N_57,N_571);
nand U4593 (N_4593,N_822,N_1075);
nor U4594 (N_4594,N_974,N_2661);
or U4595 (N_4595,N_37,N_1542);
and U4596 (N_4596,N_2147,N_1033);
xnor U4597 (N_4597,N_1348,N_929);
or U4598 (N_4598,N_360,N_2244);
nand U4599 (N_4599,N_2196,N_2260);
nand U4600 (N_4600,N_3090,N_32);
and U4601 (N_4601,N_2524,N_289);
nor U4602 (N_4602,N_336,N_2032);
nor U4603 (N_4603,N_2148,N_2552);
or U4604 (N_4604,N_2220,N_2831);
or U4605 (N_4605,N_1000,N_3060);
xnor U4606 (N_4606,N_861,N_1936);
and U4607 (N_4607,N_900,N_595);
or U4608 (N_4608,N_1314,N_394);
or U4609 (N_4609,N_3109,N_829);
nand U4610 (N_4610,N_542,N_1300);
or U4611 (N_4611,N_38,N_1074);
and U4612 (N_4612,N_1802,N_1079);
or U4613 (N_4613,N_2531,N_225);
nand U4614 (N_4614,N_2728,N_1666);
nor U4615 (N_4615,N_939,N_3054);
and U4616 (N_4616,N_2612,N_688);
or U4617 (N_4617,N_378,N_2873);
nor U4618 (N_4618,N_1501,N_2184);
and U4619 (N_4619,N_2466,N_825);
and U4620 (N_4620,N_1999,N_678);
and U4621 (N_4621,N_1663,N_1814);
nor U4622 (N_4622,N_529,N_2496);
or U4623 (N_4623,N_1384,N_2373);
nand U4624 (N_4624,N_1723,N_273);
nand U4625 (N_4625,N_1784,N_548);
nor U4626 (N_4626,N_35,N_1158);
xnor U4627 (N_4627,N_2312,N_927);
xnor U4628 (N_4628,N_1853,N_505);
or U4629 (N_4629,N_2806,N_1681);
and U4630 (N_4630,N_1266,N_2046);
or U4631 (N_4631,N_477,N_1521);
and U4632 (N_4632,N_2450,N_638);
and U4633 (N_4633,N_596,N_2230);
xor U4634 (N_4634,N_2514,N_1995);
and U4635 (N_4635,N_776,N_2);
nand U4636 (N_4636,N_342,N_1317);
or U4637 (N_4637,N_2566,N_1843);
xnor U4638 (N_4638,N_632,N_1554);
nor U4639 (N_4639,N_1806,N_1684);
and U4640 (N_4640,N_1092,N_1089);
xor U4641 (N_4641,N_281,N_255);
nand U4642 (N_4642,N_718,N_2937);
nor U4643 (N_4643,N_535,N_888);
or U4644 (N_4644,N_297,N_1688);
nor U4645 (N_4645,N_1923,N_1119);
xor U4646 (N_4646,N_1980,N_2932);
nand U4647 (N_4647,N_2587,N_1468);
nand U4648 (N_4648,N_431,N_2943);
nor U4649 (N_4649,N_2269,N_1547);
xnor U4650 (N_4650,N_2847,N_811);
nand U4651 (N_4651,N_2694,N_668);
and U4652 (N_4652,N_1492,N_1098);
and U4653 (N_4653,N_1278,N_1247);
xnor U4654 (N_4654,N_1453,N_1833);
nand U4655 (N_4655,N_1168,N_131);
or U4656 (N_4656,N_1356,N_1602);
nand U4657 (N_4657,N_2417,N_392);
or U4658 (N_4658,N_1380,N_1500);
and U4659 (N_4659,N_2139,N_1894);
and U4660 (N_4660,N_1839,N_1443);
nand U4661 (N_4661,N_79,N_1732);
or U4662 (N_4662,N_93,N_230);
nand U4663 (N_4663,N_884,N_1292);
nor U4664 (N_4664,N_14,N_1051);
xnor U4665 (N_4665,N_2707,N_3043);
and U4666 (N_4666,N_304,N_2991);
and U4667 (N_4667,N_263,N_2817);
or U4668 (N_4668,N_2008,N_179);
nand U4669 (N_4669,N_1743,N_1860);
nand U4670 (N_4670,N_648,N_544);
nor U4671 (N_4671,N_2056,N_2207);
nand U4672 (N_4672,N_1818,N_1167);
nand U4673 (N_4673,N_2933,N_3115);
nand U4674 (N_4674,N_2789,N_2934);
or U4675 (N_4675,N_1552,N_691);
nand U4676 (N_4676,N_286,N_489);
nand U4677 (N_4677,N_2185,N_1374);
nor U4678 (N_4678,N_2597,N_768);
and U4679 (N_4679,N_2234,N_11);
nand U4680 (N_4680,N_42,N_865);
xnor U4681 (N_4681,N_1215,N_2058);
and U4682 (N_4682,N_3070,N_2554);
and U4683 (N_4683,N_2963,N_622);
and U4684 (N_4684,N_2845,N_2572);
nor U4685 (N_4685,N_2140,N_349);
and U4686 (N_4686,N_2149,N_2086);
xor U4687 (N_4687,N_808,N_2459);
nand U4688 (N_4688,N_2403,N_201);
nand U4689 (N_4689,N_641,N_973);
nor U4690 (N_4690,N_2218,N_1998);
nor U4691 (N_4691,N_1717,N_3110);
nand U4692 (N_4692,N_2390,N_2336);
xnor U4693 (N_4693,N_332,N_733);
nor U4694 (N_4694,N_1954,N_1173);
xnor U4695 (N_4695,N_1656,N_2123);
and U4696 (N_4696,N_2368,N_386);
and U4697 (N_4697,N_2479,N_2979);
nor U4698 (N_4698,N_1212,N_2107);
nor U4699 (N_4699,N_880,N_86);
and U4700 (N_4700,N_2415,N_1448);
or U4701 (N_4701,N_1937,N_1815);
nand U4702 (N_4702,N_299,N_245);
or U4703 (N_4703,N_673,N_733);
nor U4704 (N_4704,N_2054,N_30);
and U4705 (N_4705,N_152,N_1293);
nand U4706 (N_4706,N_2092,N_2519);
and U4707 (N_4707,N_1396,N_2222);
nand U4708 (N_4708,N_824,N_1225);
and U4709 (N_4709,N_3121,N_1868);
nand U4710 (N_4710,N_1661,N_385);
and U4711 (N_4711,N_1815,N_1632);
nor U4712 (N_4712,N_838,N_2280);
or U4713 (N_4713,N_1838,N_615);
nand U4714 (N_4714,N_720,N_1493);
or U4715 (N_4715,N_2724,N_330);
xnor U4716 (N_4716,N_2902,N_2932);
xor U4717 (N_4717,N_2003,N_2704);
or U4718 (N_4718,N_474,N_2010);
nor U4719 (N_4719,N_2691,N_2525);
or U4720 (N_4720,N_1501,N_385);
xnor U4721 (N_4721,N_178,N_3113);
xor U4722 (N_4722,N_1196,N_2476);
and U4723 (N_4723,N_27,N_163);
xnor U4724 (N_4724,N_1335,N_1210);
nand U4725 (N_4725,N_3052,N_3017);
or U4726 (N_4726,N_1212,N_2005);
xnor U4727 (N_4727,N_2898,N_2109);
or U4728 (N_4728,N_2763,N_1157);
nand U4729 (N_4729,N_1672,N_1383);
nand U4730 (N_4730,N_121,N_2461);
nand U4731 (N_4731,N_1536,N_3052);
and U4732 (N_4732,N_2256,N_2770);
nor U4733 (N_4733,N_2108,N_2878);
or U4734 (N_4734,N_2542,N_1239);
nor U4735 (N_4735,N_1177,N_386);
nor U4736 (N_4736,N_1939,N_3098);
nand U4737 (N_4737,N_1940,N_781);
and U4738 (N_4738,N_811,N_2915);
and U4739 (N_4739,N_726,N_1447);
xnor U4740 (N_4740,N_2797,N_631);
and U4741 (N_4741,N_2325,N_1169);
and U4742 (N_4742,N_2358,N_2147);
nand U4743 (N_4743,N_356,N_3022);
nor U4744 (N_4744,N_1249,N_986);
or U4745 (N_4745,N_1911,N_1242);
xnor U4746 (N_4746,N_418,N_2808);
nand U4747 (N_4747,N_2548,N_240);
xnor U4748 (N_4748,N_1002,N_1920);
nor U4749 (N_4749,N_1848,N_169);
xor U4750 (N_4750,N_2294,N_1390);
nor U4751 (N_4751,N_2567,N_701);
and U4752 (N_4752,N_2485,N_1972);
nor U4753 (N_4753,N_2010,N_1007);
or U4754 (N_4754,N_841,N_16);
nor U4755 (N_4755,N_1372,N_163);
and U4756 (N_4756,N_1618,N_2611);
xnor U4757 (N_4757,N_300,N_46);
nand U4758 (N_4758,N_2894,N_1924);
nor U4759 (N_4759,N_1674,N_23);
and U4760 (N_4760,N_2346,N_1677);
xnor U4761 (N_4761,N_2315,N_1354);
nor U4762 (N_4762,N_3073,N_894);
or U4763 (N_4763,N_1834,N_1129);
nor U4764 (N_4764,N_1580,N_2311);
and U4765 (N_4765,N_3109,N_3041);
or U4766 (N_4766,N_353,N_7);
nor U4767 (N_4767,N_3111,N_2460);
nor U4768 (N_4768,N_2575,N_2611);
xnor U4769 (N_4769,N_2580,N_476);
and U4770 (N_4770,N_766,N_1069);
and U4771 (N_4771,N_707,N_2824);
nor U4772 (N_4772,N_2189,N_204);
nand U4773 (N_4773,N_319,N_1339);
nand U4774 (N_4774,N_1190,N_2249);
nor U4775 (N_4775,N_1736,N_2859);
xor U4776 (N_4776,N_2056,N_150);
nand U4777 (N_4777,N_2031,N_547);
nor U4778 (N_4778,N_2507,N_1764);
xnor U4779 (N_4779,N_1835,N_673);
or U4780 (N_4780,N_2556,N_2346);
xor U4781 (N_4781,N_1388,N_2980);
nor U4782 (N_4782,N_2256,N_2059);
xnor U4783 (N_4783,N_1802,N_493);
and U4784 (N_4784,N_1594,N_1168);
nand U4785 (N_4785,N_3090,N_2665);
or U4786 (N_4786,N_548,N_414);
xnor U4787 (N_4787,N_166,N_2550);
nand U4788 (N_4788,N_104,N_804);
and U4789 (N_4789,N_967,N_1062);
and U4790 (N_4790,N_560,N_714);
and U4791 (N_4791,N_1836,N_1424);
nor U4792 (N_4792,N_1246,N_691);
or U4793 (N_4793,N_284,N_1930);
or U4794 (N_4794,N_2102,N_2936);
nor U4795 (N_4795,N_344,N_2156);
or U4796 (N_4796,N_2144,N_2975);
or U4797 (N_4797,N_1196,N_82);
nand U4798 (N_4798,N_714,N_554);
nor U4799 (N_4799,N_1473,N_729);
xor U4800 (N_4800,N_486,N_245);
nand U4801 (N_4801,N_537,N_507);
and U4802 (N_4802,N_1826,N_2680);
nor U4803 (N_4803,N_1281,N_1383);
xnor U4804 (N_4804,N_999,N_1459);
nor U4805 (N_4805,N_921,N_154);
and U4806 (N_4806,N_2559,N_233);
or U4807 (N_4807,N_1028,N_652);
or U4808 (N_4808,N_1061,N_3001);
nand U4809 (N_4809,N_423,N_298);
and U4810 (N_4810,N_2817,N_1895);
nor U4811 (N_4811,N_1010,N_2287);
and U4812 (N_4812,N_933,N_1219);
nand U4813 (N_4813,N_242,N_1344);
and U4814 (N_4814,N_184,N_2098);
xor U4815 (N_4815,N_2979,N_1867);
nand U4816 (N_4816,N_2465,N_2951);
nor U4817 (N_4817,N_2757,N_1216);
nor U4818 (N_4818,N_2740,N_2201);
xnor U4819 (N_4819,N_2761,N_2889);
and U4820 (N_4820,N_2881,N_3013);
nor U4821 (N_4821,N_2476,N_1663);
nor U4822 (N_4822,N_1232,N_2793);
and U4823 (N_4823,N_792,N_646);
xor U4824 (N_4824,N_2976,N_2345);
and U4825 (N_4825,N_2497,N_2089);
xor U4826 (N_4826,N_2468,N_574);
xor U4827 (N_4827,N_1685,N_2741);
or U4828 (N_4828,N_323,N_316);
nor U4829 (N_4829,N_1083,N_803);
and U4830 (N_4830,N_212,N_325);
or U4831 (N_4831,N_1926,N_2817);
nor U4832 (N_4832,N_73,N_1625);
xnor U4833 (N_4833,N_1515,N_2805);
and U4834 (N_4834,N_586,N_1999);
xor U4835 (N_4835,N_1876,N_342);
or U4836 (N_4836,N_2083,N_465);
nor U4837 (N_4837,N_256,N_589);
nor U4838 (N_4838,N_783,N_314);
and U4839 (N_4839,N_1306,N_1538);
nor U4840 (N_4840,N_2051,N_1969);
and U4841 (N_4841,N_2679,N_2141);
nand U4842 (N_4842,N_1780,N_57);
and U4843 (N_4843,N_2206,N_2549);
nand U4844 (N_4844,N_2996,N_404);
xor U4845 (N_4845,N_1251,N_411);
nor U4846 (N_4846,N_2889,N_193);
xnor U4847 (N_4847,N_1943,N_731);
nand U4848 (N_4848,N_1801,N_3079);
or U4849 (N_4849,N_2692,N_2690);
and U4850 (N_4850,N_114,N_1951);
nand U4851 (N_4851,N_2941,N_1197);
xor U4852 (N_4852,N_2933,N_2042);
nand U4853 (N_4853,N_2031,N_1212);
nor U4854 (N_4854,N_1426,N_657);
and U4855 (N_4855,N_378,N_972);
nor U4856 (N_4856,N_2739,N_1272);
and U4857 (N_4857,N_1048,N_2090);
xnor U4858 (N_4858,N_358,N_721);
xnor U4859 (N_4859,N_941,N_1758);
nor U4860 (N_4860,N_2053,N_1416);
nand U4861 (N_4861,N_445,N_235);
xnor U4862 (N_4862,N_1518,N_2843);
nor U4863 (N_4863,N_2389,N_980);
and U4864 (N_4864,N_443,N_547);
nand U4865 (N_4865,N_2480,N_578);
xnor U4866 (N_4866,N_1491,N_541);
and U4867 (N_4867,N_2907,N_2172);
nand U4868 (N_4868,N_1223,N_267);
nor U4869 (N_4869,N_2758,N_3073);
nor U4870 (N_4870,N_1307,N_2966);
or U4871 (N_4871,N_2673,N_2304);
and U4872 (N_4872,N_1031,N_1545);
and U4873 (N_4873,N_608,N_2855);
nand U4874 (N_4874,N_627,N_2049);
nand U4875 (N_4875,N_986,N_2420);
and U4876 (N_4876,N_2725,N_1764);
or U4877 (N_4877,N_1265,N_363);
and U4878 (N_4878,N_2268,N_1707);
or U4879 (N_4879,N_402,N_1182);
xor U4880 (N_4880,N_2705,N_939);
xor U4881 (N_4881,N_2656,N_172);
xnor U4882 (N_4882,N_608,N_2441);
or U4883 (N_4883,N_583,N_1072);
xor U4884 (N_4884,N_3060,N_304);
and U4885 (N_4885,N_2598,N_2393);
nor U4886 (N_4886,N_1758,N_2686);
xor U4887 (N_4887,N_2034,N_1995);
nand U4888 (N_4888,N_584,N_2117);
or U4889 (N_4889,N_2063,N_1911);
xor U4890 (N_4890,N_2331,N_64);
and U4891 (N_4891,N_2854,N_98);
nor U4892 (N_4892,N_73,N_2460);
and U4893 (N_4893,N_2676,N_1427);
or U4894 (N_4894,N_862,N_2144);
nand U4895 (N_4895,N_672,N_1162);
nor U4896 (N_4896,N_580,N_333);
or U4897 (N_4897,N_2751,N_2006);
nor U4898 (N_4898,N_2905,N_336);
nor U4899 (N_4899,N_1001,N_1962);
and U4900 (N_4900,N_1815,N_960);
nand U4901 (N_4901,N_1766,N_1273);
and U4902 (N_4902,N_188,N_727);
or U4903 (N_4903,N_2135,N_1808);
or U4904 (N_4904,N_2859,N_1400);
xnor U4905 (N_4905,N_1190,N_1254);
nand U4906 (N_4906,N_588,N_143);
or U4907 (N_4907,N_736,N_2704);
and U4908 (N_4908,N_2492,N_1478);
and U4909 (N_4909,N_1689,N_2506);
or U4910 (N_4910,N_3026,N_2132);
nor U4911 (N_4911,N_429,N_2839);
and U4912 (N_4912,N_1073,N_2772);
nor U4913 (N_4913,N_1379,N_2398);
nor U4914 (N_4914,N_1083,N_2193);
or U4915 (N_4915,N_60,N_808);
or U4916 (N_4916,N_1953,N_1143);
and U4917 (N_4917,N_108,N_1617);
nor U4918 (N_4918,N_922,N_2982);
xnor U4919 (N_4919,N_1971,N_322);
and U4920 (N_4920,N_2206,N_215);
nor U4921 (N_4921,N_1146,N_1577);
nand U4922 (N_4922,N_2220,N_2421);
or U4923 (N_4923,N_1568,N_174);
nor U4924 (N_4924,N_1797,N_2371);
xor U4925 (N_4925,N_489,N_2929);
xnor U4926 (N_4926,N_1769,N_1081);
and U4927 (N_4927,N_2728,N_539);
xnor U4928 (N_4928,N_1290,N_2278);
or U4929 (N_4929,N_2871,N_104);
nor U4930 (N_4930,N_3081,N_1816);
and U4931 (N_4931,N_454,N_2783);
and U4932 (N_4932,N_1488,N_1359);
or U4933 (N_4933,N_1416,N_1008);
nand U4934 (N_4934,N_1714,N_1922);
nand U4935 (N_4935,N_1524,N_2220);
nand U4936 (N_4936,N_2613,N_406);
nand U4937 (N_4937,N_630,N_1380);
nor U4938 (N_4938,N_2111,N_1752);
xor U4939 (N_4939,N_2142,N_2782);
xnor U4940 (N_4940,N_391,N_1270);
or U4941 (N_4941,N_1056,N_1911);
or U4942 (N_4942,N_1640,N_2527);
nor U4943 (N_4943,N_2732,N_1500);
and U4944 (N_4944,N_876,N_1321);
nand U4945 (N_4945,N_262,N_2497);
nor U4946 (N_4946,N_1017,N_538);
nor U4947 (N_4947,N_2581,N_121);
xnor U4948 (N_4948,N_888,N_2344);
xnor U4949 (N_4949,N_2066,N_2371);
nor U4950 (N_4950,N_794,N_1384);
xor U4951 (N_4951,N_14,N_1756);
xnor U4952 (N_4952,N_467,N_1878);
nand U4953 (N_4953,N_1500,N_1791);
or U4954 (N_4954,N_1140,N_1347);
or U4955 (N_4955,N_2568,N_1810);
or U4956 (N_4956,N_921,N_2410);
nor U4957 (N_4957,N_2194,N_469);
and U4958 (N_4958,N_516,N_2374);
nor U4959 (N_4959,N_1320,N_333);
nand U4960 (N_4960,N_1832,N_1538);
xor U4961 (N_4961,N_1336,N_2811);
xor U4962 (N_4962,N_1134,N_1602);
or U4963 (N_4963,N_1955,N_789);
and U4964 (N_4964,N_2313,N_2469);
or U4965 (N_4965,N_945,N_740);
or U4966 (N_4966,N_1435,N_1899);
or U4967 (N_4967,N_503,N_384);
xor U4968 (N_4968,N_1288,N_2831);
or U4969 (N_4969,N_1202,N_575);
or U4970 (N_4970,N_2427,N_3040);
nor U4971 (N_4971,N_2741,N_2703);
nand U4972 (N_4972,N_209,N_421);
nor U4973 (N_4973,N_519,N_1262);
or U4974 (N_4974,N_2640,N_612);
xor U4975 (N_4975,N_638,N_817);
xor U4976 (N_4976,N_1998,N_2490);
nor U4977 (N_4977,N_1950,N_1393);
nand U4978 (N_4978,N_965,N_2117);
and U4979 (N_4979,N_162,N_2836);
nor U4980 (N_4980,N_1674,N_573);
or U4981 (N_4981,N_790,N_1316);
nor U4982 (N_4982,N_2140,N_2157);
and U4983 (N_4983,N_2387,N_2266);
and U4984 (N_4984,N_2770,N_1202);
and U4985 (N_4985,N_2466,N_367);
nand U4986 (N_4986,N_2106,N_990);
and U4987 (N_4987,N_1478,N_2389);
and U4988 (N_4988,N_1069,N_1522);
and U4989 (N_4989,N_2174,N_2677);
nor U4990 (N_4990,N_1736,N_719);
nand U4991 (N_4991,N_822,N_3020);
or U4992 (N_4992,N_2349,N_2115);
and U4993 (N_4993,N_1547,N_1034);
xor U4994 (N_4994,N_2992,N_735);
and U4995 (N_4995,N_1746,N_2980);
xnor U4996 (N_4996,N_225,N_2210);
and U4997 (N_4997,N_1069,N_1704);
nor U4998 (N_4998,N_1314,N_1510);
nand U4999 (N_4999,N_1532,N_1551);
or U5000 (N_5000,N_3083,N_2510);
nor U5001 (N_5001,N_2504,N_1180);
or U5002 (N_5002,N_954,N_2310);
nor U5003 (N_5003,N_114,N_943);
xnor U5004 (N_5004,N_3057,N_2687);
nand U5005 (N_5005,N_1813,N_1248);
and U5006 (N_5006,N_2231,N_1008);
nor U5007 (N_5007,N_1660,N_2979);
and U5008 (N_5008,N_58,N_1414);
nor U5009 (N_5009,N_472,N_127);
nor U5010 (N_5010,N_1211,N_1603);
nor U5011 (N_5011,N_1303,N_998);
or U5012 (N_5012,N_1604,N_2364);
or U5013 (N_5013,N_481,N_2622);
and U5014 (N_5014,N_284,N_1972);
xnor U5015 (N_5015,N_3090,N_2946);
nor U5016 (N_5016,N_525,N_2335);
nor U5017 (N_5017,N_2537,N_697);
nor U5018 (N_5018,N_307,N_137);
nand U5019 (N_5019,N_1256,N_1001);
nand U5020 (N_5020,N_1696,N_2152);
nand U5021 (N_5021,N_1866,N_1802);
and U5022 (N_5022,N_2675,N_1553);
or U5023 (N_5023,N_706,N_382);
xor U5024 (N_5024,N_2853,N_1341);
and U5025 (N_5025,N_196,N_2535);
nand U5026 (N_5026,N_980,N_2775);
and U5027 (N_5027,N_331,N_884);
nor U5028 (N_5028,N_1240,N_2219);
xnor U5029 (N_5029,N_1790,N_3025);
nor U5030 (N_5030,N_356,N_2637);
and U5031 (N_5031,N_1634,N_2113);
or U5032 (N_5032,N_2984,N_1169);
nor U5033 (N_5033,N_2285,N_595);
nand U5034 (N_5034,N_1805,N_3060);
xnor U5035 (N_5035,N_311,N_1773);
xor U5036 (N_5036,N_566,N_432);
nand U5037 (N_5037,N_707,N_313);
and U5038 (N_5038,N_108,N_1223);
or U5039 (N_5039,N_2407,N_324);
xnor U5040 (N_5040,N_2385,N_2298);
or U5041 (N_5041,N_2310,N_2814);
xnor U5042 (N_5042,N_2393,N_1571);
or U5043 (N_5043,N_49,N_992);
or U5044 (N_5044,N_2649,N_2711);
and U5045 (N_5045,N_555,N_1656);
nand U5046 (N_5046,N_1515,N_2938);
or U5047 (N_5047,N_1479,N_2582);
nand U5048 (N_5048,N_2059,N_1719);
and U5049 (N_5049,N_1258,N_1273);
nor U5050 (N_5050,N_289,N_542);
and U5051 (N_5051,N_370,N_2499);
or U5052 (N_5052,N_1122,N_288);
nand U5053 (N_5053,N_701,N_559);
nand U5054 (N_5054,N_2249,N_2316);
nor U5055 (N_5055,N_320,N_1329);
or U5056 (N_5056,N_1409,N_1366);
nor U5057 (N_5057,N_3124,N_2915);
nand U5058 (N_5058,N_547,N_2826);
xor U5059 (N_5059,N_823,N_237);
and U5060 (N_5060,N_101,N_149);
or U5061 (N_5061,N_182,N_1007);
nor U5062 (N_5062,N_188,N_2941);
nor U5063 (N_5063,N_783,N_1290);
and U5064 (N_5064,N_2628,N_1465);
nand U5065 (N_5065,N_119,N_2705);
xor U5066 (N_5066,N_2538,N_1931);
xnor U5067 (N_5067,N_1840,N_469);
nor U5068 (N_5068,N_500,N_315);
or U5069 (N_5069,N_823,N_389);
nor U5070 (N_5070,N_908,N_62);
nand U5071 (N_5071,N_1715,N_2830);
or U5072 (N_5072,N_1986,N_2259);
and U5073 (N_5073,N_172,N_351);
nor U5074 (N_5074,N_1856,N_1172);
and U5075 (N_5075,N_902,N_1189);
and U5076 (N_5076,N_1093,N_3120);
and U5077 (N_5077,N_2851,N_2978);
xor U5078 (N_5078,N_672,N_2990);
and U5079 (N_5079,N_2947,N_2582);
and U5080 (N_5080,N_1083,N_1849);
nor U5081 (N_5081,N_2560,N_1316);
or U5082 (N_5082,N_112,N_370);
or U5083 (N_5083,N_2724,N_987);
nor U5084 (N_5084,N_1786,N_718);
and U5085 (N_5085,N_1874,N_300);
and U5086 (N_5086,N_2322,N_290);
nor U5087 (N_5087,N_39,N_574);
and U5088 (N_5088,N_2970,N_2400);
nand U5089 (N_5089,N_1079,N_1558);
nand U5090 (N_5090,N_388,N_2209);
nand U5091 (N_5091,N_1401,N_2412);
or U5092 (N_5092,N_1580,N_523);
xor U5093 (N_5093,N_638,N_889);
nor U5094 (N_5094,N_928,N_1767);
xor U5095 (N_5095,N_2174,N_1118);
nor U5096 (N_5096,N_630,N_216);
nor U5097 (N_5097,N_2530,N_304);
nor U5098 (N_5098,N_1893,N_1465);
xor U5099 (N_5099,N_2444,N_1605);
nor U5100 (N_5100,N_2973,N_427);
nor U5101 (N_5101,N_2264,N_2701);
nand U5102 (N_5102,N_1520,N_556);
and U5103 (N_5103,N_2637,N_2521);
xnor U5104 (N_5104,N_2384,N_1890);
xor U5105 (N_5105,N_1178,N_900);
nor U5106 (N_5106,N_1280,N_1275);
nor U5107 (N_5107,N_1385,N_2451);
xnor U5108 (N_5108,N_1825,N_1403);
or U5109 (N_5109,N_755,N_1040);
or U5110 (N_5110,N_2565,N_1525);
nor U5111 (N_5111,N_94,N_759);
xor U5112 (N_5112,N_1620,N_1084);
or U5113 (N_5113,N_2351,N_628);
xor U5114 (N_5114,N_3075,N_2641);
nor U5115 (N_5115,N_740,N_1462);
or U5116 (N_5116,N_319,N_1877);
and U5117 (N_5117,N_844,N_1080);
nand U5118 (N_5118,N_1520,N_2070);
nand U5119 (N_5119,N_2903,N_1750);
and U5120 (N_5120,N_1858,N_3041);
nand U5121 (N_5121,N_2257,N_116);
and U5122 (N_5122,N_2310,N_605);
and U5123 (N_5123,N_2994,N_499);
xnor U5124 (N_5124,N_300,N_245);
nand U5125 (N_5125,N_2487,N_565);
xor U5126 (N_5126,N_3045,N_2083);
or U5127 (N_5127,N_1975,N_2217);
or U5128 (N_5128,N_991,N_1551);
or U5129 (N_5129,N_1106,N_217);
and U5130 (N_5130,N_637,N_1701);
xnor U5131 (N_5131,N_1099,N_2056);
or U5132 (N_5132,N_176,N_2074);
and U5133 (N_5133,N_1789,N_43);
and U5134 (N_5134,N_2543,N_3010);
nor U5135 (N_5135,N_2970,N_2395);
or U5136 (N_5136,N_33,N_2371);
nor U5137 (N_5137,N_3047,N_1356);
and U5138 (N_5138,N_703,N_2329);
and U5139 (N_5139,N_2279,N_2957);
nor U5140 (N_5140,N_2172,N_1908);
xor U5141 (N_5141,N_2557,N_1656);
nor U5142 (N_5142,N_138,N_1669);
xnor U5143 (N_5143,N_260,N_1882);
nor U5144 (N_5144,N_2332,N_840);
xor U5145 (N_5145,N_2754,N_2280);
nand U5146 (N_5146,N_2437,N_1456);
nand U5147 (N_5147,N_1330,N_1526);
and U5148 (N_5148,N_2397,N_412);
nor U5149 (N_5149,N_178,N_2176);
xor U5150 (N_5150,N_207,N_2653);
or U5151 (N_5151,N_1562,N_2338);
nand U5152 (N_5152,N_2181,N_1366);
nor U5153 (N_5153,N_2608,N_1410);
nor U5154 (N_5154,N_2616,N_1365);
or U5155 (N_5155,N_2724,N_1375);
nand U5156 (N_5156,N_1923,N_2210);
nand U5157 (N_5157,N_1065,N_1871);
and U5158 (N_5158,N_715,N_47);
or U5159 (N_5159,N_2824,N_2904);
nand U5160 (N_5160,N_1318,N_850);
nor U5161 (N_5161,N_1861,N_339);
xor U5162 (N_5162,N_940,N_2818);
and U5163 (N_5163,N_212,N_1939);
nor U5164 (N_5164,N_56,N_345);
nor U5165 (N_5165,N_2543,N_2507);
nor U5166 (N_5166,N_1654,N_31);
or U5167 (N_5167,N_2668,N_1312);
or U5168 (N_5168,N_1507,N_2884);
or U5169 (N_5169,N_1314,N_1723);
nand U5170 (N_5170,N_261,N_312);
nand U5171 (N_5171,N_3080,N_1330);
nor U5172 (N_5172,N_1008,N_1524);
xor U5173 (N_5173,N_1270,N_1715);
nand U5174 (N_5174,N_240,N_1399);
or U5175 (N_5175,N_1093,N_1172);
or U5176 (N_5176,N_212,N_2696);
nand U5177 (N_5177,N_3099,N_735);
nor U5178 (N_5178,N_2661,N_247);
nor U5179 (N_5179,N_2869,N_548);
nor U5180 (N_5180,N_1845,N_2527);
nor U5181 (N_5181,N_2083,N_1539);
nand U5182 (N_5182,N_917,N_1694);
nand U5183 (N_5183,N_2592,N_1754);
or U5184 (N_5184,N_845,N_441);
xor U5185 (N_5185,N_163,N_2516);
xnor U5186 (N_5186,N_2838,N_1898);
nor U5187 (N_5187,N_20,N_1440);
xor U5188 (N_5188,N_3093,N_1457);
nor U5189 (N_5189,N_2988,N_2449);
and U5190 (N_5190,N_1642,N_1331);
xnor U5191 (N_5191,N_826,N_453);
nand U5192 (N_5192,N_511,N_1630);
and U5193 (N_5193,N_1317,N_750);
xnor U5194 (N_5194,N_1117,N_860);
or U5195 (N_5195,N_2418,N_58);
nand U5196 (N_5196,N_2372,N_1891);
or U5197 (N_5197,N_1894,N_3053);
or U5198 (N_5198,N_1992,N_2757);
nand U5199 (N_5199,N_456,N_1429);
nand U5200 (N_5200,N_19,N_1787);
nor U5201 (N_5201,N_1416,N_695);
and U5202 (N_5202,N_689,N_1861);
and U5203 (N_5203,N_56,N_496);
nand U5204 (N_5204,N_2871,N_280);
or U5205 (N_5205,N_2987,N_1754);
xnor U5206 (N_5206,N_2114,N_2794);
and U5207 (N_5207,N_2305,N_1752);
nor U5208 (N_5208,N_1926,N_2440);
or U5209 (N_5209,N_1325,N_807);
xor U5210 (N_5210,N_817,N_1633);
nor U5211 (N_5211,N_375,N_2100);
nand U5212 (N_5212,N_1667,N_3054);
nor U5213 (N_5213,N_1877,N_1194);
and U5214 (N_5214,N_2574,N_1154);
xor U5215 (N_5215,N_2252,N_1757);
xnor U5216 (N_5216,N_383,N_1470);
and U5217 (N_5217,N_2476,N_1177);
nand U5218 (N_5218,N_2956,N_1796);
or U5219 (N_5219,N_2253,N_841);
nor U5220 (N_5220,N_1256,N_129);
or U5221 (N_5221,N_1021,N_919);
nor U5222 (N_5222,N_213,N_61);
nand U5223 (N_5223,N_2004,N_2748);
xnor U5224 (N_5224,N_1827,N_1157);
and U5225 (N_5225,N_2308,N_2101);
nand U5226 (N_5226,N_2850,N_274);
nand U5227 (N_5227,N_2956,N_702);
xor U5228 (N_5228,N_2375,N_1865);
and U5229 (N_5229,N_105,N_1786);
nor U5230 (N_5230,N_741,N_1237);
or U5231 (N_5231,N_1614,N_1121);
or U5232 (N_5232,N_782,N_2912);
nor U5233 (N_5233,N_2662,N_2456);
nor U5234 (N_5234,N_1662,N_121);
or U5235 (N_5235,N_1515,N_604);
xnor U5236 (N_5236,N_2319,N_2141);
nor U5237 (N_5237,N_1367,N_994);
xor U5238 (N_5238,N_2677,N_1923);
or U5239 (N_5239,N_12,N_2547);
or U5240 (N_5240,N_3017,N_2755);
and U5241 (N_5241,N_1596,N_2824);
nand U5242 (N_5242,N_817,N_2605);
or U5243 (N_5243,N_2609,N_1662);
or U5244 (N_5244,N_59,N_349);
xor U5245 (N_5245,N_2799,N_1952);
nand U5246 (N_5246,N_2064,N_1280);
or U5247 (N_5247,N_419,N_129);
nand U5248 (N_5248,N_3085,N_2903);
or U5249 (N_5249,N_923,N_733);
and U5250 (N_5250,N_2457,N_1514);
nand U5251 (N_5251,N_3097,N_2021);
and U5252 (N_5252,N_1167,N_2300);
xnor U5253 (N_5253,N_2819,N_2684);
nand U5254 (N_5254,N_2644,N_2121);
and U5255 (N_5255,N_1808,N_2676);
nand U5256 (N_5256,N_2324,N_1716);
or U5257 (N_5257,N_41,N_3002);
nand U5258 (N_5258,N_3064,N_974);
xnor U5259 (N_5259,N_1008,N_2706);
and U5260 (N_5260,N_1137,N_2975);
nand U5261 (N_5261,N_1372,N_2631);
xnor U5262 (N_5262,N_3112,N_939);
or U5263 (N_5263,N_2918,N_3122);
or U5264 (N_5264,N_1668,N_102);
nand U5265 (N_5265,N_1991,N_975);
xor U5266 (N_5266,N_480,N_2144);
and U5267 (N_5267,N_1885,N_1520);
xor U5268 (N_5268,N_2296,N_15);
xor U5269 (N_5269,N_1237,N_266);
nor U5270 (N_5270,N_2913,N_2862);
nand U5271 (N_5271,N_474,N_2027);
nand U5272 (N_5272,N_88,N_1216);
nand U5273 (N_5273,N_503,N_195);
nor U5274 (N_5274,N_813,N_1625);
and U5275 (N_5275,N_2398,N_2676);
xor U5276 (N_5276,N_645,N_456);
nor U5277 (N_5277,N_2245,N_810);
or U5278 (N_5278,N_1182,N_1549);
or U5279 (N_5279,N_2095,N_2906);
or U5280 (N_5280,N_1252,N_2555);
or U5281 (N_5281,N_725,N_2213);
or U5282 (N_5282,N_2958,N_858);
nand U5283 (N_5283,N_2865,N_2368);
or U5284 (N_5284,N_2553,N_2861);
nor U5285 (N_5285,N_1494,N_1698);
nor U5286 (N_5286,N_77,N_1592);
nand U5287 (N_5287,N_3092,N_2265);
nor U5288 (N_5288,N_1188,N_2694);
or U5289 (N_5289,N_2080,N_1576);
or U5290 (N_5290,N_1171,N_2950);
nand U5291 (N_5291,N_1281,N_1491);
nand U5292 (N_5292,N_1693,N_679);
and U5293 (N_5293,N_1647,N_2525);
and U5294 (N_5294,N_2894,N_2327);
and U5295 (N_5295,N_759,N_687);
and U5296 (N_5296,N_1616,N_865);
xor U5297 (N_5297,N_2741,N_30);
xor U5298 (N_5298,N_2906,N_1279);
xor U5299 (N_5299,N_287,N_1166);
or U5300 (N_5300,N_561,N_2624);
or U5301 (N_5301,N_84,N_1512);
nor U5302 (N_5302,N_892,N_737);
nor U5303 (N_5303,N_956,N_1662);
xor U5304 (N_5304,N_2710,N_733);
xnor U5305 (N_5305,N_2129,N_1852);
or U5306 (N_5306,N_1676,N_268);
or U5307 (N_5307,N_1628,N_3019);
xor U5308 (N_5308,N_2925,N_2888);
xor U5309 (N_5309,N_525,N_1263);
or U5310 (N_5310,N_125,N_545);
nor U5311 (N_5311,N_3114,N_1714);
and U5312 (N_5312,N_1360,N_1974);
or U5313 (N_5313,N_263,N_251);
nand U5314 (N_5314,N_1275,N_1732);
or U5315 (N_5315,N_2123,N_2938);
nand U5316 (N_5316,N_281,N_3023);
nand U5317 (N_5317,N_613,N_1314);
nand U5318 (N_5318,N_2235,N_862);
nor U5319 (N_5319,N_1296,N_632);
nand U5320 (N_5320,N_869,N_2230);
and U5321 (N_5321,N_2723,N_2756);
xor U5322 (N_5322,N_93,N_2509);
nand U5323 (N_5323,N_1318,N_881);
or U5324 (N_5324,N_3086,N_2767);
nor U5325 (N_5325,N_647,N_1746);
and U5326 (N_5326,N_192,N_944);
nand U5327 (N_5327,N_1455,N_505);
xnor U5328 (N_5328,N_2039,N_2537);
nor U5329 (N_5329,N_1540,N_1383);
and U5330 (N_5330,N_126,N_199);
xnor U5331 (N_5331,N_1405,N_2607);
nand U5332 (N_5332,N_1787,N_2363);
and U5333 (N_5333,N_972,N_2788);
xor U5334 (N_5334,N_1183,N_1584);
and U5335 (N_5335,N_305,N_2538);
or U5336 (N_5336,N_686,N_1640);
xnor U5337 (N_5337,N_1767,N_2486);
and U5338 (N_5338,N_2864,N_134);
nor U5339 (N_5339,N_2384,N_1270);
xor U5340 (N_5340,N_2732,N_2806);
nor U5341 (N_5341,N_1506,N_38);
or U5342 (N_5342,N_100,N_362);
nand U5343 (N_5343,N_2676,N_2113);
nand U5344 (N_5344,N_1722,N_1375);
nand U5345 (N_5345,N_1938,N_2313);
xor U5346 (N_5346,N_1390,N_1729);
xor U5347 (N_5347,N_309,N_1468);
nor U5348 (N_5348,N_1191,N_1113);
nand U5349 (N_5349,N_2904,N_2730);
nor U5350 (N_5350,N_2829,N_2921);
or U5351 (N_5351,N_2368,N_2264);
nor U5352 (N_5352,N_44,N_154);
xor U5353 (N_5353,N_510,N_1931);
nand U5354 (N_5354,N_2895,N_676);
or U5355 (N_5355,N_2911,N_333);
nor U5356 (N_5356,N_1886,N_1957);
nor U5357 (N_5357,N_2491,N_2806);
xnor U5358 (N_5358,N_1337,N_1394);
nor U5359 (N_5359,N_1821,N_380);
nand U5360 (N_5360,N_1075,N_1564);
and U5361 (N_5361,N_1235,N_2609);
xnor U5362 (N_5362,N_3013,N_1277);
nor U5363 (N_5363,N_409,N_942);
or U5364 (N_5364,N_663,N_1066);
and U5365 (N_5365,N_1753,N_1600);
and U5366 (N_5366,N_1231,N_2555);
or U5367 (N_5367,N_569,N_680);
and U5368 (N_5368,N_2429,N_2038);
xnor U5369 (N_5369,N_263,N_2442);
nor U5370 (N_5370,N_637,N_833);
and U5371 (N_5371,N_2097,N_1167);
or U5372 (N_5372,N_1498,N_2694);
and U5373 (N_5373,N_542,N_2453);
and U5374 (N_5374,N_129,N_168);
nand U5375 (N_5375,N_931,N_1866);
nand U5376 (N_5376,N_404,N_435);
or U5377 (N_5377,N_159,N_2634);
nor U5378 (N_5378,N_960,N_831);
nand U5379 (N_5379,N_745,N_2100);
and U5380 (N_5380,N_2581,N_1362);
nor U5381 (N_5381,N_1131,N_118);
nor U5382 (N_5382,N_2946,N_2649);
and U5383 (N_5383,N_526,N_2906);
nor U5384 (N_5384,N_1210,N_2174);
nor U5385 (N_5385,N_2784,N_897);
nand U5386 (N_5386,N_764,N_2153);
or U5387 (N_5387,N_1670,N_1045);
nor U5388 (N_5388,N_1392,N_1868);
nor U5389 (N_5389,N_2037,N_171);
nand U5390 (N_5390,N_866,N_1928);
and U5391 (N_5391,N_2690,N_792);
and U5392 (N_5392,N_2214,N_730);
nor U5393 (N_5393,N_2257,N_452);
or U5394 (N_5394,N_2172,N_1286);
nor U5395 (N_5395,N_1554,N_1814);
nor U5396 (N_5396,N_2068,N_1184);
and U5397 (N_5397,N_112,N_309);
nand U5398 (N_5398,N_465,N_2527);
or U5399 (N_5399,N_585,N_591);
nor U5400 (N_5400,N_2046,N_2125);
and U5401 (N_5401,N_1296,N_2148);
nand U5402 (N_5402,N_2125,N_439);
nor U5403 (N_5403,N_2682,N_465);
or U5404 (N_5404,N_836,N_2494);
and U5405 (N_5405,N_3097,N_1688);
nor U5406 (N_5406,N_164,N_2126);
xor U5407 (N_5407,N_1388,N_448);
or U5408 (N_5408,N_2747,N_107);
and U5409 (N_5409,N_2970,N_176);
nand U5410 (N_5410,N_939,N_274);
or U5411 (N_5411,N_3044,N_2809);
xor U5412 (N_5412,N_518,N_2367);
nor U5413 (N_5413,N_1399,N_2612);
nor U5414 (N_5414,N_2779,N_2105);
nor U5415 (N_5415,N_377,N_2771);
and U5416 (N_5416,N_2390,N_2693);
xor U5417 (N_5417,N_758,N_539);
nand U5418 (N_5418,N_1025,N_1386);
nand U5419 (N_5419,N_340,N_704);
xnor U5420 (N_5420,N_1211,N_2050);
nand U5421 (N_5421,N_2045,N_2178);
nand U5422 (N_5422,N_2470,N_2100);
xor U5423 (N_5423,N_2030,N_375);
nor U5424 (N_5424,N_2890,N_1270);
xnor U5425 (N_5425,N_1706,N_443);
nand U5426 (N_5426,N_1370,N_1460);
xnor U5427 (N_5427,N_205,N_134);
nor U5428 (N_5428,N_3088,N_2561);
nor U5429 (N_5429,N_1320,N_2370);
xor U5430 (N_5430,N_2906,N_1325);
xnor U5431 (N_5431,N_649,N_1244);
or U5432 (N_5432,N_3069,N_1567);
nor U5433 (N_5433,N_1498,N_2907);
xnor U5434 (N_5434,N_600,N_687);
nor U5435 (N_5435,N_2663,N_1381);
nand U5436 (N_5436,N_815,N_2777);
nor U5437 (N_5437,N_888,N_1240);
nor U5438 (N_5438,N_1162,N_2640);
xnor U5439 (N_5439,N_1268,N_2321);
and U5440 (N_5440,N_1008,N_485);
nor U5441 (N_5441,N_1107,N_1867);
or U5442 (N_5442,N_759,N_450);
and U5443 (N_5443,N_117,N_2368);
xnor U5444 (N_5444,N_579,N_525);
nor U5445 (N_5445,N_2995,N_2266);
and U5446 (N_5446,N_1531,N_925);
nand U5447 (N_5447,N_318,N_694);
nor U5448 (N_5448,N_2645,N_2523);
nand U5449 (N_5449,N_331,N_535);
xor U5450 (N_5450,N_1213,N_2871);
nor U5451 (N_5451,N_90,N_1885);
nor U5452 (N_5452,N_1,N_617);
xnor U5453 (N_5453,N_1167,N_2804);
or U5454 (N_5454,N_1761,N_1409);
xnor U5455 (N_5455,N_2628,N_1412);
nand U5456 (N_5456,N_1624,N_1001);
and U5457 (N_5457,N_990,N_2071);
nor U5458 (N_5458,N_1338,N_273);
xnor U5459 (N_5459,N_1786,N_1780);
or U5460 (N_5460,N_3021,N_2752);
nand U5461 (N_5461,N_724,N_2100);
and U5462 (N_5462,N_527,N_1652);
xnor U5463 (N_5463,N_310,N_1591);
or U5464 (N_5464,N_1508,N_2361);
nor U5465 (N_5465,N_2607,N_653);
and U5466 (N_5466,N_1295,N_783);
nor U5467 (N_5467,N_1624,N_610);
xor U5468 (N_5468,N_2026,N_1978);
xnor U5469 (N_5469,N_1939,N_2988);
nand U5470 (N_5470,N_1202,N_1767);
nor U5471 (N_5471,N_2490,N_1195);
and U5472 (N_5472,N_2066,N_2159);
and U5473 (N_5473,N_872,N_2646);
nor U5474 (N_5474,N_635,N_33);
nand U5475 (N_5475,N_55,N_2924);
xor U5476 (N_5476,N_2728,N_2262);
or U5477 (N_5477,N_2668,N_121);
nand U5478 (N_5478,N_1159,N_1804);
or U5479 (N_5479,N_1310,N_81);
nand U5480 (N_5480,N_2285,N_1879);
xnor U5481 (N_5481,N_2545,N_2290);
or U5482 (N_5482,N_923,N_2409);
and U5483 (N_5483,N_2029,N_2755);
or U5484 (N_5484,N_1523,N_1180);
nand U5485 (N_5485,N_249,N_297);
nand U5486 (N_5486,N_2297,N_2559);
nor U5487 (N_5487,N_2799,N_1267);
nand U5488 (N_5488,N_90,N_1321);
nor U5489 (N_5489,N_1960,N_1134);
or U5490 (N_5490,N_301,N_1920);
or U5491 (N_5491,N_647,N_876);
and U5492 (N_5492,N_267,N_528);
or U5493 (N_5493,N_907,N_2993);
and U5494 (N_5494,N_2770,N_2042);
or U5495 (N_5495,N_1044,N_642);
or U5496 (N_5496,N_645,N_2291);
xnor U5497 (N_5497,N_1079,N_86);
or U5498 (N_5498,N_846,N_2441);
and U5499 (N_5499,N_750,N_1644);
nand U5500 (N_5500,N_1586,N_201);
nand U5501 (N_5501,N_802,N_2760);
nor U5502 (N_5502,N_2076,N_2902);
nor U5503 (N_5503,N_2321,N_1244);
xnor U5504 (N_5504,N_2823,N_2162);
nand U5505 (N_5505,N_2924,N_404);
xor U5506 (N_5506,N_2693,N_342);
or U5507 (N_5507,N_2672,N_1413);
or U5508 (N_5508,N_693,N_1454);
nor U5509 (N_5509,N_1077,N_2210);
nor U5510 (N_5510,N_624,N_2403);
and U5511 (N_5511,N_1612,N_939);
or U5512 (N_5512,N_447,N_1450);
xor U5513 (N_5513,N_162,N_354);
nand U5514 (N_5514,N_2892,N_610);
nand U5515 (N_5515,N_2244,N_3052);
or U5516 (N_5516,N_1583,N_386);
nor U5517 (N_5517,N_2164,N_2409);
nand U5518 (N_5518,N_3099,N_1762);
nor U5519 (N_5519,N_1888,N_542);
xnor U5520 (N_5520,N_1981,N_1023);
nand U5521 (N_5521,N_113,N_1143);
xor U5522 (N_5522,N_366,N_2588);
and U5523 (N_5523,N_2893,N_2373);
and U5524 (N_5524,N_2376,N_1238);
or U5525 (N_5525,N_1532,N_2411);
nand U5526 (N_5526,N_2027,N_207);
xor U5527 (N_5527,N_1160,N_2790);
or U5528 (N_5528,N_1678,N_142);
xnor U5529 (N_5529,N_2835,N_85);
and U5530 (N_5530,N_1479,N_2640);
xnor U5531 (N_5531,N_2298,N_2091);
nand U5532 (N_5532,N_286,N_1601);
or U5533 (N_5533,N_2862,N_3109);
and U5534 (N_5534,N_1230,N_1959);
nor U5535 (N_5535,N_327,N_2582);
nand U5536 (N_5536,N_1454,N_777);
and U5537 (N_5537,N_1514,N_1035);
and U5538 (N_5538,N_3099,N_1345);
nand U5539 (N_5539,N_2548,N_3049);
nand U5540 (N_5540,N_2671,N_548);
xor U5541 (N_5541,N_297,N_1452);
xor U5542 (N_5542,N_383,N_120);
or U5543 (N_5543,N_634,N_1628);
or U5544 (N_5544,N_3090,N_2711);
or U5545 (N_5545,N_2967,N_1511);
xnor U5546 (N_5546,N_2061,N_618);
xor U5547 (N_5547,N_2986,N_2310);
nand U5548 (N_5548,N_2212,N_2932);
or U5549 (N_5549,N_146,N_1857);
xnor U5550 (N_5550,N_402,N_1083);
and U5551 (N_5551,N_23,N_253);
xnor U5552 (N_5552,N_3111,N_2110);
or U5553 (N_5553,N_585,N_2302);
xnor U5554 (N_5554,N_1532,N_2487);
and U5555 (N_5555,N_1334,N_2536);
nand U5556 (N_5556,N_293,N_1527);
or U5557 (N_5557,N_1648,N_2999);
and U5558 (N_5558,N_1488,N_789);
and U5559 (N_5559,N_2959,N_3122);
nor U5560 (N_5560,N_1190,N_910);
and U5561 (N_5561,N_195,N_2946);
xnor U5562 (N_5562,N_2540,N_1292);
nand U5563 (N_5563,N_142,N_126);
nand U5564 (N_5564,N_717,N_1622);
nor U5565 (N_5565,N_679,N_2577);
or U5566 (N_5566,N_1926,N_1999);
xor U5567 (N_5567,N_2399,N_2941);
xor U5568 (N_5568,N_2217,N_229);
or U5569 (N_5569,N_2071,N_2879);
and U5570 (N_5570,N_1034,N_2577);
xnor U5571 (N_5571,N_104,N_1918);
and U5572 (N_5572,N_667,N_904);
and U5573 (N_5573,N_440,N_345);
nor U5574 (N_5574,N_571,N_2496);
xor U5575 (N_5575,N_1171,N_2158);
nor U5576 (N_5576,N_2767,N_3011);
xnor U5577 (N_5577,N_163,N_1048);
xor U5578 (N_5578,N_2831,N_2064);
and U5579 (N_5579,N_361,N_933);
or U5580 (N_5580,N_2832,N_3005);
nand U5581 (N_5581,N_1168,N_672);
xnor U5582 (N_5582,N_279,N_299);
nor U5583 (N_5583,N_2716,N_518);
and U5584 (N_5584,N_2294,N_883);
xnor U5585 (N_5585,N_1526,N_417);
xnor U5586 (N_5586,N_518,N_602);
nand U5587 (N_5587,N_2664,N_836);
or U5588 (N_5588,N_3068,N_1265);
xnor U5589 (N_5589,N_119,N_2677);
and U5590 (N_5590,N_2762,N_911);
and U5591 (N_5591,N_83,N_2365);
and U5592 (N_5592,N_1597,N_1055);
and U5593 (N_5593,N_403,N_2890);
nor U5594 (N_5594,N_2770,N_13);
and U5595 (N_5595,N_1465,N_1495);
and U5596 (N_5596,N_778,N_238);
or U5597 (N_5597,N_1793,N_2158);
or U5598 (N_5598,N_2556,N_2575);
xnor U5599 (N_5599,N_47,N_714);
or U5600 (N_5600,N_578,N_1509);
or U5601 (N_5601,N_2556,N_756);
nor U5602 (N_5602,N_1994,N_2962);
xnor U5603 (N_5603,N_378,N_682);
nand U5604 (N_5604,N_1919,N_2022);
or U5605 (N_5605,N_1322,N_2504);
nor U5606 (N_5606,N_1919,N_883);
xnor U5607 (N_5607,N_1865,N_2300);
nor U5608 (N_5608,N_2270,N_2695);
and U5609 (N_5609,N_986,N_444);
nor U5610 (N_5610,N_569,N_1809);
nand U5611 (N_5611,N_488,N_2110);
nand U5612 (N_5612,N_608,N_1676);
xor U5613 (N_5613,N_281,N_1368);
nand U5614 (N_5614,N_452,N_1188);
or U5615 (N_5615,N_1007,N_3109);
and U5616 (N_5616,N_1539,N_3037);
nand U5617 (N_5617,N_283,N_3098);
nor U5618 (N_5618,N_839,N_2718);
and U5619 (N_5619,N_1088,N_1092);
nor U5620 (N_5620,N_1429,N_1393);
and U5621 (N_5621,N_2604,N_1788);
nor U5622 (N_5622,N_2811,N_1931);
xnor U5623 (N_5623,N_1137,N_2254);
and U5624 (N_5624,N_200,N_1371);
nand U5625 (N_5625,N_182,N_2196);
or U5626 (N_5626,N_369,N_2373);
xnor U5627 (N_5627,N_1075,N_2574);
nor U5628 (N_5628,N_2343,N_1775);
xor U5629 (N_5629,N_1701,N_1783);
xor U5630 (N_5630,N_2370,N_997);
and U5631 (N_5631,N_1251,N_2901);
xnor U5632 (N_5632,N_573,N_885);
xnor U5633 (N_5633,N_1913,N_2130);
and U5634 (N_5634,N_1843,N_2321);
and U5635 (N_5635,N_2452,N_1305);
and U5636 (N_5636,N_52,N_1640);
nor U5637 (N_5637,N_245,N_830);
and U5638 (N_5638,N_729,N_2467);
nand U5639 (N_5639,N_1224,N_2661);
xor U5640 (N_5640,N_777,N_1971);
xor U5641 (N_5641,N_18,N_937);
xnor U5642 (N_5642,N_1961,N_1951);
nand U5643 (N_5643,N_1667,N_1137);
xor U5644 (N_5644,N_1238,N_1034);
and U5645 (N_5645,N_1194,N_2049);
xnor U5646 (N_5646,N_1500,N_667);
xnor U5647 (N_5647,N_140,N_2212);
and U5648 (N_5648,N_2420,N_2583);
xnor U5649 (N_5649,N_213,N_2458);
xnor U5650 (N_5650,N_3043,N_1925);
nor U5651 (N_5651,N_344,N_2498);
or U5652 (N_5652,N_1678,N_2595);
nand U5653 (N_5653,N_1313,N_1462);
xnor U5654 (N_5654,N_1990,N_2129);
and U5655 (N_5655,N_1915,N_1672);
or U5656 (N_5656,N_1370,N_780);
nor U5657 (N_5657,N_1543,N_2656);
xnor U5658 (N_5658,N_2681,N_429);
nand U5659 (N_5659,N_1950,N_169);
nand U5660 (N_5660,N_2531,N_724);
or U5661 (N_5661,N_1546,N_1475);
and U5662 (N_5662,N_1525,N_2969);
and U5663 (N_5663,N_2079,N_1370);
xnor U5664 (N_5664,N_588,N_1223);
xnor U5665 (N_5665,N_1192,N_1427);
xnor U5666 (N_5666,N_1000,N_1400);
nor U5667 (N_5667,N_2080,N_2241);
and U5668 (N_5668,N_848,N_3107);
xnor U5669 (N_5669,N_1024,N_2080);
and U5670 (N_5670,N_2665,N_2911);
or U5671 (N_5671,N_2015,N_2829);
nand U5672 (N_5672,N_1510,N_2197);
or U5673 (N_5673,N_1913,N_97);
xnor U5674 (N_5674,N_131,N_872);
nand U5675 (N_5675,N_38,N_948);
or U5676 (N_5676,N_2249,N_607);
nor U5677 (N_5677,N_2312,N_615);
or U5678 (N_5678,N_1476,N_1845);
or U5679 (N_5679,N_2569,N_1614);
nand U5680 (N_5680,N_2992,N_3098);
and U5681 (N_5681,N_741,N_865);
xnor U5682 (N_5682,N_2669,N_2885);
nor U5683 (N_5683,N_990,N_1700);
nand U5684 (N_5684,N_200,N_961);
nand U5685 (N_5685,N_2557,N_2871);
xor U5686 (N_5686,N_2321,N_2216);
and U5687 (N_5687,N_418,N_2060);
xor U5688 (N_5688,N_442,N_112);
nand U5689 (N_5689,N_564,N_60);
nor U5690 (N_5690,N_2177,N_439);
or U5691 (N_5691,N_2369,N_2374);
nand U5692 (N_5692,N_2736,N_3010);
nand U5693 (N_5693,N_995,N_526);
and U5694 (N_5694,N_1449,N_2101);
or U5695 (N_5695,N_2283,N_2439);
or U5696 (N_5696,N_568,N_2186);
and U5697 (N_5697,N_640,N_490);
or U5698 (N_5698,N_2300,N_2637);
xnor U5699 (N_5699,N_979,N_2475);
xnor U5700 (N_5700,N_3001,N_1655);
nand U5701 (N_5701,N_1031,N_2535);
or U5702 (N_5702,N_2006,N_1596);
nand U5703 (N_5703,N_798,N_560);
nand U5704 (N_5704,N_1685,N_2904);
and U5705 (N_5705,N_1812,N_2400);
xnor U5706 (N_5706,N_2606,N_1754);
nand U5707 (N_5707,N_404,N_2426);
nor U5708 (N_5708,N_60,N_2949);
or U5709 (N_5709,N_757,N_1714);
nor U5710 (N_5710,N_1153,N_400);
nor U5711 (N_5711,N_2251,N_2764);
nand U5712 (N_5712,N_1349,N_29);
xnor U5713 (N_5713,N_2200,N_951);
xor U5714 (N_5714,N_2972,N_2484);
xnor U5715 (N_5715,N_2221,N_2244);
nor U5716 (N_5716,N_1353,N_1094);
xor U5717 (N_5717,N_2553,N_1824);
xor U5718 (N_5718,N_1276,N_1799);
nand U5719 (N_5719,N_750,N_180);
and U5720 (N_5720,N_1848,N_1423);
nand U5721 (N_5721,N_1018,N_1048);
and U5722 (N_5722,N_2861,N_234);
and U5723 (N_5723,N_1006,N_2259);
xor U5724 (N_5724,N_2270,N_1398);
xor U5725 (N_5725,N_1092,N_3111);
or U5726 (N_5726,N_2702,N_2557);
or U5727 (N_5727,N_951,N_2479);
nor U5728 (N_5728,N_2938,N_3097);
xor U5729 (N_5729,N_1005,N_849);
and U5730 (N_5730,N_1374,N_2982);
nor U5731 (N_5731,N_1484,N_420);
and U5732 (N_5732,N_1968,N_2774);
and U5733 (N_5733,N_2505,N_1461);
or U5734 (N_5734,N_2192,N_554);
and U5735 (N_5735,N_2230,N_729);
nor U5736 (N_5736,N_728,N_1455);
nand U5737 (N_5737,N_2677,N_34);
xnor U5738 (N_5738,N_2111,N_1225);
nor U5739 (N_5739,N_2738,N_565);
nand U5740 (N_5740,N_550,N_2301);
nor U5741 (N_5741,N_363,N_2333);
nand U5742 (N_5742,N_503,N_2376);
nand U5743 (N_5743,N_2176,N_2860);
or U5744 (N_5744,N_2724,N_1208);
or U5745 (N_5745,N_777,N_1383);
and U5746 (N_5746,N_3031,N_2846);
nor U5747 (N_5747,N_2351,N_1426);
or U5748 (N_5748,N_2558,N_1619);
xor U5749 (N_5749,N_490,N_3056);
or U5750 (N_5750,N_84,N_2885);
and U5751 (N_5751,N_2731,N_858);
xnor U5752 (N_5752,N_2570,N_1798);
or U5753 (N_5753,N_258,N_16);
and U5754 (N_5754,N_735,N_2411);
nor U5755 (N_5755,N_1163,N_1746);
nand U5756 (N_5756,N_684,N_1110);
nor U5757 (N_5757,N_2200,N_2693);
xor U5758 (N_5758,N_1258,N_2316);
or U5759 (N_5759,N_2144,N_449);
nor U5760 (N_5760,N_208,N_2514);
nand U5761 (N_5761,N_1608,N_630);
nand U5762 (N_5762,N_1000,N_2354);
or U5763 (N_5763,N_1359,N_1360);
nand U5764 (N_5764,N_1224,N_549);
nor U5765 (N_5765,N_1514,N_2144);
nor U5766 (N_5766,N_735,N_2947);
or U5767 (N_5767,N_2533,N_236);
xnor U5768 (N_5768,N_1335,N_1808);
xor U5769 (N_5769,N_2995,N_2064);
nor U5770 (N_5770,N_2718,N_2810);
nor U5771 (N_5771,N_2366,N_1007);
xnor U5772 (N_5772,N_2347,N_136);
or U5773 (N_5773,N_2779,N_2417);
and U5774 (N_5774,N_2966,N_838);
and U5775 (N_5775,N_540,N_88);
and U5776 (N_5776,N_2528,N_2425);
or U5777 (N_5777,N_167,N_608);
or U5778 (N_5778,N_342,N_2003);
nand U5779 (N_5779,N_2422,N_1835);
or U5780 (N_5780,N_641,N_2543);
or U5781 (N_5781,N_1989,N_163);
nand U5782 (N_5782,N_1112,N_2085);
and U5783 (N_5783,N_189,N_2356);
and U5784 (N_5784,N_642,N_529);
nand U5785 (N_5785,N_2848,N_1635);
and U5786 (N_5786,N_2128,N_2770);
xnor U5787 (N_5787,N_1811,N_134);
and U5788 (N_5788,N_2891,N_1044);
nor U5789 (N_5789,N_2107,N_1106);
nor U5790 (N_5790,N_1623,N_1803);
or U5791 (N_5791,N_1013,N_443);
nor U5792 (N_5792,N_3016,N_931);
nor U5793 (N_5793,N_1636,N_2183);
and U5794 (N_5794,N_815,N_166);
nand U5795 (N_5795,N_1015,N_1625);
xor U5796 (N_5796,N_1531,N_2719);
nor U5797 (N_5797,N_125,N_563);
and U5798 (N_5798,N_169,N_2718);
nor U5799 (N_5799,N_100,N_557);
xor U5800 (N_5800,N_1830,N_2762);
nor U5801 (N_5801,N_2650,N_2429);
and U5802 (N_5802,N_1361,N_1798);
and U5803 (N_5803,N_166,N_547);
nand U5804 (N_5804,N_681,N_2029);
nand U5805 (N_5805,N_811,N_1737);
and U5806 (N_5806,N_2699,N_2769);
nand U5807 (N_5807,N_2426,N_1938);
nor U5808 (N_5808,N_1081,N_3096);
or U5809 (N_5809,N_340,N_2838);
nor U5810 (N_5810,N_2542,N_2618);
xor U5811 (N_5811,N_1201,N_31);
nor U5812 (N_5812,N_385,N_1849);
nand U5813 (N_5813,N_2626,N_814);
nand U5814 (N_5814,N_3108,N_3073);
or U5815 (N_5815,N_1159,N_1127);
nor U5816 (N_5816,N_1863,N_2197);
xnor U5817 (N_5817,N_2363,N_1591);
nand U5818 (N_5818,N_2354,N_1954);
and U5819 (N_5819,N_2360,N_1266);
nor U5820 (N_5820,N_2857,N_162);
nor U5821 (N_5821,N_1924,N_71);
nor U5822 (N_5822,N_2797,N_1829);
nand U5823 (N_5823,N_1217,N_2283);
xnor U5824 (N_5824,N_912,N_962);
nand U5825 (N_5825,N_2955,N_1372);
xnor U5826 (N_5826,N_1705,N_1361);
nand U5827 (N_5827,N_1477,N_2486);
nand U5828 (N_5828,N_890,N_1936);
and U5829 (N_5829,N_2629,N_968);
or U5830 (N_5830,N_2076,N_598);
and U5831 (N_5831,N_1767,N_655);
or U5832 (N_5832,N_2766,N_2258);
and U5833 (N_5833,N_2991,N_48);
xnor U5834 (N_5834,N_1915,N_2062);
nor U5835 (N_5835,N_1140,N_1803);
nor U5836 (N_5836,N_618,N_2957);
xnor U5837 (N_5837,N_1897,N_726);
nor U5838 (N_5838,N_1075,N_1683);
or U5839 (N_5839,N_2095,N_107);
nand U5840 (N_5840,N_285,N_3040);
xnor U5841 (N_5841,N_799,N_2984);
or U5842 (N_5842,N_2441,N_515);
nand U5843 (N_5843,N_753,N_526);
and U5844 (N_5844,N_1711,N_2235);
nand U5845 (N_5845,N_2098,N_2176);
or U5846 (N_5846,N_273,N_1374);
or U5847 (N_5847,N_1074,N_2796);
nor U5848 (N_5848,N_1427,N_2792);
or U5849 (N_5849,N_2390,N_842);
and U5850 (N_5850,N_905,N_1142);
nand U5851 (N_5851,N_2011,N_2105);
nand U5852 (N_5852,N_2527,N_604);
and U5853 (N_5853,N_1992,N_503);
or U5854 (N_5854,N_241,N_1816);
nand U5855 (N_5855,N_2036,N_21);
or U5856 (N_5856,N_1017,N_2160);
nand U5857 (N_5857,N_2415,N_2845);
nand U5858 (N_5858,N_146,N_2439);
and U5859 (N_5859,N_2159,N_1917);
nor U5860 (N_5860,N_2794,N_2285);
and U5861 (N_5861,N_579,N_459);
xnor U5862 (N_5862,N_1246,N_1849);
xnor U5863 (N_5863,N_3076,N_416);
and U5864 (N_5864,N_838,N_937);
nor U5865 (N_5865,N_2824,N_3047);
nand U5866 (N_5866,N_2676,N_380);
or U5867 (N_5867,N_631,N_626);
nand U5868 (N_5868,N_708,N_2124);
and U5869 (N_5869,N_1041,N_695);
or U5870 (N_5870,N_986,N_1702);
nand U5871 (N_5871,N_3063,N_1471);
nand U5872 (N_5872,N_2004,N_2635);
nand U5873 (N_5873,N_1772,N_1184);
xnor U5874 (N_5874,N_111,N_1524);
and U5875 (N_5875,N_508,N_580);
xnor U5876 (N_5876,N_761,N_736);
xor U5877 (N_5877,N_651,N_214);
nor U5878 (N_5878,N_1613,N_22);
nor U5879 (N_5879,N_2360,N_74);
or U5880 (N_5880,N_1751,N_3049);
nand U5881 (N_5881,N_1912,N_1898);
or U5882 (N_5882,N_963,N_3121);
nand U5883 (N_5883,N_534,N_1339);
xnor U5884 (N_5884,N_2954,N_65);
nand U5885 (N_5885,N_1951,N_99);
or U5886 (N_5886,N_135,N_2698);
xor U5887 (N_5887,N_2469,N_2358);
xor U5888 (N_5888,N_1013,N_2462);
and U5889 (N_5889,N_1349,N_2104);
or U5890 (N_5890,N_2487,N_2003);
and U5891 (N_5891,N_494,N_1962);
and U5892 (N_5892,N_1760,N_1123);
nand U5893 (N_5893,N_916,N_2370);
nand U5894 (N_5894,N_903,N_2159);
nand U5895 (N_5895,N_1212,N_2819);
and U5896 (N_5896,N_3124,N_2856);
nand U5897 (N_5897,N_3104,N_856);
xnor U5898 (N_5898,N_2493,N_993);
nor U5899 (N_5899,N_765,N_1912);
nor U5900 (N_5900,N_1849,N_2409);
xnor U5901 (N_5901,N_1775,N_1564);
or U5902 (N_5902,N_2147,N_438);
xnor U5903 (N_5903,N_1151,N_2609);
xnor U5904 (N_5904,N_1507,N_525);
nand U5905 (N_5905,N_2002,N_129);
nor U5906 (N_5906,N_2251,N_923);
nand U5907 (N_5907,N_764,N_2210);
and U5908 (N_5908,N_668,N_254);
and U5909 (N_5909,N_2213,N_202);
or U5910 (N_5910,N_2667,N_2608);
xnor U5911 (N_5911,N_1125,N_2091);
and U5912 (N_5912,N_2364,N_2835);
or U5913 (N_5913,N_716,N_2428);
nor U5914 (N_5914,N_2414,N_1923);
nand U5915 (N_5915,N_1894,N_303);
xor U5916 (N_5916,N_1385,N_2474);
and U5917 (N_5917,N_963,N_1604);
or U5918 (N_5918,N_543,N_2528);
nor U5919 (N_5919,N_2076,N_2776);
xnor U5920 (N_5920,N_763,N_2251);
or U5921 (N_5921,N_9,N_522);
and U5922 (N_5922,N_2227,N_510);
and U5923 (N_5923,N_2613,N_2051);
xor U5924 (N_5924,N_2311,N_529);
and U5925 (N_5925,N_1420,N_1272);
xnor U5926 (N_5926,N_895,N_1574);
or U5927 (N_5927,N_520,N_738);
xor U5928 (N_5928,N_2492,N_134);
nor U5929 (N_5929,N_1549,N_3080);
and U5930 (N_5930,N_2119,N_1813);
nor U5931 (N_5931,N_943,N_2430);
nor U5932 (N_5932,N_2931,N_2091);
nand U5933 (N_5933,N_1958,N_2388);
xor U5934 (N_5934,N_1085,N_1472);
nor U5935 (N_5935,N_1882,N_2321);
nor U5936 (N_5936,N_994,N_1740);
xnor U5937 (N_5937,N_1339,N_1294);
or U5938 (N_5938,N_1595,N_265);
and U5939 (N_5939,N_2490,N_2700);
or U5940 (N_5940,N_1231,N_2251);
xor U5941 (N_5941,N_2659,N_349);
xor U5942 (N_5942,N_695,N_2285);
or U5943 (N_5943,N_1614,N_2805);
nor U5944 (N_5944,N_2946,N_1425);
or U5945 (N_5945,N_2819,N_1836);
nand U5946 (N_5946,N_239,N_440);
or U5947 (N_5947,N_1673,N_1095);
and U5948 (N_5948,N_25,N_3036);
nand U5949 (N_5949,N_126,N_1731);
and U5950 (N_5950,N_2902,N_1343);
nor U5951 (N_5951,N_1038,N_131);
and U5952 (N_5952,N_306,N_503);
nor U5953 (N_5953,N_761,N_313);
and U5954 (N_5954,N_867,N_2373);
xor U5955 (N_5955,N_1875,N_2679);
nor U5956 (N_5956,N_862,N_454);
nor U5957 (N_5957,N_1136,N_782);
xor U5958 (N_5958,N_2566,N_27);
xor U5959 (N_5959,N_1508,N_2572);
and U5960 (N_5960,N_3113,N_2387);
nor U5961 (N_5961,N_1613,N_131);
nand U5962 (N_5962,N_306,N_495);
nor U5963 (N_5963,N_798,N_3087);
nand U5964 (N_5964,N_2513,N_1132);
and U5965 (N_5965,N_392,N_140);
xnor U5966 (N_5966,N_2525,N_210);
nand U5967 (N_5967,N_198,N_828);
and U5968 (N_5968,N_2897,N_55);
or U5969 (N_5969,N_1668,N_1993);
xnor U5970 (N_5970,N_3004,N_634);
xnor U5971 (N_5971,N_2079,N_406);
or U5972 (N_5972,N_2116,N_2597);
nand U5973 (N_5973,N_6,N_357);
xor U5974 (N_5974,N_169,N_440);
and U5975 (N_5975,N_1763,N_895);
or U5976 (N_5976,N_1006,N_1239);
or U5977 (N_5977,N_1116,N_2212);
nor U5978 (N_5978,N_460,N_1859);
nand U5979 (N_5979,N_2792,N_1283);
nand U5980 (N_5980,N_725,N_832);
xor U5981 (N_5981,N_1622,N_897);
xnor U5982 (N_5982,N_1887,N_1649);
xnor U5983 (N_5983,N_2028,N_827);
and U5984 (N_5984,N_2228,N_228);
and U5985 (N_5985,N_130,N_752);
or U5986 (N_5986,N_89,N_391);
and U5987 (N_5987,N_518,N_1084);
nand U5988 (N_5988,N_1253,N_871);
or U5989 (N_5989,N_2150,N_2072);
or U5990 (N_5990,N_927,N_1110);
xnor U5991 (N_5991,N_2071,N_1368);
or U5992 (N_5992,N_2373,N_886);
nor U5993 (N_5993,N_1883,N_1771);
xor U5994 (N_5994,N_3114,N_1764);
nand U5995 (N_5995,N_1875,N_1054);
or U5996 (N_5996,N_2280,N_1511);
nand U5997 (N_5997,N_2237,N_2011);
and U5998 (N_5998,N_2353,N_1597);
or U5999 (N_5999,N_1216,N_1552);
and U6000 (N_6000,N_1745,N_2500);
and U6001 (N_6001,N_1894,N_355);
or U6002 (N_6002,N_2226,N_3088);
and U6003 (N_6003,N_1997,N_1413);
nor U6004 (N_6004,N_1990,N_406);
and U6005 (N_6005,N_2105,N_1719);
nor U6006 (N_6006,N_1590,N_831);
xor U6007 (N_6007,N_2171,N_2804);
nor U6008 (N_6008,N_94,N_965);
or U6009 (N_6009,N_1281,N_111);
or U6010 (N_6010,N_1517,N_820);
and U6011 (N_6011,N_1802,N_6);
and U6012 (N_6012,N_1531,N_62);
xor U6013 (N_6013,N_1537,N_1260);
xnor U6014 (N_6014,N_1387,N_746);
or U6015 (N_6015,N_1551,N_1966);
and U6016 (N_6016,N_2667,N_2429);
nor U6017 (N_6017,N_1006,N_2373);
nand U6018 (N_6018,N_2828,N_2086);
nand U6019 (N_6019,N_16,N_2438);
xnor U6020 (N_6020,N_1077,N_352);
xnor U6021 (N_6021,N_2122,N_2571);
and U6022 (N_6022,N_3026,N_2518);
or U6023 (N_6023,N_880,N_1156);
and U6024 (N_6024,N_2633,N_1040);
or U6025 (N_6025,N_2546,N_916);
xnor U6026 (N_6026,N_1716,N_1535);
and U6027 (N_6027,N_910,N_1435);
xor U6028 (N_6028,N_1897,N_1551);
or U6029 (N_6029,N_2155,N_3078);
and U6030 (N_6030,N_250,N_2466);
and U6031 (N_6031,N_1650,N_51);
or U6032 (N_6032,N_1255,N_1285);
and U6033 (N_6033,N_1073,N_674);
or U6034 (N_6034,N_1122,N_2426);
nor U6035 (N_6035,N_2022,N_1993);
and U6036 (N_6036,N_1859,N_3093);
nand U6037 (N_6037,N_1386,N_1858);
and U6038 (N_6038,N_2283,N_2701);
xnor U6039 (N_6039,N_1919,N_377);
and U6040 (N_6040,N_2737,N_2370);
or U6041 (N_6041,N_1176,N_2410);
or U6042 (N_6042,N_400,N_2996);
xnor U6043 (N_6043,N_430,N_390);
and U6044 (N_6044,N_1540,N_84);
and U6045 (N_6045,N_1013,N_1597);
xor U6046 (N_6046,N_2174,N_830);
or U6047 (N_6047,N_99,N_350);
and U6048 (N_6048,N_3066,N_212);
xnor U6049 (N_6049,N_1086,N_773);
and U6050 (N_6050,N_702,N_1879);
or U6051 (N_6051,N_1543,N_3119);
or U6052 (N_6052,N_3119,N_39);
or U6053 (N_6053,N_1923,N_2128);
xor U6054 (N_6054,N_2071,N_1381);
or U6055 (N_6055,N_2033,N_176);
nor U6056 (N_6056,N_2725,N_863);
xnor U6057 (N_6057,N_267,N_1533);
nand U6058 (N_6058,N_1595,N_1074);
nor U6059 (N_6059,N_1488,N_924);
nand U6060 (N_6060,N_94,N_205);
xnor U6061 (N_6061,N_1021,N_1076);
xor U6062 (N_6062,N_2667,N_2421);
nor U6063 (N_6063,N_3100,N_2200);
and U6064 (N_6064,N_283,N_1797);
nor U6065 (N_6065,N_83,N_2870);
nor U6066 (N_6066,N_507,N_2244);
nor U6067 (N_6067,N_2943,N_1643);
nor U6068 (N_6068,N_2220,N_3083);
xor U6069 (N_6069,N_2959,N_316);
xnor U6070 (N_6070,N_528,N_1586);
xor U6071 (N_6071,N_1001,N_1506);
nor U6072 (N_6072,N_2393,N_963);
and U6073 (N_6073,N_1333,N_1983);
nor U6074 (N_6074,N_222,N_2922);
xnor U6075 (N_6075,N_470,N_3079);
xnor U6076 (N_6076,N_2459,N_1942);
and U6077 (N_6077,N_2813,N_2979);
nand U6078 (N_6078,N_1535,N_2938);
xor U6079 (N_6079,N_65,N_188);
nor U6080 (N_6080,N_1339,N_2611);
nand U6081 (N_6081,N_2278,N_273);
nor U6082 (N_6082,N_2196,N_262);
nand U6083 (N_6083,N_1012,N_546);
or U6084 (N_6084,N_2907,N_1621);
nor U6085 (N_6085,N_1307,N_849);
nand U6086 (N_6086,N_2302,N_1050);
xnor U6087 (N_6087,N_977,N_1558);
xnor U6088 (N_6088,N_2640,N_843);
nor U6089 (N_6089,N_352,N_1401);
xnor U6090 (N_6090,N_2050,N_783);
or U6091 (N_6091,N_946,N_1661);
xor U6092 (N_6092,N_1091,N_2637);
nor U6093 (N_6093,N_2277,N_1235);
nand U6094 (N_6094,N_1929,N_2822);
nor U6095 (N_6095,N_2779,N_776);
or U6096 (N_6096,N_1344,N_383);
or U6097 (N_6097,N_3054,N_2030);
and U6098 (N_6098,N_889,N_651);
nand U6099 (N_6099,N_333,N_2805);
xnor U6100 (N_6100,N_1885,N_2198);
or U6101 (N_6101,N_1051,N_2082);
and U6102 (N_6102,N_2864,N_1029);
xor U6103 (N_6103,N_2386,N_311);
xnor U6104 (N_6104,N_1015,N_418);
and U6105 (N_6105,N_425,N_1510);
nor U6106 (N_6106,N_2443,N_1395);
xor U6107 (N_6107,N_2539,N_1281);
nand U6108 (N_6108,N_2596,N_2775);
xnor U6109 (N_6109,N_2912,N_2046);
or U6110 (N_6110,N_2876,N_2042);
nor U6111 (N_6111,N_1503,N_440);
xnor U6112 (N_6112,N_312,N_2760);
and U6113 (N_6113,N_162,N_26);
or U6114 (N_6114,N_1117,N_1321);
or U6115 (N_6115,N_669,N_2245);
nor U6116 (N_6116,N_2049,N_1716);
or U6117 (N_6117,N_2981,N_2607);
nor U6118 (N_6118,N_269,N_94);
and U6119 (N_6119,N_2291,N_1714);
nor U6120 (N_6120,N_3043,N_2948);
or U6121 (N_6121,N_1806,N_850);
and U6122 (N_6122,N_1660,N_248);
nand U6123 (N_6123,N_2846,N_1162);
xnor U6124 (N_6124,N_2096,N_2889);
nand U6125 (N_6125,N_2489,N_1402);
nor U6126 (N_6126,N_939,N_528);
and U6127 (N_6127,N_2652,N_1530);
nand U6128 (N_6128,N_2299,N_1186);
and U6129 (N_6129,N_2348,N_21);
nand U6130 (N_6130,N_2814,N_3099);
xor U6131 (N_6131,N_92,N_1985);
and U6132 (N_6132,N_1002,N_1051);
xnor U6133 (N_6133,N_1056,N_2671);
and U6134 (N_6134,N_3122,N_2766);
nor U6135 (N_6135,N_549,N_627);
and U6136 (N_6136,N_441,N_2549);
nand U6137 (N_6137,N_2491,N_2202);
and U6138 (N_6138,N_1059,N_1991);
nand U6139 (N_6139,N_2148,N_1163);
nand U6140 (N_6140,N_823,N_1270);
nor U6141 (N_6141,N_2242,N_1383);
and U6142 (N_6142,N_2243,N_1848);
nor U6143 (N_6143,N_38,N_511);
and U6144 (N_6144,N_1208,N_1536);
or U6145 (N_6145,N_43,N_2289);
and U6146 (N_6146,N_1487,N_1506);
and U6147 (N_6147,N_2466,N_1677);
xor U6148 (N_6148,N_1251,N_667);
and U6149 (N_6149,N_2169,N_695);
nand U6150 (N_6150,N_1699,N_261);
xor U6151 (N_6151,N_515,N_2828);
or U6152 (N_6152,N_1468,N_161);
nand U6153 (N_6153,N_2506,N_274);
or U6154 (N_6154,N_67,N_1306);
nand U6155 (N_6155,N_2937,N_2888);
or U6156 (N_6156,N_2313,N_1667);
or U6157 (N_6157,N_1709,N_1974);
xor U6158 (N_6158,N_1752,N_2992);
nor U6159 (N_6159,N_2617,N_2864);
nand U6160 (N_6160,N_2337,N_961);
and U6161 (N_6161,N_2740,N_2874);
nand U6162 (N_6162,N_783,N_2843);
or U6163 (N_6163,N_3049,N_1906);
and U6164 (N_6164,N_2516,N_2090);
or U6165 (N_6165,N_1505,N_2338);
and U6166 (N_6166,N_498,N_3097);
nor U6167 (N_6167,N_2685,N_2017);
or U6168 (N_6168,N_2261,N_2819);
nand U6169 (N_6169,N_2588,N_2129);
xor U6170 (N_6170,N_1331,N_703);
and U6171 (N_6171,N_1051,N_1940);
nor U6172 (N_6172,N_1315,N_942);
or U6173 (N_6173,N_2497,N_459);
nand U6174 (N_6174,N_5,N_587);
xor U6175 (N_6175,N_372,N_2890);
nand U6176 (N_6176,N_3116,N_871);
xor U6177 (N_6177,N_514,N_2552);
or U6178 (N_6178,N_2787,N_2648);
xnor U6179 (N_6179,N_2869,N_1434);
and U6180 (N_6180,N_827,N_1486);
xnor U6181 (N_6181,N_2663,N_2707);
or U6182 (N_6182,N_1811,N_830);
and U6183 (N_6183,N_352,N_1785);
xnor U6184 (N_6184,N_944,N_1647);
nor U6185 (N_6185,N_2026,N_1128);
nor U6186 (N_6186,N_644,N_943);
or U6187 (N_6187,N_131,N_120);
xor U6188 (N_6188,N_34,N_1144);
nor U6189 (N_6189,N_3099,N_148);
or U6190 (N_6190,N_2464,N_140);
nor U6191 (N_6191,N_1401,N_2954);
or U6192 (N_6192,N_921,N_2903);
or U6193 (N_6193,N_283,N_2867);
xor U6194 (N_6194,N_2533,N_3040);
and U6195 (N_6195,N_237,N_1099);
nor U6196 (N_6196,N_1336,N_2762);
or U6197 (N_6197,N_808,N_1188);
xor U6198 (N_6198,N_2222,N_471);
xor U6199 (N_6199,N_1077,N_2846);
nand U6200 (N_6200,N_2161,N_44);
nor U6201 (N_6201,N_2297,N_2139);
nand U6202 (N_6202,N_390,N_1601);
or U6203 (N_6203,N_656,N_2398);
nand U6204 (N_6204,N_1426,N_2327);
xor U6205 (N_6205,N_1270,N_657);
or U6206 (N_6206,N_671,N_1669);
and U6207 (N_6207,N_1673,N_454);
nor U6208 (N_6208,N_929,N_1125);
xor U6209 (N_6209,N_48,N_605);
or U6210 (N_6210,N_1191,N_460);
or U6211 (N_6211,N_2170,N_106);
xor U6212 (N_6212,N_1453,N_63);
nor U6213 (N_6213,N_2394,N_753);
nand U6214 (N_6214,N_3036,N_2507);
xnor U6215 (N_6215,N_1625,N_2373);
and U6216 (N_6216,N_2566,N_2104);
and U6217 (N_6217,N_2181,N_1431);
and U6218 (N_6218,N_2313,N_1600);
nor U6219 (N_6219,N_2719,N_2179);
and U6220 (N_6220,N_2142,N_1992);
xor U6221 (N_6221,N_526,N_1366);
nor U6222 (N_6222,N_1977,N_2687);
xnor U6223 (N_6223,N_2389,N_2345);
nand U6224 (N_6224,N_2259,N_2392);
and U6225 (N_6225,N_1859,N_1048);
nand U6226 (N_6226,N_1376,N_1360);
nor U6227 (N_6227,N_2869,N_999);
and U6228 (N_6228,N_2353,N_1529);
nand U6229 (N_6229,N_1468,N_2092);
and U6230 (N_6230,N_138,N_1481);
or U6231 (N_6231,N_197,N_76);
or U6232 (N_6232,N_1473,N_2966);
nand U6233 (N_6233,N_1647,N_293);
or U6234 (N_6234,N_542,N_258);
and U6235 (N_6235,N_1908,N_412);
and U6236 (N_6236,N_1533,N_1948);
xnor U6237 (N_6237,N_590,N_2886);
nand U6238 (N_6238,N_2718,N_1125);
and U6239 (N_6239,N_1278,N_2447);
nand U6240 (N_6240,N_1510,N_2365);
xnor U6241 (N_6241,N_2455,N_1334);
nor U6242 (N_6242,N_1578,N_2992);
and U6243 (N_6243,N_2913,N_1659);
or U6244 (N_6244,N_2499,N_953);
nand U6245 (N_6245,N_646,N_1206);
xor U6246 (N_6246,N_657,N_1157);
nor U6247 (N_6247,N_2499,N_1606);
and U6248 (N_6248,N_1753,N_2276);
nand U6249 (N_6249,N_1624,N_50);
xnor U6250 (N_6250,N_4167,N_3684);
nor U6251 (N_6251,N_3213,N_4541);
or U6252 (N_6252,N_5816,N_3214);
or U6253 (N_6253,N_5393,N_4945);
and U6254 (N_6254,N_3426,N_4833);
and U6255 (N_6255,N_3181,N_5860);
and U6256 (N_6256,N_4043,N_3869);
and U6257 (N_6257,N_5508,N_3242);
nor U6258 (N_6258,N_5991,N_5850);
xor U6259 (N_6259,N_3589,N_4728);
xor U6260 (N_6260,N_3389,N_4768);
nand U6261 (N_6261,N_4125,N_4271);
and U6262 (N_6262,N_3615,N_5800);
nand U6263 (N_6263,N_3929,N_4890);
nand U6264 (N_6264,N_3835,N_6232);
nor U6265 (N_6265,N_4574,N_3630);
xnor U6266 (N_6266,N_3241,N_4579);
xnor U6267 (N_6267,N_3330,N_5601);
nor U6268 (N_6268,N_6065,N_5896);
xor U6269 (N_6269,N_3159,N_5018);
and U6270 (N_6270,N_4030,N_4608);
or U6271 (N_6271,N_4094,N_5207);
nand U6272 (N_6272,N_5837,N_5329);
xnor U6273 (N_6273,N_6104,N_5332);
nor U6274 (N_6274,N_6137,N_6105);
nand U6275 (N_6275,N_3744,N_5311);
and U6276 (N_6276,N_4718,N_5528);
xor U6277 (N_6277,N_6006,N_4929);
nand U6278 (N_6278,N_3131,N_3656);
or U6279 (N_6279,N_4683,N_5874);
or U6280 (N_6280,N_3187,N_5989);
or U6281 (N_6281,N_3900,N_3909);
or U6282 (N_6282,N_5590,N_5302);
nand U6283 (N_6283,N_3863,N_4639);
nor U6284 (N_6284,N_4707,N_5554);
nor U6285 (N_6285,N_3260,N_5513);
or U6286 (N_6286,N_5063,N_4709);
xor U6287 (N_6287,N_5712,N_3613);
or U6288 (N_6288,N_4386,N_5765);
nand U6289 (N_6289,N_4753,N_4518);
nor U6290 (N_6290,N_3896,N_3884);
nor U6291 (N_6291,N_5367,N_4478);
xnor U6292 (N_6292,N_4018,N_5039);
or U6293 (N_6293,N_4651,N_5950);
or U6294 (N_6294,N_6239,N_3631);
xor U6295 (N_6295,N_4417,N_4534);
nor U6296 (N_6296,N_5038,N_5639);
nand U6297 (N_6297,N_5081,N_3182);
and U6298 (N_6298,N_6003,N_4046);
or U6299 (N_6299,N_5594,N_4476);
and U6300 (N_6300,N_6033,N_5410);
nand U6301 (N_6301,N_3259,N_5169);
nor U6302 (N_6302,N_3164,N_5321);
nand U6303 (N_6303,N_6139,N_4699);
nor U6304 (N_6304,N_5007,N_6014);
nor U6305 (N_6305,N_3162,N_5117);
nor U6306 (N_6306,N_6055,N_3377);
xor U6307 (N_6307,N_5012,N_4429);
xnor U6308 (N_6308,N_4860,N_3715);
xnor U6309 (N_6309,N_4242,N_4121);
nand U6310 (N_6310,N_3905,N_3697);
nor U6311 (N_6311,N_4636,N_5944);
nor U6312 (N_6312,N_3728,N_4104);
nand U6313 (N_6313,N_3165,N_5705);
and U6314 (N_6314,N_5632,N_5153);
nand U6315 (N_6315,N_5793,N_4703);
or U6316 (N_6316,N_3721,N_6138);
and U6317 (N_6317,N_4622,N_4186);
and U6318 (N_6318,N_5782,N_3899);
or U6319 (N_6319,N_4103,N_4973);
nor U6320 (N_6320,N_3366,N_3140);
or U6321 (N_6321,N_4588,N_3987);
nand U6322 (N_6322,N_5058,N_4794);
or U6323 (N_6323,N_4820,N_4040);
nor U6324 (N_6324,N_5203,N_4130);
or U6325 (N_6325,N_3901,N_4469);
or U6326 (N_6326,N_3846,N_5280);
and U6327 (N_6327,N_3271,N_3560);
nand U6328 (N_6328,N_4115,N_5602);
nor U6329 (N_6329,N_4907,N_4056);
and U6330 (N_6330,N_5664,N_5579);
xnor U6331 (N_6331,N_6000,N_3203);
and U6332 (N_6332,N_3446,N_6103);
and U6333 (N_6333,N_5562,N_4257);
and U6334 (N_6334,N_5480,N_3340);
nand U6335 (N_6335,N_4329,N_5985);
nor U6336 (N_6336,N_4602,N_4682);
nor U6337 (N_6337,N_6122,N_4733);
xnor U6338 (N_6338,N_4298,N_4615);
or U6339 (N_6339,N_4319,N_3280);
or U6340 (N_6340,N_4970,N_4077);
or U6341 (N_6341,N_5734,N_6085);
xnor U6342 (N_6342,N_4076,N_4179);
xor U6343 (N_6343,N_5478,N_4745);
nand U6344 (N_6344,N_4914,N_4238);
nor U6345 (N_6345,N_4091,N_5748);
or U6346 (N_6346,N_4049,N_3506);
and U6347 (N_6347,N_4169,N_5125);
or U6348 (N_6348,N_4510,N_5383);
xor U6349 (N_6349,N_5013,N_4882);
xnor U6350 (N_6350,N_3885,N_3368);
xnor U6351 (N_6351,N_3717,N_3765);
and U6352 (N_6352,N_5880,N_5017);
or U6353 (N_6353,N_5231,N_3387);
or U6354 (N_6354,N_3470,N_4932);
and U6355 (N_6355,N_3539,N_6154);
nor U6356 (N_6356,N_6168,N_3535);
nand U6357 (N_6357,N_5766,N_3853);
nand U6358 (N_6358,N_3382,N_5097);
nor U6359 (N_6359,N_4161,N_4010);
nand U6360 (N_6360,N_5312,N_3595);
xor U6361 (N_6361,N_5297,N_6184);
nor U6362 (N_6362,N_5413,N_3735);
xor U6363 (N_6363,N_6145,N_5261);
and U6364 (N_6364,N_3568,N_5703);
or U6365 (N_6365,N_4526,N_3665);
nand U6366 (N_6366,N_3352,N_5958);
or U6367 (N_6367,N_5627,N_3410);
nor U6368 (N_6368,N_5863,N_5300);
xor U6369 (N_6369,N_5648,N_5565);
and U6370 (N_6370,N_4689,N_4159);
nor U6371 (N_6371,N_5838,N_4552);
nand U6372 (N_6372,N_4585,N_6058);
xnor U6373 (N_6373,N_3991,N_4466);
or U6374 (N_6374,N_5202,N_3954);
and U6375 (N_6375,N_4968,N_3245);
xnor U6376 (N_6376,N_4688,N_5303);
nand U6377 (N_6377,N_4528,N_5374);
and U6378 (N_6378,N_5142,N_3264);
nand U6379 (N_6379,N_5946,N_3309);
xor U6380 (N_6380,N_3859,N_3473);
nand U6381 (N_6381,N_4821,N_5290);
nor U6382 (N_6382,N_4206,N_3325);
nor U6383 (N_6383,N_3793,N_5143);
or U6384 (N_6384,N_6019,N_5439);
xnor U6385 (N_6385,N_5737,N_5121);
or U6386 (N_6386,N_4744,N_3762);
and U6387 (N_6387,N_6045,N_3883);
nor U6388 (N_6388,N_4473,N_4392);
or U6389 (N_6389,N_3915,N_5453);
and U6390 (N_6390,N_6075,N_5882);
and U6391 (N_6391,N_6197,N_4813);
or U6392 (N_6392,N_4533,N_3633);
xor U6393 (N_6393,N_5209,N_4715);
or U6394 (N_6394,N_4201,N_3703);
and U6395 (N_6395,N_6140,N_3926);
nand U6396 (N_6396,N_3212,N_3277);
and U6397 (N_6397,N_4343,N_3167);
or U6398 (N_6398,N_6181,N_5885);
and U6399 (N_6399,N_5201,N_3946);
or U6400 (N_6400,N_5234,N_6161);
and U6401 (N_6401,N_5692,N_3985);
or U6402 (N_6402,N_4369,N_4668);
and U6403 (N_6403,N_3882,N_3658);
or U6404 (N_6404,N_5279,N_4407);
nor U6405 (N_6405,N_3579,N_5983);
and U6406 (N_6406,N_4942,N_3147);
nor U6407 (N_6407,N_4029,N_6147);
and U6408 (N_6408,N_3235,N_5357);
and U6409 (N_6409,N_5219,N_4572);
nand U6410 (N_6410,N_3827,N_5520);
nor U6411 (N_6411,N_3291,N_3622);
or U6412 (N_6412,N_4985,N_4455);
and U6413 (N_6413,N_3857,N_3937);
and U6414 (N_6414,N_4918,N_4053);
xnor U6415 (N_6415,N_4920,N_3191);
xor U6416 (N_6416,N_4583,N_4137);
nand U6417 (N_6417,N_5984,N_3781);
nor U6418 (N_6418,N_5824,N_3154);
xnor U6419 (N_6419,N_3716,N_5402);
xor U6420 (N_6420,N_3468,N_5593);
xnor U6421 (N_6421,N_3940,N_4756);
xnor U6422 (N_6422,N_6048,N_5877);
xnor U6423 (N_6423,N_4754,N_3730);
or U6424 (N_6424,N_3912,N_4354);
nand U6425 (N_6425,N_3374,N_3265);
nand U6426 (N_6426,N_5470,N_4724);
nand U6427 (N_6427,N_3526,N_3584);
xor U6428 (N_6428,N_3455,N_3585);
and U6429 (N_6429,N_3324,N_5049);
nand U6430 (N_6430,N_4274,N_5225);
xnor U6431 (N_6431,N_4562,N_5004);
or U6432 (N_6432,N_4925,N_3651);
nand U6433 (N_6433,N_3156,N_5700);
and U6434 (N_6434,N_4891,N_4923);
nor U6435 (N_6435,N_3625,N_5093);
or U6436 (N_6436,N_5629,N_6171);
or U6437 (N_6437,N_5922,N_4829);
nor U6438 (N_6438,N_3286,N_4031);
xnor U6439 (N_6439,N_5101,N_3930);
xnor U6440 (N_6440,N_6218,N_3945);
or U6441 (N_6441,N_4347,N_5879);
nand U6442 (N_6442,N_5335,N_6082);
xnor U6443 (N_6443,N_4113,N_4654);
or U6444 (N_6444,N_4864,N_3471);
and U6445 (N_6445,N_5675,N_3189);
and U6446 (N_6446,N_3327,N_4171);
nand U6447 (N_6447,N_3252,N_3565);
or U6448 (N_6448,N_4416,N_4627);
xnor U6449 (N_6449,N_5932,N_4032);
and U6450 (N_6450,N_4450,N_3641);
or U6451 (N_6451,N_3349,N_3314);
nor U6452 (N_6452,N_4126,N_4601);
and U6453 (N_6453,N_6206,N_3254);
or U6454 (N_6454,N_3461,N_4996);
xnor U6455 (N_6455,N_3807,N_4554);
or U6456 (N_6456,N_3590,N_4507);
or U6457 (N_6457,N_4906,N_5248);
or U6458 (N_6458,N_6176,N_4359);
and U6459 (N_6459,N_5835,N_3571);
and U6460 (N_6460,N_4935,N_4874);
nand U6461 (N_6461,N_3546,N_6109);
and U6462 (N_6462,N_4263,N_5843);
and U6463 (N_6463,N_5372,N_4646);
nor U6464 (N_6464,N_4247,N_4629);
nand U6465 (N_6465,N_4760,N_4513);
nand U6466 (N_6466,N_5241,N_5168);
xor U6467 (N_6467,N_4827,N_4068);
nor U6468 (N_6468,N_4940,N_4567);
nand U6469 (N_6469,N_6136,N_3424);
xor U6470 (N_6470,N_4441,N_5959);
nand U6471 (N_6471,N_4142,N_3887);
xnor U6472 (N_6472,N_3184,N_5062);
or U6473 (N_6473,N_6129,N_5795);
nor U6474 (N_6474,N_3257,N_3197);
or U6475 (N_6475,N_5543,N_4800);
nand U6476 (N_6476,N_3274,N_4494);
nand U6477 (N_6477,N_4661,N_5725);
or U6478 (N_6478,N_3823,N_6040);
xor U6479 (N_6479,N_4278,N_3889);
nand U6480 (N_6480,N_5979,N_5936);
xnor U6481 (N_6481,N_4057,N_6015);
and U6482 (N_6482,N_3984,N_5905);
nand U6483 (N_6483,N_5497,N_4938);
xor U6484 (N_6484,N_5037,N_4806);
or U6485 (N_6485,N_5555,N_4440);
or U6486 (N_6486,N_4729,N_4339);
and U6487 (N_6487,N_5130,N_4258);
or U6488 (N_6488,N_5612,N_3475);
nand U6489 (N_6489,N_4372,N_3217);
nor U6490 (N_6490,N_5432,N_3149);
xnor U6491 (N_6491,N_5380,N_4059);
and U6492 (N_6492,N_4272,N_3223);
xor U6493 (N_6493,N_3150,N_6204);
nand U6494 (N_6494,N_3190,N_5218);
and U6495 (N_6495,N_5006,N_5053);
xor U6496 (N_6496,N_3452,N_3606);
xnor U6497 (N_6497,N_5987,N_3466);
nor U6498 (N_6498,N_4796,N_5252);
nand U6499 (N_6499,N_3944,N_3799);
xnor U6500 (N_6500,N_4136,N_5047);
xnor U6501 (N_6501,N_4202,N_3752);
or U6502 (N_6502,N_3607,N_5412);
nand U6503 (N_6503,N_3636,N_5689);
and U6504 (N_6504,N_4908,N_4309);
nor U6505 (N_6505,N_5966,N_3617);
and U6506 (N_6506,N_3304,N_3856);
nor U6507 (N_6507,N_3440,N_6088);
or U6508 (N_6508,N_3422,N_5536);
nor U6509 (N_6509,N_5566,N_3688);
nor U6510 (N_6510,N_3512,N_3517);
or U6511 (N_6511,N_5861,N_5244);
nand U6512 (N_6512,N_4375,N_3811);
nand U6513 (N_6513,N_5735,N_5764);
xor U6514 (N_6514,N_5974,N_3768);
xor U6515 (N_6515,N_3971,N_3791);
and U6516 (N_6516,N_5479,N_4173);
nand U6517 (N_6517,N_4111,N_4722);
nor U6518 (N_6518,N_5730,N_5077);
or U6519 (N_6519,N_5324,N_3519);
and U6520 (N_6520,N_4519,N_5190);
and U6521 (N_6521,N_4315,N_4183);
nor U6522 (N_6522,N_3642,N_4857);
or U6523 (N_6523,N_5476,N_3146);
xor U6524 (N_6524,N_3723,N_3923);
nor U6525 (N_6525,N_5314,N_3754);
or U6526 (N_6526,N_5301,N_4460);
nor U6527 (N_6527,N_3763,N_4107);
nand U6528 (N_6528,N_4189,N_5526);
or U6529 (N_6529,N_5621,N_3219);
or U6530 (N_6530,N_3875,N_4720);
nand U6531 (N_6531,N_3787,N_4471);
nor U6532 (N_6532,N_3592,N_5890);
nand U6533 (N_6533,N_4835,N_5021);
and U6534 (N_6534,N_3640,N_5553);
and U6535 (N_6535,N_4437,N_3660);
xor U6536 (N_6536,N_5132,N_4486);
and U6537 (N_6537,N_3239,N_5733);
and U6538 (N_6538,N_4184,N_5355);
and U6539 (N_6539,N_4087,N_3614);
and U6540 (N_6540,N_3130,N_3441);
nand U6541 (N_6541,N_4358,N_3843);
xor U6542 (N_6542,N_5655,N_3982);
nand U6543 (N_6543,N_5556,N_5447);
nand U6544 (N_6544,N_4038,N_4695);
xnor U6545 (N_6545,N_5841,N_5784);
xor U6546 (N_6546,N_3710,N_3662);
nand U6547 (N_6547,N_4089,N_5030);
xor U6548 (N_6548,N_6162,N_5687);
or U6549 (N_6549,N_4606,N_3674);
or U6550 (N_6550,N_3713,N_5904);
and U6551 (N_6551,N_3193,N_4865);
nand U6552 (N_6552,N_4374,N_3145);
or U6553 (N_6553,N_5679,N_3431);
xnor U6554 (N_6554,N_6080,N_4544);
nand U6555 (N_6555,N_5490,N_4306);
nor U6556 (N_6556,N_5195,N_5173);
and U6557 (N_6557,N_4180,N_5379);
nand U6558 (N_6558,N_6099,N_3230);
or U6559 (N_6559,N_4127,N_4344);
xor U6560 (N_6560,N_3996,N_5622);
and U6561 (N_6561,N_6001,N_4809);
xnor U6562 (N_6562,N_5617,N_4066);
nand U6563 (N_6563,N_3798,N_4328);
nand U6564 (N_6564,N_5318,N_4547);
xor U6565 (N_6565,N_3370,N_4880);
nand U6566 (N_6566,N_4951,N_4879);
nor U6567 (N_6567,N_6169,N_3504);
xor U6568 (N_6568,N_3616,N_3417);
nor U6569 (N_6569,N_3933,N_3871);
and U6570 (N_6570,N_5464,N_3647);
nand U6571 (N_6571,N_3737,N_5487);
xnor U6572 (N_6572,N_5992,N_4964);
nand U6573 (N_6573,N_4168,N_5980);
or U6574 (N_6574,N_3231,N_5268);
nand U6575 (N_6575,N_5903,N_5749);
and U6576 (N_6576,N_6028,N_3559);
nand U6577 (N_6577,N_5511,N_4219);
nand U6578 (N_6578,N_4600,N_3215);
nand U6579 (N_6579,N_5886,N_3281);
and U6580 (N_6580,N_6121,N_3129);
nand U6581 (N_6581,N_6244,N_4398);
and U6582 (N_6582,N_3523,N_3652);
nand U6583 (N_6583,N_5996,N_6067);
nor U6584 (N_6584,N_4388,N_5953);
nor U6585 (N_6585,N_3232,N_4839);
or U6586 (N_6586,N_6054,N_4673);
and U6587 (N_6587,N_5845,N_4427);
nor U6588 (N_6588,N_3740,N_5282);
nor U6589 (N_6589,N_3678,N_5723);
or U6590 (N_6590,N_5570,N_5894);
and U6591 (N_6591,N_5112,N_5564);
nand U6592 (N_6592,N_4578,N_6044);
xor U6593 (N_6593,N_3518,N_4536);
xor U6594 (N_6594,N_4589,N_4342);
and U6595 (N_6595,N_4054,N_3329);
xnor U6596 (N_6596,N_5684,N_4497);
and U6597 (N_6597,N_5204,N_5605);
xor U6598 (N_6598,N_4015,N_3817);
or U6599 (N_6599,N_3877,N_6135);
nor U6600 (N_6600,N_3572,N_3602);
xor U6601 (N_6601,N_5127,N_4442);
xnor U6602 (N_6602,N_5937,N_6241);
nor U6603 (N_6603,N_4811,N_3591);
or U6604 (N_6604,N_5193,N_4904);
or U6605 (N_6605,N_4324,N_5086);
nand U6606 (N_6606,N_5309,N_3174);
xor U6607 (N_6607,N_4563,N_3675);
xor U6608 (N_6608,N_3436,N_4371);
nor U6609 (N_6609,N_5082,N_3700);
xnor U6610 (N_6610,N_4696,N_3527);
nand U6611 (N_6611,N_6102,N_3918);
and U6612 (N_6612,N_5275,N_3169);
xor U6613 (N_6613,N_3654,N_6226);
xor U6614 (N_6614,N_3224,N_5829);
nor U6615 (N_6615,N_5183,N_3433);
xnor U6616 (N_6616,N_5654,N_4525);
or U6617 (N_6617,N_5643,N_4250);
and U6618 (N_6618,N_4738,N_6125);
nor U6619 (N_6619,N_4605,N_4726);
xnor U6620 (N_6620,N_4674,N_5573);
nor U6621 (N_6621,N_5693,N_5855);
and U6622 (N_6622,N_5707,N_5444);
nand U6623 (N_6623,N_5574,N_5477);
nand U6624 (N_6624,N_5686,N_4607);
xnor U6625 (N_6625,N_3664,N_5468);
and U6626 (N_6626,N_4147,N_4260);
nor U6627 (N_6627,N_4200,N_3861);
nor U6628 (N_6628,N_5299,N_6091);
xnor U6629 (N_6629,N_5157,N_3483);
and U6630 (N_6630,N_5750,N_5229);
xnor U6631 (N_6631,N_5642,N_5438);
and U6632 (N_6632,N_5186,N_4074);
xor U6633 (N_6633,N_5095,N_5353);
nand U6634 (N_6634,N_3757,N_5771);
and U6635 (N_6635,N_4892,N_4402);
or U6636 (N_6636,N_3677,N_4373);
nand U6637 (N_6637,N_4824,N_3570);
nand U6638 (N_6638,N_4725,N_3619);
xnor U6639 (N_6639,N_3498,N_5341);
nor U6640 (N_6640,N_4414,N_3803);
or U6641 (N_6641,N_3359,N_6069);
and U6642 (N_6642,N_5074,N_3460);
and U6643 (N_6643,N_4364,N_4109);
nor U6644 (N_6644,N_5775,N_6153);
nand U6645 (N_6645,N_4766,N_4784);
nor U6646 (N_6646,N_4083,N_5015);
xnor U6647 (N_6647,N_3586,N_5338);
xor U6648 (N_6648,N_6183,N_3965);
nand U6649 (N_6649,N_5461,N_4872);
and U6650 (N_6650,N_4732,N_4296);
or U6651 (N_6651,N_4262,N_5398);
and U6652 (N_6652,N_3759,N_5113);
and U6653 (N_6653,N_5571,N_4899);
or U6654 (N_6654,N_4859,N_4735);
nor U6655 (N_6655,N_3554,N_4337);
xnor U6656 (N_6656,N_4998,N_4119);
or U6657 (N_6657,N_4524,N_4305);
nand U6658 (N_6658,N_6203,N_5939);
or U6659 (N_6659,N_6056,N_3139);
or U6660 (N_6660,N_4084,N_5714);
or U6661 (N_6661,N_4956,N_3198);
xor U6662 (N_6662,N_5681,N_3216);
or U6663 (N_6663,N_4251,N_5967);
nor U6664 (N_6664,N_4625,N_4195);
or U6665 (N_6665,N_5454,N_5706);
nand U6666 (N_6666,N_4667,N_3296);
nand U6667 (N_6667,N_3205,N_5298);
nand U6668 (N_6668,N_4152,N_4690);
or U6669 (N_6669,N_5313,N_4470);
nand U6670 (N_6670,N_5760,N_5948);
or U6671 (N_6671,N_4156,N_5931);
and U6672 (N_6672,N_4292,N_5741);
and U6673 (N_6673,N_4922,N_6178);
and U6674 (N_6674,N_5657,N_6220);
xor U6675 (N_6675,N_4840,N_4236);
nand U6676 (N_6676,N_5396,N_5893);
and U6677 (N_6677,N_3786,N_6020);
xor U6678 (N_6678,N_6225,N_4332);
and U6679 (N_6679,N_5485,N_4431);
and U6680 (N_6680,N_5080,N_3567);
and U6681 (N_6681,N_6196,N_5395);
xnor U6682 (N_6682,N_3258,N_5177);
or U6683 (N_6683,N_5167,N_5952);
nand U6684 (N_6684,N_3474,N_4546);
and U6685 (N_6685,N_3671,N_5865);
nand U6686 (N_6686,N_5065,N_5381);
nand U6687 (N_6687,N_5481,N_4816);
or U6688 (N_6688,N_3454,N_5519);
xnor U6689 (N_6689,N_4999,N_6134);
xor U6690 (N_6690,N_3620,N_3425);
nor U6691 (N_6691,N_6143,N_4436);
and U6692 (N_6692,N_4229,N_6238);
or U6693 (N_6693,N_5745,N_5133);
and U6694 (N_6694,N_5522,N_3204);
xnor U6695 (N_6695,N_5452,N_3300);
nor U6696 (N_6696,N_4118,N_3751);
xor U6697 (N_6697,N_3702,N_3893);
nor U6698 (N_6698,N_5525,N_3921);
nor U6699 (N_6699,N_3415,N_5977);
nand U6700 (N_6700,N_3880,N_3326);
xor U6701 (N_6701,N_3549,N_5633);
nor U6702 (N_6702,N_5319,N_3979);
nand U6703 (N_6703,N_3821,N_5994);
nand U6704 (N_6704,N_4868,N_3496);
nand U6705 (N_6705,N_5718,N_3743);
and U6706 (N_6706,N_5866,N_4924);
or U6707 (N_6707,N_4385,N_5405);
xnor U6708 (N_6708,N_4836,N_4791);
xnor U6709 (N_6709,N_4154,N_3952);
xnor U6710 (N_6710,N_3538,N_4687);
xnor U6711 (N_6711,N_4153,N_5220);
or U6712 (N_6712,N_3604,N_4506);
and U6713 (N_6713,N_6011,N_4336);
nand U6714 (N_6714,N_4997,N_6043);
nand U6715 (N_6715,N_3412,N_5092);
nor U6716 (N_6716,N_4477,N_5933);
or U6717 (N_6717,N_3545,N_5751);
nand U6718 (N_6718,N_5255,N_5366);
and U6719 (N_6719,N_4088,N_3298);
nor U6720 (N_6720,N_3550,N_5999);
and U6721 (N_6721,N_4082,N_4050);
xnor U6722 (N_6722,N_3188,N_5224);
or U6723 (N_6723,N_3500,N_6243);
nor U6724 (N_6724,N_3973,N_4493);
and U6725 (N_6725,N_4325,N_3854);
nand U6726 (N_6726,N_3959,N_5029);
xnor U6727 (N_6727,N_5899,N_4580);
or U6728 (N_6728,N_4656,N_5443);
xnor U6729 (N_6729,N_5502,N_3739);
and U6730 (N_6730,N_5671,N_4335);
xnor U6731 (N_6731,N_5813,N_4406);
and U6732 (N_6732,N_4955,N_6008);
nor U6733 (N_6733,N_5295,N_3769);
nor U6734 (N_6734,N_5869,N_5048);
or U6735 (N_6735,N_5662,N_3342);
or U6736 (N_6736,N_4832,N_6007);
or U6737 (N_6737,N_3967,N_3936);
or U6738 (N_6738,N_4164,N_5702);
xnor U6739 (N_6739,N_3222,N_5064);
or U6740 (N_6740,N_4789,N_3977);
nor U6741 (N_6741,N_3719,N_4395);
xnor U6742 (N_6742,N_5323,N_6199);
nor U6743 (N_6743,N_6108,N_3497);
nand U6744 (N_6744,N_6095,N_3405);
nor U6745 (N_6745,N_5728,N_5346);
or U6746 (N_6746,N_3638,N_5363);
and U6747 (N_6747,N_5673,N_3379);
and U6748 (N_6748,N_3364,N_5762);
nand U6749 (N_6749,N_5289,N_4447);
or U6750 (N_6750,N_5834,N_4543);
and U6751 (N_6751,N_3598,N_5360);
nand U6752 (N_6752,N_3593,N_3581);
nand U6753 (N_6753,N_4765,N_4190);
xor U6754 (N_6754,N_4419,N_4096);
and U6755 (N_6755,N_5499,N_5975);
or U6756 (N_6756,N_5551,N_3886);
nor U6757 (N_6757,N_3323,N_3234);
or U6758 (N_6758,N_5767,N_5292);
xor U6759 (N_6759,N_3450,N_5469);
nand U6760 (N_6760,N_3777,N_5139);
and U6761 (N_6761,N_3401,N_5839);
nand U6762 (N_6762,N_3284,N_5942);
or U6763 (N_6763,N_3731,N_3447);
xor U6764 (N_6764,N_4933,N_4931);
or U6765 (N_6765,N_3983,N_5377);
and U6766 (N_6766,N_3404,N_3419);
nand U6767 (N_6767,N_3736,N_4512);
and U6768 (N_6768,N_4937,N_5722);
nor U6769 (N_6769,N_4582,N_5900);
or U6770 (N_6770,N_5875,N_5242);
nor U6771 (N_6771,N_3238,N_5217);
nor U6772 (N_6772,N_4529,N_4098);
or U6773 (N_6773,N_4387,N_4095);
xnor U6774 (N_6774,N_6030,N_5951);
and U6775 (N_6775,N_3294,N_5666);
or U6776 (N_6776,N_3462,N_5524);
and U6777 (N_6777,N_3732,N_4828);
or U6778 (N_6778,N_5431,N_3569);
or U6779 (N_6779,N_3293,N_5009);
nor U6780 (N_6780,N_4894,N_4815);
nand U6781 (N_6781,N_4255,N_5165);
nand U6782 (N_6782,N_4128,N_4462);
or U6783 (N_6783,N_4149,N_3653);
or U6784 (N_6784,N_4830,N_3919);
nand U6785 (N_6785,N_5779,N_3542);
nor U6786 (N_6786,N_3201,N_3499);
nand U6787 (N_6787,N_5409,N_3143);
nor U6788 (N_6788,N_5315,N_4527);
and U6789 (N_6789,N_3151,N_5531);
and U6790 (N_6790,N_4716,N_5344);
or U6791 (N_6791,N_4241,N_6062);
and U6792 (N_6792,N_5802,N_5325);
or U6793 (N_6793,N_5070,N_5527);
or U6794 (N_6794,N_5175,N_6059);
xor U6795 (N_6795,N_5336,N_5756);
and U6796 (N_6796,N_3704,N_3166);
or U6797 (N_6797,N_4209,N_4261);
nor U6798 (N_6798,N_4803,N_4612);
nand U6799 (N_6799,N_4027,N_4853);
nor U6800 (N_6800,N_4210,N_3177);
nand U6801 (N_6801,N_4657,N_5720);
xnor U6802 (N_6802,N_3634,N_4215);
or U6803 (N_6803,N_3698,N_3975);
or U6804 (N_6804,N_4747,N_3482);
and U6805 (N_6805,N_3599,N_4075);
xnor U6806 (N_6806,N_6191,N_5156);
nor U6807 (N_6807,N_5957,N_5505);
xnor U6808 (N_6808,N_3211,N_5930);
nor U6809 (N_6809,N_4949,N_3333);
and U6810 (N_6810,N_3318,N_3556);
xnor U6811 (N_6811,N_3328,N_5540);
xnor U6812 (N_6812,N_5233,N_4966);
nor U6813 (N_6813,N_3953,N_5831);
xor U6814 (N_6814,N_3522,N_6240);
and U6815 (N_6815,N_3808,N_4393);
nand U6816 (N_6816,N_6126,N_4340);
xnor U6817 (N_6817,N_4649,N_5907);
and U6818 (N_6818,N_4623,N_3623);
or U6819 (N_6819,N_4897,N_3695);
xnor U6820 (N_6820,N_5397,N_4781);
xor U6821 (N_6821,N_6227,N_5079);
and U6822 (N_6822,N_5791,N_4499);
nor U6823 (N_6823,N_4067,N_3434);
nor U6824 (N_6824,N_4539,N_5184);
or U6825 (N_6825,N_3845,N_5888);
xnor U6826 (N_6826,N_3344,N_5256);
or U6827 (N_6827,N_5825,N_4143);
nor U6828 (N_6828,N_6194,N_4560);
nor U6829 (N_6829,N_5504,N_4706);
xor U6830 (N_6830,N_5103,N_5386);
xnor U6831 (N_6831,N_4614,N_3136);
or U6832 (N_6832,N_3648,N_6151);
nand U6833 (N_6833,N_3943,N_3531);
nor U6834 (N_6834,N_5471,N_4983);
or U6835 (N_6835,N_5000,N_4211);
nand U6836 (N_6836,N_5812,N_4675);
xor U6837 (N_6837,N_4736,N_4122);
or U6838 (N_6838,N_3372,N_5521);
nand U6839 (N_6839,N_5102,N_4590);
or U6840 (N_6840,N_4883,N_4301);
nor U6841 (N_6841,N_3746,N_6061);
xor U6842 (N_6842,N_5917,N_3141);
nand U6843 (N_6843,N_4762,N_5625);
nor U6844 (N_6844,N_4786,N_3770);
xnor U6845 (N_6845,N_5337,N_5213);
nor U6846 (N_6846,N_6128,N_5534);
and U6847 (N_6847,N_6046,N_3673);
or U6848 (N_6848,N_5178,N_3487);
nand U6849 (N_6849,N_3942,N_4637);
nand U6850 (N_6850,N_3494,N_3828);
nand U6851 (N_6851,N_4487,N_4222);
nor U6852 (N_6852,N_4797,N_3694);
nand U6853 (N_6853,N_4755,N_4199);
or U6854 (N_6854,N_5910,N_4253);
or U6855 (N_6855,N_6222,N_3179);
or U6856 (N_6856,N_4187,N_4341);
xnor U6857 (N_6857,N_4587,N_5390);
nand U6858 (N_6858,N_5740,N_3335);
and U6859 (N_6859,N_6159,N_3445);
xnor U6860 (N_6860,N_4299,N_5032);
and U6861 (N_6861,N_5757,N_4818);
nor U6862 (N_6862,N_5873,N_5842);
nor U6863 (N_6863,N_4802,N_4491);
or U6864 (N_6864,N_4163,N_5238);
nand U6865 (N_6865,N_5585,N_6083);
or U6866 (N_6866,N_3826,N_5407);
nand U6867 (N_6867,N_4438,N_5704);
or U6868 (N_6868,N_3851,N_5266);
nor U6869 (N_6869,N_3133,N_4737);
nor U6870 (N_6870,N_5960,N_5041);
and U6871 (N_6871,N_5307,N_4535);
nor U6872 (N_6872,N_4285,N_4484);
xor U6873 (N_6873,N_6211,N_4678);
xnor U6874 (N_6874,N_3725,N_5055);
xor U6875 (N_6875,N_4205,N_3135);
nand U6876 (N_6876,N_4194,N_4348);
nor U6877 (N_6877,N_5916,N_4975);
nor U6878 (N_6878,N_4981,N_4467);
nor U6879 (N_6879,N_4284,N_4982);
nand U6880 (N_6880,N_3505,N_3629);
or U6881 (N_6881,N_5572,N_4302);
nand U6882 (N_6882,N_5050,N_5858);
xnor U6883 (N_6883,N_3916,N_4092);
nand U6884 (N_6884,N_4172,N_5235);
nand U6885 (N_6885,N_4379,N_5116);
or U6886 (N_6886,N_3183,N_4653);
or U6887 (N_6887,N_3830,N_4283);
nor U6888 (N_6888,N_5925,N_3680);
xor U6889 (N_6889,N_5826,N_5428);
and U6890 (N_6890,N_3148,N_3564);
or U6891 (N_6891,N_4457,N_5460);
xor U6892 (N_6892,N_4871,N_5068);
nor U6893 (N_6893,N_4898,N_6177);
nor U6894 (N_6894,N_4916,N_6247);
nor U6895 (N_6895,N_4846,N_3236);
nor U6896 (N_6896,N_5550,N_3292);
nand U6897 (N_6897,N_3451,N_6224);
or U6898 (N_6898,N_3659,N_5624);
nor U6899 (N_6899,N_4788,N_3373);
xnor U6900 (N_6900,N_5440,N_4515);
xnor U6901 (N_6901,N_5777,N_4994);
nor U6902 (N_6902,N_3488,N_4175);
or U6903 (N_6903,N_5317,N_5563);
nand U6904 (N_6904,N_4779,N_4714);
or U6905 (N_6905,N_5797,N_5658);
or U6906 (N_6906,N_3790,N_5938);
xnor U6907 (N_6907,N_4408,N_3225);
xnor U6908 (N_6908,N_3345,N_3914);
and U6909 (N_6909,N_4669,N_4817);
nand U6910 (N_6910,N_5920,N_5811);
and U6911 (N_6911,N_5887,N_4459);
nand U6912 (N_6912,N_3813,N_6188);
or U6913 (N_6913,N_5088,N_3375);
or U6914 (N_6914,N_4954,N_5924);
xor U6915 (N_6915,N_4464,N_3993);
and U6916 (N_6916,N_6223,N_5544);
and U6917 (N_6917,N_5847,N_5862);
nand U6918 (N_6918,N_6124,N_5151);
and U6919 (N_6919,N_3537,N_3268);
xnor U6920 (N_6920,N_6068,N_5598);
and U6921 (N_6921,N_4220,N_3693);
nor U6922 (N_6922,N_4785,N_3511);
and U6923 (N_6923,N_6149,N_5541);
nand U6924 (N_6924,N_3667,N_6180);
or U6925 (N_6925,N_4566,N_3192);
nand U6926 (N_6926,N_4986,N_3485);
and U6927 (N_6927,N_4680,N_3794);
and U6928 (N_6928,N_5072,N_5259);
and U6929 (N_6929,N_3547,N_3776);
xor U6930 (N_6930,N_3528,N_4134);
nand U6931 (N_6931,N_4862,N_3949);
xnor U6932 (N_6932,N_3261,N_3402);
nor U6933 (N_6933,N_5210,N_5054);
and U6934 (N_6934,N_3317,N_4230);
and U6935 (N_6935,N_3683,N_5604);
or U6936 (N_6936,N_5166,N_4885);
or U6937 (N_6937,N_4719,N_4058);
xor U6938 (N_6938,N_5514,N_5090);
nand U6939 (N_6939,N_4265,N_3134);
nand U6940 (N_6940,N_4702,N_5972);
nor U6941 (N_6941,N_4227,N_5434);
nor U6942 (N_6942,N_5940,N_4514);
xnor U6943 (N_6943,N_6221,N_4322);
or U6944 (N_6944,N_4902,N_5646);
xnor U6945 (N_6945,N_4390,N_4866);
nor U6946 (N_6946,N_5044,N_5581);
or U6947 (N_6947,N_5243,N_5978);
nor U6948 (N_6948,N_3142,N_5619);
nand U6949 (N_6949,N_5736,N_4888);
or U6950 (N_6950,N_4845,N_3153);
xor U6951 (N_6951,N_5316,N_4397);
or U6952 (N_6952,N_3720,N_5988);
nor U6953 (N_6953,N_4490,N_6248);
and U6954 (N_6954,N_4645,N_5495);
nand U6955 (N_6955,N_5964,N_3849);
nor U6956 (N_6956,N_3806,N_3348);
and U6957 (N_6957,N_3319,N_3578);
and U6958 (N_6958,N_5196,N_3409);
or U6959 (N_6959,N_5919,N_5459);
and U6960 (N_6960,N_6150,N_4266);
xnor U6961 (N_6961,N_4132,N_4838);
xor U6962 (N_6962,N_5465,N_5264);
nor U6963 (N_6963,N_5537,N_5260);
or U6964 (N_6964,N_4213,N_5898);
or U6965 (N_6965,N_4599,N_4798);
xor U6966 (N_6966,N_5124,N_5584);
or U6967 (N_6967,N_4952,N_4763);
and U6968 (N_6968,N_4223,N_6041);
xnor U6969 (N_6969,N_5688,N_5792);
or U6970 (N_6970,N_4676,N_5682);
nand U6971 (N_6971,N_5591,N_5456);
and U6972 (N_6972,N_3920,N_5091);
nand U6973 (N_6973,N_4987,N_3472);
or U6974 (N_6974,N_4767,N_3534);
nor U6975 (N_6975,N_3398,N_5387);
nand U6976 (N_6976,N_4382,N_3202);
xor U6977 (N_6977,N_4004,N_3321);
nand U6978 (N_6978,N_6163,N_3897);
and U6979 (N_6979,N_4980,N_5986);
and U6980 (N_6980,N_5027,N_5160);
nand U6981 (N_6981,N_5083,N_4093);
xnor U6982 (N_6982,N_6026,N_5685);
nand U6983 (N_6983,N_4465,N_5094);
nand U6984 (N_6984,N_3307,N_3628);
or U6985 (N_6985,N_6010,N_3955);
and U6986 (N_6986,N_4297,N_5868);
nor U6987 (N_6987,N_3432,N_4114);
or U6988 (N_6988,N_5200,N_6132);
or U6989 (N_6989,N_3386,N_3395);
xor U6990 (N_6990,N_5067,N_6057);
nand U6991 (N_6991,N_5895,N_5727);
nand U6992 (N_6992,N_4456,N_4140);
nor U6993 (N_6993,N_5785,N_6142);
xnor U6994 (N_6994,N_4957,N_6200);
and U6995 (N_6995,N_5651,N_3775);
xor U6996 (N_6996,N_4584,N_5668);
or U6997 (N_6997,N_4492,N_4734);
or U6998 (N_6998,N_5251,N_5005);
and U6999 (N_6999,N_5257,N_5138);
and U7000 (N_7000,N_5949,N_4609);
xnor U7001 (N_7001,N_5118,N_3376);
or U7002 (N_7002,N_3418,N_3390);
xnor U7003 (N_7003,N_3687,N_4807);
and U7004 (N_7004,N_3381,N_5997);
and U7005 (N_7005,N_5599,N_4943);
and U7006 (N_7006,N_5352,N_4138);
or U7007 (N_7007,N_6074,N_3573);
xor U7008 (N_7008,N_6086,N_3297);
and U7009 (N_7009,N_4941,N_3714);
or U7010 (N_7010,N_3964,N_4063);
nor U7011 (N_7011,N_5378,N_3272);
xnor U7012 (N_7012,N_5135,N_5848);
nor U7013 (N_7013,N_4910,N_3263);
nand U7014 (N_7014,N_3999,N_6157);
or U7015 (N_7015,N_5721,N_3927);
nor U7016 (N_7016,N_3553,N_5236);
nand U7017 (N_7017,N_5789,N_5155);
xor U7018 (N_7018,N_4776,N_4313);
or U7019 (N_7019,N_5111,N_5161);
xnor U7020 (N_7020,N_3276,N_5631);
or U7021 (N_7021,N_3789,N_3691);
and U7022 (N_7022,N_4042,N_5884);
xor U7023 (N_7023,N_4704,N_4670);
and U7024 (N_7024,N_5976,N_5031);
nand U7025 (N_7025,N_3320,N_6190);
nand U7026 (N_7026,N_3865,N_4333);
xor U7027 (N_7027,N_5045,N_5089);
nand U7028 (N_7028,N_5119,N_4212);
xnor U7029 (N_7029,N_6034,N_6193);
and U7030 (N_7030,N_6146,N_4252);
nor U7031 (N_7031,N_5758,N_3876);
nor U7032 (N_7032,N_5445,N_6093);
and U7033 (N_7033,N_5414,N_3661);
or U7034 (N_7034,N_4008,N_6119);
xor U7035 (N_7035,N_3476,N_5222);
nand U7036 (N_7036,N_5060,N_5610);
nor U7037 (N_7037,N_5819,N_3701);
and U7038 (N_7038,N_4648,N_6036);
nand U7039 (N_7039,N_5163,N_5724);
and U7040 (N_7040,N_4400,N_4834);
or U7041 (N_7041,N_6111,N_5212);
and U7042 (N_7042,N_5227,N_4501);
nand U7043 (N_7043,N_3430,N_5359);
xnor U7044 (N_7044,N_5342,N_4041);
nand U7045 (N_7045,N_5947,N_3733);
xor U7046 (N_7046,N_5990,N_3911);
xor U7047 (N_7047,N_4367,N_3495);
nand U7048 (N_7048,N_5641,N_5628);
xnor U7049 (N_7049,N_3127,N_3650);
and U7050 (N_7050,N_6076,N_5181);
and U7051 (N_7051,N_5066,N_6023);
and U7052 (N_7052,N_5814,N_3741);
nand U7053 (N_7053,N_4145,N_4881);
or U7054 (N_7054,N_4896,N_6246);
nand U7055 (N_7055,N_4376,N_4934);
or U7056 (N_7056,N_3563,N_3925);
or U7057 (N_7057,N_5246,N_4026);
xor U7058 (N_7058,N_3760,N_4550);
nand U7059 (N_7059,N_4988,N_5539);
and U7060 (N_7060,N_5339,N_3574);
or U7061 (N_7061,N_3413,N_4568);
nor U7062 (N_7062,N_4958,N_5473);
nor U7063 (N_7063,N_6202,N_5391);
nor U7064 (N_7064,N_4001,N_3540);
nand U7065 (N_7065,N_6114,N_3644);
xnor U7066 (N_7066,N_5969,N_3339);
nand U7067 (N_7067,N_4990,N_5458);
or U7068 (N_7068,N_5022,N_3510);
nand U7069 (N_7069,N_4362,N_4557);
nand U7070 (N_7070,N_3699,N_5489);
nor U7071 (N_7071,N_5817,N_3976);
or U7072 (N_7072,N_3966,N_5179);
nor U7073 (N_7073,N_5981,N_5608);
nand U7074 (N_7074,N_5331,N_3988);
and U7075 (N_7075,N_4391,N_5560);
xor U7076 (N_7076,N_3705,N_5286);
and U7077 (N_7077,N_5437,N_4764);
xnor U7078 (N_7078,N_3492,N_5968);
nor U7079 (N_7079,N_3750,N_5016);
xnor U7080 (N_7080,N_5057,N_4700);
and U7081 (N_7081,N_3618,N_4444);
xor U7082 (N_7082,N_3525,N_5929);
or U7083 (N_7083,N_3420,N_5450);
or U7084 (N_7084,N_6120,N_5278);
nand U7085 (N_7085,N_5530,N_3639);
nor U7086 (N_7086,N_6035,N_3478);
xnor U7087 (N_7087,N_6079,N_4647);
xnor U7088 (N_7088,N_5596,N_4224);
xnor U7089 (N_7089,N_5773,N_6029);
or U7090 (N_7090,N_5310,N_3453);
nand U7091 (N_7091,N_4672,N_4630);
nand U7092 (N_7092,N_4102,N_3895);
xor U7093 (N_7093,N_4962,N_5761);
and U7094 (N_7094,N_3906,N_3520);
nor U7095 (N_7095,N_5995,N_4185);
nor U7096 (N_7096,N_5107,N_4404);
xor U7097 (N_7097,N_5287,N_4064);
nand U7098 (N_7098,N_3902,N_3458);
nor U7099 (N_7099,N_5618,N_3247);
nor U7100 (N_7100,N_3463,N_3848);
or U7101 (N_7101,N_3128,N_3246);
and U7102 (N_7102,N_4995,N_5836);
xnor U7103 (N_7103,N_3180,N_5014);
nor U7104 (N_7104,N_4321,N_4445);
nor U7105 (N_7105,N_5955,N_3290);
nor U7106 (N_7106,N_4021,N_5973);
xor U7107 (N_7107,N_4327,N_4282);
nand U7108 (N_7108,N_4979,N_4842);
nand U7109 (N_7109,N_5901,N_5897);
or U7110 (N_7110,N_5215,N_3233);
nand U7111 (N_7111,N_4155,N_5913);
and U7112 (N_7112,N_4237,N_5475);
or U7113 (N_7113,N_5284,N_5798);
or U7114 (N_7114,N_4193,N_4556);
and U7115 (N_7115,N_4502,N_4759);
nor U7116 (N_7116,N_4498,N_5144);
or U7117 (N_7117,N_4823,N_4020);
or U7118 (N_7118,N_3501,N_4575);
nand U7119 (N_7119,N_5911,N_4418);
xor U7120 (N_7120,N_5794,N_5411);
and U7121 (N_7121,N_3437,N_4804);
nand U7122 (N_7122,N_5368,N_3243);
or U7123 (N_7123,N_3870,N_5533);
xor U7124 (N_7124,N_5109,N_3668);
or U7125 (N_7125,N_3753,N_4698);
and U7126 (N_7126,N_4435,N_6112);
nor U7127 (N_7127,N_5676,N_3521);
and U7128 (N_7128,N_5586,N_4577);
nor U7129 (N_7129,N_3583,N_3341);
or U7130 (N_7130,N_4946,N_5463);
nand U7131 (N_7131,N_5388,N_6155);
nand U7132 (N_7132,N_5518,N_4717);
and U7133 (N_7133,N_3747,N_3306);
or U7134 (N_7134,N_4628,N_3712);
xor U7135 (N_7135,N_5385,N_5320);
nor U7136 (N_7136,N_3439,N_6013);
or U7137 (N_7137,N_5114,N_3138);
or U7138 (N_7138,N_4967,N_3477);
nand U7139 (N_7139,N_3682,N_4071);
xnor U7140 (N_7140,N_5369,N_4875);
and U7141 (N_7141,N_4727,N_4901);
xor U7142 (N_7142,N_3577,N_5422);
xor U7143 (N_7143,N_6107,N_3594);
nor U7144 (N_7144,N_4948,N_6195);
nand U7145 (N_7145,N_5965,N_4245);
xor U7146 (N_7146,N_6096,N_5020);
and U7147 (N_7147,N_5576,N_5696);
and U7148 (N_7148,N_3814,N_4825);
xor U7149 (N_7149,N_5909,N_3480);
and U7150 (N_7150,N_5501,N_4080);
xnor U7151 (N_7151,N_6022,N_4331);
or U7152 (N_7152,N_4405,N_5011);
and U7153 (N_7153,N_4900,N_6100);
nor U7154 (N_7154,N_3267,N_3825);
or U7155 (N_7155,N_6094,N_3672);
xor U7156 (N_7156,N_5698,N_3562);
and U7157 (N_7157,N_3986,N_5844);
or U7158 (N_7158,N_3186,N_4863);
nand U7159 (N_7159,N_5123,N_6098);
or U7160 (N_7160,N_3742,N_3396);
or U7161 (N_7161,N_3820,N_3210);
nand U7162 (N_7162,N_3288,N_3403);
or U7163 (N_7163,N_3388,N_5406);
nand U7164 (N_7164,N_5263,N_4078);
xnor U7165 (N_7165,N_5636,N_3974);
nor U7166 (N_7166,N_5881,N_5427);
nand U7167 (N_7167,N_5649,N_4551);
or U7168 (N_7168,N_5592,N_5373);
and U7169 (N_7169,N_5683,N_5425);
nand U7170 (N_7170,N_4151,N_5849);
xor U7171 (N_7171,N_4780,N_3502);
and U7172 (N_7172,N_5665,N_5024);
or U7173 (N_7173,N_3544,N_5472);
nor U7174 (N_7174,N_5799,N_5915);
or U7175 (N_7175,N_3380,N_5827);
or U7176 (N_7176,N_6131,N_4304);
or U7177 (N_7177,N_5430,N_4971);
nor U7178 (N_7178,N_5857,N_4231);
or U7179 (N_7179,N_4072,N_4293);
or U7180 (N_7180,N_5731,N_5164);
nor U7181 (N_7181,N_6209,N_5085);
nand U7182 (N_7182,N_6063,N_4055);
nor U7183 (N_7183,N_3783,N_6186);
nand U7184 (N_7184,N_5420,N_6172);
and U7185 (N_7185,N_3552,N_4869);
xor U7186 (N_7186,N_3637,N_5253);
xor U7187 (N_7187,N_3416,N_5653);
xor U7188 (N_7188,N_5451,N_3655);
nand U7189 (N_7189,N_3160,N_4805);
xnor U7190 (N_7190,N_3874,N_4424);
nand U7191 (N_7191,N_4801,N_5375);
and U7192 (N_7192,N_4003,N_3408);
nand U7193 (N_7193,N_4310,N_4503);
or U7194 (N_7194,N_5129,N_4269);
xor U7195 (N_7195,N_6060,N_5600);
and U7196 (N_7196,N_5247,N_4665);
or U7197 (N_7197,N_4758,N_5498);
xnor U7198 (N_7198,N_4959,N_4479);
and U7199 (N_7199,N_5548,N_4819);
xor U7200 (N_7200,N_5971,N_5697);
xnor U7201 (N_7201,N_5954,N_4895);
xor U7202 (N_7202,N_3429,N_5558);
nor U7203 (N_7203,N_4787,N_5921);
nor U7204 (N_7204,N_5822,N_5906);
xnor U7205 (N_7205,N_3934,N_4259);
xor U7206 (N_7206,N_3315,N_3312);
or U7207 (N_7207,N_4691,N_5354);
or U7208 (N_7208,N_4522,N_6087);
and U7209 (N_7209,N_4065,N_3864);
xor U7210 (N_7210,N_4586,N_5856);
nand U7211 (N_7211,N_4160,N_4540);
xnor U7212 (N_7212,N_4928,N_3970);
xor U7213 (N_7213,N_3868,N_5871);
nor U7214 (N_7214,N_3600,N_5345);
nand U7215 (N_7215,N_3360,N_5361);
xnor U7216 (N_7216,N_4773,N_4116);
xor U7217 (N_7217,N_6049,N_5872);
xnor U7218 (N_7218,N_4294,N_6230);
and U7219 (N_7219,N_3253,N_3172);
nand U7220 (N_7220,N_3161,N_4774);
nand U7221 (N_7221,N_4176,N_5998);
nand U7222 (N_7222,N_6236,N_4432);
or U7223 (N_7223,N_3711,N_3513);
or U7224 (N_7224,N_4953,N_4679);
nor U7225 (N_7225,N_3666,N_4616);
and U7226 (N_7226,N_5429,N_4613);
xnor U7227 (N_7227,N_5126,N_3171);
nand U7228 (N_7228,N_5547,N_3270);
xnor U7229 (N_7229,N_3343,N_5365);
or U7230 (N_7230,N_6148,N_3218);
or U7231 (N_7231,N_5019,N_3797);
nor U7232 (N_7232,N_4463,N_5801);
nand U7233 (N_7233,N_5484,N_4847);
nor U7234 (N_7234,N_3881,N_5656);
and U7235 (N_7235,N_4972,N_5546);
and U7236 (N_7236,N_5327,N_4361);
and U7237 (N_7237,N_4511,N_3670);
and U7238 (N_7238,N_3273,N_5265);
nand U7239 (N_7239,N_5003,N_5630);
and U7240 (N_7240,N_4275,N_3459);
and U7241 (N_7241,N_4481,N_3939);
xor U7242 (N_7242,N_5529,N_3301);
or U7243 (N_7243,N_4531,N_5650);
xnor U7244 (N_7244,N_4141,N_4135);
nand U7245 (N_7245,N_4182,N_5442);
or U7246 (N_7246,N_4295,N_5823);
and U7247 (N_7247,N_6066,N_4218);
nand U7248 (N_7248,N_5349,N_3626);
and U7249 (N_7249,N_4267,N_6115);
and U7250 (N_7250,N_3960,N_4969);
or U7251 (N_7251,N_3557,N_5711);
nor U7252 (N_7252,N_3338,N_3961);
nor U7253 (N_7253,N_5878,N_3336);
nand U7254 (N_7254,N_3467,N_4217);
or U7255 (N_7255,N_4323,N_3206);
and U7256 (N_7256,N_4542,N_5637);
nor U7257 (N_7257,N_6144,N_5441);
or U7258 (N_7258,N_5457,N_3289);
nor U7259 (N_7259,N_4005,N_4855);
or U7260 (N_7260,N_5902,N_3310);
nor U7261 (N_7261,N_5815,N_3779);
nor U7262 (N_7262,N_3679,N_3981);
nor U7263 (N_7263,N_4356,N_3941);
xnor U7264 (N_7264,N_4286,N_4197);
nand U7265 (N_7265,N_5423,N_5889);
nor U7266 (N_7266,N_3411,N_4039);
or U7267 (N_7267,N_6092,N_3962);
xnor U7268 (N_7268,N_4468,N_4019);
xnor U7269 (N_7269,N_3514,N_3509);
xnor U7270 (N_7270,N_5392,N_4731);
xor U7271 (N_7271,N_4790,N_5403);
nor U7272 (N_7272,N_4203,N_5701);
nand U7273 (N_7273,N_5638,N_3469);
or U7274 (N_7274,N_3400,N_3561);
nor U7275 (N_7275,N_3196,N_6245);
and U7276 (N_7276,N_3892,N_3755);
or U7277 (N_7277,N_5214,N_5035);
or U7278 (N_7278,N_5744,N_3490);
and U7279 (N_7279,N_5076,N_4624);
nor U7280 (N_7280,N_4330,N_5305);
and U7281 (N_7281,N_4401,N_4684);
nor U7282 (N_7282,N_4693,N_4453);
nand U7283 (N_7283,N_5270,N_6210);
xnor U7284 (N_7284,N_6130,N_5503);
or U7285 (N_7285,N_4394,N_5726);
or U7286 (N_7286,N_5506,N_3530);
nor U7287 (N_7287,N_5538,N_4023);
and U7288 (N_7288,N_3663,N_4363);
nor U7289 (N_7289,N_4778,N_3758);
xnor U7290 (N_7290,N_4047,N_4538);
nor U7291 (N_7291,N_5294,N_6158);
and U7292 (N_7292,N_6052,N_6025);
xnor U7293 (N_7293,N_5854,N_5634);
and U7294 (N_7294,N_3515,N_3957);
nand U7295 (N_7295,N_6032,N_4281);
and U7296 (N_7296,N_5652,N_3443);
and U7297 (N_7297,N_5230,N_5710);
or U7298 (N_7298,N_6009,N_5061);
or U7299 (N_7299,N_3302,N_4079);
xor U7300 (N_7300,N_5708,N_3738);
or U7301 (N_7301,N_5262,N_3709);
nand U7302 (N_7302,N_5492,N_4635);
and U7303 (N_7303,N_6090,N_3862);
xor U7304 (N_7304,N_3457,N_3724);
and U7305 (N_7305,N_5768,N_6050);
nor U7306 (N_7306,N_3603,N_5542);
nor U7307 (N_7307,N_3240,N_4843);
and U7308 (N_7308,N_3785,N_4848);
nor U7309 (N_7309,N_3580,N_5840);
or U7310 (N_7310,N_4711,N_6207);
nand U7311 (N_7311,N_5535,N_4659);
nor U7312 (N_7312,N_5401,N_3423);
or U7313 (N_7313,N_3322,N_5182);
or U7314 (N_7314,N_4553,N_3866);
or U7315 (N_7315,N_4006,N_4100);
and U7316 (N_7316,N_4686,N_5069);
and U7317 (N_7317,N_3773,N_5400);
xor U7318 (N_7318,N_4034,N_5100);
nand U7319 (N_7319,N_3804,N_3624);
nand U7320 (N_7320,N_4208,N_5587);
and U7321 (N_7321,N_3543,N_3951);
or U7322 (N_7322,N_4549,N_5545);
nor U7323 (N_7323,N_4244,N_5356);
xnor U7324 (N_7324,N_5328,N_4712);
or U7325 (N_7325,N_5669,N_5281);
and U7326 (N_7326,N_5833,N_4604);
and U7327 (N_7327,N_3207,N_4597);
xor U7328 (N_7328,N_3575,N_4632);
xnor U7329 (N_7329,N_4769,N_6002);
xnor U7330 (N_7330,N_5732,N_5496);
nor U7331 (N_7331,N_3555,N_3209);
or U7332 (N_7332,N_5567,N_5435);
or U7333 (N_7333,N_4960,N_6016);
nand U7334 (N_7334,N_4870,N_6071);
nor U7335 (N_7335,N_5308,N_3995);
nand U7336 (N_7336,N_4909,N_3228);
xor U7337 (N_7337,N_4939,N_6216);
xnor U7338 (N_7338,N_4926,N_4318);
or U7339 (N_7339,N_4268,N_4509);
and U7340 (N_7340,N_5228,N_4831);
xnor U7341 (N_7341,N_3299,N_4350);
nor U7342 (N_7342,N_5051,N_5075);
xnor U7343 (N_7343,N_3722,N_5171);
and U7344 (N_7344,N_4642,N_4537);
nand U7345 (N_7345,N_4877,N_3649);
nand U7346 (N_7346,N_4887,N_5941);
nor U7347 (N_7347,N_5993,N_3852);
xor U7348 (N_7348,N_3227,N_3898);
xor U7349 (N_7349,N_4850,N_4051);
and U7350 (N_7350,N_5982,N_3928);
and U7351 (N_7351,N_5810,N_4984);
xor U7352 (N_7352,N_3152,N_4192);
or U7353 (N_7353,N_4452,N_3611);
nand U7354 (N_7354,N_4254,N_3176);
nor U7355 (N_7355,N_5269,N_6165);
xor U7356 (N_7356,N_4085,N_5188);
and U7357 (N_7357,N_3406,N_3596);
nand U7358 (N_7358,N_6208,N_4300);
nor U7359 (N_7359,N_5923,N_4380);
xor U7360 (N_7360,N_3158,N_5755);
or U7361 (N_7361,N_4012,N_4120);
or U7362 (N_7362,N_5943,N_4399);
xor U7363 (N_7363,N_3392,N_3894);
xnor U7364 (N_7364,N_5046,N_5786);
or U7365 (N_7365,N_3168,N_4413);
xor U7366 (N_7366,N_3812,N_5606);
nand U7367 (N_7367,N_4617,N_5738);
and U7368 (N_7368,N_5883,N_3938);
and U7369 (N_7369,N_3428,N_4730);
or U7370 (N_7370,N_5221,N_3194);
or U7371 (N_7371,N_6234,N_4521);
or U7372 (N_7372,N_5382,N_3486);
nor U7373 (N_7373,N_5348,N_4795);
and U7374 (N_7374,N_4415,N_4287);
nand U7375 (N_7375,N_3255,N_4852);
and U7376 (N_7376,N_5597,N_3351);
nor U7377 (N_7377,N_3249,N_4799);
or U7378 (N_7378,N_4009,N_4430);
nor U7379 (N_7379,N_3279,N_3609);
xnor U7380 (N_7380,N_5807,N_6038);
or U7381 (N_7381,N_4496,N_5276);
or U7382 (N_7382,N_6164,N_5582);
or U7383 (N_7383,N_4308,N_5717);
or U7384 (N_7384,N_5025,N_4421);
nor U7385 (N_7385,N_3311,N_3879);
nand U7386 (N_7386,N_4692,N_4017);
nor U7387 (N_7387,N_5002,N_4621);
nand U7388 (N_7388,N_3832,N_5211);
xnor U7389 (N_7389,N_3358,N_4610);
and U7390 (N_7390,N_5417,N_5918);
or U7391 (N_7391,N_5148,N_4403);
or U7392 (N_7392,N_3990,N_4591);
or U7393 (N_7393,N_5763,N_4370);
xnor U7394 (N_7394,N_4694,N_6189);
nand U7395 (N_7395,N_6031,N_5695);
or U7396 (N_7396,N_3878,N_3137);
or U7397 (N_7397,N_4317,N_4086);
or U7398 (N_7398,N_3287,N_4073);
xnor U7399 (N_7399,N_3838,N_3397);
or U7400 (N_7400,N_3749,N_5523);
and U7401 (N_7401,N_4069,N_5467);
and U7402 (N_7402,N_4234,N_5408);
or U7403 (N_7403,N_5963,N_4782);
or U7404 (N_7404,N_5096,N_4884);
nor U7405 (N_7405,N_5084,N_5892);
and U7406 (N_7406,N_5575,N_3815);
xor U7407 (N_7407,N_3834,N_4037);
xor U7408 (N_7408,N_4396,N_6018);
nor U7409 (N_7409,N_5626,N_3173);
nor U7410 (N_7410,N_4307,N_4517);
nor U7411 (N_7411,N_6005,N_3676);
nor U7412 (N_7412,N_5110,N_4264);
nand U7413 (N_7413,N_4652,N_3994);
xnor U7414 (N_7414,N_5589,N_4007);
xnor U7415 (N_7415,N_5659,N_3810);
xnor U7416 (N_7416,N_4061,N_6047);
or U7417 (N_7417,N_3357,N_5772);
or U7418 (N_7418,N_5809,N_3407);
xnor U7419 (N_7419,N_5851,N_5743);
or U7420 (N_7420,N_5120,N_3689);
nand U7421 (N_7421,N_6179,N_5023);
or U7422 (N_7422,N_6152,N_4276);
xnor U7423 (N_7423,N_5042,N_5418);
or U7424 (N_7424,N_6116,N_4867);
xnor U7425 (N_7425,N_5672,N_3438);
or U7426 (N_7426,N_6039,N_4148);
nor U7427 (N_7427,N_4508,N_6051);
nand U7428 (N_7428,N_4290,N_4545);
xor U7429 (N_7429,N_5272,N_6173);
or U7430 (N_7430,N_4743,N_4638);
nor U7431 (N_7431,N_4188,N_4139);
and U7432 (N_7432,N_3587,N_6118);
nor U7433 (N_7433,N_4124,N_6214);
xnor U7434 (N_7434,N_5620,N_5208);
nor U7435 (N_7435,N_5787,N_5569);
or U7436 (N_7436,N_5970,N_5140);
and U7437 (N_7437,N_4256,N_5945);
and U7438 (N_7438,N_3481,N_3774);
nand U7439 (N_7439,N_4489,N_6175);
nor U7440 (N_7440,N_5040,N_5716);
nor U7441 (N_7441,N_3508,N_4381);
nor U7442 (N_7442,N_3978,N_5515);
nor U7443 (N_7443,N_3313,N_3935);
and U7444 (N_7444,N_4603,N_3772);
and U7445 (N_7445,N_4002,N_4748);
or U7446 (N_7446,N_3831,N_4761);
and U7447 (N_7447,N_4420,N_4425);
nand U7448 (N_7448,N_4548,N_5351);
nor U7449 (N_7449,N_3332,N_6229);
nand U7450 (N_7450,N_3605,N_4280);
or U7451 (N_7451,N_5071,N_3316);
or U7452 (N_7452,N_4793,N_3727);
and U7453 (N_7453,N_5623,N_6170);
or U7454 (N_7454,N_4446,N_4157);
nor U7455 (N_7455,N_5491,N_5449);
nand U7456 (N_7456,N_5609,N_4663);
nand U7457 (N_7457,N_4316,N_5416);
xor U7458 (N_7458,N_4214,N_5509);
nor U7459 (N_7459,N_3394,N_5507);
or U7460 (N_7460,N_6242,N_5131);
and U7461 (N_7461,N_5059,N_4170);
xor U7462 (N_7462,N_4228,N_5364);
and U7463 (N_7463,N_5056,N_5493);
nand U7464 (N_7464,N_4814,N_3484);
nand U7465 (N_7465,N_5580,N_5258);
and U7466 (N_7466,N_5249,N_3858);
nand U7467 (N_7467,N_5934,N_3414);
nand U7468 (N_7468,N_6141,N_4144);
or U7469 (N_7469,N_5180,N_4174);
or U7470 (N_7470,N_5134,N_5296);
nand U7471 (N_7471,N_6106,N_4277);
xnor U7472 (N_7472,N_4752,N_6228);
xnor U7473 (N_7473,N_3516,N_3924);
nand U7474 (N_7474,N_5852,N_4620);
or U7475 (N_7475,N_4105,N_5271);
xnor U7476 (N_7476,N_4346,N_4961);
or U7477 (N_7477,N_4658,N_5715);
nand U7478 (N_7478,N_3908,N_5162);
xnor U7479 (N_7479,N_6064,N_5828);
nor U7480 (N_7480,N_5436,N_5419);
xor U7481 (N_7481,N_3354,N_3275);
nor U7482 (N_7482,N_5486,N_5394);
or U7483 (N_7483,N_3795,N_5306);
or U7484 (N_7484,N_4461,N_5776);
nor U7485 (N_7485,N_3383,N_3597);
nand U7486 (N_7486,N_6133,N_4483);
or U7487 (N_7487,N_3867,N_5729);
or U7488 (N_7488,N_4048,N_3841);
nand U7489 (N_7489,N_3904,N_4619);
xnor U7490 (N_7490,N_5304,N_5908);
nor U7491 (N_7491,N_3847,N_5660);
xnor U7492 (N_7492,N_6123,N_4808);
nand U7493 (N_7493,N_4225,N_5223);
xor U7494 (N_7494,N_4576,N_5559);
xor U7495 (N_7495,N_4944,N_4474);
and U7496 (N_7496,N_5846,N_4936);
nor U7497 (N_7497,N_4685,N_4989);
nor U7498 (N_7498,N_3256,N_3244);
xor U7499 (N_7499,N_5197,N_4123);
or U7500 (N_7500,N_4721,N_3690);
xnor U7501 (N_7501,N_5752,N_3669);
nand U7502 (N_7502,N_5891,N_3778);
xnor U7503 (N_7503,N_3685,N_4915);
nor U7504 (N_7504,N_3465,N_4666);
or U7505 (N_7505,N_5176,N_4482);
xnor U7506 (N_7506,N_3819,N_5674);
xor U7507 (N_7507,N_3989,N_4810);
and U7508 (N_7508,N_3829,N_6117);
xnor U7509 (N_7509,N_5577,N_4011);
xor U7510 (N_7510,N_4443,N_4841);
xor U7511 (N_7511,N_5780,N_5028);
nor U7512 (N_7512,N_4565,N_5187);
or U7513 (N_7513,N_4025,N_4488);
xor U7514 (N_7514,N_5274,N_5739);
and U7515 (N_7515,N_3997,N_3331);
or U7516 (N_7516,N_5237,N_3479);
and U7517 (N_7517,N_4963,N_4516);
xor U7518 (N_7518,N_3696,N_5232);
or U7519 (N_7519,N_4303,N_3367);
and U7520 (N_7520,N_3493,N_6182);
nor U7521 (N_7521,N_3353,N_5036);
nand U7522 (N_7522,N_3221,N_5146);
and U7523 (N_7523,N_4423,N_5746);
nor U7524 (N_7524,N_3144,N_3491);
nand U7525 (N_7525,N_4233,N_4378);
nand U7526 (N_7526,N_5226,N_6037);
xor U7527 (N_7527,N_5853,N_4475);
nor U7528 (N_7528,N_3229,N_5347);
xnor U7529 (N_7529,N_3612,N_3163);
or U7530 (N_7530,N_5189,N_3175);
or U7531 (N_7531,N_3448,N_4108);
xor U7532 (N_7532,N_6215,N_4014);
nand U7533 (N_7533,N_4740,N_4351);
and U7534 (N_7534,N_4334,N_4555);
or U7535 (N_7535,N_3816,N_4530);
or U7536 (N_7536,N_3860,N_3601);
nor U7537 (N_7537,N_4207,N_5549);
xor U7538 (N_7538,N_6167,N_4365);
or U7539 (N_7539,N_3842,N_4792);
nor U7540 (N_7540,N_5152,N_4592);
nor U7541 (N_7541,N_4650,N_4226);
or U7542 (N_7542,N_3947,N_4861);
xor U7543 (N_7543,N_4713,N_4112);
nand U7544 (N_7544,N_5448,N_4741);
and U7545 (N_7545,N_5699,N_4439);
nor U7546 (N_7546,N_6070,N_3170);
and U7547 (N_7547,N_5483,N_4974);
or U7548 (N_7548,N_5927,N_4595);
and U7549 (N_7549,N_4573,N_5333);
or U7550 (N_7550,N_4196,N_3305);
nor U7551 (N_7551,N_5326,N_3844);
nor U7552 (N_7552,N_4751,N_6110);
and U7553 (N_7553,N_3980,N_3551);
or U7554 (N_7554,N_6205,N_5137);
or U7555 (N_7555,N_4593,N_6101);
xor U7556 (N_7556,N_5870,N_4349);
or U7557 (N_7557,N_5283,N_4771);
or U7558 (N_7558,N_3645,N_3399);
or U7559 (N_7559,N_3524,N_3507);
and U7560 (N_7560,N_3185,N_3761);
nor U7561 (N_7561,N_3707,N_5008);
nand U7562 (N_7562,N_3248,N_5645);
or U7563 (N_7563,N_5742,N_3771);
nor U7564 (N_7564,N_4433,N_4978);
and U7565 (N_7565,N_3378,N_3621);
nor U7566 (N_7566,N_6217,N_4249);
or U7567 (N_7567,N_4288,N_4384);
nor U7568 (N_7568,N_6017,N_4366);
xor U7569 (N_7569,N_5415,N_3766);
nand U7570 (N_7570,N_3873,N_5774);
nor U7571 (N_7571,N_4927,N_5001);
or U7572 (N_7572,N_4641,N_6113);
nor U7573 (N_7573,N_4532,N_3903);
and U7574 (N_7574,N_4893,N_4618);
and U7575 (N_7575,N_3393,N_3421);
or U7576 (N_7576,N_3442,N_5170);
nor U7577 (N_7577,N_5043,N_6156);
nand U7578 (N_7578,N_4204,N_4166);
xnor U7579 (N_7579,N_3576,N_3251);
or U7580 (N_7580,N_4177,N_5482);
xnor U7581 (N_7581,N_5615,N_3627);
nand U7582 (N_7582,N_6235,N_4314);
or U7583 (N_7583,N_3734,N_5370);
or U7584 (N_7584,N_4451,N_5611);
nand U7585 (N_7585,N_3237,N_5462);
nand U7586 (N_7586,N_5557,N_5912);
xnor U7587 (N_7587,N_3756,N_4913);
or U7588 (N_7588,N_5713,N_5115);
and U7589 (N_7589,N_6042,N_5474);
and U7590 (N_7590,N_5517,N_3308);
xnor U7591 (N_7591,N_5322,N_4570);
xnor U7592 (N_7592,N_4449,N_4681);
or U7593 (N_7593,N_4854,N_4504);
and U7594 (N_7594,N_5267,N_5803);
and U7595 (N_7595,N_4723,N_5783);
or U7596 (N_7596,N_3269,N_4036);
xor U7597 (N_7597,N_5108,N_4664);
xnor U7598 (N_7598,N_4523,N_4273);
or U7599 (N_7599,N_4770,N_5778);
xnor U7600 (N_7600,N_3283,N_6024);
nor U7601 (N_7601,N_4631,N_3334);
or U7602 (N_7602,N_5240,N_4311);
or U7603 (N_7603,N_4912,N_5245);
or U7604 (N_7604,N_4458,N_3922);
and U7605 (N_7605,N_4750,N_3632);
or U7606 (N_7606,N_3347,N_4558);
xnor U7607 (N_7607,N_4279,N_3800);
or U7608 (N_7608,N_6012,N_4248);
nor U7609 (N_7609,N_4097,N_5532);
xnor U7610 (N_7610,N_4368,N_6185);
and U7611 (N_7611,N_5709,N_4919);
xor U7612 (N_7612,N_5098,N_4045);
nand U7613 (N_7613,N_4775,N_3262);
nor U7614 (N_7614,N_6127,N_4070);
nor U7615 (N_7615,N_4596,N_5607);
nand U7616 (N_7616,N_4992,N_4357);
xnor U7617 (N_7617,N_4905,N_4106);
and U7618 (N_7618,N_5330,N_4013);
and U7619 (N_7619,N_4131,N_4917);
nand U7620 (N_7620,N_3686,N_3764);
nand U7621 (N_7621,N_4165,N_3788);
nand U7622 (N_7622,N_4520,N_5034);
nand U7623 (N_7623,N_5747,N_3363);
and U7624 (N_7624,N_5185,N_3608);
or U7625 (N_7625,N_3362,N_3355);
nand U7626 (N_7626,N_5343,N_5433);
nand U7627 (N_7627,N_4611,N_5678);
xnor U7628 (N_7628,N_5864,N_3285);
or U7629 (N_7629,N_3824,N_4886);
and U7630 (N_7630,N_3836,N_4858);
nand U7631 (N_7631,N_3266,N_4389);
xnor U7632 (N_7632,N_5677,N_5759);
nand U7633 (N_7633,N_3818,N_5149);
and U7634 (N_7634,N_4598,N_4561);
or U7635 (N_7635,N_5288,N_3391);
or U7636 (N_7636,N_3784,N_5205);
xor U7637 (N_7637,N_3805,N_3346);
and U7638 (N_7638,N_5147,N_3969);
nand U7639 (N_7639,N_3226,N_4662);
and U7640 (N_7640,N_3888,N_5832);
xor U7641 (N_7641,N_3456,N_4783);
or U7642 (N_7642,N_3533,N_3155);
nand U7643 (N_7643,N_5588,N_3958);
xnor U7644 (N_7644,N_4360,N_5719);
nor U7645 (N_7645,N_4062,N_5616);
xnor U7646 (N_7646,N_5154,N_3792);
and U7647 (N_7647,N_3385,N_6089);
nand U7648 (N_7648,N_5122,N_4640);
or U7649 (N_7649,N_5362,N_5404);
and U7650 (N_7650,N_5680,N_5277);
nand U7651 (N_7651,N_3278,N_4090);
nor U7652 (N_7652,N_5033,N_6213);
nor U7653 (N_7653,N_5568,N_4705);
nor U7654 (N_7654,N_5962,N_4500);
nand U7655 (N_7655,N_4876,N_3890);
xor U7656 (N_7656,N_4660,N_6004);
xor U7657 (N_7657,N_5466,N_4239);
or U7658 (N_7658,N_4338,N_5808);
or U7659 (N_7659,N_4052,N_5141);
nor U7660 (N_7660,N_5206,N_5928);
nor U7661 (N_7661,N_3199,N_5104);
nand U7662 (N_7662,N_5334,N_4950);
and U7663 (N_7663,N_5216,N_3801);
nor U7664 (N_7664,N_5561,N_5796);
nand U7665 (N_7665,N_4873,N_4044);
nand U7666 (N_7666,N_3200,N_4033);
and U7667 (N_7667,N_4634,N_5194);
and U7668 (N_7668,N_4976,N_4434);
nor U7669 (N_7669,N_3282,N_4448);
or U7670 (N_7670,N_4677,N_4822);
xor U7671 (N_7671,N_6160,N_5192);
nand U7672 (N_7672,N_4411,N_5661);
and U7673 (N_7673,N_4594,N_4345);
or U7674 (N_7674,N_3337,N_5239);
and U7675 (N_7675,N_5867,N_5426);
nor U7676 (N_7676,N_3371,N_6072);
nand U7677 (N_7677,N_3208,N_5198);
xnor U7678 (N_7678,N_4426,N_4826);
xnor U7679 (N_7679,N_4235,N_3582);
xnor U7680 (N_7680,N_4749,N_3384);
or U7681 (N_7681,N_4150,N_4633);
or U7682 (N_7682,N_3365,N_3796);
nor U7683 (N_7683,N_4409,N_3998);
and U7684 (N_7684,N_3427,N_4701);
xnor U7685 (N_7685,N_3726,N_5788);
and U7686 (N_7686,N_4270,N_3295);
nor U7687 (N_7687,N_5818,N_6231);
nor U7688 (N_7688,N_6027,N_3369);
xnor U7689 (N_7689,N_4480,N_3435);
and U7690 (N_7690,N_3972,N_3850);
and U7691 (N_7691,N_4947,N_5595);
and U7692 (N_7692,N_5128,N_3566);
xor U7693 (N_7693,N_4991,N_3992);
xnor U7694 (N_7694,N_5552,N_3449);
xnor U7695 (N_7695,N_3489,N_4022);
nand U7696 (N_7696,N_4129,N_4320);
nor U7697 (N_7697,N_5935,N_3361);
nand U7698 (N_7698,N_5424,N_3558);
nand U7699 (N_7699,N_4352,N_3220);
nand U7700 (N_7700,N_3718,N_3541);
nand U7701 (N_7701,N_4246,N_3635);
and U7702 (N_7702,N_4878,N_3729);
xor U7703 (N_7703,N_5500,N_6192);
and U7704 (N_7704,N_4746,N_5578);
or U7705 (N_7705,N_4739,N_5250);
xor U7706 (N_7706,N_4559,N_4993);
or U7707 (N_7707,N_5052,N_6073);
xor U7708 (N_7708,N_4016,N_3782);
nand U7709 (N_7709,N_5583,N_3536);
nand U7710 (N_7710,N_5455,N_3963);
and U7711 (N_7711,N_5754,N_4889);
xnor U7712 (N_7712,N_4289,N_6174);
and U7713 (N_7713,N_4505,N_3907);
xor U7714 (N_7714,N_5647,N_5603);
and U7715 (N_7715,N_3822,N_3250);
xor U7716 (N_7716,N_4472,N_5914);
and U7717 (N_7717,N_4412,N_4240);
nand U7718 (N_7718,N_5753,N_4428);
nand U7719 (N_7719,N_5644,N_4110);
nor U7720 (N_7720,N_4564,N_4710);
nor U7721 (N_7721,N_3917,N_5926);
or U7722 (N_7722,N_4178,N_5670);
or U7723 (N_7723,N_4000,N_5770);
xnor U7724 (N_7724,N_3840,N_4243);
xor U7725 (N_7725,N_5663,N_5159);
nand U7726 (N_7726,N_5010,N_4930);
and U7727 (N_7727,N_6233,N_4221);
nor U7728 (N_7728,N_6249,N_4643);
nand U7729 (N_7729,N_3126,N_5150);
xor U7730 (N_7730,N_4812,N_4060);
and U7731 (N_7731,N_5172,N_4158);
and U7732 (N_7732,N_3809,N_5806);
nand U7733 (N_7733,N_5421,N_5804);
xnor U7734 (N_7734,N_5512,N_6201);
xnor U7735 (N_7735,N_4485,N_6053);
and U7736 (N_7736,N_3646,N_6187);
nor U7737 (N_7737,N_4837,N_3913);
xnor U7738 (N_7738,N_4099,N_4856);
xnor U7739 (N_7739,N_5099,N_4326);
nor U7740 (N_7740,N_6077,N_5820);
nor U7741 (N_7741,N_6219,N_3195);
xnor U7742 (N_7742,N_3610,N_5446);
nand U7743 (N_7743,N_3956,N_5956);
or U7744 (N_7744,N_3681,N_3833);
or U7745 (N_7745,N_6166,N_4232);
nand U7746 (N_7746,N_6097,N_3780);
and U7747 (N_7747,N_5640,N_4569);
nor U7748 (N_7748,N_3692,N_4410);
and U7749 (N_7749,N_4081,N_5145);
nand U7750 (N_7750,N_5830,N_4383);
nand U7751 (N_7751,N_5614,N_3529);
nor U7752 (N_7752,N_5691,N_4191);
xor U7753 (N_7753,N_5285,N_3968);
nand U7754 (N_7754,N_4198,N_5516);
nand U7755 (N_7755,N_3748,N_4849);
nor U7756 (N_7756,N_4772,N_4844);
nand U7757 (N_7757,N_5350,N_5358);
nand U7758 (N_7758,N_3708,N_4024);
nand U7759 (N_7759,N_6021,N_3872);
and U7760 (N_7760,N_4851,N_3125);
nor U7761 (N_7761,N_5291,N_3950);
or U7762 (N_7762,N_3303,N_5635);
or U7763 (N_7763,N_4626,N_3356);
nand U7764 (N_7764,N_6084,N_5376);
or U7765 (N_7765,N_5087,N_3910);
nor U7766 (N_7766,N_3132,N_3444);
nor U7767 (N_7767,N_3839,N_4742);
and U7768 (N_7768,N_4708,N_5399);
or U7769 (N_7769,N_4671,N_5158);
or U7770 (N_7770,N_5769,N_4181);
nor U7771 (N_7771,N_4133,N_4921);
nand U7772 (N_7772,N_5078,N_6081);
or U7773 (N_7773,N_5191,N_3932);
nand U7774 (N_7774,N_5384,N_6198);
and U7775 (N_7775,N_4903,N_4571);
or U7776 (N_7776,N_5876,N_4101);
xor U7777 (N_7777,N_5667,N_4777);
and U7778 (N_7778,N_3157,N_5073);
and U7779 (N_7779,N_3548,N_5199);
nor U7780 (N_7780,N_5510,N_4162);
nand U7781 (N_7781,N_5488,N_5790);
or U7782 (N_7782,N_3178,N_4911);
nor U7783 (N_7783,N_3706,N_4146);
nand U7784 (N_7784,N_3948,N_4422);
or U7785 (N_7785,N_4291,N_5781);
xor U7786 (N_7786,N_4697,N_3802);
nor U7787 (N_7787,N_6237,N_5371);
xor U7788 (N_7788,N_5106,N_4581);
and U7789 (N_7789,N_3767,N_5136);
or U7790 (N_7790,N_6212,N_4965);
nor U7791 (N_7791,N_4454,N_5859);
nand U7792 (N_7792,N_3643,N_3464);
nand U7793 (N_7793,N_3837,N_5821);
or U7794 (N_7794,N_5340,N_4977);
nand U7795 (N_7795,N_4757,N_3745);
nor U7796 (N_7796,N_3532,N_4644);
or U7797 (N_7797,N_4655,N_5613);
nand U7798 (N_7798,N_4495,N_4312);
xor U7799 (N_7799,N_5494,N_5690);
or U7800 (N_7800,N_5026,N_3891);
xor U7801 (N_7801,N_4117,N_4216);
and U7802 (N_7802,N_3931,N_6078);
nand U7803 (N_7803,N_5389,N_5105);
nand U7804 (N_7804,N_5961,N_4377);
and U7805 (N_7805,N_5174,N_3503);
nand U7806 (N_7806,N_3588,N_5273);
and U7807 (N_7807,N_5694,N_3855);
or U7808 (N_7808,N_3350,N_5293);
xnor U7809 (N_7809,N_4028,N_4353);
or U7810 (N_7810,N_4355,N_3657);
xor U7811 (N_7811,N_5254,N_5805);
nand U7812 (N_7812,N_4035,N_4537);
or U7813 (N_7813,N_4869,N_5729);
and U7814 (N_7814,N_4315,N_5048);
nor U7815 (N_7815,N_5883,N_3457);
xor U7816 (N_7816,N_3292,N_5273);
xor U7817 (N_7817,N_4209,N_3476);
xnor U7818 (N_7818,N_6039,N_4688);
or U7819 (N_7819,N_5816,N_4219);
nand U7820 (N_7820,N_5944,N_5856);
and U7821 (N_7821,N_5110,N_4239);
nand U7822 (N_7822,N_6112,N_5291);
xor U7823 (N_7823,N_5730,N_4585);
or U7824 (N_7824,N_5589,N_3717);
and U7825 (N_7825,N_4024,N_3979);
or U7826 (N_7826,N_4110,N_3907);
and U7827 (N_7827,N_4175,N_3516);
nand U7828 (N_7828,N_5609,N_5572);
xor U7829 (N_7829,N_4767,N_4647);
and U7830 (N_7830,N_3587,N_5441);
xor U7831 (N_7831,N_5889,N_5253);
xnor U7832 (N_7832,N_4930,N_3927);
nor U7833 (N_7833,N_4723,N_3485);
or U7834 (N_7834,N_5068,N_3532);
and U7835 (N_7835,N_6086,N_4738);
and U7836 (N_7836,N_4578,N_5724);
nand U7837 (N_7837,N_5704,N_5097);
xnor U7838 (N_7838,N_5571,N_5507);
xor U7839 (N_7839,N_3746,N_5299);
or U7840 (N_7840,N_4651,N_4927);
and U7841 (N_7841,N_5129,N_4634);
nand U7842 (N_7842,N_4710,N_3989);
and U7843 (N_7843,N_3676,N_5943);
xnor U7844 (N_7844,N_3921,N_4024);
nand U7845 (N_7845,N_5991,N_3485);
xnor U7846 (N_7846,N_4379,N_4470);
xnor U7847 (N_7847,N_6017,N_5696);
and U7848 (N_7848,N_3784,N_4786);
and U7849 (N_7849,N_4804,N_3810);
or U7850 (N_7850,N_3786,N_3530);
xor U7851 (N_7851,N_3187,N_4854);
nor U7852 (N_7852,N_3650,N_5129);
xor U7853 (N_7853,N_4821,N_6201);
or U7854 (N_7854,N_3934,N_5913);
and U7855 (N_7855,N_5956,N_4939);
nand U7856 (N_7856,N_5604,N_4774);
xnor U7857 (N_7857,N_4847,N_5949);
nor U7858 (N_7858,N_4477,N_4795);
and U7859 (N_7859,N_3429,N_5087);
xnor U7860 (N_7860,N_3637,N_5322);
nor U7861 (N_7861,N_3555,N_3364);
nand U7862 (N_7862,N_6007,N_3603);
and U7863 (N_7863,N_3341,N_6088);
xor U7864 (N_7864,N_5024,N_3931);
xor U7865 (N_7865,N_6108,N_5138);
nor U7866 (N_7866,N_3342,N_5465);
and U7867 (N_7867,N_5001,N_3320);
nand U7868 (N_7868,N_3750,N_3627);
nor U7869 (N_7869,N_3234,N_3877);
or U7870 (N_7870,N_6211,N_4696);
nand U7871 (N_7871,N_3593,N_4365);
xor U7872 (N_7872,N_5183,N_3958);
and U7873 (N_7873,N_4642,N_3575);
and U7874 (N_7874,N_5870,N_4675);
or U7875 (N_7875,N_4636,N_3150);
nor U7876 (N_7876,N_5765,N_3362);
xor U7877 (N_7877,N_4917,N_6135);
and U7878 (N_7878,N_4289,N_5787);
nand U7879 (N_7879,N_3714,N_3973);
xnor U7880 (N_7880,N_3325,N_6224);
nor U7881 (N_7881,N_5237,N_4917);
xor U7882 (N_7882,N_4621,N_5147);
and U7883 (N_7883,N_5779,N_4803);
and U7884 (N_7884,N_4650,N_4845);
nand U7885 (N_7885,N_5679,N_5759);
nor U7886 (N_7886,N_3534,N_5786);
or U7887 (N_7887,N_4462,N_3216);
nor U7888 (N_7888,N_5519,N_4433);
xor U7889 (N_7889,N_5939,N_4447);
and U7890 (N_7890,N_5375,N_4537);
nor U7891 (N_7891,N_3722,N_5463);
xnor U7892 (N_7892,N_3735,N_5594);
or U7893 (N_7893,N_3155,N_5771);
xnor U7894 (N_7894,N_6221,N_4296);
xor U7895 (N_7895,N_3556,N_4057);
xor U7896 (N_7896,N_3639,N_5459);
and U7897 (N_7897,N_4161,N_4398);
nor U7898 (N_7898,N_5883,N_3351);
and U7899 (N_7899,N_6107,N_3722);
nor U7900 (N_7900,N_5896,N_3655);
or U7901 (N_7901,N_5900,N_3860);
nor U7902 (N_7902,N_5202,N_4135);
xnor U7903 (N_7903,N_4198,N_3460);
xor U7904 (N_7904,N_5157,N_5780);
or U7905 (N_7905,N_5724,N_3434);
xnor U7906 (N_7906,N_3277,N_4036);
nor U7907 (N_7907,N_4869,N_4695);
and U7908 (N_7908,N_3694,N_4554);
or U7909 (N_7909,N_4034,N_5260);
xor U7910 (N_7910,N_3562,N_5404);
or U7911 (N_7911,N_4488,N_3715);
nand U7912 (N_7912,N_3209,N_3156);
nor U7913 (N_7913,N_4582,N_4848);
xor U7914 (N_7914,N_3789,N_5680);
xor U7915 (N_7915,N_6001,N_5422);
xnor U7916 (N_7916,N_4737,N_4305);
xnor U7917 (N_7917,N_4176,N_5370);
xor U7918 (N_7918,N_3469,N_6109);
nand U7919 (N_7919,N_3989,N_4090);
nand U7920 (N_7920,N_4242,N_5848);
nor U7921 (N_7921,N_5913,N_5205);
and U7922 (N_7922,N_4383,N_3915);
and U7923 (N_7923,N_6117,N_5055);
or U7924 (N_7924,N_5242,N_4606);
nor U7925 (N_7925,N_3425,N_5014);
nor U7926 (N_7926,N_5140,N_5791);
nor U7927 (N_7927,N_3368,N_4620);
nor U7928 (N_7928,N_5461,N_3274);
or U7929 (N_7929,N_4925,N_3796);
or U7930 (N_7930,N_5773,N_3979);
and U7931 (N_7931,N_3751,N_5825);
or U7932 (N_7932,N_3228,N_3317);
or U7933 (N_7933,N_4772,N_3130);
and U7934 (N_7934,N_5559,N_3932);
nor U7935 (N_7935,N_3866,N_6091);
nand U7936 (N_7936,N_4428,N_4193);
or U7937 (N_7937,N_6168,N_5385);
nand U7938 (N_7938,N_5867,N_4242);
and U7939 (N_7939,N_5611,N_5031);
xnor U7940 (N_7940,N_5135,N_3190);
and U7941 (N_7941,N_6116,N_4115);
xor U7942 (N_7942,N_4787,N_3364);
or U7943 (N_7943,N_4630,N_4019);
and U7944 (N_7944,N_5433,N_3143);
nand U7945 (N_7945,N_4829,N_5690);
xor U7946 (N_7946,N_3674,N_4192);
and U7947 (N_7947,N_5514,N_5700);
xnor U7948 (N_7948,N_3282,N_3747);
nor U7949 (N_7949,N_5779,N_3980);
nand U7950 (N_7950,N_6118,N_5770);
nor U7951 (N_7951,N_5358,N_4078);
or U7952 (N_7952,N_4531,N_5021);
or U7953 (N_7953,N_3923,N_3989);
nor U7954 (N_7954,N_3747,N_3394);
nand U7955 (N_7955,N_3535,N_4791);
nor U7956 (N_7956,N_4467,N_5095);
nand U7957 (N_7957,N_5931,N_4202);
and U7958 (N_7958,N_5059,N_3615);
xnor U7959 (N_7959,N_4072,N_4655);
or U7960 (N_7960,N_4850,N_4804);
or U7961 (N_7961,N_3863,N_5612);
nand U7962 (N_7962,N_4026,N_6141);
xor U7963 (N_7963,N_5170,N_4640);
nand U7964 (N_7964,N_5347,N_4974);
and U7965 (N_7965,N_4901,N_3726);
xnor U7966 (N_7966,N_3557,N_5875);
and U7967 (N_7967,N_5764,N_5618);
and U7968 (N_7968,N_4576,N_5117);
nor U7969 (N_7969,N_4711,N_3986);
and U7970 (N_7970,N_3356,N_4311);
nand U7971 (N_7971,N_6189,N_5163);
nand U7972 (N_7972,N_5255,N_5357);
xor U7973 (N_7973,N_4162,N_4405);
or U7974 (N_7974,N_3644,N_4275);
nor U7975 (N_7975,N_5966,N_4055);
nand U7976 (N_7976,N_5991,N_6198);
and U7977 (N_7977,N_5912,N_5820);
or U7978 (N_7978,N_5685,N_4556);
nor U7979 (N_7979,N_5579,N_4608);
or U7980 (N_7980,N_5348,N_5768);
nand U7981 (N_7981,N_4922,N_3345);
and U7982 (N_7982,N_4782,N_4546);
nor U7983 (N_7983,N_4216,N_5424);
and U7984 (N_7984,N_4990,N_3743);
and U7985 (N_7985,N_4635,N_4836);
nor U7986 (N_7986,N_3831,N_5784);
nor U7987 (N_7987,N_4784,N_4080);
nor U7988 (N_7988,N_3744,N_3127);
and U7989 (N_7989,N_5985,N_3836);
and U7990 (N_7990,N_5295,N_5953);
or U7991 (N_7991,N_6248,N_3309);
nor U7992 (N_7992,N_5293,N_4604);
nor U7993 (N_7993,N_4416,N_5436);
nand U7994 (N_7994,N_5975,N_5302);
xnor U7995 (N_7995,N_6246,N_4154);
nor U7996 (N_7996,N_5979,N_5643);
nand U7997 (N_7997,N_3804,N_5767);
xnor U7998 (N_7998,N_4697,N_4173);
nor U7999 (N_7999,N_6247,N_4962);
or U8000 (N_8000,N_6056,N_6148);
or U8001 (N_8001,N_5603,N_6050);
nor U8002 (N_8002,N_5981,N_3757);
xnor U8003 (N_8003,N_4554,N_3823);
xnor U8004 (N_8004,N_4737,N_5322);
nand U8005 (N_8005,N_3219,N_3314);
xor U8006 (N_8006,N_5596,N_5483);
and U8007 (N_8007,N_5216,N_3135);
nand U8008 (N_8008,N_3644,N_3333);
nand U8009 (N_8009,N_5185,N_5160);
nand U8010 (N_8010,N_3954,N_5223);
nor U8011 (N_8011,N_5728,N_4250);
nor U8012 (N_8012,N_5115,N_5296);
and U8013 (N_8013,N_3596,N_3958);
xnor U8014 (N_8014,N_4848,N_3871);
xor U8015 (N_8015,N_6147,N_3424);
nand U8016 (N_8016,N_3689,N_4328);
nand U8017 (N_8017,N_5705,N_3396);
xnor U8018 (N_8018,N_5207,N_3968);
xnor U8019 (N_8019,N_5680,N_4519);
nand U8020 (N_8020,N_5677,N_4225);
xor U8021 (N_8021,N_3484,N_3696);
or U8022 (N_8022,N_4557,N_5933);
xnor U8023 (N_8023,N_5691,N_4596);
or U8024 (N_8024,N_5824,N_4618);
nand U8025 (N_8025,N_4464,N_5150);
and U8026 (N_8026,N_4889,N_5318);
nand U8027 (N_8027,N_3370,N_5510);
nand U8028 (N_8028,N_4583,N_3664);
nor U8029 (N_8029,N_4086,N_5944);
xor U8030 (N_8030,N_5940,N_4263);
or U8031 (N_8031,N_3282,N_5745);
nand U8032 (N_8032,N_6150,N_4550);
nand U8033 (N_8033,N_4122,N_5709);
xor U8034 (N_8034,N_4617,N_5616);
xor U8035 (N_8035,N_5529,N_4360);
xnor U8036 (N_8036,N_3429,N_4188);
nor U8037 (N_8037,N_3204,N_3298);
nand U8038 (N_8038,N_4773,N_4565);
nand U8039 (N_8039,N_4193,N_6224);
or U8040 (N_8040,N_3261,N_4785);
or U8041 (N_8041,N_4821,N_4067);
or U8042 (N_8042,N_4407,N_4233);
or U8043 (N_8043,N_5327,N_3164);
nand U8044 (N_8044,N_4191,N_5638);
nand U8045 (N_8045,N_5946,N_5731);
nor U8046 (N_8046,N_3179,N_5379);
and U8047 (N_8047,N_5823,N_6128);
and U8048 (N_8048,N_4850,N_5982);
xnor U8049 (N_8049,N_3869,N_3134);
nand U8050 (N_8050,N_6190,N_5648);
and U8051 (N_8051,N_5126,N_3178);
and U8052 (N_8052,N_3260,N_5536);
and U8053 (N_8053,N_5407,N_3156);
nand U8054 (N_8054,N_4267,N_5010);
xor U8055 (N_8055,N_5563,N_5932);
xor U8056 (N_8056,N_4537,N_5142);
nand U8057 (N_8057,N_5256,N_6027);
or U8058 (N_8058,N_6027,N_3917);
or U8059 (N_8059,N_5649,N_3186);
nor U8060 (N_8060,N_3878,N_4165);
or U8061 (N_8061,N_3769,N_4576);
nand U8062 (N_8062,N_5917,N_4601);
xnor U8063 (N_8063,N_4366,N_5249);
nor U8064 (N_8064,N_6172,N_4173);
or U8065 (N_8065,N_5351,N_4742);
nand U8066 (N_8066,N_5811,N_3913);
or U8067 (N_8067,N_3125,N_3378);
and U8068 (N_8068,N_4020,N_5473);
xor U8069 (N_8069,N_3241,N_5317);
nor U8070 (N_8070,N_4831,N_3880);
or U8071 (N_8071,N_6057,N_4271);
and U8072 (N_8072,N_4552,N_3395);
nand U8073 (N_8073,N_3739,N_5581);
or U8074 (N_8074,N_3875,N_4037);
xor U8075 (N_8075,N_3869,N_3775);
or U8076 (N_8076,N_5199,N_5358);
or U8077 (N_8077,N_5935,N_6220);
nand U8078 (N_8078,N_5252,N_4498);
nand U8079 (N_8079,N_3908,N_5770);
and U8080 (N_8080,N_4908,N_5190);
nand U8081 (N_8081,N_5835,N_3551);
or U8082 (N_8082,N_3681,N_5619);
nand U8083 (N_8083,N_5840,N_5783);
nand U8084 (N_8084,N_5504,N_3672);
nor U8085 (N_8085,N_5233,N_3742);
nor U8086 (N_8086,N_3440,N_4517);
nand U8087 (N_8087,N_5927,N_3485);
or U8088 (N_8088,N_3160,N_3468);
and U8089 (N_8089,N_4588,N_4470);
nand U8090 (N_8090,N_4060,N_5119);
nand U8091 (N_8091,N_6033,N_5742);
nor U8092 (N_8092,N_5043,N_4462);
or U8093 (N_8093,N_5237,N_6052);
or U8094 (N_8094,N_4571,N_5610);
nor U8095 (N_8095,N_6006,N_3143);
nor U8096 (N_8096,N_3881,N_3294);
xnor U8097 (N_8097,N_3308,N_5473);
nand U8098 (N_8098,N_3456,N_5465);
nand U8099 (N_8099,N_4683,N_3759);
nand U8100 (N_8100,N_4137,N_5035);
or U8101 (N_8101,N_5358,N_4522);
or U8102 (N_8102,N_5241,N_3982);
and U8103 (N_8103,N_4172,N_5555);
and U8104 (N_8104,N_4007,N_5940);
xnor U8105 (N_8105,N_4309,N_6137);
nand U8106 (N_8106,N_5403,N_6007);
nand U8107 (N_8107,N_5292,N_5926);
nand U8108 (N_8108,N_4902,N_6085);
nor U8109 (N_8109,N_5966,N_3319);
xnor U8110 (N_8110,N_3614,N_4806);
nor U8111 (N_8111,N_4298,N_4894);
and U8112 (N_8112,N_4385,N_3747);
or U8113 (N_8113,N_6248,N_5630);
nor U8114 (N_8114,N_5897,N_4327);
nor U8115 (N_8115,N_5356,N_3416);
nor U8116 (N_8116,N_5348,N_5746);
nor U8117 (N_8117,N_4324,N_5963);
or U8118 (N_8118,N_4415,N_4892);
xor U8119 (N_8119,N_3539,N_4277);
or U8120 (N_8120,N_3205,N_4395);
xnor U8121 (N_8121,N_6189,N_3336);
or U8122 (N_8122,N_6229,N_3613);
nand U8123 (N_8123,N_5804,N_4708);
nand U8124 (N_8124,N_6115,N_4499);
nor U8125 (N_8125,N_5604,N_3653);
or U8126 (N_8126,N_4742,N_5547);
and U8127 (N_8127,N_4337,N_3685);
or U8128 (N_8128,N_6211,N_4753);
and U8129 (N_8129,N_5302,N_5134);
nor U8130 (N_8130,N_4695,N_4975);
and U8131 (N_8131,N_5039,N_5082);
and U8132 (N_8132,N_4713,N_3620);
or U8133 (N_8133,N_3920,N_4651);
or U8134 (N_8134,N_3736,N_3290);
nand U8135 (N_8135,N_5195,N_5370);
nand U8136 (N_8136,N_4066,N_3277);
nor U8137 (N_8137,N_5244,N_4669);
nand U8138 (N_8138,N_3356,N_3217);
xor U8139 (N_8139,N_4242,N_5266);
nand U8140 (N_8140,N_4317,N_3300);
nand U8141 (N_8141,N_3197,N_3504);
or U8142 (N_8142,N_3903,N_3372);
or U8143 (N_8143,N_5080,N_5829);
and U8144 (N_8144,N_3919,N_4066);
nor U8145 (N_8145,N_5028,N_3505);
nand U8146 (N_8146,N_5469,N_3893);
nand U8147 (N_8147,N_5331,N_4674);
xnor U8148 (N_8148,N_5615,N_4380);
xor U8149 (N_8149,N_5387,N_6074);
or U8150 (N_8150,N_4178,N_3970);
or U8151 (N_8151,N_5534,N_5864);
xor U8152 (N_8152,N_4081,N_3198);
nand U8153 (N_8153,N_5140,N_5125);
nor U8154 (N_8154,N_5058,N_3310);
nand U8155 (N_8155,N_3995,N_6206);
xnor U8156 (N_8156,N_4986,N_4413);
and U8157 (N_8157,N_6097,N_4990);
nor U8158 (N_8158,N_4083,N_3220);
nor U8159 (N_8159,N_5382,N_3708);
nand U8160 (N_8160,N_3759,N_4841);
xor U8161 (N_8161,N_3983,N_3990);
xor U8162 (N_8162,N_4327,N_4803);
xnor U8163 (N_8163,N_3667,N_3748);
or U8164 (N_8164,N_4670,N_6066);
or U8165 (N_8165,N_4631,N_5698);
or U8166 (N_8166,N_5476,N_4675);
nand U8167 (N_8167,N_5386,N_3128);
nor U8168 (N_8168,N_4093,N_3710);
and U8169 (N_8169,N_3422,N_5730);
nand U8170 (N_8170,N_3969,N_3488);
nor U8171 (N_8171,N_4444,N_4701);
xor U8172 (N_8172,N_4742,N_3930);
and U8173 (N_8173,N_5946,N_4388);
xnor U8174 (N_8174,N_6184,N_5202);
nor U8175 (N_8175,N_5132,N_4804);
and U8176 (N_8176,N_5550,N_6143);
xnor U8177 (N_8177,N_3568,N_3644);
nor U8178 (N_8178,N_4241,N_5050);
nand U8179 (N_8179,N_4887,N_6190);
xor U8180 (N_8180,N_4603,N_5400);
nor U8181 (N_8181,N_4685,N_3814);
nand U8182 (N_8182,N_3768,N_5873);
or U8183 (N_8183,N_4398,N_5544);
nand U8184 (N_8184,N_4240,N_4308);
xor U8185 (N_8185,N_3674,N_6152);
nand U8186 (N_8186,N_5554,N_4105);
nor U8187 (N_8187,N_3999,N_3513);
xor U8188 (N_8188,N_3765,N_4613);
and U8189 (N_8189,N_4303,N_5277);
and U8190 (N_8190,N_5462,N_4224);
nor U8191 (N_8191,N_5869,N_3787);
nand U8192 (N_8192,N_5803,N_3501);
or U8193 (N_8193,N_3641,N_5815);
nor U8194 (N_8194,N_5907,N_4250);
nand U8195 (N_8195,N_5080,N_3603);
nand U8196 (N_8196,N_3747,N_3208);
nand U8197 (N_8197,N_5136,N_4488);
and U8198 (N_8198,N_4669,N_3348);
and U8199 (N_8199,N_5779,N_5306);
nor U8200 (N_8200,N_3267,N_4896);
xnor U8201 (N_8201,N_4699,N_5277);
xnor U8202 (N_8202,N_5650,N_5902);
nor U8203 (N_8203,N_4619,N_5472);
xor U8204 (N_8204,N_3380,N_5995);
nor U8205 (N_8205,N_4158,N_4113);
xor U8206 (N_8206,N_4013,N_3937);
or U8207 (N_8207,N_4383,N_4294);
xor U8208 (N_8208,N_4667,N_5425);
nor U8209 (N_8209,N_4295,N_4336);
nand U8210 (N_8210,N_4147,N_3781);
nor U8211 (N_8211,N_3385,N_6239);
nand U8212 (N_8212,N_6074,N_6054);
and U8213 (N_8213,N_3721,N_3809);
xnor U8214 (N_8214,N_5262,N_5781);
and U8215 (N_8215,N_5314,N_5891);
and U8216 (N_8216,N_5375,N_3176);
xor U8217 (N_8217,N_5720,N_4454);
nand U8218 (N_8218,N_4552,N_4690);
and U8219 (N_8219,N_4772,N_4018);
nand U8220 (N_8220,N_6108,N_5260);
or U8221 (N_8221,N_5852,N_4555);
or U8222 (N_8222,N_4486,N_3379);
nor U8223 (N_8223,N_3635,N_3378);
nor U8224 (N_8224,N_4933,N_3282);
nand U8225 (N_8225,N_5869,N_4420);
and U8226 (N_8226,N_5141,N_4713);
xor U8227 (N_8227,N_5172,N_5229);
nor U8228 (N_8228,N_4720,N_3664);
nor U8229 (N_8229,N_5715,N_5570);
xnor U8230 (N_8230,N_4580,N_5104);
nor U8231 (N_8231,N_4259,N_5922);
xor U8232 (N_8232,N_5790,N_3620);
xnor U8233 (N_8233,N_3911,N_4818);
nand U8234 (N_8234,N_5394,N_5848);
nand U8235 (N_8235,N_3436,N_4788);
or U8236 (N_8236,N_3844,N_6042);
and U8237 (N_8237,N_3560,N_6022);
and U8238 (N_8238,N_6068,N_3206);
nor U8239 (N_8239,N_3610,N_5534);
nor U8240 (N_8240,N_5661,N_5217);
xor U8241 (N_8241,N_4317,N_5121);
nand U8242 (N_8242,N_5139,N_5569);
and U8243 (N_8243,N_6171,N_5928);
xnor U8244 (N_8244,N_4595,N_4104);
or U8245 (N_8245,N_6127,N_4586);
or U8246 (N_8246,N_4155,N_3802);
xnor U8247 (N_8247,N_4582,N_5251);
or U8248 (N_8248,N_3503,N_5557);
xnor U8249 (N_8249,N_3166,N_4608);
and U8250 (N_8250,N_5849,N_4801);
xnor U8251 (N_8251,N_4723,N_4632);
and U8252 (N_8252,N_3790,N_4615);
nand U8253 (N_8253,N_4567,N_4318);
or U8254 (N_8254,N_4124,N_3626);
nand U8255 (N_8255,N_5227,N_3409);
xnor U8256 (N_8256,N_3952,N_5122);
or U8257 (N_8257,N_4025,N_4747);
nand U8258 (N_8258,N_4746,N_5712);
and U8259 (N_8259,N_5374,N_4037);
and U8260 (N_8260,N_6193,N_5807);
xnor U8261 (N_8261,N_5577,N_3372);
xor U8262 (N_8262,N_3813,N_3253);
nand U8263 (N_8263,N_3450,N_4980);
or U8264 (N_8264,N_6238,N_5095);
xnor U8265 (N_8265,N_5338,N_3666);
xor U8266 (N_8266,N_3894,N_3553);
nor U8267 (N_8267,N_4043,N_3252);
nand U8268 (N_8268,N_3284,N_5635);
or U8269 (N_8269,N_5169,N_5761);
and U8270 (N_8270,N_3249,N_5428);
nand U8271 (N_8271,N_6180,N_3951);
or U8272 (N_8272,N_6033,N_4584);
or U8273 (N_8273,N_4086,N_4122);
xor U8274 (N_8274,N_3434,N_6168);
nand U8275 (N_8275,N_4910,N_4129);
nand U8276 (N_8276,N_4137,N_5265);
and U8277 (N_8277,N_4485,N_5164);
and U8278 (N_8278,N_5579,N_5528);
xor U8279 (N_8279,N_5976,N_5346);
nand U8280 (N_8280,N_4084,N_4272);
nor U8281 (N_8281,N_4184,N_3914);
xor U8282 (N_8282,N_4612,N_3562);
or U8283 (N_8283,N_4568,N_5553);
and U8284 (N_8284,N_5627,N_3438);
nand U8285 (N_8285,N_4264,N_4346);
xor U8286 (N_8286,N_4887,N_3427);
and U8287 (N_8287,N_4904,N_3440);
xor U8288 (N_8288,N_4595,N_4288);
nand U8289 (N_8289,N_3651,N_4654);
and U8290 (N_8290,N_3954,N_5743);
xnor U8291 (N_8291,N_4046,N_4223);
xnor U8292 (N_8292,N_5508,N_5947);
xnor U8293 (N_8293,N_5524,N_3828);
nand U8294 (N_8294,N_4700,N_4552);
nand U8295 (N_8295,N_6099,N_4961);
and U8296 (N_8296,N_4875,N_5423);
nor U8297 (N_8297,N_3318,N_5996);
or U8298 (N_8298,N_3925,N_5470);
xor U8299 (N_8299,N_5358,N_3412);
and U8300 (N_8300,N_5556,N_4119);
xnor U8301 (N_8301,N_5727,N_4028);
nand U8302 (N_8302,N_3373,N_3125);
nand U8303 (N_8303,N_3670,N_5452);
nand U8304 (N_8304,N_5450,N_3564);
nor U8305 (N_8305,N_3360,N_3304);
nand U8306 (N_8306,N_5958,N_6224);
xor U8307 (N_8307,N_6206,N_4140);
xnor U8308 (N_8308,N_4711,N_5055);
or U8309 (N_8309,N_4963,N_3906);
nor U8310 (N_8310,N_3822,N_4242);
nand U8311 (N_8311,N_4437,N_4469);
and U8312 (N_8312,N_5023,N_4385);
nand U8313 (N_8313,N_3605,N_3667);
and U8314 (N_8314,N_4936,N_5443);
xnor U8315 (N_8315,N_4114,N_4548);
and U8316 (N_8316,N_4636,N_4884);
nor U8317 (N_8317,N_4849,N_4725);
nand U8318 (N_8318,N_4464,N_3927);
nor U8319 (N_8319,N_5795,N_4328);
or U8320 (N_8320,N_4985,N_3281);
and U8321 (N_8321,N_5675,N_3472);
nor U8322 (N_8322,N_4431,N_5570);
and U8323 (N_8323,N_5733,N_3414);
nor U8324 (N_8324,N_4394,N_5437);
or U8325 (N_8325,N_5099,N_4862);
and U8326 (N_8326,N_4507,N_4471);
nand U8327 (N_8327,N_3154,N_4271);
xor U8328 (N_8328,N_5475,N_3314);
and U8329 (N_8329,N_4364,N_3671);
xor U8330 (N_8330,N_4326,N_3715);
nor U8331 (N_8331,N_4503,N_5277);
and U8332 (N_8332,N_5271,N_5355);
and U8333 (N_8333,N_5580,N_3867);
nand U8334 (N_8334,N_5368,N_3128);
nand U8335 (N_8335,N_4700,N_3645);
nor U8336 (N_8336,N_3959,N_3296);
xnor U8337 (N_8337,N_5739,N_4829);
xor U8338 (N_8338,N_5544,N_5247);
nor U8339 (N_8339,N_4688,N_3994);
and U8340 (N_8340,N_3281,N_4983);
nor U8341 (N_8341,N_3862,N_6201);
xor U8342 (N_8342,N_5335,N_5304);
nor U8343 (N_8343,N_5984,N_4007);
xnor U8344 (N_8344,N_3697,N_5170);
nor U8345 (N_8345,N_6000,N_6199);
and U8346 (N_8346,N_6066,N_6182);
xor U8347 (N_8347,N_4065,N_3410);
or U8348 (N_8348,N_3441,N_3785);
nor U8349 (N_8349,N_5051,N_5204);
xor U8350 (N_8350,N_4430,N_4389);
nor U8351 (N_8351,N_3131,N_4780);
or U8352 (N_8352,N_4243,N_4147);
or U8353 (N_8353,N_4742,N_5975);
xor U8354 (N_8354,N_3149,N_4050);
xnor U8355 (N_8355,N_4306,N_5385);
nand U8356 (N_8356,N_5928,N_4685);
and U8357 (N_8357,N_4924,N_5916);
and U8358 (N_8358,N_5169,N_5162);
or U8359 (N_8359,N_4980,N_3176);
nor U8360 (N_8360,N_3903,N_5300);
xnor U8361 (N_8361,N_4747,N_5644);
xor U8362 (N_8362,N_5171,N_3368);
xnor U8363 (N_8363,N_3148,N_4522);
or U8364 (N_8364,N_3622,N_5093);
and U8365 (N_8365,N_3444,N_5497);
xnor U8366 (N_8366,N_3901,N_3313);
and U8367 (N_8367,N_3367,N_5872);
xnor U8368 (N_8368,N_4608,N_5249);
and U8369 (N_8369,N_4702,N_4661);
nand U8370 (N_8370,N_5098,N_4348);
nand U8371 (N_8371,N_5328,N_3621);
or U8372 (N_8372,N_3749,N_5368);
nand U8373 (N_8373,N_4621,N_5095);
nand U8374 (N_8374,N_6044,N_5686);
and U8375 (N_8375,N_4013,N_5882);
xnor U8376 (N_8376,N_5417,N_5129);
nor U8377 (N_8377,N_5172,N_4379);
xor U8378 (N_8378,N_4285,N_5936);
xnor U8379 (N_8379,N_3589,N_4856);
nand U8380 (N_8380,N_5032,N_5360);
xor U8381 (N_8381,N_6047,N_4853);
nand U8382 (N_8382,N_5243,N_4312);
or U8383 (N_8383,N_5331,N_4792);
nor U8384 (N_8384,N_5268,N_4977);
nand U8385 (N_8385,N_3398,N_4135);
or U8386 (N_8386,N_6220,N_4377);
xor U8387 (N_8387,N_3568,N_3512);
nand U8388 (N_8388,N_4353,N_3443);
xor U8389 (N_8389,N_4424,N_5893);
xor U8390 (N_8390,N_5540,N_5219);
or U8391 (N_8391,N_5427,N_5059);
or U8392 (N_8392,N_4964,N_4539);
and U8393 (N_8393,N_4592,N_3858);
nor U8394 (N_8394,N_4594,N_3593);
xor U8395 (N_8395,N_5430,N_5042);
nand U8396 (N_8396,N_5583,N_4208);
xnor U8397 (N_8397,N_4487,N_4211);
and U8398 (N_8398,N_3295,N_5702);
nor U8399 (N_8399,N_4112,N_3328);
nand U8400 (N_8400,N_5417,N_5738);
nand U8401 (N_8401,N_6233,N_4171);
xor U8402 (N_8402,N_5155,N_3382);
and U8403 (N_8403,N_3740,N_3343);
xnor U8404 (N_8404,N_4623,N_3938);
and U8405 (N_8405,N_4541,N_4208);
or U8406 (N_8406,N_5745,N_5247);
or U8407 (N_8407,N_5079,N_5175);
nand U8408 (N_8408,N_4134,N_5112);
nand U8409 (N_8409,N_4445,N_4606);
nand U8410 (N_8410,N_3480,N_3484);
xnor U8411 (N_8411,N_4496,N_3393);
nor U8412 (N_8412,N_3847,N_3391);
nand U8413 (N_8413,N_5453,N_5026);
nand U8414 (N_8414,N_5185,N_3759);
or U8415 (N_8415,N_5698,N_3489);
xnor U8416 (N_8416,N_6001,N_4376);
xor U8417 (N_8417,N_4905,N_4871);
or U8418 (N_8418,N_5889,N_4706);
xnor U8419 (N_8419,N_4551,N_5553);
or U8420 (N_8420,N_5737,N_4981);
xor U8421 (N_8421,N_3973,N_4110);
or U8422 (N_8422,N_4021,N_4115);
nor U8423 (N_8423,N_3566,N_4578);
and U8424 (N_8424,N_6197,N_6180);
or U8425 (N_8425,N_4126,N_3660);
xnor U8426 (N_8426,N_4427,N_5269);
xnor U8427 (N_8427,N_6008,N_5400);
nor U8428 (N_8428,N_3217,N_5432);
xor U8429 (N_8429,N_4357,N_4948);
or U8430 (N_8430,N_3296,N_4119);
nand U8431 (N_8431,N_3327,N_6192);
nor U8432 (N_8432,N_5420,N_4842);
xor U8433 (N_8433,N_5681,N_3381);
xor U8434 (N_8434,N_4303,N_3546);
or U8435 (N_8435,N_4531,N_4298);
xor U8436 (N_8436,N_3411,N_4452);
xnor U8437 (N_8437,N_4755,N_6116);
xor U8438 (N_8438,N_3242,N_4175);
nand U8439 (N_8439,N_4383,N_4410);
xor U8440 (N_8440,N_3814,N_5879);
xor U8441 (N_8441,N_4262,N_3447);
nor U8442 (N_8442,N_4789,N_4729);
and U8443 (N_8443,N_3416,N_3572);
and U8444 (N_8444,N_6057,N_5499);
and U8445 (N_8445,N_4109,N_3784);
nand U8446 (N_8446,N_4845,N_4688);
nand U8447 (N_8447,N_4428,N_3244);
and U8448 (N_8448,N_3166,N_3788);
nor U8449 (N_8449,N_3700,N_3979);
or U8450 (N_8450,N_4296,N_4622);
nor U8451 (N_8451,N_6224,N_3227);
and U8452 (N_8452,N_4862,N_5119);
xnor U8453 (N_8453,N_3674,N_4919);
or U8454 (N_8454,N_3800,N_6019);
and U8455 (N_8455,N_3530,N_5575);
or U8456 (N_8456,N_5134,N_5180);
xor U8457 (N_8457,N_4552,N_5129);
nor U8458 (N_8458,N_3765,N_4249);
and U8459 (N_8459,N_3936,N_4250);
xnor U8460 (N_8460,N_4904,N_4260);
or U8461 (N_8461,N_4151,N_3224);
or U8462 (N_8462,N_5695,N_5346);
and U8463 (N_8463,N_3304,N_5333);
or U8464 (N_8464,N_3597,N_3824);
or U8465 (N_8465,N_5908,N_3942);
and U8466 (N_8466,N_4480,N_3279);
nor U8467 (N_8467,N_4786,N_5574);
xor U8468 (N_8468,N_4481,N_3440);
xnor U8469 (N_8469,N_4773,N_6226);
nand U8470 (N_8470,N_4911,N_4398);
xnor U8471 (N_8471,N_5930,N_3185);
nand U8472 (N_8472,N_3157,N_4465);
nand U8473 (N_8473,N_4583,N_3896);
and U8474 (N_8474,N_3949,N_3347);
and U8475 (N_8475,N_5870,N_5708);
xnor U8476 (N_8476,N_6152,N_5330);
xnor U8477 (N_8477,N_5966,N_4415);
or U8478 (N_8478,N_5957,N_6020);
nor U8479 (N_8479,N_4181,N_5782);
nor U8480 (N_8480,N_5235,N_5435);
nor U8481 (N_8481,N_3597,N_5450);
nor U8482 (N_8482,N_3923,N_4045);
xor U8483 (N_8483,N_6249,N_6157);
nor U8484 (N_8484,N_4787,N_5303);
or U8485 (N_8485,N_4599,N_4662);
xnor U8486 (N_8486,N_3430,N_3183);
or U8487 (N_8487,N_3319,N_3271);
or U8488 (N_8488,N_3667,N_4107);
nand U8489 (N_8489,N_3780,N_4463);
or U8490 (N_8490,N_4267,N_5070);
and U8491 (N_8491,N_4659,N_5225);
xor U8492 (N_8492,N_3573,N_4473);
nor U8493 (N_8493,N_3919,N_6056);
nand U8494 (N_8494,N_4689,N_4079);
and U8495 (N_8495,N_6036,N_3751);
nor U8496 (N_8496,N_4378,N_5759);
xnor U8497 (N_8497,N_4150,N_5310);
and U8498 (N_8498,N_3921,N_3932);
nand U8499 (N_8499,N_4542,N_4325);
nand U8500 (N_8500,N_4454,N_4612);
nor U8501 (N_8501,N_4979,N_5524);
nand U8502 (N_8502,N_4717,N_3579);
or U8503 (N_8503,N_5894,N_5880);
or U8504 (N_8504,N_3908,N_4128);
nand U8505 (N_8505,N_4726,N_3295);
and U8506 (N_8506,N_5823,N_3776);
xnor U8507 (N_8507,N_4459,N_5796);
nand U8508 (N_8508,N_3543,N_3675);
and U8509 (N_8509,N_6046,N_4626);
xnor U8510 (N_8510,N_3496,N_4520);
nor U8511 (N_8511,N_6043,N_3812);
nand U8512 (N_8512,N_4045,N_4655);
or U8513 (N_8513,N_5596,N_4975);
xnor U8514 (N_8514,N_4740,N_5929);
or U8515 (N_8515,N_6204,N_4489);
or U8516 (N_8516,N_4911,N_3848);
and U8517 (N_8517,N_5695,N_6088);
nor U8518 (N_8518,N_4016,N_4243);
nor U8519 (N_8519,N_4927,N_5174);
and U8520 (N_8520,N_5217,N_5693);
or U8521 (N_8521,N_5313,N_4088);
nand U8522 (N_8522,N_4501,N_4848);
nand U8523 (N_8523,N_3688,N_5173);
or U8524 (N_8524,N_5482,N_3621);
and U8525 (N_8525,N_6096,N_3550);
xnor U8526 (N_8526,N_4306,N_3678);
nand U8527 (N_8527,N_6029,N_5343);
or U8528 (N_8528,N_5148,N_3354);
nor U8529 (N_8529,N_5993,N_3981);
nand U8530 (N_8530,N_3181,N_4549);
and U8531 (N_8531,N_4319,N_3496);
nor U8532 (N_8532,N_3926,N_4338);
or U8533 (N_8533,N_3877,N_3751);
nand U8534 (N_8534,N_6042,N_3744);
or U8535 (N_8535,N_4013,N_3825);
nor U8536 (N_8536,N_5760,N_5064);
or U8537 (N_8537,N_4207,N_4300);
nand U8538 (N_8538,N_5821,N_4839);
nand U8539 (N_8539,N_3794,N_4141);
xor U8540 (N_8540,N_3265,N_4205);
and U8541 (N_8541,N_4695,N_5183);
nand U8542 (N_8542,N_3897,N_3369);
xnor U8543 (N_8543,N_5028,N_4593);
or U8544 (N_8544,N_3747,N_5999);
nand U8545 (N_8545,N_4118,N_4877);
or U8546 (N_8546,N_3360,N_4393);
or U8547 (N_8547,N_6133,N_5985);
and U8548 (N_8548,N_5775,N_6199);
nand U8549 (N_8549,N_3425,N_4326);
or U8550 (N_8550,N_4292,N_3840);
nor U8551 (N_8551,N_5410,N_4835);
and U8552 (N_8552,N_4631,N_5331);
and U8553 (N_8553,N_5522,N_5749);
and U8554 (N_8554,N_3960,N_5479);
xor U8555 (N_8555,N_3760,N_4412);
nor U8556 (N_8556,N_5575,N_4712);
or U8557 (N_8557,N_3385,N_4900);
and U8558 (N_8558,N_4173,N_4124);
or U8559 (N_8559,N_5269,N_4355);
and U8560 (N_8560,N_5303,N_3396);
nor U8561 (N_8561,N_3403,N_5555);
xor U8562 (N_8562,N_4106,N_4252);
nand U8563 (N_8563,N_3747,N_4017);
nor U8564 (N_8564,N_5133,N_3702);
xor U8565 (N_8565,N_6222,N_4042);
and U8566 (N_8566,N_5025,N_3467);
nor U8567 (N_8567,N_3410,N_4382);
xnor U8568 (N_8568,N_3478,N_4837);
and U8569 (N_8569,N_5613,N_5387);
and U8570 (N_8570,N_5613,N_5929);
xnor U8571 (N_8571,N_3336,N_4508);
and U8572 (N_8572,N_4483,N_4099);
or U8573 (N_8573,N_5965,N_5099);
or U8574 (N_8574,N_4542,N_5807);
nor U8575 (N_8575,N_5994,N_4081);
nor U8576 (N_8576,N_3750,N_3343);
nor U8577 (N_8577,N_3281,N_6193);
and U8578 (N_8578,N_6162,N_3163);
and U8579 (N_8579,N_3376,N_5222);
or U8580 (N_8580,N_3839,N_4354);
or U8581 (N_8581,N_4998,N_4053);
or U8582 (N_8582,N_4641,N_3308);
or U8583 (N_8583,N_5730,N_4900);
xnor U8584 (N_8584,N_5228,N_4548);
and U8585 (N_8585,N_4210,N_3186);
xor U8586 (N_8586,N_4202,N_3787);
xor U8587 (N_8587,N_4554,N_6165);
or U8588 (N_8588,N_4200,N_4346);
nor U8589 (N_8589,N_5016,N_3320);
nor U8590 (N_8590,N_4931,N_6036);
xnor U8591 (N_8591,N_5728,N_5257);
nor U8592 (N_8592,N_4372,N_3298);
or U8593 (N_8593,N_4265,N_4855);
nand U8594 (N_8594,N_4908,N_5334);
nand U8595 (N_8595,N_3320,N_5477);
nand U8596 (N_8596,N_4007,N_4976);
or U8597 (N_8597,N_5172,N_3930);
nand U8598 (N_8598,N_3638,N_5833);
nand U8599 (N_8599,N_5497,N_5373);
nor U8600 (N_8600,N_5620,N_3515);
nor U8601 (N_8601,N_4427,N_5432);
nor U8602 (N_8602,N_5212,N_4224);
nor U8603 (N_8603,N_3422,N_4936);
nand U8604 (N_8604,N_3132,N_3912);
xor U8605 (N_8605,N_3152,N_3500);
nand U8606 (N_8606,N_4426,N_5975);
nand U8607 (N_8607,N_4299,N_5660);
nor U8608 (N_8608,N_3657,N_3945);
or U8609 (N_8609,N_5998,N_5777);
or U8610 (N_8610,N_3675,N_5007);
or U8611 (N_8611,N_6112,N_6026);
nor U8612 (N_8612,N_3259,N_4001);
or U8613 (N_8613,N_4925,N_5349);
nor U8614 (N_8614,N_5977,N_5497);
nand U8615 (N_8615,N_4086,N_3553);
or U8616 (N_8616,N_5321,N_5615);
or U8617 (N_8617,N_4935,N_4274);
and U8618 (N_8618,N_5821,N_5011);
xor U8619 (N_8619,N_4879,N_3614);
nor U8620 (N_8620,N_3741,N_5346);
and U8621 (N_8621,N_3585,N_3174);
or U8622 (N_8622,N_4165,N_3395);
and U8623 (N_8623,N_5269,N_4527);
nand U8624 (N_8624,N_3672,N_5985);
nand U8625 (N_8625,N_3629,N_5336);
nand U8626 (N_8626,N_5673,N_3781);
nand U8627 (N_8627,N_3270,N_5880);
xnor U8628 (N_8628,N_3269,N_5270);
nor U8629 (N_8629,N_3742,N_3636);
nand U8630 (N_8630,N_5377,N_5128);
or U8631 (N_8631,N_4600,N_3314);
nand U8632 (N_8632,N_4761,N_4314);
or U8633 (N_8633,N_4963,N_5699);
nand U8634 (N_8634,N_5118,N_5420);
nand U8635 (N_8635,N_3674,N_5725);
xnor U8636 (N_8636,N_5001,N_5062);
or U8637 (N_8637,N_3146,N_4966);
nor U8638 (N_8638,N_6178,N_3442);
nand U8639 (N_8639,N_5554,N_5380);
xnor U8640 (N_8640,N_3875,N_5976);
nand U8641 (N_8641,N_4820,N_5498);
or U8642 (N_8642,N_3468,N_3783);
nor U8643 (N_8643,N_3802,N_5120);
nand U8644 (N_8644,N_4759,N_3968);
nand U8645 (N_8645,N_5966,N_5714);
xor U8646 (N_8646,N_5914,N_6164);
nor U8647 (N_8647,N_4874,N_5282);
and U8648 (N_8648,N_3538,N_3572);
nand U8649 (N_8649,N_4386,N_3726);
or U8650 (N_8650,N_5853,N_3766);
and U8651 (N_8651,N_5008,N_3941);
nand U8652 (N_8652,N_5477,N_5491);
nand U8653 (N_8653,N_4063,N_5637);
nand U8654 (N_8654,N_3829,N_5323);
nor U8655 (N_8655,N_4370,N_3844);
nor U8656 (N_8656,N_5496,N_4187);
xor U8657 (N_8657,N_4451,N_3934);
nand U8658 (N_8658,N_5239,N_4524);
and U8659 (N_8659,N_4791,N_5922);
or U8660 (N_8660,N_5675,N_4274);
and U8661 (N_8661,N_4667,N_4933);
or U8662 (N_8662,N_3731,N_4650);
and U8663 (N_8663,N_4546,N_5280);
xor U8664 (N_8664,N_5368,N_5624);
or U8665 (N_8665,N_5952,N_4168);
nor U8666 (N_8666,N_3254,N_4293);
nand U8667 (N_8667,N_4968,N_3426);
or U8668 (N_8668,N_4156,N_3581);
nor U8669 (N_8669,N_3409,N_5539);
nor U8670 (N_8670,N_3838,N_4049);
nor U8671 (N_8671,N_4857,N_4582);
xor U8672 (N_8672,N_3136,N_3504);
xnor U8673 (N_8673,N_3240,N_5404);
nor U8674 (N_8674,N_5812,N_6089);
and U8675 (N_8675,N_4611,N_4923);
or U8676 (N_8676,N_3128,N_5227);
nand U8677 (N_8677,N_6237,N_4131);
and U8678 (N_8678,N_5552,N_4712);
or U8679 (N_8679,N_4315,N_4043);
xnor U8680 (N_8680,N_5098,N_4388);
nor U8681 (N_8681,N_5931,N_4528);
or U8682 (N_8682,N_5910,N_4679);
nor U8683 (N_8683,N_4253,N_5302);
nand U8684 (N_8684,N_3128,N_5564);
nand U8685 (N_8685,N_4593,N_5846);
xnor U8686 (N_8686,N_4989,N_5693);
or U8687 (N_8687,N_5727,N_5508);
or U8688 (N_8688,N_5912,N_4808);
nor U8689 (N_8689,N_6115,N_6064);
xor U8690 (N_8690,N_6217,N_3377);
and U8691 (N_8691,N_3835,N_6072);
or U8692 (N_8692,N_3812,N_6128);
xnor U8693 (N_8693,N_3998,N_3803);
or U8694 (N_8694,N_5984,N_4489);
nand U8695 (N_8695,N_5441,N_4880);
or U8696 (N_8696,N_3837,N_3944);
and U8697 (N_8697,N_4073,N_5868);
nand U8698 (N_8698,N_6006,N_5300);
and U8699 (N_8699,N_5825,N_4526);
and U8700 (N_8700,N_4471,N_5693);
nand U8701 (N_8701,N_4636,N_3558);
nor U8702 (N_8702,N_5696,N_3353);
or U8703 (N_8703,N_5377,N_4987);
or U8704 (N_8704,N_5175,N_4675);
nand U8705 (N_8705,N_4657,N_3153);
nand U8706 (N_8706,N_4901,N_6108);
xnor U8707 (N_8707,N_5172,N_5689);
nand U8708 (N_8708,N_3931,N_3824);
and U8709 (N_8709,N_3526,N_5838);
xor U8710 (N_8710,N_4653,N_4282);
and U8711 (N_8711,N_4349,N_3695);
or U8712 (N_8712,N_4153,N_5886);
and U8713 (N_8713,N_4764,N_6084);
and U8714 (N_8714,N_5176,N_4074);
and U8715 (N_8715,N_3343,N_5865);
and U8716 (N_8716,N_4032,N_3476);
or U8717 (N_8717,N_3754,N_4464);
nand U8718 (N_8718,N_5333,N_3893);
or U8719 (N_8719,N_4301,N_5816);
xor U8720 (N_8720,N_5822,N_5277);
nand U8721 (N_8721,N_4305,N_4468);
nand U8722 (N_8722,N_5471,N_5700);
nor U8723 (N_8723,N_3913,N_4322);
xnor U8724 (N_8724,N_3684,N_5693);
xor U8725 (N_8725,N_5071,N_4704);
and U8726 (N_8726,N_3722,N_3459);
or U8727 (N_8727,N_3272,N_4198);
xnor U8728 (N_8728,N_4406,N_5522);
xnor U8729 (N_8729,N_4802,N_5316);
and U8730 (N_8730,N_6038,N_3400);
nand U8731 (N_8731,N_6038,N_5244);
nand U8732 (N_8732,N_3910,N_3591);
nand U8733 (N_8733,N_3920,N_3911);
and U8734 (N_8734,N_6192,N_3336);
nand U8735 (N_8735,N_3380,N_3391);
xnor U8736 (N_8736,N_6086,N_5833);
xor U8737 (N_8737,N_5966,N_5284);
nor U8738 (N_8738,N_4831,N_4092);
xor U8739 (N_8739,N_4585,N_5557);
nor U8740 (N_8740,N_5927,N_4280);
and U8741 (N_8741,N_4728,N_4117);
or U8742 (N_8742,N_3245,N_4702);
or U8743 (N_8743,N_5460,N_5513);
or U8744 (N_8744,N_4702,N_5334);
and U8745 (N_8745,N_4419,N_5216);
xnor U8746 (N_8746,N_3920,N_3924);
nand U8747 (N_8747,N_3862,N_5451);
or U8748 (N_8748,N_5691,N_6095);
and U8749 (N_8749,N_4517,N_4810);
or U8750 (N_8750,N_5465,N_4467);
nor U8751 (N_8751,N_5195,N_4138);
or U8752 (N_8752,N_4948,N_3404);
nor U8753 (N_8753,N_3970,N_4659);
or U8754 (N_8754,N_3617,N_4696);
nor U8755 (N_8755,N_3991,N_4704);
nor U8756 (N_8756,N_3179,N_5073);
nor U8757 (N_8757,N_3629,N_6034);
nor U8758 (N_8758,N_4688,N_5557);
or U8759 (N_8759,N_5863,N_5306);
xnor U8760 (N_8760,N_4273,N_3419);
xor U8761 (N_8761,N_3175,N_4968);
nor U8762 (N_8762,N_5998,N_6180);
or U8763 (N_8763,N_5960,N_4886);
and U8764 (N_8764,N_4886,N_5131);
nor U8765 (N_8765,N_5558,N_4162);
xor U8766 (N_8766,N_3831,N_4927);
nand U8767 (N_8767,N_5518,N_6206);
and U8768 (N_8768,N_5212,N_4692);
nand U8769 (N_8769,N_5389,N_5919);
and U8770 (N_8770,N_3807,N_5282);
or U8771 (N_8771,N_5575,N_3373);
nor U8772 (N_8772,N_3264,N_5389);
nand U8773 (N_8773,N_4971,N_4686);
or U8774 (N_8774,N_3769,N_4479);
and U8775 (N_8775,N_4735,N_5401);
nand U8776 (N_8776,N_5609,N_4172);
or U8777 (N_8777,N_5333,N_3173);
xnor U8778 (N_8778,N_6071,N_5150);
xor U8779 (N_8779,N_5966,N_5277);
nand U8780 (N_8780,N_3711,N_4558);
and U8781 (N_8781,N_4712,N_5212);
xnor U8782 (N_8782,N_4100,N_5580);
nor U8783 (N_8783,N_5333,N_5307);
xor U8784 (N_8784,N_4097,N_6130);
or U8785 (N_8785,N_5015,N_4045);
xnor U8786 (N_8786,N_5794,N_5051);
and U8787 (N_8787,N_3772,N_5826);
nor U8788 (N_8788,N_4490,N_3243);
nand U8789 (N_8789,N_5658,N_3364);
or U8790 (N_8790,N_5453,N_6176);
or U8791 (N_8791,N_5629,N_3240);
xor U8792 (N_8792,N_3930,N_4051);
and U8793 (N_8793,N_5918,N_6088);
nand U8794 (N_8794,N_3251,N_4246);
nand U8795 (N_8795,N_3560,N_4312);
nor U8796 (N_8796,N_4679,N_3544);
nor U8797 (N_8797,N_5736,N_3657);
nand U8798 (N_8798,N_5263,N_6115);
and U8799 (N_8799,N_5307,N_3613);
or U8800 (N_8800,N_6188,N_4215);
and U8801 (N_8801,N_6021,N_5757);
nand U8802 (N_8802,N_5592,N_5260);
nand U8803 (N_8803,N_4454,N_4491);
nand U8804 (N_8804,N_4903,N_5343);
or U8805 (N_8805,N_3633,N_5292);
or U8806 (N_8806,N_4473,N_4674);
and U8807 (N_8807,N_3259,N_3548);
xnor U8808 (N_8808,N_3994,N_5909);
or U8809 (N_8809,N_3273,N_5790);
xor U8810 (N_8810,N_6039,N_3994);
nand U8811 (N_8811,N_5797,N_4990);
xnor U8812 (N_8812,N_5853,N_3581);
and U8813 (N_8813,N_5102,N_5503);
xnor U8814 (N_8814,N_4542,N_4633);
xor U8815 (N_8815,N_6032,N_4598);
nor U8816 (N_8816,N_4702,N_4027);
nand U8817 (N_8817,N_4113,N_4263);
nand U8818 (N_8818,N_3909,N_4185);
or U8819 (N_8819,N_4192,N_5697);
nand U8820 (N_8820,N_5760,N_6232);
or U8821 (N_8821,N_4294,N_4633);
xnor U8822 (N_8822,N_3381,N_5218);
and U8823 (N_8823,N_5951,N_3928);
or U8824 (N_8824,N_5985,N_3788);
and U8825 (N_8825,N_5555,N_3333);
or U8826 (N_8826,N_5695,N_4542);
and U8827 (N_8827,N_4918,N_5513);
xnor U8828 (N_8828,N_6188,N_4976);
nand U8829 (N_8829,N_3129,N_3333);
nor U8830 (N_8830,N_4683,N_5456);
nor U8831 (N_8831,N_4321,N_4162);
and U8832 (N_8832,N_5317,N_4904);
or U8833 (N_8833,N_4532,N_3502);
and U8834 (N_8834,N_3375,N_5343);
nand U8835 (N_8835,N_4783,N_3568);
nand U8836 (N_8836,N_4345,N_3302);
xnor U8837 (N_8837,N_5582,N_5166);
and U8838 (N_8838,N_5022,N_3770);
nand U8839 (N_8839,N_3232,N_4056);
and U8840 (N_8840,N_3330,N_6196);
xnor U8841 (N_8841,N_4679,N_4673);
and U8842 (N_8842,N_4357,N_5231);
and U8843 (N_8843,N_5983,N_5907);
xnor U8844 (N_8844,N_4891,N_3277);
xor U8845 (N_8845,N_5180,N_4327);
and U8846 (N_8846,N_4499,N_5086);
nand U8847 (N_8847,N_4757,N_4227);
and U8848 (N_8848,N_5513,N_4944);
xnor U8849 (N_8849,N_4644,N_5764);
and U8850 (N_8850,N_3148,N_3230);
xor U8851 (N_8851,N_6116,N_5926);
or U8852 (N_8852,N_4068,N_3166);
nand U8853 (N_8853,N_5709,N_3583);
xor U8854 (N_8854,N_4465,N_4048);
nand U8855 (N_8855,N_6097,N_3355);
xnor U8856 (N_8856,N_4727,N_4958);
nand U8857 (N_8857,N_4230,N_4068);
nor U8858 (N_8858,N_6111,N_5288);
and U8859 (N_8859,N_6097,N_5246);
nand U8860 (N_8860,N_5167,N_3834);
xor U8861 (N_8861,N_4253,N_4476);
or U8862 (N_8862,N_5346,N_5786);
xor U8863 (N_8863,N_3882,N_6074);
and U8864 (N_8864,N_4224,N_3509);
nor U8865 (N_8865,N_4021,N_4049);
or U8866 (N_8866,N_3514,N_4078);
or U8867 (N_8867,N_6033,N_4876);
xor U8868 (N_8868,N_4687,N_4534);
or U8869 (N_8869,N_5805,N_6060);
and U8870 (N_8870,N_4568,N_6010);
nor U8871 (N_8871,N_5752,N_6043);
or U8872 (N_8872,N_3761,N_3708);
or U8873 (N_8873,N_3294,N_3298);
nand U8874 (N_8874,N_5750,N_4489);
nand U8875 (N_8875,N_6240,N_4659);
xnor U8876 (N_8876,N_6193,N_3485);
and U8877 (N_8877,N_6001,N_5242);
nand U8878 (N_8878,N_3343,N_3560);
nor U8879 (N_8879,N_3464,N_5901);
nand U8880 (N_8880,N_5867,N_6142);
nand U8881 (N_8881,N_5088,N_4556);
and U8882 (N_8882,N_5688,N_5112);
xnor U8883 (N_8883,N_3681,N_4504);
nor U8884 (N_8884,N_6063,N_3186);
nand U8885 (N_8885,N_5376,N_3703);
and U8886 (N_8886,N_5750,N_4575);
and U8887 (N_8887,N_3785,N_4198);
nand U8888 (N_8888,N_4803,N_3146);
and U8889 (N_8889,N_5315,N_4129);
nor U8890 (N_8890,N_5188,N_3988);
nand U8891 (N_8891,N_5416,N_3632);
xor U8892 (N_8892,N_5566,N_5956);
or U8893 (N_8893,N_5047,N_4971);
or U8894 (N_8894,N_4209,N_5446);
and U8895 (N_8895,N_4900,N_4916);
and U8896 (N_8896,N_4456,N_3167);
or U8897 (N_8897,N_4156,N_5787);
or U8898 (N_8898,N_3775,N_3474);
nand U8899 (N_8899,N_5477,N_4738);
and U8900 (N_8900,N_5946,N_3614);
nand U8901 (N_8901,N_4495,N_6137);
nand U8902 (N_8902,N_3493,N_4298);
nand U8903 (N_8903,N_3251,N_4258);
xor U8904 (N_8904,N_5074,N_5889);
and U8905 (N_8905,N_3166,N_4165);
nand U8906 (N_8906,N_5243,N_5536);
nor U8907 (N_8907,N_4065,N_5364);
nand U8908 (N_8908,N_5637,N_4030);
xor U8909 (N_8909,N_3329,N_4192);
nor U8910 (N_8910,N_3504,N_4795);
or U8911 (N_8911,N_5097,N_4853);
or U8912 (N_8912,N_3801,N_3644);
or U8913 (N_8913,N_5635,N_5877);
and U8914 (N_8914,N_5987,N_5364);
and U8915 (N_8915,N_3376,N_4693);
or U8916 (N_8916,N_5128,N_4626);
nor U8917 (N_8917,N_4869,N_4991);
or U8918 (N_8918,N_5011,N_3340);
nor U8919 (N_8919,N_5123,N_5970);
xor U8920 (N_8920,N_4199,N_5973);
and U8921 (N_8921,N_5760,N_5039);
or U8922 (N_8922,N_5112,N_4742);
and U8923 (N_8923,N_5467,N_5985);
nor U8924 (N_8924,N_5722,N_3172);
and U8925 (N_8925,N_4330,N_4612);
xnor U8926 (N_8926,N_5070,N_3173);
nor U8927 (N_8927,N_5919,N_4296);
or U8928 (N_8928,N_3183,N_4963);
nor U8929 (N_8929,N_5037,N_3499);
nand U8930 (N_8930,N_4520,N_3950);
and U8931 (N_8931,N_5958,N_5977);
nand U8932 (N_8932,N_4921,N_4971);
xor U8933 (N_8933,N_3978,N_4167);
or U8934 (N_8934,N_4631,N_3230);
nand U8935 (N_8935,N_5194,N_3542);
xnor U8936 (N_8936,N_5809,N_6244);
and U8937 (N_8937,N_3715,N_5575);
nor U8938 (N_8938,N_3546,N_4919);
or U8939 (N_8939,N_5886,N_4726);
nand U8940 (N_8940,N_3753,N_5040);
xnor U8941 (N_8941,N_4688,N_3455);
and U8942 (N_8942,N_5022,N_4490);
and U8943 (N_8943,N_4329,N_5929);
and U8944 (N_8944,N_4414,N_3256);
or U8945 (N_8945,N_3375,N_5192);
nor U8946 (N_8946,N_4362,N_5529);
or U8947 (N_8947,N_4186,N_3938);
and U8948 (N_8948,N_4250,N_4803);
or U8949 (N_8949,N_6156,N_4291);
xnor U8950 (N_8950,N_3170,N_3448);
xnor U8951 (N_8951,N_4015,N_3635);
nor U8952 (N_8952,N_4237,N_5739);
nand U8953 (N_8953,N_5029,N_4391);
xor U8954 (N_8954,N_5363,N_5689);
or U8955 (N_8955,N_4021,N_3161);
nor U8956 (N_8956,N_6248,N_4690);
and U8957 (N_8957,N_3484,N_5264);
xnor U8958 (N_8958,N_4167,N_4508);
xor U8959 (N_8959,N_5245,N_5866);
nor U8960 (N_8960,N_4586,N_4924);
and U8961 (N_8961,N_3140,N_5190);
nand U8962 (N_8962,N_4405,N_3657);
and U8963 (N_8963,N_3489,N_3663);
nor U8964 (N_8964,N_5127,N_4000);
and U8965 (N_8965,N_5568,N_4514);
xor U8966 (N_8966,N_3287,N_3328);
nand U8967 (N_8967,N_6134,N_3262);
nand U8968 (N_8968,N_5035,N_4660);
xnor U8969 (N_8969,N_6168,N_5267);
nor U8970 (N_8970,N_5211,N_3381);
and U8971 (N_8971,N_3862,N_4348);
and U8972 (N_8972,N_3864,N_4599);
nand U8973 (N_8973,N_4730,N_5209);
xnor U8974 (N_8974,N_5959,N_5867);
and U8975 (N_8975,N_4917,N_6112);
or U8976 (N_8976,N_4403,N_5964);
xor U8977 (N_8977,N_3668,N_3836);
xnor U8978 (N_8978,N_3470,N_5455);
or U8979 (N_8979,N_5992,N_4330);
nor U8980 (N_8980,N_3260,N_4194);
or U8981 (N_8981,N_3955,N_5492);
or U8982 (N_8982,N_3625,N_5348);
and U8983 (N_8983,N_5976,N_5482);
and U8984 (N_8984,N_3656,N_6038);
nand U8985 (N_8985,N_3208,N_4575);
or U8986 (N_8986,N_3919,N_4219);
or U8987 (N_8987,N_5654,N_3955);
or U8988 (N_8988,N_3223,N_5112);
or U8989 (N_8989,N_4424,N_5721);
nand U8990 (N_8990,N_5797,N_5330);
or U8991 (N_8991,N_4608,N_5959);
xnor U8992 (N_8992,N_3717,N_5781);
nand U8993 (N_8993,N_4321,N_4972);
and U8994 (N_8994,N_4697,N_4764);
and U8995 (N_8995,N_5915,N_5897);
and U8996 (N_8996,N_4406,N_3506);
or U8997 (N_8997,N_3677,N_4972);
and U8998 (N_8998,N_4717,N_5910);
or U8999 (N_8999,N_4104,N_5292);
xnor U9000 (N_9000,N_4502,N_3608);
or U9001 (N_9001,N_5684,N_4067);
and U9002 (N_9002,N_5879,N_5846);
nand U9003 (N_9003,N_4377,N_3130);
or U9004 (N_9004,N_5639,N_4567);
xnor U9005 (N_9005,N_4830,N_4183);
xor U9006 (N_9006,N_5204,N_4739);
or U9007 (N_9007,N_4946,N_4649);
and U9008 (N_9008,N_4669,N_4389);
xnor U9009 (N_9009,N_6087,N_5848);
or U9010 (N_9010,N_4786,N_4449);
or U9011 (N_9011,N_3685,N_5540);
nor U9012 (N_9012,N_5524,N_6119);
nor U9013 (N_9013,N_4765,N_3306);
nand U9014 (N_9014,N_5479,N_4232);
or U9015 (N_9015,N_6092,N_5589);
and U9016 (N_9016,N_4766,N_5813);
nand U9017 (N_9017,N_3218,N_5976);
and U9018 (N_9018,N_5522,N_4285);
xor U9019 (N_9019,N_4299,N_3775);
or U9020 (N_9020,N_5634,N_5352);
xnor U9021 (N_9021,N_6235,N_5784);
and U9022 (N_9022,N_3886,N_5086);
xnor U9023 (N_9023,N_4421,N_4298);
and U9024 (N_9024,N_3283,N_6059);
xor U9025 (N_9025,N_3479,N_5055);
xor U9026 (N_9026,N_5716,N_5856);
xor U9027 (N_9027,N_4772,N_3720);
nor U9028 (N_9028,N_5543,N_4561);
nor U9029 (N_9029,N_5996,N_5786);
and U9030 (N_9030,N_4880,N_6121);
or U9031 (N_9031,N_4919,N_5313);
nand U9032 (N_9032,N_4097,N_5172);
or U9033 (N_9033,N_3331,N_5486);
or U9034 (N_9034,N_3211,N_3584);
nand U9035 (N_9035,N_5818,N_4007);
nor U9036 (N_9036,N_4201,N_5697);
and U9037 (N_9037,N_5331,N_5777);
xor U9038 (N_9038,N_5997,N_4743);
nand U9039 (N_9039,N_3778,N_3199);
and U9040 (N_9040,N_4435,N_5337);
xnor U9041 (N_9041,N_6050,N_5842);
nor U9042 (N_9042,N_4854,N_5539);
and U9043 (N_9043,N_3734,N_5579);
nor U9044 (N_9044,N_5596,N_3154);
xnor U9045 (N_9045,N_6139,N_5276);
nor U9046 (N_9046,N_4413,N_4769);
xnor U9047 (N_9047,N_3509,N_5502);
nand U9048 (N_9048,N_5182,N_5172);
nor U9049 (N_9049,N_6023,N_4823);
and U9050 (N_9050,N_5146,N_3401);
xor U9051 (N_9051,N_5307,N_3668);
xor U9052 (N_9052,N_5027,N_3408);
nor U9053 (N_9053,N_3816,N_6018);
nand U9054 (N_9054,N_4876,N_3557);
or U9055 (N_9055,N_5768,N_5325);
xor U9056 (N_9056,N_4963,N_3512);
nor U9057 (N_9057,N_4806,N_5886);
or U9058 (N_9058,N_4378,N_3436);
nor U9059 (N_9059,N_3685,N_4778);
nand U9060 (N_9060,N_5660,N_5759);
nand U9061 (N_9061,N_3846,N_3490);
nand U9062 (N_9062,N_4506,N_3467);
nor U9063 (N_9063,N_3173,N_5668);
nand U9064 (N_9064,N_3265,N_5551);
or U9065 (N_9065,N_4085,N_3919);
or U9066 (N_9066,N_4201,N_5349);
or U9067 (N_9067,N_3833,N_3238);
xnor U9068 (N_9068,N_3724,N_5816);
and U9069 (N_9069,N_3608,N_3681);
nand U9070 (N_9070,N_6074,N_4006);
xnor U9071 (N_9071,N_3888,N_4245);
and U9072 (N_9072,N_5535,N_5341);
or U9073 (N_9073,N_3944,N_5236);
nor U9074 (N_9074,N_3699,N_5303);
or U9075 (N_9075,N_5221,N_4116);
nand U9076 (N_9076,N_3994,N_4299);
nor U9077 (N_9077,N_3504,N_5747);
and U9078 (N_9078,N_4057,N_5263);
xnor U9079 (N_9079,N_6234,N_4293);
nand U9080 (N_9080,N_4726,N_5668);
nand U9081 (N_9081,N_5860,N_4393);
nor U9082 (N_9082,N_6174,N_3850);
or U9083 (N_9083,N_5630,N_4330);
or U9084 (N_9084,N_4766,N_3173);
nand U9085 (N_9085,N_4530,N_3754);
nor U9086 (N_9086,N_4025,N_5850);
nor U9087 (N_9087,N_6154,N_5186);
nand U9088 (N_9088,N_3201,N_3284);
nand U9089 (N_9089,N_6247,N_4015);
nor U9090 (N_9090,N_5358,N_4041);
xor U9091 (N_9091,N_5318,N_5325);
or U9092 (N_9092,N_5586,N_5402);
or U9093 (N_9093,N_4373,N_5208);
nor U9094 (N_9094,N_6016,N_3938);
nand U9095 (N_9095,N_5377,N_5633);
nand U9096 (N_9096,N_4463,N_4109);
and U9097 (N_9097,N_5001,N_5396);
and U9098 (N_9098,N_5963,N_5481);
and U9099 (N_9099,N_6172,N_3422);
nor U9100 (N_9100,N_4887,N_3620);
and U9101 (N_9101,N_3806,N_5638);
or U9102 (N_9102,N_5890,N_5616);
nor U9103 (N_9103,N_5453,N_3309);
nand U9104 (N_9104,N_6180,N_3646);
nor U9105 (N_9105,N_4089,N_4644);
or U9106 (N_9106,N_3836,N_5635);
xnor U9107 (N_9107,N_3325,N_3962);
xor U9108 (N_9108,N_4767,N_3920);
nand U9109 (N_9109,N_5448,N_5544);
xor U9110 (N_9110,N_4145,N_3769);
nand U9111 (N_9111,N_5204,N_3847);
nand U9112 (N_9112,N_6050,N_5745);
nand U9113 (N_9113,N_6083,N_6216);
xnor U9114 (N_9114,N_5949,N_4646);
nor U9115 (N_9115,N_5728,N_4169);
nor U9116 (N_9116,N_4466,N_4244);
or U9117 (N_9117,N_4061,N_3876);
or U9118 (N_9118,N_5908,N_5252);
nand U9119 (N_9119,N_4967,N_5966);
nor U9120 (N_9120,N_5493,N_4372);
and U9121 (N_9121,N_3891,N_6240);
nor U9122 (N_9122,N_3716,N_5866);
and U9123 (N_9123,N_6049,N_5516);
nand U9124 (N_9124,N_4512,N_5591);
nand U9125 (N_9125,N_5598,N_3370);
xnor U9126 (N_9126,N_4087,N_3731);
nor U9127 (N_9127,N_6156,N_3709);
or U9128 (N_9128,N_3553,N_3982);
and U9129 (N_9129,N_3669,N_3445);
nor U9130 (N_9130,N_4373,N_5947);
nand U9131 (N_9131,N_5424,N_3802);
xor U9132 (N_9132,N_4765,N_4398);
and U9133 (N_9133,N_3742,N_5533);
and U9134 (N_9134,N_4296,N_4241);
or U9135 (N_9135,N_5773,N_4026);
nor U9136 (N_9136,N_4077,N_4824);
and U9137 (N_9137,N_3432,N_5555);
or U9138 (N_9138,N_4337,N_6245);
xor U9139 (N_9139,N_5997,N_5017);
or U9140 (N_9140,N_3669,N_5840);
nor U9141 (N_9141,N_5565,N_5470);
nor U9142 (N_9142,N_4450,N_4764);
and U9143 (N_9143,N_4339,N_6018);
nand U9144 (N_9144,N_4988,N_4694);
or U9145 (N_9145,N_5370,N_5420);
or U9146 (N_9146,N_3503,N_5407);
and U9147 (N_9147,N_5318,N_6239);
nor U9148 (N_9148,N_5923,N_3370);
or U9149 (N_9149,N_3434,N_4554);
nand U9150 (N_9150,N_5808,N_4131);
nor U9151 (N_9151,N_5656,N_6170);
xnor U9152 (N_9152,N_5080,N_3397);
nor U9153 (N_9153,N_6200,N_4622);
and U9154 (N_9154,N_6170,N_4362);
and U9155 (N_9155,N_3203,N_5995);
nand U9156 (N_9156,N_5790,N_6040);
nor U9157 (N_9157,N_3658,N_3464);
nor U9158 (N_9158,N_5883,N_5209);
and U9159 (N_9159,N_4446,N_4008);
nor U9160 (N_9160,N_4923,N_5549);
or U9161 (N_9161,N_4736,N_4467);
nand U9162 (N_9162,N_5918,N_3574);
and U9163 (N_9163,N_5615,N_4191);
or U9164 (N_9164,N_3692,N_3630);
and U9165 (N_9165,N_4836,N_5017);
xor U9166 (N_9166,N_3211,N_5940);
or U9167 (N_9167,N_5910,N_4751);
nor U9168 (N_9168,N_3566,N_5721);
xor U9169 (N_9169,N_3489,N_3386);
and U9170 (N_9170,N_3196,N_5208);
nor U9171 (N_9171,N_4689,N_5687);
or U9172 (N_9172,N_3655,N_4066);
nand U9173 (N_9173,N_5747,N_6006);
and U9174 (N_9174,N_4559,N_3391);
and U9175 (N_9175,N_6061,N_5528);
nand U9176 (N_9176,N_5813,N_6231);
and U9177 (N_9177,N_4663,N_5680);
xor U9178 (N_9178,N_3470,N_4806);
and U9179 (N_9179,N_3667,N_3938);
and U9180 (N_9180,N_6153,N_5277);
nor U9181 (N_9181,N_5245,N_4798);
or U9182 (N_9182,N_5894,N_5727);
nor U9183 (N_9183,N_5558,N_3626);
nand U9184 (N_9184,N_5446,N_6186);
xor U9185 (N_9185,N_3999,N_5640);
nor U9186 (N_9186,N_4137,N_3395);
or U9187 (N_9187,N_6100,N_5402);
nand U9188 (N_9188,N_4051,N_3324);
nor U9189 (N_9189,N_3322,N_5500);
and U9190 (N_9190,N_3941,N_5546);
nand U9191 (N_9191,N_5857,N_4504);
xnor U9192 (N_9192,N_3340,N_4739);
nor U9193 (N_9193,N_4862,N_3399);
nand U9194 (N_9194,N_5146,N_4950);
xnor U9195 (N_9195,N_4450,N_4479);
nand U9196 (N_9196,N_4312,N_3709);
nor U9197 (N_9197,N_3346,N_4808);
nor U9198 (N_9198,N_5796,N_3347);
xor U9199 (N_9199,N_4117,N_3382);
nor U9200 (N_9200,N_5910,N_5711);
or U9201 (N_9201,N_4786,N_6148);
and U9202 (N_9202,N_5952,N_4589);
or U9203 (N_9203,N_5943,N_4771);
and U9204 (N_9204,N_3356,N_3640);
nor U9205 (N_9205,N_5566,N_3445);
nand U9206 (N_9206,N_5433,N_5639);
nor U9207 (N_9207,N_3307,N_5186);
and U9208 (N_9208,N_4245,N_3538);
or U9209 (N_9209,N_5098,N_5257);
or U9210 (N_9210,N_3460,N_4163);
nor U9211 (N_9211,N_4007,N_6034);
and U9212 (N_9212,N_4107,N_5864);
nand U9213 (N_9213,N_3196,N_3526);
or U9214 (N_9214,N_5302,N_4040);
nor U9215 (N_9215,N_4663,N_4202);
xnor U9216 (N_9216,N_3833,N_6195);
or U9217 (N_9217,N_5515,N_6051);
and U9218 (N_9218,N_5300,N_4175);
nand U9219 (N_9219,N_6170,N_4701);
nand U9220 (N_9220,N_3825,N_5254);
nor U9221 (N_9221,N_4209,N_4548);
nand U9222 (N_9222,N_3373,N_3512);
nand U9223 (N_9223,N_6061,N_3585);
or U9224 (N_9224,N_5644,N_5415);
and U9225 (N_9225,N_5626,N_6125);
and U9226 (N_9226,N_3968,N_4335);
and U9227 (N_9227,N_4514,N_5354);
and U9228 (N_9228,N_5250,N_3316);
nand U9229 (N_9229,N_4905,N_3465);
xor U9230 (N_9230,N_4299,N_5521);
xnor U9231 (N_9231,N_4056,N_6033);
or U9232 (N_9232,N_4976,N_5927);
or U9233 (N_9233,N_4253,N_4656);
xnor U9234 (N_9234,N_5494,N_5563);
nand U9235 (N_9235,N_4292,N_6053);
and U9236 (N_9236,N_5629,N_4004);
and U9237 (N_9237,N_4491,N_3160);
and U9238 (N_9238,N_3378,N_5736);
nor U9239 (N_9239,N_5651,N_5977);
nor U9240 (N_9240,N_5968,N_6247);
xnor U9241 (N_9241,N_3814,N_5676);
nor U9242 (N_9242,N_3369,N_3299);
nand U9243 (N_9243,N_5573,N_5268);
nor U9244 (N_9244,N_4478,N_3801);
nor U9245 (N_9245,N_4903,N_4886);
and U9246 (N_9246,N_5333,N_4920);
and U9247 (N_9247,N_4131,N_3455);
and U9248 (N_9248,N_5310,N_4433);
and U9249 (N_9249,N_5623,N_4837);
nor U9250 (N_9250,N_5196,N_5975);
nand U9251 (N_9251,N_4737,N_3968);
nand U9252 (N_9252,N_3521,N_4010);
or U9253 (N_9253,N_3788,N_3274);
and U9254 (N_9254,N_4145,N_5217);
or U9255 (N_9255,N_3609,N_3133);
and U9256 (N_9256,N_5247,N_4180);
xnor U9257 (N_9257,N_3275,N_5033);
nor U9258 (N_9258,N_3381,N_5606);
and U9259 (N_9259,N_4608,N_3512);
and U9260 (N_9260,N_4057,N_4449);
and U9261 (N_9261,N_4219,N_4936);
and U9262 (N_9262,N_5552,N_3392);
xnor U9263 (N_9263,N_5753,N_3269);
or U9264 (N_9264,N_5257,N_4069);
or U9265 (N_9265,N_4428,N_3801);
xnor U9266 (N_9266,N_4813,N_4691);
or U9267 (N_9267,N_4018,N_5948);
or U9268 (N_9268,N_3723,N_3125);
and U9269 (N_9269,N_6046,N_3789);
nand U9270 (N_9270,N_3950,N_3704);
nor U9271 (N_9271,N_5402,N_3224);
nor U9272 (N_9272,N_3844,N_5498);
or U9273 (N_9273,N_4828,N_3155);
and U9274 (N_9274,N_6188,N_4836);
or U9275 (N_9275,N_5983,N_4157);
or U9276 (N_9276,N_3225,N_5625);
nor U9277 (N_9277,N_5111,N_5808);
or U9278 (N_9278,N_5043,N_6035);
nor U9279 (N_9279,N_5732,N_6191);
xor U9280 (N_9280,N_5167,N_3912);
or U9281 (N_9281,N_3919,N_5432);
nor U9282 (N_9282,N_4407,N_4493);
nor U9283 (N_9283,N_4114,N_3356);
nand U9284 (N_9284,N_3542,N_6105);
nor U9285 (N_9285,N_4032,N_3274);
nand U9286 (N_9286,N_3992,N_5793);
nor U9287 (N_9287,N_3711,N_5369);
nand U9288 (N_9288,N_3795,N_4295);
xor U9289 (N_9289,N_5137,N_6127);
xnor U9290 (N_9290,N_5629,N_4814);
and U9291 (N_9291,N_3698,N_3450);
nand U9292 (N_9292,N_5310,N_6084);
or U9293 (N_9293,N_3658,N_3365);
nor U9294 (N_9294,N_4541,N_6040);
and U9295 (N_9295,N_5743,N_5241);
or U9296 (N_9296,N_4867,N_3542);
or U9297 (N_9297,N_3513,N_3855);
or U9298 (N_9298,N_5620,N_3193);
and U9299 (N_9299,N_5065,N_3343);
xor U9300 (N_9300,N_6025,N_3305);
and U9301 (N_9301,N_5416,N_3313);
and U9302 (N_9302,N_5562,N_3399);
or U9303 (N_9303,N_5632,N_3944);
xnor U9304 (N_9304,N_4467,N_6058);
xnor U9305 (N_9305,N_6066,N_4432);
nor U9306 (N_9306,N_3146,N_5882);
nand U9307 (N_9307,N_3776,N_4734);
and U9308 (N_9308,N_5652,N_5824);
xnor U9309 (N_9309,N_3793,N_3489);
or U9310 (N_9310,N_6145,N_3682);
or U9311 (N_9311,N_4044,N_3644);
nand U9312 (N_9312,N_3293,N_3719);
nand U9313 (N_9313,N_3987,N_5583);
nor U9314 (N_9314,N_5346,N_6225);
and U9315 (N_9315,N_4361,N_4619);
xnor U9316 (N_9316,N_5902,N_3455);
or U9317 (N_9317,N_4541,N_4772);
nand U9318 (N_9318,N_4930,N_5941);
or U9319 (N_9319,N_3254,N_5774);
and U9320 (N_9320,N_5310,N_4764);
xnor U9321 (N_9321,N_3712,N_6172);
nor U9322 (N_9322,N_4587,N_3280);
nor U9323 (N_9323,N_5326,N_3691);
nand U9324 (N_9324,N_3444,N_4670);
xnor U9325 (N_9325,N_3542,N_3619);
nand U9326 (N_9326,N_3503,N_3505);
and U9327 (N_9327,N_5763,N_4049);
xnor U9328 (N_9328,N_3443,N_4373);
and U9329 (N_9329,N_3136,N_5668);
xnor U9330 (N_9330,N_6025,N_4870);
and U9331 (N_9331,N_5540,N_3481);
or U9332 (N_9332,N_5842,N_5837);
xnor U9333 (N_9333,N_5266,N_3963);
and U9334 (N_9334,N_4254,N_6211);
nand U9335 (N_9335,N_4603,N_4221);
or U9336 (N_9336,N_4908,N_6069);
or U9337 (N_9337,N_3787,N_5884);
nor U9338 (N_9338,N_3152,N_5789);
xnor U9339 (N_9339,N_5309,N_3529);
nor U9340 (N_9340,N_3218,N_5204);
xor U9341 (N_9341,N_6123,N_3368);
nand U9342 (N_9342,N_3883,N_5951);
or U9343 (N_9343,N_5810,N_5327);
xor U9344 (N_9344,N_3869,N_4997);
nor U9345 (N_9345,N_5609,N_4522);
nand U9346 (N_9346,N_4230,N_3422);
nand U9347 (N_9347,N_3471,N_3996);
xor U9348 (N_9348,N_3319,N_6197);
xnor U9349 (N_9349,N_6065,N_5044);
nor U9350 (N_9350,N_4293,N_4820);
nand U9351 (N_9351,N_5108,N_5395);
xor U9352 (N_9352,N_3148,N_5065);
and U9353 (N_9353,N_3484,N_3662);
or U9354 (N_9354,N_4817,N_5769);
nor U9355 (N_9355,N_4316,N_5809);
and U9356 (N_9356,N_5224,N_5456);
and U9357 (N_9357,N_3291,N_6085);
xor U9358 (N_9358,N_5916,N_3843);
and U9359 (N_9359,N_4217,N_4104);
and U9360 (N_9360,N_5971,N_6158);
xnor U9361 (N_9361,N_4387,N_5218);
and U9362 (N_9362,N_4155,N_4684);
xor U9363 (N_9363,N_3352,N_4478);
or U9364 (N_9364,N_5539,N_4459);
and U9365 (N_9365,N_4119,N_6183);
or U9366 (N_9366,N_4768,N_5986);
nand U9367 (N_9367,N_5766,N_4752);
nor U9368 (N_9368,N_4650,N_5478);
or U9369 (N_9369,N_4479,N_4567);
nand U9370 (N_9370,N_3924,N_3793);
nor U9371 (N_9371,N_4675,N_4662);
xnor U9372 (N_9372,N_5444,N_3931);
or U9373 (N_9373,N_3491,N_4711);
or U9374 (N_9374,N_3184,N_5249);
nand U9375 (N_9375,N_8558,N_6577);
nor U9376 (N_9376,N_7381,N_8270);
and U9377 (N_9377,N_8352,N_9304);
xor U9378 (N_9378,N_8173,N_8796);
and U9379 (N_9379,N_7379,N_7889);
nand U9380 (N_9380,N_6722,N_7918);
nand U9381 (N_9381,N_7719,N_8390);
nor U9382 (N_9382,N_7455,N_7363);
nor U9383 (N_9383,N_9315,N_9138);
and U9384 (N_9384,N_6994,N_6342);
or U9385 (N_9385,N_6965,N_9020);
and U9386 (N_9386,N_7485,N_7390);
xor U9387 (N_9387,N_7953,N_6348);
xor U9388 (N_9388,N_8016,N_9357);
nor U9389 (N_9389,N_8486,N_7535);
nand U9390 (N_9390,N_8626,N_7039);
and U9391 (N_9391,N_8734,N_8949);
xor U9392 (N_9392,N_9082,N_8913);
nor U9393 (N_9393,N_8942,N_7740);
nor U9394 (N_9394,N_6907,N_7904);
xnor U9395 (N_9395,N_7433,N_8956);
nand U9396 (N_9396,N_8746,N_9210);
nand U9397 (N_9397,N_7271,N_8291);
or U9398 (N_9398,N_7632,N_6771);
nor U9399 (N_9399,N_8826,N_9229);
xnor U9400 (N_9400,N_8600,N_7623);
nand U9401 (N_9401,N_6833,N_8638);
xnor U9402 (N_9402,N_7417,N_6428);
xor U9403 (N_9403,N_8976,N_7490);
xor U9404 (N_9404,N_6708,N_8003);
nor U9405 (N_9405,N_7200,N_9206);
nor U9406 (N_9406,N_8569,N_9117);
xor U9407 (N_9407,N_8277,N_7835);
nand U9408 (N_9408,N_8218,N_8617);
or U9409 (N_9409,N_8192,N_7346);
or U9410 (N_9410,N_7681,N_6560);
nand U9411 (N_9411,N_6470,N_8762);
nor U9412 (N_9412,N_7569,N_8200);
nand U9413 (N_9413,N_8777,N_7619);
nand U9414 (N_9414,N_8404,N_8629);
nand U9415 (N_9415,N_6877,N_7182);
nand U9416 (N_9416,N_6905,N_9362);
and U9417 (N_9417,N_8232,N_8075);
nand U9418 (N_9418,N_8931,N_8407);
xnor U9419 (N_9419,N_8656,N_8363);
and U9420 (N_9420,N_8586,N_7571);
xnor U9421 (N_9421,N_7319,N_9267);
xnor U9422 (N_9422,N_6408,N_6400);
and U9423 (N_9423,N_8215,N_8310);
nand U9424 (N_9424,N_7907,N_6339);
xnor U9425 (N_9425,N_6357,N_9194);
or U9426 (N_9426,N_6576,N_7296);
xor U9427 (N_9427,N_6284,N_7176);
nor U9428 (N_9428,N_6731,N_8258);
nor U9429 (N_9429,N_8264,N_7261);
or U9430 (N_9430,N_7297,N_8188);
and U9431 (N_9431,N_6822,N_9277);
nor U9432 (N_9432,N_6613,N_6711);
xnor U9433 (N_9433,N_7664,N_7499);
xor U9434 (N_9434,N_6355,N_7680);
nand U9435 (N_9435,N_8639,N_8782);
and U9436 (N_9436,N_8707,N_8813);
nor U9437 (N_9437,N_9274,N_9182);
xnor U9438 (N_9438,N_8019,N_6785);
and U9439 (N_9439,N_7834,N_8991);
or U9440 (N_9440,N_6304,N_8533);
nand U9441 (N_9441,N_7576,N_7548);
or U9442 (N_9442,N_8353,N_6260);
nand U9443 (N_9443,N_8751,N_6287);
nor U9444 (N_9444,N_8087,N_7864);
xnor U9445 (N_9445,N_8061,N_8620);
or U9446 (N_9446,N_8437,N_7233);
nor U9447 (N_9447,N_6959,N_6475);
xor U9448 (N_9448,N_9107,N_6562);
or U9449 (N_9449,N_7057,N_7788);
or U9450 (N_9450,N_6948,N_7937);
xor U9451 (N_9451,N_8889,N_6914);
or U9452 (N_9452,N_7253,N_8424);
nand U9453 (N_9453,N_7149,N_7594);
nand U9454 (N_9454,N_7295,N_7503);
or U9455 (N_9455,N_7850,N_7803);
nand U9456 (N_9456,N_7055,N_6500);
or U9457 (N_9457,N_6601,N_6280);
and U9458 (N_9458,N_8810,N_6308);
nor U9459 (N_9459,N_8116,N_8293);
nand U9460 (N_9460,N_6430,N_6394);
xor U9461 (N_9461,N_7123,N_7066);
xor U9462 (N_9462,N_7940,N_6513);
and U9463 (N_9463,N_8550,N_8022);
and U9464 (N_9464,N_8925,N_8672);
nand U9465 (N_9465,N_7881,N_9359);
and U9466 (N_9466,N_7260,N_8175);
nand U9467 (N_9467,N_7711,N_6432);
and U9468 (N_9468,N_6866,N_8770);
or U9469 (N_9469,N_7956,N_9215);
nand U9470 (N_9470,N_8384,N_8780);
and U9471 (N_9471,N_8557,N_9333);
nor U9472 (N_9472,N_6397,N_6648);
and U9473 (N_9473,N_6952,N_9106);
nand U9474 (N_9474,N_7471,N_8104);
nor U9475 (N_9475,N_6492,N_8567);
and U9476 (N_9476,N_6688,N_6391);
nand U9477 (N_9477,N_7190,N_6756);
xnor U9478 (N_9478,N_8274,N_8530);
nor U9479 (N_9479,N_8021,N_7423);
or U9480 (N_9480,N_7321,N_8880);
nand U9481 (N_9481,N_8686,N_7194);
xor U9482 (N_9482,N_6457,N_7432);
or U9483 (N_9483,N_8864,N_8484);
nor U9484 (N_9484,N_7948,N_6401);
or U9485 (N_9485,N_9024,N_7464);
and U9486 (N_9486,N_9162,N_9166);
nor U9487 (N_9487,N_6776,N_9337);
xor U9488 (N_9488,N_8323,N_6981);
nor U9489 (N_9489,N_7345,N_8634);
nor U9490 (N_9490,N_8729,N_8189);
nand U9491 (N_9491,N_6813,N_8972);
and U9492 (N_9492,N_9156,N_9312);
nand U9493 (N_9493,N_8213,N_7896);
nand U9494 (N_9494,N_7011,N_7430);
or U9495 (N_9495,N_7515,N_6980);
xnor U9496 (N_9496,N_7671,N_7970);
xor U9497 (N_9497,N_9339,N_8472);
and U9498 (N_9498,N_8026,N_6528);
nand U9499 (N_9499,N_9064,N_8070);
nand U9500 (N_9500,N_9147,N_7702);
or U9501 (N_9501,N_7308,N_6956);
xor U9502 (N_9502,N_7924,N_8135);
xor U9503 (N_9503,N_9113,N_8236);
or U9504 (N_9504,N_8413,N_7531);
and U9505 (N_9505,N_7034,N_8932);
nand U9506 (N_9506,N_8955,N_8033);
or U9507 (N_9507,N_8903,N_7580);
and U9508 (N_9508,N_8408,N_9042);
nor U9509 (N_9509,N_8677,N_8917);
xor U9510 (N_9510,N_7400,N_8083);
or U9511 (N_9511,N_6288,N_7354);
nor U9512 (N_9512,N_9004,N_7330);
xor U9513 (N_9513,N_7765,N_9356);
and U9514 (N_9514,N_7058,N_7310);
nor U9515 (N_9515,N_9136,N_7942);
nand U9516 (N_9516,N_6379,N_7779);
nand U9517 (N_9517,N_6449,N_6422);
nor U9518 (N_9518,N_7446,N_6932);
or U9519 (N_9519,N_6552,N_9355);
xnor U9520 (N_9520,N_6325,N_6460);
or U9521 (N_9521,N_7749,N_6818);
or U9522 (N_9522,N_9114,N_7701);
or U9523 (N_9523,N_9235,N_6464);
nor U9524 (N_9524,N_7408,N_7673);
nor U9525 (N_9525,N_8082,N_8900);
xor U9526 (N_9526,N_8100,N_6774);
or U9527 (N_9527,N_9121,N_9021);
and U9528 (N_9528,N_8670,N_7715);
or U9529 (N_9529,N_7497,N_6693);
xnor U9530 (N_9530,N_8510,N_6595);
or U9531 (N_9531,N_8833,N_8548);
nor U9532 (N_9532,N_7186,N_6508);
nor U9533 (N_9533,N_7699,N_9092);
and U9534 (N_9534,N_8801,N_8092);
nor U9535 (N_9535,N_7908,N_7695);
nand U9536 (N_9536,N_6579,N_8918);
and U9537 (N_9537,N_7344,N_7537);
or U9538 (N_9538,N_9273,N_8417);
or U9539 (N_9539,N_7020,N_8679);
nor U9540 (N_9540,N_7313,N_6502);
and U9541 (N_9541,N_7006,N_7088);
or U9542 (N_9542,N_7267,N_9264);
and U9543 (N_9543,N_8910,N_8152);
and U9544 (N_9544,N_9071,N_9044);
nor U9545 (N_9545,N_8299,N_7874);
and U9546 (N_9546,N_8851,N_6714);
nand U9547 (N_9547,N_6456,N_9072);
xnor U9548 (N_9548,N_8093,N_7627);
xnor U9549 (N_9549,N_7429,N_9015);
nor U9550 (N_9550,N_6605,N_7427);
nor U9551 (N_9551,N_6939,N_8077);
and U9552 (N_9552,N_7293,N_6709);
or U9553 (N_9553,N_8978,N_9031);
xnor U9554 (N_9554,N_7744,N_8308);
nand U9555 (N_9555,N_7934,N_8845);
and U9556 (N_9556,N_6778,N_7480);
nor U9557 (N_9557,N_7553,N_8364);
nand U9558 (N_9558,N_6309,N_9151);
nor U9559 (N_9559,N_7631,N_7929);
nand U9560 (N_9560,N_7947,N_7837);
xnor U9561 (N_9561,N_7359,N_7893);
nand U9562 (N_9562,N_8186,N_8563);
or U9563 (N_9563,N_8059,N_6719);
nand U9564 (N_9564,N_9130,N_7324);
and U9565 (N_9565,N_6259,N_9100);
and U9566 (N_9566,N_7789,N_8793);
nor U9567 (N_9567,N_7726,N_7214);
and U9568 (N_9568,N_8879,N_7770);
nand U9569 (N_9569,N_6979,N_8469);
and U9570 (N_9570,N_8919,N_7759);
nor U9571 (N_9571,N_6935,N_7596);
nand U9572 (N_9572,N_7298,N_6689);
nand U9573 (N_9573,N_7349,N_7509);
and U9574 (N_9574,N_6574,N_6646);
nor U9575 (N_9575,N_7618,N_9228);
nand U9576 (N_9576,N_6406,N_7172);
or U9577 (N_9577,N_7550,N_8090);
and U9578 (N_9578,N_9211,N_8276);
or U9579 (N_9579,N_7820,N_8279);
nor U9580 (N_9580,N_8316,N_9327);
nor U9581 (N_9581,N_7243,N_9016);
xnor U9582 (N_9582,N_6992,N_8088);
or U9583 (N_9583,N_9374,N_7845);
nor U9584 (N_9584,N_9281,N_7614);
xnor U9585 (N_9585,N_9157,N_7179);
nor U9586 (N_9586,N_8724,N_7168);
or U9587 (N_9587,N_9116,N_8004);
xnor U9588 (N_9588,N_7031,N_6911);
nand U9589 (N_9589,N_7534,N_7115);
and U9590 (N_9590,N_8199,N_6323);
nor U9591 (N_9591,N_9017,N_6346);
xor U9592 (N_9592,N_8178,N_7577);
or U9593 (N_9593,N_7518,N_6593);
nand U9594 (N_9594,N_8655,N_6333);
nand U9595 (N_9595,N_6950,N_7004);
nor U9596 (N_9596,N_7582,N_7751);
xor U9597 (N_9597,N_6820,N_9124);
xnor U9598 (N_9598,N_8761,N_7668);
and U9599 (N_9599,N_6518,N_9078);
or U9600 (N_9600,N_7294,N_7292);
nand U9601 (N_9601,N_9139,N_8901);
xor U9602 (N_9602,N_8259,N_6536);
nor U9603 (N_9603,N_9291,N_7717);
xnor U9604 (N_9604,N_7470,N_8052);
or U9605 (N_9605,N_8053,N_6555);
nor U9606 (N_9606,N_8485,N_8792);
nand U9607 (N_9607,N_9296,N_7764);
nor U9608 (N_9608,N_7989,N_6766);
or U9609 (N_9609,N_8349,N_7638);
and U9610 (N_9610,N_6515,N_8504);
xor U9611 (N_9611,N_9148,N_7752);
xnor U9612 (N_9612,N_7549,N_7022);
nand U9613 (N_9613,N_7552,N_6772);
or U9614 (N_9614,N_9349,N_7921);
nor U9615 (N_9615,N_7561,N_6834);
nor U9616 (N_9616,N_7723,N_9019);
or U9617 (N_9617,N_7449,N_6807);
xor U9618 (N_9618,N_9257,N_6459);
nor U9619 (N_9619,N_7409,N_6919);
xor U9620 (N_9620,N_7683,N_6344);
and U9621 (N_9621,N_6861,N_6967);
and U9622 (N_9622,N_9321,N_7524);
xnor U9623 (N_9623,N_7257,N_7675);
and U9624 (N_9624,N_7622,N_8416);
or U9625 (N_9625,N_6694,N_8970);
and U9626 (N_9626,N_9027,N_6541);
nor U9627 (N_9627,N_7332,N_7528);
xor U9628 (N_9628,N_7091,N_8318);
and U9629 (N_9629,N_6584,N_8062);
nand U9630 (N_9630,N_9104,N_8262);
or U9631 (N_9631,N_8819,N_9090);
and U9632 (N_9632,N_7444,N_7072);
nand U9633 (N_9633,N_7670,N_6377);
nand U9634 (N_9634,N_7256,N_6479);
nand U9635 (N_9635,N_6856,N_8419);
and U9636 (N_9636,N_7096,N_8755);
nor U9637 (N_9637,N_6519,N_7230);
and U9638 (N_9638,N_8466,N_8089);
nor U9639 (N_9639,N_6496,N_6802);
or U9640 (N_9640,N_6473,N_8006);
nand U9641 (N_9641,N_8939,N_7090);
xor U9642 (N_9642,N_8676,N_7276);
or U9643 (N_9643,N_8517,N_9313);
nand U9644 (N_9644,N_8209,N_7781);
nor U9645 (N_9645,N_7236,N_6512);
and U9646 (N_9646,N_9170,N_7394);
xnor U9647 (N_9647,N_6989,N_7830);
nor U9648 (N_9648,N_8580,N_9222);
and U9649 (N_9649,N_6331,N_8072);
xor U9650 (N_9650,N_6295,N_7395);
and U9651 (N_9651,N_8643,N_8559);
xnor U9652 (N_9652,N_8314,N_7225);
or U9653 (N_9653,N_7496,N_8311);
xor U9654 (N_9654,N_7865,N_9036);
nor U9655 (N_9655,N_9133,N_7059);
nor U9656 (N_9656,N_8037,N_8776);
nand U9657 (N_9657,N_7502,N_8205);
nor U9658 (N_9658,N_9295,N_9343);
nand U9659 (N_9659,N_9174,N_6987);
nand U9660 (N_9660,N_7646,N_8301);
or U9661 (N_9661,N_6354,N_7241);
and U9662 (N_9662,N_6477,N_8275);
xor U9663 (N_9663,N_9331,N_7322);
nor U9664 (N_9664,N_8440,N_8582);
nor U9665 (N_9665,N_6817,N_6812);
and U9666 (N_9666,N_8842,N_6926);
or U9667 (N_9667,N_7911,N_6419);
nand U9668 (N_9668,N_8921,N_6871);
and U9669 (N_9669,N_8807,N_8382);
and U9670 (N_9670,N_7666,N_6891);
nand U9671 (N_9671,N_9262,N_7700);
nor U9672 (N_9672,N_7265,N_6435);
xnor U9673 (N_9673,N_6368,N_7285);
nor U9674 (N_9674,N_7076,N_8773);
or U9675 (N_9675,N_7734,N_6361);
xor U9676 (N_9676,N_8946,N_7126);
nor U9677 (N_9677,N_8476,N_8568);
nor U9678 (N_9678,N_9067,N_9176);
xnor U9679 (N_9679,N_7750,N_7971);
xor U9680 (N_9680,N_8953,N_8195);
or U9681 (N_9681,N_6307,N_6525);
xor U9682 (N_9682,N_7604,N_7574);
nor U9683 (N_9683,N_6968,N_7463);
nor U9684 (N_9684,N_7955,N_9048);
and U9685 (N_9685,N_7370,N_7676);
or U9686 (N_9686,N_9217,N_6622);
xor U9687 (N_9687,N_8696,N_8641);
xor U9688 (N_9688,N_8378,N_6250);
nor U9689 (N_9689,N_8944,N_8321);
nand U9690 (N_9690,N_8852,N_9294);
and U9691 (N_9691,N_6489,N_7800);
nand U9692 (N_9692,N_9171,N_7008);
xnor U9693 (N_9693,N_7416,N_7448);
nand U9694 (N_9694,N_8683,N_6350);
xnor U9695 (N_9695,N_7337,N_7883);
nand U9696 (N_9696,N_7768,N_6749);
xnor U9697 (N_9697,N_8391,N_6254);
xnor U9698 (N_9698,N_6626,N_8227);
or U9699 (N_9699,N_8772,N_8123);
or U9700 (N_9700,N_7647,N_9189);
nand U9701 (N_9701,N_6588,N_9317);
and U9702 (N_9702,N_8344,N_9086);
xor U9703 (N_9703,N_7218,N_9069);
or U9704 (N_9704,N_9198,N_8817);
nor U9705 (N_9705,N_6399,N_7861);
nand U9706 (N_9706,N_6970,N_8165);
nand U9707 (N_9707,N_7204,N_9224);
xor U9708 (N_9708,N_6851,N_6910);
or U9709 (N_9709,N_8487,N_7389);
and U9710 (N_9710,N_8678,N_8841);
xor U9711 (N_9711,N_9268,N_6462);
nor U9712 (N_9712,N_9325,N_6266);
nand U9713 (N_9713,N_6879,N_8861);
xor U9714 (N_9714,N_7380,N_7851);
xor U9715 (N_9715,N_7161,N_7035);
nand U9716 (N_9716,N_7650,N_8511);
nand U9717 (N_9717,N_8374,N_7262);
and U9718 (N_9718,N_8716,N_9208);
nand U9719 (N_9719,N_7517,N_6892);
nand U9720 (N_9720,N_6523,N_7049);
and U9721 (N_9721,N_6740,N_9196);
or U9722 (N_9722,N_7806,N_8140);
and U9723 (N_9723,N_8224,N_8572);
nand U9724 (N_9724,N_7897,N_7986);
or U9725 (N_9725,N_7424,N_9050);
and U9726 (N_9726,N_9115,N_7603);
xor U9727 (N_9727,N_8065,N_6691);
or U9728 (N_9728,N_7547,N_6300);
nor U9729 (N_9729,N_8884,N_6692);
or U9730 (N_9730,N_9038,N_8779);
or U9731 (N_9731,N_9289,N_8372);
nand U9732 (N_9732,N_6410,N_8589);
xor U9733 (N_9733,N_6609,N_6839);
xor U9734 (N_9734,N_6424,N_8714);
nor U9735 (N_9735,N_6286,N_9261);
or U9736 (N_9736,N_7500,N_7086);
nor U9737 (N_9737,N_7554,N_6947);
nand U9738 (N_9738,N_7320,N_8994);
or U9739 (N_9739,N_6949,N_7654);
or U9740 (N_9740,N_9328,N_8333);
nor U9741 (N_9741,N_6938,N_7141);
xor U9742 (N_9742,N_9018,N_8127);
and U9743 (N_9743,N_7142,N_7251);
nor U9744 (N_9744,N_8234,N_8534);
or U9745 (N_9745,N_9367,N_7069);
nand U9746 (N_9746,N_9122,N_6921);
and U9747 (N_9747,N_6543,N_7888);
and U9748 (N_9748,N_8605,N_9088);
xor U9749 (N_9749,N_9103,N_8957);
and U9750 (N_9750,N_7697,N_7617);
and U9751 (N_9751,N_7629,N_7613);
nor U9752 (N_9752,N_7107,N_7546);
nand U9753 (N_9753,N_8112,N_8595);
or U9754 (N_9754,N_7729,N_8074);
nand U9755 (N_9755,N_7633,N_7223);
nand U9756 (N_9756,N_9158,N_6262);
xnor U9757 (N_9757,N_6436,N_8478);
and U9758 (N_9758,N_8063,N_7121);
xor U9759 (N_9759,N_7915,N_7930);
and U9760 (N_9760,N_7189,N_8837);
xor U9761 (N_9761,N_8682,N_9146);
or U9762 (N_9762,N_8607,N_8313);
and U9763 (N_9763,N_8920,N_9282);
nor U9764 (N_9764,N_6700,N_6514);
and U9765 (N_9765,N_8536,N_6381);
and U9766 (N_9766,N_7763,N_8863);
xnor U9767 (N_9767,N_6603,N_7824);
nor U9768 (N_9768,N_6920,N_6780);
nor U9769 (N_9769,N_8376,N_7421);
nor U9770 (N_9770,N_7341,N_6864);
and U9771 (N_9771,N_7491,N_8736);
xor U9772 (N_9772,N_6794,N_6872);
xor U9773 (N_9773,N_6942,N_8969);
and U9774 (N_9774,N_7145,N_7761);
xnor U9775 (N_9775,N_9271,N_8493);
nand U9776 (N_9776,N_8035,N_7543);
nand U9777 (N_9777,N_7277,N_8386);
or U9778 (N_9778,N_8351,N_7351);
xor U9779 (N_9779,N_6825,N_8608);
and U9780 (N_9780,N_9209,N_8397);
or U9781 (N_9781,N_9056,N_6885);
nand U9782 (N_9782,N_7634,N_6697);
nand U9783 (N_9783,N_7616,N_8396);
or U9784 (N_9784,N_9254,N_9097);
nand U9785 (N_9785,N_7095,N_6695);
nand U9786 (N_9786,N_6824,N_8170);
xnor U9787 (N_9787,N_7507,N_7963);
or U9788 (N_9788,N_6608,N_6827);
or U9789 (N_9789,N_8719,N_6553);
xnor U9790 (N_9790,N_6372,N_6614);
and U9791 (N_9791,N_7544,N_7706);
and U9792 (N_9792,N_8695,N_6962);
and U9793 (N_9793,N_7157,N_8410);
or U9794 (N_9794,N_6330,N_9179);
nor U9795 (N_9795,N_8730,N_8219);
nand U9796 (N_9796,N_8666,N_9350);
xnor U9797 (N_9797,N_7884,N_7688);
nor U9798 (N_9798,N_7570,N_7590);
xor U9799 (N_9799,N_6738,N_7026);
nor U9800 (N_9800,N_6386,N_6815);
nand U9801 (N_9801,N_7775,N_7705);
or U9802 (N_9802,N_7746,N_8149);
xor U9803 (N_9803,N_7002,N_7127);
or U9804 (N_9804,N_7636,N_8541);
and U9805 (N_9805,N_6316,N_7108);
nand U9806 (N_9806,N_6918,N_6955);
xor U9807 (N_9807,N_6627,N_8768);
nor U9808 (N_9808,N_8742,N_7438);
or U9809 (N_9809,N_7643,N_7060);
nand U9810 (N_9810,N_8652,N_9256);
xnor U9811 (N_9811,N_7070,N_8139);
nor U9812 (N_9812,N_8532,N_8235);
nor U9813 (N_9813,N_6854,N_6283);
xor U9814 (N_9814,N_6638,N_7109);
nor U9815 (N_9815,N_6390,N_7945);
nand U9816 (N_9816,N_6842,N_7084);
nand U9817 (N_9817,N_6660,N_8041);
nor U9818 (N_9818,N_6612,N_7099);
nor U9819 (N_9819,N_8644,N_8373);
xnor U9820 (N_9820,N_8214,N_7626);
nor U9821 (N_9821,N_8247,N_7532);
or U9822 (N_9822,N_8324,N_7988);
or U9823 (N_9823,N_6298,N_7876);
nor U9824 (N_9824,N_7611,N_8286);
nor U9825 (N_9825,N_7027,N_8184);
nand U9826 (N_9826,N_8265,N_7335);
nor U9827 (N_9827,N_6468,N_7718);
xor U9828 (N_9828,N_8977,N_8951);
and U9829 (N_9829,N_8781,N_7826);
nor U9830 (N_9830,N_8181,N_7974);
nor U9831 (N_9831,N_6409,N_7713);
and U9832 (N_9832,N_7445,N_7239);
and U9833 (N_9833,N_7453,N_8630);
or U9834 (N_9834,N_9059,N_8565);
nand U9835 (N_9835,N_6846,N_8163);
nand U9836 (N_9836,N_7962,N_7252);
nand U9837 (N_9837,N_7735,N_8624);
xor U9838 (N_9838,N_7694,N_8549);
nand U9839 (N_9839,N_6800,N_6426);
or U9840 (N_9840,N_7756,N_8023);
and U9841 (N_9841,N_7386,N_7419);
xor U9842 (N_9842,N_6369,N_7476);
nor U9843 (N_9843,N_6299,N_7871);
or U9844 (N_9844,N_8387,N_8269);
nor U9845 (N_9845,N_8583,N_6944);
nor U9846 (N_9846,N_7198,N_8816);
or U9847 (N_9847,N_7693,N_8136);
or U9848 (N_9848,N_7965,N_6971);
or U9849 (N_9849,N_7562,N_9241);
nor U9850 (N_9850,N_6466,N_7289);
nor U9851 (N_9851,N_9276,N_7374);
nor U9852 (N_9852,N_6639,N_7103);
or U9853 (N_9853,N_7238,N_6370);
xnor U9854 (N_9854,N_8505,N_9353);
and U9855 (N_9855,N_7520,N_8432);
nor U9856 (N_9856,N_6810,N_8710);
or U9857 (N_9857,N_6685,N_6748);
or U9858 (N_9858,N_7234,N_8658);
xnor U9859 (N_9859,N_7658,N_8637);
nor U9860 (N_9860,N_8456,N_8645);
nor U9861 (N_9861,N_8046,N_8740);
xnor U9862 (N_9862,N_7958,N_8657);
or U9863 (N_9863,N_9351,N_7829);
and U9864 (N_9864,N_6592,N_8723);
nor U9865 (N_9865,N_7005,N_6654);
and U9866 (N_9866,N_7143,N_6717);
and U9867 (N_9867,N_8094,N_8718);
xor U9868 (N_9868,N_8101,N_6382);
xor U9869 (N_9869,N_6850,N_7466);
nand U9870 (N_9870,N_7221,N_8327);
and U9871 (N_9871,N_6371,N_6684);
or U9872 (N_9872,N_6253,N_8086);
nor U9873 (N_9873,N_9112,N_9183);
nor U9874 (N_9874,N_8488,N_7923);
nand U9875 (N_9875,N_9129,N_6624);
nor U9876 (N_9876,N_6427,N_8108);
or U9877 (N_9877,N_6779,N_8196);
or U9878 (N_9878,N_8687,N_6440);
nand U9879 (N_9879,N_7131,N_8744);
and U9880 (N_9880,N_6447,N_8442);
and U9881 (N_9881,N_7721,N_7707);
xnor U9882 (N_9882,N_6465,N_6874);
or U9883 (N_9883,N_7928,N_6991);
nand U9884 (N_9884,N_6568,N_6775);
or U9885 (N_9885,N_6265,N_7787);
or U9886 (N_9886,N_8650,N_8412);
and U9887 (N_9887,N_7224,N_9242);
or U9888 (N_9888,N_6486,N_8692);
nand U9889 (N_9889,N_7880,N_6602);
nand U9890 (N_9890,N_7199,N_6611);
xnor U9891 (N_9891,N_7894,N_7484);
xor U9892 (N_9892,N_7565,N_8481);
nand U9893 (N_9893,N_6929,N_8261);
nand U9894 (N_9894,N_6610,N_8519);
xor U9895 (N_9895,N_6535,N_7903);
nor U9896 (N_9896,N_8409,N_6702);
xnor U9897 (N_9897,N_7075,N_7213);
and U9898 (N_9898,N_8590,N_7376);
and U9899 (N_9899,N_8164,N_7679);
nand U9900 (N_9900,N_6777,N_8054);
nor U9901 (N_9901,N_8206,N_8706);
xnor U9902 (N_9902,N_6957,N_8296);
xnor U9903 (N_9903,N_7808,N_8524);
and U9904 (N_9904,N_6782,N_9324);
and U9905 (N_9905,N_6586,N_7101);
nor U9906 (N_9906,N_6754,N_6924);
nor U9907 (N_9907,N_6452,N_9137);
xnor U9908 (N_9908,N_6922,N_6418);
nor U9909 (N_9909,N_7600,N_7475);
xnor U9910 (N_9910,N_8475,N_8085);
and U9911 (N_9911,N_6497,N_7525);
xnor U9912 (N_9912,N_7120,N_6385);
and U9913 (N_9913,N_8787,N_8312);
and U9914 (N_9914,N_7973,N_7207);
and U9915 (N_9915,N_8506,N_7110);
xor U9916 (N_9916,N_8011,N_8553);
and U9917 (N_9917,N_6760,N_7483);
or U9918 (N_9918,N_9009,N_9040);
nor U9919 (N_9919,N_7154,N_6366);
nand U9920 (N_9920,N_6768,N_7393);
or U9921 (N_9921,N_8552,N_7169);
and U9922 (N_9922,N_8783,N_8454);
or U9923 (N_9923,N_8330,N_8434);
xor U9924 (N_9924,N_8790,N_8698);
xnor U9925 (N_9925,N_8470,N_8874);
xor U9926 (N_9926,N_8579,N_9204);
nor U9927 (N_9927,N_9223,N_8750);
and U9928 (N_9928,N_7906,N_7967);
or U9929 (N_9929,N_8320,N_8513);
nor U9930 (N_9930,N_6358,N_8223);
nor U9931 (N_9931,N_6559,N_7273);
or U9932 (N_9932,N_8893,N_7593);
and U9933 (N_9933,N_8537,N_7657);
nand U9934 (N_9934,N_7720,N_9239);
and U9935 (N_9935,N_7118,N_8522);
nand U9936 (N_9936,N_7458,N_7441);
or U9937 (N_9937,N_6889,N_8674);
or U9938 (N_9938,N_7040,N_7648);
nand U9939 (N_9939,N_7891,N_7831);
or U9940 (N_9940,N_9058,N_6450);
or U9941 (N_9941,N_7796,N_9269);
nand U9942 (N_9942,N_7291,N_6533);
or U9943 (N_9943,N_6607,N_7191);
or U9944 (N_9944,N_8797,N_8131);
xnor U9945 (N_9945,N_7226,N_6597);
xor U9946 (N_9946,N_6509,N_8025);
or U9947 (N_9947,N_6521,N_7925);
nand U9948 (N_9948,N_8615,N_8334);
and U9949 (N_9949,N_6799,N_7944);
or U9950 (N_9950,N_8172,N_9080);
nand U9951 (N_9951,N_8347,N_7556);
nor U9952 (N_9952,N_8044,N_8985);
and U9953 (N_9953,N_9041,N_6567);
nor U9954 (N_9954,N_7437,N_7357);
and U9955 (N_9955,N_6961,N_8515);
nand U9956 (N_9956,N_6630,N_7197);
or U9957 (N_9957,N_7949,N_7651);
and U9958 (N_9958,N_6665,N_7637);
nor U9959 (N_9959,N_9190,N_6291);
xor U9960 (N_9960,N_6735,N_7065);
and U9961 (N_9961,N_6364,N_7434);
nor U9962 (N_9962,N_7964,N_7817);
or U9963 (N_9963,N_9290,N_6937);
xnor U9964 (N_9964,N_8176,N_7802);
and U9965 (N_9965,N_7478,N_8272);
xnor U9966 (N_9966,N_6687,N_6977);
nand U9967 (N_9967,N_9248,N_8499);
and U9968 (N_9968,N_9293,N_9070);
nor U9969 (N_9969,N_8829,N_6642);
nand U9970 (N_9970,N_8467,N_6335);
nand U9971 (N_9971,N_8285,N_6556);
xnor U9972 (N_9972,N_8986,N_7954);
nand U9973 (N_9973,N_8007,N_7405);
nand U9974 (N_9974,N_7079,N_7979);
xor U9975 (N_9975,N_6786,N_9372);
and U9976 (N_9976,N_6471,N_7698);
and U9977 (N_9977,N_6902,N_8675);
xnor U9978 (N_9978,N_6761,N_7085);
and U9979 (N_9979,N_7809,N_8241);
xor U9980 (N_9980,N_7999,N_9087);
nand U9981 (N_9981,N_7783,N_8883);
nand U9982 (N_9982,N_7539,N_6663);
nor U9983 (N_9983,N_8317,N_6909);
nor U9984 (N_9984,N_9079,N_7209);
nor U9985 (N_9985,N_6897,N_6783);
or U9986 (N_9986,N_7813,N_6941);
and U9987 (N_9987,N_7890,N_6545);
or U9988 (N_9988,N_6988,N_8287);
nand U9989 (N_9989,N_8207,N_6867);
xor U9990 (N_9990,N_8566,N_9238);
nor U9991 (N_9991,N_6405,N_8667);
xor U9992 (N_9992,N_8663,N_6506);
or U9993 (N_9993,N_9307,N_9149);
nor U9994 (N_9994,N_8905,N_7382);
nor U9995 (N_9995,N_6281,N_7919);
xnor U9996 (N_9996,N_8873,N_8881);
nand U9997 (N_9997,N_6585,N_6458);
xor U9998 (N_9998,N_9314,N_9332);
or U9999 (N_9999,N_8963,N_8018);
or U10000 (N_10000,N_9323,N_7722);
nand U10001 (N_10001,N_9076,N_6884);
nor U10002 (N_10002,N_8989,N_8221);
and U10003 (N_10003,N_8297,N_8471);
nor U10004 (N_10004,N_8872,N_6831);
and U10005 (N_10005,N_6599,N_7208);
and U10006 (N_10006,N_7050,N_6882);
or U10007 (N_10007,N_7150,N_9192);
or U10008 (N_10008,N_9260,N_7960);
xnor U10009 (N_10009,N_7573,N_9308);
or U10010 (N_10010,N_8853,N_8886);
nor U10011 (N_10011,N_7201,N_9300);
or U10012 (N_10012,N_6395,N_8115);
xor U10013 (N_10013,N_6289,N_7385);
nand U10014 (N_10014,N_6278,N_7348);
nor U10015 (N_10015,N_6797,N_6703);
or U10016 (N_10016,N_8421,N_8614);
and U10017 (N_10017,N_7018,N_8362);
nor U10018 (N_10018,N_9259,N_8411);
or U10019 (N_10019,N_7038,N_8602);
xor U10020 (N_10020,N_7373,N_7425);
or U10021 (N_10021,N_8788,N_6946);
nor U10022 (N_10022,N_7983,N_8134);
xnor U10023 (N_10023,N_8381,N_8854);
and U10024 (N_10024,N_8907,N_6356);
or U10025 (N_10025,N_8890,N_6312);
nor U10026 (N_10026,N_6875,N_9341);
nor U10027 (N_10027,N_8616,N_7307);
or U10028 (N_10028,N_8721,N_6451);
or U10029 (N_10029,N_8067,N_7860);
and U10030 (N_10030,N_7268,N_7899);
and U10031 (N_10031,N_8594,N_8305);
nor U10032 (N_10032,N_8828,N_7976);
or U10033 (N_10033,N_7366,N_9280);
nand U10034 (N_10034,N_7579,N_9197);
xnor U10035 (N_10035,N_8665,N_7435);
or U10036 (N_10036,N_7773,N_8965);
nor U10037 (N_10037,N_7886,N_9062);
or U10038 (N_10038,N_9063,N_7966);
or U10039 (N_10039,N_6261,N_8498);
nand U10040 (N_10040,N_8030,N_8202);
and U10041 (N_10041,N_8839,N_7083);
nand U10042 (N_10042,N_9180,N_9169);
and U10043 (N_10043,N_8747,N_7170);
nor U10044 (N_10044,N_6744,N_6388);
nor U10045 (N_10045,N_7978,N_7347);
nor U10046 (N_10046,N_8243,N_8545);
nor U10047 (N_10047,N_7842,N_8341);
nand U10048 (N_10048,N_7910,N_6582);
xor U10049 (N_10049,N_8457,N_8621);
and U10050 (N_10050,N_9014,N_8906);
nand U10051 (N_10051,N_7951,N_8694);
nand U10052 (N_10052,N_9142,N_9008);
or U10053 (N_10053,N_8266,N_7935);
and U10054 (N_10054,N_7557,N_8604);
xor U10055 (N_10055,N_6631,N_7367);
and U10056 (N_10056,N_9184,N_9243);
nand U10057 (N_10057,N_8802,N_8180);
xor U10058 (N_10058,N_6444,N_7882);
or U10059 (N_10059,N_9022,N_8860);
nand U10060 (N_10060,N_8036,N_9025);
and U10061 (N_10061,N_6376,N_7092);
nand U10062 (N_10062,N_7846,N_9026);
nor U10063 (N_10063,N_7612,N_7377);
or U10064 (N_10064,N_6269,N_9152);
nand U10065 (N_10065,N_9195,N_6343);
xnor U10066 (N_10066,N_7739,N_6434);
nor U10067 (N_10067,N_7832,N_7284);
nor U10068 (N_10068,N_8823,N_8578);
nor U10069 (N_10069,N_8785,N_9134);
nand U10070 (N_10070,N_7997,N_8952);
or U10071 (N_10071,N_8526,N_6755);
or U10072 (N_10072,N_7645,N_7420);
xor U10073 (N_10073,N_6499,N_7361);
and U10074 (N_10074,N_7329,N_6633);
xnor U10075 (N_10075,N_7007,N_8882);
xnor U10076 (N_10076,N_6617,N_6495);
or U10077 (N_10077,N_6742,N_8256);
or U10078 (N_10078,N_8640,N_7229);
nor U10079 (N_10079,N_8961,N_7812);
or U10080 (N_10080,N_7311,N_6561);
or U10081 (N_10081,N_6532,N_9089);
nor U10082 (N_10082,N_6681,N_6484);
xor U10083 (N_10083,N_9029,N_7669);
or U10084 (N_10084,N_7667,N_9275);
or U10085 (N_10085,N_7384,N_8896);
nor U10086 (N_10086,N_8244,N_8848);
nand U10087 (N_10087,N_9126,N_7914);
nand U10088 (N_10088,N_8960,N_7135);
nor U10089 (N_10089,N_7828,N_8445);
or U10090 (N_10090,N_7178,N_9068);
and U10091 (N_10091,N_8335,N_8642);
or U10092 (N_10092,N_8480,N_8997);
and U10093 (N_10093,N_9244,N_6798);
nand U10094 (N_10094,N_6855,N_7331);
nor U10095 (N_10095,N_7468,N_7857);
and U10096 (N_10096,N_6791,N_8745);
xor U10097 (N_10097,N_8166,N_8468);
and U10098 (N_10098,N_9286,N_6849);
or U10099 (N_10099,N_8878,N_6563);
nand U10100 (N_10100,N_7100,N_9246);
or U10101 (N_10101,N_8885,N_8167);
nand U10102 (N_10102,N_9081,N_7663);
nor U10103 (N_10103,N_7074,N_9340);
or U10104 (N_10104,N_7443,N_8251);
nor U10105 (N_10105,N_9159,N_7456);
or U10106 (N_10106,N_7859,N_6726);
nand U10107 (N_10107,N_9368,N_7129);
nand U10108 (N_10108,N_7686,N_8280);
xor U10109 (N_10109,N_6415,N_9110);
and U10110 (N_10110,N_7212,N_6310);
nand U10111 (N_10111,N_9233,N_9083);
and U10112 (N_10112,N_9249,N_7353);
or U10113 (N_10113,N_8073,N_8651);
or U10114 (N_10114,N_8934,N_6990);
nand U10115 (N_10115,N_7714,N_7998);
xnor U10116 (N_10116,N_8805,N_8571);
or U10117 (N_10117,N_8009,N_7833);
or U10118 (N_10118,N_6759,N_7450);
or U10119 (N_10119,N_7167,N_7422);
xnor U10120 (N_10120,N_8439,N_7290);
nor U10121 (N_10121,N_8507,N_7440);
or U10122 (N_10122,N_6690,N_8119);
nand U10123 (N_10123,N_8700,N_8727);
or U10124 (N_10124,N_6472,N_8555);
and U10125 (N_10125,N_8246,N_8154);
nor U10126 (N_10126,N_9292,N_8923);
or U10127 (N_10127,N_8340,N_7938);
or U10128 (N_10128,N_8503,N_7533);
xor U10129 (N_10129,N_6540,N_6365);
and U10130 (N_10130,N_6590,N_8619);
xnor U10131 (N_10131,N_7584,N_9205);
nor U10132 (N_10132,N_7113,N_7498);
and U10133 (N_10133,N_7585,N_7474);
or U10134 (N_10134,N_6318,N_8359);
nor U10135 (N_10135,N_9108,N_8847);
nand U10136 (N_10136,N_9285,N_8474);
and U10137 (N_10137,N_8292,N_7682);
or U10138 (N_10138,N_7943,N_6656);
or U10139 (N_10139,N_8725,N_8664);
or U10140 (N_10140,N_7990,N_8928);
and U10141 (N_10141,N_8483,N_6569);
and U10142 (N_10142,N_7275,N_8013);
nand U10143 (N_10143,N_8859,N_7447);
xor U10144 (N_10144,N_8060,N_8988);
or U10145 (N_10145,N_7659,N_8446);
and U10146 (N_10146,N_9361,N_8260);
nand U10147 (N_10147,N_7356,N_7769);
and U10148 (N_10148,N_9309,N_6953);
or U10149 (N_10149,N_8584,N_8838);
and U10150 (N_10150,N_7064,N_7451);
and U10151 (N_10151,N_8850,N_8835);
nand U10152 (N_10152,N_8211,N_6683);
nor U10153 (N_10153,N_8668,N_7854);
or U10154 (N_10154,N_9207,N_6321);
or U10155 (N_10155,N_6557,N_8930);
xor U10156 (N_10156,N_7048,N_6267);
nand U10157 (N_10157,N_7665,N_7687);
nand U10158 (N_10158,N_7242,N_6538);
or U10159 (N_10159,N_7028,N_8319);
xor U10160 (N_10160,N_7398,N_6268);
nor U10161 (N_10161,N_7219,N_8701);
nor U10162 (N_10162,N_7228,N_7323);
or U10163 (N_10163,N_6913,N_7704);
nor U10164 (N_10164,N_8096,N_7309);
xnor U10165 (N_10165,N_9141,N_8754);
and U10166 (N_10166,N_7641,N_8795);
or U10167 (N_10167,N_9173,N_6662);
and U10168 (N_10168,N_8784,N_6455);
xnor U10169 (N_10169,N_7766,N_8429);
xnor U10170 (N_10170,N_9013,N_7661);
nor U10171 (N_10171,N_7875,N_8898);
nor U10172 (N_10172,N_8581,N_9095);
or U10173 (N_10173,N_8427,N_7887);
nand U10174 (N_10174,N_6803,N_6412);
or U10175 (N_10175,N_8688,N_6628);
xnor U10176 (N_10176,N_6698,N_8752);
nand U10177 (N_10177,N_6672,N_8690);
nand U10178 (N_10178,N_8753,N_8049);
and U10179 (N_10179,N_7526,N_7981);
nor U10180 (N_10180,N_8866,N_7286);
nand U10181 (N_10181,N_8428,N_8894);
xor U10182 (N_10182,N_6306,N_7724);
nor U10183 (N_10183,N_7844,N_9320);
and U10184 (N_10184,N_6963,N_7077);
and U10185 (N_10185,N_6954,N_6893);
nor U10186 (N_10186,N_7133,N_8627);
or U10187 (N_10187,N_9105,N_6301);
nor U10188 (N_10188,N_9334,N_8217);
and U10189 (N_10189,N_7542,N_6823);
xnor U10190 (N_10190,N_7266,N_9161);
or U10191 (N_10191,N_7982,N_7362);
nand U10192 (N_10192,N_7538,N_6741);
or U10193 (N_10193,N_7104,N_7708);
xnor U10194 (N_10194,N_6524,N_8109);
nand U10195 (N_10195,N_8294,N_6481);
and U10196 (N_10196,N_8452,N_6796);
nand U10197 (N_10197,N_7922,N_6320);
nand U10198 (N_10198,N_8606,N_7840);
or U10199 (N_10199,N_9125,N_7245);
and U10200 (N_10200,N_7608,N_6589);
xnor U10201 (N_10201,N_7312,N_7644);
or U10202 (N_10202,N_7564,N_8169);
nor U10203 (N_10203,N_8916,N_8857);
and U10204 (N_10204,N_9354,N_7111);
xor U10205 (N_10205,N_9225,N_6880);
and U10206 (N_10206,N_8337,N_8142);
or U10207 (N_10207,N_6581,N_6550);
nand U10208 (N_10208,N_7094,N_6566);
nand U10209 (N_10209,N_8331,N_6895);
xor U10210 (N_10210,N_7184,N_7926);
or U10211 (N_10211,N_8576,N_6894);
nor U10212 (N_10212,N_8252,N_9252);
and U10213 (N_10213,N_9251,N_7047);
xor U10214 (N_10214,N_7415,N_7607);
nor U10215 (N_10215,N_6439,N_9023);
nor U10216 (N_10216,N_9065,N_7599);
nor U10217 (N_10217,N_6404,N_6634);
and U10218 (N_10218,N_6373,N_7731);
xor U10219 (N_10219,N_7452,N_8288);
and U10220 (N_10220,N_7778,N_6467);
xor U10221 (N_10221,N_7151,N_7495);
or U10222 (N_10222,N_8102,N_6795);
and U10223 (N_10223,N_9046,N_7250);
and U10224 (N_10224,N_8249,N_7138);
nor U10225 (N_10225,N_7001,N_9219);
nand U10226 (N_10226,N_6393,N_9075);
or U10227 (N_10227,N_7082,N_8547);
nand U10228 (N_10228,N_8361,N_6285);
or U10229 (N_10229,N_7249,N_9279);
nor U10230 (N_10230,N_6931,N_6526);
or U10231 (N_10231,N_7868,N_6488);
nor U10232 (N_10232,N_6487,N_7350);
and U10233 (N_10233,N_7514,N_8844);
nor U10234 (N_10234,N_6396,N_8830);
and U10235 (N_10235,N_8654,N_6263);
nand U10236 (N_10236,N_8122,N_6701);
xor U10237 (N_10237,N_8523,N_6758);
nand U10238 (N_10238,N_9002,N_8179);
nor U10239 (N_10239,N_7853,N_9202);
or U10240 (N_10240,N_9272,N_6417);
or U10241 (N_10241,N_8904,N_7827);
nand U10242 (N_10242,N_6773,N_8161);
nor U10243 (N_10243,N_9168,N_8000);
or U10244 (N_10244,N_6983,N_8038);
nand U10245 (N_10245,N_7164,N_7021);
nand U10246 (N_10246,N_7952,N_8927);
nand U10247 (N_10247,N_7852,N_6384);
nor U10248 (N_10248,N_6539,N_7462);
and U10249 (N_10249,N_7589,N_8490);
and U10250 (N_10250,N_8821,N_9096);
or U10251 (N_10251,N_7282,N_6677);
or U10252 (N_10252,N_6852,N_8032);
and U10253 (N_10253,N_7360,N_7258);
or U10254 (N_10254,N_6403,N_8871);
nand U10255 (N_10255,N_6600,N_9039);
xnor U10256 (N_10256,N_8887,N_6686);
nand U10257 (N_10257,N_9154,N_7873);
xnor U10258 (N_10258,N_8794,N_8255);
nor U10259 (N_10259,N_6958,N_7378);
nand U10260 (N_10260,N_8342,N_8980);
or U10261 (N_10261,N_7272,N_6940);
and U10262 (N_10262,N_6619,N_8808);
or U10263 (N_10263,N_7793,N_6724);
and U10264 (N_10264,N_7794,N_6438);
xnor U10265 (N_10265,N_7112,N_8242);
xnor U10266 (N_10266,N_8107,N_7811);
nor U10267 (N_10267,N_7642,N_8014);
and U10268 (N_10268,N_8940,N_6993);
xnor U10269 (N_10269,N_7730,N_6975);
or U10270 (N_10270,N_6763,N_8632);
and U10271 (N_10271,N_7041,N_7838);
nand U10272 (N_10272,N_6367,N_6446);
nand U10273 (N_10273,N_7560,N_6715);
or U10274 (N_10274,N_7785,N_8273);
or U10275 (N_10275,N_8671,N_6943);
nor U10276 (N_10276,N_9186,N_7786);
xor U10277 (N_10277,N_8237,N_9175);
nand U10278 (N_10278,N_9298,N_8809);
xor U10279 (N_10279,N_8908,N_6313);
or U10280 (N_10280,N_7624,N_9265);
and U10281 (N_10281,N_8103,N_7984);
xor U10282 (N_10282,N_8360,N_7662);
nand U10283 (N_10283,N_7195,N_8610);
nand U10284 (N_10284,N_9278,N_8512);
or U10285 (N_10285,N_6360,N_8388);
xor U10286 (N_10286,N_9033,N_6720);
nand U10287 (N_10287,N_6303,N_8902);
xnor U10288 (N_10288,N_8201,N_9127);
and U10289 (N_10289,N_8492,N_7583);
xnor U10290 (N_10290,N_6680,N_6837);
or U10291 (N_10291,N_9073,N_8497);
and U10292 (N_10292,N_7042,N_9352);
and U10293 (N_10293,N_6598,N_7269);
xor U10294 (N_10294,N_8735,N_8091);
and U10295 (N_10295,N_7630,N_6461);
or U10296 (N_10296,N_8491,N_9232);
xor U10297 (N_10297,N_9212,N_8818);
nand U10298 (N_10298,N_7375,N_7805);
xnor U10299 (N_10299,N_9109,N_8705);
and U10300 (N_10300,N_7758,N_7757);
xor U10301 (N_10301,N_6606,N_7436);
xor U10302 (N_10302,N_7916,N_6375);
and U10303 (N_10303,N_8153,N_7568);
or U10304 (N_10304,N_8144,N_8366);
or U10305 (N_10305,N_9034,N_7372);
or U10306 (N_10306,N_6679,N_7605);
and U10307 (N_10307,N_8325,N_6442);
nand U10308 (N_10308,N_7279,N_6546);
xor U10309 (N_10309,N_7625,N_9284);
nor U10310 (N_10310,N_6338,N_8529);
and U10311 (N_10311,N_9302,N_7037);
nand U10312 (N_10312,N_7674,N_6345);
nor U10313 (N_10313,N_8463,N_9043);
or U10314 (N_10314,N_9030,N_8947);
xnor U10315 (N_10315,N_9301,N_8377);
xor U10316 (N_10316,N_7054,N_7068);
nor U10317 (N_10317,N_6675,N_6908);
nand U10318 (N_10318,N_9220,N_8105);
nand U10319 (N_10319,N_8585,N_7823);
or U10320 (N_10320,N_6733,N_6575);
and U10321 (N_10321,N_8912,N_6407);
nor U10322 (N_10322,N_8660,N_7146);
and U10323 (N_10323,N_9255,N_8371);
nor U10324 (N_10324,N_8597,N_8996);
xor U10325 (N_10325,N_8573,N_8174);
nor U10326 (N_10326,N_9099,N_8539);
xor U10327 (N_10327,N_8222,N_8609);
nor U10328 (N_10328,N_6573,N_9319);
or U10329 (N_10329,N_8459,N_6542);
nor U10330 (N_10330,N_7732,N_8081);
and U10331 (N_10331,N_8613,N_7442);
nand U10332 (N_10332,N_7776,N_7431);
or U10333 (N_10333,N_6707,N_8763);
or U10334 (N_10334,N_6480,N_7134);
nand U10335 (N_10335,N_8268,N_6296);
or U10336 (N_10336,N_8999,N_7155);
or U10337 (N_10337,N_6537,N_6668);
xor U10338 (N_10338,N_7795,N_6437);
nand U10339 (N_10339,N_7847,N_9006);
or U10340 (N_10340,N_6572,N_9310);
nand U10341 (N_10341,N_8964,N_6380);
or U10342 (N_10342,N_6317,N_8603);
nand U10343 (N_10343,N_7492,N_7901);
and U10344 (N_10344,N_8193,N_8973);
xor U10345 (N_10345,N_8915,N_8015);
and U10346 (N_10346,N_6916,N_8430);
xor U10347 (N_10347,N_6413,N_8383);
nor U10348 (N_10348,N_9164,N_9216);
or U10349 (N_10349,N_8922,N_8748);
nor U10350 (N_10350,N_8343,N_8596);
nand U10351 (N_10351,N_9091,N_6647);
nor U10352 (N_10352,N_8775,N_6340);
xor U10353 (N_10353,N_7592,N_6906);
nor U10354 (N_10354,N_6732,N_6327);
xor U10355 (N_10355,N_6620,N_8791);
nor U10356 (N_10356,N_9335,N_8525);
nand U10357 (N_10357,N_6650,N_8684);
nor U10358 (N_10358,N_7913,N_7513);
nand U10359 (N_10359,N_9111,N_6476);
or U10360 (N_10360,N_8945,N_6844);
nor U10361 (N_10361,N_7772,N_7822);
xor U10362 (N_10362,N_7506,N_9346);
or U10363 (N_10363,N_8012,N_8328);
or U10364 (N_10364,N_7235,N_8995);
or U10365 (N_10365,N_9028,N_9245);
xnor U10366 (N_10366,N_7392,N_8375);
nor U10367 (N_10367,N_9360,N_7843);
or U10368 (N_10368,N_8990,N_7477);
xnor U10369 (N_10369,N_7216,N_9236);
or U10370 (N_10370,N_6840,N_6482);
and U10371 (N_10371,N_7406,N_6972);
nor U10372 (N_10372,N_8385,N_7052);
and U10373 (N_10373,N_8728,N_8345);
or U10374 (N_10374,N_8703,N_8303);
xnor U10375 (N_10375,N_8448,N_7093);
nor U10376 (N_10376,N_7210,N_6252);
nand U10377 (N_10377,N_7980,N_6801);
xnor U10378 (N_10378,N_6337,N_6491);
and U10379 (N_10379,N_9297,N_8820);
nor U10380 (N_10380,N_8120,N_6494);
and U10381 (N_10381,N_6322,N_7174);
xor U10382 (N_10382,N_7725,N_8415);
nand U10383 (N_10383,N_8836,N_9303);
xor U10384 (N_10384,N_6792,N_7365);
xor U10385 (N_10385,N_8405,N_8554);
xor U10386 (N_10386,N_9306,N_6904);
and U10387 (N_10387,N_8825,N_8056);
or U10388 (N_10388,N_8958,N_8401);
nand U10389 (N_10389,N_8954,N_8117);
nand U10390 (N_10390,N_6673,N_8150);
nand U10391 (N_10391,N_7558,N_9032);
or U10392 (N_10392,N_7479,N_9199);
nand U10393 (N_10393,N_7089,N_8438);
or U10394 (N_10394,N_8339,N_6996);
xor U10395 (N_10395,N_7595,N_9226);
or U10396 (N_10396,N_7278,N_6276);
xor U10397 (N_10397,N_6674,N_6315);
and U10398 (N_10398,N_6402,N_7369);
nor U10399 (N_10399,N_7486,N_6764);
and U10400 (N_10400,N_7314,N_9037);
or U10401 (N_10401,N_7414,N_9132);
and U10402 (N_10402,N_7511,N_7012);
or U10403 (N_10403,N_8079,N_7051);
and U10404 (N_10404,N_6290,N_9005);
or U10405 (N_10405,N_7529,N_6767);
or U10406 (N_10406,N_9077,N_7628);
or U10407 (N_10407,N_8367,N_8680);
or U10408 (N_10408,N_8307,N_6329);
nand U10409 (N_10409,N_8422,N_7784);
nand U10410 (N_10410,N_6279,N_9283);
nor U10411 (N_10411,N_7418,N_8968);
and U10412 (N_10412,N_7128,N_8048);
xor U10413 (N_10413,N_6353,N_6669);
xor U10414 (N_10414,N_8204,N_7575);
xor U10415 (N_10415,N_6784,N_6363);
or U10416 (N_10416,N_7122,N_7597);
or U10417 (N_10417,N_7505,N_7000);
and U10418 (N_10418,N_6770,N_9084);
or U10419 (N_10419,N_7745,N_7328);
and U10420 (N_10420,N_7606,N_8601);
or U10421 (N_10421,N_7333,N_7231);
and U10422 (N_10422,N_9253,N_6425);
nor U10423 (N_10423,N_8865,N_7288);
and U10424 (N_10424,N_7396,N_6469);
or U10425 (N_10425,N_7185,N_8574);
or U10426 (N_10426,N_7741,N_8315);
nor U10427 (N_10427,N_7125,N_7411);
and U10428 (N_10428,N_9051,N_7019);
xnor U10429 (N_10429,N_6443,N_8812);
xnor U10430 (N_10430,N_7920,N_8051);
and U10431 (N_10431,N_7071,N_8598);
and U10432 (N_10432,N_9373,N_8329);
and U10433 (N_10433,N_6670,N_7160);
and U10434 (N_10434,N_8106,N_6787);
nand U10435 (N_10435,N_7488,N_7352);
nor U10436 (N_10436,N_6416,N_6264);
nand U10437 (N_10437,N_8500,N_8659);
or U10438 (N_10438,N_8047,N_8392);
nor U10439 (N_10439,N_6493,N_7340);
and U10440 (N_10440,N_8935,N_8451);
nand U10441 (N_10441,N_8423,N_7586);
and U10442 (N_10442,N_8118,N_7412);
and U10443 (N_10443,N_7081,N_8197);
or U10444 (N_10444,N_8943,N_8248);
nand U10445 (N_10445,N_6294,N_6917);
and U10446 (N_10446,N_8455,N_8216);
nand U10447 (N_10447,N_8806,N_7957);
xnor U10448 (N_10448,N_9007,N_8528);
xor U10449 (N_10449,N_6753,N_8458);
nand U10450 (N_10450,N_7407,N_8332);
or U10451 (N_10451,N_8420,N_8302);
xor U10452 (N_10452,N_8069,N_7454);
and U10453 (N_10453,N_6769,N_7710);
xnor U10454 (N_10454,N_6790,N_8760);
or U10455 (N_10455,N_8473,N_6445);
or U10456 (N_10456,N_7073,N_8591);
nand U10457 (N_10457,N_8535,N_6448);
nor U10458 (N_10458,N_9047,N_8031);
or U10459 (N_10459,N_8998,N_7132);
nand U10460 (N_10460,N_8741,N_7869);
nor U10461 (N_10461,N_7254,N_8622);
and U10462 (N_10462,N_7969,N_6655);
nand U10463 (N_10463,N_7489,N_8020);
xnor U10464 (N_10464,N_8518,N_6858);
and U10465 (N_10465,N_7080,N_7067);
and U10466 (N_10466,N_9185,N_7148);
and U10467 (N_10467,N_8336,N_8461);
nor U10468 (N_10468,N_9370,N_9240);
nor U10469 (N_10469,N_7163,N_7010);
nor U10470 (N_10470,N_8909,N_8228);
nand U10471 (N_10471,N_7114,N_6258);
nor U10472 (N_10472,N_7677,N_6554);
xnor U10473 (N_10473,N_6618,N_7193);
nand U10474 (N_10474,N_7317,N_6705);
and U10475 (N_10475,N_6548,N_7015);
and U10476 (N_10476,N_8253,N_6984);
nor U10477 (N_10477,N_8425,N_8078);
nand U10478 (N_10478,N_8295,N_6311);
nor U10479 (N_10479,N_8855,N_8693);
nor U10480 (N_10480,N_8709,N_6652);
nor U10481 (N_10481,N_8233,N_7572);
nor U10482 (N_10482,N_7848,N_9221);
and U10483 (N_10483,N_8843,N_8066);
xor U10484 (N_10484,N_8800,N_6580);
and U10485 (N_10485,N_7790,N_7274);
nor U10486 (N_10486,N_9011,N_7280);
nor U10487 (N_10487,N_6257,N_6319);
and U10488 (N_10488,N_7639,N_7205);
xor U10489 (N_10489,N_8888,N_8309);
nand U10490 (N_10490,N_8043,N_7342);
xor U10491 (N_10491,N_6857,N_7994);
or U10492 (N_10492,N_8190,N_8084);
xor U10493 (N_10493,N_8941,N_8870);
xor U10494 (N_10494,N_9287,N_7469);
nor U10495 (N_10495,N_6359,N_8098);
and U10496 (N_10496,N_7950,N_8646);
xnor U10497 (N_10497,N_7078,N_6762);
nand U10498 (N_10498,N_8895,N_6623);
and U10499 (N_10499,N_7996,N_7371);
nand U10500 (N_10500,N_6912,N_7030);
xor U10501 (N_10501,N_9364,N_6747);
nor U10502 (N_10502,N_6805,N_6292);
nand U10503 (N_10503,N_8804,N_8623);
nand U10504 (N_10504,N_8449,N_6658);
or U10505 (N_10505,N_8897,N_8283);
nor U10506 (N_10506,N_6334,N_7165);
nand U10507 (N_10507,N_8245,N_9066);
nor U10508 (N_10508,N_6876,N_7029);
nor U10509 (N_10509,N_7536,N_8356);
or U10510 (N_10510,N_8431,N_6441);
and U10511 (N_10511,N_7472,N_8587);
nand U10512 (N_10512,N_8635,N_6431);
xnor U10513 (N_10513,N_8516,N_6945);
nand U10514 (N_10514,N_6870,N_6551);
nand U10515 (N_10515,N_8508,N_8546);
xnor U10516 (N_10516,N_9200,N_8058);
or U10517 (N_10517,N_7388,N_7774);
nand U10518 (N_10518,N_8370,N_6336);
or U10519 (N_10519,N_6251,N_8298);
or U10520 (N_10520,N_6936,N_8403);
nor U10521 (N_10521,N_7814,N_9178);
xnor U10522 (N_10522,N_7551,N_6305);
or U10523 (N_10523,N_6664,N_7649);
xnor U10524 (N_10524,N_8711,N_7738);
and U10525 (N_10525,N_8441,N_7678);
or U10526 (N_10526,N_7368,N_8380);
xor U10527 (N_10527,N_7036,N_8738);
nand U10528 (N_10528,N_7555,N_7821);
xor U10529 (N_10529,N_6644,N_8540);
nor U10530 (N_10530,N_6565,N_7815);
nor U10531 (N_10531,N_7232,N_8618);
nand U10532 (N_10532,N_8543,N_9000);
nand U10533 (N_10533,N_6843,N_8368);
or U10534 (N_10534,N_8551,N_7931);
or U10535 (N_10535,N_7709,N_6845);
xnor U10536 (N_10536,N_7689,N_7587);
nor U10537 (N_10537,N_8185,N_6485);
and U10538 (N_10538,N_6848,N_6985);
nor U10539 (N_10539,N_8402,N_6821);
nand U10540 (N_10540,N_6483,N_7227);
and U10541 (N_10541,N_7905,N_8891);
nand U10542 (N_10542,N_7872,N_6743);
nor U10543 (N_10543,N_6925,N_8395);
or U10544 (N_10544,N_7222,N_7355);
and U10545 (N_10545,N_7696,N_6587);
nand U10546 (N_10546,N_7032,N_6275);
and U10547 (N_10547,N_8824,N_6835);
nor U10548 (N_10548,N_6886,N_8975);
xnor U10549 (N_10549,N_7136,N_8983);
nor U10550 (N_10550,N_8593,N_7147);
xor U10551 (N_10551,N_8138,N_8702);
nand U10552 (N_10552,N_8981,N_6596);
nor U10553 (N_10553,N_8673,N_6868);
and U10554 (N_10554,N_8071,N_8531);
or U10555 (N_10555,N_9363,N_7177);
xnor U10556 (N_10556,N_9001,N_6682);
nor U10557 (N_10557,N_8496,N_8962);
or U10558 (N_10558,N_8064,N_9120);
and U10559 (N_10559,N_7009,N_8631);
and U10560 (N_10560,N_6341,N_6583);
xnor U10561 (N_10561,N_8877,N_8399);
xor U10562 (N_10562,N_6501,N_7244);
nor U10563 (N_10563,N_8191,N_7939);
or U10564 (N_10564,N_6804,N_8418);
or U10565 (N_10565,N_7862,N_8560);
nand U10566 (N_10566,N_8479,N_7283);
nor U10567 (N_10567,N_7215,N_8414);
and U10568 (N_10568,N_6830,N_8050);
xor U10569 (N_10569,N_8326,N_7457);
xor U10570 (N_10570,N_7968,N_7933);
and U10571 (N_10571,N_6255,N_7519);
xnor U10572 (N_10572,N_7598,N_7780);
or U10573 (N_10573,N_7117,N_7566);
or U10574 (N_10574,N_6899,N_6699);
and U10575 (N_10575,N_9247,N_7439);
and U10576 (N_10576,N_9167,N_9163);
nand U10577 (N_10577,N_6389,N_7140);
nand U10578 (N_10578,N_8126,N_7767);
nand U10579 (N_10579,N_6819,N_8849);
or U10580 (N_10580,N_7753,N_8521);
nand U10581 (N_10581,N_8765,N_8157);
and U10582 (N_10582,N_8992,N_8263);
nand U10583 (N_10583,N_8225,N_8876);
xnor U10584 (N_10584,N_7043,N_8759);
nor U10585 (N_10585,N_7460,N_6896);
or U10586 (N_10586,N_8159,N_6716);
nand U10587 (N_10587,N_7426,N_6865);
nor U10588 (N_10588,N_6498,N_7995);
nor U10589 (N_10589,N_7563,N_6933);
xor U10590 (N_10590,N_6625,N_7804);
and U10591 (N_10591,N_6274,N_8322);
and U10592 (N_10592,N_8129,N_6713);
and U10593 (N_10593,N_7591,N_9270);
nor U10594 (N_10594,N_7902,N_8394);
and U10595 (N_10595,N_7403,N_8406);
nand U10596 (N_10596,N_6463,N_8538);
nor U10597 (N_10597,N_6809,N_7494);
nand U10598 (N_10598,N_9093,N_6621);
nor U10599 (N_10599,N_6721,N_7183);
or U10600 (N_10600,N_6696,N_8130);
nor U10601 (N_10601,N_8306,N_7461);
nor U10602 (N_10602,N_6712,N_6547);
and U10603 (N_10603,N_9347,N_8158);
nor U10604 (N_10604,N_8230,N_6666);
nor U10605 (N_10605,N_6517,N_9143);
xor U10606 (N_10606,N_8599,N_8649);
nand U10607 (N_10607,N_8171,N_7909);
xnor U10608 (N_10608,N_6490,N_6653);
and U10609 (N_10609,N_7246,N_6704);
xnor U10610 (N_10610,N_8357,N_8971);
or U10611 (N_10611,N_6549,N_7171);
xnor U10612 (N_10612,N_8948,N_7220);
or U10613 (N_10613,N_8867,N_6951);
xnor U10614 (N_10614,N_8097,N_6881);
nand U10615 (N_10615,N_7166,N_9305);
nor U10616 (N_10616,N_6504,N_7841);
or U10617 (N_10617,N_6788,N_6678);
nor U10618 (N_10618,N_7819,N_7465);
xnor U10619 (N_10619,N_6998,N_7799);
nor U10620 (N_10620,N_7023,N_7482);
nand U10621 (N_10621,N_6571,N_7144);
nand U10622 (N_10622,N_8137,N_7782);
nor U10623 (N_10623,N_8231,N_9187);
xnor U10624 (N_10624,N_7856,N_7523);
nor U10625 (N_10625,N_8281,N_7303);
xnor U10626 (N_10626,N_7383,N_8717);
nand U10627 (N_10627,N_6736,N_6903);
xnor U10628 (N_10628,N_7885,N_7892);
and U10629 (N_10629,N_7203,N_8786);
nand U10630 (N_10630,N_6746,N_6751);
nand U10631 (N_10631,N_7014,N_7339);
xor U10632 (N_10632,N_7863,N_6793);
or U10633 (N_10633,N_6808,N_7652);
nand U10634 (N_10634,N_8447,N_9057);
and U10635 (N_10635,N_7559,N_9311);
xnor U10636 (N_10636,N_8926,N_8914);
nand U10637 (N_10637,N_8365,N_7287);
or U10638 (N_10638,N_9177,N_9266);
or U10639 (N_10639,N_7046,N_8040);
nor U10640 (N_10640,N_8027,N_7581);
nor U10641 (N_10641,N_6271,N_7801);
or U10642 (N_10642,N_7063,N_7961);
or U10643 (N_10643,N_7621,N_9330);
or U10644 (N_10644,N_8278,N_8699);
nand U10645 (N_10645,N_6414,N_8099);
or U10646 (N_10646,N_8177,N_6454);
or U10647 (N_10647,N_8400,N_6643);
nand U10648 (N_10648,N_8495,N_7061);
xor U10649 (N_10649,N_7797,N_6930);
and U10650 (N_10650,N_8592,N_7818);
nand U10651 (N_10651,N_8834,N_8778);
or U10652 (N_10652,N_7870,N_8924);
xor U10653 (N_10653,N_7137,N_7336);
nor U10654 (N_10654,N_6282,N_7493);
nor U10655 (N_10655,N_7588,N_9010);
xor U10656 (N_10656,N_8024,N_8008);
xor U10657 (N_10657,N_7602,N_7158);
xor U10658 (N_10658,N_8254,N_7540);
nor U10659 (N_10659,N_6966,N_8938);
xor U10660 (N_10660,N_7016,N_8453);
or U10661 (N_10661,N_8194,N_7685);
or U10662 (N_10662,N_7609,N_7567);
xnor U10663 (N_10663,N_6739,N_7003);
or U10664 (N_10664,N_7946,N_9098);
and U10665 (N_10665,N_8125,N_7130);
or U10666 (N_10666,N_7013,N_6661);
or U10667 (N_10667,N_6272,N_8304);
nand U10668 (N_10668,N_6986,N_6860);
xor U10669 (N_10669,N_6997,N_8080);
and U10670 (N_10670,N_8757,N_8856);
or U10671 (N_10671,N_6928,N_7655);
and U10672 (N_10672,N_8715,N_7993);
nand U10673 (N_10673,N_9045,N_9326);
and U10674 (N_10674,N_6421,N_8198);
xnor U10675 (N_10675,N_9145,N_8832);
or U10676 (N_10676,N_8737,N_7521);
or U10677 (N_10677,N_9085,N_8113);
xor U10678 (N_10678,N_8121,N_6510);
xnor U10679 (N_10679,N_7487,N_7299);
and U10680 (N_10680,N_7255,N_6328);
nor U10681 (N_10681,N_7399,N_9128);
nand U10682 (N_10682,N_8929,N_8732);
nor U10683 (N_10683,N_6838,N_9055);
nor U10684 (N_10684,N_7912,N_6615);
or U10685 (N_10685,N_8933,N_8628);
xor U10686 (N_10686,N_7825,N_7124);
or U10687 (N_10687,N_7270,N_8443);
nand U10688 (N_10688,N_8045,N_6706);
nand U10689 (N_10689,N_7302,N_7878);
nor U10690 (N_10690,N_7987,N_7325);
and U10691 (N_10691,N_6995,N_6999);
nand U10692 (N_10692,N_7247,N_6591);
nor U10693 (N_10693,N_7807,N_7760);
nor U10694 (N_10694,N_8389,N_8028);
and U10695 (N_10695,N_6314,N_6478);
and U10696 (N_10696,N_7791,N_6637);
or U10697 (N_10697,N_7119,N_8494);
xnor U10698 (N_10698,N_7206,N_8358);
and U10699 (N_10699,N_7305,N_6651);
xnor U10700 (N_10700,N_7481,N_7777);
xnor U10701 (N_10701,N_6734,N_6277);
nor U10702 (N_10702,N_6828,N_8713);
nand U10703 (N_10703,N_9094,N_6507);
and U10704 (N_10704,N_6534,N_7816);
nand U10705 (N_10705,N_8462,N_7024);
nand U10706 (N_10706,N_9160,N_6725);
and U10707 (N_10707,N_8187,N_6505);
or U10708 (N_10708,N_6878,N_7401);
nand U10709 (N_10709,N_8798,N_8982);
and U10710 (N_10710,N_9012,N_7977);
nor U10711 (N_10711,N_8141,N_7062);
and U10712 (N_10712,N_8162,N_6750);
or U10713 (N_10713,N_8661,N_8564);
or U10714 (N_10714,N_7601,N_7017);
nor U10715 (N_10715,N_6964,N_6976);
or U10716 (N_10716,N_6982,N_9172);
xor U10717 (N_10717,N_8240,N_8346);
nand U10718 (N_10718,N_8984,N_7327);
and U10719 (N_10719,N_7836,N_8267);
nand U10720 (N_10720,N_8464,N_7992);
nand U10721 (N_10721,N_7181,N_7508);
nor U10722 (N_10722,N_8369,N_6352);
nor U10723 (N_10723,N_7578,N_8875);
nand U10724 (N_10724,N_7716,N_7932);
xnor U10725 (N_10725,N_6411,N_8739);
nand U10726 (N_10726,N_8010,N_7087);
nand U10727 (N_10727,N_7712,N_6544);
and U10728 (N_10728,N_9231,N_6578);
and U10729 (N_10729,N_6960,N_8001);
nand U10730 (N_10730,N_8633,N_6433);
xnor U10731 (N_10731,N_7691,N_9201);
nand U10732 (N_10732,N_9366,N_6530);
xnor U10733 (N_10733,N_6934,N_6326);
or U10734 (N_10734,N_9369,N_7527);
nor U10735 (N_10735,N_8846,N_8300);
nand U10736 (N_10736,N_9316,N_8704);
and U10737 (N_10737,N_7364,N_8799);
and U10738 (N_10738,N_7237,N_6558);
nor U10739 (N_10739,N_7326,N_7211);
nand U10740 (N_10740,N_9150,N_8733);
or U10741 (N_10741,N_7867,N_7413);
nand U10742 (N_10742,N_7501,N_7733);
or U10743 (N_10743,N_7771,N_7304);
nor U10744 (N_10744,N_8220,N_9358);
or U10745 (N_10745,N_8156,N_6351);
or U10746 (N_10746,N_7097,N_7300);
and U10747 (N_10747,N_9060,N_6671);
and U10748 (N_10748,N_9329,N_6520);
or U10749 (N_10749,N_7387,N_9214);
or U10750 (N_10750,N_7640,N_8450);
nor U10751 (N_10751,N_8697,N_8967);
and U10752 (N_10752,N_8756,N_7743);
nor U10753 (N_10753,N_8110,N_7512);
nor U10754 (N_10754,N_8348,N_9365);
nand U10755 (N_10755,N_7397,N_7102);
xor U10756 (N_10756,N_6718,N_6869);
nand U10757 (N_10757,N_7504,N_7316);
xnor U10758 (N_10758,N_9234,N_6832);
xor U10759 (N_10759,N_8766,N_6529);
nor U10760 (N_10760,N_7358,N_8789);
nand U10761 (N_10761,N_8271,N_8827);
xor U10762 (N_10762,N_8726,N_7098);
and U10763 (N_10763,N_8612,N_6887);
or U10764 (N_10764,N_8501,N_6256);
nor U10765 (N_10765,N_6527,N_6781);
and U10766 (N_10766,N_6737,N_7162);
nand U10767 (N_10767,N_9288,N_8133);
or U10768 (N_10768,N_8936,N_7898);
and U10769 (N_10769,N_8151,N_9074);
xnor U10770 (N_10770,N_6900,N_8743);
nor U10771 (N_10771,N_6635,N_8520);
xnor U10772 (N_10772,N_8168,N_8858);
and U10773 (N_10773,N_6429,N_8398);
nor U10774 (N_10774,N_8354,N_8444);
nor U10775 (N_10775,N_8203,N_8379);
and U10776 (N_10776,N_7755,N_6863);
nor U10777 (N_10777,N_7941,N_6383);
nand U10778 (N_10778,N_8208,N_7737);
and U10779 (N_10779,N_8338,N_8570);
xor U10780 (N_10780,N_7240,N_6659);
or U10781 (N_10781,N_7849,N_8143);
nor U10782 (N_10782,N_6873,N_8669);
or U10783 (N_10783,N_8685,N_9102);
nand U10784 (N_10784,N_9371,N_8124);
nand U10785 (N_10785,N_6516,N_8289);
or U10786 (N_10786,N_6270,N_8731);
nand U10787 (N_10787,N_7736,N_6859);
xor U10788 (N_10788,N_6570,N_6729);
and U10789 (N_10789,N_7972,N_8465);
nand U10790 (N_10790,N_9345,N_7727);
xnor U10791 (N_10791,N_8460,N_8814);
nand U10792 (N_10792,N_8029,N_8436);
xnor U10793 (N_10793,N_8899,N_7152);
nand U10794 (N_10794,N_8155,N_8284);
and U10795 (N_10795,N_8076,N_9322);
xor U10796 (N_10796,N_9061,N_6727);
nand U10797 (N_10797,N_9193,N_7541);
xor U10798 (N_10798,N_8840,N_6923);
nand U10799 (N_10799,N_8542,N_7044);
or U10800 (N_10800,N_7105,N_8068);
nor U10801 (N_10801,N_7315,N_6604);
and U10802 (N_10802,N_8509,N_6836);
xnor U10803 (N_10803,N_7684,N_7306);
nand U10804 (N_10804,N_8355,N_7656);
and U10805 (N_10805,N_7991,N_6969);
xnor U10806 (N_10806,N_6645,N_7742);
nor U10807 (N_10807,N_6293,N_9135);
xnor U10808 (N_10808,N_9153,N_6594);
nand U10809 (N_10809,N_8647,N_7192);
or U10810 (N_10810,N_8959,N_8911);
nor U10811 (N_10811,N_8950,N_6901);
nor U10812 (N_10812,N_6616,N_8160);
xnor U10813 (N_10813,N_6730,N_7635);
and U10814 (N_10814,N_6640,N_8128);
nor U10815 (N_10815,N_7180,N_8095);
or U10816 (N_10816,N_6847,N_7927);
or U10817 (N_10817,N_6273,N_7653);
or U10818 (N_10818,N_8057,N_6752);
nor U10819 (N_10819,N_6888,N_8527);
or U10820 (N_10820,N_8862,N_8148);
xor U10821 (N_10821,N_9035,N_6723);
and U10822 (N_10822,N_9348,N_7025);
or U10823 (N_10823,N_6332,N_8588);
xnor U10824 (N_10824,N_8774,N_8869);
nor U10825 (N_10825,N_6757,N_8435);
or U10826 (N_10826,N_7391,N_9338);
nor U10827 (N_10827,N_8477,N_7263);
xor U10828 (N_10828,N_8966,N_8514);
nand U10829 (N_10829,N_8811,N_6829);
xnor U10830 (N_10830,N_7839,N_9230);
xnor U10831 (N_10831,N_6978,N_6789);
or U10832 (N_10832,N_7318,N_8002);
nor U10833 (N_10833,N_9155,N_7259);
nor U10834 (N_10834,N_7985,N_7748);
xor U10835 (N_10835,N_9003,N_8681);
and U10836 (N_10836,N_9237,N_9258);
xnor U10837 (N_10837,N_9299,N_8393);
and U10838 (N_10838,N_8993,N_8250);
xor U10839 (N_10839,N_9140,N_9342);
and U10840 (N_10840,N_8229,N_8556);
nor U10841 (N_10841,N_6374,N_6297);
or U10842 (N_10842,N_7175,N_6816);
and U10843 (N_10843,N_7202,N_7620);
nor U10844 (N_10844,N_7159,N_8575);
nand U10845 (N_10845,N_7615,N_8577);
and U10846 (N_10846,N_8210,N_8350);
and U10847 (N_10847,N_9263,N_9054);
nor U10848 (N_10848,N_6826,N_7522);
nand U10849 (N_10849,N_8147,N_8489);
xor U10850 (N_10850,N_6349,N_6423);
or U10851 (N_10851,N_7866,N_9318);
nand U10852 (N_10852,N_6387,N_9119);
xnor U10853 (N_10853,N_7033,N_8987);
nor U10854 (N_10854,N_6474,N_7936);
or U10855 (N_10855,N_9165,N_7139);
and U10856 (N_10856,N_8822,N_7106);
nor U10857 (N_10857,N_7516,N_7728);
nor U10858 (N_10858,N_6636,N_8689);
or U10859 (N_10859,N_6629,N_6974);
nor U10860 (N_10860,N_8282,N_8625);
or U10861 (N_10861,N_8017,N_7217);
xnor U10862 (N_10862,N_8182,N_7116);
nand U10863 (N_10863,N_8758,N_6324);
nand U10864 (N_10864,N_8648,N_7153);
or U10865 (N_10865,N_9213,N_7510);
xor U10866 (N_10866,N_6853,N_8183);
or U10867 (N_10867,N_6898,N_7672);
and U10868 (N_10868,N_6531,N_6927);
or U10869 (N_10869,N_6814,N_7188);
nor U10870 (N_10870,N_6511,N_6676);
xor U10871 (N_10871,N_6362,N_7301);
nor U10872 (N_10872,N_7877,N_9227);
and U10873 (N_10873,N_7053,N_6392);
xnor U10874 (N_10874,N_8562,N_8937);
xor U10875 (N_10875,N_8691,N_8767);
nand U10876 (N_10876,N_6667,N_8055);
xnor U10877 (N_10877,N_6710,N_9053);
nor U10878 (N_10878,N_8111,N_8771);
nand U10879 (N_10879,N_7545,N_8979);
nor U10880 (N_10880,N_7660,N_7792);
and U10881 (N_10881,N_9344,N_7747);
nor U10882 (N_10882,N_6765,N_8034);
nand U10883 (N_10883,N_7334,N_8226);
or U10884 (N_10884,N_7754,N_8257);
and U10885 (N_10885,N_8544,N_8042);
xor U10886 (N_10886,N_7404,N_6841);
nand U10887 (N_10887,N_6649,N_6973);
or U10888 (N_10888,N_7410,N_6522);
or U10889 (N_10889,N_8712,N_7610);
nand U10890 (N_10890,N_7858,N_8749);
nand U10891 (N_10891,N_6641,N_7879);
xnor U10892 (N_10892,N_8114,N_8662);
or U10893 (N_10893,N_7530,N_7900);
xnor U10894 (N_10894,N_7402,N_7248);
and U10895 (N_10895,N_6806,N_8239);
xor U10896 (N_10896,N_6378,N_7692);
or U10897 (N_10897,N_7173,N_9131);
and U10898 (N_10898,N_7975,N_7187);
xnor U10899 (N_10899,N_6890,N_6398);
and U10900 (N_10900,N_9118,N_7281);
nand U10901 (N_10901,N_8831,N_9123);
nor U10902 (N_10902,N_7855,N_8868);
and U10903 (N_10903,N_7895,N_8722);
or U10904 (N_10904,N_8212,N_7762);
and U10905 (N_10905,N_7343,N_6745);
xnor U10906 (N_10906,N_8653,N_6453);
nor U10907 (N_10907,N_7264,N_8708);
xor U10908 (N_10908,N_9250,N_6347);
nand U10909 (N_10909,N_9191,N_7798);
or U10910 (N_10910,N_8974,N_7473);
xor U10911 (N_10911,N_7459,N_8132);
nor U10912 (N_10912,N_6915,N_7467);
or U10913 (N_10913,N_8238,N_9218);
nand U10914 (N_10914,N_7810,N_6862);
or U10915 (N_10915,N_8502,N_9144);
xnor U10916 (N_10916,N_6503,N_8636);
or U10917 (N_10917,N_7917,N_6728);
xnor U10918 (N_10918,N_7056,N_6883);
nand U10919 (N_10919,N_9336,N_8433);
xor U10920 (N_10920,N_7428,N_8482);
nand U10921 (N_10921,N_7045,N_8039);
nand U10922 (N_10922,N_6420,N_7196);
or U10923 (N_10923,N_9181,N_8005);
nand U10924 (N_10924,N_6811,N_8426);
and U10925 (N_10925,N_6632,N_9203);
and U10926 (N_10926,N_8611,N_8769);
xor U10927 (N_10927,N_7703,N_7690);
or U10928 (N_10928,N_9101,N_8764);
xor U10929 (N_10929,N_8145,N_8803);
nor U10930 (N_10930,N_7156,N_7959);
and U10931 (N_10931,N_6657,N_8815);
nor U10932 (N_10932,N_6302,N_9049);
xnor U10933 (N_10933,N_8146,N_8290);
nand U10934 (N_10934,N_9188,N_8561);
nor U10935 (N_10935,N_9052,N_6564);
xor U10936 (N_10936,N_8892,N_8720);
nor U10937 (N_10937,N_7338,N_6259);
nand U10938 (N_10938,N_9208,N_6939);
and U10939 (N_10939,N_6934,N_8240);
and U10940 (N_10940,N_9140,N_8371);
and U10941 (N_10941,N_6808,N_7504);
or U10942 (N_10942,N_7973,N_8607);
and U10943 (N_10943,N_6819,N_7792);
and U10944 (N_10944,N_8864,N_7060);
or U10945 (N_10945,N_9352,N_7017);
or U10946 (N_10946,N_8758,N_6315);
or U10947 (N_10947,N_6812,N_8807);
nor U10948 (N_10948,N_8307,N_7002);
nand U10949 (N_10949,N_7805,N_7027);
and U10950 (N_10950,N_7702,N_9186);
and U10951 (N_10951,N_6750,N_6770);
nor U10952 (N_10952,N_6496,N_9293);
and U10953 (N_10953,N_7409,N_8553);
xor U10954 (N_10954,N_7034,N_6695);
and U10955 (N_10955,N_8131,N_6389);
and U10956 (N_10956,N_6325,N_9346);
nor U10957 (N_10957,N_7873,N_6894);
and U10958 (N_10958,N_9238,N_9190);
nor U10959 (N_10959,N_6498,N_6432);
and U10960 (N_10960,N_8476,N_8087);
or U10961 (N_10961,N_7754,N_7072);
nor U10962 (N_10962,N_7263,N_7302);
nand U10963 (N_10963,N_9374,N_8220);
xor U10964 (N_10964,N_8619,N_8495);
nor U10965 (N_10965,N_8191,N_8445);
and U10966 (N_10966,N_7773,N_6885);
or U10967 (N_10967,N_6923,N_9016);
xnor U10968 (N_10968,N_7067,N_7782);
and U10969 (N_10969,N_8015,N_7676);
or U10970 (N_10970,N_8910,N_9205);
nand U10971 (N_10971,N_8924,N_9174);
nand U10972 (N_10972,N_6745,N_8981);
or U10973 (N_10973,N_9041,N_6778);
nand U10974 (N_10974,N_9137,N_7424);
nor U10975 (N_10975,N_8508,N_9283);
or U10976 (N_10976,N_7359,N_7101);
xor U10977 (N_10977,N_7963,N_8503);
or U10978 (N_10978,N_7158,N_9246);
or U10979 (N_10979,N_9328,N_6900);
nand U10980 (N_10980,N_7289,N_7288);
nand U10981 (N_10981,N_8662,N_7971);
xnor U10982 (N_10982,N_6779,N_9073);
nor U10983 (N_10983,N_8583,N_6836);
nand U10984 (N_10984,N_6687,N_7306);
nor U10985 (N_10985,N_7069,N_8098);
nor U10986 (N_10986,N_6493,N_8017);
xor U10987 (N_10987,N_6864,N_7938);
or U10988 (N_10988,N_7295,N_7934);
and U10989 (N_10989,N_6595,N_7826);
nor U10990 (N_10990,N_6976,N_8899);
and U10991 (N_10991,N_6624,N_9160);
nand U10992 (N_10992,N_8720,N_7433);
or U10993 (N_10993,N_6286,N_7474);
nor U10994 (N_10994,N_7764,N_7911);
nor U10995 (N_10995,N_8362,N_7962);
xnor U10996 (N_10996,N_7593,N_8132);
nor U10997 (N_10997,N_6747,N_7763);
nand U10998 (N_10998,N_8529,N_8028);
nand U10999 (N_10999,N_7587,N_7680);
xnor U11000 (N_11000,N_9360,N_6336);
xor U11001 (N_11001,N_6364,N_7786);
xor U11002 (N_11002,N_9074,N_9336);
xor U11003 (N_11003,N_6546,N_7206);
nand U11004 (N_11004,N_8461,N_7007);
and U11005 (N_11005,N_8618,N_6959);
or U11006 (N_11006,N_7571,N_8479);
and U11007 (N_11007,N_6738,N_8630);
xnor U11008 (N_11008,N_8113,N_6856);
nand U11009 (N_11009,N_7603,N_6895);
or U11010 (N_11010,N_9014,N_8097);
or U11011 (N_11011,N_6968,N_8904);
or U11012 (N_11012,N_6918,N_7618);
nand U11013 (N_11013,N_8860,N_7427);
xor U11014 (N_11014,N_9009,N_8333);
and U11015 (N_11015,N_6739,N_7939);
xnor U11016 (N_11016,N_9004,N_7654);
or U11017 (N_11017,N_7888,N_8591);
xor U11018 (N_11018,N_8255,N_6887);
nand U11019 (N_11019,N_8522,N_9284);
nor U11020 (N_11020,N_8476,N_7278);
xor U11021 (N_11021,N_6433,N_7752);
or U11022 (N_11022,N_9189,N_8616);
xnor U11023 (N_11023,N_7625,N_9172);
xor U11024 (N_11024,N_7609,N_9188);
xnor U11025 (N_11025,N_7722,N_9343);
xnor U11026 (N_11026,N_6959,N_7154);
xor U11027 (N_11027,N_6812,N_8607);
or U11028 (N_11028,N_7002,N_8572);
or U11029 (N_11029,N_8721,N_7711);
and U11030 (N_11030,N_6434,N_7798);
xor U11031 (N_11031,N_8424,N_7406);
or U11032 (N_11032,N_8724,N_7819);
xnor U11033 (N_11033,N_8199,N_8464);
xor U11034 (N_11034,N_6801,N_9057);
nor U11035 (N_11035,N_8236,N_7732);
nor U11036 (N_11036,N_7463,N_9154);
nand U11037 (N_11037,N_8685,N_6921);
nand U11038 (N_11038,N_8773,N_7238);
xor U11039 (N_11039,N_8550,N_6780);
or U11040 (N_11040,N_7093,N_9222);
and U11041 (N_11041,N_9219,N_8356);
and U11042 (N_11042,N_6354,N_6424);
or U11043 (N_11043,N_8679,N_7078);
and U11044 (N_11044,N_6867,N_7194);
xor U11045 (N_11045,N_6652,N_7306);
nor U11046 (N_11046,N_8459,N_7317);
xor U11047 (N_11047,N_7138,N_7936);
xnor U11048 (N_11048,N_8873,N_7705);
and U11049 (N_11049,N_8296,N_8458);
xnor U11050 (N_11050,N_7933,N_7902);
nor U11051 (N_11051,N_8885,N_8092);
or U11052 (N_11052,N_6336,N_8376);
or U11053 (N_11053,N_7635,N_8925);
xnor U11054 (N_11054,N_9175,N_6644);
nor U11055 (N_11055,N_9370,N_8730);
or U11056 (N_11056,N_6777,N_7169);
nand U11057 (N_11057,N_6319,N_6777);
and U11058 (N_11058,N_8558,N_8867);
nor U11059 (N_11059,N_7066,N_8834);
or U11060 (N_11060,N_7411,N_8642);
xnor U11061 (N_11061,N_9112,N_8527);
or U11062 (N_11062,N_7485,N_8606);
nor U11063 (N_11063,N_8664,N_6575);
nor U11064 (N_11064,N_7703,N_8782);
xor U11065 (N_11065,N_9040,N_8056);
or U11066 (N_11066,N_6674,N_7270);
nand U11067 (N_11067,N_6372,N_8214);
nor U11068 (N_11068,N_8884,N_8409);
and U11069 (N_11069,N_8195,N_6517);
xor U11070 (N_11070,N_6897,N_6474);
nand U11071 (N_11071,N_8294,N_8154);
and U11072 (N_11072,N_8230,N_7178);
nor U11073 (N_11073,N_6923,N_6897);
nor U11074 (N_11074,N_8316,N_8172);
xor U11075 (N_11075,N_7416,N_6939);
xor U11076 (N_11076,N_7142,N_7181);
and U11077 (N_11077,N_7987,N_8416);
xor U11078 (N_11078,N_7649,N_6869);
nor U11079 (N_11079,N_6768,N_8510);
or U11080 (N_11080,N_8721,N_8675);
or U11081 (N_11081,N_8880,N_8782);
nand U11082 (N_11082,N_6945,N_8411);
or U11083 (N_11083,N_9063,N_8281);
and U11084 (N_11084,N_6889,N_6973);
xnor U11085 (N_11085,N_9181,N_6610);
nor U11086 (N_11086,N_7883,N_6473);
or U11087 (N_11087,N_8464,N_8072);
nor U11088 (N_11088,N_8112,N_7249);
and U11089 (N_11089,N_8332,N_6561);
or U11090 (N_11090,N_7415,N_8229);
nand U11091 (N_11091,N_8699,N_6325);
nand U11092 (N_11092,N_8196,N_8882);
and U11093 (N_11093,N_7076,N_8153);
or U11094 (N_11094,N_6282,N_6830);
and U11095 (N_11095,N_8491,N_9063);
xor U11096 (N_11096,N_6369,N_8433);
nand U11097 (N_11097,N_7587,N_7179);
and U11098 (N_11098,N_6618,N_9218);
nor U11099 (N_11099,N_9097,N_7501);
xor U11100 (N_11100,N_8742,N_8930);
nor U11101 (N_11101,N_9282,N_6984);
nor U11102 (N_11102,N_8534,N_8559);
nor U11103 (N_11103,N_8119,N_7740);
or U11104 (N_11104,N_8660,N_8511);
or U11105 (N_11105,N_7594,N_6865);
nand U11106 (N_11106,N_7273,N_6710);
nor U11107 (N_11107,N_6385,N_8753);
or U11108 (N_11108,N_6370,N_6921);
nor U11109 (N_11109,N_8363,N_8815);
nor U11110 (N_11110,N_7611,N_7104);
nand U11111 (N_11111,N_8196,N_8018);
xnor U11112 (N_11112,N_8149,N_6337);
and U11113 (N_11113,N_8382,N_7316);
nand U11114 (N_11114,N_8478,N_7227);
nand U11115 (N_11115,N_8409,N_6484);
nand U11116 (N_11116,N_7366,N_7084);
or U11117 (N_11117,N_9116,N_6572);
and U11118 (N_11118,N_6518,N_7266);
nand U11119 (N_11119,N_6940,N_8061);
or U11120 (N_11120,N_7918,N_6887);
nor U11121 (N_11121,N_8049,N_8793);
xor U11122 (N_11122,N_7768,N_6895);
nand U11123 (N_11123,N_9095,N_8501);
or U11124 (N_11124,N_7035,N_8487);
and U11125 (N_11125,N_8502,N_6576);
xor U11126 (N_11126,N_9103,N_7199);
nand U11127 (N_11127,N_6399,N_6783);
nand U11128 (N_11128,N_8433,N_7491);
xor U11129 (N_11129,N_8123,N_6714);
nor U11130 (N_11130,N_8250,N_8677);
xnor U11131 (N_11131,N_7703,N_7926);
nor U11132 (N_11132,N_8465,N_8157);
nand U11133 (N_11133,N_8191,N_7734);
or U11134 (N_11134,N_9148,N_7909);
nand U11135 (N_11135,N_7723,N_7783);
nand U11136 (N_11136,N_6462,N_8717);
or U11137 (N_11137,N_9349,N_6337);
nand U11138 (N_11138,N_6447,N_8085);
xnor U11139 (N_11139,N_6556,N_7902);
and U11140 (N_11140,N_7582,N_6857);
xor U11141 (N_11141,N_6732,N_6952);
xnor U11142 (N_11142,N_8455,N_7877);
nand U11143 (N_11143,N_7832,N_7352);
nand U11144 (N_11144,N_7517,N_8413);
xnor U11145 (N_11145,N_7267,N_7235);
nor U11146 (N_11146,N_9259,N_7665);
nand U11147 (N_11147,N_9266,N_7605);
and U11148 (N_11148,N_8612,N_6328);
nor U11149 (N_11149,N_8053,N_6584);
xnor U11150 (N_11150,N_8842,N_8423);
xnor U11151 (N_11151,N_6373,N_7792);
or U11152 (N_11152,N_7062,N_7414);
nand U11153 (N_11153,N_9084,N_9357);
and U11154 (N_11154,N_7813,N_7263);
or U11155 (N_11155,N_8792,N_6599);
nand U11156 (N_11156,N_8766,N_9189);
or U11157 (N_11157,N_9225,N_8424);
or U11158 (N_11158,N_9351,N_7960);
or U11159 (N_11159,N_9326,N_9124);
or U11160 (N_11160,N_8480,N_8835);
nand U11161 (N_11161,N_7605,N_8626);
nor U11162 (N_11162,N_7499,N_8744);
and U11163 (N_11163,N_8346,N_6535);
and U11164 (N_11164,N_6270,N_6821);
or U11165 (N_11165,N_6553,N_8481);
nor U11166 (N_11166,N_8288,N_7890);
and U11167 (N_11167,N_8689,N_7113);
and U11168 (N_11168,N_6619,N_8886);
or U11169 (N_11169,N_8067,N_8545);
nand U11170 (N_11170,N_7410,N_7308);
or U11171 (N_11171,N_7692,N_7072);
and U11172 (N_11172,N_6789,N_7116);
xor U11173 (N_11173,N_6596,N_8164);
xnor U11174 (N_11174,N_8431,N_6646);
nor U11175 (N_11175,N_7149,N_7872);
xor U11176 (N_11176,N_8921,N_8251);
nor U11177 (N_11177,N_7426,N_8085);
and U11178 (N_11178,N_8139,N_6702);
nor U11179 (N_11179,N_9230,N_9227);
or U11180 (N_11180,N_8144,N_8719);
and U11181 (N_11181,N_8414,N_8172);
xor U11182 (N_11182,N_7606,N_8235);
or U11183 (N_11183,N_8917,N_8003);
or U11184 (N_11184,N_6653,N_8069);
xor U11185 (N_11185,N_6306,N_9284);
or U11186 (N_11186,N_8199,N_7756);
nand U11187 (N_11187,N_8767,N_6301);
xnor U11188 (N_11188,N_6286,N_6534);
or U11189 (N_11189,N_6901,N_6271);
and U11190 (N_11190,N_7079,N_6524);
nor U11191 (N_11191,N_7715,N_6734);
xnor U11192 (N_11192,N_7277,N_6448);
nor U11193 (N_11193,N_6395,N_8710);
nor U11194 (N_11194,N_6436,N_8084);
xor U11195 (N_11195,N_7740,N_7832);
or U11196 (N_11196,N_7590,N_8551);
nor U11197 (N_11197,N_8303,N_7040);
xor U11198 (N_11198,N_8369,N_7301);
xor U11199 (N_11199,N_6888,N_9361);
xor U11200 (N_11200,N_6748,N_6514);
xor U11201 (N_11201,N_8247,N_7983);
nor U11202 (N_11202,N_6942,N_8975);
xor U11203 (N_11203,N_8387,N_7958);
nor U11204 (N_11204,N_7914,N_7703);
nand U11205 (N_11205,N_8833,N_6471);
nand U11206 (N_11206,N_8198,N_7748);
nor U11207 (N_11207,N_7750,N_7947);
and U11208 (N_11208,N_7484,N_8216);
and U11209 (N_11209,N_7607,N_7501);
or U11210 (N_11210,N_7966,N_7738);
nand U11211 (N_11211,N_7262,N_8156);
and U11212 (N_11212,N_9330,N_9351);
xnor U11213 (N_11213,N_9114,N_6637);
or U11214 (N_11214,N_8152,N_8004);
or U11215 (N_11215,N_9348,N_7113);
nor U11216 (N_11216,N_6763,N_8649);
xor U11217 (N_11217,N_8333,N_8141);
xor U11218 (N_11218,N_9020,N_8711);
or U11219 (N_11219,N_6457,N_8441);
or U11220 (N_11220,N_8722,N_7275);
nor U11221 (N_11221,N_9233,N_7030);
nor U11222 (N_11222,N_6670,N_8361);
or U11223 (N_11223,N_7236,N_8259);
and U11224 (N_11224,N_6756,N_7284);
or U11225 (N_11225,N_8863,N_8578);
and U11226 (N_11226,N_7087,N_7783);
xor U11227 (N_11227,N_6888,N_6303);
or U11228 (N_11228,N_8140,N_8058);
nor U11229 (N_11229,N_6462,N_9167);
and U11230 (N_11230,N_9306,N_6479);
nand U11231 (N_11231,N_7578,N_6310);
xnor U11232 (N_11232,N_9306,N_7872);
or U11233 (N_11233,N_8598,N_8920);
nand U11234 (N_11234,N_6373,N_7183);
xnor U11235 (N_11235,N_9040,N_6584);
and U11236 (N_11236,N_6536,N_8795);
or U11237 (N_11237,N_8082,N_7195);
nor U11238 (N_11238,N_6757,N_8731);
or U11239 (N_11239,N_6839,N_8939);
nor U11240 (N_11240,N_6293,N_7840);
xnor U11241 (N_11241,N_6984,N_8757);
nor U11242 (N_11242,N_8387,N_7963);
and U11243 (N_11243,N_9104,N_8776);
xnor U11244 (N_11244,N_8535,N_8070);
or U11245 (N_11245,N_7623,N_7909);
or U11246 (N_11246,N_7557,N_7273);
and U11247 (N_11247,N_8537,N_7848);
or U11248 (N_11248,N_7720,N_7037);
nor U11249 (N_11249,N_7913,N_9061);
nand U11250 (N_11250,N_7475,N_9333);
or U11251 (N_11251,N_7280,N_6838);
nand U11252 (N_11252,N_8656,N_8275);
xnor U11253 (N_11253,N_8664,N_7764);
and U11254 (N_11254,N_7311,N_6956);
xnor U11255 (N_11255,N_7740,N_6753);
nor U11256 (N_11256,N_8502,N_6640);
and U11257 (N_11257,N_6718,N_6766);
and U11258 (N_11258,N_8130,N_9064);
xor U11259 (N_11259,N_8385,N_7359);
xor U11260 (N_11260,N_8052,N_6681);
nor U11261 (N_11261,N_7932,N_9133);
xnor U11262 (N_11262,N_6847,N_7459);
or U11263 (N_11263,N_8609,N_8637);
nor U11264 (N_11264,N_7977,N_6670);
or U11265 (N_11265,N_7350,N_6953);
or U11266 (N_11266,N_8688,N_8364);
and U11267 (N_11267,N_6981,N_7167);
or U11268 (N_11268,N_8274,N_8727);
or U11269 (N_11269,N_8011,N_8904);
and U11270 (N_11270,N_8974,N_8804);
nand U11271 (N_11271,N_7221,N_7346);
xnor U11272 (N_11272,N_8145,N_6442);
nand U11273 (N_11273,N_7279,N_8554);
and U11274 (N_11274,N_6607,N_7232);
or U11275 (N_11275,N_8235,N_9131);
and U11276 (N_11276,N_6456,N_8019);
or U11277 (N_11277,N_7559,N_6725);
nor U11278 (N_11278,N_8522,N_8008);
or U11279 (N_11279,N_6646,N_7370);
or U11280 (N_11280,N_6676,N_7771);
xor U11281 (N_11281,N_6524,N_8695);
nor U11282 (N_11282,N_6809,N_8506);
nor U11283 (N_11283,N_7350,N_7072);
nand U11284 (N_11284,N_7842,N_6508);
nand U11285 (N_11285,N_7255,N_7681);
xnor U11286 (N_11286,N_6679,N_8960);
nor U11287 (N_11287,N_8251,N_8769);
and U11288 (N_11288,N_8038,N_6332);
xor U11289 (N_11289,N_9299,N_6742);
xnor U11290 (N_11290,N_8559,N_7545);
or U11291 (N_11291,N_6279,N_7618);
or U11292 (N_11292,N_7459,N_9211);
xnor U11293 (N_11293,N_7010,N_9290);
nor U11294 (N_11294,N_8636,N_7879);
or U11295 (N_11295,N_6372,N_6442);
xor U11296 (N_11296,N_9053,N_8265);
nor U11297 (N_11297,N_8174,N_6791);
and U11298 (N_11298,N_8266,N_8526);
nor U11299 (N_11299,N_9328,N_8206);
nand U11300 (N_11300,N_9108,N_6326);
or U11301 (N_11301,N_6360,N_8989);
xnor U11302 (N_11302,N_6965,N_8202);
or U11303 (N_11303,N_8793,N_6698);
nand U11304 (N_11304,N_8890,N_9141);
and U11305 (N_11305,N_6339,N_8710);
nand U11306 (N_11306,N_7142,N_6946);
and U11307 (N_11307,N_7336,N_6941);
and U11308 (N_11308,N_9181,N_7362);
and U11309 (N_11309,N_6518,N_8249);
xor U11310 (N_11310,N_7654,N_8139);
and U11311 (N_11311,N_7754,N_8379);
and U11312 (N_11312,N_8089,N_7469);
nor U11313 (N_11313,N_8377,N_8931);
xnor U11314 (N_11314,N_6843,N_7221);
and U11315 (N_11315,N_9337,N_8499);
and U11316 (N_11316,N_6536,N_8010);
or U11317 (N_11317,N_7095,N_7647);
nor U11318 (N_11318,N_8568,N_9048);
nand U11319 (N_11319,N_6625,N_9355);
xnor U11320 (N_11320,N_7901,N_7603);
xor U11321 (N_11321,N_6869,N_7094);
and U11322 (N_11322,N_8089,N_8180);
or U11323 (N_11323,N_6556,N_8526);
and U11324 (N_11324,N_8101,N_8186);
nand U11325 (N_11325,N_8516,N_9255);
or U11326 (N_11326,N_6676,N_7984);
nor U11327 (N_11327,N_6562,N_7671);
or U11328 (N_11328,N_9003,N_7181);
or U11329 (N_11329,N_7200,N_7453);
and U11330 (N_11330,N_7771,N_6705);
xnor U11331 (N_11331,N_7196,N_6295);
xor U11332 (N_11332,N_6622,N_7144);
nor U11333 (N_11333,N_6640,N_7069);
nor U11334 (N_11334,N_8229,N_8230);
nor U11335 (N_11335,N_7053,N_6403);
and U11336 (N_11336,N_7564,N_7216);
nor U11337 (N_11337,N_7095,N_8593);
and U11338 (N_11338,N_9059,N_7383);
and U11339 (N_11339,N_8117,N_7681);
nor U11340 (N_11340,N_7599,N_8091);
nand U11341 (N_11341,N_8211,N_9242);
and U11342 (N_11342,N_6811,N_9121);
or U11343 (N_11343,N_8093,N_6395);
xnor U11344 (N_11344,N_7416,N_8462);
or U11345 (N_11345,N_8827,N_7830);
nand U11346 (N_11346,N_8323,N_8705);
xnor U11347 (N_11347,N_6736,N_8880);
or U11348 (N_11348,N_7562,N_7401);
or U11349 (N_11349,N_6716,N_7983);
or U11350 (N_11350,N_6988,N_9044);
and U11351 (N_11351,N_8666,N_8924);
nor U11352 (N_11352,N_6715,N_9022);
and U11353 (N_11353,N_8572,N_7768);
and U11354 (N_11354,N_6624,N_8054);
and U11355 (N_11355,N_7450,N_7133);
xor U11356 (N_11356,N_7395,N_6837);
and U11357 (N_11357,N_9067,N_7631);
and U11358 (N_11358,N_6827,N_9067);
or U11359 (N_11359,N_6479,N_7459);
nor U11360 (N_11360,N_6626,N_6716);
xnor U11361 (N_11361,N_8603,N_8343);
xnor U11362 (N_11362,N_8128,N_9002);
xnor U11363 (N_11363,N_8289,N_7691);
or U11364 (N_11364,N_7299,N_6599);
xor U11365 (N_11365,N_8502,N_6930);
nand U11366 (N_11366,N_6333,N_6986);
nor U11367 (N_11367,N_6494,N_8084);
nor U11368 (N_11368,N_8637,N_7489);
and U11369 (N_11369,N_7585,N_8524);
and U11370 (N_11370,N_7205,N_7891);
xor U11371 (N_11371,N_7608,N_6730);
nand U11372 (N_11372,N_7895,N_6971);
xnor U11373 (N_11373,N_7592,N_7292);
or U11374 (N_11374,N_6587,N_8660);
nand U11375 (N_11375,N_8691,N_6663);
or U11376 (N_11376,N_6882,N_8958);
nor U11377 (N_11377,N_8637,N_6853);
nor U11378 (N_11378,N_8983,N_8740);
and U11379 (N_11379,N_7414,N_8334);
nor U11380 (N_11380,N_8638,N_8202);
nor U11381 (N_11381,N_7691,N_7791);
nor U11382 (N_11382,N_6914,N_7374);
nor U11383 (N_11383,N_8237,N_6475);
and U11384 (N_11384,N_7518,N_8788);
nand U11385 (N_11385,N_7015,N_8163);
nand U11386 (N_11386,N_8588,N_6948);
nand U11387 (N_11387,N_6374,N_8917);
or U11388 (N_11388,N_6318,N_7834);
nand U11389 (N_11389,N_7296,N_7905);
or U11390 (N_11390,N_6428,N_7786);
nor U11391 (N_11391,N_8610,N_9209);
nor U11392 (N_11392,N_8241,N_7664);
xnor U11393 (N_11393,N_8145,N_7760);
or U11394 (N_11394,N_8891,N_7723);
nand U11395 (N_11395,N_8666,N_6504);
and U11396 (N_11396,N_8859,N_8127);
and U11397 (N_11397,N_8378,N_7733);
nor U11398 (N_11398,N_8593,N_8845);
or U11399 (N_11399,N_9032,N_6379);
nand U11400 (N_11400,N_8357,N_8906);
nand U11401 (N_11401,N_7326,N_8359);
nand U11402 (N_11402,N_6798,N_9210);
nand U11403 (N_11403,N_9124,N_8649);
and U11404 (N_11404,N_7682,N_8093);
or U11405 (N_11405,N_7160,N_9229);
and U11406 (N_11406,N_6664,N_8191);
nand U11407 (N_11407,N_8795,N_8102);
nor U11408 (N_11408,N_7369,N_8327);
nor U11409 (N_11409,N_8141,N_8318);
or U11410 (N_11410,N_8971,N_8290);
and U11411 (N_11411,N_8171,N_8758);
xnor U11412 (N_11412,N_7899,N_7758);
xor U11413 (N_11413,N_8479,N_7848);
or U11414 (N_11414,N_6395,N_8254);
nor U11415 (N_11415,N_6904,N_7392);
xnor U11416 (N_11416,N_8532,N_7497);
and U11417 (N_11417,N_7153,N_7522);
nand U11418 (N_11418,N_7363,N_7290);
or U11419 (N_11419,N_9359,N_6733);
or U11420 (N_11420,N_7577,N_6407);
xor U11421 (N_11421,N_8086,N_8337);
xnor U11422 (N_11422,N_6959,N_8983);
xor U11423 (N_11423,N_8169,N_7231);
or U11424 (N_11424,N_6968,N_7773);
and U11425 (N_11425,N_8280,N_6950);
nand U11426 (N_11426,N_9179,N_7166);
xor U11427 (N_11427,N_7235,N_6970);
nor U11428 (N_11428,N_6384,N_7552);
nand U11429 (N_11429,N_7385,N_8274);
and U11430 (N_11430,N_8755,N_8525);
and U11431 (N_11431,N_8662,N_7842);
nand U11432 (N_11432,N_6924,N_9167);
and U11433 (N_11433,N_8315,N_7023);
or U11434 (N_11434,N_7564,N_7578);
nand U11435 (N_11435,N_8325,N_9366);
nand U11436 (N_11436,N_9333,N_8086);
or U11437 (N_11437,N_9340,N_8881);
and U11438 (N_11438,N_7426,N_7801);
or U11439 (N_11439,N_8267,N_9157);
xnor U11440 (N_11440,N_7553,N_7941);
or U11441 (N_11441,N_7741,N_8627);
or U11442 (N_11442,N_7972,N_8521);
nor U11443 (N_11443,N_8089,N_7594);
nor U11444 (N_11444,N_8243,N_8693);
or U11445 (N_11445,N_6796,N_7357);
nand U11446 (N_11446,N_6341,N_8528);
nand U11447 (N_11447,N_6466,N_8570);
or U11448 (N_11448,N_7982,N_8433);
and U11449 (N_11449,N_9035,N_6413);
nor U11450 (N_11450,N_6895,N_8750);
and U11451 (N_11451,N_7863,N_6292);
nor U11452 (N_11452,N_6667,N_7135);
nand U11453 (N_11453,N_7452,N_8691);
nor U11454 (N_11454,N_6914,N_8053);
nor U11455 (N_11455,N_6664,N_6855);
or U11456 (N_11456,N_9052,N_7569);
nand U11457 (N_11457,N_6418,N_9212);
or U11458 (N_11458,N_8291,N_6308);
or U11459 (N_11459,N_8857,N_8145);
nand U11460 (N_11460,N_8863,N_7721);
and U11461 (N_11461,N_7769,N_8625);
nand U11462 (N_11462,N_8590,N_7812);
nand U11463 (N_11463,N_7128,N_6912);
nand U11464 (N_11464,N_6506,N_6579);
or U11465 (N_11465,N_7322,N_9105);
or U11466 (N_11466,N_6295,N_7935);
or U11467 (N_11467,N_8868,N_8048);
and U11468 (N_11468,N_8074,N_7184);
nor U11469 (N_11469,N_8974,N_8034);
nand U11470 (N_11470,N_7695,N_7776);
or U11471 (N_11471,N_8136,N_6550);
and U11472 (N_11472,N_8598,N_7942);
xnor U11473 (N_11473,N_7825,N_6667);
and U11474 (N_11474,N_8674,N_6489);
and U11475 (N_11475,N_7505,N_8764);
and U11476 (N_11476,N_8482,N_9289);
or U11477 (N_11477,N_8407,N_7725);
nand U11478 (N_11478,N_8155,N_8237);
and U11479 (N_11479,N_8433,N_7936);
xnor U11480 (N_11480,N_7464,N_8933);
nor U11481 (N_11481,N_7884,N_6857);
nor U11482 (N_11482,N_8379,N_6794);
or U11483 (N_11483,N_9323,N_6829);
xor U11484 (N_11484,N_7092,N_8332);
xnor U11485 (N_11485,N_9221,N_6838);
nor U11486 (N_11486,N_7839,N_6665);
and U11487 (N_11487,N_8536,N_8740);
and U11488 (N_11488,N_8405,N_7789);
or U11489 (N_11489,N_8441,N_8699);
nor U11490 (N_11490,N_8213,N_8889);
or U11491 (N_11491,N_7284,N_8478);
xor U11492 (N_11492,N_8870,N_6991);
xor U11493 (N_11493,N_7079,N_8976);
xor U11494 (N_11494,N_7163,N_8577);
xor U11495 (N_11495,N_8073,N_8636);
xor U11496 (N_11496,N_7076,N_6904);
nor U11497 (N_11497,N_8491,N_9292);
xor U11498 (N_11498,N_7472,N_7609);
xor U11499 (N_11499,N_8275,N_8976);
xnor U11500 (N_11500,N_7690,N_7844);
xnor U11501 (N_11501,N_8489,N_6453);
nor U11502 (N_11502,N_6923,N_6434);
nand U11503 (N_11503,N_7638,N_6277);
xnor U11504 (N_11504,N_8050,N_6999);
nand U11505 (N_11505,N_7136,N_8327);
or U11506 (N_11506,N_9237,N_8797);
xnor U11507 (N_11507,N_8983,N_8516);
nand U11508 (N_11508,N_8399,N_7948);
and U11509 (N_11509,N_6433,N_7455);
xor U11510 (N_11510,N_6863,N_9235);
nand U11511 (N_11511,N_8862,N_7223);
nand U11512 (N_11512,N_6942,N_6351);
or U11513 (N_11513,N_7151,N_8768);
nand U11514 (N_11514,N_7042,N_6391);
nand U11515 (N_11515,N_8299,N_9207);
or U11516 (N_11516,N_7095,N_6267);
xnor U11517 (N_11517,N_7628,N_8728);
xor U11518 (N_11518,N_7333,N_6571);
and U11519 (N_11519,N_6809,N_7046);
or U11520 (N_11520,N_8767,N_8806);
and U11521 (N_11521,N_7637,N_9132);
xor U11522 (N_11522,N_8783,N_8663);
xnor U11523 (N_11523,N_9207,N_8171);
nand U11524 (N_11524,N_6581,N_8560);
nand U11525 (N_11525,N_8506,N_9243);
and U11526 (N_11526,N_9061,N_8381);
nand U11527 (N_11527,N_7981,N_6373);
xor U11528 (N_11528,N_9151,N_8682);
xnor U11529 (N_11529,N_8004,N_7241);
nor U11530 (N_11530,N_9127,N_6823);
nand U11531 (N_11531,N_7134,N_7296);
and U11532 (N_11532,N_8417,N_8381);
nand U11533 (N_11533,N_7627,N_8734);
nor U11534 (N_11534,N_8434,N_8327);
nor U11535 (N_11535,N_6751,N_7366);
xnor U11536 (N_11536,N_7326,N_8235);
xor U11537 (N_11537,N_8680,N_8849);
and U11538 (N_11538,N_7753,N_6475);
and U11539 (N_11539,N_6687,N_7143);
nor U11540 (N_11540,N_7797,N_9291);
xnor U11541 (N_11541,N_7269,N_8458);
xnor U11542 (N_11542,N_6664,N_7623);
and U11543 (N_11543,N_7856,N_6616);
nor U11544 (N_11544,N_6478,N_8531);
xor U11545 (N_11545,N_7853,N_7386);
and U11546 (N_11546,N_8281,N_6495);
or U11547 (N_11547,N_9078,N_8642);
nor U11548 (N_11548,N_8156,N_7608);
xor U11549 (N_11549,N_6495,N_7347);
nand U11550 (N_11550,N_7240,N_7098);
and U11551 (N_11551,N_9373,N_7155);
nor U11552 (N_11552,N_6941,N_6982);
xor U11553 (N_11553,N_6406,N_8330);
nor U11554 (N_11554,N_8700,N_8766);
and U11555 (N_11555,N_8206,N_7299);
and U11556 (N_11556,N_9314,N_7457);
or U11557 (N_11557,N_8995,N_8596);
xor U11558 (N_11558,N_7602,N_7832);
nor U11559 (N_11559,N_7949,N_9279);
nor U11560 (N_11560,N_8743,N_8836);
or U11561 (N_11561,N_6460,N_6291);
xor U11562 (N_11562,N_6403,N_8716);
and U11563 (N_11563,N_7076,N_7236);
or U11564 (N_11564,N_7130,N_7430);
or U11565 (N_11565,N_6526,N_7652);
nor U11566 (N_11566,N_6477,N_8337);
or U11567 (N_11567,N_7255,N_7767);
or U11568 (N_11568,N_9309,N_9154);
or U11569 (N_11569,N_6423,N_6267);
or U11570 (N_11570,N_8573,N_9155);
xnor U11571 (N_11571,N_8889,N_7980);
and U11572 (N_11572,N_7397,N_7680);
nand U11573 (N_11573,N_6714,N_7292);
xnor U11574 (N_11574,N_9211,N_7404);
xor U11575 (N_11575,N_7049,N_6352);
and U11576 (N_11576,N_6259,N_6639);
or U11577 (N_11577,N_8141,N_7804);
or U11578 (N_11578,N_8619,N_9003);
and U11579 (N_11579,N_7788,N_8514);
nand U11580 (N_11580,N_6858,N_7626);
or U11581 (N_11581,N_7138,N_7509);
nor U11582 (N_11582,N_7039,N_6604);
nand U11583 (N_11583,N_9031,N_7318);
nand U11584 (N_11584,N_6851,N_7943);
or U11585 (N_11585,N_6685,N_8960);
and U11586 (N_11586,N_8949,N_6635);
xor U11587 (N_11587,N_7439,N_7128);
nand U11588 (N_11588,N_8367,N_9174);
nand U11589 (N_11589,N_6572,N_9001);
or U11590 (N_11590,N_7401,N_6799);
or U11591 (N_11591,N_9006,N_6816);
and U11592 (N_11592,N_7539,N_6882);
or U11593 (N_11593,N_8550,N_6608);
nand U11594 (N_11594,N_6730,N_9251);
nor U11595 (N_11595,N_7632,N_8515);
nor U11596 (N_11596,N_9132,N_9342);
or U11597 (N_11597,N_6279,N_8814);
and U11598 (N_11598,N_6294,N_8679);
or U11599 (N_11599,N_7332,N_9148);
and U11600 (N_11600,N_6891,N_9228);
or U11601 (N_11601,N_6878,N_7015);
xnor U11602 (N_11602,N_7926,N_6975);
nor U11603 (N_11603,N_9011,N_8866);
nor U11604 (N_11604,N_6287,N_8926);
nand U11605 (N_11605,N_6986,N_6270);
nand U11606 (N_11606,N_7929,N_7240);
nand U11607 (N_11607,N_7442,N_6613);
and U11608 (N_11608,N_8841,N_6778);
nor U11609 (N_11609,N_8299,N_6357);
nand U11610 (N_11610,N_8188,N_8101);
and U11611 (N_11611,N_8396,N_6614);
nor U11612 (N_11612,N_6278,N_7576);
nand U11613 (N_11613,N_7882,N_8510);
or U11614 (N_11614,N_7998,N_6917);
nor U11615 (N_11615,N_7411,N_7199);
or U11616 (N_11616,N_8143,N_7706);
nor U11617 (N_11617,N_9104,N_7607);
xor U11618 (N_11618,N_6350,N_6300);
and U11619 (N_11619,N_6559,N_7778);
and U11620 (N_11620,N_6791,N_7231);
nor U11621 (N_11621,N_8412,N_7327);
or U11622 (N_11622,N_6384,N_6345);
or U11623 (N_11623,N_6556,N_7037);
nor U11624 (N_11624,N_9159,N_6279);
nor U11625 (N_11625,N_9316,N_6268);
nor U11626 (N_11626,N_7882,N_8123);
nand U11627 (N_11627,N_8410,N_6679);
and U11628 (N_11628,N_8061,N_8806);
or U11629 (N_11629,N_6861,N_6322);
and U11630 (N_11630,N_8868,N_9199);
nand U11631 (N_11631,N_7344,N_7990);
nor U11632 (N_11632,N_9341,N_8737);
or U11633 (N_11633,N_6657,N_7274);
nand U11634 (N_11634,N_9219,N_8859);
and U11635 (N_11635,N_7373,N_9023);
nor U11636 (N_11636,N_8472,N_6580);
xor U11637 (N_11637,N_6600,N_8012);
and U11638 (N_11638,N_9283,N_6270);
and U11639 (N_11639,N_8247,N_9207);
xnor U11640 (N_11640,N_6667,N_8069);
nand U11641 (N_11641,N_8208,N_8217);
and U11642 (N_11642,N_6439,N_8321);
and U11643 (N_11643,N_7049,N_7111);
nor U11644 (N_11644,N_7958,N_7932);
xor U11645 (N_11645,N_6798,N_6404);
nand U11646 (N_11646,N_6769,N_8703);
xnor U11647 (N_11647,N_6446,N_8590);
or U11648 (N_11648,N_7215,N_8909);
xnor U11649 (N_11649,N_8627,N_8800);
nand U11650 (N_11650,N_6714,N_7184);
or U11651 (N_11651,N_7739,N_8004);
and U11652 (N_11652,N_8370,N_7539);
and U11653 (N_11653,N_9040,N_9110);
nor U11654 (N_11654,N_7897,N_6798);
nand U11655 (N_11655,N_6525,N_7079);
and U11656 (N_11656,N_9132,N_7436);
or U11657 (N_11657,N_8097,N_6526);
nor U11658 (N_11658,N_8773,N_8019);
nor U11659 (N_11659,N_8722,N_8317);
or U11660 (N_11660,N_6340,N_8340);
nor U11661 (N_11661,N_6688,N_9043);
and U11662 (N_11662,N_6884,N_9054);
xnor U11663 (N_11663,N_8856,N_7479);
and U11664 (N_11664,N_8014,N_7511);
nand U11665 (N_11665,N_8436,N_8324);
nor U11666 (N_11666,N_7584,N_7182);
or U11667 (N_11667,N_6317,N_7992);
or U11668 (N_11668,N_8824,N_6386);
nand U11669 (N_11669,N_6281,N_7340);
nor U11670 (N_11670,N_7315,N_8654);
or U11671 (N_11671,N_6321,N_6536);
nand U11672 (N_11672,N_7714,N_7089);
and U11673 (N_11673,N_6985,N_8284);
nand U11674 (N_11674,N_8434,N_8435);
and U11675 (N_11675,N_7749,N_7791);
nand U11676 (N_11676,N_6308,N_6938);
or U11677 (N_11677,N_8774,N_6443);
nor U11678 (N_11678,N_8321,N_7866);
nor U11679 (N_11679,N_6493,N_6507);
xor U11680 (N_11680,N_9160,N_6478);
and U11681 (N_11681,N_8369,N_8441);
xnor U11682 (N_11682,N_8623,N_8367);
nor U11683 (N_11683,N_9108,N_8999);
xor U11684 (N_11684,N_9357,N_8656);
and U11685 (N_11685,N_7939,N_8402);
nand U11686 (N_11686,N_8511,N_7133);
nand U11687 (N_11687,N_7426,N_8383);
or U11688 (N_11688,N_7682,N_6624);
or U11689 (N_11689,N_8178,N_8865);
xor U11690 (N_11690,N_6552,N_8567);
or U11691 (N_11691,N_9321,N_7801);
and U11692 (N_11692,N_8024,N_6424);
nand U11693 (N_11693,N_7542,N_9367);
and U11694 (N_11694,N_6774,N_7976);
or U11695 (N_11695,N_7737,N_7657);
nand U11696 (N_11696,N_6643,N_8666);
nor U11697 (N_11697,N_8519,N_7532);
and U11698 (N_11698,N_8197,N_8473);
or U11699 (N_11699,N_7012,N_7610);
nor U11700 (N_11700,N_8353,N_8222);
or U11701 (N_11701,N_7653,N_7397);
nor U11702 (N_11702,N_9004,N_8766);
nor U11703 (N_11703,N_6340,N_8037);
xnor U11704 (N_11704,N_6550,N_8638);
nand U11705 (N_11705,N_6877,N_8596);
xnor U11706 (N_11706,N_7465,N_6391);
and U11707 (N_11707,N_7695,N_8693);
and U11708 (N_11708,N_7458,N_7928);
and U11709 (N_11709,N_9307,N_7290);
and U11710 (N_11710,N_6932,N_7044);
xnor U11711 (N_11711,N_7674,N_6458);
nor U11712 (N_11712,N_7200,N_7975);
nand U11713 (N_11713,N_7803,N_8719);
nand U11714 (N_11714,N_6671,N_9200);
nor U11715 (N_11715,N_8769,N_6468);
and U11716 (N_11716,N_6706,N_8102);
nand U11717 (N_11717,N_9362,N_9165);
and U11718 (N_11718,N_9308,N_6358);
nor U11719 (N_11719,N_9086,N_8932);
nand U11720 (N_11720,N_6584,N_8923);
nor U11721 (N_11721,N_8182,N_8601);
and U11722 (N_11722,N_8532,N_6738);
nor U11723 (N_11723,N_7291,N_8946);
and U11724 (N_11724,N_8902,N_8745);
and U11725 (N_11725,N_8608,N_8717);
and U11726 (N_11726,N_8332,N_7593);
nor U11727 (N_11727,N_8411,N_6729);
nand U11728 (N_11728,N_9305,N_8979);
xnor U11729 (N_11729,N_6731,N_6687);
and U11730 (N_11730,N_8445,N_9298);
or U11731 (N_11731,N_7621,N_6444);
nand U11732 (N_11732,N_7438,N_6682);
nand U11733 (N_11733,N_7389,N_6633);
or U11734 (N_11734,N_6271,N_8380);
and U11735 (N_11735,N_6844,N_7471);
nand U11736 (N_11736,N_7419,N_8782);
and U11737 (N_11737,N_8076,N_7717);
nand U11738 (N_11738,N_6975,N_7816);
or U11739 (N_11739,N_6868,N_8291);
xnor U11740 (N_11740,N_8325,N_8667);
nand U11741 (N_11741,N_9185,N_9084);
or U11742 (N_11742,N_7533,N_6880);
and U11743 (N_11743,N_6720,N_6476);
or U11744 (N_11744,N_6917,N_6580);
xnor U11745 (N_11745,N_7385,N_9008);
xnor U11746 (N_11746,N_8713,N_7505);
nor U11747 (N_11747,N_8845,N_8802);
xnor U11748 (N_11748,N_7319,N_6486);
nor U11749 (N_11749,N_6974,N_7491);
and U11750 (N_11750,N_8408,N_7137);
and U11751 (N_11751,N_9237,N_9200);
or U11752 (N_11752,N_8394,N_6570);
xor U11753 (N_11753,N_6493,N_8056);
or U11754 (N_11754,N_9240,N_9295);
nor U11755 (N_11755,N_6279,N_7337);
or U11756 (N_11756,N_8076,N_8384);
and U11757 (N_11757,N_7171,N_8149);
and U11758 (N_11758,N_9194,N_7414);
nand U11759 (N_11759,N_7507,N_8824);
nand U11760 (N_11760,N_9307,N_6379);
nand U11761 (N_11761,N_7189,N_7202);
xnor U11762 (N_11762,N_8853,N_9023);
nor U11763 (N_11763,N_7980,N_9346);
nand U11764 (N_11764,N_6946,N_7520);
nor U11765 (N_11765,N_8095,N_6937);
nor U11766 (N_11766,N_7407,N_8512);
and U11767 (N_11767,N_8300,N_8209);
nor U11768 (N_11768,N_6601,N_8562);
or U11769 (N_11769,N_6766,N_6801);
xnor U11770 (N_11770,N_8582,N_6395);
and U11771 (N_11771,N_6542,N_7762);
and U11772 (N_11772,N_9312,N_8322);
nand U11773 (N_11773,N_7313,N_7515);
and U11774 (N_11774,N_7724,N_8816);
nor U11775 (N_11775,N_7414,N_6776);
nand U11776 (N_11776,N_7020,N_8555);
xor U11777 (N_11777,N_8352,N_7197);
and U11778 (N_11778,N_7871,N_7361);
nand U11779 (N_11779,N_8322,N_7672);
or U11780 (N_11780,N_7645,N_6979);
and U11781 (N_11781,N_7628,N_7789);
xnor U11782 (N_11782,N_8411,N_6705);
or U11783 (N_11783,N_9198,N_7853);
and U11784 (N_11784,N_7332,N_8156);
or U11785 (N_11785,N_7844,N_9352);
xnor U11786 (N_11786,N_8887,N_8798);
xor U11787 (N_11787,N_6715,N_8408);
nor U11788 (N_11788,N_8841,N_6264);
or U11789 (N_11789,N_6506,N_9070);
xnor U11790 (N_11790,N_7805,N_7209);
nor U11791 (N_11791,N_8568,N_7471);
nor U11792 (N_11792,N_8254,N_9161);
nor U11793 (N_11793,N_7132,N_8419);
or U11794 (N_11794,N_7398,N_8316);
or U11795 (N_11795,N_8267,N_7340);
or U11796 (N_11796,N_6953,N_8949);
xnor U11797 (N_11797,N_6461,N_7960);
nor U11798 (N_11798,N_6332,N_9253);
or U11799 (N_11799,N_6420,N_7656);
and U11800 (N_11800,N_8841,N_8329);
nand U11801 (N_11801,N_7910,N_7256);
nor U11802 (N_11802,N_6394,N_7336);
xor U11803 (N_11803,N_7207,N_8545);
and U11804 (N_11804,N_7545,N_9007);
or U11805 (N_11805,N_9060,N_6385);
nand U11806 (N_11806,N_9287,N_8925);
xor U11807 (N_11807,N_7996,N_8522);
or U11808 (N_11808,N_6603,N_6761);
xnor U11809 (N_11809,N_8813,N_9369);
nand U11810 (N_11810,N_8917,N_9287);
nand U11811 (N_11811,N_8621,N_6284);
and U11812 (N_11812,N_8114,N_9144);
nand U11813 (N_11813,N_7088,N_8050);
nand U11814 (N_11814,N_9128,N_6339);
nor U11815 (N_11815,N_6569,N_8035);
and U11816 (N_11816,N_6400,N_6688);
nor U11817 (N_11817,N_7297,N_9222);
nor U11818 (N_11818,N_7791,N_6974);
nor U11819 (N_11819,N_9137,N_9233);
nand U11820 (N_11820,N_7977,N_6646);
and U11821 (N_11821,N_6928,N_8545);
nor U11822 (N_11822,N_7784,N_8533);
xor U11823 (N_11823,N_6308,N_8141);
or U11824 (N_11824,N_6492,N_8688);
nand U11825 (N_11825,N_8545,N_6785);
nand U11826 (N_11826,N_6639,N_8167);
xnor U11827 (N_11827,N_6978,N_7075);
and U11828 (N_11828,N_8536,N_6609);
xnor U11829 (N_11829,N_6414,N_9155);
and U11830 (N_11830,N_7976,N_8384);
nor U11831 (N_11831,N_8970,N_7340);
nor U11832 (N_11832,N_8894,N_9058);
nor U11833 (N_11833,N_8862,N_9091);
xnor U11834 (N_11834,N_9318,N_7596);
and U11835 (N_11835,N_9343,N_7691);
nor U11836 (N_11836,N_8423,N_8379);
xor U11837 (N_11837,N_8492,N_6984);
xor U11838 (N_11838,N_8107,N_7538);
and U11839 (N_11839,N_9259,N_8083);
nor U11840 (N_11840,N_7631,N_8098);
nor U11841 (N_11841,N_9353,N_6351);
or U11842 (N_11842,N_7491,N_9063);
or U11843 (N_11843,N_6527,N_8964);
nand U11844 (N_11844,N_8759,N_6725);
nor U11845 (N_11845,N_9292,N_7598);
nor U11846 (N_11846,N_8328,N_6767);
xor U11847 (N_11847,N_6980,N_8480);
xnor U11848 (N_11848,N_7019,N_8548);
or U11849 (N_11849,N_9220,N_7800);
xor U11850 (N_11850,N_7769,N_6926);
nor U11851 (N_11851,N_9265,N_7725);
or U11852 (N_11852,N_8840,N_7710);
xnor U11853 (N_11853,N_6760,N_8576);
nor U11854 (N_11854,N_7130,N_7122);
or U11855 (N_11855,N_8395,N_8704);
nor U11856 (N_11856,N_7140,N_8913);
nor U11857 (N_11857,N_7855,N_8288);
nand U11858 (N_11858,N_8421,N_6879);
and U11859 (N_11859,N_6388,N_7118);
or U11860 (N_11860,N_8348,N_7314);
or U11861 (N_11861,N_6295,N_8698);
nor U11862 (N_11862,N_8679,N_7764);
nor U11863 (N_11863,N_6267,N_7035);
or U11864 (N_11864,N_8564,N_7828);
and U11865 (N_11865,N_7608,N_9373);
and U11866 (N_11866,N_9139,N_8764);
nor U11867 (N_11867,N_8800,N_8987);
nor U11868 (N_11868,N_8607,N_6294);
nor U11869 (N_11869,N_8264,N_6520);
nand U11870 (N_11870,N_8904,N_8941);
or U11871 (N_11871,N_6900,N_6970);
nand U11872 (N_11872,N_7098,N_6758);
xnor U11873 (N_11873,N_8172,N_8406);
nand U11874 (N_11874,N_8191,N_6648);
and U11875 (N_11875,N_6341,N_7246);
xor U11876 (N_11876,N_6968,N_7388);
or U11877 (N_11877,N_8862,N_7289);
xnor U11878 (N_11878,N_7788,N_7178);
or U11879 (N_11879,N_6296,N_9329);
and U11880 (N_11880,N_7906,N_6792);
nor U11881 (N_11881,N_6324,N_8650);
xor U11882 (N_11882,N_8427,N_8692);
nand U11883 (N_11883,N_8375,N_7593);
and U11884 (N_11884,N_9126,N_9326);
and U11885 (N_11885,N_7631,N_8449);
nor U11886 (N_11886,N_9190,N_6721);
or U11887 (N_11887,N_7136,N_7822);
nand U11888 (N_11888,N_6688,N_8609);
nand U11889 (N_11889,N_6815,N_7722);
or U11890 (N_11890,N_6669,N_7401);
xor U11891 (N_11891,N_7746,N_8676);
nor U11892 (N_11892,N_6376,N_7622);
or U11893 (N_11893,N_6361,N_8283);
or U11894 (N_11894,N_7867,N_7574);
nor U11895 (N_11895,N_9330,N_6279);
nor U11896 (N_11896,N_8498,N_7048);
nand U11897 (N_11897,N_7140,N_7143);
xnor U11898 (N_11898,N_7129,N_9155);
and U11899 (N_11899,N_8050,N_9002);
xor U11900 (N_11900,N_6883,N_7536);
and U11901 (N_11901,N_7606,N_9364);
xor U11902 (N_11902,N_7746,N_8411);
or U11903 (N_11903,N_8436,N_7259);
nor U11904 (N_11904,N_8406,N_8786);
nand U11905 (N_11905,N_8541,N_8244);
or U11906 (N_11906,N_7290,N_6467);
or U11907 (N_11907,N_8889,N_7353);
nand U11908 (N_11908,N_8698,N_7046);
xnor U11909 (N_11909,N_8627,N_8414);
and U11910 (N_11910,N_8169,N_8167);
nor U11911 (N_11911,N_6821,N_9008);
and U11912 (N_11912,N_6584,N_9279);
and U11913 (N_11913,N_9164,N_8422);
xor U11914 (N_11914,N_7049,N_8559);
or U11915 (N_11915,N_7930,N_6293);
and U11916 (N_11916,N_7705,N_8759);
xnor U11917 (N_11917,N_7964,N_6820);
nand U11918 (N_11918,N_8251,N_6460);
nor U11919 (N_11919,N_7648,N_7940);
and U11920 (N_11920,N_8389,N_8831);
and U11921 (N_11921,N_8990,N_6588);
nand U11922 (N_11922,N_9091,N_7533);
nand U11923 (N_11923,N_8407,N_9128);
nor U11924 (N_11924,N_6638,N_6645);
xnor U11925 (N_11925,N_8065,N_7244);
or U11926 (N_11926,N_6629,N_6891);
nor U11927 (N_11927,N_9135,N_7582);
xnor U11928 (N_11928,N_6435,N_7241);
nand U11929 (N_11929,N_6564,N_8087);
and U11930 (N_11930,N_6906,N_8206);
and U11931 (N_11931,N_8955,N_8215);
nand U11932 (N_11932,N_8250,N_7620);
and U11933 (N_11933,N_9252,N_9358);
xnor U11934 (N_11934,N_8664,N_6351);
nor U11935 (N_11935,N_8780,N_7073);
nor U11936 (N_11936,N_8291,N_7969);
nand U11937 (N_11937,N_6345,N_6535);
and U11938 (N_11938,N_7201,N_6440);
nor U11939 (N_11939,N_6523,N_8785);
nand U11940 (N_11940,N_7534,N_8232);
nor U11941 (N_11941,N_8071,N_7678);
nand U11942 (N_11942,N_7382,N_8919);
xnor U11943 (N_11943,N_8351,N_6669);
or U11944 (N_11944,N_8915,N_7663);
and U11945 (N_11945,N_7722,N_9346);
nand U11946 (N_11946,N_6427,N_8396);
xor U11947 (N_11947,N_8963,N_7073);
nor U11948 (N_11948,N_8310,N_6345);
and U11949 (N_11949,N_7266,N_7571);
nand U11950 (N_11950,N_7659,N_8120);
xor U11951 (N_11951,N_7743,N_7139);
xnor U11952 (N_11952,N_8250,N_8024);
xnor U11953 (N_11953,N_6510,N_8267);
and U11954 (N_11954,N_9342,N_6810);
nand U11955 (N_11955,N_6459,N_6668);
xor U11956 (N_11956,N_7648,N_9194);
nand U11957 (N_11957,N_8514,N_7125);
nand U11958 (N_11958,N_8199,N_7895);
nor U11959 (N_11959,N_8080,N_8662);
xnor U11960 (N_11960,N_6647,N_7519);
xnor U11961 (N_11961,N_7864,N_9044);
or U11962 (N_11962,N_8161,N_6265);
nor U11963 (N_11963,N_6764,N_7148);
or U11964 (N_11964,N_8385,N_7433);
xnor U11965 (N_11965,N_8005,N_9307);
or U11966 (N_11966,N_8853,N_8946);
and U11967 (N_11967,N_8291,N_8399);
nand U11968 (N_11968,N_8841,N_7559);
nor U11969 (N_11969,N_7753,N_6251);
nor U11970 (N_11970,N_6448,N_8565);
or U11971 (N_11971,N_7114,N_7793);
xnor U11972 (N_11972,N_7237,N_6816);
and U11973 (N_11973,N_6398,N_7917);
xor U11974 (N_11974,N_6313,N_8892);
or U11975 (N_11975,N_8674,N_6508);
xnor U11976 (N_11976,N_8025,N_7924);
and U11977 (N_11977,N_7926,N_7158);
nand U11978 (N_11978,N_6307,N_8106);
or U11979 (N_11979,N_8904,N_8346);
xor U11980 (N_11980,N_9239,N_7386);
xor U11981 (N_11981,N_8135,N_9316);
nand U11982 (N_11982,N_6903,N_8725);
nand U11983 (N_11983,N_7621,N_9074);
or U11984 (N_11984,N_8341,N_8511);
and U11985 (N_11985,N_8935,N_8348);
or U11986 (N_11986,N_9107,N_7369);
nand U11987 (N_11987,N_8324,N_9285);
or U11988 (N_11988,N_7786,N_7633);
or U11989 (N_11989,N_7366,N_8446);
nor U11990 (N_11990,N_9072,N_6645);
nand U11991 (N_11991,N_7151,N_7430);
and U11992 (N_11992,N_8530,N_7855);
and U11993 (N_11993,N_8905,N_7176);
and U11994 (N_11994,N_6640,N_6831);
and U11995 (N_11995,N_7977,N_6771);
nor U11996 (N_11996,N_8989,N_6662);
xor U11997 (N_11997,N_7911,N_7210);
and U11998 (N_11998,N_7963,N_8305);
nand U11999 (N_11999,N_7964,N_9209);
nand U12000 (N_12000,N_6391,N_8238);
nand U12001 (N_12001,N_8006,N_8633);
or U12002 (N_12002,N_6489,N_6472);
xnor U12003 (N_12003,N_6758,N_9372);
or U12004 (N_12004,N_6380,N_7772);
nand U12005 (N_12005,N_8458,N_8191);
xnor U12006 (N_12006,N_8584,N_6717);
or U12007 (N_12007,N_6946,N_6285);
nor U12008 (N_12008,N_7889,N_6526);
and U12009 (N_12009,N_7337,N_7082);
or U12010 (N_12010,N_8379,N_7503);
nor U12011 (N_12011,N_6703,N_7040);
and U12012 (N_12012,N_7634,N_6489);
nor U12013 (N_12013,N_6420,N_9042);
or U12014 (N_12014,N_6342,N_7007);
or U12015 (N_12015,N_8131,N_9115);
and U12016 (N_12016,N_7722,N_8211);
nand U12017 (N_12017,N_6863,N_8601);
nor U12018 (N_12018,N_6749,N_6823);
or U12019 (N_12019,N_7852,N_7261);
nand U12020 (N_12020,N_7205,N_7352);
xor U12021 (N_12021,N_7963,N_6490);
or U12022 (N_12022,N_7871,N_9346);
or U12023 (N_12023,N_7938,N_7070);
nand U12024 (N_12024,N_9120,N_7214);
xnor U12025 (N_12025,N_8708,N_7018);
or U12026 (N_12026,N_8829,N_6305);
xor U12027 (N_12027,N_6536,N_8400);
nor U12028 (N_12028,N_8229,N_8428);
nor U12029 (N_12029,N_6624,N_7695);
nor U12030 (N_12030,N_8429,N_8472);
nand U12031 (N_12031,N_9304,N_9116);
nand U12032 (N_12032,N_8710,N_7365);
nand U12033 (N_12033,N_7588,N_7450);
xor U12034 (N_12034,N_9150,N_8330);
and U12035 (N_12035,N_8339,N_7088);
nand U12036 (N_12036,N_6496,N_9010);
and U12037 (N_12037,N_7759,N_7783);
and U12038 (N_12038,N_8300,N_7384);
and U12039 (N_12039,N_8521,N_6922);
xnor U12040 (N_12040,N_7148,N_8122);
or U12041 (N_12041,N_7990,N_8037);
and U12042 (N_12042,N_6888,N_7790);
xnor U12043 (N_12043,N_7203,N_7948);
and U12044 (N_12044,N_9240,N_9371);
xor U12045 (N_12045,N_6250,N_7669);
nand U12046 (N_12046,N_6325,N_9084);
nor U12047 (N_12047,N_7242,N_8840);
nor U12048 (N_12048,N_8960,N_8509);
and U12049 (N_12049,N_7989,N_7612);
nor U12050 (N_12050,N_6579,N_6303);
nand U12051 (N_12051,N_8569,N_8398);
xor U12052 (N_12052,N_8812,N_7276);
nor U12053 (N_12053,N_8699,N_7073);
nand U12054 (N_12054,N_9244,N_6352);
or U12055 (N_12055,N_7386,N_8972);
xor U12056 (N_12056,N_7352,N_6533);
nand U12057 (N_12057,N_8609,N_8022);
or U12058 (N_12058,N_8119,N_8406);
nand U12059 (N_12059,N_7987,N_6573);
and U12060 (N_12060,N_8818,N_7100);
nand U12061 (N_12061,N_7902,N_9057);
and U12062 (N_12062,N_9210,N_7838);
xor U12063 (N_12063,N_6509,N_7847);
nand U12064 (N_12064,N_7878,N_7611);
nor U12065 (N_12065,N_8547,N_9290);
nand U12066 (N_12066,N_9318,N_6310);
or U12067 (N_12067,N_6669,N_8160);
or U12068 (N_12068,N_6541,N_8597);
or U12069 (N_12069,N_8642,N_7951);
nand U12070 (N_12070,N_7977,N_7150);
nor U12071 (N_12071,N_7333,N_6439);
xnor U12072 (N_12072,N_8090,N_9157);
or U12073 (N_12073,N_6557,N_8015);
and U12074 (N_12074,N_6563,N_6382);
or U12075 (N_12075,N_7435,N_8605);
nor U12076 (N_12076,N_8358,N_7999);
nor U12077 (N_12077,N_8662,N_7931);
and U12078 (N_12078,N_6868,N_6648);
or U12079 (N_12079,N_8217,N_7775);
nor U12080 (N_12080,N_8374,N_6848);
nand U12081 (N_12081,N_6304,N_8854);
xor U12082 (N_12082,N_7178,N_8761);
nor U12083 (N_12083,N_6890,N_8745);
nand U12084 (N_12084,N_8853,N_7171);
nand U12085 (N_12085,N_7641,N_6309);
and U12086 (N_12086,N_8934,N_8864);
nand U12087 (N_12087,N_8047,N_7809);
nand U12088 (N_12088,N_8208,N_6345);
and U12089 (N_12089,N_8224,N_8907);
nand U12090 (N_12090,N_7988,N_8851);
or U12091 (N_12091,N_6898,N_6983);
nor U12092 (N_12092,N_8099,N_9103);
nand U12093 (N_12093,N_6784,N_6472);
nor U12094 (N_12094,N_8204,N_8066);
and U12095 (N_12095,N_6644,N_7577);
and U12096 (N_12096,N_6943,N_7201);
xor U12097 (N_12097,N_7391,N_8303);
nand U12098 (N_12098,N_9015,N_9055);
xor U12099 (N_12099,N_6479,N_7766);
nand U12100 (N_12100,N_7388,N_6612);
and U12101 (N_12101,N_6958,N_7209);
xor U12102 (N_12102,N_7946,N_9203);
nand U12103 (N_12103,N_8690,N_6408);
and U12104 (N_12104,N_6410,N_7669);
nor U12105 (N_12105,N_7548,N_7555);
and U12106 (N_12106,N_8391,N_8890);
and U12107 (N_12107,N_7580,N_6741);
and U12108 (N_12108,N_8784,N_8658);
nor U12109 (N_12109,N_8199,N_8319);
nor U12110 (N_12110,N_6445,N_8848);
nor U12111 (N_12111,N_7075,N_8411);
and U12112 (N_12112,N_8590,N_6995);
and U12113 (N_12113,N_6726,N_8818);
xor U12114 (N_12114,N_7946,N_6332);
and U12115 (N_12115,N_7132,N_7462);
or U12116 (N_12116,N_7499,N_8647);
or U12117 (N_12117,N_7652,N_7765);
nand U12118 (N_12118,N_7663,N_7954);
nand U12119 (N_12119,N_8226,N_7625);
or U12120 (N_12120,N_8189,N_7088);
nor U12121 (N_12121,N_6908,N_6907);
and U12122 (N_12122,N_9356,N_9088);
nand U12123 (N_12123,N_8375,N_6561);
nand U12124 (N_12124,N_8641,N_7777);
nand U12125 (N_12125,N_9330,N_6867);
nand U12126 (N_12126,N_8171,N_7596);
and U12127 (N_12127,N_9323,N_9157);
xor U12128 (N_12128,N_7595,N_7328);
or U12129 (N_12129,N_6693,N_7563);
nor U12130 (N_12130,N_8365,N_9288);
or U12131 (N_12131,N_6737,N_6454);
or U12132 (N_12132,N_6632,N_9065);
nor U12133 (N_12133,N_6285,N_7346);
or U12134 (N_12134,N_6499,N_8080);
nand U12135 (N_12135,N_6719,N_9325);
or U12136 (N_12136,N_9272,N_6694);
nor U12137 (N_12137,N_8164,N_8917);
nand U12138 (N_12138,N_8623,N_7861);
nor U12139 (N_12139,N_7501,N_7764);
nor U12140 (N_12140,N_6620,N_7235);
xnor U12141 (N_12141,N_7839,N_7883);
xnor U12142 (N_12142,N_6773,N_8850);
xnor U12143 (N_12143,N_9281,N_7252);
nor U12144 (N_12144,N_7788,N_6264);
xor U12145 (N_12145,N_6649,N_8015);
nand U12146 (N_12146,N_6790,N_7232);
nand U12147 (N_12147,N_6514,N_7545);
xor U12148 (N_12148,N_6982,N_7992);
nor U12149 (N_12149,N_7725,N_6674);
nand U12150 (N_12150,N_6990,N_7065);
nor U12151 (N_12151,N_8772,N_6786);
nor U12152 (N_12152,N_8605,N_9031);
and U12153 (N_12153,N_8966,N_7844);
nand U12154 (N_12154,N_6579,N_9301);
nor U12155 (N_12155,N_9357,N_6697);
nor U12156 (N_12156,N_8908,N_7971);
xnor U12157 (N_12157,N_7408,N_6667);
or U12158 (N_12158,N_8296,N_8917);
or U12159 (N_12159,N_9064,N_6860);
nor U12160 (N_12160,N_7581,N_7068);
and U12161 (N_12161,N_6265,N_8129);
xnor U12162 (N_12162,N_8126,N_6887);
nor U12163 (N_12163,N_7930,N_9248);
xnor U12164 (N_12164,N_8661,N_8825);
and U12165 (N_12165,N_6455,N_7901);
nand U12166 (N_12166,N_8488,N_6537);
xor U12167 (N_12167,N_8237,N_7661);
or U12168 (N_12168,N_7861,N_6979);
nand U12169 (N_12169,N_9309,N_9320);
and U12170 (N_12170,N_6977,N_9137);
xnor U12171 (N_12171,N_6815,N_7429);
nand U12172 (N_12172,N_7876,N_7480);
or U12173 (N_12173,N_7856,N_8792);
nand U12174 (N_12174,N_9057,N_8944);
and U12175 (N_12175,N_7151,N_7766);
or U12176 (N_12176,N_8723,N_7370);
or U12177 (N_12177,N_8035,N_9032);
nand U12178 (N_12178,N_8610,N_7824);
nand U12179 (N_12179,N_6428,N_7809);
nor U12180 (N_12180,N_7579,N_9123);
and U12181 (N_12181,N_6375,N_6978);
and U12182 (N_12182,N_8604,N_6338);
xnor U12183 (N_12183,N_9143,N_6744);
xor U12184 (N_12184,N_7072,N_7146);
nand U12185 (N_12185,N_7506,N_6886);
xor U12186 (N_12186,N_6854,N_8601);
xor U12187 (N_12187,N_7696,N_6256);
nor U12188 (N_12188,N_8426,N_7293);
nand U12189 (N_12189,N_7348,N_8060);
or U12190 (N_12190,N_6348,N_8848);
nand U12191 (N_12191,N_7011,N_7501);
xnor U12192 (N_12192,N_9329,N_8587);
xor U12193 (N_12193,N_6862,N_8598);
xor U12194 (N_12194,N_6541,N_7333);
xnor U12195 (N_12195,N_7483,N_6594);
or U12196 (N_12196,N_8684,N_8674);
and U12197 (N_12197,N_7715,N_6392);
and U12198 (N_12198,N_8019,N_9003);
nor U12199 (N_12199,N_6866,N_7849);
xor U12200 (N_12200,N_6643,N_7352);
or U12201 (N_12201,N_8854,N_7512);
or U12202 (N_12202,N_7917,N_8942);
xnor U12203 (N_12203,N_8664,N_7837);
nor U12204 (N_12204,N_6262,N_8984);
or U12205 (N_12205,N_9191,N_7617);
nand U12206 (N_12206,N_8727,N_8147);
xnor U12207 (N_12207,N_9015,N_7783);
nor U12208 (N_12208,N_8367,N_8973);
or U12209 (N_12209,N_8542,N_6819);
nor U12210 (N_12210,N_6676,N_9368);
nor U12211 (N_12211,N_9131,N_8676);
nor U12212 (N_12212,N_6959,N_6639);
nor U12213 (N_12213,N_7030,N_7285);
xnor U12214 (N_12214,N_9239,N_7137);
and U12215 (N_12215,N_9299,N_9289);
and U12216 (N_12216,N_8731,N_8530);
nand U12217 (N_12217,N_7456,N_7150);
and U12218 (N_12218,N_9066,N_9020);
nand U12219 (N_12219,N_7392,N_6733);
nor U12220 (N_12220,N_6537,N_6559);
nor U12221 (N_12221,N_7295,N_7649);
or U12222 (N_12222,N_8487,N_7748);
xnor U12223 (N_12223,N_9021,N_7817);
and U12224 (N_12224,N_8006,N_7156);
nand U12225 (N_12225,N_8754,N_6510);
nor U12226 (N_12226,N_6962,N_8460);
xor U12227 (N_12227,N_7169,N_8414);
nor U12228 (N_12228,N_7756,N_7465);
or U12229 (N_12229,N_6724,N_7630);
or U12230 (N_12230,N_6962,N_6659);
xnor U12231 (N_12231,N_6614,N_7301);
or U12232 (N_12232,N_8941,N_6673);
and U12233 (N_12233,N_7363,N_6445);
and U12234 (N_12234,N_7970,N_9053);
or U12235 (N_12235,N_8333,N_8482);
and U12236 (N_12236,N_9097,N_7400);
nand U12237 (N_12237,N_6608,N_8770);
nor U12238 (N_12238,N_7974,N_8864);
and U12239 (N_12239,N_6420,N_7598);
xnor U12240 (N_12240,N_6265,N_8296);
nand U12241 (N_12241,N_7137,N_6655);
and U12242 (N_12242,N_7162,N_6509);
nor U12243 (N_12243,N_8495,N_6403);
nand U12244 (N_12244,N_8730,N_8980);
nand U12245 (N_12245,N_6378,N_7625);
xor U12246 (N_12246,N_7957,N_8767);
or U12247 (N_12247,N_7577,N_9314);
xnor U12248 (N_12248,N_8691,N_8763);
xnor U12249 (N_12249,N_7076,N_8726);
or U12250 (N_12250,N_7098,N_7340);
nand U12251 (N_12251,N_9055,N_9083);
nor U12252 (N_12252,N_8975,N_7945);
xor U12253 (N_12253,N_6959,N_8042);
xnor U12254 (N_12254,N_8554,N_7958);
nand U12255 (N_12255,N_7332,N_8460);
and U12256 (N_12256,N_7629,N_8346);
nor U12257 (N_12257,N_6600,N_7484);
nand U12258 (N_12258,N_9208,N_8683);
nand U12259 (N_12259,N_8140,N_9175);
xor U12260 (N_12260,N_8605,N_7578);
and U12261 (N_12261,N_9168,N_7547);
or U12262 (N_12262,N_6455,N_6658);
or U12263 (N_12263,N_7000,N_7300);
xnor U12264 (N_12264,N_7934,N_6937);
nor U12265 (N_12265,N_7239,N_6846);
or U12266 (N_12266,N_9042,N_7627);
nand U12267 (N_12267,N_7818,N_9143);
or U12268 (N_12268,N_6858,N_6968);
or U12269 (N_12269,N_9022,N_8704);
xnor U12270 (N_12270,N_7584,N_8136);
xor U12271 (N_12271,N_8360,N_8840);
nand U12272 (N_12272,N_7985,N_6545);
nor U12273 (N_12273,N_7700,N_9219);
nand U12274 (N_12274,N_7641,N_6379);
and U12275 (N_12275,N_8242,N_8977);
or U12276 (N_12276,N_7186,N_7725);
xor U12277 (N_12277,N_9336,N_6729);
or U12278 (N_12278,N_8848,N_6512);
nor U12279 (N_12279,N_7754,N_6630);
and U12280 (N_12280,N_6538,N_7153);
or U12281 (N_12281,N_8371,N_8970);
nor U12282 (N_12282,N_7180,N_7178);
xor U12283 (N_12283,N_7949,N_7835);
xnor U12284 (N_12284,N_7962,N_8288);
and U12285 (N_12285,N_7297,N_7451);
nor U12286 (N_12286,N_9234,N_6861);
nand U12287 (N_12287,N_8066,N_8286);
nor U12288 (N_12288,N_7774,N_7963);
nand U12289 (N_12289,N_6824,N_7778);
and U12290 (N_12290,N_7329,N_6842);
nand U12291 (N_12291,N_7740,N_8240);
nor U12292 (N_12292,N_8879,N_8046);
xor U12293 (N_12293,N_8722,N_9273);
nor U12294 (N_12294,N_6955,N_8206);
nand U12295 (N_12295,N_7942,N_9299);
and U12296 (N_12296,N_9133,N_6434);
or U12297 (N_12297,N_8321,N_6498);
nor U12298 (N_12298,N_6392,N_8535);
or U12299 (N_12299,N_6969,N_8269);
nor U12300 (N_12300,N_7604,N_8920);
nand U12301 (N_12301,N_7041,N_9077);
xor U12302 (N_12302,N_8693,N_7627);
nor U12303 (N_12303,N_7981,N_6937);
xor U12304 (N_12304,N_6394,N_8966);
or U12305 (N_12305,N_6279,N_8616);
and U12306 (N_12306,N_7938,N_8031);
nand U12307 (N_12307,N_7773,N_7166);
and U12308 (N_12308,N_8655,N_6296);
xor U12309 (N_12309,N_8052,N_8887);
nand U12310 (N_12310,N_8752,N_7903);
nand U12311 (N_12311,N_7583,N_9037);
xnor U12312 (N_12312,N_8389,N_6472);
nand U12313 (N_12313,N_7764,N_7006);
and U12314 (N_12314,N_7005,N_8069);
nand U12315 (N_12315,N_6666,N_7303);
nor U12316 (N_12316,N_8737,N_7912);
and U12317 (N_12317,N_6404,N_7137);
or U12318 (N_12318,N_7645,N_9349);
nor U12319 (N_12319,N_7735,N_7584);
nor U12320 (N_12320,N_7722,N_8753);
or U12321 (N_12321,N_8546,N_9307);
xor U12322 (N_12322,N_6283,N_6357);
nand U12323 (N_12323,N_7648,N_7462);
xor U12324 (N_12324,N_9273,N_8125);
nor U12325 (N_12325,N_6604,N_7500);
or U12326 (N_12326,N_8793,N_6914);
nand U12327 (N_12327,N_6773,N_9149);
or U12328 (N_12328,N_8269,N_8326);
nand U12329 (N_12329,N_7349,N_7464);
xor U12330 (N_12330,N_7502,N_7529);
and U12331 (N_12331,N_9350,N_8017);
or U12332 (N_12332,N_8088,N_7697);
nor U12333 (N_12333,N_7800,N_6669);
nor U12334 (N_12334,N_6543,N_6291);
xor U12335 (N_12335,N_8220,N_7904);
xor U12336 (N_12336,N_7412,N_7556);
xnor U12337 (N_12337,N_8304,N_6940);
nor U12338 (N_12338,N_8785,N_6286);
or U12339 (N_12339,N_9233,N_6282);
xor U12340 (N_12340,N_8304,N_8428);
xnor U12341 (N_12341,N_8257,N_7979);
or U12342 (N_12342,N_8429,N_8986);
and U12343 (N_12343,N_8582,N_7584);
or U12344 (N_12344,N_7795,N_9065);
or U12345 (N_12345,N_8628,N_7383);
or U12346 (N_12346,N_8449,N_7497);
nand U12347 (N_12347,N_9232,N_7534);
or U12348 (N_12348,N_9223,N_8916);
nand U12349 (N_12349,N_6859,N_7531);
nand U12350 (N_12350,N_6571,N_8830);
and U12351 (N_12351,N_6447,N_8130);
or U12352 (N_12352,N_7359,N_7332);
nand U12353 (N_12353,N_6939,N_6447);
and U12354 (N_12354,N_7796,N_6260);
or U12355 (N_12355,N_7090,N_9200);
or U12356 (N_12356,N_7964,N_8106);
xor U12357 (N_12357,N_7565,N_7065);
nor U12358 (N_12358,N_7065,N_8548);
and U12359 (N_12359,N_8006,N_8754);
nand U12360 (N_12360,N_6925,N_8210);
xor U12361 (N_12361,N_8488,N_7229);
nor U12362 (N_12362,N_7437,N_6425);
or U12363 (N_12363,N_6441,N_6814);
or U12364 (N_12364,N_7975,N_6801);
xor U12365 (N_12365,N_7023,N_9307);
nand U12366 (N_12366,N_7484,N_6994);
nor U12367 (N_12367,N_8613,N_8108);
nand U12368 (N_12368,N_6499,N_7448);
nor U12369 (N_12369,N_7798,N_8727);
or U12370 (N_12370,N_8465,N_6581);
nand U12371 (N_12371,N_6733,N_8340);
nand U12372 (N_12372,N_6663,N_8529);
nor U12373 (N_12373,N_9278,N_6394);
and U12374 (N_12374,N_6324,N_7811);
or U12375 (N_12375,N_8592,N_8853);
nor U12376 (N_12376,N_7313,N_6322);
xnor U12377 (N_12377,N_8689,N_9020);
nand U12378 (N_12378,N_6395,N_8546);
nand U12379 (N_12379,N_9080,N_9316);
xor U12380 (N_12380,N_6822,N_6359);
nor U12381 (N_12381,N_6408,N_8163);
nor U12382 (N_12382,N_6911,N_6634);
nand U12383 (N_12383,N_7855,N_6305);
nor U12384 (N_12384,N_6413,N_8268);
and U12385 (N_12385,N_7890,N_8856);
nand U12386 (N_12386,N_8589,N_8912);
nand U12387 (N_12387,N_6299,N_7122);
and U12388 (N_12388,N_8769,N_8396);
xnor U12389 (N_12389,N_9077,N_6297);
xnor U12390 (N_12390,N_7365,N_7218);
nor U12391 (N_12391,N_6425,N_6265);
and U12392 (N_12392,N_7202,N_7615);
nand U12393 (N_12393,N_8918,N_7226);
nor U12394 (N_12394,N_9219,N_8858);
nor U12395 (N_12395,N_8151,N_8811);
nor U12396 (N_12396,N_6788,N_7986);
nand U12397 (N_12397,N_7348,N_7484);
nor U12398 (N_12398,N_6658,N_8028);
nand U12399 (N_12399,N_6690,N_8724);
and U12400 (N_12400,N_7471,N_8369);
nor U12401 (N_12401,N_7640,N_8423);
nor U12402 (N_12402,N_9082,N_8353);
and U12403 (N_12403,N_9242,N_9159);
xnor U12404 (N_12404,N_8548,N_7209);
nor U12405 (N_12405,N_6653,N_9124);
xor U12406 (N_12406,N_6444,N_7697);
xor U12407 (N_12407,N_6638,N_9100);
nand U12408 (N_12408,N_9144,N_8843);
or U12409 (N_12409,N_8369,N_6642);
nand U12410 (N_12410,N_7306,N_7485);
or U12411 (N_12411,N_8010,N_6253);
or U12412 (N_12412,N_7500,N_8565);
xor U12413 (N_12413,N_7388,N_7709);
xor U12414 (N_12414,N_6905,N_6388);
nand U12415 (N_12415,N_7648,N_7075);
nor U12416 (N_12416,N_7347,N_7090);
nand U12417 (N_12417,N_6297,N_6970);
or U12418 (N_12418,N_8796,N_7188);
or U12419 (N_12419,N_7884,N_7096);
xnor U12420 (N_12420,N_8466,N_9010);
or U12421 (N_12421,N_7794,N_6830);
xor U12422 (N_12422,N_6271,N_7015);
or U12423 (N_12423,N_6367,N_8909);
nand U12424 (N_12424,N_6369,N_7526);
nand U12425 (N_12425,N_9320,N_8629);
xnor U12426 (N_12426,N_7659,N_7608);
nor U12427 (N_12427,N_6686,N_6551);
or U12428 (N_12428,N_8700,N_8943);
nor U12429 (N_12429,N_7170,N_8853);
and U12430 (N_12430,N_6785,N_6439);
and U12431 (N_12431,N_6545,N_7776);
xor U12432 (N_12432,N_8528,N_8336);
nand U12433 (N_12433,N_9284,N_6863);
xnor U12434 (N_12434,N_8332,N_6638);
xnor U12435 (N_12435,N_6847,N_9224);
nor U12436 (N_12436,N_9318,N_8921);
xor U12437 (N_12437,N_8923,N_8335);
and U12438 (N_12438,N_6713,N_9247);
nand U12439 (N_12439,N_9178,N_7819);
and U12440 (N_12440,N_9313,N_8870);
nor U12441 (N_12441,N_8690,N_9184);
or U12442 (N_12442,N_7442,N_7941);
or U12443 (N_12443,N_8066,N_7297);
and U12444 (N_12444,N_8231,N_6422);
or U12445 (N_12445,N_6866,N_7137);
nor U12446 (N_12446,N_8830,N_8631);
nor U12447 (N_12447,N_6564,N_7732);
and U12448 (N_12448,N_8992,N_7144);
nor U12449 (N_12449,N_6253,N_6834);
nand U12450 (N_12450,N_8232,N_6761);
nand U12451 (N_12451,N_8786,N_6343);
or U12452 (N_12452,N_8955,N_6558);
nor U12453 (N_12453,N_7085,N_6286);
or U12454 (N_12454,N_7363,N_8009);
and U12455 (N_12455,N_9014,N_7650);
and U12456 (N_12456,N_8840,N_8566);
xnor U12457 (N_12457,N_8247,N_8062);
xnor U12458 (N_12458,N_6664,N_6758);
nor U12459 (N_12459,N_8005,N_6873);
or U12460 (N_12460,N_8215,N_6691);
nor U12461 (N_12461,N_6750,N_8787);
or U12462 (N_12462,N_6867,N_9164);
and U12463 (N_12463,N_6839,N_8501);
and U12464 (N_12464,N_8933,N_8701);
nand U12465 (N_12465,N_9326,N_9351);
nand U12466 (N_12466,N_8002,N_7819);
or U12467 (N_12467,N_6864,N_7564);
nand U12468 (N_12468,N_7278,N_9063);
nor U12469 (N_12469,N_8169,N_7945);
or U12470 (N_12470,N_7432,N_7934);
or U12471 (N_12471,N_6653,N_8815);
nand U12472 (N_12472,N_8368,N_7819);
xor U12473 (N_12473,N_8820,N_8342);
nor U12474 (N_12474,N_7752,N_7744);
and U12475 (N_12475,N_8247,N_6338);
nor U12476 (N_12476,N_8949,N_7245);
nand U12477 (N_12477,N_8616,N_8574);
nand U12478 (N_12478,N_6275,N_7991);
and U12479 (N_12479,N_7058,N_7807);
or U12480 (N_12480,N_7723,N_7139);
nand U12481 (N_12481,N_9257,N_7923);
and U12482 (N_12482,N_6501,N_7784);
xnor U12483 (N_12483,N_6927,N_6759);
nand U12484 (N_12484,N_9215,N_6296);
or U12485 (N_12485,N_9317,N_7494);
and U12486 (N_12486,N_8143,N_8595);
nand U12487 (N_12487,N_7753,N_9352);
or U12488 (N_12488,N_7622,N_9070);
nand U12489 (N_12489,N_8085,N_8313);
and U12490 (N_12490,N_6474,N_7833);
nand U12491 (N_12491,N_8525,N_6509);
or U12492 (N_12492,N_7701,N_7939);
xnor U12493 (N_12493,N_6326,N_8151);
nor U12494 (N_12494,N_6591,N_7161);
nor U12495 (N_12495,N_8756,N_6582);
or U12496 (N_12496,N_6502,N_9108);
and U12497 (N_12497,N_8547,N_7869);
nand U12498 (N_12498,N_6605,N_7960);
nor U12499 (N_12499,N_8912,N_7383);
or U12500 (N_12500,N_12423,N_10000);
and U12501 (N_12501,N_9796,N_11611);
xnor U12502 (N_12502,N_11865,N_11423);
nand U12503 (N_12503,N_10483,N_11549);
and U12504 (N_12504,N_9521,N_11344);
or U12505 (N_12505,N_9606,N_10093);
and U12506 (N_12506,N_11825,N_11988);
nand U12507 (N_12507,N_10489,N_10485);
nor U12508 (N_12508,N_9994,N_11647);
nand U12509 (N_12509,N_10341,N_9765);
or U12510 (N_12510,N_11157,N_10389);
nand U12511 (N_12511,N_12003,N_10549);
nor U12512 (N_12512,N_10470,N_10421);
nand U12513 (N_12513,N_9855,N_10128);
or U12514 (N_12514,N_11883,N_9798);
or U12515 (N_12515,N_11938,N_10158);
xnor U12516 (N_12516,N_11045,N_11340);
nand U12517 (N_12517,N_11720,N_10431);
and U12518 (N_12518,N_11576,N_9624);
xnor U12519 (N_12519,N_9467,N_9492);
or U12520 (N_12520,N_10687,N_10346);
xnor U12521 (N_12521,N_9678,N_10698);
xnor U12522 (N_12522,N_11775,N_10608);
nand U12523 (N_12523,N_9518,N_11319);
xor U12524 (N_12524,N_9739,N_11718);
xnor U12525 (N_12525,N_12133,N_11134);
or U12526 (N_12526,N_11350,N_10873);
and U12527 (N_12527,N_10927,N_10875);
nand U12528 (N_12528,N_12260,N_12344);
xnor U12529 (N_12529,N_9752,N_10082);
nor U12530 (N_12530,N_11173,N_11447);
xnor U12531 (N_12531,N_10518,N_11884);
nor U12532 (N_12532,N_9968,N_11543);
or U12533 (N_12533,N_12055,N_11976);
nor U12534 (N_12534,N_11081,N_10386);
and U12535 (N_12535,N_12340,N_12446);
nand U12536 (N_12536,N_11843,N_11850);
and U12537 (N_12537,N_12225,N_9646);
and U12538 (N_12538,N_12450,N_11941);
nor U12539 (N_12539,N_9657,N_10270);
or U12540 (N_12540,N_10896,N_11547);
and U12541 (N_12541,N_11632,N_12256);
xnor U12542 (N_12542,N_12316,N_12164);
xnor U12543 (N_12543,N_10465,N_10006);
xnor U12544 (N_12544,N_11877,N_12426);
nand U12545 (N_12545,N_11180,N_12314);
nand U12546 (N_12546,N_12197,N_9864);
xnor U12547 (N_12547,N_11667,N_10350);
xnor U12548 (N_12548,N_11479,N_10318);
nand U12549 (N_12549,N_11672,N_10736);
and U12550 (N_12550,N_11221,N_11745);
nand U12551 (N_12551,N_10670,N_10028);
nor U12552 (N_12552,N_10340,N_10454);
and U12553 (N_12553,N_9986,N_9995);
and U12554 (N_12554,N_12390,N_9669);
nor U12555 (N_12555,N_11796,N_9948);
nor U12556 (N_12556,N_9918,N_9879);
xor U12557 (N_12557,N_10622,N_11737);
and U12558 (N_12558,N_9610,N_11234);
nand U12559 (N_12559,N_11087,N_10673);
and U12560 (N_12560,N_11156,N_10989);
or U12561 (N_12561,N_10111,N_10824);
xnor U12562 (N_12562,N_10576,N_10555);
or U12563 (N_12563,N_12474,N_9393);
nor U12564 (N_12564,N_10955,N_10807);
nor U12565 (N_12565,N_10027,N_10399);
or U12566 (N_12566,N_9852,N_10855);
xnor U12567 (N_12567,N_11978,N_9770);
xor U12568 (N_12568,N_11907,N_10262);
nand U12569 (N_12569,N_11658,N_11777);
and U12570 (N_12570,N_10065,N_12489);
and U12571 (N_12571,N_12192,N_9380);
and U12572 (N_12572,N_11762,N_11281);
or U12573 (N_12573,N_12351,N_9940);
xor U12574 (N_12574,N_9526,N_10564);
and U12575 (N_12575,N_11112,N_10906);
and U12576 (N_12576,N_10459,N_11058);
or U12577 (N_12577,N_11500,N_11585);
nor U12578 (N_12578,N_9885,N_10035);
and U12579 (N_12579,N_10813,N_12264);
and U12580 (N_12580,N_12274,N_11582);
and U12581 (N_12581,N_11577,N_11027);
or U12582 (N_12582,N_11609,N_12157);
or U12583 (N_12583,N_10209,N_11370);
nor U12584 (N_12584,N_10462,N_9447);
nor U12585 (N_12585,N_10204,N_10626);
nand U12586 (N_12586,N_11382,N_10393);
xor U12587 (N_12587,N_9453,N_12370);
nand U12588 (N_12588,N_12095,N_9750);
and U12589 (N_12589,N_11921,N_11627);
xor U12590 (N_12590,N_10812,N_11264);
nor U12591 (N_12591,N_11640,N_11930);
nand U12592 (N_12592,N_11397,N_12067);
or U12593 (N_12593,N_9426,N_10007);
or U12594 (N_12594,N_9621,N_11934);
and U12595 (N_12595,N_10550,N_11818);
and U12596 (N_12596,N_11636,N_10745);
or U12597 (N_12597,N_10832,N_10628);
nor U12598 (N_12598,N_11073,N_12103);
nor U12599 (N_12599,N_10806,N_11586);
nor U12600 (N_12600,N_11601,N_11455);
or U12601 (N_12601,N_10094,N_10309);
nor U12602 (N_12602,N_9910,N_9500);
nor U12603 (N_12603,N_11217,N_9830);
nor U12604 (N_12604,N_10743,N_9690);
nand U12605 (N_12605,N_12324,N_11613);
and U12606 (N_12606,N_12165,N_10566);
xor U12607 (N_12607,N_10423,N_12409);
nand U12608 (N_12608,N_11851,N_9697);
nand U12609 (N_12609,N_11761,N_9794);
or U12610 (N_12610,N_11856,N_12114);
xnor U12611 (N_12611,N_10985,N_12158);
or U12612 (N_12612,N_10468,N_10695);
nand U12613 (N_12613,N_11519,N_11629);
or U12614 (N_12614,N_9656,N_11469);
or U12615 (N_12615,N_10657,N_12288);
and U12616 (N_12616,N_11022,N_11573);
xor U12617 (N_12617,N_11411,N_12326);
or U12618 (N_12618,N_12054,N_11048);
or U12619 (N_12619,N_11853,N_12458);
nand U12620 (N_12620,N_9609,N_11969);
xor U12621 (N_12621,N_12074,N_10221);
nand U12622 (N_12622,N_11800,N_9875);
nand U12623 (N_12623,N_12081,N_10189);
nor U12624 (N_12624,N_9893,N_9441);
xnor U12625 (N_12625,N_10439,N_10026);
xor U12626 (N_12626,N_9754,N_9684);
and U12627 (N_12627,N_11278,N_9887);
nor U12628 (N_12628,N_9942,N_10900);
and U12629 (N_12629,N_10244,N_10598);
xor U12630 (N_12630,N_9615,N_9889);
and U12631 (N_12631,N_10357,N_10990);
or U12632 (N_12632,N_9776,N_11505);
nand U12633 (N_12633,N_10379,N_12290);
and U12634 (N_12634,N_11889,N_10636);
or U12635 (N_12635,N_11831,N_9861);
and U12636 (N_12636,N_9629,N_11736);
nor U12637 (N_12637,N_11915,N_12247);
nand U12638 (N_12638,N_10116,N_10764);
xor U12639 (N_12639,N_10649,N_12178);
xor U12640 (N_12640,N_9691,N_11031);
and U12641 (N_12641,N_11929,N_10982);
or U12642 (N_12642,N_11320,N_10495);
nor U12643 (N_12643,N_10652,N_10594);
and U12644 (N_12644,N_10302,N_11274);
nand U12645 (N_12645,N_11135,N_12002);
and U12646 (N_12646,N_11957,N_12477);
nand U12647 (N_12647,N_11768,N_9859);
xnor U12648 (N_12648,N_11716,N_11002);
and U12649 (N_12649,N_10269,N_9573);
or U12650 (N_12650,N_9975,N_10777);
nor U12651 (N_12651,N_11587,N_11024);
nand U12652 (N_12652,N_11171,N_9784);
and U12653 (N_12653,N_12100,N_9924);
xnor U12654 (N_12654,N_9486,N_10689);
nor U12655 (N_12655,N_11804,N_11682);
or U12656 (N_12656,N_9973,N_11291);
nand U12657 (N_12657,N_11896,N_11321);
and U12658 (N_12658,N_10690,N_11439);
nor U12659 (N_12659,N_11065,N_11757);
xor U12660 (N_12660,N_9682,N_12254);
nand U12661 (N_12661,N_9705,N_10897);
nand U12662 (N_12662,N_12308,N_11644);
xnor U12663 (N_12663,N_9632,N_11475);
nand U12664 (N_12664,N_10304,N_11289);
nand U12665 (N_12665,N_10735,N_11529);
and U12666 (N_12666,N_11679,N_10194);
nor U12667 (N_12667,N_11491,N_9804);
xor U12668 (N_12668,N_11922,N_11476);
nand U12669 (N_12669,N_9559,N_10306);
nor U12670 (N_12670,N_12377,N_10817);
nor U12671 (N_12671,N_12160,N_9555);
nor U12672 (N_12672,N_9759,N_12369);
xor U12673 (N_12673,N_9723,N_11082);
xnor U12674 (N_12674,N_11246,N_11396);
or U12675 (N_12675,N_10289,N_10208);
nor U12676 (N_12676,N_10829,N_11683);
nand U12677 (N_12677,N_10993,N_9415);
and U12678 (N_12678,N_12198,N_9671);
xor U12679 (N_12679,N_10766,N_10565);
nand U12680 (N_12680,N_12313,N_10215);
nand U12681 (N_12681,N_9626,N_10885);
nor U12682 (N_12682,N_11618,N_10863);
nor U12683 (N_12683,N_10138,N_12243);
and U12684 (N_12684,N_10883,N_10525);
xnor U12685 (N_12685,N_12478,N_11381);
and U12686 (N_12686,N_9480,N_10300);
or U12687 (N_12687,N_12154,N_10774);
nor U12688 (N_12688,N_9722,N_12436);
nand U12689 (N_12689,N_11697,N_9818);
nor U12690 (N_12690,N_11437,N_9895);
and U12691 (N_12691,N_12228,N_10298);
nand U12692 (N_12692,N_10152,N_11332);
xor U12693 (N_12693,N_12359,N_12043);
or U12694 (N_12694,N_9733,N_12123);
nand U12695 (N_12695,N_11545,N_11151);
nor U12696 (N_12696,N_11189,N_11598);
or U12697 (N_12697,N_10212,N_9542);
or U12698 (N_12698,N_11610,N_10106);
nor U12699 (N_12699,N_9886,N_9569);
nand U12700 (N_12700,N_10498,N_11981);
nor U12701 (N_12701,N_12309,N_10988);
nand U12702 (N_12702,N_10192,N_9422);
and U12703 (N_12703,N_11161,N_12498);
nand U12704 (N_12704,N_11226,N_10816);
nor U12705 (N_12705,N_10020,N_12125);
nand U12706 (N_12706,N_11528,N_11580);
nor U12707 (N_12707,N_10665,N_10014);
xnor U12708 (N_12708,N_10040,N_11669);
and U12709 (N_12709,N_9558,N_11861);
and U12710 (N_12710,N_12384,N_12296);
or U12711 (N_12711,N_10519,N_11742);
nor U12712 (N_12712,N_9915,N_11405);
nor U12713 (N_12713,N_12258,N_10281);
and U12714 (N_12714,N_11812,N_9931);
xnor U12715 (N_12715,N_11038,N_10602);
and U12716 (N_12716,N_9665,N_10995);
nand U12717 (N_12717,N_10382,N_11860);
or U12718 (N_12718,N_12315,N_9987);
xnor U12719 (N_12719,N_9427,N_9451);
or U12720 (N_12720,N_11003,N_9991);
xnor U12721 (N_12721,N_11025,N_12001);
xor U12722 (N_12722,N_11011,N_11443);
nor U12723 (N_12723,N_11122,N_10733);
xnor U12724 (N_12724,N_11449,N_10060);
and U12725 (N_12725,N_12229,N_11445);
xnor U12726 (N_12726,N_12271,N_11076);
or U12727 (N_12727,N_10137,N_11000);
xnor U12728 (N_12728,N_12008,N_11063);
xnor U12729 (N_12729,N_11402,N_11925);
nand U12730 (N_12730,N_11899,N_10823);
nor U12731 (N_12731,N_10090,N_9490);
nor U12732 (N_12732,N_10080,N_11673);
and U12733 (N_12733,N_10852,N_11385);
nand U12734 (N_12734,N_9571,N_11641);
nor U12735 (N_12735,N_11198,N_12029);
nor U12736 (N_12736,N_11318,N_10230);
nand U12737 (N_12737,N_12149,N_10238);
or U12738 (N_12738,N_11227,N_9737);
nand U12739 (N_12739,N_11743,N_9833);
xnor U12740 (N_12740,N_11079,N_10724);
xor U12741 (N_12741,N_11755,N_12028);
nor U12742 (N_12742,N_11653,N_12173);
nand U12743 (N_12743,N_10249,N_11404);
nor U12744 (N_12744,N_11815,N_10426);
nand U12745 (N_12745,N_9424,N_9382);
and U12746 (N_12746,N_10403,N_10680);
nor U12747 (N_12747,N_9772,N_10412);
or U12748 (N_12748,N_9841,N_9607);
and U12749 (N_12749,N_11124,N_11202);
xor U12750 (N_12750,N_10825,N_10157);
nor U12751 (N_12751,N_11717,N_11530);
xnor U12752 (N_12752,N_12257,N_9856);
or U12753 (N_12753,N_11193,N_11873);
nor U12754 (N_12754,N_11219,N_9799);
or U12755 (N_12755,N_10593,N_10449);
and U12756 (N_12756,N_11512,N_9988);
nand U12757 (N_12757,N_10172,N_10612);
and U12758 (N_12758,N_11563,N_11435);
and U12759 (N_12759,N_10941,N_11465);
nor U12760 (N_12760,N_9512,N_12082);
and U12761 (N_12761,N_9936,N_12382);
nand U12762 (N_12762,N_11015,N_11458);
nor U12763 (N_12763,N_10140,N_9420);
and U12764 (N_12764,N_9806,N_10641);
nor U12765 (N_12765,N_10059,N_11177);
or U12766 (N_12766,N_11758,N_9985);
and U12767 (N_12767,N_11018,N_11484);
xnor U12768 (N_12768,N_11814,N_10499);
and U12769 (N_12769,N_9557,N_12166);
and U12770 (N_12770,N_12244,N_11984);
xor U12771 (N_12771,N_11973,N_10126);
nand U12772 (N_12772,N_9658,N_10840);
nor U12773 (N_12773,N_10528,N_10229);
nand U12774 (N_12774,N_11952,N_9810);
xnor U12775 (N_12775,N_11591,N_11628);
nand U12776 (N_12776,N_9501,N_10542);
xor U12777 (N_12777,N_9548,N_12440);
xnor U12778 (N_12778,N_11971,N_11887);
nand U12779 (N_12779,N_11194,N_11571);
nand U12780 (N_12780,N_9703,N_12416);
nor U12781 (N_12781,N_10252,N_11779);
nand U12782 (N_12782,N_10540,N_10497);
and U12783 (N_12783,N_9726,N_11515);
xor U12784 (N_12784,N_9683,N_12345);
nor U12785 (N_12785,N_11313,N_10772);
nand U12786 (N_12786,N_10235,N_9633);
or U12787 (N_12787,N_10322,N_10938);
xor U12788 (N_12788,N_11798,N_11808);
xnor U12789 (N_12789,N_10992,N_10563);
xor U12790 (N_12790,N_10025,N_10307);
or U12791 (N_12791,N_11535,N_10678);
and U12792 (N_12792,N_11897,N_12253);
nand U12793 (N_12793,N_10022,N_10240);
and U12794 (N_12794,N_10672,N_9884);
or U12795 (N_12795,N_9728,N_11554);
xnor U12796 (N_12796,N_12194,N_11920);
and U12797 (N_12797,N_12062,N_10950);
nor U12798 (N_12798,N_11819,N_12325);
xor U12799 (N_12799,N_11729,N_12060);
xor U12800 (N_12800,N_11677,N_11538);
or U12801 (N_12801,N_10280,N_11365);
or U12802 (N_12802,N_10634,N_11150);
nor U12803 (N_12803,N_12145,N_11992);
nor U12804 (N_12804,N_10889,N_9568);
nand U12805 (N_12805,N_11413,N_9409);
nor U12806 (N_12806,N_10246,N_12338);
xnor U12807 (N_12807,N_11870,N_10818);
nand U12808 (N_12808,N_11725,N_11069);
xor U12809 (N_12809,N_9831,N_10871);
nand U12810 (N_12810,N_10409,N_10195);
xnor U12811 (N_12811,N_12053,N_9561);
xnor U12812 (N_12812,N_11662,N_11490);
xor U12813 (N_12813,N_11793,N_9530);
xnor U12814 (N_12814,N_10742,N_12318);
nand U12815 (N_12815,N_10492,N_9734);
nor U12816 (N_12816,N_12096,N_11652);
or U12817 (N_12817,N_12101,N_11050);
nor U12818 (N_12818,N_11533,N_10105);
xor U12819 (N_12819,N_11572,N_9820);
nor U12820 (N_12820,N_11004,N_11731);
or U12821 (N_12821,N_10952,N_10109);
or U12822 (N_12822,N_11041,N_12431);
nand U12823 (N_12823,N_11914,N_12452);
nor U12824 (N_12824,N_10477,N_9388);
or U12825 (N_12825,N_12168,N_11776);
nor U12826 (N_12826,N_11719,N_10908);
nor U12827 (N_12827,N_9470,N_11555);
nor U12828 (N_12828,N_12307,N_10384);
or U12829 (N_12829,N_11296,N_10274);
and U12830 (N_12830,N_10130,N_12201);
xor U12831 (N_12831,N_10323,N_11271);
nand U12832 (N_12832,N_10283,N_10414);
and U12833 (N_12833,N_10554,N_11136);
nand U12834 (N_12834,N_12366,N_11740);
and U12835 (N_12835,N_12089,N_10233);
and U12836 (N_12836,N_10964,N_12282);
nor U12837 (N_12837,N_11364,N_10888);
and U12838 (N_12838,N_10640,N_10044);
nor U12839 (N_12839,N_11408,N_12311);
nand U12840 (N_12840,N_11752,N_9768);
nand U12841 (N_12841,N_11649,N_11550);
xor U12842 (N_12842,N_11944,N_9466);
nand U12843 (N_12843,N_12070,N_10455);
nor U12844 (N_12844,N_10354,N_11709);
and U12845 (N_12845,N_12454,N_11966);
or U12846 (N_12846,N_12463,N_10490);
xnor U12847 (N_12847,N_12112,N_11272);
xnor U12848 (N_12848,N_9711,N_11374);
nor U12849 (N_12849,N_9954,N_11205);
nor U12850 (N_12850,N_10708,N_10308);
nor U12851 (N_12851,N_10432,N_9523);
nand U12852 (N_12852,N_11772,N_10784);
nand U12853 (N_12853,N_10599,N_10637);
and U12854 (N_12854,N_10436,N_10534);
or U12855 (N_12855,N_11149,N_10839);
or U12856 (N_12856,N_11049,N_11155);
and U12857 (N_12857,N_12215,N_10036);
nand U12858 (N_12858,N_9874,N_10174);
nor U12859 (N_12859,N_10218,N_9412);
nand U12860 (N_12860,N_10333,N_11305);
or U12861 (N_12861,N_9623,N_12039);
xor U12862 (N_12862,N_9921,N_10620);
xor U12863 (N_12863,N_9704,N_9731);
and U12864 (N_12864,N_12138,N_11108);
and U12865 (N_12865,N_10312,N_9938);
xnor U12866 (N_12866,N_11833,N_10775);
and U12867 (N_12867,N_11633,N_11287);
nor U12868 (N_12868,N_9536,N_9677);
nor U12869 (N_12869,N_10891,N_11144);
nor U12870 (N_12870,N_10630,N_11196);
nor U12871 (N_12871,N_11802,N_12073);
nor U12872 (N_12872,N_9989,N_10095);
or U12873 (N_12873,N_11336,N_11504);
and U12874 (N_12874,N_9517,N_11410);
nor U12875 (N_12875,N_11820,N_10925);
xnor U12876 (N_12876,N_10104,N_10131);
and U12877 (N_12877,N_9937,N_11960);
or U12878 (N_12878,N_10168,N_11747);
nand U12879 (N_12879,N_12167,N_12376);
or U12880 (N_12880,N_10547,N_12327);
xor U12881 (N_12881,N_10259,N_11859);
or U12882 (N_12882,N_10929,N_10255);
or U12883 (N_12883,N_10043,N_9976);
xor U12884 (N_12884,N_11078,N_11688);
and U12885 (N_12885,N_11561,N_10180);
nand U12886 (N_12886,N_11575,N_10648);
nor U12887 (N_12887,N_11551,N_12281);
or U12888 (N_12888,N_12413,N_12135);
nand U12889 (N_12889,N_9376,N_11837);
nand U12890 (N_12890,N_11212,N_11237);
or U12891 (N_12891,N_10256,N_9822);
xnor U12892 (N_12892,N_10729,N_11330);
nand U12893 (N_12893,N_11597,N_12050);
nand U12894 (N_12894,N_11308,N_10785);
and U12895 (N_12895,N_9899,N_10569);
nor U12896 (N_12896,N_11249,N_11839);
xnor U12897 (N_12897,N_10755,N_10857);
and U12898 (N_12898,N_10466,N_10344);
xor U12899 (N_12899,N_10974,N_10539);
xnor U12900 (N_12900,N_9503,N_10032);
and U12901 (N_12901,N_11461,N_11007);
nand U12902 (N_12902,N_10944,N_9552);
xnor U12903 (N_12903,N_11062,N_9418);
xnor U12904 (N_12904,N_10400,N_11084);
or U12905 (N_12905,N_9797,N_12461);
nand U12906 (N_12906,N_12321,N_9549);
and U12907 (N_12907,N_10512,N_9717);
or U12908 (N_12908,N_10385,N_11001);
or U12909 (N_12909,N_10214,N_9919);
or U12910 (N_12910,N_9745,N_12218);
nand U12911 (N_12911,N_12279,N_10753);
or U12912 (N_12912,N_12383,N_11497);
nor U12913 (N_12913,N_10515,N_10666);
and U12914 (N_12914,N_9449,N_12391);
or U12915 (N_12915,N_10050,N_11749);
xor U12916 (N_12916,N_11670,N_11399);
xor U12917 (N_12917,N_10161,N_10339);
nor U12918 (N_12918,N_9375,N_12429);
xnor U12919 (N_12919,N_10969,N_10228);
and U12920 (N_12920,N_9564,N_11692);
nor U12921 (N_12921,N_9867,N_10627);
nand U12922 (N_12922,N_10024,N_9757);
xor U12923 (N_12923,N_9625,N_11276);
nand U12924 (N_12924,N_11979,N_9904);
xor U12925 (N_12925,N_11524,N_11997);
and U12926 (N_12926,N_9967,N_10009);
or U12927 (N_12927,N_9844,N_11552);
nand U12928 (N_12928,N_12116,N_11029);
or U12929 (N_12929,N_10051,N_10031);
or U12930 (N_12930,N_11471,N_12373);
and U12931 (N_12931,N_12179,N_12221);
nor U12932 (N_12932,N_11970,N_11892);
xor U12933 (N_12933,N_10994,N_9812);
nor U12934 (N_12934,N_10019,N_9807);
and U12935 (N_12935,N_9461,N_12355);
nand U12936 (N_12936,N_10273,N_12358);
nand U12937 (N_12937,N_9958,N_10827);
or U12938 (N_12938,N_10750,N_10882);
and U12939 (N_12939,N_11603,N_11643);
nand U12940 (N_12940,N_10932,N_10790);
xnor U12941 (N_12941,N_10164,N_9850);
or U12942 (N_12942,N_9600,N_12038);
nor U12943 (N_12943,N_12386,N_12007);
xor U12944 (N_12944,N_11651,N_9709);
xnor U12945 (N_12945,N_12023,N_12346);
nand U12946 (N_12946,N_10902,N_9586);
or U12947 (N_12947,N_9576,N_12203);
nand U12948 (N_12948,N_10261,N_10848);
and U12949 (N_12949,N_11875,N_9787);
nor U12950 (N_12950,N_10746,N_11891);
nor U12951 (N_12951,N_10326,N_12083);
nand U12952 (N_12952,N_11541,N_9902);
or U12953 (N_12953,N_12206,N_11763);
nand U12954 (N_12954,N_12341,N_9680);
and U12955 (N_12955,N_11040,N_11253);
or U12956 (N_12956,N_11361,N_10844);
or U12957 (N_12957,N_10675,N_10162);
and U12958 (N_12958,N_10760,N_9716);
xor U12959 (N_12959,N_12350,N_12150);
nand U12960 (N_12960,N_12109,N_9898);
nor U12961 (N_12961,N_12335,N_12336);
nand U12962 (N_12962,N_11803,N_11834);
xnor U12963 (N_12963,N_9775,N_10702);
and U12964 (N_12964,N_9965,N_10658);
nor U12965 (N_12965,N_12414,N_10135);
and U12966 (N_12966,N_10954,N_10475);
or U12967 (N_12967,N_9990,N_10904);
and U12968 (N_12968,N_12402,N_11419);
or U12969 (N_12969,N_12273,N_12299);
or U12970 (N_12970,N_9494,N_11429);
and U12971 (N_12971,N_10311,N_9961);
and U12972 (N_12972,N_10940,N_11828);
and U12973 (N_12973,N_9592,N_10045);
or U12974 (N_12974,N_10617,N_11440);
nor U12975 (N_12975,N_12129,N_10802);
xor U12976 (N_12976,N_10072,N_10920);
xor U12977 (N_12977,N_10377,N_11666);
and U12978 (N_12978,N_11956,N_9909);
nand U12979 (N_12979,N_10008,N_11624);
xor U12980 (N_12980,N_10861,N_10717);
nand U12981 (N_12981,N_10860,N_9998);
xnor U12982 (N_12982,N_9676,N_11107);
nand U12983 (N_12983,N_10953,N_11055);
nor U12984 (N_12984,N_11895,N_11097);
nor U12985 (N_12985,N_10074,N_9992);
nand U12986 (N_12986,N_12422,N_9544);
and U12987 (N_12987,N_10038,N_9638);
xnor U12988 (N_12988,N_10797,N_10984);
xor U12989 (N_12989,N_10253,N_11844);
or U12990 (N_12990,N_10638,N_12380);
and U12991 (N_12991,N_9662,N_10623);
nor U12992 (N_12992,N_10416,N_12319);
nor U12993 (N_12993,N_11168,N_11514);
xor U12994 (N_12994,N_12151,N_11286);
or U12995 (N_12995,N_10321,N_10830);
nand U12996 (N_12996,N_12357,N_11255);
nand U12997 (N_12997,N_9802,N_11123);
and U12998 (N_12998,N_10084,N_11778);
or U12999 (N_12999,N_10338,N_11696);
nor U13000 (N_13000,N_10520,N_11511);
xor U13001 (N_13001,N_9399,N_10062);
or U13002 (N_13002,N_9378,N_11403);
nor U13003 (N_13003,N_9854,N_9878);
nand U13004 (N_13004,N_12491,N_10227);
and U13005 (N_13005,N_10912,N_10866);
and U13006 (N_13006,N_12453,N_10728);
xor U13007 (N_13007,N_10224,N_10754);
nor U13008 (N_13008,N_12022,N_11569);
nand U13009 (N_13009,N_11259,N_12122);
and U13010 (N_13010,N_9407,N_12249);
xnor U13011 (N_13011,N_12026,N_10887);
or U13012 (N_13012,N_9547,N_11166);
and U13013 (N_13013,N_11338,N_10681);
nor U13014 (N_13014,N_11903,N_10537);
nor U13015 (N_13015,N_9971,N_12111);
nand U13016 (N_13016,N_11704,N_9432);
and U13017 (N_13017,N_10266,N_11485);
or U13018 (N_13018,N_9493,N_10268);
nand U13019 (N_13019,N_11845,N_10041);
xor U13020 (N_13020,N_11996,N_9947);
and U13021 (N_13021,N_11513,N_11337);
nand U13022 (N_13022,N_9527,N_9693);
nand U13023 (N_13023,N_12052,N_11331);
nor U13024 (N_13024,N_11071,N_10363);
nand U13025 (N_13025,N_11121,N_10390);
or U13026 (N_13026,N_12387,N_12388);
nand U13027 (N_13027,N_9977,N_9773);
xnor U13028 (N_13028,N_11326,N_11939);
or U13029 (N_13029,N_12451,N_11460);
nor U13030 (N_13030,N_11866,N_11783);
nand U13031 (N_13031,N_12317,N_11111);
and U13032 (N_13032,N_9740,N_9387);
nor U13033 (N_13033,N_10487,N_10851);
nor U13034 (N_13034,N_11373,N_10267);
nand U13035 (N_13035,N_11635,N_10171);
nand U13036 (N_13036,N_11919,N_10553);
nor U13037 (N_13037,N_11314,N_11674);
xor U13038 (N_13038,N_9960,N_10585);
nand U13039 (N_13039,N_11275,N_11660);
xnor U13040 (N_13040,N_9945,N_9675);
nor U13041 (N_13041,N_10837,N_10610);
nor U13042 (N_13042,N_11239,N_10391);
nor U13043 (N_13043,N_9472,N_9386);
or U13044 (N_13044,N_10898,N_10991);
nor U13045 (N_13045,N_11295,N_10279);
nand U13046 (N_13046,N_10458,N_11926);
xnor U13047 (N_13047,N_10328,N_11280);
and U13048 (N_13048,N_12027,N_11355);
nand U13049 (N_13049,N_11659,N_9756);
nand U13050 (N_13050,N_11386,N_11315);
nand U13051 (N_13051,N_11285,N_10371);
xnor U13052 (N_13052,N_11782,N_10937);
and U13053 (N_13053,N_9984,N_11352);
or U13054 (N_13054,N_11655,N_11457);
nand U13055 (N_13055,N_10588,N_9907);
and U13056 (N_13056,N_9800,N_9406);
nand U13057 (N_13057,N_9384,N_9941);
xor U13058 (N_13058,N_9495,N_10531);
or U13059 (N_13059,N_10591,N_11544);
nor U13060 (N_13060,N_12493,N_10583);
nor U13061 (N_13061,N_11393,N_11751);
xor U13062 (N_13062,N_10590,N_9463);
or U13063 (N_13063,N_9755,N_12211);
and U13064 (N_13064,N_11523,N_10125);
xor U13065 (N_13065,N_11848,N_12204);
nor U13066 (N_13066,N_10033,N_9808);
nor U13067 (N_13067,N_9524,N_12276);
nand U13068 (N_13068,N_9613,N_10141);
and U13069 (N_13069,N_9434,N_9551);
xnor U13070 (N_13070,N_11203,N_12214);
and U13071 (N_13071,N_12481,N_11044);
or U13072 (N_13072,N_11962,N_10901);
xor U13073 (N_13073,N_9871,N_9509);
or U13074 (N_13074,N_10948,N_10376);
xor U13075 (N_13075,N_11968,N_9413);
or U13076 (N_13076,N_11821,N_12473);
or U13077 (N_13077,N_10761,N_11139);
or U13078 (N_13078,N_12196,N_11517);
xnor U13079 (N_13079,N_12411,N_9456);
xnor U13080 (N_13080,N_11868,N_9719);
or U13081 (N_13081,N_10290,N_10810);
or U13082 (N_13082,N_10099,N_10517);
xor U13083 (N_13083,N_10473,N_12360);
nor U13084 (N_13084,N_10245,N_12132);
or U13085 (N_13085,N_9581,N_11770);
xnor U13086 (N_13086,N_11738,N_9906);
nor U13087 (N_13087,N_11734,N_10453);
nand U13088 (N_13088,N_10521,N_11341);
nor U13089 (N_13089,N_12419,N_11599);
or U13090 (N_13090,N_9416,N_9643);
xnor U13091 (N_13091,N_11501,N_12140);
xor U13092 (N_13092,N_11693,N_10447);
or U13093 (N_13093,N_12010,N_11260);
nand U13094 (N_13094,N_10560,N_10700);
and U13095 (N_13095,N_11349,N_12394);
or U13096 (N_13096,N_9563,N_10175);
nand U13097 (N_13097,N_11085,N_11894);
xnor U13098 (N_13098,N_11863,N_12302);
nor U13099 (N_13099,N_12428,N_10943);
nor U13100 (N_13100,N_9751,N_10182);
or U13101 (N_13101,N_10361,N_10683);
nor U13102 (N_13102,N_12306,N_9437);
xor U13103 (N_13103,N_9648,N_12153);
xor U13104 (N_13104,N_12065,N_11060);
nand U13105 (N_13105,N_11872,N_12108);
nor U13106 (N_13106,N_9832,N_11067);
and U13107 (N_13107,N_12127,N_10086);
nand U13108 (N_13108,N_11556,N_10365);
nor U13109 (N_13109,N_9951,N_12131);
xor U13110 (N_13110,N_11256,N_11824);
nor U13111 (N_13111,N_9582,N_10139);
and U13112 (N_13112,N_10373,N_11557);
nor U13113 (N_13113,N_10085,N_12016);
nand U13114 (N_13114,N_10183,N_11233);
nand U13115 (N_13115,N_9955,N_10865);
or U13116 (N_13116,N_10410,N_12371);
and U13117 (N_13117,N_10730,N_12030);
nand U13118 (N_13118,N_11807,N_10788);
and U13119 (N_13119,N_9829,N_9901);
nand U13120 (N_13120,N_11965,N_9946);
or U13121 (N_13121,N_12275,N_9540);
nand U13122 (N_13122,N_11210,N_9611);
nor U13123 (N_13123,N_9869,N_11266);
or U13124 (N_13124,N_10314,N_12430);
nor U13125 (N_13125,N_12368,N_9777);
nand U13126 (N_13126,N_11492,N_11880);
or U13127 (N_13127,N_10366,N_10435);
nor U13128 (N_13128,N_11945,N_12406);
nor U13129 (N_13129,N_9628,N_10349);
xnor U13130 (N_13130,N_10048,N_12488);
xnor U13131 (N_13131,N_9511,N_9395);
nor U13132 (N_13132,N_10535,N_11521);
nand U13133 (N_13133,N_10508,N_12120);
nor U13134 (N_13134,N_11290,N_9949);
and U13135 (N_13135,N_10624,N_12362);
nor U13136 (N_13136,N_10383,N_10527);
nand U13137 (N_13137,N_11722,N_11127);
nand U13138 (N_13138,N_12086,N_10239);
xor U13139 (N_13139,N_10010,N_10676);
or U13140 (N_13140,N_11357,N_11181);
or U13141 (N_13141,N_12223,N_11809);
or U13142 (N_13142,N_12420,N_11304);
nor U13143 (N_13143,N_10606,N_11183);
or U13144 (N_13144,N_10939,N_11841);
nand U13145 (N_13145,N_11145,N_9452);
or U13146 (N_13146,N_10793,N_11030);
or U13147 (N_13147,N_10297,N_11878);
or U13148 (N_13148,N_12268,N_10193);
nor U13149 (N_13149,N_10607,N_12415);
nand U13150 (N_13150,N_10073,N_12438);
or U13151 (N_13151,N_12090,N_9614);
and U13152 (N_13152,N_11247,N_10958);
nor U13153 (N_13153,N_10707,N_10983);
nor U13154 (N_13154,N_9572,N_10747);
and U13155 (N_13155,N_12236,N_11430);
nand U13156 (N_13156,N_11499,N_11379);
or U13157 (N_13157,N_10881,N_9781);
xnor U13158 (N_13158,N_12298,N_11678);
xnor U13159 (N_13159,N_10644,N_11242);
and U13160 (N_13160,N_10502,N_10096);
or U13161 (N_13161,N_10826,N_9922);
nor U13162 (N_13162,N_12169,N_9398);
and U13163 (N_13163,N_11369,N_10348);
and U13164 (N_13164,N_11426,N_9764);
and U13165 (N_13165,N_10575,N_10798);
nand U13166 (N_13166,N_11104,N_11036);
nand U13167 (N_13167,N_11898,N_9430);
and U13168 (N_13168,N_10427,N_11409);
xnor U13169 (N_13169,N_11830,N_12265);
nor U13170 (N_13170,N_9531,N_11570);
xor U13171 (N_13171,N_11991,N_10185);
and U13172 (N_13172,N_10543,N_10395);
and U13173 (N_13173,N_11211,N_12460);
or U13174 (N_13174,N_9793,N_10874);
xor U13175 (N_13175,N_12331,N_10856);
nand U13176 (N_13176,N_10251,N_10005);
nand U13177 (N_13177,N_9522,N_10556);
and U13178 (N_13178,N_10117,N_10023);
or U13179 (N_13179,N_10965,N_10491);
nor U13180 (N_13180,N_9433,N_12195);
or U13181 (N_13181,N_11963,N_10408);
xor U13182 (N_13182,N_9727,N_10287);
nand U13183 (N_13183,N_9866,N_12464);
and U13184 (N_13184,N_11421,N_12234);
xnor U13185 (N_13185,N_10211,N_12364);
xnor U13186 (N_13186,N_12071,N_11905);
xnor U13187 (N_13187,N_11035,N_12014);
xor U13188 (N_13188,N_11507,N_9631);
xor U13189 (N_13189,N_9425,N_10327);
nor U13190 (N_13190,N_11283,N_11748);
nor U13191 (N_13191,N_10821,N_11453);
nor U13192 (N_13192,N_11593,N_11699);
nor U13193 (N_13193,N_11663,N_11961);
nor U13194 (N_13194,N_10356,N_10561);
and U13195 (N_13195,N_11595,N_12457);
xor U13196 (N_13196,N_11433,N_10011);
and U13197 (N_13197,N_11236,N_11020);
or U13198 (N_13198,N_11855,N_10293);
or U13199 (N_13199,N_11787,N_9795);
nand U13200 (N_13200,N_12222,N_10417);
and U13201 (N_13201,N_11546,N_10780);
xnor U13202 (N_13202,N_11927,N_11450);
or U13203 (N_13203,N_10167,N_10460);
or U13204 (N_13204,N_10178,N_11817);
and U13205 (N_13205,N_12230,N_12209);
or U13206 (N_13206,N_10703,N_9566);
or U13207 (N_13207,N_12233,N_11459);
nand U13208 (N_13208,N_9515,N_11175);
nor U13209 (N_13209,N_11431,N_11092);
and U13210 (N_13210,N_9748,N_11325);
or U13211 (N_13211,N_10004,N_9741);
and U13212 (N_13212,N_11113,N_11650);
xnor U13213 (N_13213,N_11380,N_10828);
and U13214 (N_13214,N_11689,N_10108);
and U13215 (N_13215,N_11646,N_11975);
nor U13216 (N_13216,N_12139,N_10723);
or U13217 (N_13217,N_11102,N_10030);
nand U13218 (N_13218,N_10625,N_10809);
and U13219 (N_13219,N_11312,N_11766);
nand U13220 (N_13220,N_10667,N_10042);
and U13221 (N_13221,N_9873,N_11534);
nand U13222 (N_13222,N_10671,N_10276);
and U13223 (N_13223,N_12183,N_12432);
nor U13224 (N_13224,N_9974,N_9577);
nand U13225 (N_13225,N_12072,N_9842);
xnor U13226 (N_13226,N_11026,N_10663);
nand U13227 (N_13227,N_12046,N_10794);
nand U13228 (N_13228,N_9667,N_9537);
or U13229 (N_13229,N_9894,N_11110);
xor U13230 (N_13230,N_11012,N_11977);
nand U13231 (N_13231,N_11383,N_11254);
or U13232 (N_13232,N_11080,N_9485);
nor U13233 (N_13233,N_10771,N_11240);
xor U13234 (N_13234,N_10047,N_12144);
nand U13235 (N_13235,N_10660,N_11016);
nand U13236 (N_13236,N_10068,N_10154);
or U13237 (N_13237,N_12128,N_10841);
nand U13238 (N_13238,N_12410,N_12285);
nor U13239 (N_13239,N_11310,N_10847);
and U13240 (N_13240,N_11826,N_9760);
nor U13241 (N_13241,N_12354,N_11056);
nand U13242 (N_13242,N_12495,N_10058);
or U13243 (N_13243,N_10923,N_10611);
xor U13244 (N_13244,N_9862,N_10831);
and U13245 (N_13245,N_10067,N_12106);
or U13246 (N_13246,N_10029,N_10511);
nand U13247 (N_13247,N_9604,N_10946);
or U13248 (N_13248,N_10474,N_11741);
nand U13249 (N_13249,N_11714,N_10493);
xnor U13250 (N_13250,N_12322,N_9695);
nand U13251 (N_13251,N_9550,N_9911);
nand U13252 (N_13252,N_12486,N_10718);
and U13253 (N_13253,N_10110,N_11864);
and U13254 (N_13254,N_12176,N_12076);
nand U13255 (N_13255,N_10295,N_9747);
and U13256 (N_13256,N_9890,N_11456);
nand U13257 (N_13257,N_11565,N_10107);
or U13258 (N_13258,N_12047,N_12329);
and U13259 (N_13259,N_10770,N_10573);
nand U13260 (N_13260,N_12113,N_10727);
xor U13261 (N_13261,N_9978,N_12465);
nand U13262 (N_13262,N_9778,N_11288);
xnor U13263 (N_13263,N_12213,N_12232);
nor U13264 (N_13264,N_10928,N_10979);
or U13265 (N_13265,N_11948,N_10580);
nor U13266 (N_13266,N_10419,N_10879);
nand U13267 (N_13267,N_12448,N_10406);
nor U13268 (N_13268,N_9410,N_10236);
and U13269 (N_13269,N_12013,N_11371);
and U13270 (N_13270,N_9539,N_10605);
nor U13271 (N_13271,N_10146,N_11890);
nor U13272 (N_13272,N_10078,N_9686);
nand U13273 (N_13273,N_11311,N_12427);
or U13274 (N_13274,N_9455,N_9926);
nor U13275 (N_13275,N_10910,N_10899);
nor U13276 (N_13276,N_12499,N_11142);
and U13277 (N_13277,N_10633,N_9663);
nand U13278 (N_13278,N_11487,N_11602);
nand U13279 (N_13279,N_11395,N_9860);
xor U13280 (N_13280,N_9843,N_9450);
xor U13281 (N_13281,N_9952,N_11225);
or U13282 (N_13282,N_11780,N_11631);
nor U13283 (N_13283,N_10159,N_12421);
nor U13284 (N_13284,N_11106,N_10959);
nor U13285 (N_13285,N_11959,N_9826);
nor U13286 (N_13286,N_9724,N_12434);
nand U13287 (N_13287,N_9636,N_10456);
nand U13288 (N_13288,N_10536,N_10018);
nand U13289 (N_13289,N_10579,N_10061);
nor U13290 (N_13290,N_10574,N_9627);
xnor U13291 (N_13291,N_12475,N_11277);
nand U13292 (N_13292,N_11823,N_10329);
nor U13293 (N_13293,N_11525,N_9966);
xor U13294 (N_13294,N_12033,N_9444);
or U13295 (N_13295,N_11105,N_10709);
xnor U13296 (N_13296,N_11005,N_11117);
or U13297 (N_13297,N_10744,N_12148);
or U13298 (N_13298,N_9817,N_11902);
or U13299 (N_13299,N_11216,N_11231);
xnor U13300 (N_13300,N_9596,N_9385);
nand U13301 (N_13301,N_9478,N_9729);
nor U13302 (N_13302,N_10070,N_12107);
and U13303 (N_13303,N_12485,N_10063);
nand U13304 (N_13304,N_10480,N_9762);
and U13305 (N_13305,N_11051,N_10092);
and U13306 (N_13306,N_10942,N_11438);
nand U13307 (N_13307,N_10206,N_10614);
or U13308 (N_13308,N_12036,N_11690);
xnor U13309 (N_13309,N_11190,N_9981);
xnor U13310 (N_13310,N_10231,N_11164);
or U13311 (N_13311,N_10503,N_9474);
nand U13312 (N_13312,N_11904,N_9813);
xnor U13313 (N_13313,N_11574,N_12130);
or U13314 (N_13314,N_9440,N_9672);
or U13315 (N_13315,N_10388,N_10127);
nand U13316 (N_13316,N_11083,N_10149);
or U13317 (N_13317,N_9436,N_9685);
nor U13318 (N_13318,N_10440,N_10177);
nand U13319 (N_13319,N_11098,N_12099);
nand U13320 (N_13320,N_11265,N_9661);
xnor U13321 (N_13321,N_10151,N_10446);
or U13322 (N_13322,N_11594,N_11691);
xnor U13323 (N_13323,N_9612,N_9499);
or U13324 (N_13324,N_10914,N_11936);
xnor U13325 (N_13325,N_12172,N_11222);
and U13326 (N_13326,N_11388,N_9811);
and U13327 (N_13327,N_11811,N_10210);
and U13328 (N_13328,N_10463,N_11483);
or U13329 (N_13329,N_9917,N_10163);
nand U13330 (N_13330,N_11701,N_12263);
xnor U13331 (N_13331,N_11412,N_9570);
and U13332 (N_13332,N_9601,N_11270);
nor U13333 (N_13333,N_11360,N_9732);
or U13334 (N_13334,N_10002,N_12441);
xnor U13335 (N_13335,N_10034,N_10394);
and U13336 (N_13336,N_9881,N_11068);
and U13337 (N_13337,N_9857,N_10716);
xnor U13338 (N_13338,N_10260,N_10642);
or U13339 (N_13339,N_11298,N_10961);
nor U13340 (N_13340,N_12121,N_11061);
nor U13341 (N_13341,N_9825,N_10893);
or U13342 (N_13342,N_11053,N_11795);
nor U13343 (N_13343,N_10980,N_12262);
and U13344 (N_13344,N_10118,N_10819);
nor U13345 (N_13345,N_10996,N_9713);
xnor U13346 (N_13346,N_9700,N_10037);
nand U13347 (N_13347,N_11390,N_10324);
nand U13348 (N_13348,N_11542,N_12417);
and U13349 (N_13349,N_12471,N_10368);
and U13350 (N_13350,N_11141,N_9767);
nor U13351 (N_13351,N_12210,N_11917);
nand U13352 (N_13352,N_11023,N_9914);
and U13353 (N_13353,N_12066,N_9622);
nor U13354 (N_13354,N_11668,N_10890);
or U13355 (N_13355,N_12181,N_10956);
nor U13356 (N_13356,N_12435,N_11406);
or U13357 (N_13357,N_11581,N_12470);
xnor U13358 (N_13358,N_11129,N_11424);
xor U13359 (N_13359,N_10411,N_11707);
or U13360 (N_13360,N_11206,N_9943);
or U13361 (N_13361,N_9497,N_10924);
nand U13362 (N_13362,N_11537,N_10201);
nand U13363 (N_13363,N_12437,N_9484);
xnor U13364 (N_13364,N_12119,N_10524);
nor U13365 (N_13365,N_9670,N_9487);
nor U13366 (N_13366,N_10254,N_11990);
nand U13367 (N_13367,N_9753,N_11955);
or U13368 (N_13368,N_12365,N_9923);
xor U13369 (N_13369,N_12040,N_12295);
nor U13370 (N_13370,N_11788,N_10571);
xnor U13371 (N_13371,N_10469,N_11297);
and U13372 (N_13372,N_10213,N_10544);
xor U13373 (N_13373,N_10749,N_10335);
nand U13374 (N_13374,N_10145,N_9786);
xor U13375 (N_13375,N_11584,N_10197);
or U13376 (N_13376,N_9589,N_10931);
and U13377 (N_13377,N_12291,N_11306);
or U13378 (N_13378,N_12439,N_9957);
or U13379 (N_13379,N_10842,N_9738);
nor U13380 (N_13380,N_9445,N_9725);
nor U13381 (N_13381,N_9491,N_9618);
or U13382 (N_13382,N_11091,N_11428);
nor U13383 (N_13383,N_9630,N_10442);
xor U13384 (N_13384,N_11258,N_11730);
xor U13385 (N_13385,N_9815,N_10367);
and U13386 (N_13386,N_10587,N_10776);
or U13387 (N_13387,N_10854,N_11799);
and U13388 (N_13388,N_12042,N_12056);
nor U13389 (N_13389,N_10868,N_12102);
and U13390 (N_13390,N_11148,N_11754);
xnor U13391 (N_13391,N_12069,N_12227);
nand U13392 (N_13392,N_10596,N_9546);
nand U13393 (N_13393,N_10850,N_11664);
nor U13394 (N_13394,N_11654,N_10015);
or U13395 (N_13395,N_11375,N_9982);
nor U13396 (N_13396,N_12212,N_11540);
nand U13397 (N_13397,N_10275,N_11489);
nor U13398 (N_13398,N_10013,N_11269);
nor U13399 (N_13399,N_9838,N_10604);
nor U13400 (N_13400,N_9513,N_12174);
xnor U13401 (N_13401,N_12349,N_9516);
xnor U13402 (N_13402,N_10997,N_12190);
or U13403 (N_13403,N_9506,N_11316);
nor U13404 (N_13404,N_11132,N_9620);
nor U13405 (N_13405,N_10782,N_12059);
nand U13406 (N_13406,N_12320,N_11605);
nor U13407 (N_13407,N_9482,N_9391);
or U13408 (N_13408,N_11791,N_11184);
nand U13409 (N_13409,N_10387,N_10316);
nor U13410 (N_13410,N_10264,N_11228);
nand U13411 (N_13411,N_12161,N_10557);
nand U13412 (N_13412,N_11626,N_9930);
nand U13413 (N_13413,N_10679,N_9900);
nor U13414 (N_13414,N_9541,N_12396);
nor U13415 (N_13415,N_11789,N_10795);
nor U13416 (N_13416,N_9635,N_9655);
xor U13417 (N_13417,N_11784,N_12367);
and U13418 (N_13418,N_11638,N_11918);
nor U13419 (N_13419,N_10693,N_9459);
or U13420 (N_13420,N_9939,N_10971);
xnor U13421 (N_13421,N_11014,N_10752);
xnor U13422 (N_13422,N_10773,N_9567);
nor U13423 (N_13423,N_10089,N_9591);
nand U13424 (N_13424,N_12305,N_11681);
and U13425 (N_13425,N_9839,N_11229);
or U13426 (N_13426,N_11785,N_9789);
xnor U13427 (N_13427,N_11726,N_12466);
xnor U13428 (N_13428,N_11972,N_9749);
xnor U13429 (N_13429,N_9584,N_10441);
nor U13430 (N_13430,N_10222,N_11600);
nor U13431 (N_13431,N_10849,N_11077);
nand U13432 (N_13432,N_10292,N_11913);
xnor U13433 (N_13433,N_10484,N_10836);
and U13434 (N_13434,N_11946,N_10187);
nor U13435 (N_13435,N_11661,N_10907);
or U13436 (N_13436,N_11096,N_11744);
or U13437 (N_13437,N_10696,N_10765);
or U13438 (N_13438,N_10646,N_10603);
nand U13439 (N_13439,N_10352,N_11201);
or U13440 (N_13440,N_9476,N_12051);
xnor U13441 (N_13441,N_10589,N_9598);
and U13442 (N_13442,N_12217,N_10097);
xnor U13443 (N_13443,N_12476,N_10464);
nor U13444 (N_13444,N_11810,N_10165);
nand U13445 (N_13445,N_12240,N_10494);
nand U13446 (N_13446,N_11418,N_10516);
or U13447 (N_13447,N_11685,N_11187);
and U13448 (N_13448,N_9863,N_11486);
nand U13449 (N_13449,N_11339,N_12374);
and U13450 (N_13450,N_11527,N_11531);
xnor U13451 (N_13451,N_11158,N_11033);
xor U13452 (N_13452,N_11214,N_10219);
nor U13453 (N_13453,N_12098,N_11840);
or U13454 (N_13454,N_10303,N_10160);
nor U13455 (N_13455,N_9435,N_12401);
and U13456 (N_13456,N_10562,N_9585);
or U13457 (N_13457,N_9814,N_10686);
nand U13458 (N_13458,N_11781,N_10756);
nand U13459 (N_13459,N_12343,N_11095);
nor U13460 (N_13460,N_10581,N_12084);
xor U13461 (N_13461,N_12356,N_10243);
or U13462 (N_13462,N_9496,N_10804);
xor U13463 (N_13463,N_11416,N_11153);
nand U13464 (N_13464,N_11262,N_11502);
or U13465 (N_13465,N_11937,N_11592);
nand U13466 (N_13466,N_10568,N_10286);
nand U13467 (N_13467,N_12032,N_11983);
and U13468 (N_13468,N_12407,N_10081);
xnor U13469 (N_13469,N_9928,N_11985);
nand U13470 (N_13470,N_10320,N_9574);
nor U13471 (N_13471,N_11282,N_11474);
or U13472 (N_13472,N_12250,N_9594);
xor U13473 (N_13473,N_9743,N_9761);
nor U13474 (N_13474,N_11329,N_10838);
nor U13475 (N_13475,N_11467,N_11138);
or U13476 (N_13476,N_10120,N_9556);
or U13477 (N_13477,N_12497,N_11070);
nor U13478 (N_13478,N_9714,N_11215);
nor U13479 (N_13479,N_11377,N_10199);
and U13480 (N_13480,N_10358,N_12284);
nand U13481 (N_13481,N_11713,N_9834);
and U13482 (N_13482,N_11947,N_9735);
xor U13483 (N_13483,N_10548,N_9414);
nor U13484 (N_13484,N_9534,N_10143);
and U13485 (N_13485,N_9377,N_11116);
nand U13486 (N_13486,N_10294,N_9848);
xor U13487 (N_13487,N_10424,N_9588);
xnor U13488 (N_13488,N_10859,N_9969);
and U13489 (N_13489,N_10726,N_11131);
nor U13490 (N_13490,N_10142,N_10567);
nor U13491 (N_13491,N_11954,N_10921);
or U13492 (N_13492,N_11328,N_12395);
nor U13493 (N_13493,N_11143,N_11335);
xnor U13494 (N_13494,N_9659,N_9654);
nand U13495 (N_13495,N_12186,N_10121);
xor U13496 (N_13496,N_12068,N_11869);
nand U13497 (N_13497,N_10930,N_9877);
or U13498 (N_13498,N_9419,N_9448);
or U13499 (N_13499,N_10918,N_12300);
or U13500 (N_13500,N_9934,N_10694);
or U13501 (N_13501,N_10202,N_9405);
or U13502 (N_13502,N_11508,N_11732);
or U13503 (N_13503,N_10870,N_9458);
nor U13504 (N_13504,N_12171,N_10721);
or U13505 (N_13505,N_10582,N_11876);
nand U13506 (N_13506,N_9637,N_11197);
and U13507 (N_13507,N_10616,N_9514);
xnor U13508 (N_13508,N_11637,N_10966);
nand U13509 (N_13509,N_9396,N_12399);
and U13510 (N_13510,N_10685,N_10677);
or U13511 (N_13511,N_9408,N_12185);
or U13512 (N_13512,N_11043,N_10443);
xor U13513 (N_13513,N_11642,N_11639);
or U13514 (N_13514,N_12352,N_10978);
or U13515 (N_13515,N_10375,N_9603);
nand U13516 (N_13516,N_9853,N_10706);
xor U13517 (N_13517,N_10895,N_10496);
and U13518 (N_13518,N_11590,N_12248);
and U13519 (N_13519,N_12267,N_12182);
nor U13520 (N_13520,N_10763,N_9411);
and U13521 (N_13521,N_10301,N_12034);
xor U13522 (N_13522,N_12048,N_11052);
nor U13523 (N_13523,N_10697,N_10684);
or U13524 (N_13524,N_12159,N_11715);
or U13525 (N_13525,N_12445,N_10173);
nor U13526 (N_13526,N_9816,N_11494);
and U13527 (N_13527,N_10153,N_12237);
and U13528 (N_13528,N_10822,N_11119);
and U13529 (N_13529,N_12405,N_10241);
and U13530 (N_13530,N_9562,N_11209);
and U13531 (N_13531,N_11137,N_11252);
and U13532 (N_13532,N_11074,N_11444);
and U13533 (N_13533,N_9925,N_11165);
or U13534 (N_13534,N_11273,N_11130);
xnor U13535 (N_13535,N_11665,N_9916);
xor U13536 (N_13536,N_10100,N_9827);
nor U13537 (N_13537,N_11558,N_12480);
xor U13538 (N_13538,N_11862,N_12000);
xor U13539 (N_13539,N_11376,N_10087);
xnor U13540 (N_13540,N_11836,N_10242);
xnor U13541 (N_13541,N_11101,N_11900);
nand U13542 (N_13542,N_10166,N_10088);
nor U13543 (N_13543,N_12468,N_10546);
and U13544 (N_13544,N_9870,N_11506);
xnor U13545 (N_13545,N_12077,N_10739);
or U13546 (N_13546,N_9964,N_9431);
nor U13547 (N_13547,N_9953,N_10664);
nand U13548 (N_13548,N_10584,N_9932);
or U13549 (N_13549,N_12303,N_10305);
or U13550 (N_13550,N_9712,N_9666);
xor U13551 (N_13551,N_10053,N_10071);
nor U13552 (N_13552,N_11232,N_12126);
or U13553 (N_13553,N_9400,N_10150);
nand U13554 (N_13554,N_9788,N_10402);
nand U13555 (N_13555,N_9983,N_10481);
or U13556 (N_13556,N_10632,N_11064);
nand U13557 (N_13557,N_11398,N_11324);
nand U13558 (N_13558,N_11510,N_12484);
xnor U13559 (N_13559,N_9535,N_10737);
and U13560 (N_13560,N_9483,N_12220);
or U13561 (N_13561,N_11452,N_9502);
nor U13562 (N_13562,N_11931,N_10170);
or U13563 (N_13563,N_9701,N_12482);
nand U13564 (N_13564,N_11739,N_10482);
or U13565 (N_13565,N_10425,N_12061);
xnor U13566 (N_13566,N_9381,N_11392);
nand U13567 (N_13567,N_11769,N_11790);
nor U13568 (N_13568,N_9963,N_10595);
or U13569 (N_13569,N_9647,N_10705);
or U13570 (N_13570,N_10186,N_10467);
xor U13571 (N_13571,N_10787,N_11912);
and U13572 (N_13572,N_11923,N_9903);
nand U13573 (N_13573,N_12330,N_12259);
or U13574 (N_13574,N_10786,N_12202);
nor U13575 (N_13575,N_10369,N_11813);
nand U13576 (N_13576,N_12404,N_10103);
and U13577 (N_13577,N_10310,N_10800);
xor U13578 (N_13578,N_11943,N_10343);
nand U13579 (N_13579,N_11342,N_10968);
or U13580 (N_13580,N_12472,N_11634);
nor U13581 (N_13581,N_11686,N_11401);
and U13582 (N_13582,N_12143,N_9417);
nor U13583 (N_13583,N_11924,N_9595);
xor U13584 (N_13584,N_10869,N_12490);
nand U13585 (N_13585,N_11509,N_12004);
and U13586 (N_13586,N_10843,N_9845);
nor U13587 (N_13587,N_12011,N_9438);
or U13588 (N_13588,N_11372,N_11446);
nand U13589 (N_13589,N_10541,N_10905);
or U13590 (N_13590,N_10046,N_9851);
xor U13591 (N_13591,N_11612,N_10654);
and U13592 (N_13592,N_11498,N_10123);
and U13593 (N_13593,N_10917,N_11034);
nor U13594 (N_13594,N_10609,N_10720);
nand U13595 (N_13595,N_9679,N_10661);
xnor U13596 (N_13596,N_11995,N_12278);
or U13597 (N_13597,N_12091,N_12294);
and U13598 (N_13598,N_10631,N_9504);
or U13599 (N_13599,N_11886,N_11462);
or U13600 (N_13600,N_10711,N_9580);
xnor U13601 (N_13601,N_11346,N_10207);
xnor U13602 (N_13602,N_11773,N_9979);
and U13603 (N_13603,N_11656,N_10577);
or U13604 (N_13604,N_9428,N_10653);
or U13605 (N_13605,N_10003,N_11292);
and U13606 (N_13606,N_12397,N_9996);
and U13607 (N_13607,N_9790,N_9553);
and U13608 (N_13608,N_11940,N_9692);
xor U13609 (N_13609,N_10353,N_9639);
and U13610 (N_13610,N_10179,N_11615);
or U13611 (N_13611,N_10471,N_10336);
nor U13612 (N_13612,N_11167,N_12443);
nor U13613 (N_13613,N_9443,N_10378);
or U13614 (N_13614,N_10962,N_10319);
nor U13615 (N_13615,N_11630,N_9706);
xor U13616 (N_13616,N_10374,N_10911);
or U13617 (N_13617,N_12037,N_11268);
nand U13618 (N_13618,N_9803,N_11301);
xnor U13619 (N_13619,N_10429,N_12085);
or U13620 (N_13620,N_10347,N_10872);
nor U13621 (N_13621,N_12078,N_11703);
nor U13622 (N_13622,N_10618,N_12136);
xor U13623 (N_13623,N_10986,N_11835);
and U13624 (N_13624,N_12020,N_11564);
and U13625 (N_13625,N_10514,N_12283);
nand U13626 (N_13626,N_10712,N_10551);
or U13627 (N_13627,N_12469,N_10401);
nand U13628 (N_13628,N_12301,N_10331);
or U13629 (N_13629,N_9828,N_11244);
nor U13630 (N_13630,N_10781,N_11454);
xnor U13631 (N_13631,N_12224,N_11928);
or U13632 (N_13632,N_12408,N_11998);
or U13633 (N_13633,N_11213,N_9465);
and U13634 (N_13634,N_12442,N_9650);
or U13635 (N_13635,N_11700,N_11746);
nand U13636 (N_13636,N_11442,N_12332);
and U13637 (N_13637,N_10191,N_11257);
nand U13638 (N_13638,N_11100,N_9824);
or U13639 (N_13639,N_10077,N_10433);
nor U13640 (N_13640,N_11220,N_12398);
xor U13641 (N_13641,N_10741,N_9402);
and U13642 (N_13642,N_12208,N_11916);
nor U13643 (N_13643,N_11473,N_10688);
xnor U13644 (N_13644,N_10064,N_11579);
nand U13645 (N_13645,N_12207,N_10012);
nor U13646 (N_13646,N_11774,N_10102);
nand U13647 (N_13647,N_11645,N_10858);
nand U13648 (N_13648,N_10668,N_10759);
nor U13649 (N_13649,N_11133,N_11317);
and U13650 (N_13650,N_10601,N_12012);
nor U13651 (N_13651,N_11482,N_11994);
nand U13652 (N_13652,N_10129,N_12147);
or U13653 (N_13653,N_10913,N_11794);
or U13654 (N_13654,N_10529,N_9809);
nand U13655 (N_13655,N_11208,N_9651);
or U13656 (N_13656,N_11179,N_12304);
or U13657 (N_13657,N_10523,N_10217);
xnor U13658 (N_13658,N_10909,N_11989);
nand U13659 (N_13659,N_9933,N_12019);
or U13660 (N_13660,N_10181,N_9401);
nand U13661 (N_13661,N_10176,N_11267);
nor U13662 (N_13662,N_10342,N_12239);
or U13663 (N_13663,N_11368,N_11072);
xnor U13664 (N_13664,N_10522,N_11702);
or U13665 (N_13665,N_10285,N_10325);
and U13666 (N_13666,N_11536,N_11099);
nor U13667 (N_13667,N_10196,N_10884);
or U13668 (N_13668,N_9876,N_12163);
nand U13669 (N_13669,N_11170,N_11434);
nor U13670 (N_13670,N_11596,N_10915);
xor U13671 (N_13671,N_10132,N_11204);
or U13672 (N_13672,N_11910,N_11648);
nor U13673 (N_13673,N_11159,N_9394);
nand U13674 (N_13674,N_10998,N_11322);
nand U13675 (N_13675,N_11054,N_9956);
and U13676 (N_13676,N_11750,N_11885);
nor U13677 (N_13677,N_12200,N_12064);
nor U13678 (N_13678,N_11358,N_9403);
and U13679 (N_13679,N_9468,N_12266);
nand U13680 (N_13680,N_10263,N_10532);
nor U13681 (N_13681,N_11207,N_10317);
or U13682 (N_13682,N_11867,N_10783);
xnor U13683 (N_13683,N_11496,N_11827);
and U13684 (N_13684,N_9525,N_10345);
xnor U13685 (N_13685,N_11075,N_10248);
nor U13686 (N_13686,N_10479,N_10967);
and U13687 (N_13687,N_10039,N_11838);
xnor U13688 (N_13688,N_11481,N_12193);
xnor U13689 (N_13689,N_11816,N_11154);
nor U13690 (N_13690,N_11548,N_11114);
or U13691 (N_13691,N_11146,N_11356);
and U13692 (N_13692,N_11619,N_10203);
nand U13693 (N_13693,N_12006,N_10381);
xor U13694 (N_13694,N_12017,N_11829);
or U13695 (N_13695,N_11188,N_10801);
nand U13696 (N_13696,N_11727,N_10226);
nand U13697 (N_13697,N_12292,N_10779);
and U13698 (N_13698,N_9389,N_10220);
nand U13699 (N_13699,N_11378,N_10656);
nor U13700 (N_13700,N_9587,N_12205);
xor U13701 (N_13701,N_12137,N_12156);
nand U13702 (N_13702,N_9593,N_11387);
nand U13703 (N_13703,N_10748,N_11874);
nand U13704 (N_13704,N_10452,N_10380);
or U13705 (N_13705,N_11384,N_11089);
xor U13706 (N_13706,N_9460,N_12424);
and U13707 (N_13707,N_10731,N_11710);
nand U13708 (N_13708,N_10119,N_10364);
xnor U13709 (N_13709,N_9780,N_11518);
nor U13710 (N_13710,N_9507,N_12088);
nor U13711 (N_13711,N_12189,N_10530);
nand U13712 (N_13712,N_11359,N_10056);
nand U13713 (N_13713,N_11348,N_9805);
and U13714 (N_13714,N_12381,N_9997);
and U13715 (N_13715,N_12379,N_12142);
nand U13716 (N_13716,N_10407,N_9674);
or U13717 (N_13717,N_12403,N_12246);
xor U13718 (N_13718,N_10926,N_12238);
nand U13719 (N_13719,N_9439,N_11849);
nand U13720 (N_13720,N_10878,N_11893);
or U13721 (N_13721,N_12199,N_10296);
and U13722 (N_13722,N_10655,N_11967);
nor U13723 (N_13723,N_12418,N_11284);
or U13724 (N_13724,N_10862,N_11806);
nor U13725 (N_13725,N_11733,N_11367);
or U13726 (N_13726,N_12080,N_11832);
or U13727 (N_13727,N_11477,N_11323);
xnor U13728 (N_13728,N_9664,N_9905);
xor U13729 (N_13729,N_12389,N_12242);
xor U13730 (N_13730,N_9763,N_12063);
or U13731 (N_13731,N_10977,N_9644);
nor U13732 (N_13732,N_11008,N_9689);
nor U13733 (N_13733,N_10738,N_10951);
xnor U13734 (N_13734,N_9442,N_10448);
and U13735 (N_13735,N_10188,N_9868);
and U13736 (N_13736,N_11427,N_11351);
nand U13737 (N_13737,N_11245,N_9602);
and U13738 (N_13738,N_9575,N_11109);
and U13739 (N_13739,N_9668,N_11616);
nand U13740 (N_13740,N_12162,N_11993);
xor U13741 (N_13741,N_9473,N_12025);
xnor U13742 (N_13742,N_10486,N_9699);
or U13743 (N_13743,N_12009,N_10659);
and U13744 (N_13744,N_10113,N_10122);
xor U13745 (N_13745,N_10510,N_10434);
or U13746 (N_13746,N_11712,N_11953);
and U13747 (N_13747,N_9837,N_11248);
nor U13748 (N_13748,N_9616,N_11293);
nor U13749 (N_13749,N_11160,N_10973);
or U13750 (N_13750,N_9673,N_11057);
xor U13751 (N_13751,N_12494,N_10049);
nand U13752 (N_13752,N_11932,N_9846);
nand U13753 (N_13753,N_10597,N_10225);
xnor U13754 (N_13754,N_10815,N_11066);
or U13755 (N_13755,N_10732,N_11949);
or U13756 (N_13756,N_9959,N_12093);
or U13757 (N_13757,N_9634,N_9865);
nor U13758 (N_13758,N_11263,N_10864);
nand U13759 (N_13759,N_9520,N_9660);
xor U13760 (N_13760,N_10277,N_10501);
or U13761 (N_13761,N_10934,N_9715);
nand U13762 (N_13762,N_10205,N_9742);
xor U13763 (N_13763,N_11760,N_10834);
or U13764 (N_13764,N_11705,N_10083);
and U13765 (N_13765,N_11140,N_11614);
xor U13766 (N_13766,N_11241,N_11852);
nand U13767 (N_13767,N_9475,N_11764);
nand U13768 (N_13768,N_9980,N_11711);
nor U13769 (N_13769,N_11842,N_10054);
nor U13770 (N_13770,N_11858,N_10372);
nor U13771 (N_13771,N_9479,N_11303);
nor U13772 (N_13772,N_9583,N_11986);
or U13773 (N_13773,N_10845,N_10506);
or U13774 (N_13774,N_9858,N_10355);
and U13775 (N_13775,N_10115,N_11195);
or U13776 (N_13776,N_11559,N_12392);
and U13777 (N_13777,N_11013,N_11532);
and U13778 (N_13778,N_9730,N_12455);
nor U13779 (N_13779,N_9645,N_12049);
nand U13780 (N_13780,N_11578,N_11010);
and U13781 (N_13781,N_10880,N_10184);
nand U13782 (N_13782,N_11607,N_9882);
or U13783 (N_13783,N_10397,N_9972);
and U13784 (N_13784,N_10500,N_10799);
xnor U13785 (N_13785,N_12180,N_11354);
or U13786 (N_13786,N_10662,N_11086);
xnor U13787 (N_13787,N_10526,N_11200);
nand U13788 (N_13788,N_12005,N_10757);
xnor U13789 (N_13789,N_12188,N_9758);
nand U13790 (N_13790,N_11882,N_10422);
nor U13791 (N_13791,N_11128,N_10148);
xor U13792 (N_13792,N_11021,N_10796);
xnor U13793 (N_13793,N_12079,N_10970);
and U13794 (N_13794,N_12496,N_9736);
or U13795 (N_13795,N_10769,N_10223);
or U13796 (N_13796,N_9462,N_11468);
nor U13797 (N_13797,N_9543,N_9619);
nand U13798 (N_13798,N_11118,N_9423);
nor U13799 (N_13799,N_12117,N_11568);
nand U13800 (N_13800,N_10415,N_9897);
nand U13801 (N_13801,N_9608,N_11657);
nor U13802 (N_13802,N_9792,N_11698);
nand U13803 (N_13803,N_10635,N_12348);
or U13804 (N_13804,N_10719,N_9883);
nand U13805 (N_13805,N_11243,N_10405);
xnor U13806 (N_13806,N_9640,N_12184);
nand U13807 (N_13807,N_11472,N_10976);
xnor U13808 (N_13808,N_12400,N_9783);
and U13809 (N_13809,N_11186,N_10413);
nand U13810 (N_13810,N_11797,N_9769);
nor U13811 (N_13811,N_11933,N_11120);
nor U13812 (N_13812,N_9891,N_9429);
nor U13813 (N_13813,N_12155,N_11059);
nor U13814 (N_13814,N_9597,N_10725);
nand U13815 (N_13815,N_10803,N_10428);
and U13816 (N_13816,N_10337,N_11391);
or U13817 (N_13817,N_10935,N_10578);
nand U13818 (N_13818,N_9379,N_11908);
nor U13819 (N_13819,N_10016,N_9528);
nand U13820 (N_13820,N_9560,N_12334);
nand U13821 (N_13821,N_10330,N_11250);
nand U13822 (N_13822,N_11560,N_11951);
xor U13823 (N_13823,N_12272,N_11950);
nor U13824 (N_13824,N_12462,N_10892);
or U13825 (N_13825,N_12393,N_10112);
nor U13826 (N_13826,N_11735,N_11488);
nand U13827 (N_13827,N_9653,N_11009);
nand U13828 (N_13828,N_10069,N_10762);
or U13829 (N_13829,N_10507,N_10559);
nand U13830 (N_13830,N_9710,N_10600);
and U13831 (N_13831,N_12297,N_12146);
and U13832 (N_13832,N_12226,N_10234);
nand U13833 (N_13833,N_12425,N_11309);
nor U13834 (N_13834,N_10075,N_11032);
and U13835 (N_13835,N_10351,N_12378);
or U13836 (N_13836,N_9617,N_10232);
and U13837 (N_13837,N_12287,N_12280);
or U13838 (N_13838,N_10404,N_12339);
nor U13839 (N_13839,N_11964,N_10740);
nor U13840 (N_13840,N_9823,N_9599);
xnor U13841 (N_13841,N_10124,N_11724);
or U13842 (N_13842,N_12286,N_11526);
nor U13843 (N_13843,N_10076,N_10570);
nand U13844 (N_13844,N_10833,N_9708);
and U13845 (N_13845,N_11987,N_11261);
nor U13846 (N_13846,N_11606,N_12044);
xnor U13847 (N_13847,N_11417,N_11147);
or U13848 (N_13848,N_10198,N_10299);
or U13849 (N_13849,N_12412,N_9999);
or U13850 (N_13850,N_12459,N_11553);
xor U13851 (N_13851,N_11847,N_11347);
and U13852 (N_13852,N_11906,N_11625);
and U13853 (N_13853,N_12152,N_10066);
and U13854 (N_13854,N_12353,N_12251);
xor U13855 (N_13855,N_9446,N_11042);
and U13856 (N_13856,N_11363,N_12104);
xnor U13857 (N_13857,N_9819,N_10420);
nand U13858 (N_13858,N_9698,N_12323);
xnor U13859 (N_13859,N_12097,N_10645);
xor U13860 (N_13860,N_10975,N_11771);
nand U13861 (N_13861,N_12058,N_11182);
or U13862 (N_13862,N_11420,N_10451);
xnor U13863 (N_13863,N_10669,N_11879);
xnor U13864 (N_13864,N_10701,N_9718);
nor U13865 (N_13865,N_10147,N_11389);
xor U13866 (N_13866,N_11163,N_12363);
xnor U13867 (N_13867,N_12277,N_10710);
nand U13868 (N_13868,N_10438,N_11191);
xor U13869 (N_13869,N_10021,N_11422);
nand U13870 (N_13870,N_10682,N_9840);
and U13871 (N_13871,N_9935,N_9720);
nor U13872 (N_13872,N_10835,N_11039);
nand U13873 (N_13873,N_11432,N_9545);
nor U13874 (N_13874,N_11588,N_12094);
xor U13875 (N_13875,N_10284,N_9421);
or U13876 (N_13876,N_10315,N_12124);
or U13877 (N_13877,N_11019,N_11178);
xor U13878 (N_13878,N_11846,N_12342);
and U13879 (N_13879,N_12444,N_9578);
nand U13880 (N_13880,N_9993,N_10288);
or U13881 (N_13881,N_9579,N_9464);
and U13882 (N_13882,N_10987,N_11017);
xnor U13883 (N_13883,N_9687,N_10250);
nor U13884 (N_13884,N_10552,N_10778);
nand U13885 (N_13885,N_10545,N_10957);
and U13886 (N_13886,N_10091,N_11562);
nand U13887 (N_13887,N_9590,N_9835);
nor U13888 (N_13888,N_11999,N_9529);
and U13889 (N_13889,N_9721,N_10114);
nand U13890 (N_13890,N_12141,N_11088);
nand U13891 (N_13891,N_10820,N_11706);
nor U13892 (N_13892,N_10972,N_10947);
or U13893 (N_13893,N_10619,N_10981);
nor U13894 (N_13894,N_10430,N_9766);
nand U13895 (N_13895,N_11822,N_9605);
and U13896 (N_13896,N_9641,N_12187);
and U13897 (N_13897,N_11622,N_10999);
or U13898 (N_13898,N_9779,N_11982);
and U13899 (N_13899,N_11037,N_11728);
nor U13900 (N_13900,N_12177,N_9454);
and U13901 (N_13901,N_10272,N_9744);
nor U13902 (N_13902,N_11125,N_9927);
nor U13903 (N_13903,N_12270,N_12015);
xnor U13904 (N_13904,N_10704,N_9533);
and U13905 (N_13905,N_12312,N_11028);
nor U13906 (N_13906,N_10360,N_11721);
or U13907 (N_13907,N_10282,N_11589);
or U13908 (N_13908,N_12433,N_10558);
or U13909 (N_13909,N_10057,N_10445);
nor U13910 (N_13910,N_9519,N_10513);
or U13911 (N_13911,N_9554,N_12347);
nor U13912 (N_13912,N_11169,N_11520);
nor U13913 (N_13913,N_11176,N_10359);
nand U13914 (N_13914,N_10877,N_10613);
nor U13915 (N_13915,N_11394,N_12118);
and U13916 (N_13916,N_12337,N_10418);
and U13917 (N_13917,N_10017,N_11362);
nand U13918 (N_13918,N_10169,N_10714);
and U13919 (N_13919,N_9392,N_11617);
nor U13920 (N_13920,N_12261,N_12255);
xor U13921 (N_13921,N_10478,N_11448);
xnor U13922 (N_13922,N_12191,N_10136);
nand U13923 (N_13923,N_10237,N_9801);
xor U13924 (N_13924,N_11115,N_11299);
xor U13925 (N_13925,N_10751,N_10651);
nor U13926 (N_13926,N_9896,N_11463);
nor U13927 (N_13927,N_11857,N_9782);
and U13928 (N_13928,N_11090,N_9390);
nor U13929 (N_13929,N_11480,N_12487);
and U13930 (N_13930,N_12245,N_10916);
xnor U13931 (N_13931,N_10639,N_10509);
or U13932 (N_13932,N_11334,N_11302);
nor U13933 (N_13933,N_11126,N_10876);
nor U13934 (N_13934,N_12241,N_12483);
nand U13935 (N_13935,N_11935,N_10472);
and U13936 (N_13936,N_11300,N_10791);
xor U13937 (N_13937,N_11676,N_10691);
and U13938 (N_13938,N_10457,N_10792);
nand U13939 (N_13939,N_12219,N_11425);
nand U13940 (N_13940,N_9944,N_9649);
and U13941 (N_13941,N_11759,N_11353);
or U13942 (N_13942,N_11539,N_10814);
nand U13943 (N_13943,N_11307,N_12447);
nor U13944 (N_13944,N_11251,N_11414);
and U13945 (N_13945,N_9481,N_12372);
nor U13946 (N_13946,N_11516,N_10650);
nand U13947 (N_13947,N_10257,N_12087);
nand U13948 (N_13948,N_10572,N_9508);
xor U13949 (N_13949,N_11400,N_11218);
or U13950 (N_13950,N_12170,N_10621);
nand U13951 (N_13951,N_11503,N_12216);
nor U13952 (N_13952,N_11942,N_9477);
xnor U13953 (N_13953,N_11466,N_10615);
nor U13954 (N_13954,N_11675,N_11522);
nor U13955 (N_13955,N_10258,N_10533);
and U13956 (N_13956,N_10647,N_10362);
nor U13957 (N_13957,N_12235,N_11199);
xnor U13958 (N_13958,N_11909,N_12293);
or U13959 (N_13959,N_11723,N_9488);
and U13960 (N_13960,N_10370,N_9696);
and U13961 (N_13961,N_12031,N_12021);
nor U13962 (N_13962,N_9821,N_11223);
xnor U13963 (N_13963,N_12041,N_11046);
xnor U13964 (N_13964,N_12449,N_11888);
and U13965 (N_13965,N_9774,N_9702);
nand U13966 (N_13966,N_11451,N_11103);
xnor U13967 (N_13967,N_9652,N_11980);
nor U13968 (N_13968,N_9642,N_11881);
or U13969 (N_13969,N_9505,N_12134);
nand U13970 (N_13970,N_9888,N_11006);
nor U13971 (N_13971,N_9913,N_11238);
or U13972 (N_13972,N_10476,N_11958);
nor U13973 (N_13973,N_12105,N_11621);
and U13974 (N_13974,N_12045,N_9892);
and U13975 (N_13975,N_10674,N_12333);
nor U13976 (N_13976,N_11786,N_12269);
or U13977 (N_13977,N_11327,N_10079);
or U13978 (N_13978,N_10334,N_10945);
and U13979 (N_13979,N_10919,N_11478);
nor U13980 (N_13980,N_9457,N_10332);
or U13981 (N_13981,N_11047,N_10247);
and U13982 (N_13982,N_11911,N_11623);
xor U13983 (N_13983,N_11172,N_10592);
nor U13984 (N_13984,N_10933,N_12075);
xor U13985 (N_13985,N_10538,N_11801);
xnor U13986 (N_13986,N_12310,N_10629);
nor U13987 (N_13987,N_10444,N_12492);
and U13988 (N_13988,N_11583,N_10313);
nor U13989 (N_13989,N_10144,N_10692);
nand U13990 (N_13990,N_9565,N_9849);
xor U13991 (N_13991,N_9404,N_11294);
xnor U13992 (N_13992,N_11152,N_11279);
nor U13993 (N_13993,N_12175,N_11333);
nand U13994 (N_13994,N_10808,N_10101);
nor U13995 (N_13995,N_12231,N_12057);
or U13996 (N_13996,N_9489,N_11684);
or U13997 (N_13997,N_10271,N_11224);
and U13998 (N_13998,N_9510,N_10461);
nor U13999 (N_13999,N_10450,N_11708);
xnor U14000 (N_14000,N_10586,N_10278);
xor U14001 (N_14001,N_11415,N_11470);
nor U14002 (N_14002,N_9694,N_10156);
and U14003 (N_14003,N_9929,N_9970);
nor U14004 (N_14004,N_10894,N_9681);
xor U14005 (N_14005,N_10488,N_11671);
and U14006 (N_14006,N_12024,N_10001);
or U14007 (N_14007,N_10133,N_10134);
and U14008 (N_14008,N_9836,N_11687);
nor U14009 (N_14009,N_11192,N_12092);
xnor U14010 (N_14010,N_11756,N_9688);
nand U14011 (N_14011,N_10052,N_11753);
or U14012 (N_14012,N_10758,N_9791);
xor U14013 (N_14013,N_9872,N_12456);
nand U14014 (N_14014,N_10922,N_10846);
and U14015 (N_14015,N_12252,N_11094);
and U14016 (N_14016,N_11235,N_11407);
nor U14017 (N_14017,N_12361,N_10265);
xnor U14018 (N_14018,N_9962,N_10713);
and U14019 (N_14019,N_12289,N_12479);
nand U14020 (N_14020,N_10505,N_9908);
or U14021 (N_14021,N_9397,N_11495);
and U14022 (N_14022,N_9498,N_11174);
nor U14023 (N_14023,N_11493,N_11366);
or U14024 (N_14024,N_9746,N_11871);
nand U14025 (N_14025,N_11805,N_9771);
or U14026 (N_14026,N_9383,N_9950);
xnor U14027 (N_14027,N_10768,N_10949);
or U14028 (N_14028,N_11680,N_10190);
xnor U14029 (N_14029,N_10853,N_10200);
and U14030 (N_14030,N_10963,N_11608);
nand U14031 (N_14031,N_9880,N_10886);
xor U14032 (N_14032,N_10437,N_9469);
nor U14033 (N_14033,N_9847,N_12467);
or U14034 (N_14034,N_9912,N_9471);
and U14035 (N_14035,N_11854,N_11441);
and U14036 (N_14036,N_10767,N_10789);
or U14037 (N_14037,N_10699,N_10398);
xor U14038 (N_14038,N_10867,N_12115);
nand U14039 (N_14039,N_11436,N_10216);
nor U14040 (N_14040,N_10396,N_9920);
nand U14041 (N_14041,N_10643,N_11765);
and U14042 (N_14042,N_11185,N_10155);
and U14043 (N_14043,N_9707,N_9532);
and U14044 (N_14044,N_10055,N_12035);
xor U14045 (N_14045,N_12375,N_11604);
nand U14046 (N_14046,N_11694,N_12328);
or U14047 (N_14047,N_10392,N_11345);
nor U14048 (N_14048,N_11767,N_11567);
nor U14049 (N_14049,N_11695,N_10291);
or U14050 (N_14050,N_11162,N_10715);
nor U14051 (N_14051,N_11464,N_10734);
and U14052 (N_14052,N_10936,N_10504);
nor U14053 (N_14053,N_10722,N_10903);
xnor U14054 (N_14054,N_11901,N_10811);
or U14055 (N_14055,N_11974,N_11343);
nor U14056 (N_14056,N_9785,N_12385);
nand U14057 (N_14057,N_10098,N_11792);
nor U14058 (N_14058,N_11566,N_10960);
nand U14059 (N_14059,N_11093,N_12018);
nor U14060 (N_14060,N_11230,N_11620);
nand U14061 (N_14061,N_12110,N_9538);
nand U14062 (N_14062,N_10805,N_12374);
or U14063 (N_14063,N_9702,N_11748);
and U14064 (N_14064,N_12357,N_11661);
or U14065 (N_14065,N_9437,N_11906);
nand U14066 (N_14066,N_12103,N_11663);
nand U14067 (N_14067,N_10754,N_11435);
and U14068 (N_14068,N_10975,N_10599);
or U14069 (N_14069,N_10210,N_11589);
nor U14070 (N_14070,N_12088,N_9689);
and U14071 (N_14071,N_12442,N_10336);
or U14072 (N_14072,N_11791,N_12433);
xnor U14073 (N_14073,N_10163,N_9519);
and U14074 (N_14074,N_10787,N_11269);
nor U14075 (N_14075,N_11768,N_11780);
nand U14076 (N_14076,N_11737,N_12061);
and U14077 (N_14077,N_9662,N_11868);
and U14078 (N_14078,N_10523,N_11456);
and U14079 (N_14079,N_10088,N_10093);
and U14080 (N_14080,N_9755,N_11902);
and U14081 (N_14081,N_9508,N_10310);
or U14082 (N_14082,N_11252,N_9411);
nand U14083 (N_14083,N_11281,N_12397);
xor U14084 (N_14084,N_10406,N_12439);
nand U14085 (N_14085,N_10569,N_10227);
xnor U14086 (N_14086,N_10463,N_12035);
xnor U14087 (N_14087,N_12106,N_10311);
and U14088 (N_14088,N_11832,N_12380);
xor U14089 (N_14089,N_11239,N_10826);
and U14090 (N_14090,N_10727,N_12125);
and U14091 (N_14091,N_11632,N_10904);
or U14092 (N_14092,N_10132,N_12209);
and U14093 (N_14093,N_9737,N_9906);
or U14094 (N_14094,N_10610,N_11512);
and U14095 (N_14095,N_11501,N_10983);
nor U14096 (N_14096,N_10267,N_9853);
nor U14097 (N_14097,N_11591,N_9456);
or U14098 (N_14098,N_10032,N_9689);
nand U14099 (N_14099,N_11838,N_11256);
nor U14100 (N_14100,N_12323,N_9635);
or U14101 (N_14101,N_9873,N_12428);
nand U14102 (N_14102,N_9848,N_10185);
or U14103 (N_14103,N_12271,N_10088);
nor U14104 (N_14104,N_10989,N_9739);
nand U14105 (N_14105,N_12260,N_12073);
xnor U14106 (N_14106,N_10797,N_12191);
and U14107 (N_14107,N_11909,N_11694);
and U14108 (N_14108,N_10508,N_10697);
or U14109 (N_14109,N_12368,N_9509);
nor U14110 (N_14110,N_9436,N_10521);
nand U14111 (N_14111,N_10364,N_11918);
nor U14112 (N_14112,N_12128,N_11140);
nor U14113 (N_14113,N_11619,N_12357);
or U14114 (N_14114,N_12273,N_11068);
nor U14115 (N_14115,N_10798,N_11698);
and U14116 (N_14116,N_11843,N_10897);
xnor U14117 (N_14117,N_11464,N_11115);
nand U14118 (N_14118,N_9498,N_11770);
xor U14119 (N_14119,N_10492,N_12154);
xor U14120 (N_14120,N_11997,N_12227);
xnor U14121 (N_14121,N_10500,N_10141);
or U14122 (N_14122,N_11123,N_10762);
or U14123 (N_14123,N_9605,N_10230);
xnor U14124 (N_14124,N_9843,N_10485);
nand U14125 (N_14125,N_10488,N_10392);
and U14126 (N_14126,N_10670,N_10098);
and U14127 (N_14127,N_11305,N_10705);
and U14128 (N_14128,N_11023,N_10732);
nor U14129 (N_14129,N_10963,N_9579);
xnor U14130 (N_14130,N_10692,N_9957);
nor U14131 (N_14131,N_9999,N_12372);
or U14132 (N_14132,N_9896,N_11625);
nor U14133 (N_14133,N_9999,N_9932);
xnor U14134 (N_14134,N_9814,N_11895);
nand U14135 (N_14135,N_10207,N_11151);
nor U14136 (N_14136,N_12062,N_9462);
xor U14137 (N_14137,N_11112,N_12421);
xnor U14138 (N_14138,N_11709,N_10241);
nor U14139 (N_14139,N_10191,N_10637);
xnor U14140 (N_14140,N_9414,N_11339);
and U14141 (N_14141,N_12427,N_10561);
nand U14142 (N_14142,N_12175,N_11147);
xnor U14143 (N_14143,N_12266,N_9533);
and U14144 (N_14144,N_11161,N_9764);
xnor U14145 (N_14145,N_10633,N_12178);
nor U14146 (N_14146,N_10080,N_10459);
and U14147 (N_14147,N_9890,N_11946);
and U14148 (N_14148,N_10155,N_9517);
and U14149 (N_14149,N_10722,N_11411);
and U14150 (N_14150,N_11908,N_11607);
nand U14151 (N_14151,N_11841,N_12283);
nand U14152 (N_14152,N_9773,N_11041);
nor U14153 (N_14153,N_9823,N_10056);
or U14154 (N_14154,N_10103,N_11602);
nor U14155 (N_14155,N_10814,N_11815);
or U14156 (N_14156,N_10930,N_10157);
or U14157 (N_14157,N_11825,N_12051);
and U14158 (N_14158,N_10016,N_9968);
and U14159 (N_14159,N_12247,N_10816);
and U14160 (N_14160,N_10473,N_10394);
or U14161 (N_14161,N_11090,N_10422);
or U14162 (N_14162,N_11628,N_10115);
nand U14163 (N_14163,N_12381,N_12139);
xor U14164 (N_14164,N_9696,N_11388);
and U14165 (N_14165,N_9434,N_12471);
and U14166 (N_14166,N_11657,N_11006);
nand U14167 (N_14167,N_10828,N_11607);
xnor U14168 (N_14168,N_9879,N_9784);
or U14169 (N_14169,N_10460,N_9804);
or U14170 (N_14170,N_9391,N_12341);
and U14171 (N_14171,N_11557,N_11926);
or U14172 (N_14172,N_11596,N_11496);
nand U14173 (N_14173,N_12267,N_10832);
xor U14174 (N_14174,N_10078,N_10134);
and U14175 (N_14175,N_11196,N_11319);
or U14176 (N_14176,N_11255,N_11776);
and U14177 (N_14177,N_10624,N_11048);
xor U14178 (N_14178,N_11076,N_9924);
and U14179 (N_14179,N_11153,N_12337);
nor U14180 (N_14180,N_10702,N_11904);
xor U14181 (N_14181,N_10664,N_12489);
or U14182 (N_14182,N_12216,N_10188);
nor U14183 (N_14183,N_10779,N_10605);
nor U14184 (N_14184,N_11632,N_9715);
and U14185 (N_14185,N_9635,N_9822);
nand U14186 (N_14186,N_10820,N_11297);
or U14187 (N_14187,N_9492,N_10152);
nand U14188 (N_14188,N_10410,N_10070);
or U14189 (N_14189,N_9488,N_9854);
or U14190 (N_14190,N_10475,N_10314);
xnor U14191 (N_14191,N_10111,N_11510);
nand U14192 (N_14192,N_10182,N_11075);
nand U14193 (N_14193,N_11530,N_11677);
xnor U14194 (N_14194,N_11113,N_10748);
or U14195 (N_14195,N_9713,N_10526);
xor U14196 (N_14196,N_10853,N_11808);
nor U14197 (N_14197,N_11957,N_11501);
or U14198 (N_14198,N_11533,N_10420);
and U14199 (N_14199,N_12312,N_10458);
nand U14200 (N_14200,N_9730,N_10664);
nand U14201 (N_14201,N_11396,N_11452);
or U14202 (N_14202,N_10968,N_12071);
or U14203 (N_14203,N_11615,N_9871);
xnor U14204 (N_14204,N_11748,N_11552);
or U14205 (N_14205,N_11719,N_11452);
or U14206 (N_14206,N_10700,N_10863);
nand U14207 (N_14207,N_11369,N_9772);
nand U14208 (N_14208,N_10906,N_12375);
nor U14209 (N_14209,N_10543,N_9718);
nand U14210 (N_14210,N_11970,N_10858);
and U14211 (N_14211,N_11890,N_10267);
nand U14212 (N_14212,N_11498,N_11996);
nand U14213 (N_14213,N_11654,N_12105);
xnor U14214 (N_14214,N_11923,N_11743);
xor U14215 (N_14215,N_11827,N_11736);
nand U14216 (N_14216,N_11348,N_12467);
or U14217 (N_14217,N_10404,N_10169);
nor U14218 (N_14218,N_9562,N_11285);
xnor U14219 (N_14219,N_10523,N_9839);
nand U14220 (N_14220,N_10824,N_11619);
or U14221 (N_14221,N_11152,N_11938);
or U14222 (N_14222,N_11820,N_9989);
nor U14223 (N_14223,N_9880,N_11059);
or U14224 (N_14224,N_10416,N_11893);
and U14225 (N_14225,N_11449,N_11319);
xnor U14226 (N_14226,N_10596,N_10095);
or U14227 (N_14227,N_10717,N_12429);
xnor U14228 (N_14228,N_11576,N_11480);
or U14229 (N_14229,N_9701,N_9759);
xor U14230 (N_14230,N_10611,N_12052);
xor U14231 (N_14231,N_12299,N_10456);
nor U14232 (N_14232,N_10672,N_12173);
nor U14233 (N_14233,N_10068,N_10315);
xor U14234 (N_14234,N_9803,N_10665);
or U14235 (N_14235,N_12231,N_11494);
nand U14236 (N_14236,N_12416,N_9428);
and U14237 (N_14237,N_12337,N_11259);
and U14238 (N_14238,N_9424,N_9459);
and U14239 (N_14239,N_10307,N_9947);
nand U14240 (N_14240,N_9975,N_9817);
nor U14241 (N_14241,N_9946,N_11856);
nor U14242 (N_14242,N_11018,N_12050);
nand U14243 (N_14243,N_9796,N_9537);
nand U14244 (N_14244,N_10865,N_9929);
or U14245 (N_14245,N_11745,N_9470);
and U14246 (N_14246,N_10582,N_10849);
xor U14247 (N_14247,N_9624,N_11722);
and U14248 (N_14248,N_9997,N_11623);
and U14249 (N_14249,N_11350,N_12456);
nand U14250 (N_14250,N_11627,N_10119);
and U14251 (N_14251,N_9706,N_10261);
xnor U14252 (N_14252,N_10510,N_11122);
and U14253 (N_14253,N_10029,N_9767);
nor U14254 (N_14254,N_12494,N_10555);
xnor U14255 (N_14255,N_9714,N_10868);
or U14256 (N_14256,N_11159,N_9851);
nand U14257 (N_14257,N_12154,N_10429);
or U14258 (N_14258,N_10722,N_9710);
xor U14259 (N_14259,N_11026,N_11557);
and U14260 (N_14260,N_11727,N_11183);
and U14261 (N_14261,N_11446,N_11221);
nand U14262 (N_14262,N_9918,N_11467);
nand U14263 (N_14263,N_9683,N_11404);
xnor U14264 (N_14264,N_11297,N_11581);
and U14265 (N_14265,N_12004,N_11596);
or U14266 (N_14266,N_10799,N_11010);
xor U14267 (N_14267,N_9881,N_11796);
nor U14268 (N_14268,N_12026,N_10030);
and U14269 (N_14269,N_10757,N_10364);
nand U14270 (N_14270,N_11015,N_11941);
xor U14271 (N_14271,N_12233,N_10582);
nand U14272 (N_14272,N_10623,N_10940);
xnor U14273 (N_14273,N_10597,N_11973);
and U14274 (N_14274,N_12488,N_10845);
xnor U14275 (N_14275,N_12140,N_9806);
nand U14276 (N_14276,N_9407,N_11802);
or U14277 (N_14277,N_11085,N_11148);
xor U14278 (N_14278,N_11143,N_10696);
or U14279 (N_14279,N_9899,N_10180);
xnor U14280 (N_14280,N_11924,N_11820);
xnor U14281 (N_14281,N_11238,N_12437);
and U14282 (N_14282,N_11241,N_11010);
nor U14283 (N_14283,N_11218,N_11158);
xnor U14284 (N_14284,N_11069,N_9677);
or U14285 (N_14285,N_11920,N_10871);
and U14286 (N_14286,N_11003,N_9747);
nand U14287 (N_14287,N_10687,N_11529);
xor U14288 (N_14288,N_9560,N_11594);
xor U14289 (N_14289,N_9610,N_10262);
and U14290 (N_14290,N_11487,N_11381);
nand U14291 (N_14291,N_12455,N_12250);
nor U14292 (N_14292,N_11158,N_11486);
nor U14293 (N_14293,N_9743,N_11298);
xnor U14294 (N_14294,N_11281,N_10984);
and U14295 (N_14295,N_11367,N_10152);
nor U14296 (N_14296,N_11551,N_10070);
xor U14297 (N_14297,N_10399,N_12499);
xnor U14298 (N_14298,N_9464,N_10215);
nand U14299 (N_14299,N_10103,N_12109);
xnor U14300 (N_14300,N_12175,N_11088);
nor U14301 (N_14301,N_9547,N_12309);
nor U14302 (N_14302,N_11982,N_9676);
nor U14303 (N_14303,N_10136,N_9990);
or U14304 (N_14304,N_11114,N_12210);
or U14305 (N_14305,N_9494,N_9647);
and U14306 (N_14306,N_11292,N_9801);
nand U14307 (N_14307,N_9550,N_10000);
nand U14308 (N_14308,N_9924,N_11916);
or U14309 (N_14309,N_11391,N_11784);
nor U14310 (N_14310,N_10357,N_12023);
nor U14311 (N_14311,N_10062,N_9483);
xor U14312 (N_14312,N_10113,N_12320);
or U14313 (N_14313,N_11584,N_11446);
nor U14314 (N_14314,N_12274,N_11032);
and U14315 (N_14315,N_10067,N_9869);
xor U14316 (N_14316,N_12124,N_10625);
or U14317 (N_14317,N_10823,N_12230);
and U14318 (N_14318,N_11815,N_10410);
nand U14319 (N_14319,N_10863,N_10576);
nand U14320 (N_14320,N_11642,N_11832);
and U14321 (N_14321,N_9413,N_10328);
xor U14322 (N_14322,N_11041,N_11805);
xor U14323 (N_14323,N_9763,N_10411);
nand U14324 (N_14324,N_10713,N_12218);
nor U14325 (N_14325,N_9754,N_11463);
xor U14326 (N_14326,N_12192,N_12008);
or U14327 (N_14327,N_9616,N_10780);
nand U14328 (N_14328,N_10135,N_11265);
or U14329 (N_14329,N_9817,N_11264);
nand U14330 (N_14330,N_11224,N_10560);
and U14331 (N_14331,N_10425,N_10055);
nor U14332 (N_14332,N_11070,N_10820);
or U14333 (N_14333,N_12207,N_11919);
nor U14334 (N_14334,N_10312,N_9970);
nand U14335 (N_14335,N_11315,N_11686);
nand U14336 (N_14336,N_10280,N_10246);
xor U14337 (N_14337,N_11606,N_11683);
nor U14338 (N_14338,N_11527,N_12132);
and U14339 (N_14339,N_9600,N_10139);
xnor U14340 (N_14340,N_10728,N_10933);
nand U14341 (N_14341,N_12191,N_9389);
and U14342 (N_14342,N_10028,N_12134);
nor U14343 (N_14343,N_10821,N_10977);
xnor U14344 (N_14344,N_9760,N_10812);
nor U14345 (N_14345,N_10180,N_11092);
and U14346 (N_14346,N_12369,N_9926);
nor U14347 (N_14347,N_10221,N_10578);
xor U14348 (N_14348,N_10093,N_11159);
or U14349 (N_14349,N_12176,N_9841);
nor U14350 (N_14350,N_10805,N_10532);
xor U14351 (N_14351,N_9755,N_11016);
xnor U14352 (N_14352,N_11078,N_11803);
xnor U14353 (N_14353,N_11047,N_9589);
nor U14354 (N_14354,N_10850,N_9941);
and U14355 (N_14355,N_11014,N_11793);
xor U14356 (N_14356,N_11692,N_12002);
xnor U14357 (N_14357,N_11396,N_10259);
and U14358 (N_14358,N_12447,N_12384);
nor U14359 (N_14359,N_12091,N_11566);
or U14360 (N_14360,N_11905,N_10023);
nor U14361 (N_14361,N_9913,N_10799);
xor U14362 (N_14362,N_10750,N_10682);
nand U14363 (N_14363,N_11939,N_11956);
or U14364 (N_14364,N_12184,N_11210);
nor U14365 (N_14365,N_10613,N_9863);
xnor U14366 (N_14366,N_10986,N_11611);
xnor U14367 (N_14367,N_10234,N_11502);
xor U14368 (N_14368,N_9471,N_10850);
or U14369 (N_14369,N_11855,N_11896);
nand U14370 (N_14370,N_12316,N_11144);
xnor U14371 (N_14371,N_9983,N_10937);
nor U14372 (N_14372,N_11659,N_9782);
nor U14373 (N_14373,N_10686,N_9751);
xnor U14374 (N_14374,N_12340,N_11746);
or U14375 (N_14375,N_11600,N_11378);
or U14376 (N_14376,N_9449,N_10408);
and U14377 (N_14377,N_10425,N_11416);
or U14378 (N_14378,N_10001,N_9758);
xnor U14379 (N_14379,N_10730,N_11607);
nor U14380 (N_14380,N_11948,N_9522);
nand U14381 (N_14381,N_10976,N_9445);
or U14382 (N_14382,N_9732,N_12231);
and U14383 (N_14383,N_11306,N_10961);
nor U14384 (N_14384,N_9866,N_9725);
xnor U14385 (N_14385,N_12102,N_10782);
and U14386 (N_14386,N_12219,N_9545);
nand U14387 (N_14387,N_12340,N_11093);
xor U14388 (N_14388,N_11084,N_11417);
nor U14389 (N_14389,N_10105,N_11645);
or U14390 (N_14390,N_9513,N_9797);
xnor U14391 (N_14391,N_10179,N_10877);
or U14392 (N_14392,N_10081,N_11789);
xor U14393 (N_14393,N_11561,N_12201);
and U14394 (N_14394,N_10651,N_10970);
or U14395 (N_14395,N_11248,N_11490);
and U14396 (N_14396,N_9457,N_11865);
nor U14397 (N_14397,N_9472,N_9754);
nand U14398 (N_14398,N_12390,N_11185);
nor U14399 (N_14399,N_10824,N_10119);
or U14400 (N_14400,N_9398,N_10168);
and U14401 (N_14401,N_9434,N_9396);
nand U14402 (N_14402,N_11503,N_11025);
and U14403 (N_14403,N_9659,N_11298);
nor U14404 (N_14404,N_9608,N_9430);
or U14405 (N_14405,N_11332,N_10405);
and U14406 (N_14406,N_10252,N_10443);
and U14407 (N_14407,N_9585,N_11845);
nand U14408 (N_14408,N_11724,N_10657);
xnor U14409 (N_14409,N_11474,N_10449);
nand U14410 (N_14410,N_10866,N_9496);
and U14411 (N_14411,N_11207,N_12343);
xor U14412 (N_14412,N_9661,N_12032);
and U14413 (N_14413,N_11085,N_10828);
xor U14414 (N_14414,N_10551,N_10963);
nand U14415 (N_14415,N_10666,N_11070);
or U14416 (N_14416,N_11347,N_10432);
and U14417 (N_14417,N_11463,N_11264);
and U14418 (N_14418,N_10896,N_10155);
or U14419 (N_14419,N_10358,N_11530);
nor U14420 (N_14420,N_11963,N_9668);
xnor U14421 (N_14421,N_11667,N_10249);
and U14422 (N_14422,N_11653,N_11699);
nand U14423 (N_14423,N_12325,N_11660);
nand U14424 (N_14424,N_11619,N_12478);
and U14425 (N_14425,N_10277,N_11858);
or U14426 (N_14426,N_11451,N_9794);
nor U14427 (N_14427,N_11168,N_11639);
or U14428 (N_14428,N_10123,N_9894);
nand U14429 (N_14429,N_12210,N_11807);
nor U14430 (N_14430,N_11982,N_11421);
xor U14431 (N_14431,N_10282,N_11534);
xnor U14432 (N_14432,N_11868,N_11153);
xor U14433 (N_14433,N_12108,N_11564);
and U14434 (N_14434,N_11000,N_10051);
nor U14435 (N_14435,N_10694,N_11718);
xor U14436 (N_14436,N_12024,N_10941);
nand U14437 (N_14437,N_12073,N_9820);
nor U14438 (N_14438,N_10641,N_11682);
nor U14439 (N_14439,N_11253,N_9720);
or U14440 (N_14440,N_10083,N_9628);
and U14441 (N_14441,N_11072,N_11558);
nor U14442 (N_14442,N_9587,N_9865);
nand U14443 (N_14443,N_9555,N_11139);
and U14444 (N_14444,N_11164,N_9744);
or U14445 (N_14445,N_11798,N_12041);
nor U14446 (N_14446,N_11771,N_9970);
and U14447 (N_14447,N_11107,N_9408);
xnor U14448 (N_14448,N_12370,N_11328);
nand U14449 (N_14449,N_11245,N_11161);
nand U14450 (N_14450,N_11490,N_10064);
nand U14451 (N_14451,N_11764,N_11401);
nand U14452 (N_14452,N_12324,N_9446);
nor U14453 (N_14453,N_12349,N_10925);
or U14454 (N_14454,N_12320,N_9702);
or U14455 (N_14455,N_11586,N_10226);
and U14456 (N_14456,N_10976,N_11723);
nor U14457 (N_14457,N_12290,N_10997);
nor U14458 (N_14458,N_11984,N_11987);
nor U14459 (N_14459,N_9911,N_9446);
and U14460 (N_14460,N_10756,N_12013);
nand U14461 (N_14461,N_10197,N_11086);
xor U14462 (N_14462,N_9491,N_11852);
xnor U14463 (N_14463,N_10514,N_11672);
xor U14464 (N_14464,N_11149,N_11638);
nor U14465 (N_14465,N_12368,N_11646);
nor U14466 (N_14466,N_10870,N_10707);
nor U14467 (N_14467,N_9823,N_10131);
xnor U14468 (N_14468,N_9909,N_9618);
nor U14469 (N_14469,N_11254,N_10898);
nand U14470 (N_14470,N_9833,N_10159);
and U14471 (N_14471,N_9812,N_12122);
nand U14472 (N_14472,N_11959,N_9944);
nor U14473 (N_14473,N_9827,N_10668);
nor U14474 (N_14474,N_10091,N_11998);
nand U14475 (N_14475,N_11473,N_12177);
nor U14476 (N_14476,N_11529,N_11265);
and U14477 (N_14477,N_12488,N_12003);
xor U14478 (N_14478,N_10353,N_10388);
nand U14479 (N_14479,N_10920,N_10318);
nand U14480 (N_14480,N_11150,N_10577);
nand U14481 (N_14481,N_11975,N_9969);
xor U14482 (N_14482,N_9408,N_12289);
or U14483 (N_14483,N_11251,N_9511);
or U14484 (N_14484,N_11197,N_12210);
or U14485 (N_14485,N_10872,N_10013);
nand U14486 (N_14486,N_10694,N_11972);
and U14487 (N_14487,N_10645,N_11706);
nor U14488 (N_14488,N_9824,N_10529);
xnor U14489 (N_14489,N_11598,N_12035);
or U14490 (N_14490,N_10276,N_10546);
or U14491 (N_14491,N_11291,N_12446);
and U14492 (N_14492,N_12206,N_11798);
nand U14493 (N_14493,N_10451,N_10675);
or U14494 (N_14494,N_10443,N_12015);
nand U14495 (N_14495,N_10339,N_11621);
nand U14496 (N_14496,N_10523,N_9781);
nand U14497 (N_14497,N_9441,N_9757);
nand U14498 (N_14498,N_10891,N_12378);
xor U14499 (N_14499,N_12312,N_9556);
nor U14500 (N_14500,N_10146,N_10361);
nor U14501 (N_14501,N_10519,N_10679);
or U14502 (N_14502,N_12076,N_12421);
xnor U14503 (N_14503,N_11468,N_9582);
and U14504 (N_14504,N_11278,N_10563);
xor U14505 (N_14505,N_11057,N_12316);
or U14506 (N_14506,N_10326,N_12021);
xor U14507 (N_14507,N_11301,N_9709);
nor U14508 (N_14508,N_12220,N_11974);
nand U14509 (N_14509,N_12363,N_10840);
nor U14510 (N_14510,N_10144,N_9379);
xor U14511 (N_14511,N_11039,N_12249);
or U14512 (N_14512,N_12186,N_11309);
and U14513 (N_14513,N_11671,N_11669);
and U14514 (N_14514,N_10946,N_10914);
and U14515 (N_14515,N_10313,N_9726);
nor U14516 (N_14516,N_10848,N_11044);
xnor U14517 (N_14517,N_9456,N_10504);
or U14518 (N_14518,N_11999,N_11323);
and U14519 (N_14519,N_11074,N_9605);
xor U14520 (N_14520,N_11127,N_9702);
nor U14521 (N_14521,N_11615,N_10312);
and U14522 (N_14522,N_10434,N_12435);
or U14523 (N_14523,N_10702,N_10539);
xnor U14524 (N_14524,N_11047,N_11993);
and U14525 (N_14525,N_12387,N_11169);
or U14526 (N_14526,N_11675,N_9405);
and U14527 (N_14527,N_11146,N_10426);
nand U14528 (N_14528,N_10853,N_9500);
and U14529 (N_14529,N_10587,N_10802);
and U14530 (N_14530,N_11115,N_9913);
and U14531 (N_14531,N_10981,N_10611);
and U14532 (N_14532,N_10356,N_10403);
or U14533 (N_14533,N_9454,N_9394);
nor U14534 (N_14534,N_11040,N_11638);
nor U14535 (N_14535,N_10627,N_11679);
nand U14536 (N_14536,N_11032,N_11435);
or U14537 (N_14537,N_9946,N_11499);
or U14538 (N_14538,N_11182,N_10731);
and U14539 (N_14539,N_10493,N_9905);
and U14540 (N_14540,N_9688,N_12068);
or U14541 (N_14541,N_10863,N_11095);
or U14542 (N_14542,N_11568,N_10009);
xor U14543 (N_14543,N_10992,N_11341);
xnor U14544 (N_14544,N_9446,N_12116);
and U14545 (N_14545,N_10179,N_11787);
and U14546 (N_14546,N_10950,N_11875);
or U14547 (N_14547,N_10496,N_11946);
or U14548 (N_14548,N_12267,N_9533);
xnor U14549 (N_14549,N_11443,N_9927);
xor U14550 (N_14550,N_11606,N_9404);
nand U14551 (N_14551,N_10551,N_11435);
nand U14552 (N_14552,N_12054,N_11313);
and U14553 (N_14553,N_11737,N_12092);
and U14554 (N_14554,N_10578,N_9400);
xnor U14555 (N_14555,N_10285,N_11235);
or U14556 (N_14556,N_11598,N_9948);
nand U14557 (N_14557,N_11289,N_10528);
nand U14558 (N_14558,N_11381,N_11083);
nand U14559 (N_14559,N_12041,N_10245);
nand U14560 (N_14560,N_11669,N_11409);
nor U14561 (N_14561,N_11048,N_9610);
nand U14562 (N_14562,N_10899,N_9793);
nor U14563 (N_14563,N_12274,N_12327);
and U14564 (N_14564,N_11092,N_11227);
and U14565 (N_14565,N_10307,N_10845);
or U14566 (N_14566,N_10704,N_11348);
nor U14567 (N_14567,N_12244,N_11563);
nor U14568 (N_14568,N_10644,N_10090);
xnor U14569 (N_14569,N_9891,N_11009);
or U14570 (N_14570,N_12075,N_10643);
nand U14571 (N_14571,N_12179,N_10319);
and U14572 (N_14572,N_11142,N_12035);
nand U14573 (N_14573,N_9712,N_9843);
nor U14574 (N_14574,N_12442,N_10614);
nand U14575 (N_14575,N_9707,N_11171);
nor U14576 (N_14576,N_10236,N_9867);
nand U14577 (N_14577,N_12081,N_10027);
xor U14578 (N_14578,N_9576,N_9408);
nand U14579 (N_14579,N_11992,N_10470);
nor U14580 (N_14580,N_11820,N_12307);
xnor U14581 (N_14581,N_11802,N_12221);
nor U14582 (N_14582,N_11826,N_11545);
nand U14583 (N_14583,N_9625,N_10444);
nand U14584 (N_14584,N_9627,N_10781);
nand U14585 (N_14585,N_9391,N_11214);
or U14586 (N_14586,N_10567,N_9681);
and U14587 (N_14587,N_10870,N_11709);
nand U14588 (N_14588,N_10070,N_11736);
xnor U14589 (N_14589,N_10527,N_12047);
nand U14590 (N_14590,N_12157,N_11313);
nand U14591 (N_14591,N_12488,N_10268);
and U14592 (N_14592,N_11405,N_9469);
nor U14593 (N_14593,N_9995,N_10623);
nand U14594 (N_14594,N_10529,N_11506);
nor U14595 (N_14595,N_11389,N_11596);
and U14596 (N_14596,N_10942,N_11318);
and U14597 (N_14597,N_10958,N_10293);
nor U14598 (N_14598,N_10010,N_11944);
nand U14599 (N_14599,N_9404,N_10108);
nand U14600 (N_14600,N_10067,N_11311);
nor U14601 (N_14601,N_9686,N_11915);
or U14602 (N_14602,N_10633,N_12078);
xor U14603 (N_14603,N_10013,N_11288);
nand U14604 (N_14604,N_12324,N_10893);
nor U14605 (N_14605,N_12329,N_10258);
or U14606 (N_14606,N_10667,N_11952);
xor U14607 (N_14607,N_9749,N_9699);
xor U14608 (N_14608,N_12375,N_10563);
nor U14609 (N_14609,N_10838,N_10989);
xnor U14610 (N_14610,N_9418,N_12197);
nand U14611 (N_14611,N_11815,N_11276);
xor U14612 (N_14612,N_12235,N_9962);
nor U14613 (N_14613,N_12257,N_12058);
or U14614 (N_14614,N_9943,N_11940);
nand U14615 (N_14615,N_10023,N_12040);
nor U14616 (N_14616,N_10960,N_10562);
nor U14617 (N_14617,N_9710,N_10258);
nand U14618 (N_14618,N_9785,N_10389);
xor U14619 (N_14619,N_11474,N_10999);
nor U14620 (N_14620,N_9924,N_11063);
xnor U14621 (N_14621,N_12036,N_11936);
nor U14622 (N_14622,N_12435,N_10461);
nor U14623 (N_14623,N_10384,N_10176);
nand U14624 (N_14624,N_12352,N_9637);
nor U14625 (N_14625,N_10383,N_10710);
and U14626 (N_14626,N_11421,N_10205);
nor U14627 (N_14627,N_10598,N_12435);
and U14628 (N_14628,N_10070,N_11666);
xor U14629 (N_14629,N_11616,N_10127);
nor U14630 (N_14630,N_10944,N_9459);
nor U14631 (N_14631,N_11176,N_12275);
xor U14632 (N_14632,N_10802,N_10719);
or U14633 (N_14633,N_10569,N_9988);
or U14634 (N_14634,N_9440,N_11030);
xor U14635 (N_14635,N_10078,N_11283);
or U14636 (N_14636,N_10333,N_11036);
nand U14637 (N_14637,N_11973,N_9489);
nor U14638 (N_14638,N_9692,N_11257);
nand U14639 (N_14639,N_10657,N_11080);
or U14640 (N_14640,N_11181,N_11346);
nand U14641 (N_14641,N_10506,N_11654);
nand U14642 (N_14642,N_11756,N_9483);
nand U14643 (N_14643,N_9574,N_11444);
nor U14644 (N_14644,N_9565,N_10246);
xor U14645 (N_14645,N_11768,N_10207);
nand U14646 (N_14646,N_11311,N_11558);
and U14647 (N_14647,N_10520,N_11509);
xnor U14648 (N_14648,N_11021,N_11669);
nand U14649 (N_14649,N_10890,N_12417);
and U14650 (N_14650,N_10644,N_9922);
and U14651 (N_14651,N_11799,N_11674);
nand U14652 (N_14652,N_12190,N_12284);
nor U14653 (N_14653,N_10396,N_11289);
or U14654 (N_14654,N_10025,N_9814);
or U14655 (N_14655,N_9917,N_11494);
xor U14656 (N_14656,N_11644,N_10808);
xnor U14657 (N_14657,N_9451,N_12007);
or U14658 (N_14658,N_10343,N_11031);
nor U14659 (N_14659,N_9465,N_11878);
or U14660 (N_14660,N_11886,N_10666);
and U14661 (N_14661,N_10814,N_9846);
xnor U14662 (N_14662,N_12455,N_11657);
xor U14663 (N_14663,N_9691,N_10980);
nor U14664 (N_14664,N_10744,N_12199);
or U14665 (N_14665,N_10249,N_10464);
or U14666 (N_14666,N_10771,N_10844);
nor U14667 (N_14667,N_9801,N_9486);
nand U14668 (N_14668,N_12382,N_11470);
xor U14669 (N_14669,N_12407,N_12239);
and U14670 (N_14670,N_11240,N_10326);
nor U14671 (N_14671,N_9858,N_10406);
nor U14672 (N_14672,N_10735,N_12462);
and U14673 (N_14673,N_11597,N_9668);
xnor U14674 (N_14674,N_9567,N_11348);
or U14675 (N_14675,N_10257,N_10283);
or U14676 (N_14676,N_10623,N_9813);
and U14677 (N_14677,N_10917,N_12321);
nor U14678 (N_14678,N_11358,N_11598);
and U14679 (N_14679,N_10008,N_11041);
xor U14680 (N_14680,N_9557,N_11392);
and U14681 (N_14681,N_9980,N_9899);
and U14682 (N_14682,N_9519,N_11877);
or U14683 (N_14683,N_11833,N_11578);
nor U14684 (N_14684,N_10947,N_12176);
nor U14685 (N_14685,N_11226,N_11544);
nor U14686 (N_14686,N_10708,N_11974);
xnor U14687 (N_14687,N_11671,N_11411);
or U14688 (N_14688,N_9669,N_11133);
and U14689 (N_14689,N_10835,N_10162);
xor U14690 (N_14690,N_9459,N_11387);
nor U14691 (N_14691,N_11522,N_10379);
nor U14692 (N_14692,N_10002,N_9734);
or U14693 (N_14693,N_10098,N_11872);
or U14694 (N_14694,N_12217,N_10928);
xor U14695 (N_14695,N_11721,N_11790);
nor U14696 (N_14696,N_11204,N_12036);
or U14697 (N_14697,N_10114,N_9991);
nand U14698 (N_14698,N_11284,N_10662);
or U14699 (N_14699,N_11600,N_11700);
or U14700 (N_14700,N_9648,N_11819);
nor U14701 (N_14701,N_12410,N_9704);
and U14702 (N_14702,N_12189,N_12055);
and U14703 (N_14703,N_10283,N_12311);
and U14704 (N_14704,N_9869,N_10101);
nand U14705 (N_14705,N_10759,N_11197);
nand U14706 (N_14706,N_10971,N_10681);
xor U14707 (N_14707,N_11647,N_9999);
and U14708 (N_14708,N_10648,N_10026);
nor U14709 (N_14709,N_10004,N_11592);
xor U14710 (N_14710,N_9662,N_11954);
and U14711 (N_14711,N_11974,N_9611);
or U14712 (N_14712,N_12062,N_9895);
and U14713 (N_14713,N_10482,N_9669);
xor U14714 (N_14714,N_11350,N_9639);
or U14715 (N_14715,N_11785,N_11004);
xnor U14716 (N_14716,N_11750,N_9590);
or U14717 (N_14717,N_9511,N_10374);
or U14718 (N_14718,N_11650,N_9527);
xnor U14719 (N_14719,N_9989,N_11560);
xnor U14720 (N_14720,N_12357,N_12269);
and U14721 (N_14721,N_10851,N_12424);
xnor U14722 (N_14722,N_11350,N_10189);
nand U14723 (N_14723,N_11171,N_12457);
nand U14724 (N_14724,N_9882,N_10474);
nand U14725 (N_14725,N_12458,N_12189);
xor U14726 (N_14726,N_12473,N_10967);
or U14727 (N_14727,N_10843,N_11082);
or U14728 (N_14728,N_9438,N_9559);
xor U14729 (N_14729,N_10819,N_9721);
and U14730 (N_14730,N_10142,N_9466);
and U14731 (N_14731,N_10620,N_10611);
and U14732 (N_14732,N_10840,N_12376);
xor U14733 (N_14733,N_10056,N_9860);
and U14734 (N_14734,N_9718,N_12403);
and U14735 (N_14735,N_9428,N_10044);
or U14736 (N_14736,N_12462,N_11320);
and U14737 (N_14737,N_9893,N_10936);
nand U14738 (N_14738,N_12234,N_12422);
and U14739 (N_14739,N_9942,N_12162);
nand U14740 (N_14740,N_11617,N_11142);
xor U14741 (N_14741,N_11925,N_9620);
nor U14742 (N_14742,N_11535,N_9599);
nand U14743 (N_14743,N_12281,N_10050);
or U14744 (N_14744,N_10023,N_12294);
nand U14745 (N_14745,N_10001,N_10823);
xor U14746 (N_14746,N_11392,N_10749);
nor U14747 (N_14747,N_10354,N_10906);
or U14748 (N_14748,N_9408,N_12206);
nand U14749 (N_14749,N_10273,N_11574);
nor U14750 (N_14750,N_11971,N_10282);
nor U14751 (N_14751,N_9848,N_11613);
nor U14752 (N_14752,N_10037,N_10023);
or U14753 (N_14753,N_9664,N_9773);
nor U14754 (N_14754,N_10764,N_9568);
nor U14755 (N_14755,N_12456,N_10242);
and U14756 (N_14756,N_9750,N_10034);
or U14757 (N_14757,N_12388,N_10052);
xnor U14758 (N_14758,N_11172,N_11954);
nor U14759 (N_14759,N_12318,N_9458);
nor U14760 (N_14760,N_11914,N_9413);
nand U14761 (N_14761,N_10612,N_12265);
nor U14762 (N_14762,N_10047,N_12170);
xor U14763 (N_14763,N_10980,N_11495);
nor U14764 (N_14764,N_11149,N_9502);
nand U14765 (N_14765,N_10222,N_10071);
xor U14766 (N_14766,N_11930,N_11265);
or U14767 (N_14767,N_9553,N_12363);
and U14768 (N_14768,N_11466,N_9976);
nor U14769 (N_14769,N_10256,N_11355);
or U14770 (N_14770,N_11395,N_10760);
nand U14771 (N_14771,N_10300,N_9389);
xor U14772 (N_14772,N_10602,N_10036);
nor U14773 (N_14773,N_10701,N_11158);
nand U14774 (N_14774,N_11540,N_9552);
xnor U14775 (N_14775,N_11863,N_11435);
and U14776 (N_14776,N_10236,N_9613);
or U14777 (N_14777,N_11222,N_10642);
nor U14778 (N_14778,N_10195,N_9687);
nor U14779 (N_14779,N_10600,N_11519);
and U14780 (N_14780,N_9585,N_12068);
nor U14781 (N_14781,N_10451,N_12066);
nand U14782 (N_14782,N_11390,N_12343);
or U14783 (N_14783,N_10962,N_11583);
xnor U14784 (N_14784,N_10468,N_10993);
or U14785 (N_14785,N_12380,N_10218);
and U14786 (N_14786,N_11213,N_11461);
nand U14787 (N_14787,N_10360,N_10643);
nor U14788 (N_14788,N_10706,N_11886);
or U14789 (N_14789,N_10291,N_10032);
nor U14790 (N_14790,N_10174,N_10976);
or U14791 (N_14791,N_10842,N_12322);
xor U14792 (N_14792,N_10089,N_11276);
xnor U14793 (N_14793,N_11651,N_9680);
nor U14794 (N_14794,N_11340,N_9996);
and U14795 (N_14795,N_11312,N_11677);
and U14796 (N_14796,N_9487,N_12472);
xnor U14797 (N_14797,N_10230,N_10388);
or U14798 (N_14798,N_11487,N_10313);
and U14799 (N_14799,N_10443,N_10455);
nand U14800 (N_14800,N_11400,N_10806);
or U14801 (N_14801,N_11573,N_11264);
xor U14802 (N_14802,N_12097,N_11027);
nor U14803 (N_14803,N_11133,N_9809);
nor U14804 (N_14804,N_9745,N_10914);
xnor U14805 (N_14805,N_9947,N_10546);
and U14806 (N_14806,N_12056,N_9510);
and U14807 (N_14807,N_10175,N_11260);
xor U14808 (N_14808,N_10104,N_10442);
nor U14809 (N_14809,N_10399,N_12298);
xnor U14810 (N_14810,N_11665,N_10256);
or U14811 (N_14811,N_11607,N_12396);
or U14812 (N_14812,N_9839,N_10654);
and U14813 (N_14813,N_11353,N_11746);
and U14814 (N_14814,N_11921,N_10117);
nand U14815 (N_14815,N_11329,N_10600);
or U14816 (N_14816,N_10198,N_11532);
or U14817 (N_14817,N_12232,N_11182);
nand U14818 (N_14818,N_10821,N_10371);
xor U14819 (N_14819,N_11946,N_12301);
xnor U14820 (N_14820,N_10347,N_11123);
nor U14821 (N_14821,N_11308,N_9978);
nor U14822 (N_14822,N_12261,N_11138);
xor U14823 (N_14823,N_11878,N_11979);
nand U14824 (N_14824,N_10171,N_9826);
and U14825 (N_14825,N_11968,N_11981);
xor U14826 (N_14826,N_10047,N_9518);
nor U14827 (N_14827,N_9832,N_11707);
and U14828 (N_14828,N_10860,N_9952);
xnor U14829 (N_14829,N_10769,N_10326);
nor U14830 (N_14830,N_10121,N_12438);
and U14831 (N_14831,N_10562,N_11246);
nor U14832 (N_14832,N_10086,N_12255);
and U14833 (N_14833,N_10762,N_9840);
xnor U14834 (N_14834,N_12418,N_11155);
and U14835 (N_14835,N_11346,N_11516);
xnor U14836 (N_14836,N_12340,N_10410);
or U14837 (N_14837,N_11777,N_10492);
or U14838 (N_14838,N_12159,N_11348);
nand U14839 (N_14839,N_11496,N_11719);
nor U14840 (N_14840,N_10703,N_10141);
nand U14841 (N_14841,N_10394,N_11999);
nand U14842 (N_14842,N_11101,N_9966);
nand U14843 (N_14843,N_12225,N_11686);
and U14844 (N_14844,N_10939,N_9435);
nand U14845 (N_14845,N_11991,N_11370);
xnor U14846 (N_14846,N_9660,N_9776);
xor U14847 (N_14847,N_12103,N_10710);
and U14848 (N_14848,N_10986,N_9541);
nand U14849 (N_14849,N_11536,N_12237);
nand U14850 (N_14850,N_9710,N_9833);
nor U14851 (N_14851,N_11195,N_9554);
and U14852 (N_14852,N_10344,N_9392);
nor U14853 (N_14853,N_11430,N_10866);
nand U14854 (N_14854,N_10113,N_12447);
or U14855 (N_14855,N_10254,N_11153);
xnor U14856 (N_14856,N_9824,N_10263);
or U14857 (N_14857,N_11241,N_10573);
xor U14858 (N_14858,N_11405,N_11270);
xnor U14859 (N_14859,N_9765,N_10357);
nand U14860 (N_14860,N_11093,N_9714);
and U14861 (N_14861,N_11212,N_9976);
or U14862 (N_14862,N_10123,N_11221);
or U14863 (N_14863,N_9600,N_9961);
nand U14864 (N_14864,N_12224,N_11347);
or U14865 (N_14865,N_12323,N_9628);
xnor U14866 (N_14866,N_12064,N_12016);
nor U14867 (N_14867,N_10625,N_9854);
or U14868 (N_14868,N_12215,N_10069);
or U14869 (N_14869,N_11375,N_10297);
nand U14870 (N_14870,N_10502,N_10698);
xor U14871 (N_14871,N_10269,N_10432);
or U14872 (N_14872,N_12473,N_9964);
nand U14873 (N_14873,N_12430,N_9844);
xor U14874 (N_14874,N_12126,N_9892);
nor U14875 (N_14875,N_10342,N_10357);
nor U14876 (N_14876,N_12260,N_10439);
nor U14877 (N_14877,N_10441,N_10644);
or U14878 (N_14878,N_9793,N_9606);
nand U14879 (N_14879,N_12471,N_10021);
or U14880 (N_14880,N_11895,N_11398);
xnor U14881 (N_14881,N_12329,N_10131);
nor U14882 (N_14882,N_10130,N_10597);
and U14883 (N_14883,N_10921,N_10751);
xor U14884 (N_14884,N_12076,N_10399);
xnor U14885 (N_14885,N_9579,N_10550);
nand U14886 (N_14886,N_10716,N_9391);
nor U14887 (N_14887,N_9523,N_11716);
nand U14888 (N_14888,N_9789,N_12049);
xor U14889 (N_14889,N_11743,N_11831);
xnor U14890 (N_14890,N_10640,N_10238);
or U14891 (N_14891,N_12422,N_10668);
nor U14892 (N_14892,N_11327,N_11635);
xnor U14893 (N_14893,N_10023,N_11151);
nand U14894 (N_14894,N_10923,N_10904);
and U14895 (N_14895,N_10365,N_10853);
xnor U14896 (N_14896,N_10250,N_9715);
nand U14897 (N_14897,N_9850,N_9781);
or U14898 (N_14898,N_10280,N_9890);
xor U14899 (N_14899,N_10631,N_12238);
xor U14900 (N_14900,N_12205,N_10446);
xor U14901 (N_14901,N_10644,N_12167);
and U14902 (N_14902,N_10614,N_9847);
nand U14903 (N_14903,N_10797,N_11508);
nor U14904 (N_14904,N_10902,N_12499);
nor U14905 (N_14905,N_10724,N_9381);
or U14906 (N_14906,N_9645,N_9924);
nand U14907 (N_14907,N_11603,N_9465);
xor U14908 (N_14908,N_11740,N_10912);
nand U14909 (N_14909,N_11447,N_11786);
or U14910 (N_14910,N_10800,N_11971);
nor U14911 (N_14911,N_11429,N_11472);
nand U14912 (N_14912,N_12162,N_10683);
nor U14913 (N_14913,N_9978,N_9772);
and U14914 (N_14914,N_11789,N_10734);
or U14915 (N_14915,N_9991,N_11508);
xnor U14916 (N_14916,N_10745,N_9876);
xnor U14917 (N_14917,N_11865,N_10998);
xnor U14918 (N_14918,N_11231,N_9526);
xnor U14919 (N_14919,N_10551,N_9995);
nand U14920 (N_14920,N_11490,N_9704);
and U14921 (N_14921,N_10351,N_9868);
and U14922 (N_14922,N_9762,N_11382);
and U14923 (N_14923,N_10107,N_10685);
nor U14924 (N_14924,N_11024,N_11729);
or U14925 (N_14925,N_12210,N_11952);
and U14926 (N_14926,N_12304,N_11263);
nand U14927 (N_14927,N_9525,N_12379);
nand U14928 (N_14928,N_12213,N_9744);
nor U14929 (N_14929,N_9586,N_10182);
or U14930 (N_14930,N_10739,N_11009);
and U14931 (N_14931,N_10977,N_11980);
or U14932 (N_14932,N_10240,N_9813);
and U14933 (N_14933,N_11156,N_11672);
or U14934 (N_14934,N_9662,N_11755);
or U14935 (N_14935,N_11210,N_9720);
xnor U14936 (N_14936,N_10599,N_11192);
and U14937 (N_14937,N_9797,N_11691);
or U14938 (N_14938,N_11884,N_11848);
or U14939 (N_14939,N_9656,N_10338);
or U14940 (N_14940,N_9626,N_10221);
and U14941 (N_14941,N_11487,N_10682);
nor U14942 (N_14942,N_9500,N_11696);
nand U14943 (N_14943,N_12025,N_12375);
and U14944 (N_14944,N_10230,N_11657);
xor U14945 (N_14945,N_11896,N_10187);
nand U14946 (N_14946,N_10048,N_9491);
and U14947 (N_14947,N_12231,N_10220);
or U14948 (N_14948,N_10241,N_10449);
and U14949 (N_14949,N_10416,N_12193);
or U14950 (N_14950,N_10169,N_9428);
or U14951 (N_14951,N_12306,N_12255);
xnor U14952 (N_14952,N_10457,N_11671);
nand U14953 (N_14953,N_12438,N_10600);
and U14954 (N_14954,N_9639,N_9990);
or U14955 (N_14955,N_10304,N_11572);
nor U14956 (N_14956,N_10166,N_12383);
and U14957 (N_14957,N_9393,N_11217);
or U14958 (N_14958,N_11268,N_12171);
nand U14959 (N_14959,N_11663,N_9382);
nor U14960 (N_14960,N_12400,N_12458);
and U14961 (N_14961,N_9712,N_9873);
nor U14962 (N_14962,N_10211,N_11604);
xor U14963 (N_14963,N_9597,N_10906);
and U14964 (N_14964,N_11181,N_10488);
or U14965 (N_14965,N_11760,N_9654);
or U14966 (N_14966,N_11143,N_12316);
or U14967 (N_14967,N_11268,N_11692);
and U14968 (N_14968,N_9440,N_11549);
xor U14969 (N_14969,N_11876,N_11223);
xnor U14970 (N_14970,N_10218,N_12289);
and U14971 (N_14971,N_11603,N_11950);
or U14972 (N_14972,N_10683,N_12154);
nand U14973 (N_14973,N_10577,N_11164);
nand U14974 (N_14974,N_10502,N_10460);
xnor U14975 (N_14975,N_9515,N_11561);
or U14976 (N_14976,N_9796,N_10037);
nor U14977 (N_14977,N_11481,N_10893);
nand U14978 (N_14978,N_11527,N_10992);
xor U14979 (N_14979,N_11517,N_11299);
xnor U14980 (N_14980,N_11867,N_10011);
xor U14981 (N_14981,N_11905,N_11026);
or U14982 (N_14982,N_10751,N_9651);
and U14983 (N_14983,N_10024,N_11568);
and U14984 (N_14984,N_11442,N_10765);
and U14985 (N_14985,N_9639,N_10487);
xor U14986 (N_14986,N_10555,N_9432);
and U14987 (N_14987,N_11203,N_11193);
nand U14988 (N_14988,N_9528,N_10387);
xnor U14989 (N_14989,N_12004,N_11152);
nor U14990 (N_14990,N_11447,N_12406);
xor U14991 (N_14991,N_10006,N_10354);
nand U14992 (N_14992,N_10826,N_10975);
and U14993 (N_14993,N_12008,N_10319);
nand U14994 (N_14994,N_9423,N_10777);
or U14995 (N_14995,N_10205,N_10739);
xnor U14996 (N_14996,N_11419,N_11944);
xnor U14997 (N_14997,N_11473,N_10828);
or U14998 (N_14998,N_10154,N_9384);
or U14999 (N_14999,N_11123,N_11084);
or U15000 (N_15000,N_9972,N_12233);
or U15001 (N_15001,N_11665,N_9517);
or U15002 (N_15002,N_9584,N_10162);
nor U15003 (N_15003,N_9885,N_12039);
or U15004 (N_15004,N_11064,N_10346);
xnor U15005 (N_15005,N_11242,N_10061);
and U15006 (N_15006,N_9941,N_9663);
or U15007 (N_15007,N_11832,N_11895);
nand U15008 (N_15008,N_10169,N_9929);
and U15009 (N_15009,N_11542,N_9549);
nor U15010 (N_15010,N_11230,N_10827);
and U15011 (N_15011,N_12448,N_12400);
nand U15012 (N_15012,N_10224,N_11229);
nor U15013 (N_15013,N_10701,N_9642);
xnor U15014 (N_15014,N_11192,N_10776);
nor U15015 (N_15015,N_9569,N_9643);
xor U15016 (N_15016,N_9619,N_10246);
xnor U15017 (N_15017,N_9434,N_9796);
nand U15018 (N_15018,N_12009,N_11857);
and U15019 (N_15019,N_9905,N_10865);
and U15020 (N_15020,N_10960,N_11468);
or U15021 (N_15021,N_12458,N_10329);
xnor U15022 (N_15022,N_12124,N_10262);
and U15023 (N_15023,N_11797,N_11117);
xor U15024 (N_15024,N_11046,N_9795);
xor U15025 (N_15025,N_10244,N_11912);
xor U15026 (N_15026,N_12420,N_12257);
nor U15027 (N_15027,N_10395,N_11969);
nand U15028 (N_15028,N_10406,N_11958);
xor U15029 (N_15029,N_10497,N_9831);
xor U15030 (N_15030,N_12070,N_11316);
and U15031 (N_15031,N_10575,N_10271);
and U15032 (N_15032,N_10794,N_11257);
nor U15033 (N_15033,N_12106,N_9991);
nor U15034 (N_15034,N_12075,N_10022);
nand U15035 (N_15035,N_11225,N_11001);
xor U15036 (N_15036,N_10726,N_9483);
and U15037 (N_15037,N_10255,N_11720);
nand U15038 (N_15038,N_11367,N_10615);
nor U15039 (N_15039,N_11040,N_10422);
nor U15040 (N_15040,N_12204,N_9820);
or U15041 (N_15041,N_11611,N_10792);
xnor U15042 (N_15042,N_11325,N_10766);
nor U15043 (N_15043,N_9780,N_12446);
and U15044 (N_15044,N_10980,N_9988);
or U15045 (N_15045,N_12320,N_9790);
and U15046 (N_15046,N_11484,N_10686);
and U15047 (N_15047,N_9796,N_10472);
xnor U15048 (N_15048,N_12361,N_11618);
xor U15049 (N_15049,N_12377,N_11877);
or U15050 (N_15050,N_10770,N_10435);
or U15051 (N_15051,N_10776,N_10112);
and U15052 (N_15052,N_9423,N_9974);
nor U15053 (N_15053,N_9604,N_9772);
nand U15054 (N_15054,N_11388,N_11572);
xnor U15055 (N_15055,N_10258,N_9633);
and U15056 (N_15056,N_10072,N_10093);
nand U15057 (N_15057,N_11738,N_10174);
nand U15058 (N_15058,N_12103,N_10805);
nor U15059 (N_15059,N_11872,N_9979);
or U15060 (N_15060,N_9525,N_10370);
nand U15061 (N_15061,N_9995,N_12279);
xnor U15062 (N_15062,N_9706,N_9778);
and U15063 (N_15063,N_10423,N_9750);
xnor U15064 (N_15064,N_9479,N_11797);
nor U15065 (N_15065,N_10828,N_10657);
nand U15066 (N_15066,N_9594,N_10586);
xnor U15067 (N_15067,N_11310,N_12429);
or U15068 (N_15068,N_11519,N_12295);
xor U15069 (N_15069,N_9404,N_10667);
nor U15070 (N_15070,N_12011,N_10442);
or U15071 (N_15071,N_10962,N_11430);
or U15072 (N_15072,N_10279,N_12314);
xor U15073 (N_15073,N_10412,N_11095);
nand U15074 (N_15074,N_10455,N_9859);
nand U15075 (N_15075,N_12260,N_11567);
and U15076 (N_15076,N_9587,N_10704);
and U15077 (N_15077,N_11317,N_11425);
and U15078 (N_15078,N_11152,N_11170);
and U15079 (N_15079,N_11347,N_11951);
nor U15080 (N_15080,N_9377,N_10895);
nor U15081 (N_15081,N_10079,N_11872);
or U15082 (N_15082,N_11962,N_10831);
xnor U15083 (N_15083,N_11938,N_12406);
and U15084 (N_15084,N_11609,N_11982);
xor U15085 (N_15085,N_10599,N_10895);
or U15086 (N_15086,N_10493,N_10214);
and U15087 (N_15087,N_11102,N_11251);
nand U15088 (N_15088,N_10195,N_10885);
xor U15089 (N_15089,N_11929,N_9718);
nor U15090 (N_15090,N_10871,N_10538);
nand U15091 (N_15091,N_11735,N_9721);
and U15092 (N_15092,N_12232,N_11900);
nor U15093 (N_15093,N_11070,N_12045);
and U15094 (N_15094,N_11766,N_10856);
nor U15095 (N_15095,N_11774,N_9427);
nand U15096 (N_15096,N_10606,N_11059);
nand U15097 (N_15097,N_11159,N_10554);
or U15098 (N_15098,N_10957,N_9399);
nand U15099 (N_15099,N_10181,N_9778);
or U15100 (N_15100,N_12401,N_9418);
or U15101 (N_15101,N_10510,N_10962);
xor U15102 (N_15102,N_9423,N_11745);
nor U15103 (N_15103,N_12286,N_10558);
xor U15104 (N_15104,N_9940,N_10133);
xnor U15105 (N_15105,N_11659,N_11902);
nand U15106 (N_15106,N_10113,N_9811);
xnor U15107 (N_15107,N_11155,N_9510);
or U15108 (N_15108,N_9949,N_10124);
and U15109 (N_15109,N_10536,N_9564);
or U15110 (N_15110,N_9998,N_9447);
xnor U15111 (N_15111,N_9414,N_12160);
xnor U15112 (N_15112,N_10557,N_10383);
and U15113 (N_15113,N_10309,N_10217);
nand U15114 (N_15114,N_9435,N_9625);
and U15115 (N_15115,N_9601,N_10616);
or U15116 (N_15116,N_11889,N_10317);
nor U15117 (N_15117,N_9383,N_12422);
nand U15118 (N_15118,N_11461,N_12434);
nor U15119 (N_15119,N_12157,N_10137);
and U15120 (N_15120,N_11174,N_11262);
nor U15121 (N_15121,N_12216,N_11766);
and U15122 (N_15122,N_10910,N_11232);
xnor U15123 (N_15123,N_11277,N_9433);
nor U15124 (N_15124,N_11127,N_9964);
and U15125 (N_15125,N_9550,N_10896);
and U15126 (N_15126,N_10438,N_10647);
nor U15127 (N_15127,N_10892,N_9876);
nand U15128 (N_15128,N_10935,N_11301);
nor U15129 (N_15129,N_11782,N_10847);
xnor U15130 (N_15130,N_9906,N_11759);
nor U15131 (N_15131,N_11585,N_11404);
xnor U15132 (N_15132,N_10285,N_11516);
or U15133 (N_15133,N_10456,N_11829);
nand U15134 (N_15134,N_12272,N_11618);
xor U15135 (N_15135,N_12113,N_9873);
and U15136 (N_15136,N_12256,N_10083);
or U15137 (N_15137,N_11206,N_9518);
or U15138 (N_15138,N_12165,N_11565);
nand U15139 (N_15139,N_12491,N_10564);
nor U15140 (N_15140,N_12208,N_11964);
nand U15141 (N_15141,N_10903,N_11773);
and U15142 (N_15142,N_9903,N_11968);
or U15143 (N_15143,N_11845,N_11554);
nand U15144 (N_15144,N_12424,N_10709);
nor U15145 (N_15145,N_10465,N_11270);
nand U15146 (N_15146,N_11734,N_9793);
or U15147 (N_15147,N_10154,N_10204);
or U15148 (N_15148,N_12102,N_9451);
or U15149 (N_15149,N_12369,N_11962);
xor U15150 (N_15150,N_12173,N_10199);
nor U15151 (N_15151,N_10436,N_11969);
xor U15152 (N_15152,N_12456,N_10908);
or U15153 (N_15153,N_10683,N_9619);
nand U15154 (N_15154,N_10779,N_10171);
or U15155 (N_15155,N_10730,N_12402);
xor U15156 (N_15156,N_11745,N_9730);
and U15157 (N_15157,N_12013,N_11979);
xnor U15158 (N_15158,N_9555,N_12474);
nand U15159 (N_15159,N_11141,N_10520);
and U15160 (N_15160,N_9612,N_11700);
or U15161 (N_15161,N_12452,N_11516);
or U15162 (N_15162,N_12030,N_10140);
or U15163 (N_15163,N_11465,N_12307);
xnor U15164 (N_15164,N_10569,N_11105);
and U15165 (N_15165,N_10808,N_9664);
and U15166 (N_15166,N_10047,N_10879);
or U15167 (N_15167,N_9621,N_9542);
nand U15168 (N_15168,N_11182,N_11726);
nand U15169 (N_15169,N_10067,N_9762);
xnor U15170 (N_15170,N_10037,N_10891);
nand U15171 (N_15171,N_11288,N_10315);
or U15172 (N_15172,N_10803,N_11107);
and U15173 (N_15173,N_12002,N_11244);
nand U15174 (N_15174,N_9967,N_9661);
xor U15175 (N_15175,N_9643,N_11345);
xor U15176 (N_15176,N_10154,N_11345);
nand U15177 (N_15177,N_10211,N_11869);
nor U15178 (N_15178,N_12011,N_10679);
nor U15179 (N_15179,N_12348,N_10025);
or U15180 (N_15180,N_10731,N_9658);
or U15181 (N_15181,N_12373,N_12328);
nor U15182 (N_15182,N_11447,N_10171);
or U15183 (N_15183,N_12262,N_10832);
nand U15184 (N_15184,N_12270,N_11862);
nor U15185 (N_15185,N_11018,N_12175);
or U15186 (N_15186,N_12372,N_10981);
and U15187 (N_15187,N_11340,N_9544);
nor U15188 (N_15188,N_12384,N_10955);
xnor U15189 (N_15189,N_9594,N_11741);
nand U15190 (N_15190,N_11048,N_11927);
nand U15191 (N_15191,N_9551,N_10609);
and U15192 (N_15192,N_12474,N_11804);
or U15193 (N_15193,N_10018,N_10325);
and U15194 (N_15194,N_11995,N_10245);
and U15195 (N_15195,N_11128,N_11379);
nand U15196 (N_15196,N_11300,N_10514);
xor U15197 (N_15197,N_10810,N_9504);
nor U15198 (N_15198,N_11098,N_9389);
and U15199 (N_15199,N_9737,N_9819);
or U15200 (N_15200,N_9954,N_10741);
nor U15201 (N_15201,N_11775,N_9676);
or U15202 (N_15202,N_10081,N_11399);
and U15203 (N_15203,N_11204,N_10540);
nand U15204 (N_15204,N_9991,N_12455);
nor U15205 (N_15205,N_11467,N_12416);
xnor U15206 (N_15206,N_11323,N_11819);
or U15207 (N_15207,N_11319,N_12445);
and U15208 (N_15208,N_12322,N_9697);
and U15209 (N_15209,N_12440,N_11326);
xnor U15210 (N_15210,N_11169,N_9524);
and U15211 (N_15211,N_10768,N_11489);
or U15212 (N_15212,N_10065,N_9824);
xor U15213 (N_15213,N_9945,N_11334);
and U15214 (N_15214,N_11361,N_11486);
nor U15215 (N_15215,N_9473,N_11489);
nor U15216 (N_15216,N_12156,N_11909);
and U15217 (N_15217,N_11442,N_10706);
or U15218 (N_15218,N_12015,N_12205);
xor U15219 (N_15219,N_9699,N_11042);
and U15220 (N_15220,N_11924,N_10724);
nand U15221 (N_15221,N_12236,N_10818);
xor U15222 (N_15222,N_9742,N_11999);
nor U15223 (N_15223,N_12192,N_9470);
nor U15224 (N_15224,N_10999,N_9746);
or U15225 (N_15225,N_11263,N_11125);
or U15226 (N_15226,N_11805,N_10791);
or U15227 (N_15227,N_9628,N_10429);
xor U15228 (N_15228,N_11026,N_10205);
xor U15229 (N_15229,N_10349,N_12450);
xor U15230 (N_15230,N_11077,N_11011);
or U15231 (N_15231,N_11223,N_10594);
xor U15232 (N_15232,N_11609,N_10393);
and U15233 (N_15233,N_10928,N_10031);
xor U15234 (N_15234,N_10253,N_10920);
nand U15235 (N_15235,N_10476,N_12272);
or U15236 (N_15236,N_11292,N_11039);
nor U15237 (N_15237,N_10171,N_10696);
and U15238 (N_15238,N_11882,N_11528);
nand U15239 (N_15239,N_11747,N_11620);
nand U15240 (N_15240,N_12126,N_10428);
nand U15241 (N_15241,N_11423,N_11730);
xor U15242 (N_15242,N_12285,N_9683);
or U15243 (N_15243,N_9810,N_10135);
and U15244 (N_15244,N_10154,N_10665);
nand U15245 (N_15245,N_9775,N_11865);
nand U15246 (N_15246,N_10090,N_10559);
nand U15247 (N_15247,N_11383,N_11332);
nand U15248 (N_15248,N_11738,N_11125);
xor U15249 (N_15249,N_10483,N_10666);
xnor U15250 (N_15250,N_10342,N_11753);
or U15251 (N_15251,N_9971,N_11620);
and U15252 (N_15252,N_12460,N_10499);
xnor U15253 (N_15253,N_9978,N_11552);
xor U15254 (N_15254,N_11904,N_12380);
nand U15255 (N_15255,N_12293,N_10171);
nand U15256 (N_15256,N_12222,N_11996);
xor U15257 (N_15257,N_10939,N_12422);
nor U15258 (N_15258,N_11291,N_10690);
and U15259 (N_15259,N_12012,N_11041);
nor U15260 (N_15260,N_10480,N_11778);
nor U15261 (N_15261,N_9500,N_11074);
nor U15262 (N_15262,N_11319,N_9452);
nand U15263 (N_15263,N_12388,N_10332);
and U15264 (N_15264,N_10194,N_12048);
nand U15265 (N_15265,N_12445,N_12340);
nand U15266 (N_15266,N_9733,N_12164);
or U15267 (N_15267,N_12280,N_11526);
nand U15268 (N_15268,N_10843,N_9582);
or U15269 (N_15269,N_10314,N_12296);
nand U15270 (N_15270,N_9596,N_12144);
nor U15271 (N_15271,N_9644,N_10880);
nand U15272 (N_15272,N_10854,N_10383);
and U15273 (N_15273,N_11090,N_10902);
xor U15274 (N_15274,N_11298,N_10216);
nor U15275 (N_15275,N_10493,N_11755);
xor U15276 (N_15276,N_9969,N_9668);
nand U15277 (N_15277,N_10565,N_10977);
and U15278 (N_15278,N_10375,N_9508);
nand U15279 (N_15279,N_9687,N_9915);
or U15280 (N_15280,N_11938,N_10582);
xor U15281 (N_15281,N_11691,N_11426);
nand U15282 (N_15282,N_10279,N_9527);
nand U15283 (N_15283,N_10685,N_9861);
xor U15284 (N_15284,N_10736,N_10994);
nor U15285 (N_15285,N_12432,N_9518);
xor U15286 (N_15286,N_9760,N_11876);
nand U15287 (N_15287,N_12358,N_10009);
nor U15288 (N_15288,N_12379,N_10451);
and U15289 (N_15289,N_10007,N_11020);
or U15290 (N_15290,N_11054,N_10373);
and U15291 (N_15291,N_12259,N_11216);
and U15292 (N_15292,N_10696,N_12469);
nor U15293 (N_15293,N_12033,N_10129);
xnor U15294 (N_15294,N_11052,N_11392);
and U15295 (N_15295,N_9983,N_9561);
and U15296 (N_15296,N_9718,N_10907);
nand U15297 (N_15297,N_11744,N_12178);
and U15298 (N_15298,N_9945,N_12298);
nand U15299 (N_15299,N_11641,N_10920);
nor U15300 (N_15300,N_10356,N_10613);
and U15301 (N_15301,N_9792,N_11476);
nand U15302 (N_15302,N_11741,N_10679);
nand U15303 (N_15303,N_10917,N_10759);
nor U15304 (N_15304,N_9611,N_9397);
xnor U15305 (N_15305,N_11913,N_9699);
xor U15306 (N_15306,N_11037,N_11744);
nor U15307 (N_15307,N_12163,N_10364);
and U15308 (N_15308,N_10294,N_10366);
xor U15309 (N_15309,N_9498,N_12035);
or U15310 (N_15310,N_11385,N_10473);
nand U15311 (N_15311,N_10767,N_11577);
xor U15312 (N_15312,N_10505,N_9385);
and U15313 (N_15313,N_9576,N_9679);
and U15314 (N_15314,N_11492,N_11652);
xor U15315 (N_15315,N_10693,N_10546);
or U15316 (N_15316,N_10371,N_9809);
xnor U15317 (N_15317,N_11275,N_11199);
and U15318 (N_15318,N_10028,N_9781);
nand U15319 (N_15319,N_11937,N_10098);
nor U15320 (N_15320,N_12147,N_10897);
or U15321 (N_15321,N_10847,N_10844);
or U15322 (N_15322,N_9616,N_12026);
nand U15323 (N_15323,N_11726,N_10211);
or U15324 (N_15324,N_10071,N_11939);
nand U15325 (N_15325,N_10791,N_12199);
xor U15326 (N_15326,N_9858,N_10531);
xnor U15327 (N_15327,N_11918,N_9689);
or U15328 (N_15328,N_10266,N_10912);
nor U15329 (N_15329,N_10473,N_10663);
and U15330 (N_15330,N_10639,N_11069);
xor U15331 (N_15331,N_11021,N_10737);
xor U15332 (N_15332,N_12083,N_10105);
xor U15333 (N_15333,N_10812,N_11638);
or U15334 (N_15334,N_9781,N_11721);
nor U15335 (N_15335,N_10829,N_12032);
nand U15336 (N_15336,N_10099,N_9605);
or U15337 (N_15337,N_11884,N_9715);
and U15338 (N_15338,N_11251,N_10427);
nand U15339 (N_15339,N_10140,N_10582);
or U15340 (N_15340,N_10373,N_12150);
xor U15341 (N_15341,N_11139,N_9911);
or U15342 (N_15342,N_9891,N_11121);
nor U15343 (N_15343,N_12478,N_11181);
or U15344 (N_15344,N_11555,N_10288);
nor U15345 (N_15345,N_10041,N_10318);
nor U15346 (N_15346,N_10103,N_11506);
or U15347 (N_15347,N_10496,N_10227);
nor U15348 (N_15348,N_12153,N_10588);
xor U15349 (N_15349,N_10509,N_11530);
xnor U15350 (N_15350,N_12419,N_12270);
and U15351 (N_15351,N_12190,N_11531);
nand U15352 (N_15352,N_10847,N_10281);
xor U15353 (N_15353,N_10900,N_12068);
nand U15354 (N_15354,N_12245,N_10805);
and U15355 (N_15355,N_9958,N_11518);
nand U15356 (N_15356,N_10714,N_9429);
nor U15357 (N_15357,N_9397,N_9568);
nand U15358 (N_15358,N_10659,N_11630);
or U15359 (N_15359,N_11161,N_12020);
or U15360 (N_15360,N_9467,N_9884);
or U15361 (N_15361,N_10050,N_11745);
nand U15362 (N_15362,N_10283,N_9552);
xnor U15363 (N_15363,N_10935,N_10220);
xnor U15364 (N_15364,N_10854,N_9633);
nand U15365 (N_15365,N_9464,N_10014);
nor U15366 (N_15366,N_11834,N_12168);
nand U15367 (N_15367,N_10572,N_10364);
nor U15368 (N_15368,N_10607,N_12409);
or U15369 (N_15369,N_10949,N_10315);
or U15370 (N_15370,N_9956,N_11949);
nor U15371 (N_15371,N_9418,N_12319);
and U15372 (N_15372,N_11214,N_11522);
and U15373 (N_15373,N_10742,N_12170);
and U15374 (N_15374,N_10947,N_11432);
or U15375 (N_15375,N_9664,N_12073);
xor U15376 (N_15376,N_10986,N_10101);
and U15377 (N_15377,N_11767,N_10230);
nor U15378 (N_15378,N_12124,N_10867);
nand U15379 (N_15379,N_10279,N_9394);
and U15380 (N_15380,N_12297,N_10178);
nand U15381 (N_15381,N_10504,N_12082);
or U15382 (N_15382,N_9662,N_10718);
nor U15383 (N_15383,N_11694,N_10428);
nor U15384 (N_15384,N_11971,N_11267);
nor U15385 (N_15385,N_9504,N_10744);
and U15386 (N_15386,N_10612,N_10685);
nand U15387 (N_15387,N_10333,N_11596);
or U15388 (N_15388,N_11449,N_10850);
nor U15389 (N_15389,N_11462,N_11669);
or U15390 (N_15390,N_11093,N_12491);
or U15391 (N_15391,N_10012,N_10147);
or U15392 (N_15392,N_10941,N_10522);
nand U15393 (N_15393,N_11325,N_12069);
and U15394 (N_15394,N_10679,N_9574);
nand U15395 (N_15395,N_10570,N_9777);
and U15396 (N_15396,N_11460,N_11761);
nand U15397 (N_15397,N_10201,N_11715);
xor U15398 (N_15398,N_10670,N_12137);
or U15399 (N_15399,N_12041,N_11909);
and U15400 (N_15400,N_10637,N_10150);
nor U15401 (N_15401,N_11323,N_10944);
nand U15402 (N_15402,N_9584,N_11198);
xor U15403 (N_15403,N_9965,N_9817);
nor U15404 (N_15404,N_10732,N_12160);
nor U15405 (N_15405,N_11615,N_9787);
nor U15406 (N_15406,N_12315,N_9887);
nor U15407 (N_15407,N_9963,N_11581);
nand U15408 (N_15408,N_10040,N_10036);
nand U15409 (N_15409,N_10900,N_10191);
nand U15410 (N_15410,N_10945,N_9907);
nor U15411 (N_15411,N_10155,N_10901);
and U15412 (N_15412,N_9380,N_12292);
nand U15413 (N_15413,N_11656,N_10347);
xnor U15414 (N_15414,N_11185,N_10672);
xnor U15415 (N_15415,N_10621,N_12187);
or U15416 (N_15416,N_11157,N_11026);
and U15417 (N_15417,N_11275,N_10194);
xnor U15418 (N_15418,N_9718,N_11697);
nand U15419 (N_15419,N_10637,N_10752);
or U15420 (N_15420,N_10789,N_11608);
nand U15421 (N_15421,N_11648,N_9882);
nor U15422 (N_15422,N_9715,N_11265);
xor U15423 (N_15423,N_10819,N_11358);
or U15424 (N_15424,N_11383,N_9398);
nor U15425 (N_15425,N_9579,N_12247);
xor U15426 (N_15426,N_11739,N_11531);
xnor U15427 (N_15427,N_10958,N_11241);
xnor U15428 (N_15428,N_11879,N_12083);
or U15429 (N_15429,N_9502,N_11379);
nand U15430 (N_15430,N_9451,N_11496);
nor U15431 (N_15431,N_10431,N_10219);
xnor U15432 (N_15432,N_9433,N_12486);
or U15433 (N_15433,N_10589,N_10897);
and U15434 (N_15434,N_10658,N_11087);
nor U15435 (N_15435,N_11169,N_10894);
or U15436 (N_15436,N_11781,N_12406);
or U15437 (N_15437,N_12127,N_10163);
xor U15438 (N_15438,N_10395,N_11518);
nand U15439 (N_15439,N_10959,N_11323);
nand U15440 (N_15440,N_9497,N_12445);
xor U15441 (N_15441,N_10542,N_10886);
nand U15442 (N_15442,N_11301,N_11152);
nand U15443 (N_15443,N_10511,N_10013);
xnor U15444 (N_15444,N_11703,N_10992);
xnor U15445 (N_15445,N_10386,N_9692);
nor U15446 (N_15446,N_9664,N_9817);
nand U15447 (N_15447,N_10470,N_11813);
nand U15448 (N_15448,N_11326,N_10823);
xor U15449 (N_15449,N_11518,N_9971);
xnor U15450 (N_15450,N_9769,N_11364);
and U15451 (N_15451,N_11474,N_10945);
xor U15452 (N_15452,N_12311,N_10534);
nor U15453 (N_15453,N_12132,N_11102);
or U15454 (N_15454,N_12014,N_12297);
nor U15455 (N_15455,N_9798,N_10476);
nor U15456 (N_15456,N_9815,N_9689);
nand U15457 (N_15457,N_11341,N_10990);
or U15458 (N_15458,N_11370,N_10333);
or U15459 (N_15459,N_10619,N_10624);
and U15460 (N_15460,N_10067,N_9935);
nor U15461 (N_15461,N_9650,N_10851);
nor U15462 (N_15462,N_11512,N_11339);
xor U15463 (N_15463,N_10395,N_10236);
or U15464 (N_15464,N_9489,N_11049);
or U15465 (N_15465,N_10650,N_10543);
and U15466 (N_15466,N_11763,N_10531);
or U15467 (N_15467,N_11547,N_10682);
xnor U15468 (N_15468,N_10222,N_10794);
nand U15469 (N_15469,N_10521,N_9991);
or U15470 (N_15470,N_11429,N_11253);
xor U15471 (N_15471,N_12038,N_10796);
nor U15472 (N_15472,N_11015,N_9731);
or U15473 (N_15473,N_12209,N_11950);
and U15474 (N_15474,N_11116,N_10397);
or U15475 (N_15475,N_12121,N_10998);
nor U15476 (N_15476,N_12256,N_10315);
and U15477 (N_15477,N_10490,N_11492);
xnor U15478 (N_15478,N_12072,N_10788);
and U15479 (N_15479,N_11165,N_11254);
xor U15480 (N_15480,N_11256,N_10869);
nand U15481 (N_15481,N_12088,N_9755);
nor U15482 (N_15482,N_10343,N_9854);
nor U15483 (N_15483,N_10041,N_9992);
or U15484 (N_15484,N_10396,N_9633);
xnor U15485 (N_15485,N_9492,N_11298);
nand U15486 (N_15486,N_11241,N_10750);
xor U15487 (N_15487,N_9737,N_12286);
xnor U15488 (N_15488,N_10056,N_9867);
or U15489 (N_15489,N_11931,N_10035);
nor U15490 (N_15490,N_10760,N_10362);
nor U15491 (N_15491,N_12371,N_10761);
nor U15492 (N_15492,N_10809,N_10026);
or U15493 (N_15493,N_9553,N_10784);
xor U15494 (N_15494,N_10233,N_10912);
nor U15495 (N_15495,N_9721,N_11717);
xnor U15496 (N_15496,N_10981,N_11100);
or U15497 (N_15497,N_12096,N_12110);
nand U15498 (N_15498,N_10993,N_9499);
nand U15499 (N_15499,N_10189,N_11459);
nor U15500 (N_15500,N_11426,N_11842);
nor U15501 (N_15501,N_10974,N_11159);
or U15502 (N_15502,N_10909,N_9940);
or U15503 (N_15503,N_10121,N_9639);
or U15504 (N_15504,N_10394,N_12214);
and U15505 (N_15505,N_11316,N_10608);
nor U15506 (N_15506,N_10472,N_10925);
nor U15507 (N_15507,N_9598,N_10251);
or U15508 (N_15508,N_10506,N_9494);
and U15509 (N_15509,N_11917,N_11004);
xnor U15510 (N_15510,N_12288,N_10265);
or U15511 (N_15511,N_9552,N_11055);
nor U15512 (N_15512,N_11133,N_10988);
and U15513 (N_15513,N_12442,N_10352);
nor U15514 (N_15514,N_11669,N_11815);
xnor U15515 (N_15515,N_11684,N_10582);
nor U15516 (N_15516,N_10489,N_10593);
xnor U15517 (N_15517,N_12419,N_11645);
nor U15518 (N_15518,N_9637,N_11313);
and U15519 (N_15519,N_10009,N_10273);
nand U15520 (N_15520,N_12209,N_9944);
xor U15521 (N_15521,N_10926,N_10430);
nand U15522 (N_15522,N_10788,N_11460);
nor U15523 (N_15523,N_12048,N_10181);
xor U15524 (N_15524,N_10244,N_9621);
and U15525 (N_15525,N_11821,N_10360);
nand U15526 (N_15526,N_10054,N_9494);
xnor U15527 (N_15527,N_9591,N_9771);
or U15528 (N_15528,N_11025,N_12147);
nand U15529 (N_15529,N_12176,N_11054);
nand U15530 (N_15530,N_11291,N_11829);
nand U15531 (N_15531,N_12111,N_9525);
or U15532 (N_15532,N_9597,N_12414);
and U15533 (N_15533,N_10927,N_9580);
nand U15534 (N_15534,N_11561,N_9379);
and U15535 (N_15535,N_11621,N_11721);
nor U15536 (N_15536,N_11893,N_11435);
and U15537 (N_15537,N_12402,N_11300);
or U15538 (N_15538,N_11313,N_10308);
or U15539 (N_15539,N_9687,N_11084);
nand U15540 (N_15540,N_10773,N_11120);
xnor U15541 (N_15541,N_11133,N_12163);
or U15542 (N_15542,N_10524,N_10576);
nand U15543 (N_15543,N_10657,N_9924);
or U15544 (N_15544,N_12131,N_11578);
nor U15545 (N_15545,N_10729,N_12095);
nor U15546 (N_15546,N_10043,N_12043);
nor U15547 (N_15547,N_12237,N_11413);
nand U15548 (N_15548,N_9540,N_9395);
xor U15549 (N_15549,N_11385,N_12279);
xnor U15550 (N_15550,N_9718,N_12210);
xor U15551 (N_15551,N_10416,N_10461);
nor U15552 (N_15552,N_10672,N_10239);
or U15553 (N_15553,N_9626,N_11859);
or U15554 (N_15554,N_10958,N_9907);
nand U15555 (N_15555,N_10047,N_12073);
and U15556 (N_15556,N_9553,N_9789);
and U15557 (N_15557,N_10219,N_10969);
nand U15558 (N_15558,N_11203,N_9625);
xor U15559 (N_15559,N_9491,N_10547);
or U15560 (N_15560,N_9827,N_10969);
nand U15561 (N_15561,N_11971,N_12056);
or U15562 (N_15562,N_9931,N_11848);
nand U15563 (N_15563,N_11644,N_11294);
or U15564 (N_15564,N_10844,N_11099);
and U15565 (N_15565,N_10419,N_11328);
or U15566 (N_15566,N_10732,N_12164);
nand U15567 (N_15567,N_10034,N_11440);
and U15568 (N_15568,N_10309,N_11560);
xor U15569 (N_15569,N_10680,N_12402);
xnor U15570 (N_15570,N_11153,N_10536);
nor U15571 (N_15571,N_10810,N_11707);
xor U15572 (N_15572,N_11514,N_10180);
or U15573 (N_15573,N_9966,N_11386);
xor U15574 (N_15574,N_11940,N_11937);
nor U15575 (N_15575,N_9691,N_9557);
nor U15576 (N_15576,N_12004,N_10306);
nand U15577 (N_15577,N_11603,N_9620);
xnor U15578 (N_15578,N_10014,N_11439);
and U15579 (N_15579,N_9626,N_12494);
and U15580 (N_15580,N_11941,N_11148);
nand U15581 (N_15581,N_9429,N_12214);
nand U15582 (N_15582,N_9758,N_12170);
or U15583 (N_15583,N_12128,N_9879);
nor U15584 (N_15584,N_11237,N_11734);
nor U15585 (N_15585,N_9937,N_11797);
or U15586 (N_15586,N_11821,N_10194);
and U15587 (N_15587,N_11674,N_12165);
nor U15588 (N_15588,N_12238,N_12183);
and U15589 (N_15589,N_11886,N_10463);
or U15590 (N_15590,N_11748,N_9812);
or U15591 (N_15591,N_10429,N_10033);
xor U15592 (N_15592,N_11744,N_10969);
nand U15593 (N_15593,N_9383,N_11311);
and U15594 (N_15594,N_9407,N_10102);
and U15595 (N_15595,N_9573,N_12085);
and U15596 (N_15596,N_11529,N_12490);
and U15597 (N_15597,N_12325,N_10571);
or U15598 (N_15598,N_10156,N_10226);
and U15599 (N_15599,N_10210,N_10677);
xnor U15600 (N_15600,N_9451,N_11575);
xor U15601 (N_15601,N_10834,N_12436);
xor U15602 (N_15602,N_9568,N_9425);
nor U15603 (N_15603,N_11570,N_10745);
xor U15604 (N_15604,N_11648,N_10012);
or U15605 (N_15605,N_11999,N_12449);
and U15606 (N_15606,N_12327,N_10221);
nor U15607 (N_15607,N_11165,N_10444);
or U15608 (N_15608,N_12450,N_9497);
nand U15609 (N_15609,N_11254,N_12206);
or U15610 (N_15610,N_10642,N_9631);
or U15611 (N_15611,N_12081,N_12446);
and U15612 (N_15612,N_11522,N_10290);
and U15613 (N_15613,N_10809,N_11994);
nor U15614 (N_15614,N_11941,N_9827);
and U15615 (N_15615,N_9844,N_12298);
xnor U15616 (N_15616,N_10544,N_11739);
or U15617 (N_15617,N_10361,N_12292);
or U15618 (N_15618,N_9782,N_10786);
nand U15619 (N_15619,N_10279,N_11541);
or U15620 (N_15620,N_10699,N_11263);
xnor U15621 (N_15621,N_11499,N_10388);
xnor U15622 (N_15622,N_12202,N_11923);
or U15623 (N_15623,N_10556,N_9576);
xor U15624 (N_15624,N_11666,N_10628);
or U15625 (N_15625,N_12838,N_13238);
nor U15626 (N_15626,N_14100,N_14731);
nand U15627 (N_15627,N_15602,N_14290);
nand U15628 (N_15628,N_12965,N_13943);
or U15629 (N_15629,N_15229,N_12910);
nand U15630 (N_15630,N_13522,N_14691);
xnor U15631 (N_15631,N_14980,N_13135);
nand U15632 (N_15632,N_12699,N_14490);
or U15633 (N_15633,N_14115,N_14024);
nor U15634 (N_15634,N_14149,N_14217);
nor U15635 (N_15635,N_14665,N_13773);
and U15636 (N_15636,N_14930,N_12668);
or U15637 (N_15637,N_15512,N_14752);
xor U15638 (N_15638,N_15015,N_13167);
or U15639 (N_15639,N_13023,N_14406);
and U15640 (N_15640,N_15542,N_14921);
or U15641 (N_15641,N_13936,N_12878);
nand U15642 (N_15642,N_12616,N_12879);
and U15643 (N_15643,N_12964,N_15483);
nand U15644 (N_15644,N_14122,N_14689);
and U15645 (N_15645,N_14247,N_13810);
nand U15646 (N_15646,N_14883,N_14028);
and U15647 (N_15647,N_13470,N_12714);
and U15648 (N_15648,N_14979,N_13892);
or U15649 (N_15649,N_12969,N_12722);
xor U15650 (N_15650,N_13896,N_12899);
nand U15651 (N_15651,N_15258,N_13493);
or U15652 (N_15652,N_13545,N_12933);
xnor U15653 (N_15653,N_14938,N_13814);
nand U15654 (N_15654,N_13580,N_14204);
or U15655 (N_15655,N_13374,N_13663);
xnor U15656 (N_15656,N_12773,N_12537);
and U15657 (N_15657,N_14117,N_14165);
nor U15658 (N_15658,N_13624,N_15329);
xnor U15659 (N_15659,N_14700,N_15442);
and U15660 (N_15660,N_14532,N_14348);
nor U15661 (N_15661,N_14225,N_12974);
xnor U15662 (N_15662,N_15234,N_15008);
xor U15663 (N_15663,N_14120,N_13334);
or U15664 (N_15664,N_13932,N_13190);
or U15665 (N_15665,N_13213,N_14947);
nor U15666 (N_15666,N_13784,N_12562);
xor U15667 (N_15667,N_13536,N_12880);
nor U15668 (N_15668,N_15577,N_13022);
and U15669 (N_15669,N_13154,N_15197);
nand U15670 (N_15670,N_12634,N_13860);
and U15671 (N_15671,N_14517,N_14672);
nand U15672 (N_15672,N_12510,N_14419);
xor U15673 (N_15673,N_13954,N_14956);
and U15674 (N_15674,N_14832,N_13298);
nor U15675 (N_15675,N_14297,N_15279);
or U15676 (N_15676,N_14879,N_13286);
nor U15677 (N_15677,N_15511,N_12750);
and U15678 (N_15678,N_14656,N_14670);
nor U15679 (N_15679,N_13696,N_12882);
nand U15680 (N_15680,N_14260,N_14594);
nor U15681 (N_15681,N_14516,N_13911);
or U15682 (N_15682,N_12914,N_14345);
xnor U15683 (N_15683,N_14417,N_14040);
nor U15684 (N_15684,N_15464,N_14151);
or U15685 (N_15685,N_15290,N_14943);
nor U15686 (N_15686,N_13611,N_13109);
nand U15687 (N_15687,N_14513,N_14279);
and U15688 (N_15688,N_13137,N_13080);
xor U15689 (N_15689,N_15020,N_15477);
xnor U15690 (N_15690,N_14212,N_15334);
or U15691 (N_15691,N_14363,N_12854);
nand U15692 (N_15692,N_14944,N_15605);
and U15693 (N_15693,N_14164,N_13568);
nand U15694 (N_15694,N_15022,N_13273);
or U15695 (N_15695,N_14300,N_12960);
nand U15696 (N_15696,N_14551,N_15176);
xor U15697 (N_15697,N_12583,N_15308);
nor U15698 (N_15698,N_12558,N_14505);
nor U15699 (N_15699,N_12855,N_12520);
nor U15700 (N_15700,N_13788,N_12825);
and U15701 (N_15701,N_12777,N_12962);
xor U15702 (N_15702,N_14992,N_13234);
xnor U15703 (N_15703,N_14144,N_13822);
nand U15704 (N_15704,N_14008,N_15569);
xnor U15705 (N_15705,N_14892,N_13661);
nor U15706 (N_15706,N_15058,N_14064);
nor U15707 (N_15707,N_12966,N_15275);
and U15708 (N_15708,N_14186,N_15622);
or U15709 (N_15709,N_12612,N_14336);
nor U15710 (N_15710,N_14628,N_14463);
nor U15711 (N_15711,N_13224,N_14801);
xor U15712 (N_15712,N_12509,N_14588);
nor U15713 (N_15713,N_13774,N_13508);
xnor U15714 (N_15714,N_14367,N_15076);
and U15715 (N_15715,N_14231,N_14006);
xor U15716 (N_15716,N_15053,N_14312);
or U15717 (N_15717,N_14773,N_12840);
nor U15718 (N_15718,N_15405,N_13990);
or U15719 (N_15719,N_14677,N_13305);
or U15720 (N_15720,N_13703,N_13254);
nor U15721 (N_15721,N_12533,N_13680);
xor U15722 (N_15722,N_13420,N_12913);
xor U15723 (N_15723,N_14566,N_13079);
or U15724 (N_15724,N_15557,N_13887);
nor U15725 (N_15725,N_13863,N_15547);
or U15726 (N_15726,N_14882,N_13743);
nor U15727 (N_15727,N_12704,N_13592);
nor U15728 (N_15728,N_13581,N_14420);
nand U15729 (N_15729,N_14510,N_15374);
nor U15730 (N_15730,N_14473,N_15516);
and U15731 (N_15731,N_12522,N_15583);
nor U15732 (N_15732,N_12918,N_13162);
or U15733 (N_15733,N_13113,N_14994);
nand U15734 (N_15734,N_14386,N_13296);
nand U15735 (N_15735,N_12903,N_14527);
nor U15736 (N_15736,N_13692,N_13565);
nor U15737 (N_15737,N_15340,N_13124);
and U15738 (N_15738,N_13546,N_12700);
nand U15739 (N_15739,N_12919,N_12824);
nand U15740 (N_15740,N_13978,N_14894);
xor U15741 (N_15741,N_12666,N_15530);
and U15742 (N_15742,N_15142,N_13176);
and U15743 (N_15743,N_12861,N_14397);
and U15744 (N_15744,N_14612,N_13654);
nor U15745 (N_15745,N_14817,N_14910);
or U15746 (N_15746,N_12850,N_12967);
nand U15747 (N_15747,N_12954,N_14605);
nand U15748 (N_15748,N_13045,N_15227);
nor U15749 (N_15749,N_14499,N_13391);
nor U15750 (N_15750,N_15415,N_14307);
and U15751 (N_15751,N_14041,N_13052);
xor U15752 (N_15752,N_14922,N_13159);
nand U15753 (N_15753,N_13626,N_12846);
xnor U15754 (N_15754,N_13761,N_14423);
and U15755 (N_15755,N_14998,N_12888);
and U15756 (N_15756,N_13389,N_15387);
xnor U15757 (N_15757,N_14427,N_14716);
xnor U15758 (N_15758,N_13709,N_14553);
and U15759 (N_15759,N_14522,N_12772);
xor U15760 (N_15760,N_13153,N_13132);
nand U15761 (N_15761,N_13304,N_14826);
nor U15762 (N_15762,N_14990,N_13476);
nand U15763 (N_15763,N_12895,N_13034);
xnor U15764 (N_15764,N_13101,N_13477);
xor U15765 (N_15765,N_14767,N_15230);
or U15766 (N_15766,N_14074,N_13384);
nor U15767 (N_15767,N_15225,N_15216);
or U15768 (N_15768,N_15170,N_14641);
or U15769 (N_15769,N_13363,N_13938);
nor U15770 (N_15770,N_13123,N_14368);
xor U15771 (N_15771,N_14845,N_12638);
or U15772 (N_15772,N_14294,N_14190);
nor U15773 (N_15773,N_12743,N_13729);
nor U15774 (N_15774,N_15438,N_12552);
nand U15775 (N_15775,N_14021,N_13591);
nor U15776 (N_15776,N_14802,N_12872);
xor U15777 (N_15777,N_13248,N_13647);
nor U15778 (N_15778,N_12950,N_13292);
nor U15779 (N_15779,N_13940,N_14133);
nor U15780 (N_15780,N_15260,N_15404);
nor U15781 (N_15781,N_14026,N_15322);
nand U15782 (N_15782,N_13882,N_13408);
xor U15783 (N_15783,N_13745,N_14985);
and U15784 (N_15784,N_15193,N_13695);
nor U15785 (N_15785,N_13084,N_12911);
nand U15786 (N_15786,N_14210,N_15503);
or U15787 (N_15787,N_15039,N_13199);
nor U15788 (N_15788,N_14687,N_13561);
or U15789 (N_15789,N_13942,N_14774);
nand U15790 (N_15790,N_13429,N_12740);
and U15791 (N_15791,N_13619,N_14476);
xor U15792 (N_15792,N_15526,N_13212);
nand U15793 (N_15793,N_15292,N_12993);
xor U15794 (N_15794,N_14342,N_13371);
nand U15795 (N_15795,N_15467,N_14441);
and U15796 (N_15796,N_15502,N_14760);
and U15797 (N_15797,N_13988,N_14431);
or U15798 (N_15798,N_12547,N_13783);
and U15799 (N_15799,N_14808,N_15388);
or U15800 (N_15800,N_14014,N_15561);
nor U15801 (N_15801,N_12805,N_13419);
xor U15802 (N_15802,N_14283,N_14614);
xor U15803 (N_15803,N_14685,N_14791);
and U15804 (N_15804,N_14373,N_14253);
xnor U15805 (N_15805,N_13404,N_14137);
nand U15806 (N_15806,N_14055,N_13240);
nand U15807 (N_15807,N_15504,N_13732);
xnor U15808 (N_15808,N_14452,N_13142);
or U15809 (N_15809,N_13461,N_13157);
or U15810 (N_15810,N_14207,N_12618);
nor U15811 (N_15811,N_12756,N_14914);
or U15812 (N_15812,N_14303,N_15499);
nor U15813 (N_15813,N_14743,N_15124);
nand U15814 (N_15814,N_12736,N_12717);
nor U15815 (N_15815,N_14177,N_13505);
and U15816 (N_15816,N_13852,N_14183);
or U15817 (N_15817,N_13338,N_15281);
or U15818 (N_15818,N_14061,N_12671);
xnor U15819 (N_15819,N_12904,N_15167);
xnor U15820 (N_15820,N_14255,N_12694);
xor U15821 (N_15821,N_12594,N_14491);
or U15822 (N_15822,N_13350,N_12534);
and U15823 (N_15823,N_13434,N_12749);
or U15824 (N_15824,N_15276,N_13438);
nor U15825 (N_15825,N_14907,N_13141);
nor U15826 (N_15826,N_13617,N_15121);
or U15827 (N_15827,N_13782,N_13638);
nor U15828 (N_15828,N_14382,N_13598);
or U15829 (N_15829,N_13950,N_13516);
xnor U15830 (N_15830,N_14310,N_13051);
nand U15831 (N_15831,N_15253,N_13143);
or U15832 (N_15832,N_13453,N_13726);
xor U15833 (N_15833,N_14284,N_12818);
nor U15834 (N_15834,N_12713,N_14898);
xnor U15835 (N_15835,N_13679,N_15574);
nand U15836 (N_15836,N_15109,N_12663);
and U15837 (N_15837,N_14509,N_13741);
nand U15838 (N_15838,N_13651,N_13466);
nor U15839 (N_15839,N_12997,N_12893);
or U15840 (N_15840,N_14782,N_14748);
and U15841 (N_15841,N_15386,N_12782);
or U15842 (N_15842,N_15420,N_15435);
nor U15843 (N_15843,N_15609,N_13605);
xor U15844 (N_15844,N_15558,N_14459);
xnor U15845 (N_15845,N_14970,N_12864);
nor U15846 (N_15846,N_14957,N_13055);
xnor U15847 (N_15847,N_13287,N_15389);
xnor U15848 (N_15848,N_15168,N_14200);
or U15849 (N_15849,N_13697,N_15338);
or U15850 (N_15850,N_14319,N_14197);
or U15851 (N_15851,N_13720,N_13173);
or U15852 (N_15852,N_12747,N_14591);
nor U15853 (N_15853,N_15231,N_14624);
nor U15854 (N_15854,N_14796,N_13980);
nor U15855 (N_15855,N_15597,N_14188);
xnor U15856 (N_15856,N_12984,N_13976);
and U15857 (N_15857,N_13275,N_15521);
nand U15858 (N_15858,N_13897,N_12513);
nand U15859 (N_15859,N_14704,N_15576);
nor U15860 (N_15860,N_13129,N_14178);
xnor U15861 (N_15861,N_14753,N_14318);
xnor U15862 (N_15862,N_14585,N_15088);
nor U15863 (N_15863,N_15552,N_13362);
xor U15864 (N_15864,N_14453,N_12801);
and U15865 (N_15865,N_15102,N_12688);
and U15866 (N_15866,N_14698,N_12842);
xnor U15867 (N_15867,N_12902,N_13417);
or U15868 (N_15868,N_15246,N_15449);
nor U15869 (N_15869,N_12590,N_15037);
nand U15870 (N_15870,N_15339,N_12991);
xnor U15871 (N_15871,N_12819,N_14366);
xnor U15872 (N_15872,N_14781,N_15257);
nand U15873 (N_15873,N_12517,N_14145);
nor U15874 (N_15874,N_15592,N_12557);
nor U15875 (N_15875,N_15301,N_12889);
and U15876 (N_15876,N_12602,N_13138);
xor U15877 (N_15877,N_15612,N_13884);
xnor U15878 (N_15878,N_15402,N_14350);
nand U15879 (N_15879,N_13594,N_14906);
xnor U15880 (N_15880,N_15151,N_14933);
xnor U15881 (N_15881,N_15615,N_14592);
nand U15882 (N_15882,N_14409,N_14011);
and U15883 (N_15883,N_13635,N_14820);
xor U15884 (N_15884,N_14926,N_15127);
and U15885 (N_15885,N_14126,N_15436);
nand U15886 (N_15886,N_13603,N_13103);
xor U15887 (N_15887,N_13541,N_13291);
or U15888 (N_15888,N_14548,N_14436);
nand U15889 (N_15889,N_14602,N_13195);
nor U15890 (N_15890,N_13295,N_13755);
nor U15891 (N_15891,N_13785,N_15345);
and U15892 (N_15892,N_14264,N_13431);
nand U15893 (N_15893,N_15224,N_13722);
and U15894 (N_15894,N_15537,N_14084);
and U15895 (N_15895,N_15610,N_14972);
or U15896 (N_15896,N_14315,N_15122);
nand U15897 (N_15897,N_14642,N_12501);
nor U15898 (N_15898,N_15366,N_14187);
nor U15899 (N_15899,N_13798,N_15298);
nand U15900 (N_15900,N_13922,N_13615);
nand U15901 (N_15901,N_13805,N_14056);
nor U15902 (N_15902,N_12812,N_12833);
nor U15903 (N_15903,N_15238,N_13705);
and U15904 (N_15904,N_12909,N_14552);
nand U15905 (N_15905,N_14201,N_12523);
or U15906 (N_15906,N_13192,N_13490);
and U15907 (N_15907,N_14042,N_15129);
or U15908 (N_15908,N_14757,N_15103);
or U15909 (N_15909,N_13025,N_15481);
xor U15910 (N_15910,N_13027,N_13584);
xor U15911 (N_15911,N_15300,N_14269);
and U15912 (N_15912,N_13993,N_14376);
or U15913 (N_15913,N_13119,N_13105);
or U15914 (N_15914,N_12932,N_13083);
xnor U15915 (N_15915,N_12761,N_14384);
or U15916 (N_15916,N_13958,N_13155);
and U15917 (N_15917,N_12892,N_14309);
nand U15918 (N_15918,N_14439,N_13693);
xor U15919 (N_15919,N_12944,N_12857);
xor U15920 (N_15920,N_13198,N_13320);
or U15921 (N_15921,N_15429,N_13847);
nor U15922 (N_15922,N_12669,N_13258);
nand U15923 (N_15923,N_15051,N_13222);
nand U15924 (N_15924,N_13998,N_15307);
xor U15925 (N_15925,N_15443,N_14523);
xnor U15926 (N_15926,N_15492,N_12640);
nor U15927 (N_15927,N_15033,N_13539);
nand U15928 (N_15928,N_12647,N_13011);
or U15929 (N_15929,N_13145,N_15045);
and U15930 (N_15930,N_12516,N_15446);
nor U15931 (N_15931,N_12572,N_12614);
and U15932 (N_15932,N_12844,N_13855);
and U15933 (N_15933,N_13944,N_15517);
xor U15934 (N_15934,N_13432,N_15140);
and U15935 (N_15935,N_13948,N_14037);
or U15936 (N_15936,N_13514,N_13507);
nor U15937 (N_15937,N_13524,N_12692);
nor U15938 (N_15938,N_14541,N_14596);
nand U15939 (N_15939,N_14285,N_15038);
xnor U15940 (N_15940,N_15553,N_13657);
nand U15941 (N_15941,N_13989,N_15028);
nand U15942 (N_15942,N_14736,N_13040);
and U15943 (N_15943,N_15453,N_13242);
nor U15944 (N_15944,N_14728,N_13671);
nor U15945 (N_15945,N_13383,N_14827);
and U15946 (N_15946,N_13941,N_12752);
and U15947 (N_15947,N_14220,N_14720);
and U15948 (N_15948,N_13961,N_15589);
nand U15949 (N_15949,N_14680,N_12582);
or U15950 (N_15950,N_15191,N_14920);
nand U15951 (N_15951,N_14132,N_12847);
nand U15952 (N_15952,N_13409,N_13844);
or U15953 (N_15953,N_15575,N_12983);
nand U15954 (N_15954,N_14697,N_14901);
nor U15955 (N_15955,N_13228,N_12672);
xor U15956 (N_15956,N_14400,N_13444);
nor U15957 (N_15957,N_15562,N_13381);
and U15958 (N_15958,N_13837,N_13136);
nor U15959 (N_15959,N_13426,N_14338);
nor U15960 (N_15960,N_13365,N_14891);
nand U15961 (N_15961,N_12813,N_12644);
nand U15962 (N_15962,N_15336,N_13920);
and U15963 (N_15963,N_14182,N_13796);
xnor U15964 (N_15964,N_12765,N_14829);
nor U15965 (N_15965,N_12649,N_14945);
or U15966 (N_15966,N_12768,N_15536);
nor U15967 (N_15967,N_14525,N_13956);
nor U15968 (N_15968,N_12780,N_15331);
nand U15969 (N_15969,N_13098,N_15243);
or U15970 (N_15970,N_14424,N_14657);
xor U15971 (N_15971,N_14324,N_12724);
or U15972 (N_15972,N_12887,N_14948);
and U15973 (N_15973,N_15207,N_13612);
and U15974 (N_15974,N_13537,N_12566);
or U15975 (N_15975,N_15035,N_14568);
nand U15976 (N_15976,N_12698,N_14590);
and U15977 (N_15977,N_12968,N_13010);
xnor U15978 (N_15978,N_14460,N_15280);
xnor U15979 (N_15979,N_13166,N_13962);
or U15980 (N_15980,N_15498,N_14719);
and U15981 (N_15981,N_13193,N_14851);
or U15982 (N_15982,N_13202,N_13152);
nand U15983 (N_15983,N_12697,N_14821);
nand U15984 (N_15984,N_14834,N_13757);
xnor U15985 (N_15985,N_15508,N_14763);
and U15986 (N_15986,N_15115,N_14196);
nor U15987 (N_15987,N_12972,N_15391);
or U15988 (N_15988,N_14241,N_14029);
nand U15989 (N_15989,N_14222,N_15206);
nor U15990 (N_15990,N_13309,N_15242);
and U15991 (N_15991,N_14722,N_15304);
or U15992 (N_15992,N_15482,N_13313);
nand U15993 (N_15993,N_13555,N_14542);
and U15994 (N_15994,N_14616,N_12925);
nand U15995 (N_15995,N_14414,N_15384);
and U15996 (N_15996,N_13842,N_13549);
nor U15997 (N_15997,N_13256,N_15540);
nand U15998 (N_15998,N_14941,N_14637);
xor U15999 (N_15999,N_12580,N_15613);
xor U16000 (N_16000,N_13096,N_13596);
xnor U16001 (N_16001,N_13778,N_14579);
or U16002 (N_16002,N_15024,N_13436);
nor U16003 (N_16003,N_14580,N_14261);
or U16004 (N_16004,N_13411,N_15198);
and U16005 (N_16005,N_13092,N_13239);
xnor U16006 (N_16006,N_13845,N_12657);
or U16007 (N_16007,N_13877,N_14160);
xor U16008 (N_16008,N_15289,N_15172);
and U16009 (N_16009,N_12860,N_13464);
nand U16010 (N_16010,N_14908,N_12735);
nor U16011 (N_16011,N_14359,N_14504);
xor U16012 (N_16012,N_14876,N_12524);
nor U16013 (N_16013,N_14009,N_14089);
and U16014 (N_16014,N_13415,N_14226);
xnor U16015 (N_16015,N_14238,N_14482);
or U16016 (N_16016,N_14887,N_12998);
nor U16017 (N_16017,N_13351,N_14135);
nor U16018 (N_16018,N_12908,N_15259);
nor U16019 (N_16019,N_14379,N_14618);
or U16020 (N_16020,N_13353,N_13232);
or U16021 (N_16021,N_13104,N_12792);
nand U16022 (N_16022,N_15185,N_12605);
xor U16023 (N_16023,N_13414,N_14198);
xnor U16024 (N_16024,N_13968,N_15011);
and U16025 (N_16025,N_15541,N_14508);
and U16026 (N_16026,N_14375,N_14022);
xor U16027 (N_16027,N_13893,N_15531);
nor U16028 (N_16028,N_13634,N_15457);
nand U16029 (N_16029,N_15594,N_14583);
nor U16030 (N_16030,N_15459,N_12883);
and U16031 (N_16031,N_15302,N_14136);
xor U16032 (N_16032,N_14265,N_13346);
nor U16033 (N_16033,N_13945,N_12858);
and U16034 (N_16034,N_12507,N_15196);
nor U16035 (N_16035,N_15312,N_13853);
xor U16036 (N_16036,N_15554,N_15488);
nor U16037 (N_16037,N_13174,N_13871);
and U16038 (N_16038,N_13526,N_14357);
or U16039 (N_16039,N_15458,N_14570);
xor U16040 (N_16040,N_14962,N_15044);
nor U16041 (N_16041,N_12529,N_12601);
nand U16042 (N_16042,N_12521,N_14125);
and U16043 (N_16043,N_14848,N_15461);
xnor U16044 (N_16044,N_14617,N_15082);
nand U16045 (N_16045,N_13704,N_14789);
xor U16046 (N_16046,N_14867,N_14988);
nand U16047 (N_16047,N_14754,N_15532);
nor U16048 (N_16048,N_12905,N_15318);
nor U16049 (N_16049,N_15327,N_15523);
xnor U16050 (N_16050,N_12624,N_13220);
and U16051 (N_16051,N_14604,N_14804);
or U16052 (N_16052,N_14387,N_12835);
and U16053 (N_16053,N_14337,N_14783);
nand U16054 (N_16054,N_12691,N_15556);
xnor U16055 (N_16055,N_14272,N_13700);
nand U16056 (N_16056,N_15041,N_14912);
nand U16057 (N_16057,N_13099,N_13227);
nand U16058 (N_16058,N_13768,N_13898);
or U16059 (N_16059,N_14521,N_14790);
and U16060 (N_16060,N_14835,N_13107);
xnor U16061 (N_16061,N_14816,N_15217);
nor U16062 (N_16062,N_15179,N_12870);
and U16063 (N_16063,N_15248,N_15272);
or U16064 (N_16064,N_15424,N_15199);
nand U16065 (N_16065,N_13312,N_14786);
and U16066 (N_16066,N_15305,N_12575);
xnor U16067 (N_16067,N_13209,N_13604);
and U16068 (N_16068,N_14072,N_14809);
nor U16069 (N_16069,N_12979,N_13369);
or U16070 (N_16070,N_15428,N_14667);
nand U16071 (N_16071,N_13714,N_14440);
and U16072 (N_16072,N_13759,N_15125);
and U16073 (N_16073,N_13525,N_15614);
xor U16074 (N_16074,N_14062,N_13347);
or U16075 (N_16075,N_14445,N_14299);
or U16076 (N_16076,N_15204,N_15286);
xor U16077 (N_16077,N_13779,N_13380);
xnor U16078 (N_16078,N_14960,N_13412);
xnor U16079 (N_16079,N_12631,N_13225);
nor U16080 (N_16080,N_13684,N_15515);
xnor U16081 (N_16081,N_14167,N_13762);
xnor U16082 (N_16082,N_14039,N_13327);
xnor U16083 (N_16083,N_15178,N_13053);
nand U16084 (N_16084,N_12674,N_14044);
and U16085 (N_16085,N_14323,N_13252);
xor U16086 (N_16086,N_13026,N_14799);
and U16087 (N_16087,N_12753,N_13170);
xor U16088 (N_16088,N_12748,N_13515);
xnor U16089 (N_16089,N_13054,N_13971);
nand U16090 (N_16090,N_13205,N_15138);
and U16091 (N_16091,N_15171,N_13725);
or U16092 (N_16092,N_12865,N_14215);
and U16093 (N_16093,N_15518,N_13959);
nor U16094 (N_16094,N_12937,N_15578);
nand U16095 (N_16095,N_14154,N_12951);
xor U16096 (N_16096,N_12896,N_13314);
nand U16097 (N_16097,N_14717,N_14865);
xnor U16098 (N_16098,N_14636,N_13068);
and U16099 (N_16099,N_15529,N_13396);
xor U16100 (N_16100,N_15346,N_12931);
nor U16101 (N_16101,N_13475,N_14462);
nand U16102 (N_16102,N_13609,N_12900);
and U16103 (N_16103,N_15432,N_14124);
nand U16104 (N_16104,N_12938,N_13278);
nand U16105 (N_16105,N_12538,N_14356);
and U16106 (N_16106,N_14733,N_14905);
nand U16107 (N_16107,N_12577,N_14601);
nand U16108 (N_16108,N_13879,N_15007);
xnor U16109 (N_16109,N_14096,N_14537);
and U16110 (N_16110,N_14959,N_13229);
nor U16111 (N_16111,N_13572,N_14239);
xnor U16112 (N_16112,N_13169,N_14295);
xnor U16113 (N_16113,N_13751,N_12586);
or U16114 (N_16114,N_14402,N_12681);
and U16115 (N_16115,N_13593,N_13102);
nand U16116 (N_16116,N_15430,N_12550);
nor U16117 (N_16117,N_14507,N_14986);
or U16118 (N_16118,N_15116,N_14951);
nor U16119 (N_16119,N_12626,N_13498);
xor U16120 (N_16120,N_15315,N_12930);
nor U16121 (N_16121,N_15239,N_12915);
nor U16122 (N_16122,N_14437,N_13035);
nand U16123 (N_16123,N_13835,N_12957);
and U16124 (N_16124,N_15616,N_14169);
or U16125 (N_16125,N_12936,N_13557);
xnor U16126 (N_16126,N_12721,N_12662);
and U16127 (N_16127,N_14180,N_12596);
nor U16128 (N_16128,N_12771,N_13403);
and U16129 (N_16129,N_13405,N_13446);
and U16130 (N_16130,N_13738,N_14900);
and U16131 (N_16131,N_14846,N_12973);
or U16132 (N_16132,N_15455,N_13358);
nor U16133 (N_16133,N_13857,N_14455);
and U16134 (N_16134,N_12994,N_14586);
and U16135 (N_16135,N_14143,N_14091);
nor U16136 (N_16136,N_13008,N_13342);
xnor U16137 (N_16137,N_12738,N_15325);
and U16138 (N_16138,N_14610,N_13284);
and U16139 (N_16139,N_13550,N_15373);
nor U16140 (N_16140,N_13724,N_15363);
nor U16141 (N_16141,N_15066,N_14870);
and U16142 (N_16142,N_12784,N_14621);
nand U16143 (N_16143,N_12619,N_12708);
or U16144 (N_16144,N_13813,N_15228);
or U16145 (N_16145,N_15087,N_13185);
or U16146 (N_16146,N_15359,N_15150);
nand U16147 (N_16147,N_13375,N_12703);
nor U16148 (N_16148,N_15072,N_14822);
xor U16149 (N_16149,N_13646,N_13535);
xor U16150 (N_16150,N_15156,N_14221);
nor U16151 (N_16151,N_13901,N_13039);
and U16152 (N_16152,N_14405,N_14328);
nand U16153 (N_16153,N_12544,N_13236);
and U16154 (N_16154,N_15548,N_14007);
nor U16155 (N_16155,N_14082,N_13607);
and U16156 (N_16156,N_15251,N_15016);
nor U16157 (N_16157,N_12808,N_13370);
nor U16158 (N_16158,N_15570,N_15032);
or U16159 (N_16159,N_13015,N_12928);
or U16160 (N_16160,N_13097,N_14129);
or U16161 (N_16161,N_12953,N_15287);
nor U16162 (N_16162,N_13792,N_14545);
nor U16163 (N_16163,N_14780,N_13033);
xnor U16164 (N_16164,N_15113,N_15264);
and U16165 (N_16165,N_14113,N_14744);
nor U16166 (N_16166,N_13937,N_15568);
or U16167 (N_16167,N_13175,N_12633);
nand U16168 (N_16168,N_13050,N_15463);
nand U16169 (N_16169,N_12775,N_13172);
nand U16170 (N_16170,N_13064,N_14426);
xor U16171 (N_16171,N_15462,N_14712);
nand U16172 (N_16172,N_14561,N_14795);
and U16173 (N_16173,N_14885,N_15046);
xor U16174 (N_16174,N_13538,N_13471);
and U16175 (N_16175,N_12757,N_13093);
xor U16176 (N_16176,N_12881,N_13326);
or U16177 (N_16177,N_13566,N_13487);
nor U16178 (N_16178,N_14755,N_14528);
xor U16179 (N_16179,N_15510,N_14889);
and U16180 (N_16180,N_12710,N_12584);
nand U16181 (N_16181,N_14107,N_13427);
nor U16182 (N_16182,N_14498,N_13613);
or U16183 (N_16183,N_12670,N_13583);
and U16184 (N_16184,N_13637,N_14584);
nand U16185 (N_16185,N_13349,N_15050);
or U16186 (N_16186,N_13544,N_12642);
and U16187 (N_16187,N_13691,N_13623);
nor U16188 (N_16188,N_13717,N_15095);
xor U16189 (N_16189,N_13300,N_15064);
xor U16190 (N_16190,N_15273,N_15468);
nor U16191 (N_16191,N_13484,N_14195);
xnor U16192 (N_16192,N_13865,N_13977);
xnor U16193 (N_16193,N_14997,N_13401);
xor U16194 (N_16194,N_14475,N_13648);
or U16195 (N_16195,N_15250,N_13189);
nor U16196 (N_16196,N_12766,N_12981);
or U16197 (N_16197,N_13460,N_15081);
nand U16198 (N_16198,N_15379,N_13642);
xor U16199 (N_16199,N_15268,N_14157);
nand U16200 (N_16200,N_12573,N_14692);
xnor U16201 (N_16201,N_14916,N_14214);
or U16202 (N_16202,N_13085,N_13548);
nand U16203 (N_16203,N_14886,N_14138);
nand U16204 (N_16204,N_12891,N_15559);
and U16205 (N_16205,N_15369,N_14571);
and U16206 (N_16206,N_15586,N_13823);
nor U16207 (N_16207,N_12656,N_13125);
nand U16208 (N_16208,N_13249,N_13269);
and U16209 (N_16209,N_13708,N_12762);
nand U16210 (N_16210,N_13710,N_14114);
or U16211 (N_16211,N_13824,N_14660);
and U16212 (N_16212,N_15147,N_14560);
or U16213 (N_16213,N_13688,N_12725);
xnor U16214 (N_16214,N_14751,N_13231);
xnor U16215 (N_16215,N_14340,N_15539);
and U16216 (N_16216,N_14965,N_13206);
or U16217 (N_16217,N_15148,N_13909);
and U16218 (N_16218,N_13066,N_14654);
nand U16219 (N_16219,N_13770,N_15527);
nand U16220 (N_16220,N_14470,N_13818);
xnor U16221 (N_16221,N_14577,N_14448);
or U16222 (N_16222,N_13983,N_14381);
and U16223 (N_16223,N_12845,N_13216);
xor U16224 (N_16224,N_13888,N_12600);
nor U16225 (N_16225,N_14083,N_12591);
or U16226 (N_16226,N_13277,N_12543);
nand U16227 (N_16227,N_12728,N_15358);
and U16228 (N_16228,N_13267,N_15452);
and U16229 (N_16229,N_12648,N_13502);
xnor U16230 (N_16230,N_14018,N_13450);
nor U16231 (N_16231,N_14171,N_12791);
nand U16232 (N_16232,N_12961,N_12916);
nor U16233 (N_16233,N_15326,N_15343);
xnor U16234 (N_16234,N_14842,N_15143);
xnor U16235 (N_16235,N_15608,N_13850);
and U16236 (N_16236,N_13171,N_14394);
nor U16237 (N_16237,N_14308,N_13921);
or U16238 (N_16238,N_12853,N_14245);
and U16239 (N_16239,N_15174,N_14057);
or U16240 (N_16240,N_13018,N_15068);
and U16241 (N_16241,N_13707,N_12958);
nand U16242 (N_16242,N_14727,N_15310);
xor U16243 (N_16243,N_13780,N_14488);
xor U16244 (N_16244,N_14049,N_13866);
or U16245 (N_16245,N_13440,N_13194);
nand U16246 (N_16246,N_14678,N_13794);
nand U16247 (N_16247,N_12675,N_14016);
xnor U16248 (N_16248,N_14703,N_13633);
nor U16249 (N_16249,N_14502,N_14288);
nor U16250 (N_16250,N_14973,N_13931);
nand U16251 (N_16251,N_14838,N_13244);
or U16252 (N_16252,N_15454,N_12821);
and U16253 (N_16253,N_12707,N_14468);
or U16254 (N_16254,N_14099,N_14877);
and U16255 (N_16255,N_12632,N_12588);
xnor U16256 (N_16256,N_13081,N_13147);
xnor U16257 (N_16257,N_13433,N_12837);
nor U16258 (N_16258,N_14408,N_13203);
nor U16259 (N_16259,N_13279,N_14742);
xor U16260 (N_16260,N_13260,N_14811);
and U16261 (N_16261,N_15077,N_13595);
and U16262 (N_16262,N_15263,N_13658);
and U16263 (N_16263,N_14306,N_14098);
and U16264 (N_16264,N_15434,N_15110);
and U16265 (N_16265,N_15414,N_14749);
or U16266 (N_16266,N_13789,N_12680);
nand U16267 (N_16267,N_13563,N_13582);
xor U16268 (N_16268,N_15347,N_15490);
nand U16269 (N_16269,N_13333,N_15019);
nor U16270 (N_16270,N_14480,N_13044);
xnor U16271 (N_16271,N_14534,N_15117);
xor U16272 (N_16272,N_12554,N_15190);
or U16273 (N_16273,N_14179,N_12830);
nor U16274 (N_16274,N_13873,N_14170);
nand U16275 (N_16275,N_15514,N_12530);
and U16276 (N_16276,N_13131,N_12797);
nand U16277 (N_16277,N_12923,N_14412);
or U16278 (N_16278,N_15126,N_14981);
nor U16279 (N_16279,N_14159,N_13042);
and U16280 (N_16280,N_14158,N_13458);
nor U16281 (N_16281,N_14554,N_14068);
and U16282 (N_16282,N_14707,N_14747);
or U16283 (N_16283,N_14766,N_15057);
xor U16284 (N_16284,N_14902,N_14569);
nand U16285 (N_16285,N_14954,N_13418);
xor U16286 (N_16286,N_15328,N_15383);
nand U16287 (N_16287,N_12701,N_12571);
nor U16288 (N_16288,N_12511,N_14163);
nor U16289 (N_16289,N_15152,N_15118);
and U16290 (N_16290,N_14034,N_14166);
nand U16291 (N_16291,N_13685,N_14139);
xnor U16292 (N_16292,N_13151,N_13430);
xnor U16293 (N_16293,N_14193,N_15031);
or U16294 (N_16294,N_15071,N_13058);
and U16295 (N_16295,N_14395,N_14219);
nor U16296 (N_16296,N_13766,N_15299);
xor U16297 (N_16297,N_15219,N_14369);
and U16298 (N_16298,N_14088,N_13919);
or U16299 (N_16299,N_13821,N_13924);
and U16300 (N_16300,N_15293,N_13812);
or U16301 (N_16301,N_13144,N_15220);
nor U16302 (N_16302,N_15399,N_14705);
nand U16303 (N_16303,N_12679,N_15069);
or U16304 (N_16304,N_15445,N_12852);
nand U16305 (N_16305,N_14257,N_13880);
and U16306 (N_16306,N_14688,N_14273);
xor U16307 (N_16307,N_14365,N_13673);
and U16308 (N_16308,N_14244,N_14729);
and U16309 (N_16309,N_13062,N_15247);
nand U16310 (N_16310,N_12732,N_14547);
xnor U16311 (N_16311,N_14830,N_14076);
or U16312 (N_16312,N_14803,N_12690);
nor U16313 (N_16313,N_13521,N_13979);
or U16314 (N_16314,N_15226,N_14519);
nand U16315 (N_16315,N_14168,N_12659);
or U16316 (N_16316,N_13421,N_13527);
xor U16317 (N_16317,N_14772,N_13974);
nand U16318 (N_16318,N_15098,N_15471);
and U16319 (N_16319,N_15545,N_14355);
or U16320 (N_16320,N_12621,N_14370);
nand U16321 (N_16321,N_14694,N_15397);
nor U16322 (N_16322,N_15040,N_14105);
and U16323 (N_16323,N_13764,N_14485);
nor U16324 (N_16324,N_14927,N_14478);
nand U16325 (N_16325,N_12832,N_13311);
xor U16326 (N_16326,N_15385,N_14185);
xor U16327 (N_16327,N_14002,N_12744);
and U16328 (N_16328,N_13639,N_14343);
xnor U16329 (N_16329,N_13997,N_14233);
or U16330 (N_16330,N_13072,N_13985);
and U16331 (N_16331,N_15200,N_12542);
and U16332 (N_16332,N_13758,N_12992);
nand U16333 (N_16333,N_13043,N_12924);
or U16334 (N_16334,N_14422,N_14818);
xnor U16335 (N_16335,N_13870,N_14352);
nand U16336 (N_16336,N_14659,N_14112);
and U16337 (N_16337,N_14155,N_12935);
xor U16338 (N_16338,N_13463,N_14477);
or U16339 (N_16339,N_15215,N_14676);
xnor U16340 (N_16340,N_15593,N_12764);
or U16341 (N_16341,N_15381,N_14347);
xnor U16342 (N_16342,N_12652,N_12603);
nor U16343 (N_16343,N_15018,N_14924);
xor U16344 (N_16344,N_15354,N_13868);
nand U16345 (N_16345,N_13881,N_14715);
nor U16346 (N_16346,N_15145,N_14329);
or U16347 (N_16347,N_13439,N_14953);
and U16348 (N_16348,N_12898,N_15321);
or U16349 (N_16349,N_13664,N_13361);
or U16350 (N_16350,N_13059,N_12767);
and U16351 (N_16351,N_13235,N_13087);
nand U16352 (N_16352,N_12686,N_13553);
or U16353 (N_16353,N_13219,N_14732);
nand U16354 (N_16354,N_14010,N_14649);
or U16355 (N_16355,N_13982,N_15323);
xor U16356 (N_16356,N_13200,N_14249);
nand U16357 (N_16357,N_13090,N_14223);
nor U16358 (N_16358,N_15564,N_13395);
xnor U16359 (N_16359,N_14466,N_13073);
nand U16360 (N_16360,N_13492,N_14013);
xor U16361 (N_16361,N_14110,N_14538);
or U16362 (N_16362,N_14630,N_12592);
nor U16363 (N_16363,N_13221,N_15036);
and U16364 (N_16364,N_14880,N_15094);
nand U16365 (N_16365,N_13112,N_14267);
or U16366 (N_16366,N_14919,N_15450);
nor U16367 (N_16367,N_14853,N_14101);
or U16368 (N_16368,N_15390,N_14486);
nand U16369 (N_16369,N_15367,N_14067);
or U16370 (N_16370,N_13503,N_13100);
or U16371 (N_16371,N_14798,N_15427);
xor U16372 (N_16372,N_12715,N_13727);
xnor U16373 (N_16373,N_14492,N_13406);
xnor U16374 (N_16374,N_13315,N_13832);
and U16375 (N_16375,N_15086,N_13655);
nor U16376 (N_16376,N_12587,N_13070);
nor U16377 (N_16377,N_14974,N_14847);
or U16378 (N_16378,N_13781,N_14805);
and U16379 (N_16379,N_14866,N_15062);
and U16380 (N_16380,N_12866,N_13261);
nor U16381 (N_16381,N_13289,N_15624);
nand U16382 (N_16382,N_15324,N_14001);
and U16383 (N_16383,N_12929,N_13478);
nand U16384 (N_16384,N_14861,N_15401);
nand U16385 (N_16385,N_14695,N_13578);
nand U16386 (N_16386,N_13337,N_13666);
nor U16387 (N_16387,N_14479,N_12595);
or U16388 (N_16388,N_12682,N_13184);
nor U16389 (N_16389,N_14806,N_15074);
nand U16390 (N_16390,N_12977,N_12739);
and U16391 (N_16391,N_14940,N_15104);
and U16392 (N_16392,N_13069,N_13322);
xnor U16393 (N_16393,N_12863,N_13264);
nand U16394 (N_16394,N_12598,N_15470);
xnor U16395 (N_16395,N_14711,N_12635);
xor U16396 (N_16396,N_15099,N_13891);
and U16397 (N_16397,N_14918,N_15212);
xor U16398 (N_16398,N_15617,N_13335);
xor U16399 (N_16399,N_15368,N_15350);
nor U16400 (N_16400,N_14884,N_13451);
nor U16401 (N_16401,N_12886,N_13698);
nand U16402 (N_16402,N_14615,N_15180);
or U16403 (N_16403,N_14176,N_14864);
and U16404 (N_16404,N_13364,N_13579);
nor U16405 (N_16405,N_13268,N_13283);
and U16406 (N_16406,N_14635,N_15528);
xnor U16407 (N_16407,N_12561,N_12826);
and U16408 (N_16408,N_14669,N_12607);
or U16409 (N_16409,N_14425,N_14031);
xor U16410 (N_16410,N_14116,N_14093);
nand U16411 (N_16411,N_13182,N_13856);
xnor U16412 (N_16412,N_13777,N_14194);
nor U16413 (N_16413,N_13377,N_14844);
and U16414 (N_16414,N_14825,N_15283);
and U16415 (N_16415,N_14520,N_12630);
nor U16416 (N_16416,N_13946,N_15210);
nand U16417 (N_16417,N_13771,N_15267);
and U16418 (N_16418,N_13890,N_15131);
nand U16419 (N_16419,N_12693,N_15572);
nand U16420 (N_16420,N_14597,N_14052);
and U16421 (N_16421,N_15364,N_15146);
or U16422 (N_16422,N_15413,N_13914);
nand U16423 (N_16423,N_13007,N_12987);
or U16424 (N_16424,N_14765,N_13543);
and U16425 (N_16425,N_12959,N_15566);
xnor U16426 (N_16426,N_12848,N_14511);
xnor U16427 (N_16427,N_14392,N_15271);
or U16428 (N_16428,N_14005,N_14030);
and U16429 (N_16429,N_14917,N_14737);
xnor U16430 (N_16430,N_14092,N_12664);
nor U16431 (N_16431,N_13271,N_14671);
nand U16432 (N_16432,N_12939,N_14690);
nor U16433 (N_16433,N_15571,N_12658);
or U16434 (N_16434,N_13290,N_14467);
nor U16435 (N_16435,N_12651,N_13843);
xnor U16436 (N_16436,N_14487,N_14268);
nand U16437 (N_16437,N_14587,N_13558);
nand U16438 (N_16438,N_13479,N_15491);
nand U16439 (N_16439,N_15601,N_15192);
nand U16440 (N_16440,N_13904,N_13618);
nor U16441 (N_16441,N_12941,N_13500);
nand U16442 (N_16442,N_14543,N_12528);
and U16443 (N_16443,N_13319,N_15378);
nor U16444 (N_16444,N_12559,N_14332);
nand U16445 (N_16445,N_14077,N_13689);
nand U16446 (N_16446,N_13742,N_13573);
xor U16447 (N_16447,N_12654,N_14483);
nand U16448 (N_16448,N_15061,N_15371);
nor U16449 (N_16449,N_13293,N_13833);
and U16450 (N_16450,N_13303,N_12641);
or U16451 (N_16451,N_12661,N_13127);
nor U16452 (N_16452,N_15560,N_13749);
xnor U16453 (N_16453,N_12795,N_13294);
nand U16454 (N_16454,N_12548,N_15133);
xor U16455 (N_16455,N_14097,N_13122);
nand U16456 (N_16456,N_15565,N_15254);
xnor U16457 (N_16457,N_14003,N_12999);
and U16458 (N_16458,N_14289,N_14859);
and U16459 (N_16459,N_15352,N_13009);
and U16460 (N_16460,N_14501,N_12677);
and U16461 (N_16461,N_12629,N_14327);
nand U16462 (N_16462,N_14070,N_13963);
xor U16463 (N_16463,N_13376,N_14073);
or U16464 (N_16464,N_14161,N_15112);
xor U16465 (N_16465,N_12985,N_14824);
nand U16466 (N_16466,N_13343,N_13325);
nor U16467 (N_16467,N_14065,N_14415);
xor U16468 (N_16468,N_14147,N_15149);
nand U16469 (N_16469,N_13399,N_13281);
nor U16470 (N_16470,N_14721,N_13285);
nor U16471 (N_16471,N_14228,N_13265);
nand U16472 (N_16472,N_13263,N_15473);
nor U16473 (N_16473,N_14874,N_13656);
nand U16474 (N_16474,N_14411,N_14058);
and U16475 (N_16475,N_12986,N_14360);
and U16476 (N_16476,N_13041,N_13006);
xor U16477 (N_16477,N_13448,N_13622);
and U16478 (N_16478,N_12549,N_13282);
or U16479 (N_16479,N_14681,N_14211);
xor U16480 (N_16480,N_14606,N_15155);
nand U16481 (N_16481,N_13061,N_12871);
and U16482 (N_16482,N_13340,N_12789);
nand U16483 (N_16483,N_14046,N_14647);
or U16484 (N_16484,N_13786,N_13753);
or U16485 (N_16485,N_15288,N_14536);
xor U16486 (N_16486,N_12926,N_15159);
or U16487 (N_16487,N_12877,N_14103);
or U16488 (N_16488,N_14761,N_15089);
and U16489 (N_16489,N_13462,N_14813);
nor U16490 (N_16490,N_12741,N_14526);
and U16491 (N_16491,N_13902,N_13973);
or U16492 (N_16492,N_13672,N_14762);
and U16493 (N_16493,N_13014,N_12869);
xor U16494 (N_16494,N_15361,N_14334);
xor U16495 (N_16495,N_13715,N_15509);
or U16496 (N_16496,N_15422,N_12535);
xnor U16497 (N_16497,N_14608,N_14150);
xnor U16498 (N_16498,N_15222,N_14828);
or U16499 (N_16499,N_14109,N_13825);
or U16500 (N_16500,N_14620,N_13237);
or U16501 (N_16501,N_12796,N_15187);
or U16502 (N_16502,N_13804,N_15221);
or U16503 (N_16503,N_13191,N_13274);
and U16504 (N_16504,N_14033,N_12689);
or U16505 (N_16505,N_13564,N_13630);
nor U16506 (N_16506,N_15451,N_13772);
nand U16507 (N_16507,N_14256,N_12996);
and U16508 (N_16508,N_15080,N_15484);
nor U16509 (N_16509,N_15441,N_14683);
xnor U16510 (N_16510,N_13393,N_14248);
xor U16511 (N_16511,N_15489,N_15500);
nor U16512 (N_16512,N_15456,N_14633);
xor U16513 (N_16513,N_13272,N_15418);
or U16514 (N_16514,N_13597,N_13629);
nand U16515 (N_16515,N_15203,N_14442);
xnor U16516 (N_16516,N_14745,N_13024);
nand U16517 (N_16517,N_14661,N_13829);
or U16518 (N_16518,N_13964,N_13299);
xnor U16519 (N_16519,N_15375,N_14966);
and U16520 (N_16520,N_12611,N_12849);
and U16521 (N_16521,N_14925,N_15407);
xor U16522 (N_16522,N_14915,N_15606);
and U16523 (N_16523,N_15400,N_13036);
and U16524 (N_16524,N_13266,N_14831);
xnor U16525 (N_16525,N_14020,N_15353);
nand U16526 (N_16526,N_14443,N_14121);
nand U16527 (N_16527,N_13590,N_13848);
or U16528 (N_16528,N_15421,N_13894);
and U16529 (N_16529,N_14181,N_14085);
nand U16530 (N_16530,N_14060,N_15431);
or U16531 (N_16531,N_15396,N_14934);
nand U16532 (N_16532,N_14819,N_12508);
and U16533 (N_16533,N_14048,N_13385);
or U16534 (N_16534,N_13110,N_15169);
xor U16535 (N_16535,N_13934,N_13165);
nand U16536 (N_16536,N_13716,N_12531);
nor U16537 (N_16537,N_14982,N_13049);
nor U16538 (N_16538,N_13454,N_14576);
nor U16539 (N_16539,N_15590,N_13747);
nand U16540 (N_16540,N_15009,N_12859);
or U16541 (N_16541,N_13793,N_14075);
xnor U16542 (N_16542,N_15621,N_13791);
nor U16543 (N_16543,N_14559,N_13841);
nand U16544 (N_16544,N_14156,N_14380);
nand U16545 (N_16545,N_13872,N_14993);
nand U16546 (N_16546,N_15507,N_13731);
and U16547 (N_16547,N_14709,N_12545);
xor U16548 (N_16548,N_14458,N_14609);
xnor U16549 (N_16549,N_12716,N_13201);
nand U16550 (N_16550,N_13907,N_14837);
or U16551 (N_16551,N_14404,N_12807);
nand U16552 (N_16552,N_15620,N_13628);
nand U16553 (N_16553,N_14344,N_13065);
or U16554 (N_16554,N_15004,N_12706);
nor U16555 (N_16555,N_13329,N_13316);
xnor U16556 (N_16556,N_13106,N_15412);
nand U16557 (N_16557,N_14652,N_13317);
xor U16558 (N_16558,N_12546,N_14778);
or U16559 (N_16559,N_15505,N_13676);
nand U16560 (N_16560,N_12995,N_14270);
nor U16561 (N_16561,N_15021,N_13760);
nor U16562 (N_16562,N_12822,N_15465);
or U16563 (N_16563,N_14639,N_13095);
nor U16564 (N_16564,N_13970,N_15487);
or U16565 (N_16565,N_13859,N_15538);
or U16566 (N_16566,N_13551,N_15108);
nand U16567 (N_16567,N_14999,N_13217);
nor U16568 (N_16568,N_13331,N_14769);
and U16569 (N_16569,N_12800,N_13074);
nor U16570 (N_16570,N_12532,N_15245);
and U16571 (N_16571,N_13037,N_13667);
nand U16572 (N_16572,N_15284,N_13556);
or U16573 (N_16573,N_12769,N_15047);
and U16574 (N_16574,N_13991,N_15130);
and U16575 (N_16575,N_14027,N_13575);
xnor U16576 (N_16576,N_13839,N_13992);
and U16577 (N_16577,N_14714,N_13449);
and U16578 (N_16578,N_13883,N_15596);
xnor U16579 (N_16579,N_14302,N_14435);
nor U16580 (N_16580,N_12809,N_14758);
and U16581 (N_16581,N_13455,N_15184);
and U16582 (N_16582,N_13645,N_13318);
nor U16583 (N_16583,N_13223,N_14472);
nand U16584 (N_16584,N_14189,N_14674);
and U16585 (N_16585,N_15360,N_14326);
xnor U16586 (N_16586,N_13465,N_14713);
nor U16587 (N_16587,N_12685,N_14396);
nor U16588 (N_16588,N_15002,N_14909);
xnor U16589 (N_16589,N_13257,N_14550);
nand U16590 (N_16590,N_12581,N_13571);
nand U16591 (N_16591,N_14493,N_14465);
and U16592 (N_16592,N_15162,N_14939);
xnor U16593 (N_16593,N_12945,N_13903);
nand U16594 (N_16594,N_13957,N_14054);
nand U16595 (N_16595,N_12971,N_13017);
and U16596 (N_16596,N_13437,N_13912);
or U16597 (N_16597,N_15078,N_14234);
xnor U16598 (N_16598,N_15588,N_15580);
nor U16599 (N_16599,N_15380,N_13588);
or U16600 (N_16600,N_15282,N_15333);
or U16601 (N_16601,N_13495,N_15144);
or U16602 (N_16602,N_13483,N_13999);
nor U16603 (N_16603,N_14710,N_14625);
or U16604 (N_16604,N_15202,N_14658);
nand U16605 (N_16605,N_14388,N_13621);
nand U16606 (N_16606,N_12578,N_14873);
xnor U16607 (N_16607,N_15106,N_14418);
and U16608 (N_16608,N_13750,N_13734);
and U16609 (N_16609,N_13456,N_14632);
nand U16610 (N_16610,N_14942,N_14371);
xor U16611 (N_16611,N_13348,N_14385);
xor U16612 (N_16612,N_14815,N_15134);
xor U16613 (N_16613,N_13763,N_13012);
and U16614 (N_16614,N_15355,N_13179);
nor U16615 (N_16615,N_14975,N_12660);
and U16616 (N_16616,N_13831,N_14878);
nand U16617 (N_16617,N_14282,N_15274);
or U16618 (N_16618,N_14146,N_14514);
xor U16619 (N_16619,N_13056,N_13886);
nand U16620 (N_16620,N_13809,N_14724);
or U16621 (N_16621,N_15398,N_15291);
xor U16622 (N_16622,N_14372,N_15165);
nor U16623 (N_16623,N_14850,N_13719);
or U16624 (N_16624,N_13382,N_14123);
and U16625 (N_16625,N_12514,N_14929);
nor U16626 (N_16626,N_13413,N_13965);
nand U16627 (N_16627,N_14274,N_14792);
nor U16628 (N_16628,N_15524,N_15411);
or U16629 (N_16629,N_12650,N_13208);
or U16630 (N_16630,N_12851,N_13574);
and U16631 (N_16631,N_13885,N_14863);
nand U16632 (N_16632,N_15551,N_14764);
or U16633 (N_16633,N_12505,N_12802);
nor U16634 (N_16634,N_14192,N_12628);
nand U16635 (N_16635,N_12684,N_13801);
nor U16636 (N_16636,N_13233,N_13576);
and U16637 (N_16637,N_13827,N_13730);
nand U16638 (N_16638,N_13030,N_14741);
nor U16639 (N_16639,N_12949,N_15567);
nor U16640 (N_16640,N_13935,N_15269);
nand U16641 (N_16641,N_12645,N_12867);
xor U16642 (N_16642,N_13060,N_12841);
xor U16643 (N_16643,N_14206,N_15409);
and U16644 (N_16644,N_12563,N_13735);
and U16645 (N_16645,N_12737,N_14969);
nand U16646 (N_16646,N_15049,N_14613);
nor U16647 (N_16647,N_14893,N_15372);
xor U16648 (N_16648,N_13262,N_14770);
nand U16649 (N_16649,N_12885,N_14810);
nor U16650 (N_16650,N_13297,N_14469);
xnor U16651 (N_16651,N_13469,N_13746);
nor U16652 (N_16652,N_12574,N_14726);
nor U16653 (N_16653,N_13394,N_14489);
nand U16654 (N_16654,N_13474,N_15223);
or U16655 (N_16655,N_13706,N_14686);
or U16656 (N_16656,N_15425,N_14258);
xnor U16657 (N_16657,N_12873,N_13631);
or U16658 (N_16658,N_15493,N_13864);
nand U16659 (N_16659,N_15297,N_15213);
or U16660 (N_16660,N_15209,N_14946);
or U16661 (N_16661,N_14153,N_14961);
nand U16662 (N_16662,N_14254,N_14535);
and U16663 (N_16663,N_15067,N_12553);
or U16664 (N_16664,N_14619,N_14506);
and U16665 (N_16665,N_14421,N_13740);
xnor U16666 (N_16666,N_13560,N_14203);
and U16667 (N_16667,N_14235,N_13599);
nor U16668 (N_16668,N_13803,N_15303);
and U16669 (N_16669,N_13862,N_15351);
and U16670 (N_16670,N_12613,N_13230);
xnor U16671 (N_16671,N_14708,N_15314);
nor U16672 (N_16672,N_13620,N_12810);
nand U16673 (N_16673,N_14032,N_15137);
nor U16674 (N_16674,N_14080,N_13150);
and U16675 (N_16675,N_14524,N_15091);
xnor U16676 (N_16676,N_13302,N_15123);
or U16677 (N_16677,N_14756,N_12978);
or U16678 (N_16678,N_14495,N_14531);
nand U16679 (N_16679,N_15479,N_12597);
xor U16680 (N_16680,N_15097,N_13306);
nor U16681 (N_16681,N_13250,N_13995);
and U16682 (N_16682,N_14043,N_15501);
xor U16683 (N_16683,N_12665,N_13410);
nand U16684 (N_16684,N_15604,N_14503);
xnor U16685 (N_16685,N_13452,N_14036);
and U16686 (N_16686,N_14673,N_14645);
nand U16687 (N_16687,N_12525,N_13797);
nand U16688 (N_16688,N_12823,N_14856);
nor U16689 (N_16689,N_13214,N_13916);
or U16690 (N_16690,N_14012,N_13869);
nor U16691 (N_16691,N_13372,N_15278);
nor U16692 (N_16692,N_13939,N_13918);
xor U16693 (N_16693,N_14246,N_13161);
nor U16694 (N_16694,N_13926,N_14936);
xor U16695 (N_16695,N_14775,N_14015);
or U16696 (N_16696,N_15466,N_13435);
nor U16697 (N_16697,N_15319,N_13259);
or U16698 (N_16698,N_12733,N_12673);
nor U16699 (N_16699,N_14964,N_13513);
xor U16700 (N_16700,N_15083,N_15013);
xor U16701 (N_16701,N_14623,N_14852);
nand U16702 (N_16702,N_12907,N_14679);
xor U16703 (N_16703,N_12519,N_13702);
xor U16704 (N_16704,N_14401,N_14322);
and U16705 (N_16705,N_14025,N_15177);
or U16706 (N_16706,N_13899,N_15211);
and U16707 (N_16707,N_15525,N_14325);
xor U16708 (N_16708,N_12667,N_14152);
and U16709 (N_16709,N_14209,N_15603);
nand U16710 (N_16710,N_14800,N_13765);
nor U16711 (N_16711,N_14567,N_13519);
nor U16712 (N_16712,N_15555,N_12702);
nor U16713 (N_16713,N_13641,N_14895);
nand U16714 (N_16714,N_12615,N_14682);
nand U16715 (N_16715,N_14995,N_12901);
or U16716 (N_16716,N_12980,N_14638);
xnor U16717 (N_16717,N_14759,N_12518);
or U16718 (N_16718,N_12897,N_12787);
nor U16719 (N_16719,N_13215,N_15029);
xor U16720 (N_16720,N_13984,N_12610);
and U16721 (N_16721,N_13114,N_15595);
nor U16722 (N_16722,N_12604,N_15335);
xnor U16723 (N_16723,N_14237,N_12876);
and U16724 (N_16724,N_15160,N_14291);
nor U16725 (N_16725,N_13799,N_14454);
nor U16726 (N_16726,N_13494,N_14872);
xnor U16727 (N_16727,N_14565,N_13602);
or U16728 (N_16728,N_13321,N_13387);
xnor U16729 (N_16729,N_13851,N_12804);
nand U16730 (N_16730,N_14640,N_14836);
nand U16731 (N_16731,N_13836,N_12839);
and U16732 (N_16732,N_12500,N_15584);
or U16733 (N_16733,N_13530,N_12720);
or U16734 (N_16734,N_13134,N_12589);
and U16735 (N_16735,N_12751,N_13830);
or U16736 (N_16736,N_14059,N_14963);
and U16737 (N_16737,N_13003,N_13601);
xor U16738 (N_16738,N_14869,N_13028);
or U16739 (N_16739,N_14130,N_13632);
nand U16740 (N_16740,N_15188,N_14298);
nand U16741 (N_16741,N_15017,N_15232);
xnor U16742 (N_16742,N_14131,N_14949);
and U16743 (N_16743,N_12709,N_13344);
nor U16744 (N_16744,N_13067,N_12970);
nand U16745 (N_16745,N_14281,N_14461);
or U16746 (N_16746,N_12829,N_14141);
or U16747 (N_16747,N_13518,N_13981);
nand U16748 (N_16748,N_15100,N_14971);
and U16749 (N_16749,N_13366,N_13802);
nor U16750 (N_16750,N_14913,N_14897);
nand U16751 (N_16751,N_15520,N_14967);
or U16752 (N_16752,N_13674,N_14118);
xnor U16753 (N_16753,N_13690,N_13108);
nand U16754 (N_16754,N_14321,N_14296);
and U16755 (N_16755,N_13485,N_12947);
nand U16756 (N_16756,N_13048,N_14389);
or U16757 (N_16757,N_13808,N_14562);
xnor U16758 (N_16758,N_12828,N_15376);
and U16759 (N_16759,N_12758,N_14430);
or U16760 (N_16760,N_14862,N_14293);
and U16761 (N_16761,N_13341,N_15205);
and U16762 (N_16762,N_13834,N_12731);
and U16763 (N_16763,N_13441,N_14339);
or U16764 (N_16764,N_12946,N_15052);
and U16765 (N_16765,N_13071,N_15092);
and U16766 (N_16766,N_14218,N_15342);
nand U16767 (N_16767,N_14446,N_14304);
nor U16768 (N_16768,N_14840,N_14911);
or U16769 (N_16769,N_13531,N_14529);
or U16770 (N_16770,N_13875,N_15447);
or U16771 (N_16771,N_12922,N_13736);
and U16772 (N_16772,N_13447,N_13849);
nor U16773 (N_16773,N_14081,N_12955);
nand U16774 (N_16774,N_14718,N_13967);
nor U16775 (N_16775,N_12606,N_14354);
xnor U16776 (N_16776,N_14311,N_12565);
xnor U16777 (N_16777,N_14349,N_12920);
xnor U16778 (N_16778,N_12526,N_12742);
or U16779 (N_16779,N_14320,N_15533);
xnor U16780 (N_16780,N_13499,N_15444);
and U16781 (N_16781,N_15316,N_13330);
and U16782 (N_16782,N_13826,N_13373);
xor U16783 (N_16783,N_12502,N_12759);
nand U16784 (N_16784,N_14540,N_13146);
or U16785 (N_16785,N_14793,N_13790);
and U16786 (N_16786,N_13874,N_14230);
nand U16787 (N_16787,N_13356,N_14797);
nand U16788 (N_16788,N_12912,N_12678);
nand U16789 (N_16789,N_15395,N_14038);
and U16790 (N_16790,N_13368,N_13721);
and U16791 (N_16791,N_13308,N_13481);
xor U16792 (N_16792,N_14662,N_14199);
nand U16793 (N_16793,N_14983,N_13128);
nor U16794 (N_16794,N_13677,N_14629);
or U16795 (N_16795,N_14004,N_15120);
and U16796 (N_16796,N_13712,N_14978);
or U16797 (N_16797,N_13816,N_13168);
or U16798 (N_16798,N_12940,N_14931);
or U16799 (N_16799,N_12637,N_13775);
xor U16800 (N_16800,N_13276,N_14000);
xor U16801 (N_16801,N_14627,N_15320);
nand U16802 (N_16802,N_13528,N_13610);
xor U16803 (N_16803,N_14047,N_15534);
nand U16804 (N_16804,N_13923,N_13955);
and U16805 (N_16805,N_13211,N_12541);
or U16806 (N_16806,N_12730,N_13386);
nand U16807 (N_16807,N_13354,N_13226);
and U16808 (N_16808,N_14317,N_14768);
nand U16809 (N_16809,N_15012,N_14148);
or U16810 (N_16810,N_14626,N_14428);
nor U16811 (N_16811,N_13585,N_13925);
and U16812 (N_16812,N_14140,N_12786);
nor U16813 (N_16813,N_14871,N_13744);
nor U16814 (N_16814,N_15014,N_13542);
and U16815 (N_16815,N_14868,N_15153);
and U16816 (N_16816,N_15119,N_14305);
or U16817 (N_16817,N_15591,N_13270);
and U16818 (N_16818,N_13148,N_14335);
and U16819 (N_16819,N_15285,N_14471);
or U16820 (N_16820,N_14497,N_15496);
and U16821 (N_16821,N_15256,N_14173);
nand U16822 (N_16822,N_14860,N_13352);
nand U16823 (N_16823,N_13650,N_13126);
and U16824 (N_16824,N_13795,N_14019);
and U16825 (N_16825,N_15296,N_15475);
or U16826 (N_16826,N_12843,N_13687);
nand U16827 (N_16827,N_14890,N_12579);
or U16828 (N_16828,N_14563,N_14833);
or U16829 (N_16829,N_15277,N_12794);
and U16830 (N_16830,N_12655,N_12956);
nand U16831 (N_16831,N_15042,N_12536);
or U16832 (N_16832,N_14589,N_14858);
xnor U16833 (N_16833,N_13207,N_15309);
or U16834 (N_16834,N_14812,N_15084);
or U16835 (N_16835,N_14243,N_15270);
and U16836 (N_16836,N_12781,N_12503);
or U16837 (N_16837,N_14725,N_13187);
or U16838 (N_16838,N_15581,N_14572);
nand U16839 (N_16839,N_14341,N_14017);
nand U16840 (N_16840,N_14881,N_15195);
nand U16841 (N_16841,N_13552,N_14555);
or U16842 (N_16842,N_13094,N_15485);
or U16843 (N_16843,N_14557,N_13913);
and U16844 (N_16844,N_15495,N_13895);
nor U16845 (N_16845,N_12695,N_13908);
nand U16846 (N_16846,N_13288,N_15494);
or U16847 (N_16847,N_13016,N_14750);
nor U16848 (N_16848,N_15513,N_13559);
or U16849 (N_16849,N_13004,N_15550);
or U16850 (N_16850,N_15128,N_13713);
nand U16851 (N_16851,N_13390,N_12990);
nand U16852 (N_16852,N_14278,N_12687);
nand U16853 (N_16853,N_15101,N_14693);
nor U16854 (N_16854,N_13840,N_14854);
nor U16855 (N_16855,N_15476,N_13047);
nand U16856 (N_16856,N_13665,N_12894);
nor U16857 (N_16857,N_13718,N_14191);
nor U16858 (N_16858,N_14390,N_13905);
nand U16859 (N_16859,N_13442,N_13360);
or U16860 (N_16860,N_14202,N_13088);
nand U16861 (N_16861,N_13139,N_15252);
and U16862 (N_16862,N_14481,N_14875);
or U16863 (N_16863,N_13517,N_14904);
nand U16864 (N_16864,N_13486,N_15026);
or U16865 (N_16865,N_13310,N_14740);
xnor U16866 (N_16866,N_14134,N_13388);
nor U16867 (N_16867,N_12729,N_13817);
and U16868 (N_16868,N_15023,N_15201);
and U16869 (N_16869,N_15419,N_15111);
nor U16870 (N_16870,N_13345,N_14666);
xnor U16871 (N_16871,N_13459,N_14262);
or U16872 (N_16872,N_13425,N_14227);
nor U16873 (N_16873,N_14079,N_14069);
nand U16874 (N_16874,N_15048,N_12567);
or U16875 (N_16875,N_12814,N_13828);
nor U16876 (N_16876,N_14573,N_14603);
and U16877 (N_16877,N_12705,N_14776);
and U16878 (N_16878,N_14364,N_13038);
or U16879 (N_16879,N_14205,N_14250);
xnor U16880 (N_16880,N_15085,N_15600);
or U16881 (N_16881,N_13457,N_12836);
and U16882 (N_16882,N_13117,N_15006);
nor U16883 (N_16883,N_14383,N_13861);
or U16884 (N_16884,N_15073,N_13529);
or U16885 (N_16885,N_13280,N_13660);
and U16886 (N_16886,N_15237,N_13407);
or U16887 (N_16887,N_14450,N_14558);
or U16888 (N_16888,N_14301,N_15549);
xnor U16889 (N_16889,N_13614,N_12834);
nand U16890 (N_16890,N_13378,N_14251);
nand U16891 (N_16891,N_12811,N_13398);
xor U16892 (N_16892,N_14631,N_15437);
nand U16893 (N_16893,N_13497,N_13889);
nand U16894 (N_16894,N_15235,N_14843);
nor U16895 (N_16895,N_12719,N_15611);
nor U16896 (N_16896,N_14784,N_14643);
or U16897 (N_16897,N_15295,N_13756);
nand U16898 (N_16898,N_15543,N_14413);
and U16899 (N_16899,N_14730,N_15416);
and U16900 (N_16900,N_14407,N_13002);
xor U16901 (N_16901,N_15317,N_13534);
and U16902 (N_16902,N_15619,N_13737);
nand U16903 (N_16903,N_12576,N_13445);
nand U16904 (N_16904,N_12609,N_15472);
xor U16905 (N_16905,N_14346,N_12608);
nand U16906 (N_16906,N_14968,N_14581);
nand U16907 (N_16907,N_13723,N_15341);
or U16908 (N_16908,N_14398,N_14622);
or U16909 (N_16909,N_12982,N_12874);
xnor U16910 (N_16910,N_13523,N_14292);
and U16911 (N_16911,N_12568,N_14823);
or U16912 (N_16912,N_14556,N_12646);
or U16913 (N_16913,N_14699,N_13986);
nand U16914 (N_16914,N_14236,N_14275);
xor U16915 (N_16915,N_12783,N_14444);
and U16916 (N_16916,N_14111,N_12617);
nor U16917 (N_16917,N_14849,N_13728);
nor U16918 (N_16918,N_13013,N_14106);
nor U16919 (N_16919,N_13301,N_12988);
nand U16920 (N_16920,N_13197,N_13339);
or U16921 (N_16921,N_12639,N_12820);
nand U16922 (N_16922,N_13247,N_12774);
xor U16923 (N_16923,N_15075,N_15186);
xor U16924 (N_16924,N_14996,N_13636);
and U16925 (N_16925,N_15349,N_15163);
or U16926 (N_16926,N_13509,N_13854);
xor U16927 (N_16927,N_15544,N_13307);
nand U16928 (N_16928,N_15382,N_12989);
and U16929 (N_16929,N_14935,N_15469);
nand U16930 (N_16930,N_14474,N_13586);
nor U16931 (N_16931,N_13019,N_14500);
nor U16932 (N_16932,N_15460,N_15255);
nand U16933 (N_16933,N_14287,N_15262);
xnor U16934 (N_16934,N_14280,N_15005);
nor U16935 (N_16935,N_12622,N_14391);
or U16936 (N_16936,N_14575,N_13678);
or U16937 (N_16937,N_15392,N_13082);
or U16938 (N_16938,N_14984,N_13748);
or U16939 (N_16939,N_14361,N_13767);
or U16940 (N_16940,N_14484,N_13020);
and U16941 (N_16941,N_14664,N_13424);
nand U16942 (N_16942,N_14701,N_13468);
nand U16943 (N_16943,N_15266,N_12627);
and U16944 (N_16944,N_13616,N_14051);
or U16945 (N_16945,N_14574,N_13160);
xor U16946 (N_16946,N_14172,N_15055);
and U16947 (N_16947,N_12696,N_15618);
or U16948 (N_16948,N_15607,N_13218);
xnor U16949 (N_16949,N_14696,N_12760);
xnor U16950 (N_16950,N_14899,N_15579);
nand U16951 (N_16951,N_15135,N_13652);
or U16952 (N_16952,N_12512,N_14286);
or U16953 (N_16953,N_15294,N_12815);
or U16954 (N_16954,N_12593,N_12754);
or U16955 (N_16955,N_13906,N_14449);
nor U16956 (N_16956,N_13987,N_13811);
and U16957 (N_16957,N_13929,N_15070);
or U16958 (N_16958,N_13379,N_13089);
xnor U16959 (N_16959,N_15377,N_15535);
or U16960 (N_16960,N_12952,N_13953);
nor U16961 (N_16961,N_13917,N_14600);
xnor U16962 (N_16962,N_13422,N_12653);
nand U16963 (N_16963,N_15208,N_14438);
nor U16964 (N_16964,N_15000,N_14544);
xnor U16965 (N_16965,N_15344,N_13467);
or U16966 (N_16966,N_15439,N_12776);
nand U16967 (N_16967,N_14648,N_14378);
and U16968 (N_16968,N_13210,N_15236);
xor U16969 (N_16969,N_12798,N_14102);
and U16970 (N_16970,N_13482,N_14358);
nor U16971 (N_16971,N_14515,N_15059);
nand U16972 (N_16972,N_13659,N_14787);
nand U16973 (N_16973,N_13951,N_13186);
and U16974 (N_16974,N_12831,N_14403);
xnor U16975 (N_16975,N_12942,N_14094);
xnor U16976 (N_16976,N_15474,N_15365);
nor U16977 (N_16977,N_15261,N_13668);
and U16978 (N_16978,N_13683,N_13858);
and U16979 (N_16979,N_15486,N_15010);
or U16980 (N_16980,N_13681,N_15173);
and U16981 (N_16981,N_13443,N_14494);
nand U16982 (N_16982,N_13243,N_13878);
nor U16983 (N_16983,N_14333,N_15060);
and U16984 (N_16984,N_13662,N_14429);
nor U16985 (N_16985,N_13776,N_13332);
or U16986 (N_16986,N_14668,N_14127);
or U16987 (N_16987,N_12683,N_14950);
and U16988 (N_16988,N_14841,N_15478);
nor U16989 (N_16989,N_14582,N_13063);
and U16990 (N_16990,N_13204,N_13078);
nand U16991 (N_16991,N_12779,N_15079);
or U16992 (N_16992,N_14162,N_15027);
xor U16993 (N_16993,N_14432,N_12976);
xor U16994 (N_16994,N_14451,N_12564);
nand U16995 (N_16995,N_14653,N_14777);
or U16996 (N_16996,N_14045,N_13787);
nand U16997 (N_16997,N_14634,N_14224);
xnor U16998 (N_16998,N_13140,N_15241);
nor U16999 (N_16999,N_15519,N_15182);
nor U17000 (N_17000,N_13682,N_14955);
nand U17001 (N_17001,N_14937,N_13994);
or U17002 (N_17002,N_15063,N_15337);
nor U17003 (N_17003,N_14128,N_15141);
nor U17004 (N_17004,N_15598,N_13183);
and U17005 (N_17005,N_14456,N_13752);
nand U17006 (N_17006,N_15332,N_13488);
xnor U17007 (N_17007,N_14599,N_13357);
and U17008 (N_17008,N_14651,N_14987);
and U17009 (N_17009,N_14071,N_14464);
nor U17010 (N_17010,N_13031,N_15164);
nand U17011 (N_17011,N_12975,N_14794);
xnor U17012 (N_17012,N_15043,N_14174);
or U17013 (N_17013,N_15417,N_13819);
or U17014 (N_17014,N_13933,N_12799);
nor U17015 (N_17015,N_15330,N_12948);
xor U17016 (N_17016,N_14702,N_14184);
and U17017 (N_17017,N_14416,N_14232);
and U17018 (N_17018,N_13754,N_14663);
nand U17019 (N_17019,N_12884,N_13181);
nand U17020 (N_17020,N_15175,N_14242);
xnor U17021 (N_17021,N_13846,N_15585);
nor U17022 (N_17022,N_13606,N_15370);
xor U17023 (N_17023,N_14903,N_15025);
and U17024 (N_17024,N_14104,N_13397);
and U17025 (N_17025,N_15161,N_12927);
nor U17026 (N_17026,N_13711,N_14952);
and U17027 (N_17027,N_13915,N_13699);
or U17028 (N_17028,N_14434,N_13504);
or U17029 (N_17029,N_13820,N_14814);
or U17030 (N_17030,N_13640,N_14734);
nand U17031 (N_17031,N_14142,N_13569);
nand U17032 (N_17032,N_13966,N_15265);
nand U17033 (N_17033,N_13512,N_14546);
or U17034 (N_17034,N_15158,N_12746);
and U17035 (N_17035,N_12827,N_13075);
nor U17036 (N_17036,N_13806,N_14313);
xnor U17037 (N_17037,N_14771,N_12934);
xor U17038 (N_17038,N_13876,N_15394);
nor U17039 (N_17039,N_13669,N_13402);
nor U17040 (N_17040,N_13554,N_13323);
and U17041 (N_17041,N_13927,N_12560);
nand U17042 (N_17042,N_12711,N_15356);
or U17043 (N_17043,N_14539,N_14330);
nor U17044 (N_17044,N_13670,N_12943);
xnor U17045 (N_17045,N_12862,N_12816);
nand U17046 (N_17046,N_12745,N_15410);
and U17047 (N_17047,N_15423,N_13975);
xor U17048 (N_17048,N_14650,N_15136);
nor U17049 (N_17049,N_14229,N_14063);
or U17050 (N_17050,N_13496,N_14393);
nand U17051 (N_17051,N_15240,N_13532);
and U17052 (N_17052,N_12778,N_14706);
xnor U17053 (N_17053,N_12790,N_12555);
nand U17054 (N_17054,N_13587,N_14977);
xor U17055 (N_17055,N_15054,N_12763);
nor U17056 (N_17056,N_13501,N_13949);
or U17057 (N_17057,N_13029,N_15139);
nand U17058 (N_17058,N_13739,N_15480);
xnor U17059 (N_17059,N_13245,N_12623);
xor U17060 (N_17060,N_14035,N_13130);
and U17061 (N_17061,N_15157,N_12921);
and U17062 (N_17062,N_13800,N_14598);
nor U17063 (N_17063,N_12539,N_13608);
and U17064 (N_17064,N_15065,N_15623);
and U17065 (N_17065,N_13164,N_15194);
nor U17066 (N_17066,N_15582,N_14086);
xor U17067 (N_17067,N_14362,N_14785);
and U17068 (N_17068,N_13077,N_15003);
or U17069 (N_17069,N_14277,N_15107);
or U17070 (N_17070,N_13838,N_13428);
xor U17071 (N_17071,N_13111,N_15105);
nand U17072 (N_17072,N_15181,N_13032);
nor U17073 (N_17073,N_14410,N_12718);
and U17074 (N_17074,N_14593,N_12506);
or U17075 (N_17075,N_14259,N_14316);
xor U17076 (N_17076,N_13589,N_12726);
nor U17077 (N_17077,N_12636,N_15362);
xor U17078 (N_17078,N_14213,N_15093);
or U17079 (N_17079,N_15448,N_13489);
or U17080 (N_17080,N_12856,N_13567);
xor U17081 (N_17081,N_15311,N_13867);
nand U17082 (N_17082,N_12817,N_12770);
or U17083 (N_17083,N_13900,N_14090);
or U17084 (N_17084,N_13996,N_13241);
nor U17085 (N_17085,N_13021,N_14739);
and U17086 (N_17086,N_12788,N_15132);
nor U17087 (N_17087,N_13000,N_15406);
nand U17088 (N_17088,N_13177,N_15408);
xor U17089 (N_17089,N_15433,N_13156);
or U17090 (N_17090,N_14928,N_13005);
or U17091 (N_17091,N_13091,N_14723);
nor U17092 (N_17092,N_12515,N_12599);
and U17093 (N_17093,N_13355,N_13149);
nand U17094 (N_17094,N_14857,N_14108);
nor U17095 (N_17095,N_14738,N_13562);
nand U17096 (N_17096,N_14989,N_13960);
nor U17097 (N_17097,N_13769,N_13675);
or U17098 (N_17098,N_14644,N_13969);
nor U17099 (N_17099,N_15249,N_15189);
nand U17100 (N_17100,N_15348,N_13807);
nand U17101 (N_17101,N_13473,N_13686);
xor U17102 (N_17102,N_14549,N_13643);
nand U17103 (N_17103,N_14023,N_14240);
and U17104 (N_17104,N_13178,N_13116);
or U17105 (N_17105,N_13694,N_12868);
xor U17106 (N_17106,N_15001,N_13246);
xnor U17107 (N_17107,N_13392,N_14896);
xor U17108 (N_17108,N_13520,N_13952);
and U17109 (N_17109,N_13577,N_12569);
and U17110 (N_17110,N_14607,N_13701);
and U17111 (N_17111,N_15218,N_15403);
nand U17112 (N_17112,N_15096,N_12551);
or U17113 (N_17113,N_14263,N_15546);
nor U17114 (N_17114,N_14646,N_14684);
or U17115 (N_17115,N_14271,N_13253);
nand U17116 (N_17116,N_15426,N_14655);
nand U17117 (N_17117,N_15313,N_15587);
xor U17118 (N_17118,N_14512,N_13367);
and U17119 (N_17119,N_13086,N_14331);
or U17120 (N_17120,N_14496,N_12504);
nor U17121 (N_17121,N_13472,N_14788);
xor U17122 (N_17122,N_13196,N_14276);
nor U17123 (N_17123,N_13653,N_12963);
xnor U17124 (N_17124,N_12755,N_12803);
or U17125 (N_17125,N_14175,N_12570);
nand U17126 (N_17126,N_14746,N_12556);
and U17127 (N_17127,N_14530,N_12917);
nor U17128 (N_17128,N_13001,N_13328);
nand U17129 (N_17129,N_13491,N_13416);
xor U17130 (N_17130,N_13540,N_12793);
or U17131 (N_17131,N_13644,N_14374);
and U17132 (N_17132,N_13158,N_13255);
nand U17133 (N_17133,N_13930,N_14888);
xnor U17134 (N_17134,N_13733,N_15030);
nand U17135 (N_17135,N_14932,N_12527);
xnor U17136 (N_17136,N_14976,N_13649);
nor U17137 (N_17137,N_15090,N_14578);
xor U17138 (N_17138,N_14119,N_12625);
nand U17139 (N_17139,N_12620,N_14735);
xnor U17140 (N_17140,N_13625,N_14095);
nand U17141 (N_17141,N_13570,N_13251);
nand U17142 (N_17142,N_13076,N_14433);
or U17143 (N_17143,N_13336,N_14353);
and U17144 (N_17144,N_14377,N_12785);
nor U17145 (N_17145,N_15244,N_14314);
xnor U17146 (N_17146,N_12712,N_13188);
and U17147 (N_17147,N_14779,N_14447);
xor U17148 (N_17148,N_12540,N_13118);
nor U17149 (N_17149,N_13120,N_15599);
or U17150 (N_17150,N_13163,N_13324);
xor U17151 (N_17151,N_14208,N_13115);
nand U17152 (N_17152,N_15166,N_14675);
or U17153 (N_17153,N_12906,N_14807);
nor U17154 (N_17154,N_12890,N_14066);
xnor U17155 (N_17155,N_13947,N_14078);
nand U17156 (N_17156,N_12806,N_14266);
nor U17157 (N_17157,N_13359,N_14457);
and U17158 (N_17158,N_15214,N_13121);
xor U17159 (N_17159,N_13815,N_15573);
or U17160 (N_17160,N_13547,N_14564);
nor U17161 (N_17161,N_12875,N_13400);
xnor U17162 (N_17162,N_15497,N_14216);
nor U17163 (N_17163,N_14855,N_14252);
or U17164 (N_17164,N_15522,N_15357);
nor U17165 (N_17165,N_13057,N_13480);
and U17166 (N_17166,N_12643,N_12734);
nand U17167 (N_17167,N_13600,N_14991);
xor U17168 (N_17168,N_15183,N_13180);
nand U17169 (N_17169,N_13506,N_14351);
nor U17170 (N_17170,N_14533,N_15056);
nor U17171 (N_17171,N_12585,N_13133);
nor U17172 (N_17172,N_14053,N_13510);
or U17173 (N_17173,N_14839,N_13910);
or U17174 (N_17174,N_15393,N_14518);
nor U17175 (N_17175,N_13627,N_13511);
xnor U17176 (N_17176,N_15506,N_15034);
xnor U17177 (N_17177,N_14958,N_13533);
nor U17178 (N_17178,N_14611,N_15306);
or U17179 (N_17179,N_14399,N_15440);
nand U17180 (N_17180,N_15114,N_14595);
or U17181 (N_17181,N_13972,N_15233);
nand U17182 (N_17182,N_12723,N_12727);
or U17183 (N_17183,N_13928,N_14087);
nor U17184 (N_17184,N_15563,N_13046);
and U17185 (N_17185,N_14923,N_13423);
xor U17186 (N_17186,N_15154,N_14050);
or U17187 (N_17187,N_12676,N_14313);
and U17188 (N_17188,N_15231,N_15606);
nor U17189 (N_17189,N_14133,N_15193);
nor U17190 (N_17190,N_14645,N_15593);
xnor U17191 (N_17191,N_14880,N_15597);
and U17192 (N_17192,N_13058,N_13851);
nor U17193 (N_17193,N_14942,N_14519);
nor U17194 (N_17194,N_13229,N_14079);
or U17195 (N_17195,N_15390,N_12864);
xor U17196 (N_17196,N_12856,N_13155);
or U17197 (N_17197,N_13723,N_12938);
and U17198 (N_17198,N_14925,N_14637);
xnor U17199 (N_17199,N_14803,N_15503);
or U17200 (N_17200,N_14875,N_12522);
or U17201 (N_17201,N_13884,N_13422);
nor U17202 (N_17202,N_14189,N_15158);
or U17203 (N_17203,N_14585,N_15366);
and U17204 (N_17204,N_13037,N_12829);
nand U17205 (N_17205,N_14766,N_13935);
nor U17206 (N_17206,N_15365,N_14939);
and U17207 (N_17207,N_13173,N_14459);
xor U17208 (N_17208,N_12921,N_13449);
xnor U17209 (N_17209,N_13668,N_13218);
and U17210 (N_17210,N_13206,N_15246);
nor U17211 (N_17211,N_13626,N_15048);
and U17212 (N_17212,N_13957,N_12975);
or U17213 (N_17213,N_13354,N_13953);
and U17214 (N_17214,N_12756,N_12892);
or U17215 (N_17215,N_13091,N_15416);
nor U17216 (N_17216,N_15177,N_14633);
nor U17217 (N_17217,N_12905,N_15174);
and U17218 (N_17218,N_13580,N_13355);
nand U17219 (N_17219,N_14784,N_14589);
xor U17220 (N_17220,N_15185,N_14655);
nor U17221 (N_17221,N_13943,N_14974);
nor U17222 (N_17222,N_13197,N_13417);
or U17223 (N_17223,N_13120,N_12550);
nand U17224 (N_17224,N_14442,N_14553);
and U17225 (N_17225,N_15035,N_14762);
and U17226 (N_17226,N_14007,N_15096);
or U17227 (N_17227,N_15439,N_14029);
and U17228 (N_17228,N_13601,N_14275);
nand U17229 (N_17229,N_13128,N_14572);
and U17230 (N_17230,N_13518,N_15389);
and U17231 (N_17231,N_14714,N_14020);
nor U17232 (N_17232,N_13095,N_13078);
and U17233 (N_17233,N_12846,N_13434);
and U17234 (N_17234,N_14430,N_12802);
and U17235 (N_17235,N_13447,N_14494);
xor U17236 (N_17236,N_13158,N_15438);
and U17237 (N_17237,N_12584,N_13399);
nor U17238 (N_17238,N_13670,N_15324);
nand U17239 (N_17239,N_12707,N_13070);
and U17240 (N_17240,N_13188,N_12622);
xnor U17241 (N_17241,N_15195,N_12683);
nor U17242 (N_17242,N_12785,N_15434);
nand U17243 (N_17243,N_13320,N_13871);
or U17244 (N_17244,N_12849,N_15472);
or U17245 (N_17245,N_15283,N_13266);
or U17246 (N_17246,N_13448,N_13942);
nor U17247 (N_17247,N_13943,N_14201);
nor U17248 (N_17248,N_14474,N_14015);
nand U17249 (N_17249,N_15162,N_14102);
xor U17250 (N_17250,N_13844,N_13600);
nor U17251 (N_17251,N_15329,N_14087);
or U17252 (N_17252,N_14156,N_12831);
nor U17253 (N_17253,N_13896,N_15080);
nor U17254 (N_17254,N_15129,N_12570);
nand U17255 (N_17255,N_15502,N_14831);
nand U17256 (N_17256,N_15073,N_14075);
and U17257 (N_17257,N_14718,N_15032);
and U17258 (N_17258,N_15293,N_15071);
and U17259 (N_17259,N_13268,N_14731);
and U17260 (N_17260,N_14665,N_13038);
and U17261 (N_17261,N_13225,N_14251);
or U17262 (N_17262,N_13836,N_13567);
or U17263 (N_17263,N_13685,N_13937);
nor U17264 (N_17264,N_14975,N_14945);
and U17265 (N_17265,N_14418,N_14330);
and U17266 (N_17266,N_15019,N_13597);
xnor U17267 (N_17267,N_14081,N_12808);
and U17268 (N_17268,N_14877,N_13868);
and U17269 (N_17269,N_13460,N_12615);
nand U17270 (N_17270,N_14792,N_14278);
or U17271 (N_17271,N_14378,N_15048);
and U17272 (N_17272,N_12625,N_12680);
nor U17273 (N_17273,N_13870,N_13542);
nand U17274 (N_17274,N_12651,N_15577);
nand U17275 (N_17275,N_15196,N_13343);
and U17276 (N_17276,N_14373,N_12674);
nor U17277 (N_17277,N_15245,N_15575);
and U17278 (N_17278,N_13630,N_15030);
or U17279 (N_17279,N_14013,N_15092);
or U17280 (N_17280,N_14080,N_15254);
and U17281 (N_17281,N_14960,N_15127);
or U17282 (N_17282,N_14831,N_12749);
or U17283 (N_17283,N_15107,N_13323);
nand U17284 (N_17284,N_14476,N_13767);
or U17285 (N_17285,N_13210,N_14655);
xor U17286 (N_17286,N_15134,N_12971);
xnor U17287 (N_17287,N_12832,N_14890);
and U17288 (N_17288,N_12908,N_14756);
nor U17289 (N_17289,N_13658,N_13457);
nor U17290 (N_17290,N_14155,N_14149);
nor U17291 (N_17291,N_13865,N_14925);
nand U17292 (N_17292,N_12528,N_12628);
or U17293 (N_17293,N_13425,N_15447);
nand U17294 (N_17294,N_12655,N_13592);
nand U17295 (N_17295,N_12737,N_15624);
or U17296 (N_17296,N_14714,N_12966);
nor U17297 (N_17297,N_15394,N_14347);
nand U17298 (N_17298,N_13745,N_13040);
or U17299 (N_17299,N_13386,N_14298);
or U17300 (N_17300,N_12857,N_15401);
or U17301 (N_17301,N_14294,N_14926);
and U17302 (N_17302,N_13169,N_13065);
nor U17303 (N_17303,N_14213,N_14398);
and U17304 (N_17304,N_14053,N_14181);
or U17305 (N_17305,N_14858,N_12559);
or U17306 (N_17306,N_14045,N_13623);
nand U17307 (N_17307,N_13500,N_14185);
nand U17308 (N_17308,N_15169,N_15269);
and U17309 (N_17309,N_14024,N_13469);
nand U17310 (N_17310,N_13477,N_13188);
and U17311 (N_17311,N_15407,N_14994);
nand U17312 (N_17312,N_12762,N_15297);
or U17313 (N_17313,N_14991,N_13425);
nor U17314 (N_17314,N_15080,N_14857);
nor U17315 (N_17315,N_15407,N_15000);
and U17316 (N_17316,N_14147,N_14836);
nand U17317 (N_17317,N_14299,N_12527);
nand U17318 (N_17318,N_12915,N_15102);
nand U17319 (N_17319,N_12598,N_13287);
nor U17320 (N_17320,N_12673,N_15376);
or U17321 (N_17321,N_13767,N_13996);
and U17322 (N_17322,N_14686,N_14840);
nor U17323 (N_17323,N_15367,N_14920);
nand U17324 (N_17324,N_12979,N_13204);
nand U17325 (N_17325,N_13630,N_12885);
xnor U17326 (N_17326,N_13356,N_14492);
nand U17327 (N_17327,N_14387,N_13789);
or U17328 (N_17328,N_13880,N_13989);
nand U17329 (N_17329,N_15528,N_13962);
and U17330 (N_17330,N_13697,N_13448);
nor U17331 (N_17331,N_12834,N_13704);
nor U17332 (N_17332,N_13439,N_15432);
or U17333 (N_17333,N_14725,N_13436);
nor U17334 (N_17334,N_15471,N_14105);
and U17335 (N_17335,N_14061,N_15354);
xor U17336 (N_17336,N_13147,N_14068);
or U17337 (N_17337,N_12913,N_13368);
nor U17338 (N_17338,N_13346,N_14230);
nand U17339 (N_17339,N_12522,N_15362);
or U17340 (N_17340,N_13492,N_13084);
nand U17341 (N_17341,N_14005,N_15166);
nand U17342 (N_17342,N_14548,N_14231);
or U17343 (N_17343,N_13765,N_13352);
nor U17344 (N_17344,N_12751,N_13130);
and U17345 (N_17345,N_14985,N_13614);
xnor U17346 (N_17346,N_12712,N_14641);
or U17347 (N_17347,N_15301,N_13651);
nor U17348 (N_17348,N_13204,N_13028);
xor U17349 (N_17349,N_13860,N_12889);
nand U17350 (N_17350,N_15392,N_13781);
and U17351 (N_17351,N_12715,N_13295);
nand U17352 (N_17352,N_12503,N_13767);
xnor U17353 (N_17353,N_14377,N_13915);
nand U17354 (N_17354,N_13723,N_14544);
nand U17355 (N_17355,N_15564,N_15403);
nand U17356 (N_17356,N_12992,N_14678);
and U17357 (N_17357,N_13984,N_12579);
and U17358 (N_17358,N_14738,N_12643);
or U17359 (N_17359,N_15198,N_14465);
or U17360 (N_17360,N_12909,N_14669);
and U17361 (N_17361,N_13962,N_15152);
xnor U17362 (N_17362,N_15505,N_13790);
and U17363 (N_17363,N_15176,N_13316);
nand U17364 (N_17364,N_14043,N_14562);
nor U17365 (N_17365,N_12966,N_13956);
nand U17366 (N_17366,N_14074,N_14679);
xnor U17367 (N_17367,N_13834,N_15151);
or U17368 (N_17368,N_14816,N_15279);
nand U17369 (N_17369,N_13859,N_15233);
and U17370 (N_17370,N_13654,N_13398);
and U17371 (N_17371,N_15554,N_14874);
and U17372 (N_17372,N_15353,N_13942);
nor U17373 (N_17373,N_14682,N_14585);
or U17374 (N_17374,N_14572,N_14237);
and U17375 (N_17375,N_12574,N_12858);
xor U17376 (N_17376,N_15429,N_15032);
or U17377 (N_17377,N_13487,N_14437);
xor U17378 (N_17378,N_14576,N_14767);
nor U17379 (N_17379,N_12979,N_15087);
or U17380 (N_17380,N_13426,N_15000);
and U17381 (N_17381,N_13100,N_14693);
nor U17382 (N_17382,N_13859,N_14975);
nand U17383 (N_17383,N_14714,N_13024);
or U17384 (N_17384,N_14497,N_14449);
or U17385 (N_17385,N_13593,N_13628);
nor U17386 (N_17386,N_13436,N_13460);
or U17387 (N_17387,N_14826,N_12580);
and U17388 (N_17388,N_15503,N_13253);
and U17389 (N_17389,N_15123,N_13439);
nand U17390 (N_17390,N_14667,N_14916);
or U17391 (N_17391,N_15345,N_13574);
xor U17392 (N_17392,N_12642,N_15567);
nand U17393 (N_17393,N_14108,N_13504);
or U17394 (N_17394,N_14359,N_14822);
nand U17395 (N_17395,N_14311,N_13025);
xnor U17396 (N_17396,N_12679,N_14155);
or U17397 (N_17397,N_13990,N_13047);
or U17398 (N_17398,N_14477,N_12724);
xnor U17399 (N_17399,N_13783,N_12556);
nand U17400 (N_17400,N_14876,N_13539);
and U17401 (N_17401,N_12941,N_13551);
xor U17402 (N_17402,N_13858,N_13274);
or U17403 (N_17403,N_14015,N_14326);
and U17404 (N_17404,N_14475,N_15006);
and U17405 (N_17405,N_14709,N_14498);
nand U17406 (N_17406,N_14426,N_13851);
nand U17407 (N_17407,N_12603,N_14276);
or U17408 (N_17408,N_12723,N_14775);
nor U17409 (N_17409,N_15088,N_13838);
and U17410 (N_17410,N_15447,N_15467);
and U17411 (N_17411,N_12807,N_13365);
nand U17412 (N_17412,N_15513,N_15160);
and U17413 (N_17413,N_14613,N_13355);
xnor U17414 (N_17414,N_14860,N_14342);
and U17415 (N_17415,N_13954,N_14623);
nand U17416 (N_17416,N_14605,N_14608);
or U17417 (N_17417,N_14854,N_14872);
nand U17418 (N_17418,N_15607,N_13922);
nor U17419 (N_17419,N_13321,N_12906);
nor U17420 (N_17420,N_13104,N_14674);
nand U17421 (N_17421,N_15533,N_13605);
and U17422 (N_17422,N_14997,N_13940);
nor U17423 (N_17423,N_14536,N_14431);
or U17424 (N_17424,N_13801,N_13546);
or U17425 (N_17425,N_14695,N_15238);
nand U17426 (N_17426,N_12687,N_15619);
or U17427 (N_17427,N_12544,N_14527);
nor U17428 (N_17428,N_15031,N_14946);
and U17429 (N_17429,N_14664,N_12774);
nand U17430 (N_17430,N_15546,N_14748);
or U17431 (N_17431,N_13507,N_13719);
and U17432 (N_17432,N_13690,N_13124);
nand U17433 (N_17433,N_15098,N_12849);
and U17434 (N_17434,N_13702,N_14076);
and U17435 (N_17435,N_15280,N_14233);
or U17436 (N_17436,N_15276,N_13026);
nor U17437 (N_17437,N_15432,N_13025);
nand U17438 (N_17438,N_13419,N_14910);
and U17439 (N_17439,N_15586,N_14021);
nand U17440 (N_17440,N_14426,N_13006);
xor U17441 (N_17441,N_13644,N_15480);
xor U17442 (N_17442,N_14497,N_15597);
nor U17443 (N_17443,N_13201,N_14009);
or U17444 (N_17444,N_14906,N_13445);
nor U17445 (N_17445,N_12973,N_12862);
and U17446 (N_17446,N_13849,N_14462);
and U17447 (N_17447,N_14034,N_13835);
or U17448 (N_17448,N_14894,N_13446);
and U17449 (N_17449,N_13340,N_13073);
nor U17450 (N_17450,N_13773,N_14603);
nor U17451 (N_17451,N_13330,N_12740);
xnor U17452 (N_17452,N_14957,N_13020);
nand U17453 (N_17453,N_13583,N_14061);
nor U17454 (N_17454,N_13397,N_13068);
or U17455 (N_17455,N_12677,N_14920);
nor U17456 (N_17456,N_15316,N_14738);
or U17457 (N_17457,N_15059,N_13061);
and U17458 (N_17458,N_14246,N_12943);
or U17459 (N_17459,N_13359,N_13242);
and U17460 (N_17460,N_13629,N_13090);
nor U17461 (N_17461,N_12846,N_15181);
xor U17462 (N_17462,N_14399,N_12673);
or U17463 (N_17463,N_14407,N_15044);
nand U17464 (N_17464,N_13512,N_15559);
nand U17465 (N_17465,N_15308,N_15163);
nor U17466 (N_17466,N_12529,N_15513);
or U17467 (N_17467,N_12683,N_12946);
or U17468 (N_17468,N_12943,N_13045);
and U17469 (N_17469,N_13552,N_14518);
nand U17470 (N_17470,N_15302,N_14197);
nand U17471 (N_17471,N_12564,N_14434);
nor U17472 (N_17472,N_15574,N_13812);
nand U17473 (N_17473,N_12543,N_14218);
and U17474 (N_17474,N_13730,N_15045);
and U17475 (N_17475,N_14990,N_13084);
nand U17476 (N_17476,N_15535,N_15154);
or U17477 (N_17477,N_15348,N_13176);
or U17478 (N_17478,N_14359,N_14040);
or U17479 (N_17479,N_12697,N_13014);
xor U17480 (N_17480,N_14234,N_14866);
or U17481 (N_17481,N_13473,N_15383);
nor U17482 (N_17482,N_14339,N_13702);
xor U17483 (N_17483,N_13699,N_13853);
and U17484 (N_17484,N_13123,N_13163);
or U17485 (N_17485,N_15604,N_12960);
or U17486 (N_17486,N_14736,N_14768);
or U17487 (N_17487,N_13904,N_14012);
and U17488 (N_17488,N_15100,N_15105);
or U17489 (N_17489,N_13376,N_15055);
xor U17490 (N_17490,N_15510,N_13813);
and U17491 (N_17491,N_13867,N_13252);
nor U17492 (N_17492,N_12877,N_12682);
nor U17493 (N_17493,N_12611,N_14420);
and U17494 (N_17494,N_15339,N_15202);
or U17495 (N_17495,N_14498,N_15040);
and U17496 (N_17496,N_13880,N_15279);
xnor U17497 (N_17497,N_14787,N_13675);
nand U17498 (N_17498,N_12851,N_15384);
and U17499 (N_17499,N_15474,N_14766);
and U17500 (N_17500,N_15503,N_14050);
nor U17501 (N_17501,N_14863,N_13211);
or U17502 (N_17502,N_15136,N_12850);
nor U17503 (N_17503,N_14218,N_15456);
and U17504 (N_17504,N_13637,N_14342);
or U17505 (N_17505,N_13808,N_12627);
nor U17506 (N_17506,N_14399,N_14302);
xnor U17507 (N_17507,N_13622,N_13507);
nand U17508 (N_17508,N_12718,N_14975);
xnor U17509 (N_17509,N_14322,N_14422);
nand U17510 (N_17510,N_12992,N_12768);
and U17511 (N_17511,N_14459,N_13081);
nand U17512 (N_17512,N_14598,N_14609);
xnor U17513 (N_17513,N_14373,N_12539);
or U17514 (N_17514,N_13477,N_15159);
xnor U17515 (N_17515,N_13715,N_14510);
and U17516 (N_17516,N_13745,N_13075);
xnor U17517 (N_17517,N_13374,N_14915);
nand U17518 (N_17518,N_13604,N_15162);
or U17519 (N_17519,N_12809,N_12935);
and U17520 (N_17520,N_12638,N_13311);
or U17521 (N_17521,N_13464,N_15053);
xnor U17522 (N_17522,N_13070,N_15432);
xnor U17523 (N_17523,N_14885,N_14195);
nor U17524 (N_17524,N_14188,N_13279);
nand U17525 (N_17525,N_15155,N_12668);
xnor U17526 (N_17526,N_15385,N_13049);
xnor U17527 (N_17527,N_13665,N_14603);
or U17528 (N_17528,N_13418,N_15283);
or U17529 (N_17529,N_14889,N_15622);
nor U17530 (N_17530,N_13720,N_13002);
xor U17531 (N_17531,N_14194,N_14620);
nor U17532 (N_17532,N_12819,N_15150);
xor U17533 (N_17533,N_12601,N_14020);
nand U17534 (N_17534,N_15382,N_14991);
nand U17535 (N_17535,N_15139,N_15171);
nand U17536 (N_17536,N_15011,N_14680);
xor U17537 (N_17537,N_13411,N_12717);
nor U17538 (N_17538,N_15430,N_14754);
nand U17539 (N_17539,N_13130,N_15590);
and U17540 (N_17540,N_12619,N_13975);
or U17541 (N_17541,N_13163,N_13723);
or U17542 (N_17542,N_13039,N_13808);
xor U17543 (N_17543,N_13153,N_12733);
xnor U17544 (N_17544,N_15027,N_14505);
or U17545 (N_17545,N_15482,N_14892);
nand U17546 (N_17546,N_15349,N_14435);
xnor U17547 (N_17547,N_12950,N_13394);
or U17548 (N_17548,N_14271,N_12735);
and U17549 (N_17549,N_15598,N_13555);
and U17550 (N_17550,N_14250,N_12646);
nand U17551 (N_17551,N_14614,N_15419);
and U17552 (N_17552,N_13983,N_14883);
nand U17553 (N_17553,N_14170,N_13821);
nor U17554 (N_17554,N_14225,N_13523);
or U17555 (N_17555,N_14680,N_15544);
xor U17556 (N_17556,N_14908,N_13511);
xor U17557 (N_17557,N_14982,N_13767);
nand U17558 (N_17558,N_14910,N_13894);
xnor U17559 (N_17559,N_13865,N_15454);
nor U17560 (N_17560,N_12912,N_13967);
and U17561 (N_17561,N_14998,N_13564);
xnor U17562 (N_17562,N_15352,N_12757);
nor U17563 (N_17563,N_12569,N_13784);
xnor U17564 (N_17564,N_12556,N_15049);
and U17565 (N_17565,N_13888,N_13405);
and U17566 (N_17566,N_14912,N_12758);
nand U17567 (N_17567,N_14775,N_13023);
and U17568 (N_17568,N_13682,N_14349);
or U17569 (N_17569,N_14320,N_15518);
xnor U17570 (N_17570,N_15223,N_14515);
nor U17571 (N_17571,N_14554,N_13470);
and U17572 (N_17572,N_12930,N_13973);
and U17573 (N_17573,N_14999,N_12947);
nor U17574 (N_17574,N_15363,N_12930);
or U17575 (N_17575,N_12812,N_13886);
or U17576 (N_17576,N_13720,N_13026);
xnor U17577 (N_17577,N_15518,N_13077);
or U17578 (N_17578,N_14344,N_13051);
and U17579 (N_17579,N_14353,N_12599);
xnor U17580 (N_17580,N_12540,N_14029);
nand U17581 (N_17581,N_14416,N_13465);
or U17582 (N_17582,N_13607,N_15578);
or U17583 (N_17583,N_13208,N_13387);
xor U17584 (N_17584,N_15290,N_14683);
and U17585 (N_17585,N_15097,N_12708);
xor U17586 (N_17586,N_15383,N_15341);
nand U17587 (N_17587,N_12522,N_15069);
and U17588 (N_17588,N_15603,N_15489);
xnor U17589 (N_17589,N_15553,N_14072);
xor U17590 (N_17590,N_14594,N_13427);
and U17591 (N_17591,N_15623,N_13019);
and U17592 (N_17592,N_13758,N_12693);
xnor U17593 (N_17593,N_14237,N_14210);
and U17594 (N_17594,N_12942,N_13992);
nor U17595 (N_17595,N_13273,N_15522);
and U17596 (N_17596,N_15279,N_13483);
and U17597 (N_17597,N_14515,N_13335);
nand U17598 (N_17598,N_13376,N_14072);
or U17599 (N_17599,N_13942,N_13867);
and U17600 (N_17600,N_14868,N_12913);
nand U17601 (N_17601,N_15370,N_12650);
xnor U17602 (N_17602,N_15122,N_14202);
or U17603 (N_17603,N_13537,N_14304);
nor U17604 (N_17604,N_12994,N_12946);
nor U17605 (N_17605,N_13389,N_12787);
xnor U17606 (N_17606,N_14093,N_13879);
or U17607 (N_17607,N_12555,N_12988);
and U17608 (N_17608,N_15544,N_13835);
nand U17609 (N_17609,N_14155,N_13788);
xnor U17610 (N_17610,N_13501,N_12983);
xnor U17611 (N_17611,N_12717,N_14113);
nor U17612 (N_17612,N_14001,N_13831);
nand U17613 (N_17613,N_14809,N_13249);
nand U17614 (N_17614,N_12613,N_13116);
xnor U17615 (N_17615,N_12772,N_13041);
nor U17616 (N_17616,N_14603,N_15133);
nor U17617 (N_17617,N_13390,N_15497);
nand U17618 (N_17618,N_13388,N_14214);
nand U17619 (N_17619,N_15360,N_12775);
and U17620 (N_17620,N_13481,N_15446);
nor U17621 (N_17621,N_14889,N_13408);
xnor U17622 (N_17622,N_14290,N_14716);
or U17623 (N_17623,N_15074,N_14869);
nor U17624 (N_17624,N_14450,N_14682);
and U17625 (N_17625,N_14242,N_12711);
nor U17626 (N_17626,N_14090,N_14775);
nand U17627 (N_17627,N_13005,N_14033);
nor U17628 (N_17628,N_13541,N_13484);
nor U17629 (N_17629,N_12829,N_12731);
or U17630 (N_17630,N_14400,N_12830);
nor U17631 (N_17631,N_14271,N_15117);
or U17632 (N_17632,N_14781,N_14980);
or U17633 (N_17633,N_14462,N_15238);
xor U17634 (N_17634,N_14800,N_13675);
nand U17635 (N_17635,N_15083,N_14206);
and U17636 (N_17636,N_12545,N_12905);
and U17637 (N_17637,N_14471,N_13439);
xnor U17638 (N_17638,N_12670,N_14088);
nor U17639 (N_17639,N_14968,N_12556);
nor U17640 (N_17640,N_13670,N_14086);
nand U17641 (N_17641,N_14861,N_14139);
nor U17642 (N_17642,N_13552,N_15256);
nor U17643 (N_17643,N_12672,N_14395);
xor U17644 (N_17644,N_14714,N_15166);
nor U17645 (N_17645,N_13819,N_15119);
nor U17646 (N_17646,N_14377,N_14283);
nand U17647 (N_17647,N_13097,N_14919);
and U17648 (N_17648,N_13212,N_12657);
or U17649 (N_17649,N_15349,N_14145);
or U17650 (N_17650,N_13019,N_15184);
and U17651 (N_17651,N_15158,N_14056);
xnor U17652 (N_17652,N_14183,N_15222);
and U17653 (N_17653,N_15198,N_15489);
nor U17654 (N_17654,N_14856,N_14212);
nor U17655 (N_17655,N_14936,N_14415);
and U17656 (N_17656,N_12525,N_13496);
nand U17657 (N_17657,N_15358,N_15615);
nor U17658 (N_17658,N_15578,N_13340);
nand U17659 (N_17659,N_13138,N_13272);
or U17660 (N_17660,N_15275,N_15247);
xor U17661 (N_17661,N_14569,N_15214);
and U17662 (N_17662,N_13490,N_15502);
xnor U17663 (N_17663,N_14369,N_14778);
nor U17664 (N_17664,N_13093,N_14599);
or U17665 (N_17665,N_13659,N_12842);
and U17666 (N_17666,N_13230,N_12665);
nand U17667 (N_17667,N_13032,N_15385);
nand U17668 (N_17668,N_15129,N_15353);
nand U17669 (N_17669,N_14003,N_13844);
xnor U17670 (N_17670,N_13375,N_13622);
xnor U17671 (N_17671,N_14768,N_13952);
xnor U17672 (N_17672,N_14165,N_13884);
and U17673 (N_17673,N_14664,N_13210);
xnor U17674 (N_17674,N_13362,N_14913);
or U17675 (N_17675,N_15025,N_12978);
nor U17676 (N_17676,N_15383,N_15158);
or U17677 (N_17677,N_14820,N_13550);
nor U17678 (N_17678,N_13429,N_12920);
and U17679 (N_17679,N_13964,N_12581);
or U17680 (N_17680,N_14787,N_14161);
nand U17681 (N_17681,N_14218,N_14393);
xnor U17682 (N_17682,N_13038,N_13773);
nand U17683 (N_17683,N_13495,N_12768);
or U17684 (N_17684,N_14940,N_12740);
xnor U17685 (N_17685,N_15617,N_14877);
and U17686 (N_17686,N_14449,N_12922);
nand U17687 (N_17687,N_14579,N_14997);
nand U17688 (N_17688,N_13328,N_14997);
and U17689 (N_17689,N_12515,N_14844);
and U17690 (N_17690,N_13968,N_12993);
xor U17691 (N_17691,N_12528,N_13518);
and U17692 (N_17692,N_14698,N_12597);
or U17693 (N_17693,N_13574,N_15355);
or U17694 (N_17694,N_13978,N_13141);
and U17695 (N_17695,N_14721,N_15389);
and U17696 (N_17696,N_14895,N_15157);
nor U17697 (N_17697,N_15020,N_14149);
nor U17698 (N_17698,N_14244,N_12530);
nand U17699 (N_17699,N_15481,N_15499);
xor U17700 (N_17700,N_12671,N_14464);
nor U17701 (N_17701,N_14306,N_13974);
xor U17702 (N_17702,N_14298,N_14602);
nor U17703 (N_17703,N_13671,N_14089);
nor U17704 (N_17704,N_13486,N_15312);
and U17705 (N_17705,N_14850,N_15370);
and U17706 (N_17706,N_12711,N_14794);
and U17707 (N_17707,N_13686,N_13833);
xor U17708 (N_17708,N_14349,N_13450);
nand U17709 (N_17709,N_14906,N_13603);
or U17710 (N_17710,N_12865,N_15176);
and U17711 (N_17711,N_14557,N_14386);
xor U17712 (N_17712,N_14586,N_13754);
or U17713 (N_17713,N_12840,N_14506);
nand U17714 (N_17714,N_13115,N_12520);
or U17715 (N_17715,N_12924,N_13454);
nor U17716 (N_17716,N_13852,N_13815);
nor U17717 (N_17717,N_13762,N_12938);
nand U17718 (N_17718,N_13006,N_13875);
xor U17719 (N_17719,N_12624,N_15383);
or U17720 (N_17720,N_14535,N_13702);
xnor U17721 (N_17721,N_15038,N_13723);
and U17722 (N_17722,N_13881,N_13723);
nor U17723 (N_17723,N_15624,N_12827);
and U17724 (N_17724,N_14427,N_13795);
nor U17725 (N_17725,N_13272,N_14384);
or U17726 (N_17726,N_13225,N_12544);
xnor U17727 (N_17727,N_13121,N_12699);
nand U17728 (N_17728,N_12935,N_12783);
or U17729 (N_17729,N_13831,N_13392);
xnor U17730 (N_17730,N_15569,N_13894);
and U17731 (N_17731,N_15530,N_14195);
nor U17732 (N_17732,N_14687,N_14426);
xnor U17733 (N_17733,N_14074,N_15061);
xnor U17734 (N_17734,N_13890,N_14845);
nand U17735 (N_17735,N_14276,N_14531);
or U17736 (N_17736,N_13499,N_14101);
and U17737 (N_17737,N_15201,N_13169);
nand U17738 (N_17738,N_14850,N_13972);
or U17739 (N_17739,N_15094,N_13667);
xnor U17740 (N_17740,N_14353,N_14459);
and U17741 (N_17741,N_14714,N_12587);
nor U17742 (N_17742,N_14801,N_12555);
xor U17743 (N_17743,N_12865,N_13525);
nor U17744 (N_17744,N_15089,N_14826);
nand U17745 (N_17745,N_15349,N_15520);
nor U17746 (N_17746,N_15525,N_14604);
nor U17747 (N_17747,N_15199,N_13009);
nand U17748 (N_17748,N_13840,N_15042);
and U17749 (N_17749,N_12762,N_14138);
nor U17750 (N_17750,N_14342,N_13049);
or U17751 (N_17751,N_15530,N_15328);
xor U17752 (N_17752,N_12924,N_14536);
xor U17753 (N_17753,N_14813,N_14073);
or U17754 (N_17754,N_13174,N_15436);
or U17755 (N_17755,N_14273,N_13712);
nor U17756 (N_17756,N_13852,N_13732);
and U17757 (N_17757,N_13386,N_13646);
or U17758 (N_17758,N_13277,N_14596);
nand U17759 (N_17759,N_12588,N_13514);
xnor U17760 (N_17760,N_14731,N_13466);
or U17761 (N_17761,N_13433,N_12878);
nand U17762 (N_17762,N_12677,N_12768);
nand U17763 (N_17763,N_14044,N_14293);
nor U17764 (N_17764,N_12525,N_12697);
or U17765 (N_17765,N_15443,N_12927);
nor U17766 (N_17766,N_14462,N_12852);
and U17767 (N_17767,N_12538,N_15555);
xor U17768 (N_17768,N_12509,N_13090);
nand U17769 (N_17769,N_13027,N_14246);
xor U17770 (N_17770,N_13170,N_13063);
nand U17771 (N_17771,N_15387,N_14163);
nor U17772 (N_17772,N_13492,N_13607);
nor U17773 (N_17773,N_15271,N_15549);
or U17774 (N_17774,N_14981,N_14275);
nand U17775 (N_17775,N_12960,N_13668);
nand U17776 (N_17776,N_15490,N_15576);
or U17777 (N_17777,N_14297,N_15208);
nand U17778 (N_17778,N_14744,N_14605);
and U17779 (N_17779,N_14849,N_15049);
nand U17780 (N_17780,N_15566,N_13251);
xor U17781 (N_17781,N_12696,N_14785);
nand U17782 (N_17782,N_14080,N_14038);
or U17783 (N_17783,N_13435,N_13115);
nand U17784 (N_17784,N_14736,N_13820);
or U17785 (N_17785,N_13850,N_12791);
xnor U17786 (N_17786,N_15335,N_15172);
nand U17787 (N_17787,N_14047,N_15331);
nand U17788 (N_17788,N_13401,N_13075);
nor U17789 (N_17789,N_14068,N_13982);
and U17790 (N_17790,N_12951,N_14638);
nor U17791 (N_17791,N_14986,N_13438);
and U17792 (N_17792,N_15204,N_13652);
xor U17793 (N_17793,N_13435,N_13355);
nor U17794 (N_17794,N_14644,N_12509);
nand U17795 (N_17795,N_14355,N_13448);
nor U17796 (N_17796,N_13092,N_12623);
nand U17797 (N_17797,N_12632,N_13775);
nand U17798 (N_17798,N_12782,N_14099);
nand U17799 (N_17799,N_14957,N_15182);
nand U17800 (N_17800,N_14685,N_15589);
xor U17801 (N_17801,N_13013,N_13384);
and U17802 (N_17802,N_15286,N_14933);
and U17803 (N_17803,N_15335,N_15510);
or U17804 (N_17804,N_13421,N_14726);
nand U17805 (N_17805,N_15174,N_14282);
or U17806 (N_17806,N_14253,N_13180);
or U17807 (N_17807,N_12814,N_12999);
nor U17808 (N_17808,N_13642,N_13452);
or U17809 (N_17809,N_13677,N_14926);
nand U17810 (N_17810,N_14457,N_14426);
nor U17811 (N_17811,N_14309,N_12891);
or U17812 (N_17812,N_13459,N_14279);
or U17813 (N_17813,N_14656,N_14152);
and U17814 (N_17814,N_12732,N_15221);
xnor U17815 (N_17815,N_14215,N_14627);
or U17816 (N_17816,N_14859,N_14535);
nor U17817 (N_17817,N_15061,N_15157);
and U17818 (N_17818,N_13575,N_14668);
or U17819 (N_17819,N_13574,N_14550);
nor U17820 (N_17820,N_12944,N_14636);
xor U17821 (N_17821,N_15214,N_15437);
nor U17822 (N_17822,N_13657,N_14919);
and U17823 (N_17823,N_15529,N_15204);
or U17824 (N_17824,N_13077,N_15612);
xor U17825 (N_17825,N_14868,N_13094);
nand U17826 (N_17826,N_13097,N_13181);
nor U17827 (N_17827,N_12500,N_14057);
nor U17828 (N_17828,N_14964,N_14706);
or U17829 (N_17829,N_13542,N_13318);
xnor U17830 (N_17830,N_14452,N_12805);
xor U17831 (N_17831,N_12524,N_12606);
or U17832 (N_17832,N_13662,N_14209);
or U17833 (N_17833,N_14650,N_13356);
xnor U17834 (N_17834,N_15241,N_12677);
nand U17835 (N_17835,N_12909,N_14457);
and U17836 (N_17836,N_14667,N_15560);
nor U17837 (N_17837,N_15524,N_13066);
and U17838 (N_17838,N_12936,N_12525);
xor U17839 (N_17839,N_13572,N_15595);
or U17840 (N_17840,N_13430,N_14397);
nor U17841 (N_17841,N_12670,N_14310);
and U17842 (N_17842,N_13187,N_14662);
xor U17843 (N_17843,N_14565,N_13241);
xor U17844 (N_17844,N_12537,N_13877);
nor U17845 (N_17845,N_13030,N_13934);
nor U17846 (N_17846,N_14615,N_12707);
and U17847 (N_17847,N_15068,N_12995);
nor U17848 (N_17848,N_12686,N_14276);
nor U17849 (N_17849,N_12789,N_13500);
nor U17850 (N_17850,N_14605,N_14808);
nand U17851 (N_17851,N_15151,N_13183);
nand U17852 (N_17852,N_13547,N_15375);
nor U17853 (N_17853,N_13595,N_14479);
nand U17854 (N_17854,N_14662,N_14513);
nand U17855 (N_17855,N_12921,N_14607);
and U17856 (N_17856,N_13500,N_13003);
and U17857 (N_17857,N_12845,N_14096);
and U17858 (N_17858,N_13202,N_12698);
nor U17859 (N_17859,N_15358,N_13500);
or U17860 (N_17860,N_15020,N_14288);
and U17861 (N_17861,N_14820,N_12634);
xnor U17862 (N_17862,N_12779,N_14399);
or U17863 (N_17863,N_12518,N_13484);
or U17864 (N_17864,N_12994,N_15541);
or U17865 (N_17865,N_14576,N_13612);
or U17866 (N_17866,N_13957,N_14267);
nor U17867 (N_17867,N_13749,N_14316);
nand U17868 (N_17868,N_13250,N_13991);
nand U17869 (N_17869,N_12973,N_12861);
or U17870 (N_17870,N_15150,N_13213);
and U17871 (N_17871,N_15028,N_15222);
nand U17872 (N_17872,N_14763,N_14594);
nor U17873 (N_17873,N_12832,N_13835);
and U17874 (N_17874,N_15052,N_13448);
or U17875 (N_17875,N_12693,N_15000);
and U17876 (N_17876,N_15148,N_14099);
or U17877 (N_17877,N_13232,N_13342);
and U17878 (N_17878,N_12870,N_14522);
xor U17879 (N_17879,N_13024,N_12838);
and U17880 (N_17880,N_13162,N_14016);
nor U17881 (N_17881,N_13261,N_13701);
or U17882 (N_17882,N_12643,N_13729);
nand U17883 (N_17883,N_13475,N_13199);
or U17884 (N_17884,N_13231,N_15387);
nor U17885 (N_17885,N_13670,N_15494);
xor U17886 (N_17886,N_14517,N_15116);
and U17887 (N_17887,N_15204,N_12658);
nand U17888 (N_17888,N_14584,N_15035);
nand U17889 (N_17889,N_13227,N_14525);
and U17890 (N_17890,N_12586,N_13545);
and U17891 (N_17891,N_13831,N_14268);
and U17892 (N_17892,N_13182,N_14681);
xor U17893 (N_17893,N_14504,N_14060);
nand U17894 (N_17894,N_15125,N_13384);
nand U17895 (N_17895,N_12711,N_13944);
or U17896 (N_17896,N_13353,N_12833);
nor U17897 (N_17897,N_15300,N_12679);
nand U17898 (N_17898,N_13288,N_14810);
xnor U17899 (N_17899,N_14419,N_12787);
and U17900 (N_17900,N_14160,N_13588);
and U17901 (N_17901,N_14157,N_14774);
and U17902 (N_17902,N_13391,N_12678);
xnor U17903 (N_17903,N_14501,N_13541);
or U17904 (N_17904,N_15402,N_13499);
and U17905 (N_17905,N_12718,N_13393);
nand U17906 (N_17906,N_14398,N_15603);
xor U17907 (N_17907,N_13708,N_15176);
nand U17908 (N_17908,N_14914,N_13779);
nor U17909 (N_17909,N_12883,N_14559);
or U17910 (N_17910,N_14586,N_13585);
xor U17911 (N_17911,N_12823,N_12795);
or U17912 (N_17912,N_13025,N_12642);
nor U17913 (N_17913,N_13705,N_13948);
nor U17914 (N_17914,N_14459,N_14532);
or U17915 (N_17915,N_13488,N_12527);
nor U17916 (N_17916,N_14532,N_15533);
nor U17917 (N_17917,N_15467,N_14030);
xor U17918 (N_17918,N_12580,N_15122);
or U17919 (N_17919,N_14480,N_12721);
nor U17920 (N_17920,N_12625,N_15611);
xor U17921 (N_17921,N_12693,N_12704);
nor U17922 (N_17922,N_14266,N_15383);
nor U17923 (N_17923,N_13407,N_13195);
xor U17924 (N_17924,N_14252,N_14036);
xor U17925 (N_17925,N_14435,N_14656);
and U17926 (N_17926,N_13740,N_15318);
xnor U17927 (N_17927,N_15548,N_15189);
nor U17928 (N_17928,N_13270,N_13289);
nor U17929 (N_17929,N_15485,N_15177);
and U17930 (N_17930,N_14600,N_14854);
and U17931 (N_17931,N_13321,N_12843);
nand U17932 (N_17932,N_14739,N_13982);
and U17933 (N_17933,N_13921,N_13791);
and U17934 (N_17934,N_14619,N_15465);
or U17935 (N_17935,N_14803,N_14018);
and U17936 (N_17936,N_13431,N_12654);
nor U17937 (N_17937,N_12568,N_15224);
nand U17938 (N_17938,N_13874,N_15427);
xor U17939 (N_17939,N_14293,N_13477);
nor U17940 (N_17940,N_12999,N_14773);
xor U17941 (N_17941,N_13881,N_15067);
and U17942 (N_17942,N_15011,N_13427);
or U17943 (N_17943,N_15471,N_13612);
or U17944 (N_17944,N_14194,N_13026);
and U17945 (N_17945,N_15552,N_12585);
nand U17946 (N_17946,N_12586,N_13032);
or U17947 (N_17947,N_15062,N_14418);
xnor U17948 (N_17948,N_15208,N_13049);
nor U17949 (N_17949,N_15582,N_13422);
nand U17950 (N_17950,N_14051,N_13999);
and U17951 (N_17951,N_14191,N_14105);
nor U17952 (N_17952,N_13700,N_15536);
or U17953 (N_17953,N_14124,N_15608);
and U17954 (N_17954,N_12566,N_14672);
nand U17955 (N_17955,N_13956,N_13880);
and U17956 (N_17956,N_13256,N_13701);
xnor U17957 (N_17957,N_13948,N_13795);
or U17958 (N_17958,N_14005,N_12579);
nor U17959 (N_17959,N_14869,N_14971);
nor U17960 (N_17960,N_13222,N_13103);
nor U17961 (N_17961,N_14108,N_14385);
or U17962 (N_17962,N_14408,N_14992);
xnor U17963 (N_17963,N_14965,N_12824);
nor U17964 (N_17964,N_14128,N_14661);
and U17965 (N_17965,N_14381,N_14405);
nor U17966 (N_17966,N_14098,N_13970);
xnor U17967 (N_17967,N_14812,N_15104);
or U17968 (N_17968,N_15561,N_14332);
nand U17969 (N_17969,N_14968,N_13424);
xor U17970 (N_17970,N_14833,N_15296);
and U17971 (N_17971,N_14571,N_12723);
or U17972 (N_17972,N_15422,N_13579);
and U17973 (N_17973,N_15527,N_15585);
or U17974 (N_17974,N_14035,N_15538);
or U17975 (N_17975,N_14935,N_15592);
and U17976 (N_17976,N_12976,N_14769);
nor U17977 (N_17977,N_13201,N_15110);
nor U17978 (N_17978,N_14281,N_14566);
or U17979 (N_17979,N_15230,N_15420);
nor U17980 (N_17980,N_12984,N_12732);
nor U17981 (N_17981,N_12900,N_15279);
nand U17982 (N_17982,N_12566,N_15021);
nor U17983 (N_17983,N_15359,N_12715);
nor U17984 (N_17984,N_14253,N_14268);
or U17985 (N_17985,N_13571,N_14340);
and U17986 (N_17986,N_15234,N_15144);
nand U17987 (N_17987,N_14515,N_13735);
and U17988 (N_17988,N_14777,N_13546);
xor U17989 (N_17989,N_12901,N_15342);
or U17990 (N_17990,N_13236,N_14434);
nand U17991 (N_17991,N_15140,N_12819);
nand U17992 (N_17992,N_14055,N_12929);
and U17993 (N_17993,N_13031,N_14553);
or U17994 (N_17994,N_15127,N_13014);
nor U17995 (N_17995,N_14560,N_13804);
xor U17996 (N_17996,N_13113,N_13930);
xor U17997 (N_17997,N_14870,N_15064);
xnor U17998 (N_17998,N_13646,N_13856);
nand U17999 (N_17999,N_15411,N_13435);
nand U18000 (N_18000,N_12736,N_14092);
nor U18001 (N_18001,N_13430,N_14241);
nor U18002 (N_18002,N_12920,N_14618);
xnor U18003 (N_18003,N_15223,N_12984);
nor U18004 (N_18004,N_14870,N_12755);
and U18005 (N_18005,N_14110,N_13082);
and U18006 (N_18006,N_14300,N_14549);
and U18007 (N_18007,N_12799,N_12571);
and U18008 (N_18008,N_12559,N_15511);
nor U18009 (N_18009,N_12629,N_13598);
and U18010 (N_18010,N_14004,N_13181);
or U18011 (N_18011,N_13202,N_12686);
or U18012 (N_18012,N_14160,N_14271);
nand U18013 (N_18013,N_12771,N_13652);
nor U18014 (N_18014,N_13945,N_13805);
nor U18015 (N_18015,N_13437,N_14123);
nor U18016 (N_18016,N_15201,N_15004);
nor U18017 (N_18017,N_13862,N_15557);
nor U18018 (N_18018,N_14093,N_14416);
or U18019 (N_18019,N_14260,N_14436);
nand U18020 (N_18020,N_13177,N_14017);
nand U18021 (N_18021,N_14585,N_15090);
nor U18022 (N_18022,N_12767,N_13868);
nor U18023 (N_18023,N_15551,N_14537);
or U18024 (N_18024,N_13959,N_12995);
or U18025 (N_18025,N_13595,N_12852);
nor U18026 (N_18026,N_13146,N_13598);
and U18027 (N_18027,N_15574,N_15055);
nor U18028 (N_18028,N_14190,N_12914);
nand U18029 (N_18029,N_13643,N_15406);
nor U18030 (N_18030,N_12572,N_14592);
nor U18031 (N_18031,N_14517,N_13403);
xor U18032 (N_18032,N_12565,N_12996);
or U18033 (N_18033,N_14294,N_15535);
nor U18034 (N_18034,N_12940,N_15475);
or U18035 (N_18035,N_15292,N_15479);
nor U18036 (N_18036,N_13993,N_14217);
nor U18037 (N_18037,N_13203,N_13435);
nand U18038 (N_18038,N_15332,N_13566);
xor U18039 (N_18039,N_15038,N_14796);
and U18040 (N_18040,N_12989,N_15505);
nor U18041 (N_18041,N_12778,N_12692);
xnor U18042 (N_18042,N_13445,N_14811);
nand U18043 (N_18043,N_12654,N_12566);
xnor U18044 (N_18044,N_15088,N_15577);
nand U18045 (N_18045,N_15037,N_13974);
or U18046 (N_18046,N_15456,N_14442);
nand U18047 (N_18047,N_14537,N_13505);
or U18048 (N_18048,N_14944,N_14664);
nor U18049 (N_18049,N_14646,N_15359);
or U18050 (N_18050,N_15601,N_14384);
or U18051 (N_18051,N_14939,N_13046);
and U18052 (N_18052,N_13296,N_13532);
xnor U18053 (N_18053,N_14056,N_14959);
nand U18054 (N_18054,N_12641,N_13340);
and U18055 (N_18055,N_13978,N_15266);
xor U18056 (N_18056,N_12719,N_12949);
nor U18057 (N_18057,N_12845,N_13857);
nand U18058 (N_18058,N_14755,N_15623);
xor U18059 (N_18059,N_15153,N_14909);
xnor U18060 (N_18060,N_15009,N_14070);
and U18061 (N_18061,N_12963,N_15096);
nand U18062 (N_18062,N_15345,N_13418);
xor U18063 (N_18063,N_14675,N_13237);
xnor U18064 (N_18064,N_12834,N_15253);
nand U18065 (N_18065,N_15157,N_14873);
nand U18066 (N_18066,N_14629,N_14326);
or U18067 (N_18067,N_13652,N_13034);
and U18068 (N_18068,N_13825,N_12775);
or U18069 (N_18069,N_13055,N_12691);
and U18070 (N_18070,N_15623,N_12527);
xnor U18071 (N_18071,N_15438,N_12879);
and U18072 (N_18072,N_14545,N_12698);
or U18073 (N_18073,N_13495,N_15482);
or U18074 (N_18074,N_14835,N_14232);
xnor U18075 (N_18075,N_13947,N_13931);
nand U18076 (N_18076,N_14913,N_12822);
and U18077 (N_18077,N_14598,N_12734);
and U18078 (N_18078,N_15404,N_12989);
nor U18079 (N_18079,N_13585,N_14864);
xnor U18080 (N_18080,N_13459,N_14133);
xnor U18081 (N_18081,N_13410,N_12714);
nand U18082 (N_18082,N_13819,N_15331);
or U18083 (N_18083,N_13860,N_15213);
xor U18084 (N_18084,N_13593,N_13552);
or U18085 (N_18085,N_12879,N_15238);
nand U18086 (N_18086,N_13178,N_12877);
and U18087 (N_18087,N_15287,N_12901);
or U18088 (N_18088,N_13124,N_12647);
nor U18089 (N_18089,N_15254,N_12796);
or U18090 (N_18090,N_13220,N_13924);
nor U18091 (N_18091,N_13845,N_14793);
nor U18092 (N_18092,N_14080,N_12630);
nor U18093 (N_18093,N_13785,N_15005);
nor U18094 (N_18094,N_13272,N_14436);
xor U18095 (N_18095,N_14612,N_13144);
nand U18096 (N_18096,N_15007,N_13534);
nand U18097 (N_18097,N_14299,N_13398);
and U18098 (N_18098,N_13531,N_15590);
nor U18099 (N_18099,N_14961,N_15351);
nand U18100 (N_18100,N_15141,N_14030);
nand U18101 (N_18101,N_14766,N_12967);
nand U18102 (N_18102,N_13255,N_14974);
or U18103 (N_18103,N_14751,N_13587);
nor U18104 (N_18104,N_12748,N_13123);
or U18105 (N_18105,N_15317,N_12878);
xnor U18106 (N_18106,N_13477,N_14216);
xor U18107 (N_18107,N_13870,N_15070);
or U18108 (N_18108,N_12743,N_13860);
or U18109 (N_18109,N_15249,N_14410);
or U18110 (N_18110,N_12718,N_13150);
and U18111 (N_18111,N_14887,N_14833);
nand U18112 (N_18112,N_13139,N_15159);
nor U18113 (N_18113,N_13789,N_12814);
nor U18114 (N_18114,N_12711,N_13620);
nor U18115 (N_18115,N_12568,N_15570);
nand U18116 (N_18116,N_15156,N_13852);
or U18117 (N_18117,N_14891,N_12650);
xor U18118 (N_18118,N_13660,N_13362);
nor U18119 (N_18119,N_13120,N_14234);
nand U18120 (N_18120,N_13781,N_14090);
and U18121 (N_18121,N_13215,N_14555);
and U18122 (N_18122,N_12685,N_13888);
xor U18123 (N_18123,N_12624,N_13606);
nand U18124 (N_18124,N_13036,N_15346);
nand U18125 (N_18125,N_14778,N_15156);
and U18126 (N_18126,N_14102,N_13603);
xor U18127 (N_18127,N_13070,N_13935);
nor U18128 (N_18128,N_12563,N_13736);
nand U18129 (N_18129,N_14819,N_12748);
xnor U18130 (N_18130,N_15303,N_12645);
nand U18131 (N_18131,N_13555,N_13214);
or U18132 (N_18132,N_14060,N_13515);
or U18133 (N_18133,N_15613,N_14568);
or U18134 (N_18134,N_14486,N_13907);
nor U18135 (N_18135,N_15448,N_13076);
or U18136 (N_18136,N_14478,N_15492);
or U18137 (N_18137,N_12863,N_14420);
or U18138 (N_18138,N_14556,N_14686);
or U18139 (N_18139,N_12657,N_14684);
nand U18140 (N_18140,N_13869,N_14422);
and U18141 (N_18141,N_14036,N_13275);
and U18142 (N_18142,N_14050,N_14255);
xnor U18143 (N_18143,N_13159,N_15188);
xnor U18144 (N_18144,N_12657,N_13546);
and U18145 (N_18145,N_14489,N_15376);
nand U18146 (N_18146,N_13312,N_14242);
nand U18147 (N_18147,N_15332,N_13311);
or U18148 (N_18148,N_14892,N_13531);
nand U18149 (N_18149,N_14491,N_14060);
nand U18150 (N_18150,N_13924,N_15467);
nand U18151 (N_18151,N_13571,N_13148);
nand U18152 (N_18152,N_14566,N_14013);
xnor U18153 (N_18153,N_15420,N_13243);
or U18154 (N_18154,N_14860,N_12500);
nand U18155 (N_18155,N_14274,N_13691);
nor U18156 (N_18156,N_14966,N_13397);
or U18157 (N_18157,N_15150,N_13461);
or U18158 (N_18158,N_14517,N_14518);
and U18159 (N_18159,N_13545,N_14369);
nand U18160 (N_18160,N_13974,N_14718);
xnor U18161 (N_18161,N_13534,N_13219);
nor U18162 (N_18162,N_13606,N_15401);
xor U18163 (N_18163,N_14645,N_13595);
xnor U18164 (N_18164,N_13727,N_14667);
or U18165 (N_18165,N_15498,N_14442);
nor U18166 (N_18166,N_13847,N_12939);
nand U18167 (N_18167,N_12977,N_12944);
or U18168 (N_18168,N_14359,N_12843);
nor U18169 (N_18169,N_14714,N_15061);
and U18170 (N_18170,N_15303,N_13242);
nand U18171 (N_18171,N_14869,N_15312);
or U18172 (N_18172,N_14720,N_13577);
or U18173 (N_18173,N_13008,N_12870);
nand U18174 (N_18174,N_12577,N_12831);
nand U18175 (N_18175,N_13112,N_14006);
nand U18176 (N_18176,N_12571,N_13157);
or U18177 (N_18177,N_15265,N_15139);
xor U18178 (N_18178,N_15101,N_12567);
or U18179 (N_18179,N_14796,N_14241);
or U18180 (N_18180,N_13536,N_12735);
xnor U18181 (N_18181,N_14482,N_15566);
nor U18182 (N_18182,N_14080,N_15208);
or U18183 (N_18183,N_15325,N_13042);
xnor U18184 (N_18184,N_12572,N_13721);
and U18185 (N_18185,N_13729,N_14777);
nor U18186 (N_18186,N_14135,N_12888);
or U18187 (N_18187,N_15576,N_13512);
nor U18188 (N_18188,N_14704,N_14993);
nor U18189 (N_18189,N_15196,N_15496);
nand U18190 (N_18190,N_12726,N_12756);
and U18191 (N_18191,N_14415,N_14255);
and U18192 (N_18192,N_14252,N_14046);
nor U18193 (N_18193,N_13304,N_12551);
and U18194 (N_18194,N_12592,N_14235);
xnor U18195 (N_18195,N_12580,N_15116);
and U18196 (N_18196,N_12687,N_15184);
xor U18197 (N_18197,N_14178,N_13854);
nor U18198 (N_18198,N_14590,N_13678);
and U18199 (N_18199,N_13101,N_14783);
xnor U18200 (N_18200,N_13344,N_13548);
and U18201 (N_18201,N_12827,N_13804);
and U18202 (N_18202,N_15147,N_13168);
xor U18203 (N_18203,N_15261,N_14862);
nor U18204 (N_18204,N_13565,N_12825);
nor U18205 (N_18205,N_14317,N_13362);
or U18206 (N_18206,N_14999,N_12761);
nand U18207 (N_18207,N_13377,N_13944);
nor U18208 (N_18208,N_15244,N_13018);
nor U18209 (N_18209,N_12685,N_15620);
nor U18210 (N_18210,N_14697,N_14096);
nor U18211 (N_18211,N_13691,N_12639);
nor U18212 (N_18212,N_13542,N_14109);
and U18213 (N_18213,N_14151,N_13992);
or U18214 (N_18214,N_12653,N_13792);
nand U18215 (N_18215,N_13888,N_13587);
nor U18216 (N_18216,N_13887,N_12618);
nor U18217 (N_18217,N_14920,N_14603);
xor U18218 (N_18218,N_13886,N_15041);
nand U18219 (N_18219,N_13216,N_14342);
nor U18220 (N_18220,N_12682,N_14496);
and U18221 (N_18221,N_13989,N_14181);
or U18222 (N_18222,N_14955,N_13510);
nor U18223 (N_18223,N_15481,N_13515);
nand U18224 (N_18224,N_14108,N_13030);
and U18225 (N_18225,N_12806,N_12724);
xnor U18226 (N_18226,N_14990,N_14255);
nor U18227 (N_18227,N_14102,N_13473);
xnor U18228 (N_18228,N_14870,N_13322);
nand U18229 (N_18229,N_15042,N_15616);
or U18230 (N_18230,N_14742,N_13589);
and U18231 (N_18231,N_13382,N_14244);
or U18232 (N_18232,N_13572,N_13995);
nor U18233 (N_18233,N_13927,N_15418);
or U18234 (N_18234,N_13297,N_13658);
and U18235 (N_18235,N_13693,N_13275);
and U18236 (N_18236,N_13446,N_15144);
nor U18237 (N_18237,N_15334,N_13084);
and U18238 (N_18238,N_13064,N_13296);
and U18239 (N_18239,N_15261,N_13719);
and U18240 (N_18240,N_13309,N_13795);
or U18241 (N_18241,N_15434,N_13418);
xnor U18242 (N_18242,N_12998,N_13573);
or U18243 (N_18243,N_14106,N_12726);
and U18244 (N_18244,N_14097,N_12979);
nand U18245 (N_18245,N_13010,N_14404);
and U18246 (N_18246,N_14638,N_14735);
and U18247 (N_18247,N_14941,N_12693);
nor U18248 (N_18248,N_14239,N_13026);
xnor U18249 (N_18249,N_13243,N_13110);
xnor U18250 (N_18250,N_14129,N_15623);
nor U18251 (N_18251,N_12690,N_14700);
and U18252 (N_18252,N_14245,N_13467);
or U18253 (N_18253,N_12769,N_15323);
and U18254 (N_18254,N_12921,N_12784);
nor U18255 (N_18255,N_14121,N_13176);
or U18256 (N_18256,N_15176,N_15130);
or U18257 (N_18257,N_13501,N_14605);
nor U18258 (N_18258,N_13627,N_12927);
nand U18259 (N_18259,N_15578,N_14960);
xnor U18260 (N_18260,N_14174,N_14018);
nand U18261 (N_18261,N_14166,N_13212);
nor U18262 (N_18262,N_12689,N_14959);
or U18263 (N_18263,N_13796,N_15288);
and U18264 (N_18264,N_14457,N_15402);
and U18265 (N_18265,N_15484,N_13741);
or U18266 (N_18266,N_13155,N_15583);
nor U18267 (N_18267,N_14937,N_14981);
or U18268 (N_18268,N_13794,N_13408);
xor U18269 (N_18269,N_12811,N_14826);
or U18270 (N_18270,N_15600,N_15003);
or U18271 (N_18271,N_15022,N_13748);
nand U18272 (N_18272,N_13157,N_14191);
xor U18273 (N_18273,N_13472,N_15175);
xnor U18274 (N_18274,N_14163,N_14750);
and U18275 (N_18275,N_15258,N_14902);
nand U18276 (N_18276,N_13745,N_14714);
and U18277 (N_18277,N_14042,N_14353);
or U18278 (N_18278,N_12871,N_14435);
nand U18279 (N_18279,N_14751,N_13394);
and U18280 (N_18280,N_14888,N_15448);
or U18281 (N_18281,N_12696,N_13707);
or U18282 (N_18282,N_13456,N_15453);
nor U18283 (N_18283,N_15589,N_13393);
nor U18284 (N_18284,N_14254,N_14698);
and U18285 (N_18285,N_14697,N_13936);
nor U18286 (N_18286,N_13881,N_13927);
nor U18287 (N_18287,N_12925,N_14680);
or U18288 (N_18288,N_13064,N_14250);
nor U18289 (N_18289,N_15418,N_15279);
or U18290 (N_18290,N_14786,N_14972);
and U18291 (N_18291,N_13345,N_14960);
nor U18292 (N_18292,N_12959,N_13666);
or U18293 (N_18293,N_12562,N_13558);
and U18294 (N_18294,N_13144,N_13335);
nor U18295 (N_18295,N_14898,N_14934);
and U18296 (N_18296,N_13234,N_13562);
or U18297 (N_18297,N_12887,N_14054);
xor U18298 (N_18298,N_12629,N_15369);
xnor U18299 (N_18299,N_13757,N_13058);
nor U18300 (N_18300,N_12637,N_14216);
xor U18301 (N_18301,N_13398,N_14556);
xor U18302 (N_18302,N_13108,N_13358);
xnor U18303 (N_18303,N_13640,N_14241);
nand U18304 (N_18304,N_14766,N_14263);
xor U18305 (N_18305,N_14219,N_14433);
xnor U18306 (N_18306,N_12832,N_13858);
nand U18307 (N_18307,N_13188,N_14668);
nor U18308 (N_18308,N_12869,N_12930);
xnor U18309 (N_18309,N_14269,N_12700);
xnor U18310 (N_18310,N_13944,N_12978);
and U18311 (N_18311,N_14723,N_14690);
nor U18312 (N_18312,N_14886,N_14752);
nor U18313 (N_18313,N_14575,N_15541);
xnor U18314 (N_18314,N_15293,N_15324);
nor U18315 (N_18315,N_12822,N_15308);
nand U18316 (N_18316,N_14092,N_15281);
nand U18317 (N_18317,N_14534,N_13069);
nor U18318 (N_18318,N_14513,N_14984);
or U18319 (N_18319,N_14308,N_13451);
or U18320 (N_18320,N_12861,N_13908);
or U18321 (N_18321,N_14421,N_15220);
xor U18322 (N_18322,N_12918,N_12681);
or U18323 (N_18323,N_13582,N_12518);
nor U18324 (N_18324,N_14838,N_15342);
xor U18325 (N_18325,N_15081,N_14773);
or U18326 (N_18326,N_14609,N_12904);
and U18327 (N_18327,N_14219,N_13390);
nor U18328 (N_18328,N_14067,N_14237);
xor U18329 (N_18329,N_15049,N_12922);
nand U18330 (N_18330,N_12904,N_13167);
nor U18331 (N_18331,N_13404,N_14150);
xnor U18332 (N_18332,N_13368,N_15282);
nand U18333 (N_18333,N_12809,N_12556);
xnor U18334 (N_18334,N_14469,N_15584);
nor U18335 (N_18335,N_12818,N_12737);
and U18336 (N_18336,N_13986,N_14255);
nor U18337 (N_18337,N_13298,N_13055);
and U18338 (N_18338,N_15382,N_13709);
xor U18339 (N_18339,N_13825,N_13350);
nor U18340 (N_18340,N_13283,N_14294);
or U18341 (N_18341,N_14417,N_13137);
nor U18342 (N_18342,N_13799,N_13258);
nand U18343 (N_18343,N_14005,N_13240);
and U18344 (N_18344,N_13960,N_13156);
and U18345 (N_18345,N_12756,N_14418);
or U18346 (N_18346,N_14280,N_12974);
nand U18347 (N_18347,N_15378,N_14027);
nor U18348 (N_18348,N_14221,N_14532);
nor U18349 (N_18349,N_15447,N_12588);
nand U18350 (N_18350,N_12857,N_13814);
nor U18351 (N_18351,N_14713,N_14070);
nor U18352 (N_18352,N_14750,N_14873);
or U18353 (N_18353,N_12911,N_14620);
nand U18354 (N_18354,N_15226,N_15074);
nor U18355 (N_18355,N_13572,N_14833);
nand U18356 (N_18356,N_15554,N_12673);
nand U18357 (N_18357,N_15597,N_14807);
xnor U18358 (N_18358,N_13059,N_15360);
or U18359 (N_18359,N_13280,N_14794);
nor U18360 (N_18360,N_15262,N_12715);
xor U18361 (N_18361,N_13055,N_12528);
and U18362 (N_18362,N_14912,N_15335);
or U18363 (N_18363,N_12648,N_14699);
xnor U18364 (N_18364,N_13714,N_15298);
or U18365 (N_18365,N_13901,N_13756);
or U18366 (N_18366,N_14469,N_14571);
nand U18367 (N_18367,N_12974,N_13838);
nand U18368 (N_18368,N_12987,N_13218);
nand U18369 (N_18369,N_15262,N_13094);
xor U18370 (N_18370,N_14327,N_13465);
xnor U18371 (N_18371,N_13200,N_15271);
xnor U18372 (N_18372,N_13915,N_13101);
nand U18373 (N_18373,N_14255,N_14329);
and U18374 (N_18374,N_13123,N_13436);
and U18375 (N_18375,N_13198,N_14406);
nand U18376 (N_18376,N_15383,N_15022);
or U18377 (N_18377,N_12516,N_15167);
nand U18378 (N_18378,N_14158,N_14980);
nor U18379 (N_18379,N_14709,N_12566);
nor U18380 (N_18380,N_13071,N_15578);
nor U18381 (N_18381,N_15124,N_14760);
nand U18382 (N_18382,N_15220,N_13816);
xor U18383 (N_18383,N_14477,N_12553);
nor U18384 (N_18384,N_13419,N_14478);
or U18385 (N_18385,N_14177,N_13948);
nor U18386 (N_18386,N_13919,N_15246);
and U18387 (N_18387,N_14306,N_13377);
and U18388 (N_18388,N_14085,N_15347);
nand U18389 (N_18389,N_14352,N_12918);
nand U18390 (N_18390,N_13687,N_13779);
nand U18391 (N_18391,N_13758,N_12967);
and U18392 (N_18392,N_13275,N_12663);
and U18393 (N_18393,N_15025,N_13140);
and U18394 (N_18394,N_14937,N_13772);
or U18395 (N_18395,N_13302,N_13381);
or U18396 (N_18396,N_15400,N_14037);
and U18397 (N_18397,N_12626,N_15189);
xnor U18398 (N_18398,N_13560,N_13755);
nor U18399 (N_18399,N_12738,N_13960);
nor U18400 (N_18400,N_14995,N_14116);
xor U18401 (N_18401,N_15238,N_14110);
and U18402 (N_18402,N_13260,N_12851);
or U18403 (N_18403,N_14740,N_14577);
nor U18404 (N_18404,N_14653,N_13544);
nand U18405 (N_18405,N_13989,N_14517);
and U18406 (N_18406,N_13714,N_14306);
or U18407 (N_18407,N_14063,N_13384);
or U18408 (N_18408,N_15092,N_13600);
or U18409 (N_18409,N_13721,N_13323);
nor U18410 (N_18410,N_13823,N_15074);
nor U18411 (N_18411,N_15523,N_15005);
nor U18412 (N_18412,N_12550,N_14295);
nor U18413 (N_18413,N_13924,N_12949);
and U18414 (N_18414,N_15020,N_15131);
or U18415 (N_18415,N_12789,N_13882);
nand U18416 (N_18416,N_13600,N_13276);
nand U18417 (N_18417,N_12582,N_14569);
nor U18418 (N_18418,N_12941,N_14321);
or U18419 (N_18419,N_13550,N_14141);
or U18420 (N_18420,N_15025,N_13268);
nor U18421 (N_18421,N_14980,N_14866);
nor U18422 (N_18422,N_15485,N_14540);
and U18423 (N_18423,N_13688,N_14862);
or U18424 (N_18424,N_14997,N_13012);
xor U18425 (N_18425,N_15448,N_15581);
nand U18426 (N_18426,N_13546,N_13237);
and U18427 (N_18427,N_12889,N_14964);
nor U18428 (N_18428,N_13362,N_13513);
nand U18429 (N_18429,N_14530,N_15543);
xnor U18430 (N_18430,N_14318,N_13738);
or U18431 (N_18431,N_14094,N_15370);
nor U18432 (N_18432,N_13198,N_13705);
and U18433 (N_18433,N_14707,N_14366);
nor U18434 (N_18434,N_12511,N_14467);
nor U18435 (N_18435,N_14295,N_15363);
nand U18436 (N_18436,N_12937,N_15588);
nor U18437 (N_18437,N_15106,N_14223);
and U18438 (N_18438,N_15096,N_14482);
or U18439 (N_18439,N_12518,N_14633);
and U18440 (N_18440,N_13230,N_13277);
nor U18441 (N_18441,N_12995,N_13336);
and U18442 (N_18442,N_13318,N_15381);
or U18443 (N_18443,N_14584,N_14295);
xor U18444 (N_18444,N_15546,N_15001);
and U18445 (N_18445,N_14075,N_13028);
nand U18446 (N_18446,N_14707,N_13292);
or U18447 (N_18447,N_14384,N_12805);
nand U18448 (N_18448,N_13831,N_13956);
nor U18449 (N_18449,N_13425,N_14703);
and U18450 (N_18450,N_14874,N_14104);
and U18451 (N_18451,N_13760,N_15295);
and U18452 (N_18452,N_14439,N_14925);
nor U18453 (N_18453,N_13062,N_13748);
and U18454 (N_18454,N_15483,N_14868);
and U18455 (N_18455,N_14708,N_14246);
nand U18456 (N_18456,N_14620,N_15038);
and U18457 (N_18457,N_14710,N_14846);
nor U18458 (N_18458,N_13141,N_13874);
or U18459 (N_18459,N_15048,N_12647);
or U18460 (N_18460,N_14207,N_12664);
nor U18461 (N_18461,N_13760,N_12561);
nand U18462 (N_18462,N_14952,N_12549);
nor U18463 (N_18463,N_12516,N_13744);
or U18464 (N_18464,N_14560,N_13576);
xnor U18465 (N_18465,N_14701,N_14245);
nor U18466 (N_18466,N_15142,N_13061);
and U18467 (N_18467,N_14853,N_15237);
nand U18468 (N_18468,N_14238,N_14441);
xnor U18469 (N_18469,N_14953,N_14956);
and U18470 (N_18470,N_14346,N_15365);
and U18471 (N_18471,N_13730,N_15231);
and U18472 (N_18472,N_13861,N_15041);
nand U18473 (N_18473,N_14795,N_12927);
or U18474 (N_18474,N_15215,N_12707);
or U18475 (N_18475,N_13148,N_12957);
nand U18476 (N_18476,N_14140,N_14918);
nand U18477 (N_18477,N_14018,N_14157);
or U18478 (N_18478,N_12564,N_14049);
nor U18479 (N_18479,N_12866,N_12896);
xnor U18480 (N_18480,N_15254,N_12679);
and U18481 (N_18481,N_12660,N_13882);
nand U18482 (N_18482,N_13710,N_15140);
or U18483 (N_18483,N_13184,N_15488);
or U18484 (N_18484,N_14874,N_15527);
xor U18485 (N_18485,N_13656,N_13401);
nor U18486 (N_18486,N_14654,N_14684);
nor U18487 (N_18487,N_12950,N_14958);
nor U18488 (N_18488,N_14445,N_13829);
nor U18489 (N_18489,N_15616,N_14638);
or U18490 (N_18490,N_13415,N_12566);
or U18491 (N_18491,N_14324,N_13352);
or U18492 (N_18492,N_14633,N_13877);
or U18493 (N_18493,N_14401,N_14303);
nor U18494 (N_18494,N_15296,N_13529);
xnor U18495 (N_18495,N_13334,N_15040);
nor U18496 (N_18496,N_12596,N_13769);
xor U18497 (N_18497,N_13775,N_13469);
or U18498 (N_18498,N_15126,N_14232);
xnor U18499 (N_18499,N_13568,N_12921);
or U18500 (N_18500,N_14216,N_12616);
or U18501 (N_18501,N_12541,N_13893);
nor U18502 (N_18502,N_14598,N_13199);
or U18503 (N_18503,N_13068,N_15612);
or U18504 (N_18504,N_13910,N_14374);
or U18505 (N_18505,N_12851,N_13848);
nand U18506 (N_18506,N_13670,N_14158);
and U18507 (N_18507,N_12986,N_12998);
and U18508 (N_18508,N_15499,N_12630);
nor U18509 (N_18509,N_14217,N_12722);
xor U18510 (N_18510,N_14121,N_13630);
xnor U18511 (N_18511,N_13486,N_15387);
nand U18512 (N_18512,N_13352,N_13777);
xor U18513 (N_18513,N_15538,N_14690);
nor U18514 (N_18514,N_13009,N_14145);
nand U18515 (N_18515,N_13190,N_13409);
nor U18516 (N_18516,N_13416,N_13587);
or U18517 (N_18517,N_15251,N_15483);
and U18518 (N_18518,N_15200,N_15420);
xnor U18519 (N_18519,N_12634,N_15362);
nand U18520 (N_18520,N_15613,N_12874);
or U18521 (N_18521,N_12625,N_13123);
xnor U18522 (N_18522,N_13120,N_14057);
nor U18523 (N_18523,N_13422,N_14333);
nor U18524 (N_18524,N_12644,N_14825);
and U18525 (N_18525,N_14905,N_14481);
xnor U18526 (N_18526,N_15130,N_13049);
nor U18527 (N_18527,N_14563,N_12532);
and U18528 (N_18528,N_15148,N_13771);
xnor U18529 (N_18529,N_12632,N_14944);
nor U18530 (N_18530,N_14620,N_13061);
nor U18531 (N_18531,N_14440,N_13092);
nand U18532 (N_18532,N_14258,N_14181);
nand U18533 (N_18533,N_14267,N_13017);
or U18534 (N_18534,N_13721,N_13925);
nand U18535 (N_18535,N_12718,N_12580);
nor U18536 (N_18536,N_14290,N_15458);
nor U18537 (N_18537,N_15028,N_14064);
nor U18538 (N_18538,N_13688,N_14505);
nor U18539 (N_18539,N_12701,N_15576);
nor U18540 (N_18540,N_12654,N_13854);
nand U18541 (N_18541,N_15011,N_13127);
and U18542 (N_18542,N_13608,N_13685);
xor U18543 (N_18543,N_14476,N_14460);
and U18544 (N_18544,N_15021,N_13424);
and U18545 (N_18545,N_13149,N_14326);
nand U18546 (N_18546,N_13657,N_15295);
nor U18547 (N_18547,N_13653,N_15133);
nor U18548 (N_18548,N_14092,N_14946);
nand U18549 (N_18549,N_13686,N_13267);
or U18550 (N_18550,N_15163,N_14959);
or U18551 (N_18551,N_15221,N_13067);
xor U18552 (N_18552,N_13779,N_12735);
xor U18553 (N_18553,N_14586,N_14108);
nor U18554 (N_18554,N_13997,N_14385);
nand U18555 (N_18555,N_14253,N_12685);
and U18556 (N_18556,N_13635,N_12850);
xor U18557 (N_18557,N_13172,N_12839);
or U18558 (N_18558,N_14279,N_14711);
xor U18559 (N_18559,N_13426,N_13868);
nand U18560 (N_18560,N_14559,N_13769);
and U18561 (N_18561,N_13760,N_12820);
and U18562 (N_18562,N_14624,N_13781);
nor U18563 (N_18563,N_14690,N_13381);
or U18564 (N_18564,N_13401,N_14942);
and U18565 (N_18565,N_15621,N_15303);
and U18566 (N_18566,N_14010,N_13403);
nor U18567 (N_18567,N_13332,N_12905);
nand U18568 (N_18568,N_12558,N_13335);
or U18569 (N_18569,N_13995,N_15151);
nor U18570 (N_18570,N_13237,N_14172);
and U18571 (N_18571,N_13867,N_14218);
nand U18572 (N_18572,N_14221,N_14924);
xnor U18573 (N_18573,N_14996,N_15359);
and U18574 (N_18574,N_15387,N_13613);
xnor U18575 (N_18575,N_14958,N_14957);
and U18576 (N_18576,N_13077,N_14557);
or U18577 (N_18577,N_15053,N_12855);
nand U18578 (N_18578,N_13898,N_12723);
xnor U18579 (N_18579,N_13713,N_15477);
and U18580 (N_18580,N_13412,N_12637);
nand U18581 (N_18581,N_14311,N_13336);
nand U18582 (N_18582,N_14098,N_12883);
and U18583 (N_18583,N_13847,N_15442);
xnor U18584 (N_18584,N_12993,N_13640);
nand U18585 (N_18585,N_13564,N_12742);
nor U18586 (N_18586,N_13271,N_15176);
nand U18587 (N_18587,N_13309,N_14504);
and U18588 (N_18588,N_13290,N_12577);
nand U18589 (N_18589,N_14000,N_12521);
xor U18590 (N_18590,N_13639,N_13314);
nand U18591 (N_18591,N_14341,N_14238);
or U18592 (N_18592,N_14844,N_14893);
xnor U18593 (N_18593,N_12689,N_14374);
or U18594 (N_18594,N_14759,N_12564);
and U18595 (N_18595,N_14082,N_12646);
and U18596 (N_18596,N_15016,N_13746);
xnor U18597 (N_18597,N_15279,N_12834);
or U18598 (N_18598,N_14307,N_12620);
or U18599 (N_18599,N_14372,N_14671);
nand U18600 (N_18600,N_13776,N_12699);
xor U18601 (N_18601,N_15193,N_14713);
nand U18602 (N_18602,N_14274,N_14242);
nand U18603 (N_18603,N_12895,N_13526);
nand U18604 (N_18604,N_14332,N_13891);
nor U18605 (N_18605,N_15165,N_14380);
or U18606 (N_18606,N_12519,N_13556);
and U18607 (N_18607,N_14107,N_12943);
and U18608 (N_18608,N_14026,N_15476);
and U18609 (N_18609,N_14284,N_13849);
and U18610 (N_18610,N_13828,N_14792);
and U18611 (N_18611,N_14709,N_15217);
nor U18612 (N_18612,N_14621,N_15478);
and U18613 (N_18613,N_14840,N_13675);
or U18614 (N_18614,N_13291,N_14588);
and U18615 (N_18615,N_14091,N_13043);
nand U18616 (N_18616,N_13775,N_14659);
nor U18617 (N_18617,N_15438,N_13793);
and U18618 (N_18618,N_13166,N_13159);
or U18619 (N_18619,N_13910,N_14666);
xor U18620 (N_18620,N_12926,N_14785);
and U18621 (N_18621,N_15349,N_14632);
or U18622 (N_18622,N_13574,N_15153);
nand U18623 (N_18623,N_15110,N_13579);
and U18624 (N_18624,N_13616,N_12557);
nor U18625 (N_18625,N_14445,N_12553);
and U18626 (N_18626,N_15038,N_12839);
and U18627 (N_18627,N_12556,N_12958);
and U18628 (N_18628,N_14718,N_13134);
nor U18629 (N_18629,N_14764,N_12692);
and U18630 (N_18630,N_14653,N_13493);
or U18631 (N_18631,N_14401,N_13162);
or U18632 (N_18632,N_14342,N_14201);
nand U18633 (N_18633,N_12821,N_14012);
nand U18634 (N_18634,N_13420,N_14390);
xnor U18635 (N_18635,N_14495,N_12929);
nor U18636 (N_18636,N_15275,N_14811);
nor U18637 (N_18637,N_15409,N_12810);
nand U18638 (N_18638,N_15527,N_13917);
nor U18639 (N_18639,N_13479,N_14342);
or U18640 (N_18640,N_12803,N_14214);
xor U18641 (N_18641,N_13711,N_14766);
and U18642 (N_18642,N_12973,N_15293);
nand U18643 (N_18643,N_14012,N_15054);
nor U18644 (N_18644,N_15494,N_12912);
nand U18645 (N_18645,N_13313,N_13157);
nor U18646 (N_18646,N_13897,N_12580);
or U18647 (N_18647,N_13934,N_12767);
and U18648 (N_18648,N_14786,N_15054);
nor U18649 (N_18649,N_13314,N_14427);
xor U18650 (N_18650,N_14839,N_13542);
nand U18651 (N_18651,N_14240,N_15551);
or U18652 (N_18652,N_14486,N_15588);
nand U18653 (N_18653,N_12693,N_13335);
xnor U18654 (N_18654,N_14387,N_13712);
nand U18655 (N_18655,N_15509,N_12628);
or U18656 (N_18656,N_15225,N_14098);
or U18657 (N_18657,N_12665,N_15384);
or U18658 (N_18658,N_14056,N_14238);
nand U18659 (N_18659,N_14614,N_12921);
nor U18660 (N_18660,N_14522,N_14026);
and U18661 (N_18661,N_14790,N_14414);
nor U18662 (N_18662,N_15555,N_14124);
nand U18663 (N_18663,N_12824,N_12967);
xor U18664 (N_18664,N_13885,N_13790);
or U18665 (N_18665,N_14807,N_13922);
xnor U18666 (N_18666,N_13993,N_15603);
xnor U18667 (N_18667,N_13297,N_12543);
nor U18668 (N_18668,N_13634,N_15097);
nor U18669 (N_18669,N_13593,N_14445);
or U18670 (N_18670,N_12611,N_12617);
nand U18671 (N_18671,N_15548,N_13600);
xor U18672 (N_18672,N_15339,N_15376);
or U18673 (N_18673,N_15104,N_14566);
xor U18674 (N_18674,N_13065,N_12519);
xnor U18675 (N_18675,N_14565,N_15537);
nand U18676 (N_18676,N_13607,N_14884);
xnor U18677 (N_18677,N_12554,N_13169);
or U18678 (N_18678,N_12655,N_13400);
nand U18679 (N_18679,N_13339,N_14221);
nand U18680 (N_18680,N_14765,N_12641);
nor U18681 (N_18681,N_14403,N_15527);
nand U18682 (N_18682,N_14002,N_12853);
nand U18683 (N_18683,N_14233,N_15164);
xor U18684 (N_18684,N_15108,N_14631);
and U18685 (N_18685,N_13045,N_15041);
or U18686 (N_18686,N_15335,N_14858);
nor U18687 (N_18687,N_13721,N_15589);
xor U18688 (N_18688,N_14767,N_12823);
xnor U18689 (N_18689,N_14646,N_14125);
xnor U18690 (N_18690,N_13675,N_12622);
or U18691 (N_18691,N_14745,N_15582);
or U18692 (N_18692,N_14760,N_14679);
nand U18693 (N_18693,N_13505,N_12532);
xnor U18694 (N_18694,N_12613,N_13955);
nand U18695 (N_18695,N_12706,N_14555);
xor U18696 (N_18696,N_14439,N_14343);
nor U18697 (N_18697,N_15152,N_14075);
nand U18698 (N_18698,N_15305,N_13709);
or U18699 (N_18699,N_13946,N_15595);
xnor U18700 (N_18700,N_14636,N_14544);
nand U18701 (N_18701,N_14543,N_14898);
xnor U18702 (N_18702,N_15033,N_14038);
nand U18703 (N_18703,N_13876,N_14302);
xnor U18704 (N_18704,N_13087,N_12701);
nor U18705 (N_18705,N_15034,N_13403);
nor U18706 (N_18706,N_15415,N_13724);
and U18707 (N_18707,N_13851,N_14116);
xor U18708 (N_18708,N_14282,N_15269);
nand U18709 (N_18709,N_15045,N_12722);
and U18710 (N_18710,N_13261,N_15038);
xnor U18711 (N_18711,N_15127,N_15483);
nor U18712 (N_18712,N_14030,N_13608);
nor U18713 (N_18713,N_13098,N_13440);
xor U18714 (N_18714,N_15406,N_13051);
nand U18715 (N_18715,N_13012,N_14176);
or U18716 (N_18716,N_14379,N_14668);
nor U18717 (N_18717,N_13615,N_13748);
and U18718 (N_18718,N_14370,N_13526);
nor U18719 (N_18719,N_13031,N_14050);
nor U18720 (N_18720,N_12535,N_13504);
nand U18721 (N_18721,N_14205,N_13310);
nand U18722 (N_18722,N_13203,N_12542);
or U18723 (N_18723,N_13344,N_15113);
nand U18724 (N_18724,N_13280,N_14065);
and U18725 (N_18725,N_12675,N_14177);
or U18726 (N_18726,N_12790,N_12636);
or U18727 (N_18727,N_14098,N_14679);
xor U18728 (N_18728,N_14091,N_13034);
nor U18729 (N_18729,N_12799,N_12681);
xnor U18730 (N_18730,N_14917,N_13202);
nand U18731 (N_18731,N_14970,N_13878);
and U18732 (N_18732,N_13549,N_14650);
nor U18733 (N_18733,N_13817,N_14838);
or U18734 (N_18734,N_13821,N_14835);
nand U18735 (N_18735,N_13693,N_13065);
nand U18736 (N_18736,N_13119,N_13387);
nand U18737 (N_18737,N_12719,N_13658);
or U18738 (N_18738,N_12642,N_13244);
nand U18739 (N_18739,N_13302,N_14394);
xor U18740 (N_18740,N_12583,N_15364);
xor U18741 (N_18741,N_13015,N_14507);
xnor U18742 (N_18742,N_12688,N_15355);
xor U18743 (N_18743,N_12823,N_14816);
or U18744 (N_18744,N_12859,N_14550);
or U18745 (N_18745,N_12886,N_14883);
nand U18746 (N_18746,N_13446,N_13607);
xor U18747 (N_18747,N_12550,N_14647);
or U18748 (N_18748,N_13954,N_15188);
nand U18749 (N_18749,N_13716,N_14993);
nor U18750 (N_18750,N_17415,N_18726);
nor U18751 (N_18751,N_17638,N_16238);
nor U18752 (N_18752,N_17962,N_16602);
xnor U18753 (N_18753,N_16034,N_15967);
or U18754 (N_18754,N_15912,N_15666);
nor U18755 (N_18755,N_18156,N_17056);
or U18756 (N_18756,N_18434,N_18550);
and U18757 (N_18757,N_16245,N_16356);
nand U18758 (N_18758,N_17584,N_16333);
nand U18759 (N_18759,N_17966,N_17728);
and U18760 (N_18760,N_17526,N_18725);
nor U18761 (N_18761,N_18112,N_17971);
xor U18762 (N_18762,N_17177,N_17620);
nand U18763 (N_18763,N_17276,N_17023);
nor U18764 (N_18764,N_17983,N_17268);
or U18765 (N_18765,N_15829,N_16263);
nand U18766 (N_18766,N_18212,N_17514);
and U18767 (N_18767,N_16858,N_18515);
nor U18768 (N_18768,N_16061,N_18409);
nor U18769 (N_18769,N_15853,N_17853);
xor U18770 (N_18770,N_17501,N_16708);
and U18771 (N_18771,N_17847,N_17167);
xor U18772 (N_18772,N_17884,N_16272);
nor U18773 (N_18773,N_16766,N_15845);
or U18774 (N_18774,N_17903,N_17445);
nand U18775 (N_18775,N_16660,N_15635);
nor U18776 (N_18776,N_16531,N_18296);
nand U18777 (N_18777,N_16881,N_17690);
nand U18778 (N_18778,N_16995,N_17367);
or U18779 (N_18779,N_18604,N_18500);
nor U18780 (N_18780,N_16822,N_17945);
nand U18781 (N_18781,N_16889,N_17979);
xnor U18782 (N_18782,N_18440,N_17138);
xor U18783 (N_18783,N_15837,N_15766);
nor U18784 (N_18784,N_18307,N_16933);
nand U18785 (N_18785,N_16295,N_17927);
nand U18786 (N_18786,N_17398,N_16131);
xor U18787 (N_18787,N_17472,N_17730);
nand U18788 (N_18788,N_17057,N_16247);
nor U18789 (N_18789,N_17529,N_15753);
nand U18790 (N_18790,N_17310,N_17609);
or U18791 (N_18791,N_18319,N_16824);
nand U18792 (N_18792,N_18048,N_16224);
nand U18793 (N_18793,N_15781,N_18000);
or U18794 (N_18794,N_18313,N_15906);
or U18795 (N_18795,N_18659,N_18126);
or U18796 (N_18796,N_17121,N_17131);
or U18797 (N_18797,N_17928,N_16310);
and U18798 (N_18798,N_18258,N_16629);
nand U18799 (N_18799,N_16994,N_15651);
or U18800 (N_18800,N_17001,N_17206);
or U18801 (N_18801,N_16320,N_18261);
nand U18802 (N_18802,N_18374,N_17916);
nand U18803 (N_18803,N_16783,N_17758);
xor U18804 (N_18804,N_18579,N_15726);
or U18805 (N_18805,N_18344,N_18616);
nor U18806 (N_18806,N_16405,N_16433);
or U18807 (N_18807,N_17414,N_17286);
or U18808 (N_18808,N_16371,N_18358);
nor U18809 (N_18809,N_17798,N_17570);
nor U18810 (N_18810,N_17302,N_18591);
and U18811 (N_18811,N_18366,N_17608);
and U18812 (N_18812,N_16427,N_15755);
nand U18813 (N_18813,N_16361,N_18511);
nand U18814 (N_18814,N_16284,N_18165);
nor U18815 (N_18815,N_18325,N_16450);
xnor U18816 (N_18816,N_15884,N_15970);
nand U18817 (N_18817,N_18477,N_16618);
nor U18818 (N_18818,N_16920,N_18394);
nor U18819 (N_18819,N_18180,N_15687);
nor U18820 (N_18820,N_18179,N_18147);
nor U18821 (N_18821,N_16759,N_15846);
or U18822 (N_18822,N_16138,N_17672);
xnor U18823 (N_18823,N_18004,N_15953);
xnor U18824 (N_18824,N_16236,N_16244);
and U18825 (N_18825,N_18581,N_16538);
or U18826 (N_18826,N_18299,N_16078);
and U18827 (N_18827,N_16515,N_15814);
nand U18828 (N_18828,N_16655,N_18494);
xor U18829 (N_18829,N_17532,N_17565);
and U18830 (N_18830,N_17178,N_17038);
or U18831 (N_18831,N_15863,N_18610);
nand U18832 (N_18832,N_17336,N_17790);
or U18833 (N_18833,N_17017,N_18486);
or U18834 (N_18834,N_17677,N_17273);
and U18835 (N_18835,N_15770,N_17186);
xnor U18836 (N_18836,N_16147,N_17282);
xor U18837 (N_18837,N_18082,N_18019);
and U18838 (N_18838,N_17588,N_15739);
xor U18839 (N_18839,N_16052,N_18640);
nor U18840 (N_18840,N_16909,N_17817);
xor U18841 (N_18841,N_16283,N_17073);
xnor U18842 (N_18842,N_18588,N_17419);
xnor U18843 (N_18843,N_16966,N_18586);
or U18844 (N_18844,N_16019,N_18392);
nand U18845 (N_18845,N_18499,N_16622);
nand U18846 (N_18846,N_16376,N_15757);
xnor U18847 (N_18847,N_16859,N_17292);
nand U18848 (N_18848,N_18736,N_17099);
and U18849 (N_18849,N_16491,N_16617);
nand U18850 (N_18850,N_18678,N_17520);
and U18851 (N_18851,N_17942,N_17880);
and U18852 (N_18852,N_16720,N_17881);
and U18853 (N_18853,N_16937,N_16146);
nor U18854 (N_18854,N_17072,N_16342);
xnor U18855 (N_18855,N_18110,N_16586);
nand U18856 (N_18856,N_16688,N_18593);
and U18857 (N_18857,N_18315,N_15668);
nor U18858 (N_18858,N_15659,N_18514);
nor U18859 (N_18859,N_17270,N_18176);
nor U18860 (N_18860,N_18701,N_15838);
xor U18861 (N_18861,N_16728,N_15657);
xor U18862 (N_18862,N_17841,N_17865);
nand U18863 (N_18863,N_18424,N_15835);
xor U18864 (N_18864,N_17750,N_15998);
nor U18865 (N_18865,N_17059,N_17124);
nand U18866 (N_18866,N_16239,N_17946);
xnor U18867 (N_18867,N_18119,N_17350);
nor U18868 (N_18868,N_18362,N_17811);
nand U18869 (N_18869,N_18158,N_15852);
and U18870 (N_18870,N_16861,N_18471);
nor U18871 (N_18871,N_16643,N_17639);
or U18872 (N_18872,N_16013,N_15678);
nand U18873 (N_18873,N_17870,N_17151);
or U18874 (N_18874,N_17778,N_18537);
or U18875 (N_18875,N_15937,N_17201);
nand U18876 (N_18876,N_17901,N_17523);
nand U18877 (N_18877,N_15729,N_16420);
xnor U18878 (N_18878,N_16888,N_16860);
and U18879 (N_18879,N_18340,N_17670);
and U18880 (N_18880,N_18252,N_17699);
xor U18881 (N_18881,N_18692,N_16004);
or U18882 (N_18882,N_18557,N_16476);
nand U18883 (N_18883,N_17914,N_17162);
or U18884 (N_18884,N_18033,N_17855);
or U18885 (N_18885,N_16950,N_15861);
and U18886 (N_18886,N_18094,N_16821);
xor U18887 (N_18887,N_18445,N_16784);
nor U18888 (N_18888,N_17256,N_17524);
and U18889 (N_18889,N_16524,N_15960);
xor U18890 (N_18890,N_17625,N_16558);
nand U18891 (N_18891,N_17566,N_16388);
or U18892 (N_18892,N_18534,N_16792);
or U18893 (N_18893,N_17999,N_18519);
and U18894 (N_18894,N_15819,N_15707);
xor U18895 (N_18895,N_17298,N_18492);
or U18896 (N_18896,N_15875,N_18411);
nand U18897 (N_18897,N_18364,N_17450);
or U18898 (N_18898,N_16401,N_18051);
nor U18899 (N_18899,N_18631,N_18136);
or U18900 (N_18900,N_16581,N_17908);
and U18901 (N_18901,N_18723,N_18143);
and U18902 (N_18902,N_16207,N_16040);
xor U18903 (N_18903,N_17637,N_18247);
nor U18904 (N_18904,N_16422,N_17198);
or U18905 (N_18905,N_17607,N_16158);
nand U18906 (N_18906,N_18259,N_17732);
or U18907 (N_18907,N_18086,N_15705);
and U18908 (N_18908,N_16169,N_18318);
xor U18909 (N_18909,N_16248,N_15716);
and U18910 (N_18910,N_18219,N_16517);
xor U18911 (N_18911,N_16605,N_17560);
or U18912 (N_18912,N_18287,N_16639);
or U18913 (N_18913,N_18383,N_17030);
xnor U18914 (N_18914,N_17838,N_16693);
nor U18915 (N_18915,N_15754,N_17851);
nor U18916 (N_18916,N_18468,N_16938);
and U18917 (N_18917,N_17071,N_17327);
nor U18918 (N_18918,N_17809,N_15921);
or U18919 (N_18919,N_17561,N_17402);
xnor U18920 (N_18920,N_17269,N_16678);
nand U18921 (N_18921,N_17305,N_16760);
nor U18922 (N_18922,N_16752,N_18023);
nor U18923 (N_18923,N_17102,N_16150);
and U18924 (N_18924,N_15832,N_17378);
and U18925 (N_18925,N_18602,N_18712);
nor U18926 (N_18926,N_17528,N_17813);
xnor U18927 (N_18927,N_17940,N_16296);
and U18928 (N_18928,N_16627,N_17895);
and U18929 (N_18929,N_18675,N_17875);
nor U18930 (N_18930,N_15639,N_16606);
or U18931 (N_18931,N_16638,N_17107);
nand U18932 (N_18932,N_17964,N_17370);
nor U18933 (N_18933,N_18160,N_17573);
or U18934 (N_18934,N_16211,N_15680);
nand U18935 (N_18935,N_18728,N_16216);
and U18936 (N_18936,N_18636,N_17209);
nand U18937 (N_18937,N_17082,N_16649);
and U18938 (N_18938,N_16345,N_15689);
xnor U18939 (N_18939,N_16363,N_16585);
nor U18940 (N_18940,N_17096,N_18217);
nor U18941 (N_18941,N_17887,N_16114);
nand U18942 (N_18942,N_17824,N_15812);
and U18943 (N_18943,N_17120,N_16520);
nor U18944 (N_18944,N_15848,N_17444);
nand U18945 (N_18945,N_16869,N_16336);
or U18946 (N_18946,N_18233,N_16458);
nor U18947 (N_18947,N_17169,N_16033);
or U18948 (N_18948,N_16805,N_17103);
and U18949 (N_18949,N_16056,N_18229);
or U18950 (N_18950,N_16790,N_17163);
xor U18951 (N_18951,N_16195,N_17645);
nand U18952 (N_18952,N_18559,N_16924);
or U18953 (N_18953,N_18702,N_16576);
xnor U18954 (N_18954,N_15656,N_15762);
or U18955 (N_18955,N_16079,N_17727);
or U18956 (N_18956,N_17068,N_17165);
nand U18957 (N_18957,N_16441,N_18495);
xor U18958 (N_18958,N_17599,N_16563);
xnor U18959 (N_18959,N_17461,N_15650);
or U18960 (N_18960,N_17430,N_17743);
xnor U18961 (N_18961,N_16703,N_17821);
and U18962 (N_18962,N_18053,N_15719);
or U18963 (N_18963,N_15866,N_16782);
xnor U18964 (N_18964,N_18128,N_16561);
or U18965 (N_18965,N_16142,N_18300);
and U18966 (N_18966,N_17788,N_18237);
xnor U18967 (N_18967,N_15785,N_17128);
xnor U18968 (N_18968,N_18303,N_16952);
xnor U18969 (N_18969,N_17510,N_17381);
and U18970 (N_18970,N_16091,N_17231);
or U18971 (N_18971,N_18360,N_18352);
xnor U18972 (N_18972,N_17541,N_15697);
nor U18973 (N_18973,N_16096,N_17271);
xor U18974 (N_18974,N_16624,N_16358);
xor U18975 (N_18975,N_17950,N_17656);
or U18976 (N_18976,N_15756,N_18647);
or U18977 (N_18977,N_17990,N_17458);
nand U18978 (N_18978,N_18115,N_16178);
or U18979 (N_18979,N_18677,N_17933);
or U18980 (N_18980,N_18510,N_18547);
or U18981 (N_18981,N_16452,N_17399);
or U18982 (N_18982,N_15767,N_17116);
and U18983 (N_18983,N_17390,N_16032);
or U18984 (N_18984,N_16574,N_17919);
and U18985 (N_18985,N_17605,N_15975);
and U18986 (N_18986,N_18524,N_16771);
nor U18987 (N_18987,N_17987,N_18085);
nor U18988 (N_18988,N_18011,N_17230);
nand U18989 (N_18989,N_16701,N_15750);
and U18990 (N_18990,N_17519,N_18443);
nand U18991 (N_18991,N_15879,N_15946);
and U18992 (N_18992,N_16212,N_18669);
nand U18993 (N_18993,N_16803,N_16447);
or U18994 (N_18994,N_16521,N_18649);
or U18995 (N_18995,N_16832,N_17185);
or U18996 (N_18996,N_15727,N_17077);
nand U18997 (N_18997,N_16732,N_17886);
or U18998 (N_18998,N_17626,N_15714);
or U18999 (N_18999,N_16875,N_16025);
nor U19000 (N_19000,N_16282,N_15942);
nand U19001 (N_19001,N_18665,N_16189);
xor U19002 (N_19002,N_17036,N_18455);
nor U19003 (N_19003,N_18517,N_17591);
nand U19004 (N_19004,N_17534,N_15712);
and U19005 (N_19005,N_17006,N_17334);
xor U19006 (N_19006,N_16497,N_16095);
and U19007 (N_19007,N_17024,N_17667);
nor U19008 (N_19008,N_16121,N_16262);
and U19009 (N_19009,N_18575,N_16974);
nand U19010 (N_19010,N_18533,N_18473);
nand U19011 (N_19011,N_17243,N_16955);
or U19012 (N_19012,N_18484,N_17234);
or U19013 (N_19013,N_17848,N_17705);
nand U19014 (N_19014,N_16003,N_16555);
xnor U19015 (N_19015,N_17470,N_16680);
nand U19016 (N_19016,N_18620,N_18312);
xnor U19017 (N_19017,N_16945,N_17545);
nand U19018 (N_19018,N_18731,N_16528);
and U19019 (N_19019,N_16038,N_15971);
xor U19020 (N_19020,N_17580,N_15646);
nor U19021 (N_19021,N_15868,N_17578);
and U19022 (N_19022,N_18069,N_16428);
nand U19023 (N_19023,N_16896,N_18410);
xnor U19024 (N_19024,N_16082,N_18555);
nor U19025 (N_19025,N_17833,N_15911);
and U19026 (N_19026,N_18348,N_18071);
or U19027 (N_19027,N_16468,N_17015);
nor U19028 (N_19028,N_16818,N_18232);
or U19029 (N_19029,N_17819,N_16650);
xnor U19030 (N_19030,N_18190,N_17547);
or U19031 (N_19031,N_16823,N_16508);
and U19032 (N_19032,N_16511,N_17299);
nand U19033 (N_19033,N_17597,N_16939);
xnor U19034 (N_19034,N_15817,N_18099);
or U19035 (N_19035,N_17823,N_15901);
nand U19036 (N_19036,N_16046,N_17248);
nand U19037 (N_19037,N_15824,N_18483);
nand U19038 (N_19038,N_15790,N_18422);
and U19039 (N_19039,N_18187,N_17630);
or U19040 (N_19040,N_17041,N_15815);
xnor U19041 (N_19041,N_16200,N_17330);
nand U19042 (N_19042,N_18626,N_16795);
and U19043 (N_19043,N_18166,N_15782);
xor U19044 (N_19044,N_16537,N_17301);
xnor U19045 (N_19045,N_18090,N_16946);
xor U19046 (N_19046,N_18558,N_15918);
xor U19047 (N_19047,N_18629,N_16291);
nand U19048 (N_19048,N_15944,N_16856);
or U19049 (N_19049,N_16741,N_18059);
nor U19050 (N_19050,N_17619,N_16704);
nor U19051 (N_19051,N_15673,N_17181);
nand U19052 (N_19052,N_15694,N_17957);
xor U19053 (N_19053,N_18530,N_17156);
and U19054 (N_19054,N_17757,N_18188);
nand U19055 (N_19055,N_17127,N_17548);
nor U19056 (N_19056,N_16827,N_16462);
xor U19057 (N_19057,N_17318,N_16658);
and U19058 (N_19058,N_16380,N_18606);
and U19059 (N_19059,N_18384,N_16503);
xnor U19060 (N_19060,N_17012,N_18087);
nor U19061 (N_19061,N_16877,N_16948);
and U19062 (N_19062,N_18706,N_16763);
or U19063 (N_19063,N_18039,N_18722);
xor U19064 (N_19064,N_15703,N_17438);
nor U19065 (N_19065,N_18135,N_17467);
and U19066 (N_19066,N_16011,N_18423);
nand U19067 (N_19067,N_18234,N_16979);
xnor U19068 (N_19068,N_18657,N_16314);
or U19069 (N_19069,N_16707,N_17644);
nor U19070 (N_19070,N_18216,N_18152);
nor U19071 (N_19071,N_18682,N_18482);
nand U19072 (N_19072,N_18578,N_18120);
and U19073 (N_19073,N_15671,N_17679);
or U19074 (N_19074,N_17039,N_17618);
nor U19075 (N_19075,N_17180,N_16059);
nor U19076 (N_19076,N_18028,N_18041);
and U19077 (N_19077,N_18161,N_16724);
xor U19078 (N_19078,N_17351,N_17382);
or U19079 (N_19079,N_15948,N_17258);
nand U19080 (N_19080,N_18543,N_18379);
xnor U19081 (N_19081,N_16712,N_16237);
or U19082 (N_19082,N_15919,N_18243);
or U19083 (N_19083,N_17417,N_16964);
and U19084 (N_19084,N_16328,N_15821);
and U19085 (N_19085,N_18407,N_15632);
and U19086 (N_19086,N_18076,N_16073);
nand U19087 (N_19087,N_16855,N_18042);
xor U19088 (N_19088,N_16005,N_16334);
xor U19089 (N_19089,N_16097,N_18615);
nand U19090 (N_19090,N_16365,N_16906);
nor U19091 (N_19091,N_17452,N_17907);
and U19092 (N_19092,N_17155,N_17818);
nor U19093 (N_19093,N_16066,N_17160);
nand U19094 (N_19094,N_17998,N_16738);
and U19095 (N_19095,N_18406,N_17556);
and U19096 (N_19096,N_15935,N_18412);
and U19097 (N_19097,N_18589,N_17852);
and U19098 (N_19098,N_18623,N_15990);
nand U19099 (N_19099,N_18202,N_17188);
or U19100 (N_19100,N_16665,N_18369);
xor U19101 (N_19101,N_16136,N_18248);
xnor U19102 (N_19102,N_17700,N_17291);
xor U19103 (N_19103,N_16852,N_16303);
and U19104 (N_19104,N_16842,N_16434);
nand U19105 (N_19105,N_15931,N_17965);
or U19106 (N_19106,N_16304,N_17506);
xor U19107 (N_19107,N_15813,N_15945);
xor U19108 (N_19108,N_17641,N_16265);
or U19109 (N_19109,N_16182,N_16299);
nand U19110 (N_19110,N_17263,N_18331);
nor U19111 (N_19111,N_16149,N_16446);
nor U19112 (N_19112,N_17683,N_16560);
xor U19113 (N_19113,N_17736,N_18679);
xor U19114 (N_19114,N_18465,N_18672);
or U19115 (N_19115,N_18159,N_17183);
and U19116 (N_19116,N_16064,N_15642);
xor U19117 (N_19117,N_17721,N_18005);
xnor U19118 (N_19118,N_18189,N_15980);
nand U19119 (N_19119,N_18246,N_17312);
nand U19120 (N_19120,N_16915,N_16975);
xnor U19121 (N_19121,N_16849,N_17320);
or U19122 (N_19122,N_18175,N_17388);
and U19123 (N_19123,N_18435,N_17911);
nand U19124 (N_19124,N_17371,N_18498);
xor U19125 (N_19125,N_16353,N_16958);
xor U19126 (N_19126,N_16865,N_16438);
or U19127 (N_19127,N_15749,N_15818);
or U19128 (N_19128,N_16396,N_16051);
xnor U19129 (N_19129,N_16267,N_18061);
xor U19130 (N_19130,N_16435,N_18502);
nor U19131 (N_19131,N_17617,N_16443);
or U19132 (N_19132,N_17376,N_17518);
or U19133 (N_19133,N_16928,N_17432);
and U19134 (N_19134,N_17577,N_16523);
nor U19135 (N_19135,N_17385,N_18538);
nor U19136 (N_19136,N_16437,N_18413);
xnor U19137 (N_19137,N_18717,N_17266);
and U19138 (N_19138,N_15677,N_18178);
nor U19139 (N_19139,N_16596,N_17315);
or U19140 (N_19140,N_16749,N_17344);
or U19141 (N_19141,N_15934,N_18562);
and U19142 (N_19142,N_17353,N_15696);
xor U19143 (N_19143,N_17693,N_17132);
or U19144 (N_19144,N_18463,N_18153);
or U19145 (N_19145,N_15828,N_15924);
or U19146 (N_19146,N_18145,N_18236);
nor U19147 (N_19147,N_16999,N_18316);
and U19148 (N_19148,N_16312,N_18345);
xnor U19149 (N_19149,N_18414,N_17706);
nor U19150 (N_19150,N_18386,N_15709);
nor U19151 (N_19151,N_18356,N_18021);
and U19152 (N_19152,N_17869,N_16120);
and U19153 (N_19153,N_18391,N_15905);
and U19154 (N_19154,N_17765,N_16455);
and U19155 (N_19155,N_17251,N_17595);
or U19156 (N_19156,N_17631,N_16816);
nor U19157 (N_19157,N_16758,N_15954);
xor U19158 (N_19158,N_17589,N_18551);
nor U19159 (N_19159,N_18196,N_18585);
xor U19160 (N_19160,N_15896,N_18129);
or U19161 (N_19161,N_16807,N_15904);
xnor U19162 (N_19162,N_16921,N_18351);
and U19163 (N_19163,N_16961,N_18680);
nand U19164 (N_19164,N_16645,N_16393);
or U19165 (N_19165,N_17592,N_16479);
xnor U19166 (N_19166,N_16084,N_16904);
xor U19167 (N_19167,N_18661,N_18609);
nand U19168 (N_19168,N_15856,N_17931);
nand U19169 (N_19169,N_17718,N_17719);
xnor U19170 (N_19170,N_16722,N_16871);
nand U19171 (N_19171,N_16395,N_16220);
nor U19172 (N_19172,N_16251,N_17303);
xor U19173 (N_19173,N_17982,N_16554);
nor U19174 (N_19174,N_16197,N_18720);
or U19175 (N_19175,N_16647,N_17832);
or U19176 (N_19176,N_16810,N_17433);
nand U19177 (N_19177,N_16868,N_18685);
nand U19178 (N_19178,N_16294,N_17440);
nand U19179 (N_19179,N_16113,N_18563);
nor U19180 (N_19180,N_18614,N_17558);
xnor U19181 (N_19181,N_17738,N_17489);
xnor U19182 (N_19182,N_17374,N_17816);
nand U19183 (N_19183,N_15734,N_16156);
nor U19184 (N_19184,N_18503,N_15955);
or U19185 (N_19185,N_16652,N_16199);
nand U19186 (N_19186,N_16954,N_16481);
nand U19187 (N_19187,N_18169,N_17929);
and U19188 (N_19188,N_16362,N_18026);
or U19189 (N_19189,N_16186,N_18047);
nor U19190 (N_19190,N_17511,N_17717);
or U19191 (N_19191,N_17492,N_17660);
nor U19192 (N_19192,N_15893,N_16599);
xor U19193 (N_19193,N_16743,N_17060);
nand U19194 (N_19194,N_16851,N_18138);
nor U19195 (N_19195,N_16054,N_16431);
xor U19196 (N_19196,N_17405,N_16746);
xnor U19197 (N_19197,N_17702,N_17742);
or U19198 (N_19198,N_17361,N_15735);
nand U19199 (N_19199,N_17002,N_17954);
or U19200 (N_19200,N_16525,N_18148);
xnor U19201 (N_19201,N_15798,N_17710);
nand U19202 (N_19202,N_18070,N_16735);
xor U19203 (N_19203,N_17642,N_18225);
xor U19204 (N_19204,N_16470,N_15839);
or U19205 (N_19205,N_18350,N_17878);
nand U19206 (N_19206,N_16773,N_17439);
xnor U19207 (N_19207,N_17250,N_17569);
or U19208 (N_19208,N_16067,N_17583);
and U19209 (N_19209,N_16550,N_18127);
xor U19210 (N_19210,N_17355,N_18083);
or U19211 (N_19211,N_16667,N_17471);
and U19212 (N_19212,N_18073,N_18240);
and U19213 (N_19213,N_16566,N_16202);
and U19214 (N_19214,N_18030,N_16072);
or U19215 (N_19215,N_17496,N_18607);
nor U19216 (N_19216,N_16278,N_17171);
xor U19217 (N_19217,N_17640,N_16159);
nand U19218 (N_19218,N_17770,N_16163);
nor U19219 (N_19219,N_17820,N_16375);
xor U19220 (N_19220,N_18522,N_16731);
nor U19221 (N_19221,N_17386,N_16213);
xnor U19222 (N_19222,N_18744,N_16632);
xnor U19223 (N_19223,N_16109,N_16473);
nor U19224 (N_19224,N_16960,N_15880);
nor U19225 (N_19225,N_15862,N_18686);
xor U19226 (N_19226,N_17070,N_18269);
or U19227 (N_19227,N_16190,N_16379);
xor U19228 (N_19228,N_16196,N_16718);
nand U19229 (N_19229,N_15995,N_17150);
nand U19230 (N_19230,N_16943,N_16165);
or U19231 (N_19231,N_16486,N_16534);
xor U19232 (N_19232,N_17055,N_16762);
nand U19233 (N_19233,N_17760,N_18116);
and U19234 (N_19234,N_15807,N_16167);
nand U19235 (N_19235,N_17600,N_16008);
or U19236 (N_19236,N_15993,N_17993);
or U19237 (N_19237,N_16171,N_18108);
and U19238 (N_19238,N_17707,N_17741);
xnor U19239 (N_19239,N_17604,N_15987);
xnor U19240 (N_19240,N_18441,N_15864);
and U19241 (N_19241,N_18485,N_17142);
and U19242 (N_19242,N_16919,N_16817);
and U19243 (N_19243,N_18065,N_16828);
xor U19244 (N_19244,N_16918,N_18564);
nor U19245 (N_19245,N_18684,N_16706);
or U19246 (N_19246,N_17125,N_17239);
or U19247 (N_19247,N_16876,N_15764);
xor U19248 (N_19248,N_15725,N_18638);
nor U19249 (N_19249,N_16118,N_17633);
or U19250 (N_19250,N_17807,N_18480);
nand U19251 (N_19251,N_18613,N_16309);
or U19252 (N_19252,N_17687,N_18057);
xnor U19253 (N_19253,N_17843,N_16739);
and U19254 (N_19254,N_16887,N_16671);
and U19255 (N_19255,N_16983,N_16297);
nor U19256 (N_19256,N_15951,N_17771);
or U19257 (N_19257,N_16498,N_16591);
nand U19258 (N_19258,N_18705,N_17035);
xor U19259 (N_19259,N_16543,N_15810);
and U19260 (N_19260,N_18676,N_16289);
and U19261 (N_19261,N_16778,N_16206);
nor U19262 (N_19262,N_18658,N_18054);
nor U19263 (N_19263,N_17428,N_16302);
xor U19264 (N_19264,N_17751,N_17013);
or U19265 (N_19265,N_16496,N_17245);
and U19266 (N_19266,N_18460,N_17348);
nor U19267 (N_19267,N_15913,N_17010);
nor U19268 (N_19268,N_17825,N_15676);
nand U19269 (N_19269,N_16987,N_16108);
xnor U19270 (N_19270,N_15702,N_17685);
nor U19271 (N_19271,N_18298,N_17499);
nand U19272 (N_19272,N_17277,N_15752);
nor U19273 (N_19273,N_15661,N_17767);
and U19274 (N_19274,N_16180,N_18710);
or U19275 (N_19275,N_17969,N_17252);
or U19276 (N_19276,N_18306,N_18222);
or U19277 (N_19277,N_15902,N_16661);
or U19278 (N_19278,N_18560,N_15688);
xnor U19279 (N_19279,N_18608,N_16094);
and U19280 (N_19280,N_15776,N_17549);
xnor U19281 (N_19281,N_18737,N_15916);
and U19282 (N_19282,N_18645,N_17483);
and U19283 (N_19283,N_17948,N_18375);
or U19284 (N_19284,N_18539,N_16410);
and U19285 (N_19285,N_18184,N_15701);
and U19286 (N_19286,N_17507,N_16233);
xnor U19287 (N_19287,N_17352,N_17321);
and U19288 (N_19288,N_16747,N_15732);
nand U19289 (N_19289,N_18239,N_17182);
nand U19290 (N_19290,N_16648,N_18475);
or U19291 (N_19291,N_17655,N_17574);
or U19292 (N_19292,N_17293,N_15965);
or U19293 (N_19293,N_15758,N_18183);
xor U19294 (N_19294,N_16311,N_15669);
or U19295 (N_19295,N_18355,N_16811);
nand U19296 (N_19296,N_18545,N_16886);
or U19297 (N_19297,N_16769,N_16258);
or U19298 (N_19298,N_17897,N_17482);
or U19299 (N_19299,N_16161,N_18611);
and U19300 (N_19300,N_18735,N_17246);
xor U19301 (N_19301,N_17341,N_17290);
and U19302 (N_19302,N_16480,N_18077);
and U19303 (N_19303,N_15647,N_16494);
nand U19304 (N_19304,N_17844,N_15898);
and U19305 (N_19305,N_15724,N_17362);
xnor U19306 (N_19306,N_17731,N_17196);
xor U19307 (N_19307,N_16836,N_17554);
and U19308 (N_19308,N_17422,N_16902);
nand U19309 (N_19309,N_15691,N_15690);
xnor U19310 (N_19310,N_17890,N_16429);
or U19311 (N_19311,N_17349,N_17648);
nand U19312 (N_19312,N_18742,N_18452);
and U19313 (N_19313,N_16100,N_15722);
nand U19314 (N_19314,N_16271,N_17020);
and U19315 (N_19315,N_16997,N_18566);
or U19316 (N_19316,N_18489,N_18031);
nand U19317 (N_19317,N_16215,N_18730);
nand U19318 (N_19318,N_15961,N_17759);
nor U19319 (N_19319,N_17708,N_18403);
or U19320 (N_19320,N_16255,N_16039);
and U19321 (N_19321,N_18734,N_16474);
nor U19322 (N_19322,N_17447,N_17190);
and U19323 (N_19323,N_17118,N_17505);
or U19324 (N_19324,N_16612,N_17335);
nor U19325 (N_19325,N_18683,N_18323);
nand U19326 (N_19326,N_15761,N_15741);
xnor U19327 (N_19327,N_17210,N_16557);
or U19328 (N_19328,N_18721,N_16081);
nor U19329 (N_19329,N_16872,N_17840);
and U19330 (N_19330,N_16959,N_17046);
nor U19331 (N_19331,N_17084,N_18198);
or U19332 (N_19332,N_16857,N_16878);
or U19333 (N_19333,N_16717,N_18436);
or U19334 (N_19334,N_17473,N_16484);
xnor U19335 (N_19335,N_16360,N_16007);
nand U19336 (N_19336,N_16510,N_18072);
and U19337 (N_19337,N_15823,N_16330);
xor U19338 (N_19338,N_17217,N_17042);
nor U19339 (N_19339,N_17537,N_18377);
xnor U19340 (N_19340,N_18091,N_17410);
and U19341 (N_19341,N_16409,N_17704);
nor U19342 (N_19342,N_17011,N_16913);
or U19343 (N_19343,N_15799,N_18400);
and U19344 (N_19344,N_16699,N_17725);
nand U19345 (N_19345,N_15738,N_17508);
nor U19346 (N_19346,N_16035,N_18621);
and U19347 (N_19347,N_16736,N_18182);
xor U19348 (N_19348,N_16323,N_17387);
xor U19349 (N_19349,N_16293,N_17225);
nand U19350 (N_19350,N_15740,N_18210);
nand U19351 (N_19351,N_18448,N_17654);
or U19352 (N_19352,N_18421,N_16306);
or U19353 (N_19353,N_17661,N_16093);
xor U19354 (N_19354,N_18218,N_16145);
or U19355 (N_19355,N_18396,N_15984);
xor U19356 (N_19356,N_17115,N_16589);
xnor U19357 (N_19357,N_18556,N_18235);
and U19358 (N_19358,N_18038,N_18474);
nand U19359 (N_19359,N_16594,N_15867);
or U19360 (N_19360,N_18253,N_17005);
nor U19361 (N_19361,N_16742,N_15991);
or U19362 (N_19362,N_16991,N_18288);
and U19363 (N_19363,N_17883,N_16932);
nor U19364 (N_19364,N_17559,N_18426);
nor U19365 (N_19365,N_16259,N_17590);
and U19366 (N_19366,N_18429,N_18535);
xnor U19367 (N_19367,N_16426,N_18745);
and U19368 (N_19368,N_18304,N_16050);
nand U19369 (N_19369,N_17476,N_17572);
nand U19370 (N_19370,N_15977,N_15663);
nand U19371 (N_19371,N_16727,N_17359);
nand U19372 (N_19372,N_16063,N_18174);
nand U19373 (N_19373,N_17674,N_16116);
or U19374 (N_19374,N_18513,N_17977);
and U19375 (N_19375,N_18294,N_16471);
xnor U19376 (N_19376,N_18724,N_16088);
nor U19377 (N_19377,N_16014,N_15728);
nor U19378 (N_19378,N_16631,N_16935);
and U19379 (N_19379,N_18141,N_17682);
nand U19380 (N_19380,N_17061,N_17996);
or U19381 (N_19381,N_15685,N_17793);
and U19382 (N_19382,N_15858,N_18220);
and U19383 (N_19383,N_17229,N_16616);
nand U19384 (N_19384,N_15908,N_17598);
and U19385 (N_19385,N_16275,N_16526);
or U19386 (N_19386,N_17935,N_18648);
or U19387 (N_19387,N_16001,N_17610);
nand U19388 (N_19388,N_17100,N_18329);
nor U19389 (N_19389,N_18670,N_18097);
and U19390 (N_19390,N_16595,N_17435);
and U19391 (N_19391,N_17274,N_18226);
xnor U19392 (N_19392,N_15800,N_17646);
xnor U19393 (N_19393,N_17981,N_17022);
xor U19394 (N_19394,N_17949,N_16608);
or U19395 (N_19395,N_17713,N_17129);
or U19396 (N_19396,N_15857,N_18181);
nor U19397 (N_19397,N_18472,N_16848);
nand U19398 (N_19398,N_16290,N_17431);
xnor U19399 (N_19399,N_16148,N_17338);
or U19400 (N_19400,N_18376,N_17856);
xnor U19401 (N_19401,N_18493,N_18633);
nor U19402 (N_19402,N_16685,N_16620);
nand U19403 (N_19403,N_16579,N_16490);
nor U19404 (N_19404,N_18273,N_15637);
or U19405 (N_19405,N_18532,N_16235);
nor U19406 (N_19406,N_16231,N_16780);
xnor U19407 (N_19407,N_17834,N_18442);
and U19408 (N_19408,N_15723,N_15943);
xor U19409 (N_19409,N_15806,N_17086);
and U19410 (N_19410,N_17249,N_17284);
nand U19411 (N_19411,N_17923,N_18584);
nor U19412 (N_19412,N_16164,N_17285);
or U19413 (N_19413,N_15649,N_17986);
nor U19414 (N_19414,N_18297,N_15759);
nand U19415 (N_19415,N_16814,N_18089);
xor U19416 (N_19416,N_17393,N_16440);
nor U19417 (N_19417,N_17941,N_18518);
nand U19418 (N_19418,N_15760,N_17579);
nor U19419 (N_19419,N_18167,N_17093);
nor U19420 (N_19420,N_17722,N_16536);
and U19421 (N_19421,N_17067,N_17004);
nand U19422 (N_19422,N_18671,N_17307);
xor U19423 (N_19423,N_16144,N_17653);
nor U19424 (N_19424,N_16664,N_18203);
or U19425 (N_19425,N_17300,N_15957);
or U19426 (N_19426,N_17546,N_18317);
or U19427 (N_19427,N_15897,N_18095);
xnor U19428 (N_19428,N_17502,N_16825);
xor U19429 (N_19429,N_16076,N_18531);
or U19430 (N_19430,N_16768,N_17392);
nor U19431 (N_19431,N_17976,N_17028);
xnor U19432 (N_19432,N_17533,N_16941);
xnor U19433 (N_19433,N_18012,N_18496);
xor U19434 (N_19434,N_16908,N_16062);
nor U19435 (N_19435,N_18244,N_17744);
or U19436 (N_19436,N_17275,N_16316);
nand U19437 (N_19437,N_16253,N_15772);
xor U19438 (N_19438,N_16575,N_17289);
nor U19439 (N_19439,N_16969,N_17323);
nand U19440 (N_19440,N_17215,N_17401);
or U19441 (N_19441,N_16493,N_17888);
xnor U19442 (N_19442,N_18464,N_18650);
nand U19443 (N_19443,N_16366,N_16653);
and U19444 (N_19444,N_18016,N_17316);
and U19445 (N_19445,N_17689,N_16126);
and U19446 (N_19446,N_16514,N_16748);
or U19447 (N_19447,N_16412,N_16725);
nand U19448 (N_19448,N_16670,N_16286);
or U19449 (N_19449,N_17262,N_17621);
nand U19450 (N_19450,N_17045,N_16377);
xnor U19451 (N_19451,N_15627,N_17459);
nand U19452 (N_19452,N_17539,N_18066);
nor U19453 (N_19453,N_16368,N_17074);
and U19454 (N_19454,N_18249,N_17154);
and U19455 (N_19455,N_16339,N_16143);
or U19456 (N_19456,N_15804,N_18043);
or U19457 (N_19457,N_17389,N_18428);
or U19458 (N_19458,N_17157,N_17238);
and U19459 (N_19459,N_16341,N_16972);
or U19460 (N_19460,N_15972,N_18321);
and U19461 (N_19461,N_16389,N_18404);
nor U19462 (N_19462,N_16914,N_17535);
nor U19463 (N_19463,N_18271,N_17531);
nor U19464 (N_19464,N_16549,N_18250);
nand U19465 (N_19465,N_16590,N_16134);
or U19466 (N_19466,N_18003,N_17885);
xnor U19467 (N_19467,N_17343,N_17850);
and U19468 (N_19468,N_16565,N_16022);
or U19469 (N_19469,N_18642,N_16765);
xor U19470 (N_19470,N_18326,N_15801);
xor U19471 (N_19471,N_17446,N_18096);
nand U19472 (N_19472,N_17090,N_18748);
xnor U19473 (N_19473,N_17221,N_18060);
nor U19474 (N_19474,N_15736,N_17455);
and U19475 (N_19475,N_18105,N_17003);
and U19476 (N_19476,N_18393,N_17799);
and U19477 (N_19477,N_17668,N_16676);
nand U19478 (N_19478,N_16249,N_17220);
xnor U19479 (N_19479,N_17783,N_15888);
nor U19480 (N_19480,N_16252,N_17781);
nor U19481 (N_19481,N_16241,N_16850);
or U19482 (N_19482,N_18367,N_16137);
nor U19483 (N_19483,N_16578,N_17065);
or U19484 (N_19484,N_15885,N_15927);
xnor U19485 (N_19485,N_17830,N_18416);
nor U19486 (N_19486,N_15830,N_16980);
or U19487 (N_19487,N_18270,N_17575);
nor U19488 (N_19488,N_18700,N_18612);
xnor U19489 (N_19489,N_17029,N_16281);
and U19490 (N_19490,N_15662,N_17874);
or U19491 (N_19491,N_16166,N_18281);
nand U19492 (N_19492,N_17170,N_17106);
nor U19493 (N_19493,N_17716,N_15748);
xor U19494 (N_19494,N_16018,N_17873);
or U19495 (N_19495,N_15826,N_16442);
xnor U19496 (N_19496,N_18173,N_17536);
and U19497 (N_19497,N_15730,N_18015);
or U19498 (N_19498,N_15938,N_18687);
or U19499 (N_19499,N_17465,N_17191);
and U19500 (N_19500,N_15715,N_16646);
nand U19501 (N_19501,N_17416,N_15877);
nand U19502 (N_19502,N_16404,N_16439);
nor U19503 (N_19503,N_15941,N_16416);
nand U19504 (N_19504,N_16628,N_17568);
nor U19505 (N_19505,N_18006,N_17542);
xnor U19506 (N_19506,N_16568,N_18525);
and U19507 (N_19507,N_16879,N_16614);
nor U19508 (N_19508,N_17772,N_18101);
nor U19509 (N_19509,N_16288,N_15909);
xnor U19510 (N_19510,N_16321,N_18652);
nor U19511 (N_19511,N_18655,N_16414);
and U19512 (N_19512,N_15859,N_16976);
xnor U19513 (N_19513,N_16268,N_17089);
nand U19514 (N_19514,N_15889,N_16598);
xor U19515 (N_19515,N_17200,N_16102);
and U19516 (N_19516,N_18282,N_17080);
xnor U19517 (N_19517,N_16923,N_17787);
nor U19518 (N_19518,N_16600,N_18634);
or U19519 (N_19519,N_16630,N_18521);
and U19520 (N_19520,N_17763,N_17696);
nand U19521 (N_19521,N_16112,N_17984);
and U19522 (N_19522,N_18568,N_17857);
nor U19523 (N_19523,N_17345,N_17469);
nor U19524 (N_19524,N_18314,N_16124);
nor U19525 (N_19525,N_16540,N_17516);
xor U19526 (N_19526,N_17628,N_18272);
nor U19527 (N_19527,N_18279,N_17317);
nand U19528 (N_19528,N_16198,N_15720);
xor U19529 (N_19529,N_16413,N_18337);
and U19530 (N_19530,N_18328,N_17810);
xnor U19531 (N_19531,N_17538,N_18438);
nor U19532 (N_19532,N_16744,N_16770);
and U19533 (N_19533,N_17159,N_17427);
or U19534 (N_19534,N_18231,N_17714);
nor U19535 (N_19535,N_15774,N_17420);
and U19536 (N_19536,N_17457,N_16812);
and U19537 (N_19537,N_17601,N_17904);
nand U19538 (N_19538,N_18334,N_15847);
and U19539 (N_19539,N_16776,N_16478);
nand U19540 (N_19540,N_17963,N_17384);
xnor U19541 (N_19541,N_18264,N_17479);
xnor U19542 (N_19542,N_17497,N_17236);
and U19543 (N_19543,N_16755,N_18497);
and U19544 (N_19544,N_18122,N_17715);
and U19545 (N_19545,N_16068,N_16392);
nand U19546 (N_19546,N_17441,N_17280);
or U19547 (N_19547,N_18201,N_18079);
xor U19548 (N_19548,N_18388,N_17139);
nor U19549 (N_19549,N_18274,N_17166);
or U19550 (N_19550,N_18646,N_17522);
nand U19551 (N_19551,N_16787,N_16463);
nor U19552 (N_19552,N_16500,N_17650);
or U19553 (N_19553,N_17729,N_16710);
nor U19554 (N_19554,N_16642,N_18570);
and U19555 (N_19555,N_17846,N_16421);
nor U19556 (N_19556,N_15874,N_16507);
or U19557 (N_19557,N_18408,N_15683);
nor U19558 (N_19558,N_17462,N_17571);
nor U19559 (N_19559,N_17795,N_16936);
or U19560 (N_19560,N_18439,N_15952);
xor U19561 (N_19561,N_18078,N_17204);
nor U19562 (N_19562,N_16250,N_16193);
xor U19563 (N_19563,N_16070,N_16354);
nor U19564 (N_19564,N_16835,N_16157);
or U19565 (N_19565,N_18466,N_16107);
nor U19566 (N_19566,N_15778,N_17801);
and U19567 (N_19567,N_18208,N_18707);
nand U19568 (N_19568,N_16609,N_18009);
xnor U19569 (N_19569,N_17669,N_16260);
nand U19570 (N_19570,N_17512,N_18154);
and U19571 (N_19571,N_17253,N_16571);
xor U19572 (N_19572,N_18123,N_16403);
and U19573 (N_19573,N_16829,N_16625);
nand U19574 (N_19574,N_17959,N_16559);
or U19575 (N_19575,N_16929,N_17110);
nand U19576 (N_19576,N_16357,N_16372);
nor U19577 (N_19577,N_16570,N_17956);
and U19578 (N_19578,N_17033,N_16218);
xnor U19579 (N_19579,N_17866,N_18280);
nor U19580 (N_19580,N_16700,N_15820);
xnor U19581 (N_19581,N_15773,N_16217);
nor U19582 (N_19582,N_16890,N_17365);
and U19583 (N_19583,N_16779,N_17775);
and U19584 (N_19584,N_18668,N_16384);
nor U19585 (N_19585,N_16682,N_16234);
or U19586 (N_19586,N_16951,N_16185);
nand U19587 (N_19587,N_17400,N_17329);
nand U19588 (N_19588,N_18656,N_17456);
and U19589 (N_19589,N_16352,N_15860);
and U19590 (N_19590,N_18215,N_16662);
or U19591 (N_19591,N_17478,N_16122);
nand U19592 (N_19592,N_15881,N_17208);
xnor U19593 (N_19593,N_18008,N_16899);
or U19594 (N_19594,N_17596,N_18104);
nand U19595 (N_19595,N_17686,N_16423);
xor U19596 (N_19596,N_17488,N_16583);
xor U19597 (N_19597,N_16327,N_18200);
nor U19598 (N_19598,N_17148,N_18191);
xor U19599 (N_19599,N_15765,N_15660);
and U19600 (N_19600,N_17521,N_18142);
or U19601 (N_19601,N_16716,N_17197);
xnor U19602 (N_19602,N_15932,N_18137);
nor U19603 (N_19603,N_16804,N_18689);
nand U19604 (N_19604,N_15992,N_15737);
and U19605 (N_19605,N_16080,N_15692);
and U19606 (N_19606,N_16695,N_16172);
or U19607 (N_19607,N_18703,N_17527);
or U19608 (N_19608,N_16506,N_16449);
or U19609 (N_19609,N_18446,N_17487);
or U19610 (N_19610,N_15962,N_18690);
xor U19611 (N_19611,N_18107,N_18046);
xnor U19612 (N_19612,N_17481,N_18738);
nand U19613 (N_19613,N_18305,N_16436);
nand U19614 (N_19614,N_17356,N_17943);
nor U19615 (N_19615,N_18283,N_16673);
or U19616 (N_19616,N_18293,N_18098);
nor U19617 (N_19617,N_18125,N_15854);
nor U19618 (N_19618,N_17363,N_16326);
xnor U19619 (N_19619,N_17244,N_16679);
nor U19620 (N_19620,N_17133,N_17854);
nor U19621 (N_19621,N_16895,N_18164);
nand U19622 (N_19622,N_18330,N_18583);
or U19623 (N_19623,N_18052,N_16518);
xnor U19624 (N_19624,N_16737,N_15929);
nand U19625 (N_19625,N_15779,N_15850);
and U19626 (N_19626,N_16378,N_18478);
nand U19627 (N_19627,N_16666,N_16794);
or U19628 (N_19628,N_18322,N_18343);
xor U19629 (N_19629,N_18625,N_17586);
nand U19630 (N_19630,N_16367,N_16119);
or U19631 (N_19631,N_18205,N_17153);
nand U19632 (N_19632,N_18363,N_17712);
xnor U19633 (N_19633,N_18749,N_17449);
nand U19634 (N_19634,N_17484,N_16292);
or U19635 (N_19635,N_17627,N_17134);
or U19636 (N_19636,N_18295,N_16337);
nand U19637 (N_19637,N_17164,N_18554);
xnor U19638 (N_19638,N_17491,N_17550);
xor U19639 (N_19639,N_17808,N_17216);
nand U19640 (N_19640,N_17937,N_16808);
nand U19641 (N_19641,N_15718,N_17726);
and U19642 (N_19642,N_16977,N_16188);
or U19643 (N_19643,N_16154,N_17517);
and U19644 (N_19644,N_15843,N_17283);
xnor U19645 (N_19645,N_16175,N_16228);
and U19646 (N_19646,N_17425,N_17991);
nor U19647 (N_19647,N_17495,N_16151);
nand U19648 (N_19648,N_18713,N_18587);
xnor U19649 (N_19649,N_15658,N_17814);
xor U19650 (N_19650,N_17676,N_18168);
nand U19651 (N_19651,N_17161,N_16499);
xnor U19652 (N_19652,N_16152,N_15968);
and U19653 (N_19653,N_16529,N_18688);
xnor U19654 (N_19654,N_17032,N_17649);
nand U19655 (N_19655,N_15733,N_16194);
or U19656 (N_19656,N_16788,N_16777);
xnor U19657 (N_19657,N_16489,N_15686);
and U19658 (N_19658,N_17173,N_18193);
nand U19659 (N_19659,N_16677,N_16277);
nand U19660 (N_19660,N_16340,N_17053);
and U19661 (N_19661,N_17369,N_16603);
and U19662 (N_19662,N_16210,N_16187);
and U19663 (N_19663,N_18622,N_17494);
or U19664 (N_19664,N_17709,N_18599);
nor U19665 (N_19665,N_16382,N_18401);
or U19666 (N_19666,N_16269,N_16015);
nor U19667 (N_19667,N_17924,N_16839);
nand U19668 (N_19668,N_16922,N_17872);
nor U19669 (N_19669,N_15842,N_17773);
xor U19670 (N_19670,N_17697,N_16456);
or U19671 (N_19671,N_15981,N_17900);
or U19672 (N_19672,N_17769,N_18102);
or U19673 (N_19673,N_18034,N_18594);
xnor U19674 (N_19674,N_16815,N_16556);
nand U19675 (N_19675,N_16225,N_17593);
nor U19676 (N_19676,N_17746,N_17831);
nor U19677 (N_19677,N_17920,N_18130);
and U19678 (N_19678,N_18567,N_15922);
nor U19679 (N_19679,N_15876,N_16044);
nand U19680 (N_19680,N_18509,N_16359);
xor U19681 (N_19681,N_17678,N_16800);
and U19682 (N_19682,N_17576,N_18398);
nand U19683 (N_19683,N_18417,N_17098);
and U19684 (N_19684,N_16483,N_15887);
and U19685 (N_19685,N_18447,N_16230);
nand U19686 (N_19686,N_16512,N_18195);
nor U19687 (N_19687,N_16105,N_17007);
nand U19688 (N_19688,N_15644,N_16021);
and U19689 (N_19689,N_16335,N_17968);
nand U19690 (N_19690,N_16485,N_16564);
and U19691 (N_19691,N_16892,N_15751);
or U19692 (N_19692,N_16846,N_16691);
and U19693 (N_19693,N_17913,N_18124);
xor U19694 (N_19694,N_17779,N_16785);
nand U19695 (N_19695,N_18501,N_16049);
or U19696 (N_19696,N_17822,N_18711);
or U19697 (N_19697,N_17265,N_16854);
nand U19698 (N_19698,N_16893,N_18662);
nand U19699 (N_19699,N_17958,N_18462);
and U19700 (N_19700,N_18427,N_17406);
nand U19701 (N_19701,N_16833,N_16065);
nor U19702 (N_19702,N_17994,N_17485);
and U19703 (N_19703,N_17179,N_16604);
xor U19704 (N_19704,N_17314,N_17849);
and U19705 (N_19705,N_15629,N_17614);
and U19706 (N_19706,N_17862,N_16417);
and U19707 (N_19707,N_16074,N_17651);
nor U19708 (N_19708,N_17143,N_15667);
nor U19709 (N_19709,N_15783,N_17168);
xor U19710 (N_19710,N_15704,N_15693);
or U19711 (N_19711,N_18549,N_16764);
nand U19712 (N_19712,N_16862,N_18619);
or U19713 (N_19713,N_18292,N_18162);
xnor U19714 (N_19714,N_17975,N_18359);
nand U19715 (N_19715,N_15746,N_15793);
nor U19716 (N_19716,N_17634,N_16419);
xnor U19717 (N_19717,N_15986,N_18456);
nor U19718 (N_19718,N_17974,N_15664);
nand U19719 (N_19719,N_17694,N_15964);
xnor U19720 (N_19720,N_18327,N_15674);
nor U19721 (N_19721,N_16592,N_16968);
or U19722 (N_19722,N_16753,N_16826);
xor U19723 (N_19723,N_18415,N_15771);
xnor U19724 (N_19724,N_16644,N_16910);
nand U19725 (N_19725,N_16873,N_17733);
xor U19726 (N_19726,N_17992,N_18320);
or U19727 (N_19727,N_16996,N_17845);
xor U19728 (N_19728,N_18603,N_17278);
nand U19729 (N_19729,N_18093,N_16373);
nand U19730 (N_19730,N_15855,N_17666);
or U19731 (N_19731,N_17812,N_18336);
and U19732 (N_19732,N_18600,N_17205);
xnor U19733 (N_19733,N_18081,N_17720);
nand U19734 (N_19734,N_18018,N_15869);
nor U19735 (N_19735,N_18699,N_16477);
and U19736 (N_19736,N_15684,N_15763);
or U19737 (N_19737,N_18378,N_17768);
xnor U19738 (N_19738,N_17894,N_18572);
nor U19739 (N_19739,N_17411,N_17014);
and U19740 (N_19740,N_16221,N_17175);
and U19741 (N_19741,N_16934,N_15899);
and U19742 (N_19742,N_17394,N_16318);
and U19743 (N_19743,N_18420,N_17172);
nand U19744 (N_19744,N_18035,N_18146);
nor U19745 (N_19745,N_17326,N_16786);
and U19746 (N_19746,N_15936,N_17202);
nand U19747 (N_19747,N_17552,N_16569);
and U19748 (N_19748,N_16687,N_16469);
xnor U19749 (N_19749,N_18488,N_17868);
and U19750 (N_19750,N_17509,N_16698);
or U19751 (N_19751,N_17031,N_18260);
and U19752 (N_19752,N_15816,N_16845);
nand U19753 (N_19753,N_17635,N_18577);
xor U19754 (N_19754,N_17871,N_16408);
nor U19755 (N_19755,N_17126,N_16229);
xor U19756 (N_19756,N_18630,N_17346);
xor U19757 (N_19757,N_16092,N_18674);
and U19758 (N_19758,N_18242,N_17858);
xor U19759 (N_19759,N_16402,N_17094);
or U19760 (N_19760,N_15994,N_16551);
nand U19761 (N_19761,N_16903,N_18133);
and U19762 (N_19762,N_16313,N_17939);
nand U19763 (N_19763,N_18192,N_18526);
and U19764 (N_19764,N_17052,N_16548);
and U19765 (N_19765,N_17681,N_15786);
and U19766 (N_19766,N_17562,N_18353);
nand U19767 (N_19767,N_16988,N_17602);
xor U19768 (N_19768,N_16775,N_15892);
nor U19769 (N_19769,N_16399,N_15956);
nand U19770 (N_19770,N_18693,N_17815);
nand U19771 (N_19771,N_18425,N_17044);
or U19772 (N_19772,N_18719,N_16465);
or U19773 (N_19773,N_16880,N_16973);
xnor U19774 (N_19774,N_18291,N_18418);
nor U19775 (N_19775,N_17581,N_17827);
and U19776 (N_19776,N_17564,N_17985);
nor U19777 (N_19777,N_17279,N_17149);
nor U19778 (N_19778,N_16801,N_17069);
xor U19779 (N_19779,N_18653,N_15988);
nand U19780 (N_19780,N_18691,N_15947);
xor U19781 (N_19781,N_15655,N_15871);
xnor U19782 (N_19782,N_15933,N_17978);
or U19783 (N_19783,N_17606,N_18139);
nand U19784 (N_19784,N_17095,N_17734);
or U19785 (N_19785,N_17257,N_15717);
nand U19786 (N_19786,N_15788,N_16944);
or U19787 (N_19787,N_18716,N_16866);
nor U19788 (N_19788,N_15706,N_16257);
nand U19789 (N_19789,N_17739,N_17259);
or U19790 (N_19790,N_17691,N_17424);
xor U19791 (N_19791,N_15654,N_18553);
or U19792 (N_19792,N_16110,N_15743);
xor U19793 (N_19793,N_18523,N_18074);
nand U19794 (N_19794,N_18529,N_17837);
nand U19795 (N_19795,N_15958,N_17786);
and U19796 (N_19796,N_17785,N_16024);
xnor U19797 (N_19797,N_18049,N_16370);
or U19798 (N_19798,N_15989,N_15742);
nand U19799 (N_19799,N_16058,N_17932);
and U19800 (N_19800,N_16640,N_17297);
xnor U19801 (N_19801,N_17088,N_16274);
and U19802 (N_19802,N_17530,N_18062);
nand U19803 (N_19803,N_18565,N_16942);
or U19804 (N_19804,N_17141,N_16751);
and U19805 (N_19805,N_16522,N_17762);
nand U19806 (N_19806,N_16301,N_16111);
and U19807 (N_19807,N_18263,N_18370);
nand U19808 (N_19808,N_16103,N_16115);
nand U19809 (N_19809,N_15966,N_17860);
and U19810 (N_19810,N_17896,N_18213);
nand U19811 (N_19811,N_17189,N_18037);
nand U19812 (N_19812,N_18666,N_16083);
or U19813 (N_19813,N_17114,N_16243);
nand U19814 (N_19814,N_15802,N_15675);
or U19815 (N_19815,N_16885,N_18569);
nor U19816 (N_19816,N_16023,N_16053);
nor U19817 (N_19817,N_18106,N_16745);
nor U19818 (N_19818,N_17776,N_16319);
nand U19819 (N_19819,N_16002,N_18199);
nand U19820 (N_19820,N_18708,N_18387);
xor U19821 (N_19821,N_15811,N_15747);
nor U19822 (N_19822,N_18746,N_18651);
nor U19823 (N_19823,N_16809,N_17421);
nand U19824 (N_19824,N_18211,N_15974);
nor U19825 (N_19825,N_18381,N_17136);
xor U19826 (N_19826,N_16432,N_16513);
nor U19827 (N_19827,N_16300,N_17412);
nand U19828 (N_19828,N_18390,N_16077);
or U19829 (N_19829,N_15996,N_17101);
xor U19830 (N_19830,N_17064,N_16867);
nand U19831 (N_19831,N_17078,N_17085);
or U19832 (N_19832,N_17104,N_17213);
nand U19833 (N_19833,N_18068,N_17658);
xnor U19834 (N_19834,N_18357,N_16205);
nor U19835 (N_19835,N_15886,N_17091);
or U19836 (N_19836,N_17135,N_16697);
xnor U19837 (N_19837,N_16347,N_16911);
nand U19838 (N_19838,N_17754,N_16613);
nand U19839 (N_19839,N_16461,N_15745);
xnor U19840 (N_19840,N_17863,N_18056);
nor U19841 (N_19841,N_17026,N_16573);
and U19842 (N_19842,N_18277,N_16183);
nor U19843 (N_19843,N_15796,N_16174);
or U19844 (N_19844,N_18617,N_16454);
xnor U19845 (N_19845,N_17212,N_18432);
or U19846 (N_19846,N_18667,N_18278);
nor U19847 (N_19847,N_18437,N_15803);
xnor U19848 (N_19848,N_17953,N_18469);
or U19849 (N_19849,N_15985,N_16089);
xor U19850 (N_19850,N_17021,N_16696);
and U19851 (N_19851,N_16069,N_16037);
nor U19852 (N_19852,N_17408,N_16394);
and U19853 (N_19853,N_17475,N_16125);
nor U19854 (N_19854,N_16398,N_17480);
and U19855 (N_19855,N_18032,N_16387);
nor U19856 (N_19856,N_16488,N_16907);
or U19857 (N_19857,N_17224,N_15873);
and U19858 (N_19858,N_17066,N_18729);
or U19859 (N_19859,N_17917,N_15939);
or U19860 (N_19860,N_16087,N_17105);
or U19861 (N_19861,N_17951,N_15834);
and U19862 (N_19862,N_17322,N_15926);
nor U19863 (N_19863,N_17585,N_18024);
xor U19864 (N_19864,N_16905,N_15805);
or U19865 (N_19865,N_18241,N_16659);
or U19866 (N_19866,N_18092,N_18520);
nor U19867 (N_19867,N_17436,N_16270);
and U19868 (N_19868,N_16891,N_18709);
nand U19869 (N_19869,N_18301,N_16155);
and U19870 (N_19870,N_18111,N_17451);
and U19871 (N_19871,N_16242,N_17882);
nand U19872 (N_19872,N_17232,N_16501);
nor U19873 (N_19873,N_17938,N_17879);
or U19874 (N_19874,N_17227,N_16381);
and U19875 (N_19875,N_18149,N_15895);
nand U19876 (N_19876,N_18598,N_17500);
or U19877 (N_19877,N_15999,N_17671);
and U19878 (N_19878,N_16981,N_16898);
or U19879 (N_19879,N_16947,N_18405);
xor U19880 (N_19880,N_18663,N_18681);
nor U19881 (N_19881,N_16582,N_16317);
nor U19882 (N_19882,N_16374,N_16668);
nor U19883 (N_19883,N_16767,N_15791);
or U19884 (N_19884,N_18402,N_17503);
and U19885 (N_19885,N_16681,N_16900);
xor U19886 (N_19886,N_15625,N_17889);
or U19887 (N_19887,N_17944,N_16457);
xor U19888 (N_19888,N_17753,N_17313);
nand U19889 (N_19889,N_17947,N_16931);
or U19890 (N_19890,N_18194,N_18632);
and U19891 (N_19891,N_18335,N_17755);
nand U19892 (N_19892,N_18382,N_16390);
nor U19893 (N_19893,N_15914,N_18479);
nor U19894 (N_19894,N_15969,N_15825);
or U19895 (N_19895,N_17267,N_16411);
nand U19896 (N_19896,N_16656,N_15891);
xor U19897 (N_19897,N_16684,N_17553);
xor U19898 (N_19898,N_17332,N_16734);
and U19899 (N_19899,N_17794,N_16036);
or U19900 (N_19900,N_17372,N_16048);
or U19901 (N_19901,N_16332,N_16611);
or U19902 (N_19902,N_15827,N_17921);
nand U19903 (N_19903,N_15878,N_17934);
nand U19904 (N_19904,N_17176,N_16593);
and U19905 (N_19905,N_15777,N_17936);
nor U19906 (N_19906,N_15731,N_16071);
and U19907 (N_19907,N_16123,N_17613);
and U19908 (N_19908,N_18673,N_17972);
nor U19909 (N_19909,N_17752,N_18001);
and U19910 (N_19910,N_18419,N_16287);
nor U19911 (N_19911,N_16689,N_17805);
nor U19912 (N_19912,N_17504,N_15634);
nor U19913 (N_19913,N_16030,N_16504);
and U19914 (N_19914,N_17498,N_16219);
xor U19915 (N_19915,N_15768,N_17366);
and U19916 (N_19916,N_18286,N_17774);
nor U19917 (N_19917,N_15626,N_18309);
or U19918 (N_19918,N_15700,N_17203);
xnor U19919 (N_19919,N_15711,N_17877);
and U19920 (N_19920,N_16406,N_16006);
nor U19921 (N_19921,N_16240,N_15797);
nand U19922 (N_19922,N_17240,N_18040);
nor U19923 (N_19923,N_17616,N_17567);
xor U19924 (N_19924,N_17861,N_18214);
xor U19925 (N_19925,N_18347,N_18644);
xnor U19926 (N_19926,N_16475,N_18064);
or U19927 (N_19927,N_16305,N_18302);
or U19928 (N_19928,N_17695,N_15809);
nand U19929 (N_19929,N_18641,N_17146);
and U19930 (N_19930,N_17112,N_17784);
nor U19931 (N_19931,N_18571,N_16962);
xor U19932 (N_19932,N_16280,N_17254);
xor U19933 (N_19933,N_16654,N_17460);
nand U19934 (N_19934,N_17804,N_18508);
nor U19935 (N_19935,N_15653,N_18341);
xnor U19936 (N_19936,N_17454,N_17152);
nand U19937 (N_19937,N_16338,N_16424);
xor U19938 (N_19938,N_17636,N_16351);
and U19939 (N_19939,N_16177,N_17448);
or U19940 (N_19940,N_16940,N_17199);
nand U19941 (N_19941,N_18150,N_18654);
and U19942 (N_19942,N_16128,N_17383);
nand U19943 (N_19943,N_17223,N_18338);
and U19944 (N_19944,N_17147,N_16675);
or U19945 (N_19945,N_16055,N_16400);
xnor U19946 (N_19946,N_17659,N_17288);
xnor U19947 (N_19947,N_15982,N_17789);
nand U19948 (N_19948,N_18453,N_16990);
nor U19949 (N_19949,N_18002,N_16509);
and U19950 (N_19950,N_18461,N_16031);
or U19951 (N_19951,N_15640,N_18601);
nand U19952 (N_19952,N_18163,N_17434);
nor U19953 (N_19953,N_18221,N_16184);
and U19954 (N_19954,N_17040,N_16168);
nand U19955 (N_19955,N_16884,N_17193);
xnor U19956 (N_19956,N_16254,N_18457);
and U19957 (N_19957,N_15794,N_17902);
or U19958 (N_19958,N_18582,N_15978);
and U19959 (N_19959,N_15721,N_17130);
or U19960 (N_19960,N_18014,N_18540);
nand U19961 (N_19961,N_16459,N_17563);
or U19962 (N_19962,N_17723,N_17097);
nand U19963 (N_19963,N_18747,N_16139);
xnor U19964 (N_19964,N_15915,N_18289);
xor U19965 (N_19965,N_17328,N_16978);
nor U19966 (N_19966,N_17407,N_18267);
nor U19967 (N_19967,N_17409,N_15792);
and U19968 (N_19968,N_17490,N_17281);
and U19969 (N_19969,N_15831,N_16204);
and U19970 (N_19970,N_17043,N_16723);
nor U19971 (N_19971,N_16702,N_17242);
or U19972 (N_19972,N_17235,N_15641);
nor U19973 (N_19973,N_16502,N_17058);
nor U19974 (N_19974,N_16897,N_17062);
and U19975 (N_19975,N_15840,N_16209);
nor U19976 (N_19976,N_17782,N_17397);
nand U19977 (N_19977,N_17083,N_18118);
xor U19978 (N_19978,N_18505,N_18186);
or U19979 (N_19979,N_18346,N_18285);
nor U19980 (N_19980,N_15917,N_17662);
or U19981 (N_19981,N_17241,N_17915);
nor U19982 (N_19982,N_17325,N_18022);
nand U19983 (N_19983,N_15645,N_15744);
nor U19984 (N_19984,N_17311,N_16385);
xor U19985 (N_19985,N_17379,N_16047);
and U19986 (N_19986,N_17339,N_15710);
xnor U19987 (N_19987,N_15652,N_17766);
nor U19988 (N_19988,N_16641,N_16173);
or U19989 (N_19989,N_17891,N_15699);
or U19990 (N_19990,N_16170,N_17926);
and U19991 (N_19991,N_16010,N_18084);
and U19992 (N_19992,N_17612,N_16539);
or U19993 (N_19993,N_16754,N_16017);
nand U19994 (N_19994,N_16674,N_18741);
nand U19995 (N_19995,N_17684,N_18660);
or U19996 (N_19996,N_18171,N_16407);
nor U19997 (N_19997,N_17443,N_16730);
or U19998 (N_19998,N_16482,N_16799);
or U19999 (N_19999,N_18595,N_18373);
xor U20000 (N_20000,N_17603,N_18528);
nand U20001 (N_20001,N_16201,N_16162);
and U20002 (N_20002,N_17261,N_18027);
xor U20003 (N_20003,N_17797,N_16901);
or U20004 (N_20004,N_16043,N_17377);
or U20005 (N_20005,N_17309,N_16601);
or U20006 (N_20006,N_18332,N_17800);
xnor U20007 (N_20007,N_17009,N_16542);
nor U20008 (N_20008,N_18385,N_15851);
xor U20009 (N_20009,N_16615,N_16383);
and U20010 (N_20010,N_17087,N_18389);
and U20011 (N_20011,N_16547,N_17442);
or U20012 (N_20012,N_17075,N_16772);
and U20013 (N_20013,N_18311,N_17144);
and U20014 (N_20014,N_17395,N_17747);
nand U20015 (N_20015,N_16223,N_18354);
and U20016 (N_20016,N_17905,N_17663);
xor U20017 (N_20017,N_17342,N_17540);
xnor U20018 (N_20018,N_18254,N_16530);
and U20019 (N_20019,N_18399,N_18144);
nor U20020 (N_20020,N_16386,N_16057);
xnor U20021 (N_20021,N_16993,N_15682);
or U20022 (N_20022,N_16714,N_17802);
and U20023 (N_20023,N_17555,N_16544);
and U20024 (N_20024,N_17018,N_16588);
nor U20025 (N_20025,N_17247,N_16349);
xnor U20026 (N_20026,N_18739,N_15695);
or U20027 (N_20027,N_16090,N_17912);
nand U20028 (N_20028,N_15940,N_15903);
nor U20029 (N_20029,N_15882,N_18113);
and U20030 (N_20030,N_16492,N_16104);
nor U20031 (N_20031,N_16705,N_18372);
or U20032 (N_20032,N_18491,N_18451);
or U20033 (N_20033,N_18664,N_18257);
xnor U20034 (N_20034,N_17111,N_16487);
nor U20035 (N_20035,N_17791,N_17623);
and U20036 (N_20036,N_18349,N_17828);
nand U20037 (N_20037,N_18007,N_15787);
and U20038 (N_20038,N_16953,N_16791);
nor U20039 (N_20039,N_15670,N_16757);
or U20040 (N_20040,N_18238,N_16545);
or U20041 (N_20041,N_16160,N_16448);
or U20042 (N_20042,N_15883,N_18454);
nor U20043 (N_20043,N_18481,N_17357);
and U20044 (N_20044,N_17260,N_18487);
xor U20045 (N_20045,N_16020,N_16636);
and U20046 (N_20046,N_18574,N_17737);
nor U20047 (N_20047,N_18025,N_17892);
or U20048 (N_20048,N_18695,N_16864);
nand U20049 (N_20049,N_16256,N_16912);
or U20050 (N_20050,N_18131,N_16967);
nor U20051 (N_20051,N_15976,N_16519);
xor U20052 (N_20052,N_17050,N_16467);
nand U20053 (N_20053,N_18643,N_17745);
or U20054 (N_20054,N_15836,N_18266);
and U20055 (N_20055,N_17113,N_17037);
or U20056 (N_20056,N_18230,N_18714);
and U20057 (N_20057,N_18512,N_16285);
and U20058 (N_20058,N_18704,N_16651);
nand U20059 (N_20059,N_17918,N_16715);
nor U20060 (N_20060,N_17864,N_17380);
nor U20061 (N_20061,N_16391,N_16874);
nor U20062 (N_20062,N_17680,N_16965);
and U20063 (N_20063,N_17092,N_18157);
xnor U20064 (N_20064,N_17027,N_17019);
and U20065 (N_20065,N_17237,N_16726);
nor U20066 (N_20066,N_16546,N_16882);
nor U20067 (N_20067,N_16028,N_16535);
or U20068 (N_20068,N_16098,N_15925);
or U20069 (N_20069,N_16298,N_18544);
nand U20070 (N_20070,N_17632,N_18592);
nand U20071 (N_20071,N_16597,N_16425);
nor U20072 (N_20072,N_18017,N_17952);
and U20073 (N_20073,N_17551,N_15822);
or U20074 (N_20074,N_18044,N_16466);
nor U20075 (N_20075,N_16982,N_17324);
nor U20076 (N_20076,N_15894,N_17054);
and U20077 (N_20077,N_17218,N_17493);
or U20078 (N_20078,N_17228,N_18088);
nand U20079 (N_20079,N_16009,N_17429);
nor U20080 (N_20080,N_15636,N_16041);
or U20081 (N_20081,N_16998,N_16266);
nor U20082 (N_20082,N_18224,N_17391);
nor U20083 (N_20083,N_16329,N_16086);
and U20084 (N_20084,N_16830,N_16307);
nor U20085 (N_20085,N_18228,N_18697);
and U20086 (N_20086,N_17211,N_17735);
or U20087 (N_20087,N_18597,N_18618);
nand U20088 (N_20088,N_16621,N_17756);
nor U20089 (N_20089,N_18080,N_17296);
and U20090 (N_20090,N_17796,N_16820);
nand U20091 (N_20091,N_17906,N_17543);
and U20092 (N_20092,N_18696,N_17893);
xnor U20093 (N_20093,N_17294,N_17331);
nor U20094 (N_20094,N_16129,N_18380);
and U20095 (N_20095,N_16637,N_17624);
nor U20096 (N_20096,N_18036,N_17622);
xnor U20097 (N_20097,N_18172,N_17544);
nand U20098 (N_20098,N_17740,N_18548);
nor U20099 (N_20099,N_15979,N_16577);
and U20100 (N_20100,N_17675,N_16844);
nand U20101 (N_20101,N_17145,N_17692);
and U20102 (N_20102,N_16099,N_16853);
and U20103 (N_20103,N_17910,N_18276);
and U20104 (N_20104,N_16445,N_16140);
nor U20105 (N_20105,N_17034,N_17304);
nor U20106 (N_20106,N_16847,N_17876);
nor U20107 (N_20107,N_17333,N_16324);
xnor U20108 (N_20108,N_15643,N_16721);
or U20109 (N_20109,N_18010,N_15630);
xnor U20110 (N_20110,N_17486,N_16464);
xnor U20111 (N_20111,N_18368,N_18639);
and U20112 (N_20112,N_18516,N_16016);
or U20113 (N_20113,N_15784,N_15808);
nand U20114 (N_20114,N_15708,N_15775);
and U20115 (N_20115,N_16181,N_17008);
xnor U20116 (N_20116,N_15769,N_15795);
or U20117 (N_20117,N_17295,N_16719);
nor U20118 (N_20118,N_16870,N_16101);
or U20119 (N_20119,N_16584,N_18536);
nor U20120 (N_20120,N_17792,N_16626);
or U20121 (N_20121,N_18310,N_16863);
nand U20122 (N_20122,N_17995,N_17643);
nor U20123 (N_20123,N_18596,N_15833);
and U20124 (N_20124,N_16325,N_17025);
xor U20125 (N_20125,N_15872,N_17629);
and U20126 (N_20126,N_16541,N_18140);
or U20127 (N_20127,N_18134,N_17360);
and U20128 (N_20128,N_17806,N_15713);
nand U20129 (N_20129,N_16355,N_18151);
or U20130 (N_20130,N_16179,N_17673);
xnor U20131 (N_20131,N_16430,N_17123);
or U20132 (N_20132,N_16709,N_15633);
nor U20133 (N_20133,N_16460,N_16516);
nand U20134 (N_20134,N_18197,N_16346);
xor U20135 (N_20135,N_18470,N_15959);
xor U20136 (N_20136,N_18170,N_16793);
nor U20137 (N_20137,N_18361,N_16261);
nor U20138 (N_20138,N_15923,N_18459);
or U20139 (N_20139,N_16619,N_18605);
nor U20140 (N_20140,N_16505,N_17255);
or U20141 (N_20141,N_16957,N_15865);
nand U20142 (N_20142,N_17899,N_17652);
and U20143 (N_20143,N_16831,N_17922);
nor U20144 (N_20144,N_16085,N_17437);
or U20145 (N_20145,N_17925,N_17347);
nand U20146 (N_20146,N_16796,N_15665);
and U20147 (N_20147,N_16153,N_18155);
nand U20148 (N_20148,N_15780,N_16970);
xor U20149 (N_20149,N_15631,N_16567);
and U20150 (N_20150,N_15849,N_16133);
or U20151 (N_20151,N_16683,N_15928);
nor U20152 (N_20152,N_17375,N_17703);
nand U20153 (N_20153,N_15910,N_17117);
nor U20154 (N_20154,N_16364,N_16106);
nor U20155 (N_20155,N_16750,N_16203);
nand U20156 (N_20156,N_17525,N_16397);
and U20157 (N_20157,N_18290,N_16672);
and U20158 (N_20158,N_18527,N_17158);
nand U20159 (N_20159,N_16694,N_16925);
xnor U20160 (N_20160,N_17463,N_16841);
and U20161 (N_20161,N_16927,N_15997);
and U20162 (N_20162,N_18029,N_16042);
nand U20163 (N_20163,N_18450,N_17337);
and U20164 (N_20164,N_16587,N_17867);
xnor U20165 (N_20165,N_16532,N_18308);
or U20166 (N_20166,N_17764,N_16246);
nand U20167 (N_20167,N_17468,N_16322);
or U20168 (N_20168,N_15841,N_16657);
nor U20169 (N_20169,N_17308,N_16843);
nand U20170 (N_20170,N_18063,N_18204);
nand U20171 (N_20171,N_18627,N_17761);
nor U20172 (N_20172,N_16610,N_18013);
or U20173 (N_20173,N_17051,N_16415);
and U20174 (N_20174,N_16176,N_17970);
nand U20175 (N_20175,N_15628,N_17909);
and U20176 (N_20176,N_17207,N_18371);
xor U20177 (N_20177,N_15950,N_18732);
or U20178 (N_20178,N_16308,N_17233);
or U20179 (N_20179,N_18490,N_17306);
nand U20180 (N_20180,N_16273,N_16633);
and U20181 (N_20181,N_18576,N_17358);
nor U20182 (N_20182,N_17513,N_16926);
nor U20183 (N_20183,N_17396,N_18552);
xnor U20184 (N_20184,N_16027,N_17980);
and U20185 (N_20185,N_17930,N_17665);
nor U20186 (N_20186,N_18255,N_16774);
or U20187 (N_20187,N_16711,N_17664);
or U20188 (N_20188,N_15789,N_18624);
nand U20189 (N_20189,N_17364,N_17835);
xor U20190 (N_20190,N_16029,N_18431);
nand U20191 (N_20191,N_15648,N_17047);
nand U20192 (N_20192,N_18209,N_16132);
or U20193 (N_20193,N_16012,N_17724);
nand U20194 (N_20194,N_16819,N_17839);
nand U20195 (N_20195,N_17701,N_16343);
or U20196 (N_20196,N_16552,N_16135);
or U20197 (N_20197,N_16060,N_18206);
nor U20198 (N_20198,N_17988,N_17464);
nor U20199 (N_20199,N_16806,N_17319);
nor U20200 (N_20200,N_17174,N_16075);
and U20201 (N_20201,N_16813,N_17859);
or U20202 (N_20202,N_16026,N_18476);
nor U20203 (N_20203,N_15890,N_16130);
xor U20204 (N_20204,N_17611,N_18132);
nand U20205 (N_20205,N_18058,N_17615);
or U20206 (N_20206,N_18430,N_18715);
and U20207 (N_20207,N_16686,N_18268);
nor U20208 (N_20208,N_17109,N_15949);
nor U20209 (N_20209,N_17474,N_18055);
nand U20210 (N_20210,N_18546,N_16789);
and U20211 (N_20211,N_16802,N_17418);
and U20212 (N_20212,N_16276,N_16222);
xnor U20213 (N_20213,N_18733,N_17582);
or U20214 (N_20214,N_16634,N_18114);
or U20215 (N_20215,N_18045,N_16985);
nand U20216 (N_20216,N_16141,N_18504);
xnor U20217 (N_20217,N_16635,N_16690);
xnor U20218 (N_20218,N_18109,N_16949);
xor U20219 (N_20219,N_18284,N_16917);
xnor U20220 (N_20220,N_16916,N_15963);
and U20221 (N_20221,N_17403,N_17373);
xor U20222 (N_20222,N_16444,N_18628);
or U20223 (N_20223,N_18580,N_18365);
xnor U20224 (N_20224,N_17967,N_16000);
xor U20225 (N_20225,N_16756,N_16127);
and U20226 (N_20226,N_16692,N_17195);
nor U20227 (N_20227,N_17264,N_16562);
and U20228 (N_20228,N_16963,N_17140);
xor U20229 (N_20229,N_18050,N_17515);
or U20230 (N_20230,N_17657,N_18573);
nand U20231 (N_20231,N_17826,N_16838);
and U20232 (N_20232,N_18542,N_18207);
or U20233 (N_20233,N_17647,N_18561);
nor U20234 (N_20234,N_17081,N_17079);
nand U20235 (N_20235,N_17184,N_16192);
xor U20236 (N_20236,N_17426,N_17594);
nor U20237 (N_20237,N_16992,N_16930);
nand U20238 (N_20238,N_17466,N_15920);
nand U20239 (N_20239,N_15983,N_18743);
or U20240 (N_20240,N_16331,N_17076);
or U20241 (N_20241,N_17587,N_18223);
and U20242 (N_20242,N_16834,N_18397);
xnor U20243 (N_20243,N_18541,N_18262);
and U20244 (N_20244,N_17836,N_16989);
xnor U20245 (N_20245,N_17973,N_17354);
and U20246 (N_20246,N_16232,N_16117);
nor U20247 (N_20247,N_17063,N_15900);
and U20248 (N_20248,N_17000,N_15698);
nor U20249 (N_20249,N_16840,N_16607);
nor U20250 (N_20250,N_18395,N_17780);
and U20251 (N_20251,N_16191,N_16971);
nor U20252 (N_20252,N_16663,N_16984);
nor U20253 (N_20253,N_16208,N_16761);
and U20254 (N_20254,N_18265,N_16418);
nand U20255 (N_20255,N_18718,N_17477);
nand U20256 (N_20256,N_17829,N_17997);
or U20257 (N_20257,N_17226,N_18449);
or U20258 (N_20258,N_17711,N_17122);
or U20259 (N_20259,N_17187,N_17049);
or U20260 (N_20260,N_17404,N_18185);
xor U20261 (N_20261,N_18103,N_16369);
or U20262 (N_20262,N_15907,N_18121);
xor U20263 (N_20263,N_16279,N_17423);
xor U20264 (N_20264,N_17960,N_18117);
nand U20265 (N_20265,N_18727,N_17955);
xor U20266 (N_20266,N_18506,N_16348);
and U20267 (N_20267,N_15844,N_18275);
nor U20268 (N_20268,N_18590,N_16315);
and U20269 (N_20269,N_18698,N_15679);
or U20270 (N_20270,N_17961,N_18433);
nand U20271 (N_20271,N_17413,N_17108);
nor U20272 (N_20272,N_16623,N_18740);
nand U20273 (N_20273,N_18020,N_17048);
xor U20274 (N_20274,N_17749,N_18458);
or U20275 (N_20275,N_16894,N_16713);
nor U20276 (N_20276,N_17192,N_16227);
and U20277 (N_20277,N_16798,N_16669);
and U20278 (N_20278,N_18256,N_18507);
xnor U20279 (N_20279,N_16986,N_18635);
xnor U20280 (N_20280,N_16533,N_17453);
and U20281 (N_20281,N_15973,N_18342);
xor U20282 (N_20282,N_18333,N_18694);
nor U20283 (N_20283,N_17557,N_17748);
nor U20284 (N_20284,N_17368,N_17016);
nand U20285 (N_20285,N_17698,N_17287);
and U20286 (N_20286,N_16344,N_15672);
or U20287 (N_20287,N_16451,N_17222);
nand U20288 (N_20288,N_17688,N_18251);
nor U20289 (N_20289,N_18444,N_16495);
nand U20290 (N_20290,N_16527,N_16837);
or U20291 (N_20291,N_17842,N_16045);
and U20292 (N_20292,N_16733,N_17194);
nand U20293 (N_20293,N_18324,N_16797);
or U20294 (N_20294,N_17137,N_18245);
or U20295 (N_20295,N_17989,N_16956);
xnor U20296 (N_20296,N_15870,N_16553);
xor U20297 (N_20297,N_17214,N_18467);
or U20298 (N_20298,N_15930,N_17272);
nand U20299 (N_20299,N_18227,N_18177);
nand U20300 (N_20300,N_17119,N_17777);
and U20301 (N_20301,N_16740,N_16264);
nor U20302 (N_20302,N_16883,N_17803);
nand U20303 (N_20303,N_15681,N_15638);
nor U20304 (N_20304,N_16350,N_18067);
nor U20305 (N_20305,N_18637,N_16472);
xor U20306 (N_20306,N_18075,N_17219);
and U20307 (N_20307,N_16580,N_18339);
nor U20308 (N_20308,N_16214,N_16453);
nor U20309 (N_20309,N_16572,N_17340);
xnor U20310 (N_20310,N_16781,N_18100);
nor U20311 (N_20311,N_16729,N_16226);
nand U20312 (N_20312,N_17898,N_16648);
or U20313 (N_20313,N_18126,N_15813);
nor U20314 (N_20314,N_17689,N_15666);
nand U20315 (N_20315,N_18133,N_16164);
nand U20316 (N_20316,N_17343,N_17425);
xor U20317 (N_20317,N_16171,N_16844);
and U20318 (N_20318,N_18242,N_18345);
or U20319 (N_20319,N_17882,N_16201);
and U20320 (N_20320,N_18000,N_16542);
xnor U20321 (N_20321,N_17136,N_16808);
and U20322 (N_20322,N_18158,N_17925);
or U20323 (N_20323,N_16426,N_18495);
nor U20324 (N_20324,N_18174,N_17985);
nand U20325 (N_20325,N_16516,N_17044);
nor U20326 (N_20326,N_15696,N_16211);
nand U20327 (N_20327,N_17990,N_16717);
and U20328 (N_20328,N_16847,N_18592);
nor U20329 (N_20329,N_16814,N_16057);
or U20330 (N_20330,N_17442,N_16854);
xnor U20331 (N_20331,N_17158,N_17000);
xnor U20332 (N_20332,N_15968,N_17619);
nand U20333 (N_20333,N_16436,N_15792);
or U20334 (N_20334,N_18403,N_16680);
nor U20335 (N_20335,N_15634,N_17908);
nor U20336 (N_20336,N_17067,N_18508);
and U20337 (N_20337,N_17783,N_16739);
nand U20338 (N_20338,N_17195,N_18745);
nor U20339 (N_20339,N_18674,N_17253);
xnor U20340 (N_20340,N_16565,N_16472);
nand U20341 (N_20341,N_17640,N_16228);
nor U20342 (N_20342,N_18267,N_17104);
nor U20343 (N_20343,N_16723,N_17529);
nand U20344 (N_20344,N_16944,N_16615);
nand U20345 (N_20345,N_16698,N_17968);
and U20346 (N_20346,N_18749,N_18261);
or U20347 (N_20347,N_16176,N_16654);
nand U20348 (N_20348,N_16196,N_17779);
xnor U20349 (N_20349,N_18074,N_16044);
and U20350 (N_20350,N_16020,N_17392);
xnor U20351 (N_20351,N_18040,N_17644);
xor U20352 (N_20352,N_18620,N_16855);
nand U20353 (N_20353,N_17729,N_16989);
or U20354 (N_20354,N_16676,N_15763);
xnor U20355 (N_20355,N_17069,N_17152);
or U20356 (N_20356,N_15759,N_18025);
xor U20357 (N_20357,N_16966,N_16628);
nand U20358 (N_20358,N_18014,N_16103);
nor U20359 (N_20359,N_18252,N_17841);
nor U20360 (N_20360,N_18438,N_17128);
or U20361 (N_20361,N_18063,N_18566);
nor U20362 (N_20362,N_17686,N_15836);
nand U20363 (N_20363,N_16710,N_18480);
nor U20364 (N_20364,N_16653,N_17297);
and U20365 (N_20365,N_16766,N_16806);
nand U20366 (N_20366,N_18324,N_15758);
nand U20367 (N_20367,N_18280,N_17089);
xor U20368 (N_20368,N_16003,N_16240);
or U20369 (N_20369,N_16616,N_15649);
nand U20370 (N_20370,N_18584,N_16044);
nand U20371 (N_20371,N_15955,N_18048);
or U20372 (N_20372,N_17576,N_16620);
nand U20373 (N_20373,N_17901,N_16146);
and U20374 (N_20374,N_15675,N_17201);
and U20375 (N_20375,N_16365,N_16728);
nor U20376 (N_20376,N_17359,N_17814);
and U20377 (N_20377,N_18273,N_18159);
xnor U20378 (N_20378,N_16541,N_17794);
nor U20379 (N_20379,N_16597,N_17270);
and U20380 (N_20380,N_16828,N_16227);
nor U20381 (N_20381,N_16827,N_17189);
or U20382 (N_20382,N_17557,N_16411);
and U20383 (N_20383,N_16893,N_16910);
nor U20384 (N_20384,N_18384,N_16162);
nand U20385 (N_20385,N_16898,N_17440);
or U20386 (N_20386,N_15921,N_17928);
nand U20387 (N_20387,N_17003,N_18463);
nor U20388 (N_20388,N_16334,N_16020);
xor U20389 (N_20389,N_16766,N_16222);
nand U20390 (N_20390,N_15778,N_17271);
nand U20391 (N_20391,N_16443,N_18558);
xnor U20392 (N_20392,N_16625,N_18249);
and U20393 (N_20393,N_17427,N_16770);
xor U20394 (N_20394,N_15679,N_18307);
nor U20395 (N_20395,N_16002,N_16913);
or U20396 (N_20396,N_16908,N_15826);
nand U20397 (N_20397,N_15763,N_16972);
xnor U20398 (N_20398,N_17256,N_17765);
nand U20399 (N_20399,N_18604,N_16218);
or U20400 (N_20400,N_16234,N_16788);
xor U20401 (N_20401,N_16771,N_17990);
nand U20402 (N_20402,N_16412,N_17177);
nand U20403 (N_20403,N_16754,N_17776);
xnor U20404 (N_20404,N_17929,N_17182);
or U20405 (N_20405,N_16234,N_18169);
nand U20406 (N_20406,N_16122,N_15632);
or U20407 (N_20407,N_16872,N_16843);
nor U20408 (N_20408,N_18652,N_17243);
nand U20409 (N_20409,N_18319,N_17801);
and U20410 (N_20410,N_17042,N_15834);
nor U20411 (N_20411,N_17994,N_16326);
or U20412 (N_20412,N_17800,N_17025);
xor U20413 (N_20413,N_17372,N_16116);
or U20414 (N_20414,N_18240,N_16971);
nor U20415 (N_20415,N_17536,N_18619);
nor U20416 (N_20416,N_16056,N_16284);
xor U20417 (N_20417,N_16380,N_17051);
xnor U20418 (N_20418,N_18614,N_17596);
xnor U20419 (N_20419,N_15759,N_15872);
nor U20420 (N_20420,N_16413,N_18523);
and U20421 (N_20421,N_18591,N_18550);
nor U20422 (N_20422,N_17127,N_15965);
nor U20423 (N_20423,N_18150,N_16192);
nor U20424 (N_20424,N_18517,N_16731);
nor U20425 (N_20425,N_18245,N_15902);
nand U20426 (N_20426,N_18419,N_17178);
or U20427 (N_20427,N_18612,N_17748);
nand U20428 (N_20428,N_17340,N_17116);
xnor U20429 (N_20429,N_16304,N_17487);
and U20430 (N_20430,N_16991,N_18328);
or U20431 (N_20431,N_16481,N_16434);
or U20432 (N_20432,N_15778,N_17180);
nor U20433 (N_20433,N_16983,N_17057);
xor U20434 (N_20434,N_17662,N_17131);
and U20435 (N_20435,N_18554,N_16411);
or U20436 (N_20436,N_16772,N_18081);
or U20437 (N_20437,N_18253,N_15830);
xor U20438 (N_20438,N_18294,N_17468);
xnor U20439 (N_20439,N_15666,N_17411);
and U20440 (N_20440,N_18116,N_17559);
nand U20441 (N_20441,N_17842,N_17296);
and U20442 (N_20442,N_18543,N_18086);
nand U20443 (N_20443,N_15910,N_18669);
and U20444 (N_20444,N_17378,N_16274);
or U20445 (N_20445,N_17398,N_15891);
or U20446 (N_20446,N_17675,N_17356);
xnor U20447 (N_20447,N_16115,N_15926);
or U20448 (N_20448,N_17471,N_16868);
nand U20449 (N_20449,N_18073,N_17562);
and U20450 (N_20450,N_16432,N_17164);
xnor U20451 (N_20451,N_18132,N_18525);
and U20452 (N_20452,N_18046,N_18183);
xor U20453 (N_20453,N_15719,N_17915);
nand U20454 (N_20454,N_18506,N_16480);
and U20455 (N_20455,N_18426,N_16786);
xnor U20456 (N_20456,N_16309,N_17752);
nor U20457 (N_20457,N_17096,N_18582);
nand U20458 (N_20458,N_16569,N_17386);
nor U20459 (N_20459,N_15860,N_17633);
xnor U20460 (N_20460,N_17344,N_18121);
nor U20461 (N_20461,N_16709,N_16266);
and U20462 (N_20462,N_18467,N_18098);
or U20463 (N_20463,N_15833,N_17479);
nor U20464 (N_20464,N_16406,N_16728);
nor U20465 (N_20465,N_16184,N_17478);
or U20466 (N_20466,N_18385,N_16508);
nor U20467 (N_20467,N_16706,N_17270);
nand U20468 (N_20468,N_16989,N_16890);
xor U20469 (N_20469,N_15740,N_15976);
or U20470 (N_20470,N_15914,N_17693);
and U20471 (N_20471,N_17748,N_15968);
xnor U20472 (N_20472,N_16847,N_17288);
xnor U20473 (N_20473,N_18335,N_16166);
nor U20474 (N_20474,N_16874,N_18522);
nand U20475 (N_20475,N_15976,N_15955);
and U20476 (N_20476,N_16095,N_16620);
nand U20477 (N_20477,N_17756,N_16829);
nor U20478 (N_20478,N_16129,N_15995);
nor U20479 (N_20479,N_17279,N_18444);
xor U20480 (N_20480,N_17637,N_15673);
nor U20481 (N_20481,N_18499,N_17832);
xor U20482 (N_20482,N_16205,N_16112);
nand U20483 (N_20483,N_17811,N_17568);
nand U20484 (N_20484,N_16983,N_18332);
or U20485 (N_20485,N_18031,N_17202);
or U20486 (N_20486,N_16026,N_18377);
xor U20487 (N_20487,N_17072,N_17803);
nor U20488 (N_20488,N_17338,N_16386);
nand U20489 (N_20489,N_15920,N_17661);
xor U20490 (N_20490,N_18122,N_17295);
and U20491 (N_20491,N_17413,N_16415);
nor U20492 (N_20492,N_16221,N_18709);
xnor U20493 (N_20493,N_16508,N_16418);
nor U20494 (N_20494,N_15847,N_17996);
xnor U20495 (N_20495,N_18422,N_16803);
xor U20496 (N_20496,N_18041,N_16835);
or U20497 (N_20497,N_15809,N_17283);
xnor U20498 (N_20498,N_16542,N_18046);
and U20499 (N_20499,N_17366,N_16903);
nand U20500 (N_20500,N_16619,N_15743);
nor U20501 (N_20501,N_15765,N_16505);
or U20502 (N_20502,N_16558,N_17952);
or U20503 (N_20503,N_18482,N_16020);
nand U20504 (N_20504,N_16950,N_17731);
and U20505 (N_20505,N_15921,N_16162);
nand U20506 (N_20506,N_18710,N_18690);
or U20507 (N_20507,N_18559,N_17513);
or U20508 (N_20508,N_16976,N_16853);
nor U20509 (N_20509,N_18424,N_17377);
nor U20510 (N_20510,N_17752,N_16939);
or U20511 (N_20511,N_17613,N_16837);
nor U20512 (N_20512,N_16583,N_16806);
and U20513 (N_20513,N_18272,N_17991);
or U20514 (N_20514,N_17233,N_15909);
or U20515 (N_20515,N_16396,N_16805);
and U20516 (N_20516,N_16894,N_18173);
nor U20517 (N_20517,N_16535,N_18697);
xnor U20518 (N_20518,N_15857,N_16312);
xnor U20519 (N_20519,N_16711,N_16312);
xnor U20520 (N_20520,N_15788,N_17264);
nor U20521 (N_20521,N_18315,N_16940);
xor U20522 (N_20522,N_16764,N_16914);
nand U20523 (N_20523,N_18008,N_17717);
or U20524 (N_20524,N_16368,N_16117);
xor U20525 (N_20525,N_18290,N_17374);
xor U20526 (N_20526,N_18735,N_18111);
xnor U20527 (N_20527,N_17507,N_15719);
nand U20528 (N_20528,N_18501,N_17536);
or U20529 (N_20529,N_16951,N_17454);
nor U20530 (N_20530,N_18150,N_18706);
nor U20531 (N_20531,N_17639,N_17832);
nand U20532 (N_20532,N_16008,N_18120);
or U20533 (N_20533,N_17022,N_17901);
xor U20534 (N_20534,N_17046,N_16289);
or U20535 (N_20535,N_15642,N_17573);
and U20536 (N_20536,N_18521,N_18205);
xor U20537 (N_20537,N_18305,N_16488);
nor U20538 (N_20538,N_16855,N_15900);
nand U20539 (N_20539,N_17893,N_15771);
and U20540 (N_20540,N_17521,N_15874);
xnor U20541 (N_20541,N_15782,N_18537);
and U20542 (N_20542,N_17453,N_16781);
and U20543 (N_20543,N_18110,N_17468);
or U20544 (N_20544,N_15648,N_16638);
or U20545 (N_20545,N_17338,N_16435);
or U20546 (N_20546,N_16239,N_15635);
nand U20547 (N_20547,N_18515,N_15788);
and U20548 (N_20548,N_16778,N_16963);
or U20549 (N_20549,N_17363,N_17452);
xor U20550 (N_20550,N_18540,N_15747);
or U20551 (N_20551,N_15673,N_16767);
or U20552 (N_20552,N_15720,N_17097);
xor U20553 (N_20553,N_17097,N_18025);
nor U20554 (N_20554,N_18566,N_18561);
nand U20555 (N_20555,N_17312,N_18281);
and U20556 (N_20556,N_17348,N_16041);
xnor U20557 (N_20557,N_18448,N_18227);
or U20558 (N_20558,N_16451,N_18233);
nand U20559 (N_20559,N_16699,N_16761);
nor U20560 (N_20560,N_18202,N_18669);
nand U20561 (N_20561,N_18033,N_17773);
or U20562 (N_20562,N_18574,N_15955);
xnor U20563 (N_20563,N_18397,N_16464);
or U20564 (N_20564,N_15790,N_18376);
xor U20565 (N_20565,N_16786,N_16395);
nor U20566 (N_20566,N_15765,N_17706);
or U20567 (N_20567,N_17774,N_16252);
nor U20568 (N_20568,N_16132,N_17332);
and U20569 (N_20569,N_18049,N_17350);
and U20570 (N_20570,N_17657,N_16978);
xor U20571 (N_20571,N_17115,N_18228);
nand U20572 (N_20572,N_16882,N_18548);
and U20573 (N_20573,N_18096,N_17264);
nor U20574 (N_20574,N_16918,N_16593);
or U20575 (N_20575,N_16354,N_16431);
or U20576 (N_20576,N_16243,N_17115);
xor U20577 (N_20577,N_16346,N_16646);
xnor U20578 (N_20578,N_18130,N_17035);
and U20579 (N_20579,N_16304,N_15648);
nand U20580 (N_20580,N_16621,N_18323);
or U20581 (N_20581,N_15786,N_15919);
and U20582 (N_20582,N_15863,N_17719);
or U20583 (N_20583,N_18417,N_17953);
nor U20584 (N_20584,N_17360,N_18025);
nor U20585 (N_20585,N_18074,N_17901);
nand U20586 (N_20586,N_18291,N_16568);
nor U20587 (N_20587,N_15840,N_16134);
nor U20588 (N_20588,N_17662,N_17490);
and U20589 (N_20589,N_18092,N_18207);
and U20590 (N_20590,N_16683,N_17564);
and U20591 (N_20591,N_15936,N_18235);
nand U20592 (N_20592,N_16136,N_18271);
or U20593 (N_20593,N_16013,N_16157);
nand U20594 (N_20594,N_16016,N_17007);
and U20595 (N_20595,N_16543,N_17558);
or U20596 (N_20596,N_15663,N_16015);
and U20597 (N_20597,N_17609,N_18643);
or U20598 (N_20598,N_16890,N_18190);
nand U20599 (N_20599,N_16388,N_18684);
nand U20600 (N_20600,N_17559,N_18603);
or U20601 (N_20601,N_18676,N_16597);
and U20602 (N_20602,N_17870,N_17811);
nand U20603 (N_20603,N_17898,N_18553);
xor U20604 (N_20604,N_18644,N_15788);
nand U20605 (N_20605,N_18135,N_15654);
nand U20606 (N_20606,N_18238,N_17376);
nor U20607 (N_20607,N_17471,N_17544);
and U20608 (N_20608,N_16239,N_18279);
xor U20609 (N_20609,N_18261,N_17033);
nand U20610 (N_20610,N_17987,N_18659);
and U20611 (N_20611,N_17979,N_18275);
and U20612 (N_20612,N_17243,N_16853);
or U20613 (N_20613,N_15704,N_15790);
xnor U20614 (N_20614,N_18541,N_16090);
xor U20615 (N_20615,N_18504,N_15628);
or U20616 (N_20616,N_16795,N_17424);
or U20617 (N_20617,N_18166,N_16896);
nand U20618 (N_20618,N_18743,N_18138);
xnor U20619 (N_20619,N_18387,N_17496);
and U20620 (N_20620,N_16302,N_17087);
and U20621 (N_20621,N_18558,N_18496);
nor U20622 (N_20622,N_18262,N_16081);
and U20623 (N_20623,N_16367,N_17346);
nand U20624 (N_20624,N_16168,N_17075);
and U20625 (N_20625,N_16886,N_15695);
nor U20626 (N_20626,N_16968,N_15661);
and U20627 (N_20627,N_17753,N_15944);
nand U20628 (N_20628,N_15840,N_18074);
xor U20629 (N_20629,N_17127,N_17673);
xor U20630 (N_20630,N_18137,N_16724);
or U20631 (N_20631,N_16642,N_16380);
and U20632 (N_20632,N_16923,N_16595);
and U20633 (N_20633,N_15932,N_16917);
xnor U20634 (N_20634,N_18738,N_18414);
or U20635 (N_20635,N_17186,N_17934);
xor U20636 (N_20636,N_16184,N_16120);
and U20637 (N_20637,N_17495,N_16491);
nand U20638 (N_20638,N_16394,N_16243);
and U20639 (N_20639,N_17637,N_18175);
and U20640 (N_20640,N_17235,N_16322);
and U20641 (N_20641,N_17849,N_15747);
xor U20642 (N_20642,N_18012,N_17147);
nand U20643 (N_20643,N_16285,N_15651);
nor U20644 (N_20644,N_17763,N_18094);
xor U20645 (N_20645,N_15745,N_17111);
or U20646 (N_20646,N_15836,N_16641);
nand U20647 (N_20647,N_16359,N_15658);
nand U20648 (N_20648,N_17615,N_17061);
xor U20649 (N_20649,N_17640,N_16508);
nor U20650 (N_20650,N_17196,N_16226);
nor U20651 (N_20651,N_16347,N_18617);
or U20652 (N_20652,N_18542,N_18366);
nand U20653 (N_20653,N_16239,N_15811);
xnor U20654 (N_20654,N_16103,N_15691);
nand U20655 (N_20655,N_17037,N_16273);
and U20656 (N_20656,N_17992,N_18568);
nor U20657 (N_20657,N_17675,N_17317);
or U20658 (N_20658,N_16829,N_18280);
nor U20659 (N_20659,N_16789,N_18282);
or U20660 (N_20660,N_18718,N_15751);
and U20661 (N_20661,N_16671,N_16707);
xor U20662 (N_20662,N_16903,N_15775);
nand U20663 (N_20663,N_16342,N_16336);
nand U20664 (N_20664,N_17501,N_17849);
nor U20665 (N_20665,N_16257,N_17152);
or U20666 (N_20666,N_17956,N_18561);
nand U20667 (N_20667,N_16840,N_16716);
nand U20668 (N_20668,N_18322,N_18428);
or U20669 (N_20669,N_18251,N_16664);
or U20670 (N_20670,N_17936,N_18090);
and U20671 (N_20671,N_17568,N_16197);
nor U20672 (N_20672,N_16769,N_17222);
or U20673 (N_20673,N_16274,N_16434);
or U20674 (N_20674,N_18620,N_16830);
xor U20675 (N_20675,N_17880,N_15683);
and U20676 (N_20676,N_16666,N_17582);
nand U20677 (N_20677,N_18402,N_17902);
xnor U20678 (N_20678,N_17704,N_16451);
nor U20679 (N_20679,N_18179,N_16511);
nor U20680 (N_20680,N_17456,N_17826);
and U20681 (N_20681,N_16824,N_18016);
or U20682 (N_20682,N_16663,N_17092);
nor U20683 (N_20683,N_16129,N_17220);
nor U20684 (N_20684,N_18364,N_17261);
and U20685 (N_20685,N_15801,N_17840);
or U20686 (N_20686,N_18301,N_17065);
xnor U20687 (N_20687,N_18191,N_16446);
xnor U20688 (N_20688,N_15893,N_16031);
and U20689 (N_20689,N_16318,N_18562);
nand U20690 (N_20690,N_17861,N_18490);
nor U20691 (N_20691,N_17954,N_17498);
xor U20692 (N_20692,N_17947,N_18664);
xor U20693 (N_20693,N_15669,N_18346);
nand U20694 (N_20694,N_17109,N_18357);
nand U20695 (N_20695,N_15869,N_15773);
and U20696 (N_20696,N_16291,N_16087);
and U20697 (N_20697,N_16020,N_18058);
and U20698 (N_20698,N_16088,N_17360);
nor U20699 (N_20699,N_15692,N_17435);
and U20700 (N_20700,N_18450,N_16330);
nand U20701 (N_20701,N_17619,N_17063);
nor U20702 (N_20702,N_17924,N_17466);
nor U20703 (N_20703,N_16615,N_17771);
xnor U20704 (N_20704,N_18655,N_17046);
or U20705 (N_20705,N_15918,N_15886);
nand U20706 (N_20706,N_16956,N_16825);
xor U20707 (N_20707,N_17272,N_18554);
or U20708 (N_20708,N_18255,N_17265);
nor U20709 (N_20709,N_16824,N_15871);
and U20710 (N_20710,N_16519,N_16493);
or U20711 (N_20711,N_15759,N_16323);
nor U20712 (N_20712,N_16842,N_17427);
nor U20713 (N_20713,N_18009,N_18565);
nor U20714 (N_20714,N_18485,N_16577);
and U20715 (N_20715,N_16879,N_15901);
and U20716 (N_20716,N_18340,N_16787);
xor U20717 (N_20717,N_17348,N_17448);
or U20718 (N_20718,N_17423,N_17476);
or U20719 (N_20719,N_17353,N_16700);
and U20720 (N_20720,N_15869,N_17078);
or U20721 (N_20721,N_16794,N_16665);
or U20722 (N_20722,N_16815,N_16607);
and U20723 (N_20723,N_17281,N_18502);
xnor U20724 (N_20724,N_18104,N_18153);
xnor U20725 (N_20725,N_17843,N_17424);
xor U20726 (N_20726,N_18489,N_17973);
or U20727 (N_20727,N_17996,N_16155);
xor U20728 (N_20728,N_18256,N_17710);
nor U20729 (N_20729,N_18580,N_15930);
nor U20730 (N_20730,N_16398,N_17646);
nand U20731 (N_20731,N_18141,N_17938);
nand U20732 (N_20732,N_16150,N_17009);
or U20733 (N_20733,N_17689,N_15781);
nor U20734 (N_20734,N_16542,N_17246);
or U20735 (N_20735,N_17129,N_16605);
or U20736 (N_20736,N_17424,N_16729);
xnor U20737 (N_20737,N_16065,N_16183);
nor U20738 (N_20738,N_16325,N_17775);
nand U20739 (N_20739,N_17143,N_16495);
xnor U20740 (N_20740,N_17100,N_17489);
and U20741 (N_20741,N_16819,N_18143);
nor U20742 (N_20742,N_18178,N_16724);
or U20743 (N_20743,N_17368,N_16169);
or U20744 (N_20744,N_18572,N_16526);
nand U20745 (N_20745,N_15925,N_18521);
and U20746 (N_20746,N_16217,N_15661);
and U20747 (N_20747,N_16159,N_16956);
nor U20748 (N_20748,N_16731,N_15646);
and U20749 (N_20749,N_18711,N_17480);
xor U20750 (N_20750,N_17810,N_16544);
and U20751 (N_20751,N_18727,N_16120);
xnor U20752 (N_20752,N_16160,N_16407);
and U20753 (N_20753,N_18454,N_16207);
or U20754 (N_20754,N_16682,N_18728);
xnor U20755 (N_20755,N_15909,N_16018);
nor U20756 (N_20756,N_16931,N_16531);
nand U20757 (N_20757,N_18227,N_16496);
nor U20758 (N_20758,N_17345,N_16733);
nand U20759 (N_20759,N_17047,N_17472);
or U20760 (N_20760,N_17878,N_18571);
xor U20761 (N_20761,N_17749,N_18501);
nand U20762 (N_20762,N_16112,N_15780);
nor U20763 (N_20763,N_16026,N_15651);
and U20764 (N_20764,N_16692,N_17239);
nand U20765 (N_20765,N_16287,N_16303);
and U20766 (N_20766,N_16810,N_16909);
or U20767 (N_20767,N_16021,N_16712);
nor U20768 (N_20768,N_17801,N_18127);
xnor U20769 (N_20769,N_18028,N_18389);
xnor U20770 (N_20770,N_18133,N_16239);
or U20771 (N_20771,N_18240,N_15921);
and U20772 (N_20772,N_17446,N_15689);
or U20773 (N_20773,N_17646,N_16714);
xor U20774 (N_20774,N_18730,N_17957);
nor U20775 (N_20775,N_15767,N_18095);
xor U20776 (N_20776,N_17581,N_16824);
or U20777 (N_20777,N_17728,N_17674);
xnor U20778 (N_20778,N_17441,N_17168);
or U20779 (N_20779,N_16153,N_17538);
xnor U20780 (N_20780,N_18740,N_18236);
xnor U20781 (N_20781,N_17683,N_18160);
nor U20782 (N_20782,N_17288,N_15716);
xor U20783 (N_20783,N_18373,N_18556);
and U20784 (N_20784,N_16025,N_16495);
nor U20785 (N_20785,N_16419,N_17745);
nand U20786 (N_20786,N_17595,N_17436);
xnor U20787 (N_20787,N_18065,N_16566);
xnor U20788 (N_20788,N_17520,N_18299);
xor U20789 (N_20789,N_16069,N_18340);
and U20790 (N_20790,N_17883,N_18387);
and U20791 (N_20791,N_16309,N_16100);
xnor U20792 (N_20792,N_16651,N_17122);
xnor U20793 (N_20793,N_15855,N_18350);
or U20794 (N_20794,N_16287,N_16971);
xnor U20795 (N_20795,N_17128,N_16112);
nor U20796 (N_20796,N_17359,N_18410);
nand U20797 (N_20797,N_16626,N_15990);
nor U20798 (N_20798,N_17010,N_17564);
nand U20799 (N_20799,N_16138,N_16067);
or U20800 (N_20800,N_17708,N_16261);
or U20801 (N_20801,N_17509,N_17909);
and U20802 (N_20802,N_16156,N_17493);
nand U20803 (N_20803,N_18566,N_17728);
nand U20804 (N_20804,N_15962,N_17968);
nand U20805 (N_20805,N_17392,N_16548);
or U20806 (N_20806,N_16130,N_17237);
nor U20807 (N_20807,N_16159,N_17578);
and U20808 (N_20808,N_16399,N_17775);
or U20809 (N_20809,N_17526,N_17467);
or U20810 (N_20810,N_15766,N_15701);
xnor U20811 (N_20811,N_18729,N_16245);
nor U20812 (N_20812,N_18025,N_16040);
xor U20813 (N_20813,N_16998,N_18651);
xor U20814 (N_20814,N_16312,N_17765);
and U20815 (N_20815,N_15970,N_17123);
xor U20816 (N_20816,N_16126,N_16923);
nor U20817 (N_20817,N_18291,N_18298);
xor U20818 (N_20818,N_16493,N_15692);
nand U20819 (N_20819,N_17691,N_17476);
xor U20820 (N_20820,N_17966,N_18559);
nor U20821 (N_20821,N_15772,N_16809);
nor U20822 (N_20822,N_18624,N_15960);
or U20823 (N_20823,N_17083,N_17440);
and U20824 (N_20824,N_18739,N_16984);
or U20825 (N_20825,N_18022,N_16664);
nand U20826 (N_20826,N_16416,N_17058);
nor U20827 (N_20827,N_16724,N_16307);
and U20828 (N_20828,N_17321,N_17038);
nor U20829 (N_20829,N_16230,N_18489);
or U20830 (N_20830,N_17541,N_17841);
and U20831 (N_20831,N_17049,N_17040);
nor U20832 (N_20832,N_16758,N_18130);
or U20833 (N_20833,N_18598,N_18516);
and U20834 (N_20834,N_16587,N_16669);
xnor U20835 (N_20835,N_16676,N_18497);
and U20836 (N_20836,N_17878,N_16424);
nor U20837 (N_20837,N_18009,N_15649);
or U20838 (N_20838,N_15647,N_18117);
xnor U20839 (N_20839,N_16785,N_18410);
nor U20840 (N_20840,N_17121,N_16703);
xnor U20841 (N_20841,N_16785,N_17288);
or U20842 (N_20842,N_15780,N_17457);
or U20843 (N_20843,N_18393,N_15630);
nor U20844 (N_20844,N_18203,N_18305);
nand U20845 (N_20845,N_15727,N_16463);
or U20846 (N_20846,N_16728,N_16585);
xor U20847 (N_20847,N_15666,N_16620);
nor U20848 (N_20848,N_15650,N_16880);
nand U20849 (N_20849,N_17553,N_17879);
and U20850 (N_20850,N_17922,N_18279);
or U20851 (N_20851,N_17075,N_16707);
nor U20852 (N_20852,N_15693,N_16076);
or U20853 (N_20853,N_15794,N_18309);
nand U20854 (N_20854,N_16249,N_17599);
nor U20855 (N_20855,N_16108,N_17117);
nor U20856 (N_20856,N_17952,N_17969);
xnor U20857 (N_20857,N_18540,N_16337);
and U20858 (N_20858,N_17502,N_16075);
and U20859 (N_20859,N_18380,N_18585);
xnor U20860 (N_20860,N_18293,N_16879);
xnor U20861 (N_20861,N_15835,N_15673);
nor U20862 (N_20862,N_15653,N_17518);
xnor U20863 (N_20863,N_16242,N_17226);
and U20864 (N_20864,N_17083,N_16087);
and U20865 (N_20865,N_16880,N_17782);
nand U20866 (N_20866,N_18730,N_18319);
xor U20867 (N_20867,N_17198,N_17767);
or U20868 (N_20868,N_18422,N_17612);
and U20869 (N_20869,N_16773,N_16040);
xnor U20870 (N_20870,N_17165,N_16655);
nand U20871 (N_20871,N_18134,N_16352);
xnor U20872 (N_20872,N_17031,N_17230);
and U20873 (N_20873,N_18063,N_17427);
nand U20874 (N_20874,N_15664,N_16260);
nor U20875 (N_20875,N_16747,N_17445);
nand U20876 (N_20876,N_16821,N_18496);
or U20877 (N_20877,N_18247,N_15784);
nand U20878 (N_20878,N_18122,N_17738);
xnor U20879 (N_20879,N_18222,N_18469);
nand U20880 (N_20880,N_16589,N_17844);
nor U20881 (N_20881,N_15928,N_16420);
and U20882 (N_20882,N_18088,N_16520);
or U20883 (N_20883,N_15638,N_16273);
or U20884 (N_20884,N_17362,N_18159);
or U20885 (N_20885,N_16573,N_17690);
nand U20886 (N_20886,N_16275,N_18120);
nor U20887 (N_20887,N_17117,N_18080);
or U20888 (N_20888,N_17567,N_15902);
nand U20889 (N_20889,N_17876,N_17200);
xnor U20890 (N_20890,N_18443,N_17959);
nand U20891 (N_20891,N_16031,N_18020);
xor U20892 (N_20892,N_17827,N_15872);
xor U20893 (N_20893,N_16924,N_15718);
and U20894 (N_20894,N_15884,N_17014);
or U20895 (N_20895,N_16705,N_16425);
nor U20896 (N_20896,N_16203,N_17173);
or U20897 (N_20897,N_16443,N_16422);
and U20898 (N_20898,N_16607,N_16018);
xor U20899 (N_20899,N_16716,N_17451);
xor U20900 (N_20900,N_15625,N_17906);
nand U20901 (N_20901,N_18641,N_16511);
nand U20902 (N_20902,N_16169,N_16796);
nand U20903 (N_20903,N_16296,N_16996);
xor U20904 (N_20904,N_18087,N_15893);
or U20905 (N_20905,N_16802,N_16793);
or U20906 (N_20906,N_16751,N_16897);
xor U20907 (N_20907,N_18024,N_16295);
xnor U20908 (N_20908,N_16411,N_17452);
nand U20909 (N_20909,N_18682,N_16550);
and U20910 (N_20910,N_18545,N_16594);
xnor U20911 (N_20911,N_18651,N_15942);
xnor U20912 (N_20912,N_16194,N_18467);
nand U20913 (N_20913,N_15719,N_17380);
and U20914 (N_20914,N_18173,N_17584);
and U20915 (N_20915,N_18313,N_17287);
xor U20916 (N_20916,N_16501,N_18020);
and U20917 (N_20917,N_17213,N_16034);
and U20918 (N_20918,N_17395,N_16407);
nor U20919 (N_20919,N_18353,N_16158);
nand U20920 (N_20920,N_16213,N_15675);
nor U20921 (N_20921,N_16025,N_17950);
nor U20922 (N_20922,N_18268,N_16627);
nand U20923 (N_20923,N_16256,N_18573);
xor U20924 (N_20924,N_17983,N_15667);
nor U20925 (N_20925,N_16495,N_18211);
xor U20926 (N_20926,N_16166,N_16404);
nor U20927 (N_20927,N_16154,N_15741);
and U20928 (N_20928,N_15855,N_16774);
xnor U20929 (N_20929,N_16106,N_17675);
xor U20930 (N_20930,N_16847,N_17493);
nand U20931 (N_20931,N_16574,N_17528);
xor U20932 (N_20932,N_16478,N_16113);
or U20933 (N_20933,N_16925,N_15982);
and U20934 (N_20934,N_18098,N_16358);
and U20935 (N_20935,N_17511,N_15923);
or U20936 (N_20936,N_17449,N_16432);
nor U20937 (N_20937,N_16356,N_17949);
xnor U20938 (N_20938,N_18404,N_18536);
or U20939 (N_20939,N_16281,N_16810);
and U20940 (N_20940,N_17095,N_16450);
nand U20941 (N_20941,N_18519,N_17308);
or U20942 (N_20942,N_17505,N_16932);
nand U20943 (N_20943,N_18274,N_15939);
or U20944 (N_20944,N_15689,N_16436);
or U20945 (N_20945,N_18674,N_15940);
and U20946 (N_20946,N_15654,N_17787);
and U20947 (N_20947,N_15694,N_17979);
nand U20948 (N_20948,N_15670,N_17480);
or U20949 (N_20949,N_16486,N_16283);
or U20950 (N_20950,N_16375,N_17495);
xor U20951 (N_20951,N_16764,N_16644);
xor U20952 (N_20952,N_17875,N_18280);
and U20953 (N_20953,N_18426,N_16489);
nor U20954 (N_20954,N_18455,N_18351);
xnor U20955 (N_20955,N_17039,N_15804);
xor U20956 (N_20956,N_16518,N_16795);
and U20957 (N_20957,N_17665,N_16010);
or U20958 (N_20958,N_18064,N_17857);
or U20959 (N_20959,N_16451,N_16016);
nor U20960 (N_20960,N_16987,N_16954);
and U20961 (N_20961,N_17992,N_16163);
or U20962 (N_20962,N_16921,N_17728);
nor U20963 (N_20963,N_16813,N_17050);
nand U20964 (N_20964,N_16843,N_16647);
or U20965 (N_20965,N_17703,N_18265);
xnor U20966 (N_20966,N_15915,N_18672);
and U20967 (N_20967,N_18424,N_16214);
xor U20968 (N_20968,N_16097,N_16139);
nor U20969 (N_20969,N_18378,N_16763);
nand U20970 (N_20970,N_16297,N_15939);
or U20971 (N_20971,N_16687,N_16894);
or U20972 (N_20972,N_16879,N_17941);
nor U20973 (N_20973,N_16127,N_17321);
xnor U20974 (N_20974,N_18684,N_17888);
xnor U20975 (N_20975,N_17153,N_17258);
xor U20976 (N_20976,N_16241,N_18501);
nor U20977 (N_20977,N_18412,N_16220);
nor U20978 (N_20978,N_17966,N_16368);
or U20979 (N_20979,N_17674,N_16780);
and U20980 (N_20980,N_15701,N_17370);
and U20981 (N_20981,N_18633,N_17052);
xor U20982 (N_20982,N_17787,N_15917);
nor U20983 (N_20983,N_17587,N_16222);
nand U20984 (N_20984,N_18350,N_15836);
and U20985 (N_20985,N_15999,N_17794);
nor U20986 (N_20986,N_17545,N_17176);
xnor U20987 (N_20987,N_15701,N_17840);
xor U20988 (N_20988,N_16001,N_16522);
nor U20989 (N_20989,N_18351,N_17527);
xnor U20990 (N_20990,N_16027,N_16342);
xor U20991 (N_20991,N_17835,N_18098);
and U20992 (N_20992,N_15858,N_15998);
and U20993 (N_20993,N_17737,N_17886);
nand U20994 (N_20994,N_16808,N_18607);
xnor U20995 (N_20995,N_17740,N_17150);
nor U20996 (N_20996,N_17868,N_16361);
and U20997 (N_20997,N_16402,N_15686);
nand U20998 (N_20998,N_17916,N_15784);
nand U20999 (N_20999,N_17114,N_15640);
xnor U21000 (N_21000,N_16547,N_17376);
nand U21001 (N_21001,N_15936,N_17413);
or U21002 (N_21002,N_16090,N_15743);
and U21003 (N_21003,N_15910,N_15739);
xnor U21004 (N_21004,N_17009,N_17882);
and U21005 (N_21005,N_17718,N_18533);
nor U21006 (N_21006,N_15713,N_16582);
nor U21007 (N_21007,N_15864,N_17311);
nand U21008 (N_21008,N_16739,N_18663);
nand U21009 (N_21009,N_18741,N_16358);
nor U21010 (N_21010,N_17203,N_17819);
or U21011 (N_21011,N_18267,N_18630);
nor U21012 (N_21012,N_18133,N_17520);
and U21013 (N_21013,N_16213,N_15820);
xnor U21014 (N_21014,N_17809,N_18581);
nor U21015 (N_21015,N_15963,N_17437);
xor U21016 (N_21016,N_15903,N_16946);
and U21017 (N_21017,N_18293,N_18167);
nor U21018 (N_21018,N_15882,N_17208);
or U21019 (N_21019,N_17937,N_18336);
and U21020 (N_21020,N_18413,N_18534);
xor U21021 (N_21021,N_15792,N_18425);
nand U21022 (N_21022,N_18734,N_17255);
xnor U21023 (N_21023,N_17419,N_17129);
nor U21024 (N_21024,N_18132,N_17147);
and U21025 (N_21025,N_18490,N_17321);
nand U21026 (N_21026,N_16214,N_17502);
nor U21027 (N_21027,N_16443,N_16399);
nand U21028 (N_21028,N_18532,N_18701);
and U21029 (N_21029,N_17808,N_18440);
nand U21030 (N_21030,N_17272,N_15999);
or U21031 (N_21031,N_18397,N_17402);
xor U21032 (N_21032,N_18359,N_17358);
nor U21033 (N_21033,N_17245,N_16490);
xor U21034 (N_21034,N_16073,N_16983);
xnor U21035 (N_21035,N_16677,N_16880);
xor U21036 (N_21036,N_18599,N_18556);
xnor U21037 (N_21037,N_18696,N_15891);
nand U21038 (N_21038,N_17486,N_16793);
or U21039 (N_21039,N_18639,N_18023);
and U21040 (N_21040,N_18381,N_17048);
or U21041 (N_21041,N_18074,N_16338);
or U21042 (N_21042,N_18699,N_16723);
and U21043 (N_21043,N_17287,N_17938);
xor U21044 (N_21044,N_15944,N_16779);
or U21045 (N_21045,N_15694,N_15973);
nor U21046 (N_21046,N_17266,N_15833);
or U21047 (N_21047,N_18677,N_16343);
nand U21048 (N_21048,N_16529,N_18076);
or U21049 (N_21049,N_17983,N_16635);
xor U21050 (N_21050,N_18005,N_15971);
and U21051 (N_21051,N_16557,N_18479);
nand U21052 (N_21052,N_18620,N_18127);
or U21053 (N_21053,N_16619,N_16966);
xnor U21054 (N_21054,N_18720,N_18574);
xor U21055 (N_21055,N_16225,N_18658);
and U21056 (N_21056,N_17988,N_15969);
nor U21057 (N_21057,N_17131,N_17692);
nand U21058 (N_21058,N_16551,N_17887);
nand U21059 (N_21059,N_16389,N_17672);
nand U21060 (N_21060,N_17274,N_17618);
nor U21061 (N_21061,N_18183,N_18562);
nor U21062 (N_21062,N_15849,N_16554);
xor U21063 (N_21063,N_15660,N_17080);
nand U21064 (N_21064,N_16152,N_16019);
xor U21065 (N_21065,N_17626,N_18425);
nand U21066 (N_21066,N_16117,N_18321);
nand U21067 (N_21067,N_18228,N_18248);
xnor U21068 (N_21068,N_18528,N_15879);
nor U21069 (N_21069,N_16041,N_17743);
xnor U21070 (N_21070,N_17464,N_17137);
nand U21071 (N_21071,N_16098,N_16161);
xor U21072 (N_21072,N_17288,N_18664);
or U21073 (N_21073,N_18592,N_17216);
xor U21074 (N_21074,N_17717,N_17972);
or U21075 (N_21075,N_16034,N_16100);
nor U21076 (N_21076,N_15640,N_18515);
or U21077 (N_21077,N_18149,N_16202);
or U21078 (N_21078,N_15887,N_17708);
and U21079 (N_21079,N_18724,N_17304);
xor U21080 (N_21080,N_17804,N_15689);
and U21081 (N_21081,N_17802,N_15902);
or U21082 (N_21082,N_17157,N_15991);
nor U21083 (N_21083,N_17167,N_17899);
nor U21084 (N_21084,N_17544,N_16971);
and U21085 (N_21085,N_18173,N_15900);
or U21086 (N_21086,N_16508,N_16923);
or U21087 (N_21087,N_16085,N_17796);
or U21088 (N_21088,N_18107,N_15984);
and U21089 (N_21089,N_18645,N_15943);
nor U21090 (N_21090,N_16226,N_17403);
and U21091 (N_21091,N_18094,N_16490);
and U21092 (N_21092,N_16548,N_16353);
xnor U21093 (N_21093,N_16829,N_16631);
or U21094 (N_21094,N_18564,N_16823);
nor U21095 (N_21095,N_16024,N_17465);
or U21096 (N_21096,N_16390,N_16061);
nand U21097 (N_21097,N_17419,N_16109);
and U21098 (N_21098,N_17509,N_16080);
nand U21099 (N_21099,N_18040,N_18384);
or U21100 (N_21100,N_17662,N_16818);
nor U21101 (N_21101,N_17798,N_17475);
nand U21102 (N_21102,N_16615,N_17495);
or U21103 (N_21103,N_15847,N_16284);
nor U21104 (N_21104,N_17155,N_17281);
xnor U21105 (N_21105,N_16940,N_16626);
and U21106 (N_21106,N_17487,N_17316);
and U21107 (N_21107,N_16147,N_16233);
and U21108 (N_21108,N_16344,N_16252);
and U21109 (N_21109,N_17846,N_16937);
nand U21110 (N_21110,N_16153,N_18130);
nand U21111 (N_21111,N_17841,N_16074);
and U21112 (N_21112,N_15655,N_15776);
nor U21113 (N_21113,N_17638,N_15956);
and U21114 (N_21114,N_17765,N_17083);
or U21115 (N_21115,N_15920,N_15963);
and U21116 (N_21116,N_18540,N_18446);
xnor U21117 (N_21117,N_16243,N_16224);
or U21118 (N_21118,N_15817,N_17604);
or U21119 (N_21119,N_18102,N_16461);
xor U21120 (N_21120,N_17519,N_17665);
or U21121 (N_21121,N_18096,N_17157);
or U21122 (N_21122,N_16686,N_17169);
xor U21123 (N_21123,N_16151,N_15652);
nor U21124 (N_21124,N_17193,N_15709);
and U21125 (N_21125,N_18413,N_16160);
and U21126 (N_21126,N_16897,N_15986);
and U21127 (N_21127,N_15694,N_17622);
xnor U21128 (N_21128,N_16844,N_17105);
nor U21129 (N_21129,N_16264,N_16745);
nand U21130 (N_21130,N_17006,N_18563);
xnor U21131 (N_21131,N_15936,N_16451);
or U21132 (N_21132,N_18548,N_17834);
xnor U21133 (N_21133,N_17452,N_17060);
or U21134 (N_21134,N_16289,N_16922);
and U21135 (N_21135,N_18510,N_17987);
nor U21136 (N_21136,N_15667,N_17538);
nor U21137 (N_21137,N_17718,N_18124);
and U21138 (N_21138,N_16674,N_18144);
nand U21139 (N_21139,N_17320,N_16739);
and U21140 (N_21140,N_16276,N_16628);
xor U21141 (N_21141,N_18264,N_17082);
or U21142 (N_21142,N_18343,N_17061);
nand U21143 (N_21143,N_17235,N_18717);
and U21144 (N_21144,N_16155,N_18257);
or U21145 (N_21145,N_18731,N_17606);
or U21146 (N_21146,N_15962,N_17798);
nand U21147 (N_21147,N_17820,N_15714);
and U21148 (N_21148,N_17972,N_18266);
nand U21149 (N_21149,N_17427,N_16046);
or U21150 (N_21150,N_16736,N_17363);
or U21151 (N_21151,N_17277,N_15783);
or U21152 (N_21152,N_15649,N_18463);
nand U21153 (N_21153,N_16241,N_16311);
or U21154 (N_21154,N_18706,N_17279);
and U21155 (N_21155,N_16506,N_16257);
or U21156 (N_21156,N_17789,N_17142);
or U21157 (N_21157,N_16187,N_16612);
nand U21158 (N_21158,N_16217,N_17695);
or U21159 (N_21159,N_17868,N_18226);
and U21160 (N_21160,N_17383,N_17857);
and U21161 (N_21161,N_18571,N_15995);
or U21162 (N_21162,N_16837,N_15788);
and U21163 (N_21163,N_18510,N_16918);
xor U21164 (N_21164,N_18316,N_15732);
nand U21165 (N_21165,N_15983,N_18228);
xnor U21166 (N_21166,N_18587,N_16064);
or U21167 (N_21167,N_16615,N_18464);
nand U21168 (N_21168,N_18375,N_15875);
nor U21169 (N_21169,N_15960,N_17233);
nor U21170 (N_21170,N_16066,N_17708);
or U21171 (N_21171,N_17597,N_16667);
and U21172 (N_21172,N_15906,N_15992);
or U21173 (N_21173,N_16933,N_16376);
xnor U21174 (N_21174,N_15760,N_17053);
or U21175 (N_21175,N_15706,N_15876);
nand U21176 (N_21176,N_16408,N_17529);
xnor U21177 (N_21177,N_17757,N_16395);
and U21178 (N_21178,N_16691,N_16579);
and U21179 (N_21179,N_17590,N_17569);
xor U21180 (N_21180,N_18439,N_15636);
nor U21181 (N_21181,N_18078,N_15892);
nand U21182 (N_21182,N_16998,N_18208);
xnor U21183 (N_21183,N_17680,N_16630);
and U21184 (N_21184,N_15641,N_18465);
nor U21185 (N_21185,N_17556,N_15950);
or U21186 (N_21186,N_17432,N_16123);
nor U21187 (N_21187,N_17323,N_17238);
xor U21188 (N_21188,N_18091,N_18418);
nand U21189 (N_21189,N_16929,N_17758);
and U21190 (N_21190,N_16441,N_16119);
or U21191 (N_21191,N_18685,N_15849);
or U21192 (N_21192,N_18073,N_15785);
and U21193 (N_21193,N_18518,N_17523);
xnor U21194 (N_21194,N_18394,N_15753);
and U21195 (N_21195,N_17518,N_16187);
nor U21196 (N_21196,N_18050,N_17932);
or U21197 (N_21197,N_18630,N_16035);
nand U21198 (N_21198,N_16575,N_16015);
nand U21199 (N_21199,N_17362,N_15708);
and U21200 (N_21200,N_16561,N_18204);
nand U21201 (N_21201,N_16019,N_17957);
and U21202 (N_21202,N_17144,N_16245);
or U21203 (N_21203,N_16109,N_16660);
xnor U21204 (N_21204,N_16114,N_15988);
xor U21205 (N_21205,N_18018,N_17420);
nand U21206 (N_21206,N_15702,N_16245);
and U21207 (N_21207,N_16839,N_17243);
nand U21208 (N_21208,N_17636,N_17739);
nand U21209 (N_21209,N_17816,N_17924);
or U21210 (N_21210,N_18158,N_16510);
or U21211 (N_21211,N_17476,N_18137);
or U21212 (N_21212,N_16981,N_16686);
nand U21213 (N_21213,N_17968,N_17796);
nor U21214 (N_21214,N_16681,N_17293);
xnor U21215 (N_21215,N_16724,N_17065);
xor U21216 (N_21216,N_18707,N_17271);
and U21217 (N_21217,N_18133,N_17474);
nand U21218 (N_21218,N_18433,N_17646);
nor U21219 (N_21219,N_18355,N_17588);
xor U21220 (N_21220,N_17325,N_18438);
or U21221 (N_21221,N_17364,N_17931);
or U21222 (N_21222,N_17286,N_18103);
and U21223 (N_21223,N_17769,N_16205);
and U21224 (N_21224,N_16953,N_17402);
xor U21225 (N_21225,N_17315,N_17419);
nor U21226 (N_21226,N_15714,N_18210);
or U21227 (N_21227,N_18141,N_16876);
xnor U21228 (N_21228,N_18719,N_17015);
nand U21229 (N_21229,N_16780,N_16944);
nand U21230 (N_21230,N_18113,N_17837);
xnor U21231 (N_21231,N_18616,N_17018);
and U21232 (N_21232,N_16491,N_16892);
xnor U21233 (N_21233,N_16324,N_16097);
and U21234 (N_21234,N_16628,N_16437);
and U21235 (N_21235,N_18632,N_16442);
xnor U21236 (N_21236,N_17363,N_15686);
nor U21237 (N_21237,N_16529,N_17802);
and U21238 (N_21238,N_16876,N_16442);
nor U21239 (N_21239,N_17210,N_18417);
xnor U21240 (N_21240,N_16666,N_17761);
or U21241 (N_21241,N_16710,N_18600);
or U21242 (N_21242,N_17352,N_17586);
xnor U21243 (N_21243,N_17570,N_16320);
and U21244 (N_21244,N_16843,N_17512);
nand U21245 (N_21245,N_16815,N_17895);
xor U21246 (N_21246,N_16541,N_17919);
nand U21247 (N_21247,N_17348,N_16106);
or U21248 (N_21248,N_18651,N_16003);
nand U21249 (N_21249,N_16258,N_15706);
nor U21250 (N_21250,N_16089,N_16873);
or U21251 (N_21251,N_16660,N_17361);
or U21252 (N_21252,N_17218,N_16796);
nand U21253 (N_21253,N_18570,N_17586);
xnor U21254 (N_21254,N_18252,N_18738);
and U21255 (N_21255,N_15779,N_16079);
xnor U21256 (N_21256,N_16107,N_17628);
xnor U21257 (N_21257,N_17417,N_15635);
nor U21258 (N_21258,N_18353,N_16228);
xor U21259 (N_21259,N_16675,N_18670);
and U21260 (N_21260,N_17865,N_17182);
and U21261 (N_21261,N_16731,N_17098);
nand U21262 (N_21262,N_15923,N_17086);
nand U21263 (N_21263,N_18635,N_17600);
nor U21264 (N_21264,N_17102,N_15784);
nand U21265 (N_21265,N_17526,N_15919);
nor U21266 (N_21266,N_16762,N_16595);
xnor U21267 (N_21267,N_18659,N_16596);
and U21268 (N_21268,N_16547,N_15866);
xnor U21269 (N_21269,N_15891,N_16173);
or U21270 (N_21270,N_16666,N_17215);
nand U21271 (N_21271,N_17215,N_17379);
xnor U21272 (N_21272,N_17742,N_18203);
nand U21273 (N_21273,N_17225,N_18649);
and U21274 (N_21274,N_17477,N_18632);
nor U21275 (N_21275,N_16765,N_17631);
or U21276 (N_21276,N_16750,N_18016);
xnor U21277 (N_21277,N_16185,N_17166);
xor U21278 (N_21278,N_16198,N_18367);
or U21279 (N_21279,N_17096,N_18640);
or U21280 (N_21280,N_16903,N_18497);
nor U21281 (N_21281,N_17205,N_17035);
nand U21282 (N_21282,N_15714,N_17186);
nand U21283 (N_21283,N_17871,N_16894);
nor U21284 (N_21284,N_18468,N_17535);
xor U21285 (N_21285,N_17268,N_17542);
nor U21286 (N_21286,N_16823,N_17694);
nand U21287 (N_21287,N_15869,N_15630);
xnor U21288 (N_21288,N_17727,N_16623);
or U21289 (N_21289,N_16964,N_16513);
or U21290 (N_21290,N_18217,N_16362);
nor U21291 (N_21291,N_18407,N_17545);
nand U21292 (N_21292,N_16539,N_16163);
nand U21293 (N_21293,N_16416,N_16934);
nor U21294 (N_21294,N_16029,N_18543);
nand U21295 (N_21295,N_17062,N_16039);
and U21296 (N_21296,N_16866,N_16886);
nand U21297 (N_21297,N_15985,N_17392);
nor U21298 (N_21298,N_15645,N_16853);
xor U21299 (N_21299,N_15704,N_17764);
nor U21300 (N_21300,N_17881,N_17994);
and U21301 (N_21301,N_16441,N_17212);
and U21302 (N_21302,N_16574,N_17646);
nand U21303 (N_21303,N_16457,N_17824);
nand U21304 (N_21304,N_17371,N_18184);
nand U21305 (N_21305,N_18523,N_16239);
nor U21306 (N_21306,N_15632,N_17524);
nor U21307 (N_21307,N_18595,N_17013);
xnor U21308 (N_21308,N_15695,N_15706);
nor U21309 (N_21309,N_15837,N_17165);
nor U21310 (N_21310,N_17728,N_17680);
nor U21311 (N_21311,N_17864,N_16314);
xor U21312 (N_21312,N_17687,N_16805);
and U21313 (N_21313,N_18032,N_17902);
xnor U21314 (N_21314,N_17611,N_18225);
nor U21315 (N_21315,N_18129,N_17251);
xnor U21316 (N_21316,N_16493,N_16717);
xor U21317 (N_21317,N_17888,N_18348);
and U21318 (N_21318,N_17831,N_18501);
nand U21319 (N_21319,N_16454,N_15913);
nand U21320 (N_21320,N_17259,N_17684);
nor U21321 (N_21321,N_18579,N_16164);
or U21322 (N_21322,N_17880,N_16395);
or U21323 (N_21323,N_16883,N_16562);
or U21324 (N_21324,N_16531,N_16843);
and U21325 (N_21325,N_16376,N_16571);
nor U21326 (N_21326,N_17910,N_16383);
nand U21327 (N_21327,N_16295,N_16847);
nand U21328 (N_21328,N_18319,N_16535);
xnor U21329 (N_21329,N_15723,N_16493);
or U21330 (N_21330,N_16955,N_16612);
xnor U21331 (N_21331,N_16323,N_16343);
nand U21332 (N_21332,N_15916,N_17194);
nor U21333 (N_21333,N_16068,N_18387);
xor U21334 (N_21334,N_18478,N_18505);
xor U21335 (N_21335,N_17128,N_18525);
xnor U21336 (N_21336,N_17318,N_17433);
nor U21337 (N_21337,N_17074,N_16304);
and U21338 (N_21338,N_17208,N_18054);
nor U21339 (N_21339,N_15872,N_16135);
nand U21340 (N_21340,N_18699,N_17323);
xnor U21341 (N_21341,N_16236,N_17013);
or U21342 (N_21342,N_15710,N_18610);
nor U21343 (N_21343,N_15949,N_17296);
nor U21344 (N_21344,N_17278,N_16623);
or U21345 (N_21345,N_16678,N_15683);
xnor U21346 (N_21346,N_18303,N_15712);
and U21347 (N_21347,N_16791,N_16353);
and U21348 (N_21348,N_17598,N_15866);
and U21349 (N_21349,N_18098,N_16355);
or U21350 (N_21350,N_17837,N_18465);
nand U21351 (N_21351,N_16277,N_18613);
or U21352 (N_21352,N_17077,N_16634);
and U21353 (N_21353,N_16963,N_16038);
nor U21354 (N_21354,N_15965,N_15979);
nand U21355 (N_21355,N_18519,N_17713);
or U21356 (N_21356,N_18370,N_15683);
nand U21357 (N_21357,N_17702,N_16764);
nor U21358 (N_21358,N_16641,N_15815);
or U21359 (N_21359,N_16540,N_18538);
nand U21360 (N_21360,N_17538,N_15961);
or U21361 (N_21361,N_16762,N_17713);
nor U21362 (N_21362,N_16296,N_18232);
nor U21363 (N_21363,N_16557,N_17304);
nand U21364 (N_21364,N_17885,N_18482);
nor U21365 (N_21365,N_16218,N_16372);
or U21366 (N_21366,N_18301,N_15822);
or U21367 (N_21367,N_18111,N_15846);
nand U21368 (N_21368,N_16468,N_17183);
and U21369 (N_21369,N_17587,N_17961);
or U21370 (N_21370,N_18694,N_18101);
and U21371 (N_21371,N_16151,N_17303);
or U21372 (N_21372,N_15973,N_17512);
nand U21373 (N_21373,N_17128,N_16537);
and U21374 (N_21374,N_16074,N_18318);
and U21375 (N_21375,N_18420,N_17065);
nand U21376 (N_21376,N_16370,N_16971);
xnor U21377 (N_21377,N_18405,N_18264);
nand U21378 (N_21378,N_16962,N_17133);
nor U21379 (N_21379,N_15645,N_16312);
or U21380 (N_21380,N_17132,N_15741);
nor U21381 (N_21381,N_16602,N_15730);
xor U21382 (N_21382,N_18504,N_16774);
nand U21383 (N_21383,N_17152,N_15870);
nor U21384 (N_21384,N_18643,N_18257);
nor U21385 (N_21385,N_18318,N_17285);
xnor U21386 (N_21386,N_16517,N_16774);
or U21387 (N_21387,N_18346,N_15944);
and U21388 (N_21388,N_17441,N_15876);
nand U21389 (N_21389,N_18738,N_17971);
nor U21390 (N_21390,N_17076,N_16692);
xnor U21391 (N_21391,N_18501,N_16361);
or U21392 (N_21392,N_17306,N_16262);
nand U21393 (N_21393,N_18399,N_16400);
nor U21394 (N_21394,N_16584,N_18353);
xnor U21395 (N_21395,N_18463,N_16406);
and U21396 (N_21396,N_15803,N_17011);
nand U21397 (N_21397,N_17624,N_18489);
or U21398 (N_21398,N_16958,N_16974);
nor U21399 (N_21399,N_17900,N_16489);
or U21400 (N_21400,N_17665,N_17829);
nand U21401 (N_21401,N_17526,N_17759);
xor U21402 (N_21402,N_16740,N_17548);
xor U21403 (N_21403,N_16166,N_17759);
nand U21404 (N_21404,N_18230,N_16445);
nor U21405 (N_21405,N_18631,N_16538);
nand U21406 (N_21406,N_18289,N_17383);
or U21407 (N_21407,N_17545,N_15698);
nand U21408 (N_21408,N_17579,N_17144);
and U21409 (N_21409,N_18538,N_17228);
xor U21410 (N_21410,N_15712,N_15811);
nor U21411 (N_21411,N_17543,N_17878);
or U21412 (N_21412,N_17457,N_18227);
nand U21413 (N_21413,N_16575,N_18076);
nand U21414 (N_21414,N_17833,N_17522);
and U21415 (N_21415,N_16793,N_18000);
and U21416 (N_21416,N_16624,N_17162);
xnor U21417 (N_21417,N_16828,N_16444);
xor U21418 (N_21418,N_16786,N_17256);
xnor U21419 (N_21419,N_17014,N_17543);
xor U21420 (N_21420,N_18261,N_18529);
xnor U21421 (N_21421,N_18080,N_16796);
and U21422 (N_21422,N_16631,N_18362);
and U21423 (N_21423,N_17365,N_16339);
nand U21424 (N_21424,N_17679,N_18735);
xor U21425 (N_21425,N_17969,N_16512);
and U21426 (N_21426,N_17488,N_15792);
and U21427 (N_21427,N_16354,N_16770);
xnor U21428 (N_21428,N_17829,N_18279);
or U21429 (N_21429,N_17959,N_17810);
xnor U21430 (N_21430,N_15713,N_17377);
and U21431 (N_21431,N_17306,N_18426);
or U21432 (N_21432,N_16935,N_15735);
or U21433 (N_21433,N_17036,N_16152);
or U21434 (N_21434,N_16929,N_18234);
xnor U21435 (N_21435,N_16738,N_16028);
xor U21436 (N_21436,N_17443,N_17687);
nand U21437 (N_21437,N_16778,N_16131);
nand U21438 (N_21438,N_18107,N_17592);
xor U21439 (N_21439,N_15939,N_18128);
nand U21440 (N_21440,N_16866,N_16057);
nor U21441 (N_21441,N_16585,N_17367);
or U21442 (N_21442,N_18447,N_17348);
nand U21443 (N_21443,N_17086,N_16195);
nand U21444 (N_21444,N_17432,N_17919);
or U21445 (N_21445,N_18138,N_17714);
nor U21446 (N_21446,N_16708,N_17452);
and U21447 (N_21447,N_17096,N_18575);
nand U21448 (N_21448,N_18111,N_15775);
nand U21449 (N_21449,N_18182,N_18205);
or U21450 (N_21450,N_17356,N_17475);
and U21451 (N_21451,N_15993,N_17005);
or U21452 (N_21452,N_15808,N_18390);
and U21453 (N_21453,N_18682,N_18245);
nor U21454 (N_21454,N_15907,N_17361);
or U21455 (N_21455,N_16987,N_17478);
nand U21456 (N_21456,N_16908,N_18223);
nor U21457 (N_21457,N_16903,N_16776);
nor U21458 (N_21458,N_18563,N_17701);
xnor U21459 (N_21459,N_17549,N_16722);
xnor U21460 (N_21460,N_16276,N_16058);
xor U21461 (N_21461,N_16661,N_17878);
and U21462 (N_21462,N_16305,N_18332);
xnor U21463 (N_21463,N_16482,N_17975);
xor U21464 (N_21464,N_15720,N_17462);
and U21465 (N_21465,N_17477,N_16571);
and U21466 (N_21466,N_18677,N_18732);
or U21467 (N_21467,N_17723,N_18267);
or U21468 (N_21468,N_17856,N_17124);
nand U21469 (N_21469,N_18660,N_18423);
xnor U21470 (N_21470,N_17670,N_15999);
or U21471 (N_21471,N_18114,N_18638);
nor U21472 (N_21472,N_18647,N_17361);
nor U21473 (N_21473,N_17768,N_17550);
and U21474 (N_21474,N_17614,N_17413);
and U21475 (N_21475,N_17582,N_17062);
xor U21476 (N_21476,N_15896,N_15648);
nor U21477 (N_21477,N_18192,N_16520);
and U21478 (N_21478,N_15995,N_16395);
nor U21479 (N_21479,N_17641,N_17036);
nand U21480 (N_21480,N_18171,N_18532);
xnor U21481 (N_21481,N_18193,N_17187);
nor U21482 (N_21482,N_16193,N_17117);
xor U21483 (N_21483,N_18115,N_17392);
nor U21484 (N_21484,N_18471,N_17263);
nor U21485 (N_21485,N_17832,N_16323);
nor U21486 (N_21486,N_18422,N_17821);
and U21487 (N_21487,N_16848,N_18179);
nor U21488 (N_21488,N_16108,N_18549);
or U21489 (N_21489,N_16072,N_17735);
nor U21490 (N_21490,N_16986,N_16710);
nor U21491 (N_21491,N_17991,N_17813);
nand U21492 (N_21492,N_17702,N_15721);
xnor U21493 (N_21493,N_17984,N_17700);
xor U21494 (N_21494,N_17810,N_18494);
xnor U21495 (N_21495,N_17852,N_15755);
or U21496 (N_21496,N_16281,N_16538);
nor U21497 (N_21497,N_18532,N_16617);
nor U21498 (N_21498,N_18036,N_16066);
or U21499 (N_21499,N_16118,N_16716);
nor U21500 (N_21500,N_17401,N_16132);
nor U21501 (N_21501,N_18724,N_16869);
and U21502 (N_21502,N_15780,N_17483);
nand U21503 (N_21503,N_18076,N_18051);
or U21504 (N_21504,N_17660,N_16604);
xor U21505 (N_21505,N_17920,N_17605);
and U21506 (N_21506,N_16818,N_16914);
or U21507 (N_21507,N_17527,N_16037);
and U21508 (N_21508,N_16400,N_17296);
xor U21509 (N_21509,N_17116,N_16659);
and U21510 (N_21510,N_15719,N_17719);
and U21511 (N_21511,N_17034,N_16248);
and U21512 (N_21512,N_17320,N_18555);
nor U21513 (N_21513,N_18642,N_17104);
xnor U21514 (N_21514,N_16946,N_17473);
nand U21515 (N_21515,N_17547,N_17335);
nor U21516 (N_21516,N_18181,N_17379);
xor U21517 (N_21517,N_18357,N_17064);
and U21518 (N_21518,N_17702,N_17359);
and U21519 (N_21519,N_17312,N_18507);
or U21520 (N_21520,N_15784,N_17281);
xnor U21521 (N_21521,N_17831,N_16476);
and U21522 (N_21522,N_16419,N_16468);
xor U21523 (N_21523,N_15765,N_16902);
or U21524 (N_21524,N_17449,N_18476);
or U21525 (N_21525,N_17222,N_17457);
and U21526 (N_21526,N_18297,N_17069);
or U21527 (N_21527,N_17777,N_15725);
and U21528 (N_21528,N_17093,N_16490);
nand U21529 (N_21529,N_18748,N_18028);
nor U21530 (N_21530,N_17718,N_17056);
nor U21531 (N_21531,N_17904,N_18051);
nor U21532 (N_21532,N_18171,N_15807);
nor U21533 (N_21533,N_18584,N_17597);
or U21534 (N_21534,N_16808,N_16698);
and U21535 (N_21535,N_16933,N_15775);
and U21536 (N_21536,N_18223,N_18161);
and U21537 (N_21537,N_17812,N_16155);
xor U21538 (N_21538,N_16464,N_17738);
or U21539 (N_21539,N_18052,N_17784);
nor U21540 (N_21540,N_16947,N_16965);
xor U21541 (N_21541,N_16935,N_16677);
nor U21542 (N_21542,N_16240,N_17148);
xnor U21543 (N_21543,N_16118,N_16348);
nor U21544 (N_21544,N_18385,N_17374);
or U21545 (N_21545,N_16927,N_18588);
nand U21546 (N_21546,N_18085,N_18193);
nor U21547 (N_21547,N_17358,N_15891);
and U21548 (N_21548,N_16354,N_15877);
nand U21549 (N_21549,N_15882,N_16428);
or U21550 (N_21550,N_18654,N_18547);
and U21551 (N_21551,N_16487,N_15979);
or U21552 (N_21552,N_16777,N_18159);
nand U21553 (N_21553,N_16314,N_15853);
nand U21554 (N_21554,N_16376,N_16468);
nor U21555 (N_21555,N_16104,N_17252);
or U21556 (N_21556,N_16393,N_18500);
and U21557 (N_21557,N_17529,N_15779);
nand U21558 (N_21558,N_17317,N_16088);
and U21559 (N_21559,N_15937,N_17518);
nor U21560 (N_21560,N_17209,N_16509);
nor U21561 (N_21561,N_15667,N_18212);
or U21562 (N_21562,N_17097,N_18267);
nor U21563 (N_21563,N_16126,N_16534);
xor U21564 (N_21564,N_18065,N_16795);
or U21565 (N_21565,N_16026,N_17297);
nand U21566 (N_21566,N_18698,N_15721);
and U21567 (N_21567,N_15926,N_18192);
or U21568 (N_21568,N_17278,N_18192);
nor U21569 (N_21569,N_18386,N_18264);
and U21570 (N_21570,N_18212,N_16486);
or U21571 (N_21571,N_18095,N_16646);
xor U21572 (N_21572,N_16399,N_16432);
xor U21573 (N_21573,N_17204,N_16533);
and U21574 (N_21574,N_16643,N_16950);
nor U21575 (N_21575,N_16357,N_17971);
nor U21576 (N_21576,N_17078,N_16894);
or U21577 (N_21577,N_16526,N_15801);
and U21578 (N_21578,N_16132,N_16147);
or U21579 (N_21579,N_16574,N_16812);
and U21580 (N_21580,N_15793,N_18437);
and U21581 (N_21581,N_16756,N_17579);
xor U21582 (N_21582,N_15779,N_18159);
nand U21583 (N_21583,N_17393,N_18314);
and U21584 (N_21584,N_17682,N_17779);
nand U21585 (N_21585,N_16217,N_18395);
nand U21586 (N_21586,N_18115,N_15926);
nor U21587 (N_21587,N_15720,N_16365);
or U21588 (N_21588,N_15647,N_17864);
and U21589 (N_21589,N_18201,N_17976);
xor U21590 (N_21590,N_15844,N_17284);
nor U21591 (N_21591,N_18555,N_17725);
xnor U21592 (N_21592,N_18093,N_16853);
or U21593 (N_21593,N_18439,N_18021);
xor U21594 (N_21594,N_18406,N_17920);
nor U21595 (N_21595,N_17474,N_18011);
and U21596 (N_21596,N_17799,N_15933);
or U21597 (N_21597,N_16634,N_17253);
nand U21598 (N_21598,N_18097,N_18678);
xnor U21599 (N_21599,N_18060,N_18555);
or U21600 (N_21600,N_16675,N_16836);
or U21601 (N_21601,N_18328,N_18107);
xor U21602 (N_21602,N_18052,N_16913);
and U21603 (N_21603,N_15927,N_17524);
or U21604 (N_21604,N_18267,N_18098);
nor U21605 (N_21605,N_15704,N_17634);
or U21606 (N_21606,N_17440,N_17605);
xor U21607 (N_21607,N_18322,N_15641);
or U21608 (N_21608,N_17934,N_16813);
nor U21609 (N_21609,N_18732,N_17812);
and U21610 (N_21610,N_18613,N_17391);
nand U21611 (N_21611,N_18321,N_16198);
nor U21612 (N_21612,N_17944,N_17713);
xnor U21613 (N_21613,N_17504,N_15757);
or U21614 (N_21614,N_16041,N_17994);
nor U21615 (N_21615,N_18618,N_15643);
or U21616 (N_21616,N_16623,N_15685);
nor U21617 (N_21617,N_16276,N_15693);
nand U21618 (N_21618,N_15775,N_18648);
nand U21619 (N_21619,N_17544,N_16320);
or U21620 (N_21620,N_17746,N_16202);
nand U21621 (N_21621,N_18289,N_18133);
and U21622 (N_21622,N_17630,N_18151);
xor U21623 (N_21623,N_16259,N_18120);
xnor U21624 (N_21624,N_16816,N_17296);
nand U21625 (N_21625,N_15978,N_17959);
nand U21626 (N_21626,N_17831,N_18738);
and U21627 (N_21627,N_16822,N_17276);
and U21628 (N_21628,N_15886,N_15911);
and U21629 (N_21629,N_16717,N_17871);
or U21630 (N_21630,N_18522,N_17427);
and U21631 (N_21631,N_16084,N_17529);
nor U21632 (N_21632,N_16928,N_16566);
and U21633 (N_21633,N_16448,N_17828);
nand U21634 (N_21634,N_17896,N_18525);
and U21635 (N_21635,N_16624,N_15844);
nor U21636 (N_21636,N_16541,N_17082);
and U21637 (N_21637,N_16214,N_18680);
nor U21638 (N_21638,N_17763,N_16422);
or U21639 (N_21639,N_16120,N_17108);
nand U21640 (N_21640,N_16671,N_16648);
nand U21641 (N_21641,N_18462,N_17748);
nand U21642 (N_21642,N_15972,N_18334);
nand U21643 (N_21643,N_16621,N_15716);
or U21644 (N_21644,N_17702,N_18306);
nand U21645 (N_21645,N_17317,N_18638);
or U21646 (N_21646,N_18081,N_16759);
or U21647 (N_21647,N_17222,N_18058);
xnor U21648 (N_21648,N_17297,N_18160);
and U21649 (N_21649,N_16947,N_17107);
nor U21650 (N_21650,N_17906,N_18371);
nand U21651 (N_21651,N_18523,N_15788);
xor U21652 (N_21652,N_16403,N_17498);
or U21653 (N_21653,N_17003,N_16710);
nand U21654 (N_21654,N_16009,N_18727);
or U21655 (N_21655,N_17571,N_17860);
nand U21656 (N_21656,N_18551,N_18078);
or U21657 (N_21657,N_16166,N_18215);
nand U21658 (N_21658,N_18737,N_18613);
or U21659 (N_21659,N_17260,N_17953);
and U21660 (N_21660,N_18553,N_16770);
nand U21661 (N_21661,N_18382,N_16810);
and U21662 (N_21662,N_16551,N_17356);
xor U21663 (N_21663,N_16724,N_16219);
or U21664 (N_21664,N_17875,N_16988);
or U21665 (N_21665,N_16808,N_18133);
and U21666 (N_21666,N_17109,N_16738);
or U21667 (N_21667,N_17080,N_16835);
nand U21668 (N_21668,N_18489,N_17732);
or U21669 (N_21669,N_16519,N_18542);
xor U21670 (N_21670,N_16269,N_18647);
xor U21671 (N_21671,N_18579,N_15711);
nand U21672 (N_21672,N_17340,N_15909);
nor U21673 (N_21673,N_17449,N_15660);
xor U21674 (N_21674,N_15628,N_16081);
xnor U21675 (N_21675,N_18586,N_16377);
xor U21676 (N_21676,N_18531,N_16891);
or U21677 (N_21677,N_16697,N_15822);
or U21678 (N_21678,N_15827,N_17493);
nand U21679 (N_21679,N_17570,N_16381);
nor U21680 (N_21680,N_18491,N_16295);
xnor U21681 (N_21681,N_18613,N_16137);
or U21682 (N_21682,N_17204,N_15941);
and U21683 (N_21683,N_16328,N_18116);
and U21684 (N_21684,N_18106,N_16252);
xnor U21685 (N_21685,N_17754,N_15836);
or U21686 (N_21686,N_17260,N_18518);
nand U21687 (N_21687,N_15853,N_18125);
and U21688 (N_21688,N_18443,N_18739);
nand U21689 (N_21689,N_18076,N_16299);
nand U21690 (N_21690,N_17047,N_15817);
xnor U21691 (N_21691,N_17238,N_15755);
or U21692 (N_21692,N_18351,N_18042);
nor U21693 (N_21693,N_16307,N_17047);
xnor U21694 (N_21694,N_16369,N_16752);
xnor U21695 (N_21695,N_16323,N_18676);
nor U21696 (N_21696,N_16643,N_15727);
nand U21697 (N_21697,N_17817,N_16327);
nand U21698 (N_21698,N_18702,N_18422);
and U21699 (N_21699,N_18575,N_17054);
and U21700 (N_21700,N_18520,N_17045);
and U21701 (N_21701,N_16608,N_17018);
and U21702 (N_21702,N_18227,N_16059);
and U21703 (N_21703,N_17703,N_16143);
nand U21704 (N_21704,N_15884,N_18205);
or U21705 (N_21705,N_17722,N_17235);
nand U21706 (N_21706,N_18592,N_16882);
or U21707 (N_21707,N_16674,N_17545);
nand U21708 (N_21708,N_18364,N_16923);
xor U21709 (N_21709,N_18749,N_16004);
or U21710 (N_21710,N_16090,N_17374);
nor U21711 (N_21711,N_15638,N_18066);
nand U21712 (N_21712,N_17426,N_16306);
or U21713 (N_21713,N_15663,N_18580);
nor U21714 (N_21714,N_15726,N_16205);
nor U21715 (N_21715,N_15818,N_17888);
and U21716 (N_21716,N_16693,N_18354);
and U21717 (N_21717,N_18340,N_17056);
or U21718 (N_21718,N_17236,N_18079);
nor U21719 (N_21719,N_16924,N_16839);
nand U21720 (N_21720,N_18484,N_15897);
nand U21721 (N_21721,N_18644,N_16777);
and U21722 (N_21722,N_16216,N_17336);
and U21723 (N_21723,N_15694,N_16187);
xnor U21724 (N_21724,N_15798,N_15939);
nor U21725 (N_21725,N_17812,N_16412);
or U21726 (N_21726,N_17322,N_17679);
nor U21727 (N_21727,N_17288,N_15864);
and U21728 (N_21728,N_18596,N_18172);
nand U21729 (N_21729,N_15910,N_17845);
and U21730 (N_21730,N_17476,N_17380);
xnor U21731 (N_21731,N_18153,N_17942);
or U21732 (N_21732,N_16016,N_16594);
xor U21733 (N_21733,N_15747,N_16084);
nand U21734 (N_21734,N_17977,N_16980);
nand U21735 (N_21735,N_16129,N_16328);
or U21736 (N_21736,N_18497,N_18329);
nor U21737 (N_21737,N_16594,N_15853);
nand U21738 (N_21738,N_16881,N_18665);
or U21739 (N_21739,N_16820,N_18261);
nor U21740 (N_21740,N_16183,N_17927);
nor U21741 (N_21741,N_18571,N_18103);
nand U21742 (N_21742,N_16541,N_17173);
xor U21743 (N_21743,N_17059,N_17891);
or U21744 (N_21744,N_16899,N_15984);
and U21745 (N_21745,N_18713,N_17149);
nand U21746 (N_21746,N_16162,N_16317);
and U21747 (N_21747,N_18029,N_17281);
xnor U21748 (N_21748,N_16982,N_16947);
and U21749 (N_21749,N_16582,N_18101);
nand U21750 (N_21750,N_15885,N_15916);
or U21751 (N_21751,N_16180,N_17264);
nor U21752 (N_21752,N_17557,N_18548);
or U21753 (N_21753,N_18634,N_17372);
xnor U21754 (N_21754,N_18118,N_17902);
xor U21755 (N_21755,N_17812,N_16851);
or U21756 (N_21756,N_17400,N_16639);
xnor U21757 (N_21757,N_18313,N_18065);
and U21758 (N_21758,N_17524,N_18392);
or U21759 (N_21759,N_18186,N_15884);
or U21760 (N_21760,N_17368,N_17631);
nand U21761 (N_21761,N_18067,N_18544);
xor U21762 (N_21762,N_17630,N_17793);
or U21763 (N_21763,N_18720,N_17294);
or U21764 (N_21764,N_17909,N_16713);
nand U21765 (N_21765,N_16352,N_17260);
and U21766 (N_21766,N_17961,N_17437);
and U21767 (N_21767,N_16613,N_17138);
or U21768 (N_21768,N_17222,N_17085);
and U21769 (N_21769,N_18376,N_16534);
or U21770 (N_21770,N_17786,N_16121);
nand U21771 (N_21771,N_16654,N_16467);
nor U21772 (N_21772,N_15978,N_16073);
nor U21773 (N_21773,N_15986,N_18299);
and U21774 (N_21774,N_16395,N_17229);
nand U21775 (N_21775,N_15698,N_18623);
nand U21776 (N_21776,N_16761,N_18411);
xor U21777 (N_21777,N_17205,N_18657);
and U21778 (N_21778,N_16075,N_18619);
nor U21779 (N_21779,N_16557,N_17238);
nand U21780 (N_21780,N_17470,N_16821);
and U21781 (N_21781,N_16529,N_15694);
and U21782 (N_21782,N_17754,N_18050);
or U21783 (N_21783,N_17764,N_16276);
nand U21784 (N_21784,N_17245,N_18176);
or U21785 (N_21785,N_17518,N_17033);
xnor U21786 (N_21786,N_16798,N_18039);
xnor U21787 (N_21787,N_17485,N_15999);
nand U21788 (N_21788,N_17072,N_18203);
or U21789 (N_21789,N_16201,N_18482);
nor U21790 (N_21790,N_16637,N_18566);
and U21791 (N_21791,N_18685,N_17258);
or U21792 (N_21792,N_17344,N_17087);
or U21793 (N_21793,N_18459,N_15778);
and U21794 (N_21794,N_16723,N_15950);
and U21795 (N_21795,N_16255,N_18163);
xor U21796 (N_21796,N_18327,N_16776);
nor U21797 (N_21797,N_18120,N_17347);
xor U21798 (N_21798,N_16268,N_17695);
xnor U21799 (N_21799,N_16779,N_16226);
and U21800 (N_21800,N_15679,N_16525);
nand U21801 (N_21801,N_16478,N_16238);
and U21802 (N_21802,N_16283,N_16291);
nand U21803 (N_21803,N_17282,N_15714);
and U21804 (N_21804,N_16484,N_18113);
or U21805 (N_21805,N_18693,N_18744);
nand U21806 (N_21806,N_15651,N_18575);
xor U21807 (N_21807,N_17424,N_16731);
nand U21808 (N_21808,N_17792,N_16388);
nor U21809 (N_21809,N_17347,N_18469);
or U21810 (N_21810,N_16194,N_15922);
or U21811 (N_21811,N_16100,N_18593);
xor U21812 (N_21812,N_16618,N_18507);
nor U21813 (N_21813,N_15965,N_16842);
and U21814 (N_21814,N_17146,N_16994);
xor U21815 (N_21815,N_15755,N_17964);
nand U21816 (N_21816,N_17241,N_18711);
and U21817 (N_21817,N_17924,N_17139);
xnor U21818 (N_21818,N_18457,N_16095);
nand U21819 (N_21819,N_18388,N_16947);
and U21820 (N_21820,N_16081,N_16208);
nor U21821 (N_21821,N_16996,N_16385);
or U21822 (N_21822,N_17791,N_17631);
xnor U21823 (N_21823,N_16400,N_17728);
and U21824 (N_21824,N_17262,N_18206);
nand U21825 (N_21825,N_16816,N_15948);
xor U21826 (N_21826,N_18580,N_17558);
xor U21827 (N_21827,N_17580,N_17342);
nor U21828 (N_21828,N_17854,N_17772);
nor U21829 (N_21829,N_17345,N_15872);
and U21830 (N_21830,N_16993,N_16278);
or U21831 (N_21831,N_17609,N_16969);
or U21832 (N_21832,N_17001,N_17004);
nand U21833 (N_21833,N_18453,N_15697);
and U21834 (N_21834,N_17744,N_15953);
nor U21835 (N_21835,N_16129,N_18253);
nand U21836 (N_21836,N_17507,N_18350);
xnor U21837 (N_21837,N_18585,N_15833);
xor U21838 (N_21838,N_18663,N_15795);
or U21839 (N_21839,N_16272,N_16004);
xor U21840 (N_21840,N_17523,N_16287);
or U21841 (N_21841,N_17935,N_17247);
nor U21842 (N_21842,N_17212,N_17145);
nor U21843 (N_21843,N_17173,N_18368);
nand U21844 (N_21844,N_16413,N_17537);
and U21845 (N_21845,N_18062,N_18212);
nor U21846 (N_21846,N_18527,N_17246);
or U21847 (N_21847,N_16837,N_17921);
and U21848 (N_21848,N_16017,N_16306);
or U21849 (N_21849,N_17916,N_18097);
and U21850 (N_21850,N_16504,N_16688);
nor U21851 (N_21851,N_16762,N_15939);
nand U21852 (N_21852,N_16802,N_17284);
or U21853 (N_21853,N_15639,N_17377);
xor U21854 (N_21854,N_18604,N_16236);
xor U21855 (N_21855,N_16691,N_18723);
and U21856 (N_21856,N_17089,N_16281);
nand U21857 (N_21857,N_16111,N_18188);
nand U21858 (N_21858,N_16661,N_17177);
nand U21859 (N_21859,N_15761,N_16442);
nor U21860 (N_21860,N_16949,N_17410);
xnor U21861 (N_21861,N_17270,N_17043);
nor U21862 (N_21862,N_16378,N_17652);
nand U21863 (N_21863,N_15787,N_16212);
and U21864 (N_21864,N_15960,N_16991);
and U21865 (N_21865,N_16529,N_17808);
xor U21866 (N_21866,N_17382,N_17361);
nand U21867 (N_21867,N_18604,N_15859);
nor U21868 (N_21868,N_17029,N_16871);
and U21869 (N_21869,N_16862,N_16380);
nand U21870 (N_21870,N_18393,N_17459);
and U21871 (N_21871,N_16417,N_17886);
or U21872 (N_21872,N_17550,N_17723);
xor U21873 (N_21873,N_17646,N_17455);
and U21874 (N_21874,N_18645,N_18451);
or U21875 (N_21875,N_20849,N_20452);
xor U21876 (N_21876,N_21560,N_18849);
and U21877 (N_21877,N_19700,N_19298);
xnor U21878 (N_21878,N_21671,N_20818);
and U21879 (N_21879,N_18769,N_18880);
xor U21880 (N_21880,N_20722,N_20817);
or U21881 (N_21881,N_21468,N_19390);
and U21882 (N_21882,N_18902,N_19706);
nand U21883 (N_21883,N_19697,N_20512);
and U21884 (N_21884,N_19045,N_20247);
and U21885 (N_21885,N_20243,N_21840);
nor U21886 (N_21886,N_19403,N_19516);
nand U21887 (N_21887,N_20836,N_19432);
and U21888 (N_21888,N_18955,N_21508);
and U21889 (N_21889,N_20059,N_19581);
xnor U21890 (N_21890,N_19209,N_18835);
nand U21891 (N_21891,N_19717,N_19069);
and U21892 (N_21892,N_19551,N_21190);
and U21893 (N_21893,N_20188,N_20414);
xor U21894 (N_21894,N_18804,N_20946);
and U21895 (N_21895,N_19804,N_20474);
nand U21896 (N_21896,N_21013,N_18855);
nor U21897 (N_21897,N_19994,N_21293);
and U21898 (N_21898,N_20829,N_20027);
or U21899 (N_21899,N_19903,N_21309);
and U21900 (N_21900,N_21195,N_20528);
nand U21901 (N_21901,N_20736,N_21786);
and U21902 (N_21902,N_21062,N_18911);
xor U21903 (N_21903,N_19479,N_18825);
or U21904 (N_21904,N_20403,N_19875);
or U21905 (N_21905,N_19812,N_21721);
nor U21906 (N_21906,N_20071,N_19671);
nor U21907 (N_21907,N_20886,N_20412);
and U21908 (N_21908,N_19270,N_21594);
xnor U21909 (N_21909,N_19984,N_18999);
nor U21910 (N_21910,N_19441,N_19970);
and U21911 (N_21911,N_19594,N_20928);
nand U21912 (N_21912,N_21718,N_18973);
and U21913 (N_21913,N_20418,N_20563);
and U21914 (N_21914,N_18815,N_21524);
nand U21915 (N_21915,N_19330,N_20174);
and U21916 (N_21916,N_20982,N_19019);
or U21917 (N_21917,N_21503,N_20601);
or U21918 (N_21918,N_20715,N_19345);
or U21919 (N_21919,N_19016,N_18766);
nor U21920 (N_21920,N_19112,N_21868);
nand U21921 (N_21921,N_21550,N_20887);
nor U21922 (N_21922,N_21192,N_20094);
xor U21923 (N_21923,N_20519,N_21079);
or U21924 (N_21924,N_19549,N_20926);
or U21925 (N_21925,N_20054,N_21541);
or U21926 (N_21926,N_21490,N_19872);
xnor U21927 (N_21927,N_21326,N_19187);
nand U21928 (N_21928,N_19325,N_21830);
nand U21929 (N_21929,N_19603,N_21793);
nor U21930 (N_21930,N_19078,N_20822);
and U21931 (N_21931,N_21536,N_21675);
nor U21932 (N_21932,N_20402,N_20776);
nor U21933 (N_21933,N_21015,N_18957);
or U21934 (N_21934,N_19795,N_20870);
and U21935 (N_21935,N_21530,N_20043);
or U21936 (N_21936,N_20156,N_21331);
nand U21937 (N_21937,N_19997,N_19742);
and U21938 (N_21938,N_20202,N_21515);
or U21939 (N_21939,N_21211,N_21574);
xor U21940 (N_21940,N_21736,N_21225);
nand U21941 (N_21941,N_19553,N_20598);
or U21942 (N_21942,N_21040,N_20303);
and U21943 (N_21943,N_21308,N_19168);
nand U21944 (N_21944,N_20577,N_19393);
nand U21945 (N_21945,N_21411,N_19021);
xor U21946 (N_21946,N_19018,N_21083);
nand U21947 (N_21947,N_21425,N_21036);
and U21948 (N_21948,N_21858,N_19362);
nor U21949 (N_21949,N_19965,N_21837);
or U21950 (N_21950,N_21711,N_19440);
or U21951 (N_21951,N_21813,N_20649);
nor U21952 (N_21952,N_20665,N_19499);
nand U21953 (N_21953,N_18762,N_21029);
and U21954 (N_21954,N_21654,N_21733);
nand U21955 (N_21955,N_19445,N_20718);
nor U21956 (N_21956,N_21754,N_20237);
nand U21957 (N_21957,N_19975,N_20793);
and U21958 (N_21958,N_21204,N_21597);
xnor U21959 (N_21959,N_20292,N_21621);
or U21960 (N_21960,N_20786,N_20281);
xor U21961 (N_21961,N_18851,N_19121);
xnor U21962 (N_21962,N_21347,N_21471);
nand U21963 (N_21963,N_19958,N_19250);
and U21964 (N_21964,N_21239,N_19404);
nand U21965 (N_21965,N_19331,N_19099);
xnor U21966 (N_21966,N_19686,N_19025);
nor U21967 (N_21967,N_19720,N_20175);
and U21968 (N_21968,N_21473,N_21410);
xnor U21969 (N_21969,N_19847,N_20290);
or U21970 (N_21970,N_19616,N_21361);
and U21971 (N_21971,N_21500,N_21861);
xnor U21972 (N_21972,N_19329,N_19514);
or U21973 (N_21973,N_20002,N_21540);
nand U21974 (N_21974,N_18790,N_21852);
and U21975 (N_21975,N_20666,N_20589);
and U21976 (N_21976,N_20357,N_20972);
nand U21977 (N_21977,N_20834,N_20686);
nor U21978 (N_21978,N_21212,N_21283);
nand U21979 (N_21979,N_20896,N_19973);
xnor U21980 (N_21980,N_21593,N_20398);
nand U21981 (N_21981,N_20255,N_20087);
nor U21982 (N_21982,N_20646,N_21526);
xnor U21983 (N_21983,N_21420,N_20148);
nand U21984 (N_21984,N_20384,N_19027);
xor U21985 (N_21985,N_21244,N_21796);
and U21986 (N_21986,N_21379,N_20510);
xnor U21987 (N_21987,N_20272,N_18822);
nor U21988 (N_21988,N_21340,N_20289);
xnor U21989 (N_21989,N_18939,N_20841);
xor U21990 (N_21990,N_21088,N_21798);
and U21991 (N_21991,N_21205,N_20737);
nand U21992 (N_21992,N_20436,N_19768);
and U21993 (N_21993,N_20074,N_20652);
xnor U21994 (N_21994,N_21517,N_19035);
nand U21995 (N_21995,N_19396,N_20688);
and U21996 (N_21996,N_21185,N_18823);
xnor U21997 (N_21997,N_20101,N_20354);
or U21998 (N_21998,N_20008,N_18863);
xor U21999 (N_21999,N_19119,N_18961);
or U22000 (N_22000,N_20534,N_18960);
xor U22001 (N_22001,N_21601,N_21566);
xor U22002 (N_22002,N_20491,N_21169);
nand U22003 (N_22003,N_19429,N_19370);
xnor U22004 (N_22004,N_19261,N_21563);
nand U22005 (N_22005,N_18892,N_20034);
xnor U22006 (N_22006,N_21787,N_21374);
and U22007 (N_22007,N_19465,N_19899);
and U22008 (N_22008,N_21290,N_21196);
xnor U22009 (N_22009,N_20932,N_20805);
xnor U22010 (N_22010,N_19637,N_21569);
and U22011 (N_22011,N_19456,N_18990);
xnor U22012 (N_22012,N_18874,N_20687);
nor U22013 (N_22013,N_20373,N_20558);
nand U22014 (N_22014,N_19427,N_18967);
and U22015 (N_22015,N_21870,N_19070);
and U22016 (N_22016,N_21071,N_21218);
xnor U22017 (N_22017,N_18765,N_18925);
nand U22018 (N_22018,N_19386,N_18768);
or U22019 (N_22019,N_19013,N_21392);
or U22020 (N_22020,N_20988,N_20544);
and U22021 (N_22021,N_19148,N_20977);
nor U22022 (N_22022,N_21068,N_21737);
and U22023 (N_22023,N_21389,N_19601);
and U22024 (N_22024,N_21806,N_20151);
xnor U22025 (N_22025,N_20518,N_21727);
and U22026 (N_22026,N_21258,N_19780);
xor U22027 (N_22027,N_19234,N_18839);
xnor U22028 (N_22028,N_19416,N_20731);
nand U22029 (N_22029,N_19868,N_19857);
or U22030 (N_22030,N_20604,N_21484);
or U22031 (N_22031,N_21148,N_18982);
nand U22032 (N_22032,N_19494,N_21778);
xor U22033 (N_22033,N_20937,N_21682);
xor U22034 (N_22034,N_19892,N_18884);
or U22035 (N_22035,N_21485,N_19106);
nor U22036 (N_22036,N_19712,N_19472);
nand U22037 (N_22037,N_19764,N_19627);
or U22038 (N_22038,N_21302,N_19898);
or U22039 (N_22039,N_20205,N_18980);
or U22040 (N_22040,N_19424,N_20443);
nor U22041 (N_22041,N_19096,N_20991);
nand U22042 (N_22042,N_19305,N_19876);
xor U22043 (N_22043,N_19798,N_20444);
or U22044 (N_22044,N_20061,N_21208);
or U22045 (N_22045,N_20236,N_20976);
or U22046 (N_22046,N_18778,N_21803);
nor U22047 (N_22047,N_19259,N_19782);
nor U22048 (N_22048,N_21871,N_20322);
xor U22049 (N_22049,N_19587,N_19655);
xnor U22050 (N_22050,N_20949,N_19648);
nand U22051 (N_22051,N_21329,N_18786);
nor U22052 (N_22052,N_20533,N_21241);
or U22053 (N_22053,N_19458,N_21203);
or U22054 (N_22054,N_19446,N_19247);
nand U22055 (N_22055,N_20620,N_18837);
nand U22056 (N_22056,N_19461,N_20249);
xnor U22057 (N_22057,N_19705,N_20233);
nand U22058 (N_22058,N_21305,N_20407);
nand U22059 (N_22059,N_18818,N_21125);
nand U22060 (N_22060,N_20635,N_21081);
and U22061 (N_22061,N_19092,N_21284);
nand U22062 (N_22062,N_20521,N_19090);
nor U22063 (N_22063,N_19274,N_18841);
and U22064 (N_22064,N_20933,N_19038);
nand U22065 (N_22065,N_20192,N_19521);
xnor U22066 (N_22066,N_19232,N_21140);
nor U22067 (N_22067,N_21095,N_19267);
nor U22068 (N_22068,N_19995,N_19545);
nand U22069 (N_22069,N_21470,N_19156);
or U22070 (N_22070,N_19091,N_20241);
nor U22071 (N_22071,N_20593,N_18757);
or U22072 (N_22072,N_20103,N_20750);
nand U22073 (N_22073,N_19583,N_20800);
nor U22074 (N_22074,N_19349,N_21461);
nand U22075 (N_22075,N_19423,N_20930);
xor U22076 (N_22076,N_19029,N_19186);
xnor U22077 (N_22077,N_20531,N_19398);
nor U22078 (N_22078,N_20874,N_20942);
nor U22079 (N_22079,N_19490,N_18983);
xnor U22080 (N_22080,N_20166,N_19867);
and U22081 (N_22081,N_20127,N_18972);
nor U22082 (N_22082,N_20179,N_21367);
and U22083 (N_22083,N_20647,N_19529);
nor U22084 (N_22084,N_19421,N_21055);
xnor U22085 (N_22085,N_18928,N_21653);
xor U22086 (N_22086,N_21514,N_19546);
nand U22087 (N_22087,N_18929,N_20177);
nor U22088 (N_22088,N_21368,N_20807);
and U22089 (N_22089,N_21343,N_19557);
xnor U22090 (N_22090,N_19065,N_19179);
or U22091 (N_22091,N_19877,N_19100);
nand U22092 (N_22092,N_20012,N_21327);
nand U22093 (N_22093,N_19208,N_20803);
and U22094 (N_22094,N_20376,N_21706);
xnor U22095 (N_22095,N_19203,N_19328);
nor U22096 (N_22096,N_21090,N_19149);
nor U22097 (N_22097,N_21557,N_19891);
or U22098 (N_22098,N_19771,N_20456);
xor U22099 (N_22099,N_20015,N_21763);
or U22100 (N_22100,N_21223,N_20092);
xor U22101 (N_22101,N_21679,N_20682);
or U22102 (N_22102,N_21109,N_19881);
nor U22103 (N_22103,N_21131,N_19037);
and U22104 (N_22104,N_19792,N_20337);
xor U22105 (N_22105,N_18787,N_21224);
and U22106 (N_22106,N_21664,N_18801);
and U22107 (N_22107,N_18792,N_20634);
nand U22108 (N_22108,N_18795,N_20910);
nand U22109 (N_22109,N_18881,N_20399);
nor U22110 (N_22110,N_19064,N_19559);
xor U22111 (N_22111,N_19354,N_19218);
nor U22112 (N_22112,N_18989,N_21116);
nand U22113 (N_22113,N_20743,N_19852);
or U22114 (N_22114,N_19944,N_20323);
xor U22115 (N_22115,N_19590,N_20921);
nor U22116 (N_22116,N_21611,N_19348);
xor U22117 (N_22117,N_20216,N_18821);
xnor U22118 (N_22118,N_20908,N_19838);
or U22119 (N_22119,N_18836,N_20245);
xor U22120 (N_22120,N_19911,N_21264);
nand U22121 (N_22121,N_19196,N_18860);
or U22122 (N_22122,N_21547,N_21027);
xor U22123 (N_22123,N_19443,N_20432);
and U22124 (N_22124,N_21720,N_21233);
xnor U22125 (N_22125,N_21623,N_21110);
nor U22126 (N_22126,N_20338,N_19957);
nor U22127 (N_22127,N_18824,N_19871);
nand U22128 (N_22128,N_21427,N_20501);
nor U22129 (N_22129,N_19097,N_21390);
nand U22130 (N_22130,N_19063,N_20833);
xor U22131 (N_22131,N_19579,N_19048);
or U22132 (N_22132,N_21377,N_20111);
xnor U22133 (N_22133,N_21094,N_19605);
or U22134 (N_22134,N_20602,N_20080);
nor U22135 (N_22135,N_21318,N_19762);
nand U22136 (N_22136,N_19139,N_20548);
or U22137 (N_22137,N_18754,N_20696);
nand U22138 (N_22138,N_18949,N_18842);
nor U22139 (N_22139,N_20150,N_18771);
or U22140 (N_22140,N_20324,N_19629);
nor U22141 (N_22141,N_19542,N_20332);
nor U22142 (N_22142,N_21700,N_19055);
nand U22143 (N_22143,N_21455,N_19102);
and U22144 (N_22144,N_20535,N_19310);
and U22145 (N_22145,N_19041,N_20819);
nand U22146 (N_22146,N_18820,N_18913);
xor U22147 (N_22147,N_20614,N_19428);
xnor U22148 (N_22148,N_19816,N_21004);
nand U22149 (N_22149,N_20451,N_19083);
nand U22150 (N_22150,N_20371,N_20215);
nand U22151 (N_22151,N_20542,N_19582);
and U22152 (N_22152,N_21467,N_20405);
nor U22153 (N_22153,N_21638,N_19455);
nor U22154 (N_22154,N_19086,N_21710);
nand U22155 (N_22155,N_19913,N_20306);
and U22156 (N_22156,N_19978,N_20339);
xor U22157 (N_22157,N_20391,N_21435);
nor U22158 (N_22158,N_21122,N_21126);
and U22159 (N_22159,N_20994,N_20137);
and U22160 (N_22160,N_19580,N_21141);
xnor U22161 (N_22161,N_20482,N_21408);
and U22162 (N_22162,N_20437,N_19910);
or U22163 (N_22163,N_20098,N_19785);
xnor U22164 (N_22164,N_21422,N_19089);
nand U22165 (N_22165,N_19547,N_20547);
xor U22166 (N_22166,N_20349,N_20091);
or U22167 (N_22167,N_19111,N_20845);
nand U22168 (N_22168,N_21089,N_20663);
xor U22169 (N_22169,N_20035,N_19578);
nand U22170 (N_22170,N_20507,N_21760);
xnor U22171 (N_22171,N_19945,N_19359);
nand U22172 (N_22172,N_19003,N_18873);
nand U22173 (N_22173,N_19756,N_20782);
or U22174 (N_22174,N_20499,N_19217);
or U22175 (N_22175,N_20107,N_20479);
and U22176 (N_22176,N_19734,N_20721);
xor U22177 (N_22177,N_19220,N_18878);
nor U22178 (N_22178,N_18763,N_19663);
nand U22179 (N_22179,N_21277,N_21246);
and U22180 (N_22180,N_19495,N_21824);
xor U22181 (N_22181,N_19185,N_21429);
and U22182 (N_22182,N_20990,N_20729);
nand U22183 (N_22183,N_19260,N_21385);
and U22184 (N_22184,N_20346,N_19878);
xnor U22185 (N_22185,N_19776,N_21098);
and U22186 (N_22186,N_19618,N_18853);
and U22187 (N_22187,N_20254,N_19971);
xor U22188 (N_22188,N_19548,N_19485);
nor U22189 (N_22189,N_19550,N_21627);
or U22190 (N_22190,N_21034,N_19586);
xor U22191 (N_22191,N_19539,N_21259);
nand U22192 (N_22192,N_21193,N_20844);
nor U22193 (N_22193,N_20893,N_19888);
xnor U22194 (N_22194,N_19650,N_20423);
or U22195 (N_22195,N_19120,N_21074);
nor U22196 (N_22196,N_19730,N_20132);
xor U22197 (N_22197,N_18974,N_21655);
nor U22198 (N_22198,N_21297,N_19468);
or U22199 (N_22199,N_19759,N_19905);
or U22200 (N_22200,N_19813,N_18894);
nor U22201 (N_22201,N_19500,N_21119);
nand U22202 (N_22202,N_19940,N_19230);
and U22203 (N_22203,N_19854,N_19193);
nor U22204 (N_22204,N_19453,N_21712);
and U22205 (N_22205,N_20367,N_19739);
xor U22206 (N_22206,N_21644,N_20057);
xor U22207 (N_22207,N_21132,N_19135);
nor U22208 (N_22208,N_21358,N_21482);
nor U22209 (N_22209,N_20697,N_20457);
or U22210 (N_22210,N_21634,N_20867);
nor U22211 (N_22211,N_20725,N_19841);
or U22212 (N_22212,N_19794,N_21016);
or U22213 (N_22213,N_21771,N_18813);
nor U22214 (N_22214,N_21802,N_20873);
nand U22215 (N_22215,N_21512,N_18898);
xor U22216 (N_22216,N_19028,N_19433);
nand U22217 (N_22217,N_19192,N_18917);
nand U22218 (N_22218,N_21618,N_20072);
or U22219 (N_22219,N_20345,N_20540);
or U22220 (N_22220,N_21757,N_21166);
or U22221 (N_22221,N_19502,N_20515);
nor U22222 (N_22222,N_18998,N_20550);
and U22223 (N_22223,N_18829,N_19471);
nor U22224 (N_22224,N_20230,N_20333);
and U22225 (N_22225,N_20843,N_19426);
or U22226 (N_22226,N_19022,N_20472);
or U22227 (N_22227,N_19840,N_19746);
or U22228 (N_22228,N_18903,N_21165);
nor U22229 (N_22229,N_20777,N_20251);
nor U22230 (N_22230,N_21534,N_19319);
and U22231 (N_22231,N_21740,N_19757);
nand U22232 (N_22232,N_21439,N_19672);
xnor U22233 (N_22233,N_21171,N_19374);
nand U22234 (N_22234,N_19302,N_20710);
and U22235 (N_22235,N_21050,N_20892);
or U22236 (N_22236,N_20252,N_19195);
nand U22237 (N_22237,N_20850,N_21525);
or U22238 (N_22238,N_19425,N_19729);
xnor U22239 (N_22239,N_20855,N_19077);
nand U22240 (N_22240,N_20895,N_19749);
or U22241 (N_22241,N_19636,N_19569);
and U22242 (N_22242,N_18844,N_20705);
or U22243 (N_22243,N_21502,N_18830);
nor U22244 (N_22244,N_19436,N_21873);
xnor U22245 (N_22245,N_19842,N_18991);
nand U22246 (N_22246,N_20314,N_21337);
or U22247 (N_22247,N_20827,N_19343);
xor U22248 (N_22248,N_21279,N_21100);
or U22249 (N_22249,N_21457,N_19538);
nor U22250 (N_22250,N_21307,N_20446);
and U22251 (N_22251,N_20438,N_20397);
or U22252 (N_22252,N_19412,N_20038);
and U22253 (N_22253,N_21505,N_20861);
nor U22254 (N_22254,N_21579,N_18887);
xnor U22255 (N_22255,N_19080,N_20851);
nand U22256 (N_22256,N_19667,N_19365);
or U22257 (N_22257,N_20749,N_19522);
nand U22258 (N_22258,N_19543,N_19384);
or U22259 (N_22259,N_20212,N_20020);
xor U22260 (N_22260,N_19900,N_20773);
nor U22261 (N_22261,N_19023,N_21105);
and U22262 (N_22262,N_18807,N_19418);
and U22263 (N_22263,N_20370,N_20018);
nor U22264 (N_22264,N_19544,N_20470);
xor U22265 (N_22265,N_19138,N_19624);
xor U22266 (N_22266,N_21826,N_19383);
or U22267 (N_22267,N_20271,N_21481);
or U22268 (N_22268,N_20473,N_18946);
nor U22269 (N_22269,N_19473,N_21103);
and U22270 (N_22270,N_21501,N_19810);
or U22271 (N_22271,N_21699,N_18859);
or U22272 (N_22272,N_20159,N_19199);
nor U22273 (N_22273,N_18755,N_20033);
or U22274 (N_22274,N_19174,N_20651);
and U22275 (N_22275,N_21206,N_21030);
xor U22276 (N_22276,N_18833,N_21322);
and U22277 (N_22277,N_19718,N_19145);
xor U22278 (N_22278,N_19926,N_21397);
and U22279 (N_22279,N_19056,N_19000);
nand U22280 (N_22280,N_19879,N_20006);
nand U22281 (N_22281,N_19666,N_20619);
and U22282 (N_22282,N_19257,N_21046);
nand U22283 (N_22283,N_19134,N_20305);
nor U22284 (N_22284,N_20846,N_20450);
nand U22285 (N_22285,N_19464,N_20664);
nor U22286 (N_22286,N_19266,N_20335);
or U22287 (N_22287,N_19882,N_21646);
xnor U22288 (N_22288,N_20935,N_21145);
and U22289 (N_22289,N_19397,N_21051);
nor U22290 (N_22290,N_21044,N_19001);
nand U22291 (N_22291,N_21529,N_19561);
and U22292 (N_22292,N_21747,N_20366);
or U22293 (N_22293,N_20865,N_19075);
nor U22294 (N_22294,N_19366,N_21099);
nor U22295 (N_22295,N_20939,N_20069);
nand U22296 (N_22296,N_20142,N_18979);
nor U22297 (N_22297,N_18896,N_18936);
xor U22298 (N_22298,N_19962,N_20783);
nand U22299 (N_22299,N_19269,N_19239);
or U22300 (N_22300,N_21780,N_21564);
nor U22301 (N_22301,N_21197,N_21556);
xnor U22302 (N_22302,N_18919,N_19444);
or U22303 (N_22303,N_20523,N_19231);
xor U22304 (N_22304,N_21795,N_21306);
or U22305 (N_22305,N_19219,N_21217);
nand U22306 (N_22306,N_19588,N_19311);
or U22307 (N_22307,N_20832,N_21553);
and U22308 (N_22308,N_20285,N_21513);
nor U22309 (N_22309,N_20350,N_20866);
nor U22310 (N_22310,N_18905,N_18850);
xor U22311 (N_22311,N_19858,N_20759);
nor U22312 (N_22312,N_20459,N_19689);
xnor U22313 (N_22313,N_18994,N_19564);
or U22314 (N_22314,N_21386,N_21854);
nor U22315 (N_22315,N_20692,N_20965);
and U22316 (N_22316,N_19039,N_21693);
nand U22317 (N_22317,N_20429,N_19415);
and U22318 (N_22318,N_20812,N_19407);
or U22319 (N_22319,N_19562,N_21292);
nor U22320 (N_22320,N_20740,N_21829);
nor U22321 (N_22321,N_21022,N_21257);
xor U22322 (N_22322,N_19535,N_21555);
nand U22323 (N_22323,N_21592,N_19118);
nand U22324 (N_22324,N_21366,N_19336);
or U22325 (N_22325,N_20197,N_21111);
or U22326 (N_22326,N_20300,N_19692);
nand U22327 (N_22327,N_18914,N_20707);
xor U22328 (N_22328,N_20073,N_21383);
and U22329 (N_22329,N_21261,N_20716);
nand U22330 (N_22330,N_19612,N_20198);
nor U22331 (N_22331,N_19074,N_19837);
nand U22332 (N_22332,N_20621,N_20878);
and U22333 (N_22333,N_19941,N_20848);
nor U22334 (N_22334,N_20562,N_18816);
or U22335 (N_22335,N_18798,N_20204);
nor U22336 (N_22336,N_20263,N_19435);
nor U22337 (N_22337,N_21493,N_20109);
or U22338 (N_22338,N_19046,N_19641);
nor U22339 (N_22339,N_21767,N_19631);
or U22340 (N_22340,N_18760,N_19665);
or U22341 (N_22341,N_21701,N_19701);
nor U22342 (N_22342,N_19492,N_21694);
nand U22343 (N_22343,N_20426,N_21188);
or U22344 (N_22344,N_18770,N_21207);
nand U22345 (N_22345,N_21458,N_20684);
xnor U22346 (N_22346,N_20169,N_20210);
and U22347 (N_22347,N_19113,N_20623);
and U22348 (N_22348,N_20014,N_19952);
nor U22349 (N_22349,N_20269,N_20853);
nand U22350 (N_22350,N_19358,N_20108);
xor U22351 (N_22351,N_20701,N_19357);
or U22352 (N_22352,N_19806,N_19800);
nor U22353 (N_22353,N_19049,N_21542);
and U22354 (N_22354,N_19177,N_20775);
nand U22355 (N_22355,N_20505,N_19674);
xnor U22356 (N_22356,N_19575,N_20195);
nand U22357 (N_22357,N_20223,N_20102);
or U22358 (N_22358,N_19737,N_19921);
or U22359 (N_22359,N_20171,N_20100);
xnor U22360 (N_22360,N_20309,N_20941);
xnor U22361 (N_22361,N_20821,N_20751);
nor U22362 (N_22362,N_21250,N_21067);
xnor U22363 (N_22363,N_20395,N_20712);
and U22364 (N_22364,N_18885,N_21652);
or U22365 (N_22365,N_19205,N_19181);
and U22366 (N_22366,N_20901,N_21375);
and U22367 (N_22367,N_18806,N_20516);
xor U22368 (N_22368,N_19823,N_19608);
and U22369 (N_22369,N_18930,N_19030);
xnor U22370 (N_22370,N_18956,N_21150);
nand U22371 (N_22371,N_21092,N_20597);
nor U22372 (N_22372,N_20170,N_20557);
nand U22373 (N_22373,N_19537,N_21313);
nand U22374 (N_22374,N_19703,N_21114);
xnor U22375 (N_22375,N_21235,N_21643);
xnor U22376 (N_22376,N_19153,N_21731);
nand U22377 (N_22377,N_20968,N_21742);
or U22378 (N_22378,N_20160,N_19402);
nor U22379 (N_22379,N_20961,N_20068);
xnor U22380 (N_22380,N_21848,N_21444);
xnor U22381 (N_22381,N_19606,N_18772);
nor U22382 (N_22382,N_20058,N_20218);
nand U22383 (N_22383,N_19738,N_21202);
or U22384 (N_22384,N_20719,N_21049);
nor U22385 (N_22385,N_20224,N_20430);
and U22386 (N_22386,N_20375,N_21174);
and U22387 (N_22387,N_20084,N_21670);
nand U22388 (N_22388,N_21093,N_18971);
or U22389 (N_22389,N_19934,N_21756);
xor U22390 (N_22390,N_19241,N_21538);
xnor U22391 (N_22391,N_20257,N_21139);
nand U22392 (N_22392,N_19147,N_19755);
nand U22393 (N_22393,N_20386,N_20922);
nand U22394 (N_22394,N_21507,N_19459);
xor U22395 (N_22395,N_21299,N_21748);
nand U22396 (N_22396,N_20139,N_21118);
xor U22397 (N_22397,N_18981,N_21342);
and U22398 (N_22398,N_20268,N_21777);
nand U22399 (N_22399,N_21511,N_20876);
nand U22400 (N_22400,N_19598,N_19043);
xor U22401 (N_22401,N_20798,N_20966);
nor U22402 (N_22402,N_20462,N_19133);
nor U22403 (N_22403,N_21372,N_20206);
nor U22404 (N_22404,N_18756,N_19287);
and U22405 (N_22405,N_21052,N_21781);
xnor U22406 (N_22406,N_21242,N_19811);
xnor U22407 (N_22407,N_19291,N_19299);
nor U22408 (N_22408,N_18848,N_20641);
xor U22409 (N_22409,N_20530,N_18857);
xnor U22410 (N_22410,N_21038,N_21228);
nand U22411 (N_22411,N_21384,N_21158);
xnor U22412 (N_22412,N_20779,N_20624);
nor U22413 (N_22413,N_19904,N_19236);
nand U22414 (N_22414,N_21019,N_20724);
nor U22415 (N_22415,N_19924,N_19604);
xnor U22416 (N_22416,N_20097,N_20787);
nor U22417 (N_22417,N_20476,N_20001);
xor U22418 (N_22418,N_19818,N_20467);
nand U22419 (N_22419,N_18845,N_19796);
nand U22420 (N_22420,N_18924,N_20117);
or U22421 (N_22421,N_18776,N_21715);
nor U22422 (N_22422,N_20978,N_20608);
nand U22423 (N_22423,N_21412,N_21483);
xor U22424 (N_22424,N_21466,N_19897);
nor U22425 (N_22425,N_20622,N_21488);
or U22426 (N_22426,N_21519,N_20755);
xor U22427 (N_22427,N_19364,N_19363);
nor U22428 (N_22428,N_21163,N_19142);
or U22429 (N_22429,N_19886,N_19990);
and U22430 (N_22430,N_19724,N_19072);
xor U22431 (N_22431,N_20653,N_21032);
nor U22432 (N_22432,N_20970,N_21187);
or U22433 (N_22433,N_20596,N_19640);
nor U22434 (N_22434,N_21102,N_20794);
and U22435 (N_22435,N_19062,N_20477);
nand U22436 (N_22436,N_21134,N_19741);
and U22437 (N_22437,N_20607,N_20276);
nor U22438 (N_22438,N_19127,N_19752);
nand U22439 (N_22439,N_20211,N_20037);
nand U22440 (N_22440,N_21161,N_20095);
or U22441 (N_22441,N_21130,N_20984);
nand U22442 (N_22442,N_21006,N_20957);
and U22443 (N_22443,N_19457,N_20924);
and U22444 (N_22444,N_18895,N_19262);
nand U22445 (N_22445,N_21296,N_20422);
xor U22446 (N_22446,N_21863,N_20960);
and U22447 (N_22447,N_21023,N_19413);
nor U22448 (N_22448,N_21234,N_20260);
nand U22449 (N_22449,N_19894,N_21590);
nor U22450 (N_22450,N_20019,N_21008);
nor U22451 (N_22451,N_20590,N_19988);
or U22452 (N_22452,N_19229,N_18975);
xor U22453 (N_22453,N_20668,N_18858);
or U22454 (N_22454,N_20904,N_19323);
nand U22455 (N_22455,N_20685,N_21024);
or U22456 (N_22456,N_21516,N_19394);
and U22457 (N_22457,N_19530,N_20187);
and U22458 (N_22458,N_20454,N_19060);
nand U22459 (N_22459,N_21214,N_18797);
nor U22460 (N_22460,N_20178,N_20576);
nand U22461 (N_22461,N_20278,N_18918);
or U22462 (N_22462,N_21790,N_21474);
xor U22463 (N_22463,N_21647,N_21520);
nand U22464 (N_22464,N_18777,N_19853);
and U22465 (N_22465,N_21822,N_19695);
nor U22466 (N_22466,N_20173,N_20028);
nand U22467 (N_22467,N_18758,N_19275);
nor U22468 (N_22468,N_19885,N_21685);
nand U22469 (N_22469,N_19600,N_20588);
or U22470 (N_22470,N_20181,N_20980);
and U22471 (N_22471,N_20385,N_20363);
nor U22472 (N_22472,N_18817,N_20918);
nand U22473 (N_22473,N_21179,N_20790);
or U22474 (N_22474,N_19508,N_19344);
or U22475 (N_22475,N_19558,N_21237);
or U22476 (N_22476,N_19356,N_20083);
and U22477 (N_22477,N_18827,N_21801);
nor U22478 (N_22478,N_19909,N_20795);
nor U22479 (N_22479,N_19293,N_21333);
or U22480 (N_22480,N_19770,N_19983);
nor U22481 (N_22481,N_19836,N_19371);
or U22482 (N_22482,N_19215,N_19844);
nor U22483 (N_22483,N_20382,N_19565);
xor U22484 (N_22484,N_20307,N_20567);
or U22485 (N_22485,N_21613,N_19314);
or U22486 (N_22486,N_20408,N_21320);
nand U22487 (N_22487,N_21460,N_19948);
nand U22488 (N_22488,N_21120,N_20129);
nand U22489 (N_22489,N_20869,N_19540);
and U22490 (N_22490,N_20964,N_19577);
nor U22491 (N_22491,N_18814,N_19908);
or U22492 (N_22492,N_21614,N_20760);
or U22493 (N_22493,N_20944,N_19381);
xnor U22494 (N_22494,N_18893,N_19942);
nand U22495 (N_22495,N_21451,N_21716);
or U22496 (N_22496,N_21245,N_20756);
nor U22497 (N_22497,N_20056,N_21807);
or U22498 (N_22498,N_20642,N_20545);
or U22499 (N_22499,N_21576,N_18890);
nand U22500 (N_22500,N_18869,N_19188);
nor U22501 (N_22501,N_21595,N_19728);
nand U22502 (N_22502,N_21047,N_20203);
nor U22503 (N_22503,N_18826,N_19292);
xnor U22504 (N_22504,N_18788,N_20671);
nand U22505 (N_22505,N_20162,N_21096);
and U22506 (N_22506,N_21831,N_19602);
xnor U22507 (N_22507,N_19377,N_19515);
xnor U22508 (N_22508,N_20079,N_20952);
xor U22509 (N_22509,N_19680,N_20772);
nor U22510 (N_22510,N_21464,N_21121);
nor U22511 (N_22511,N_19802,N_19342);
xnor U22512 (N_22512,N_21144,N_20656);
nand U22513 (N_22513,N_20618,N_19974);
xnor U22514 (N_22514,N_20190,N_20655);
nor U22515 (N_22515,N_21359,N_21356);
and U22516 (N_22516,N_20063,N_19375);
or U22517 (N_22517,N_19303,N_19711);
nand U22518 (N_22518,N_20830,N_21612);
nand U22519 (N_22519,N_21726,N_19778);
xnor U22520 (N_22520,N_19301,N_18947);
and U22521 (N_22521,N_21452,N_21423);
nand U22522 (N_22522,N_21764,N_19527);
nor U22523 (N_22523,N_19439,N_21572);
xor U22524 (N_22524,N_21632,N_21229);
and U22525 (N_22525,N_20086,N_19726);
and U22526 (N_22526,N_20336,N_20288);
nor U22527 (N_22527,N_19808,N_21298);
or U22528 (N_22528,N_21328,N_19057);
nor U22529 (N_22529,N_20050,N_20796);
nand U22530 (N_22530,N_19180,N_21248);
xnor U22531 (N_22531,N_19306,N_21663);
nand U22532 (N_22532,N_19024,N_19654);
nor U22533 (N_22533,N_20648,N_19890);
nor U22534 (N_22534,N_20234,N_21396);
xor U22535 (N_22535,N_19555,N_20122);
nor U22536 (N_22536,N_19727,N_21463);
nand U22537 (N_22537,N_20131,N_20556);
and U22538 (N_22538,N_19162,N_19679);
and U22539 (N_22539,N_19207,N_20090);
nand U22540 (N_22540,N_21442,N_19475);
nand U22541 (N_22541,N_20788,N_19534);
nand U22542 (N_22542,N_20560,N_21459);
nor U22543 (N_22543,N_20010,N_20877);
and U22544 (N_22544,N_18809,N_20738);
nor U22545 (N_22545,N_18846,N_21360);
or U22546 (N_22546,N_18978,N_18907);
xor U22547 (N_22547,N_20258,N_20898);
nor U22548 (N_22548,N_21522,N_19228);
xnor U22549 (N_22549,N_20388,N_21836);
and U22550 (N_22550,N_20326,N_19675);
nor U22551 (N_22551,N_19085,N_20321);
nor U22552 (N_22552,N_19685,N_21636);
nand U22553 (N_22553,N_18838,N_21070);
or U22554 (N_22554,N_20575,N_20527);
or U22555 (N_22555,N_20574,N_21509);
and U22556 (N_22556,N_20155,N_21172);
nand U22557 (N_22557,N_21661,N_19296);
nor U22558 (N_22558,N_20082,N_21434);
or U22559 (N_22559,N_18868,N_18968);
nor U22560 (N_22560,N_21713,N_20026);
and U22561 (N_22561,N_19657,N_20717);
or U22562 (N_22562,N_20469,N_18854);
xor U22563 (N_22563,N_20815,N_21380);
or U22564 (N_22564,N_19201,N_20536);
xor U22565 (N_22565,N_20319,N_21544);
and U22566 (N_22566,N_19332,N_21053);
xor U22567 (N_22567,N_21773,N_21265);
xor U22568 (N_22568,N_21853,N_21596);
nand U22569 (N_22569,N_21369,N_20040);
nor U22570 (N_22570,N_19406,N_19949);
nor U22571 (N_22571,N_21506,N_19864);
and U22572 (N_22572,N_18899,N_21057);
or U22573 (N_22573,N_19449,N_20958);
nor U22574 (N_22574,N_19827,N_20085);
and U22575 (N_22575,N_18952,N_20514);
or U22576 (N_22576,N_19480,N_21617);
or U22577 (N_22577,N_20905,N_18781);
nor U22578 (N_22578,N_20912,N_19783);
nor U22579 (N_22579,N_19175,N_20120);
or U22580 (N_22580,N_19987,N_19324);
nor U22581 (N_22581,N_19008,N_20636);
or U22582 (N_22582,N_20780,N_19566);
xnor U22583 (N_22583,N_19171,N_20951);
or U22584 (N_22584,N_20448,N_21113);
nor U22585 (N_22585,N_19634,N_20325);
and U22586 (N_22586,N_20744,N_19985);
nor U22587 (N_22587,N_19979,N_20439);
or U22588 (N_22588,N_19136,N_21734);
nand U22589 (N_22589,N_20902,N_19087);
nor U22590 (N_22590,N_19474,N_21862);
xor U22591 (N_22591,N_21091,N_20267);
nand U22592 (N_22592,N_19227,N_19125);
or U22593 (N_22593,N_20802,N_19519);
xnor U22594 (N_22594,N_21448,N_20248);
nand U22595 (N_22595,N_19032,N_19609);
xnor U22596 (N_22596,N_19684,N_21310);
xor U22597 (N_22597,N_20193,N_19845);
or U22598 (N_22598,N_21548,N_19651);
or U22599 (N_22599,N_18773,N_20945);
or U22600 (N_22600,N_20266,N_21842);
and U22601 (N_22601,N_20311,N_18920);
or U22602 (N_22602,N_19116,N_19743);
and U22603 (N_22603,N_20199,N_20610);
nand U22604 (N_22604,N_19714,N_19033);
or U22605 (N_22605,N_20232,N_20694);
xor U22606 (N_22606,N_19664,N_20565);
nand U22607 (N_22607,N_21332,N_20067);
xnor U22608 (N_22608,N_19843,N_21209);
xnor U22609 (N_22609,N_19850,N_21319);
nor U22610 (N_22610,N_19623,N_20741);
or U22611 (N_22611,N_21414,N_21240);
or U22612 (N_22612,N_18953,N_20262);
or U22613 (N_22613,N_20883,N_18927);
xnor U22614 (N_22614,N_19312,N_19777);
nor U22615 (N_22615,N_19411,N_20963);
nand U22616 (N_22616,N_19202,N_19933);
or U22617 (N_22617,N_19387,N_20125);
or U22618 (N_22618,N_21035,N_20416);
nand U22619 (N_22619,N_19420,N_18761);
nor U22620 (N_22620,N_21262,N_21355);
and U22621 (N_22621,N_21725,N_21584);
nor U22622 (N_22622,N_20299,N_20702);
xor U22623 (N_22623,N_18831,N_21176);
nor U22624 (N_22624,N_20146,N_20541);
or U22625 (N_22625,N_20214,N_20691);
nand U22626 (N_22626,N_21147,N_19677);
nand U22627 (N_22627,N_19595,N_20679);
nand U22628 (N_22628,N_18852,N_21752);
nor U22629 (N_22629,N_19437,N_20164);
and U22630 (N_22630,N_19477,N_20334);
nor U22631 (N_22631,N_19880,N_21048);
xor U22632 (N_22632,N_20730,N_20566);
or U22633 (N_22633,N_21376,N_21005);
and U22634 (N_22634,N_19484,N_20105);
nand U22635 (N_22635,N_21838,N_19567);
or U22636 (N_22636,N_20769,N_18799);
nor U22637 (N_22637,N_20956,N_19702);
nor U22638 (N_22638,N_20427,N_21128);
xnor U22639 (N_22639,N_20923,N_20568);
xor U22640 (N_22640,N_19754,N_19493);
or U22641 (N_22641,N_19912,N_21669);
and U22642 (N_22642,N_20280,N_19034);
xor U22643 (N_22643,N_20351,N_19339);
and U22644 (N_22644,N_20579,N_19831);
xor U22645 (N_22645,N_20167,N_19799);
nand U22646 (N_22646,N_19954,N_20513);
nand U22647 (N_22647,N_21681,N_19378);
or U22648 (N_22648,N_18932,N_21789);
or U22649 (N_22649,N_20485,N_20753);
xnor U22650 (N_22650,N_19715,N_21850);
or U22651 (N_22651,N_21758,N_21723);
or U22652 (N_22652,N_21431,N_18941);
xor U22653 (N_22653,N_20785,N_19972);
nand U22654 (N_22654,N_19893,N_20906);
and U22655 (N_22655,N_18796,N_19327);
or U22656 (N_22656,N_20287,N_21056);
or U22657 (N_22657,N_19690,N_21728);
nor U22658 (N_22658,N_18782,N_19814);
and U22659 (N_22659,N_20369,N_21689);
xor U22660 (N_22660,N_20594,N_21363);
and U22661 (N_22661,N_20194,N_19401);
and U22662 (N_22662,N_19863,N_21865);
and U22663 (N_22663,N_19733,N_20981);
or U22664 (N_22664,N_21243,N_19395);
nand U22665 (N_22665,N_19829,N_19385);
nor U22666 (N_22666,N_21177,N_19736);
and U22667 (N_22667,N_20383,N_21475);
nor U22668 (N_22668,N_21812,N_19273);
xor U22669 (N_22669,N_20110,N_19167);
xnor U22670 (N_22670,N_21404,N_20360);
or U22671 (N_22671,N_21856,N_20811);
or U22672 (N_22672,N_20631,N_19373);
xor U22673 (N_22673,N_21167,N_20104);
nand U22674 (N_22674,N_20064,N_21494);
and U22675 (N_22675,N_18871,N_21839);
or U22676 (N_22676,N_20184,N_20907);
nor U22677 (N_22677,N_21588,N_19212);
and U22678 (N_22678,N_19709,N_19197);
nor U22679 (N_22679,N_19015,N_21339);
xor U22680 (N_22680,N_20340,N_20708);
nor U22681 (N_22681,N_21266,N_19004);
nand U22682 (N_22682,N_19172,N_21213);
or U22683 (N_22683,N_20434,N_19763);
nor U22684 (N_22684,N_21575,N_21254);
xnor U22685 (N_22685,N_20468,N_21750);
and U22686 (N_22686,N_19498,N_19889);
nor U22687 (N_22687,N_19190,N_18958);
nor U22688 (N_22688,N_19006,N_21287);
nor U22689 (N_22689,N_21808,N_20081);
nand U22690 (N_22690,N_19182,N_19747);
xnor U22691 (N_22691,N_20049,N_20606);
nand U22692 (N_22692,N_19315,N_21817);
nand U22693 (N_22693,N_19213,N_21178);
xor U22694 (N_22694,N_19820,N_20406);
nand U22695 (N_22695,N_21275,N_20112);
nor U22696 (N_22696,N_18933,N_19981);
xor U22697 (N_22697,N_19379,N_19194);
xnor U22698 (N_22698,N_21650,N_20754);
nor U22699 (N_22699,N_20720,N_21666);
nor U22700 (N_22700,N_20176,N_19788);
and U22701 (N_22701,N_20706,N_21751);
nand U22702 (N_22702,N_20938,N_20698);
nor U22703 (N_22703,N_19980,N_20356);
xnor U22704 (N_22704,N_20133,N_21504);
xnor U22705 (N_22705,N_20235,N_18910);
nand U22706 (N_22706,N_20954,N_19044);
or U22707 (N_22707,N_20676,N_19649);
xor U22708 (N_22708,N_19335,N_20825);
nor U22709 (N_22709,N_20914,N_18759);
and U22710 (N_22710,N_19163,N_20637);
xnor U22711 (N_22711,N_21269,N_21487);
or U22712 (N_22712,N_19920,N_19214);
and U22713 (N_22713,N_18995,N_18996);
nand U22714 (N_22714,N_19884,N_19895);
nand U22715 (N_22715,N_20480,N_21274);
or U22716 (N_22716,N_21041,N_19688);
nand U22717 (N_22717,N_20526,N_21772);
and U22718 (N_22718,N_21249,N_21252);
xnor U22719 (N_22719,N_21558,N_20244);
or U22720 (N_22720,N_19626,N_21717);
nor U22721 (N_22721,N_21352,N_21344);
xor U22722 (N_22722,N_18872,N_21295);
and U22723 (N_22723,N_19146,N_20265);
or U22724 (N_22724,N_20711,N_19067);
xor U22725 (N_22725,N_19042,N_21373);
xor U22726 (N_22726,N_21338,N_19501);
and U22727 (N_22727,N_21799,N_20967);
nand U22728 (N_22728,N_21215,N_18922);
and U22729 (N_22729,N_18915,N_21138);
and U22730 (N_22730,N_20256,N_20699);
nor U22731 (N_22731,N_21708,N_20654);
and U22732 (N_22732,N_21518,N_21409);
nand U22733 (N_22733,N_20275,N_20767);
nor U22734 (N_22734,N_21424,N_20872);
xnor U22735 (N_22735,N_19531,N_19824);
or U22736 (N_22736,N_20207,N_19447);
xor U22737 (N_22737,N_21453,N_20343);
or U22738 (N_22738,N_20329,N_21353);
nor U22739 (N_22739,N_20380,N_21658);
or U22740 (N_22740,N_19740,N_21495);
and U22741 (N_22741,N_20657,N_21626);
xnor U22742 (N_22742,N_20838,N_21194);
nand U22743 (N_22743,N_19572,N_20017);
and U22744 (N_22744,N_20983,N_20025);
and U22745 (N_22745,N_19860,N_21591);
and U22746 (N_22746,N_19389,N_19668);
xor U22747 (N_22747,N_21746,N_21341);
xor U22748 (N_22748,N_21164,N_20331);
and U22749 (N_22749,N_21827,N_20704);
nor U22750 (N_22750,N_20153,N_20660);
xnor U22751 (N_22751,N_20494,N_20771);
xnor U22752 (N_22752,N_19935,N_20458);
or U22753 (N_22753,N_21755,N_19108);
nand U22754 (N_22754,N_18948,N_19160);
and U22755 (N_22755,N_20778,N_19245);
and U22756 (N_22756,N_19036,N_20240);
or U22757 (N_22757,N_20291,N_19819);
and U22758 (N_22758,N_20683,N_19012);
and U22759 (N_22759,N_21438,N_19169);
nand U22760 (N_22760,N_19614,N_20899);
xnor U22761 (N_22761,N_20700,N_18843);
nand U22762 (N_22762,N_19896,N_21075);
nand U22763 (N_22763,N_20039,N_19969);
nor U22764 (N_22764,N_20879,N_19570);
nor U22765 (N_22765,N_21739,N_20934);
nor U22766 (N_22766,N_19846,N_21162);
xor U22767 (N_22767,N_19340,N_20465);
or U22768 (N_22768,N_19059,N_19647);
nand U22769 (N_22769,N_19376,N_21009);
nand U22770 (N_22770,N_20242,N_19731);
nand U22771 (N_22771,N_19278,N_20419);
nand U22772 (N_22772,N_21687,N_20561);
nand U22773 (N_22773,N_20552,N_18779);
nand U22774 (N_22774,N_19927,N_20353);
or U22775 (N_22775,N_21156,N_20312);
and U22776 (N_22776,N_20628,N_19638);
xor U22777 (N_22777,N_21189,N_20009);
xor U22778 (N_22778,N_19722,N_21394);
or U22779 (N_22779,N_20042,N_19613);
xnor U22780 (N_22780,N_20974,N_19721);
and U22781 (N_22781,N_19951,N_20897);
nand U22782 (N_22782,N_20466,N_20612);
or U22783 (N_22783,N_20191,N_20789);
nor U22784 (N_22784,N_20044,N_19244);
xor U22785 (N_22785,N_21770,N_21580);
nand U22786 (N_22786,N_21449,N_21026);
xor U22787 (N_22787,N_20302,N_20030);
xor U22788 (N_22788,N_20820,N_19622);
xor U22789 (N_22789,N_21683,N_19322);
or U22790 (N_22790,N_19047,N_20609);
and U22791 (N_22791,N_21220,N_20487);
and U22792 (N_22792,N_19388,N_20361);
xor U22793 (N_22793,N_19422,N_20396);
xnor U22794 (N_22794,N_20739,N_18950);
nor U22795 (N_22795,N_18954,N_20999);
or U22796 (N_22796,N_21168,N_19497);
and U22797 (N_22797,N_21869,N_20229);
xnor U22798 (N_22798,N_20294,N_21133);
nand U22799 (N_22799,N_21286,N_21859);
nand U22800 (N_22800,N_19704,N_20124);
nor U22801 (N_22801,N_21407,N_19968);
nand U22802 (N_22802,N_21738,N_21866);
nor U22803 (N_22803,N_21413,N_21805);
or U22804 (N_22804,N_19321,N_21447);
xnor U22805 (N_22805,N_19937,N_20219);
nor U22806 (N_22806,N_20273,N_21774);
nor U22807 (N_22807,N_18976,N_18800);
nor U22808 (N_22808,N_20411,N_21762);
xnor U22809 (N_22809,N_19938,N_19683);
nand U22810 (N_22810,N_21561,N_19786);
xnor U22811 (N_22811,N_20119,N_20503);
and U22812 (N_22812,N_19887,N_20126);
nand U22813 (N_22813,N_21628,N_21749);
nor U22814 (N_22814,N_20047,N_21020);
nand U22815 (N_22815,N_19998,N_19964);
and U22816 (N_22816,N_20298,N_19052);
nor U22817 (N_22817,N_20228,N_21418);
xnor U22818 (N_22818,N_19489,N_20709);
nor U22819 (N_22819,N_20070,N_19463);
nand U22820 (N_22820,N_20831,N_20605);
or U22821 (N_22821,N_19351,N_21382);
xnor U22822 (N_22822,N_20135,N_21462);
and U22823 (N_22823,N_19977,N_19932);
nand U22824 (N_22824,N_18937,N_21000);
or U22825 (N_22825,N_19790,N_20183);
and U22826 (N_22826,N_18940,N_18861);
nand U22827 (N_22827,N_19235,N_20441);
or U22828 (N_22828,N_21785,N_20992);
and U22829 (N_22829,N_19643,N_19775);
nand U22830 (N_22830,N_19991,N_21117);
xor U22831 (N_22831,N_21676,N_20186);
and U22832 (N_22832,N_20486,N_21605);
nor U22833 (N_22833,N_20613,N_19512);
or U22834 (N_22834,N_21031,N_18962);
or U22835 (N_22835,N_21270,N_20209);
nor U22836 (N_22836,N_19693,N_20860);
nor U22837 (N_22837,N_20890,N_20746);
and U22838 (N_22838,N_20837,N_20633);
nand U22839 (N_22839,N_19859,N_21845);
and U22840 (N_22840,N_19173,N_19901);
xor U22841 (N_22841,N_20626,N_19222);
xor U22842 (N_22842,N_20424,N_20348);
and U22843 (N_22843,N_21137,N_19915);
nor U22844 (N_22844,N_21465,N_21219);
or U22845 (N_22845,N_20587,N_20804);
nand U22846 (N_22846,N_20500,N_18912);
xor U22847 (N_22847,N_21454,N_20840);
xor U22848 (N_22848,N_19902,N_20506);
nor U22849 (N_22849,N_20862,N_20520);
nand U22850 (N_22850,N_21479,N_19642);
nor U22851 (N_22851,N_18767,N_20400);
or U22852 (N_22852,N_21315,N_18780);
or U22853 (N_22853,N_19589,N_20182);
or U22854 (N_22854,N_18791,N_20021);
and U22855 (N_22855,N_21381,N_20714);
or U22856 (N_22856,N_19673,N_19682);
or U22857 (N_22857,N_21112,N_21765);
and U22858 (N_22858,N_20675,N_21672);
nand U22859 (N_22859,N_18923,N_18828);
xor U22860 (N_22860,N_19137,N_21533);
nand U22861 (N_22861,N_20762,N_20185);
xnor U22862 (N_22862,N_19791,N_19254);
nor U22863 (N_22863,N_18945,N_20639);
and U22864 (N_22864,N_19454,N_21860);
nor U22865 (N_22865,N_21562,N_20013);
nor U22866 (N_22866,N_21702,N_20374);
xor U22867 (N_22867,N_20282,N_20672);
nor U22868 (N_22868,N_20149,N_19552);
and U22869 (N_22869,N_19178,N_19068);
nor U22870 (N_22870,N_18775,N_20824);
xor U22871 (N_22871,N_21084,N_19341);
and U22872 (N_22872,N_20784,N_19835);
and U22873 (N_22873,N_19855,N_20225);
xnor U22874 (N_22874,N_21619,N_20365);
nor U22875 (N_22875,N_21058,N_21849);
nand U22876 (N_22876,N_19591,N_21844);
nor U22877 (N_22877,N_21391,N_19956);
xor U22878 (N_22878,N_20296,N_21753);
xor U22879 (N_22879,N_20078,N_19630);
or U22880 (N_22880,N_21272,N_20630);
xor U22881 (N_22881,N_18965,N_21280);
or U22882 (N_22882,N_20492,N_21061);
nor U22883 (N_22883,N_18862,N_21820);
and U22884 (N_22884,N_19161,N_21581);
or U22885 (N_22885,N_21186,N_21828);
nand U22886 (N_22886,N_18879,N_20460);
nand U22887 (N_22887,N_21314,N_21794);
nor U22888 (N_22888,N_19264,N_21857);
nor U22889 (N_22889,N_21456,N_20163);
nor U22890 (N_22890,N_21523,N_19928);
nand U22891 (N_22891,N_21154,N_20643);
nand U22892 (N_22892,N_21800,N_19669);
nor U22893 (N_22893,N_21582,N_21797);
and U22894 (N_22894,N_21744,N_20669);
nand U22895 (N_22895,N_20856,N_19105);
nand U22896 (N_22896,N_19243,N_20659);
or U22897 (N_22897,N_18992,N_21657);
nor U22898 (N_22898,N_20752,N_19694);
nor U22899 (N_22899,N_20387,N_19109);
nor U22900 (N_22900,N_20681,N_19005);
and U22901 (N_22901,N_20537,N_19246);
or U22902 (N_22902,N_21175,N_20920);
or U22903 (N_22903,N_21735,N_20911);
nor U22904 (N_22904,N_21804,N_19233);
nor U22905 (N_22905,N_20539,N_21843);
xor U22906 (N_22906,N_18900,N_18832);
nor U22907 (N_22907,N_19532,N_19476);
nor U22908 (N_22908,N_19825,N_21625);
or U22909 (N_22909,N_19633,N_20509);
and U22910 (N_22910,N_21010,N_20936);
or U22911 (N_22911,N_20863,N_19141);
nand U22912 (N_22912,N_19431,N_21085);
nand U22913 (N_22913,N_20342,N_21232);
nand U22914 (N_22914,N_18750,N_20442);
and U22915 (N_22915,N_21432,N_18908);
xor U22916 (N_22916,N_21696,N_20297);
xnor U22917 (N_22917,N_19482,N_20661);
or U22918 (N_22918,N_19670,N_19801);
or U22919 (N_22919,N_21768,N_20404);
or U22920 (N_22920,N_19617,N_19088);
or U22921 (N_22921,N_21478,N_18926);
xor U22922 (N_22922,N_19874,N_20564);
and U22923 (N_22923,N_20658,N_21399);
or U22924 (N_22924,N_19518,N_20238);
and U22925 (N_22925,N_21732,N_21782);
nor U22926 (N_22926,N_20522,N_18751);
and U22927 (N_22927,N_18964,N_19955);
nor U22928 (N_22928,N_21349,N_19392);
xor U22929 (N_22929,N_21640,N_19288);
and U22930 (N_22930,N_21065,N_21251);
nand U22931 (N_22931,N_20004,N_21039);
nor U22932 (N_22932,N_19206,N_19434);
xor U22933 (N_22933,N_20440,N_20734);
nor U22934 (N_22934,N_19826,N_20055);
nor U22935 (N_22935,N_18876,N_19223);
nand U22936 (N_22936,N_21325,N_20884);
and U22937 (N_22937,N_19644,N_20496);
nor U22938 (N_22938,N_21497,N_19150);
nand U22939 (N_22939,N_20532,N_19408);
nor U22940 (N_22940,N_19767,N_19803);
or U22941 (N_22941,N_20549,N_21437);
or U22942 (N_22942,N_19071,N_21271);
or U22943 (N_22943,N_19766,N_19976);
nand U22944 (N_22944,N_20859,N_20022);
or U22945 (N_22945,N_21722,N_20810);
and U22946 (N_22946,N_21665,N_19525);
or U22947 (N_22947,N_21651,N_19723);
nand U22948 (N_22948,N_19708,N_21469);
and U22949 (N_22949,N_19176,N_20368);
and U22950 (N_22950,N_18808,N_21072);
xor U22951 (N_22951,N_19996,N_19992);
nand U22952 (N_22952,N_20435,N_19054);
nand U22953 (N_22953,N_19076,N_19350);
xnor U22954 (N_22954,N_19249,N_20261);
nor U22955 (N_22955,N_20315,N_18774);
xnor U22956 (N_22956,N_18944,N_20925);
xor U22957 (N_22957,N_20313,N_20421);
and U22958 (N_22958,N_19805,N_21792);
xor U22959 (N_22959,N_19645,N_21324);
and U22960 (N_22960,N_20678,N_21028);
and U22961 (N_22961,N_21054,N_18783);
nor U22962 (N_22962,N_19917,N_21323);
and U22963 (N_22963,N_19098,N_21043);
nor U22964 (N_22964,N_21761,N_19526);
nand U22965 (N_22965,N_18753,N_20768);
and U22966 (N_22966,N_20227,N_21692);
and U22967 (N_22967,N_21151,N_18794);
and U22968 (N_22968,N_18865,N_21745);
or U22969 (N_22969,N_21697,N_20003);
nor U22970 (N_22970,N_19916,N_21589);
xnor U22971 (N_22971,N_19020,N_20377);
nor U22972 (N_22972,N_19283,N_20581);
xor U22973 (N_22973,N_21648,N_19238);
or U22974 (N_22974,N_21527,N_21086);
xnor U22975 (N_22975,N_20484,N_20060);
or U22976 (N_22976,N_19123,N_21551);
nand U22977 (N_22977,N_20264,N_19930);
or U22978 (N_22978,N_20147,N_19774);
nor U22979 (N_22979,N_19621,N_20625);
or U22980 (N_22980,N_20455,N_19126);
or U22981 (N_22981,N_18802,N_20781);
nand U22982 (N_22982,N_19183,N_19773);
and U22983 (N_22983,N_18901,N_21076);
and U22984 (N_22984,N_19661,N_21285);
nand U22985 (N_22985,N_19095,N_21191);
and U22986 (N_22986,N_21157,N_21059);
nand U22987 (N_22987,N_21489,N_21025);
nor U22988 (N_22988,N_21231,N_19509);
nor U22989 (N_22989,N_19560,N_20947);
xor U22990 (N_22990,N_20381,N_19870);
nand U22991 (N_22991,N_20975,N_21864);
and U22992 (N_22992,N_19289,N_18988);
xor U22993 (N_22993,N_19610,N_19360);
nor U22994 (N_22994,N_20554,N_21395);
nand U22995 (N_22995,N_21609,N_19662);
xor U22996 (N_22996,N_20875,N_21436);
nand U22997 (N_22997,N_20953,N_18805);
or U22998 (N_22998,N_20948,N_19050);
or U22999 (N_22999,N_19946,N_21388);
and U23000 (N_23000,N_20328,N_21256);
and U23001 (N_23001,N_20996,N_19576);
or U23002 (N_23002,N_20213,N_19130);
and U23003 (N_23003,N_21686,N_21531);
nor U23004 (N_23004,N_21846,N_21598);
or U23005 (N_23005,N_21335,N_20584);
nor U23006 (N_23006,N_20498,N_19817);
nand U23007 (N_23007,N_21063,N_20761);
and U23008 (N_23008,N_21624,N_20616);
and U23009 (N_23009,N_21350,N_19832);
xnor U23010 (N_23010,N_20582,N_19352);
nand U23011 (N_23011,N_19919,N_19698);
nor U23012 (N_23012,N_20138,N_19347);
or U23013 (N_23013,N_21719,N_20894);
nand U23014 (N_23014,N_21199,N_21668);
or U23015 (N_23015,N_19787,N_20882);
nor U23016 (N_23016,N_21680,N_20585);
or U23017 (N_23017,N_20979,N_19520);
nand U23018 (N_23018,N_19789,N_20226);
or U23019 (N_23019,N_19625,N_20379);
or U23020 (N_23020,N_20546,N_20962);
or U23021 (N_23021,N_19584,N_20880);
nor U23022 (N_23022,N_20005,N_21704);
or U23023 (N_23023,N_19862,N_21707);
and U23024 (N_23024,N_21573,N_20814);
or U23025 (N_23025,N_19469,N_18856);
nor U23026 (N_23026,N_19503,N_20940);
nor U23027 (N_23027,N_19159,N_19784);
nand U23028 (N_23028,N_20118,N_19993);
nand U23029 (N_23029,N_19822,N_20099);
nor U23030 (N_23030,N_21282,N_19999);
and U23031 (N_23031,N_20538,N_21357);
and U23032 (N_23032,N_20362,N_21607);
or U23033 (N_23033,N_20950,N_21779);
nor U23034 (N_23034,N_19593,N_19619);
nand U23035 (N_23035,N_21387,N_19568);
nor U23036 (N_23036,N_21198,N_21629);
and U23037 (N_23037,N_21587,N_21649);
or U23038 (N_23038,N_20813,N_21631);
or U23039 (N_23039,N_19009,N_21406);
xor U23040 (N_23040,N_20449,N_20106);
nor U23041 (N_23041,N_21021,N_21741);
and U23042 (N_23042,N_21370,N_19732);
nand U23043 (N_23043,N_20586,N_18866);
nor U23044 (N_23044,N_20917,N_18789);
nand U23045 (N_23045,N_19839,N_20640);
nor U23046 (N_23046,N_19807,N_19462);
xnor U23047 (N_23047,N_19073,N_20310);
or U23048 (N_23048,N_21823,N_19611);
or U23049 (N_23049,N_19797,N_19696);
xnor U23050 (N_23050,N_20555,N_20024);
xnor U23051 (N_23051,N_20393,N_19507);
or U23052 (N_23052,N_20680,N_21181);
and U23053 (N_23053,N_19923,N_18969);
xor U23054 (N_23054,N_19833,N_20903);
xor U23055 (N_23055,N_19152,N_21769);
nand U23056 (N_23056,N_18934,N_21011);
xnor U23057 (N_23057,N_18966,N_20543);
or U23058 (N_23058,N_18931,N_19279);
or U23059 (N_23059,N_19496,N_21586);
nand U23060 (N_23060,N_19184,N_20511);
nor U23061 (N_23061,N_20595,N_20341);
nand U23062 (N_23062,N_21155,N_21201);
xnor U23063 (N_23063,N_20096,N_19285);
and U23064 (N_23064,N_20401,N_19639);
xor U23065 (N_23065,N_21703,N_19659);
or U23066 (N_23066,N_20168,N_19760);
and U23067 (N_23067,N_19253,N_21210);
and U23068 (N_23068,N_19031,N_18891);
nor U23069 (N_23069,N_20797,N_19660);
nand U23070 (N_23070,N_21847,N_19656);
and U23071 (N_23071,N_20517,N_19297);
xor U23072 (N_23072,N_20475,N_21419);
nand U23073 (N_23073,N_21440,N_20274);
nor U23074 (N_23074,N_21400,N_20852);
nand U23075 (N_23075,N_19779,N_20318);
nor U23076 (N_23076,N_19597,N_21253);
and U23077 (N_23077,N_20330,N_19166);
and U23078 (N_23078,N_20358,N_19628);
nand U23079 (N_23079,N_20478,N_21311);
nand U23080 (N_23080,N_19225,N_19251);
nor U23081 (N_23081,N_20747,N_21107);
nand U23082 (N_23082,N_19248,N_20989);
nor U23083 (N_23083,N_20158,N_19467);
xor U23084 (N_23084,N_21656,N_21615);
and U23085 (N_23085,N_21226,N_19966);
xor U23086 (N_23086,N_20413,N_20114);
or U23087 (N_23087,N_20045,N_19430);
nor U23088 (N_23088,N_21608,N_21645);
nand U23089 (N_23089,N_19240,N_21874);
and U23090 (N_23090,N_20464,N_18959);
or U23091 (N_23091,N_20732,N_21571);
nor U23092 (N_23092,N_18864,N_20495);
xor U23093 (N_23093,N_21364,N_21002);
xor U23094 (N_23094,N_18847,N_19950);
xnor U23095 (N_23095,N_19268,N_21060);
nand U23096 (N_23096,N_21698,N_21610);
nor U23097 (N_23097,N_20816,N_19486);
xor U23098 (N_23098,N_21677,N_20765);
nand U23099 (N_23099,N_19093,N_19405);
nand U23100 (N_23100,N_20662,N_18943);
xor U23101 (N_23101,N_20611,N_21776);
nor U23102 (N_23102,N_21851,N_21815);
nand U23103 (N_23103,N_19906,N_18977);
nor U23104 (N_23104,N_19725,N_21336);
nand U23105 (N_23105,N_20644,N_21160);
nor U23106 (N_23106,N_19713,N_18840);
or U23107 (N_23107,N_21401,N_21365);
nand U23108 (N_23108,N_19361,N_19592);
nor U23109 (N_23109,N_19687,N_20208);
and U23110 (N_23110,N_21622,N_19367);
nor U23111 (N_23111,N_21268,N_21818);
nand U23112 (N_23112,N_20051,N_19256);
nor U23113 (N_23113,N_20463,N_19107);
nand U23114 (N_23114,N_19907,N_18993);
nand U23115 (N_23115,N_19632,N_19699);
xor U23116 (N_23116,N_20842,N_20075);
nor U23117 (N_23117,N_20123,N_21142);
nor U23118 (N_23118,N_21123,N_21559);
and U23119 (N_23119,N_19265,N_19947);
and U23120 (N_23120,N_20048,N_21227);
nand U23121 (N_23121,N_19960,N_21814);
nand U23122 (N_23122,N_21568,N_18906);
nand U23123 (N_23123,N_20115,N_19170);
and U23124 (N_23124,N_21152,N_20909);
and U23125 (N_23125,N_20041,N_20603);
xor U23126 (N_23126,N_21825,N_19007);
nand U23127 (N_23127,N_20140,N_20673);
xnor U23128 (N_23128,N_20670,N_20200);
and U23129 (N_23129,N_20489,N_19419);
and U23130 (N_23130,N_20293,N_19082);
and U23131 (N_23131,N_20969,N_19337);
nand U23132 (N_23132,N_20728,N_20093);
nor U23133 (N_23133,N_19989,N_20493);
nand U23134 (N_23134,N_18875,N_19599);
or U23135 (N_23135,N_21546,N_20076);
or U23136 (N_23136,N_21097,N_19691);
and U23137 (N_23137,N_19368,N_20161);
nand U23138 (N_23138,N_20378,N_19014);
nor U23139 (N_23139,N_19164,N_19943);
xor U23140 (N_23140,N_19620,N_19536);
and U23141 (N_23141,N_21018,N_19748);
and U23142 (N_23142,N_21405,N_19511);
xnor U23143 (N_23143,N_20995,N_21378);
nand U23144 (N_23144,N_19355,N_20283);
nand U23145 (N_23145,N_21334,N_21078);
nand U23146 (N_23146,N_20592,N_21714);
and U23147 (N_23147,N_21603,N_18984);
or U23148 (N_23148,N_19338,N_19716);
nand U23149 (N_23149,N_21001,N_20998);
nor U23150 (N_23150,N_21834,N_20295);
xor U23151 (N_23151,N_19294,N_18811);
and U23152 (N_23152,N_20231,N_19280);
or U23153 (N_23153,N_20286,N_20871);
and U23154 (N_23154,N_19011,N_20525);
and U23155 (N_23155,N_21783,N_21273);
nand U23156 (N_23156,N_21403,N_20570);
nand U23157 (N_23157,N_19745,N_19571);
nor U23158 (N_23158,N_19986,N_21267);
nor U23159 (N_23159,N_20143,N_19216);
nand U23160 (N_23160,N_21069,N_21835);
nand U23161 (N_23161,N_20246,N_21003);
or U23162 (N_23162,N_20927,N_19117);
nor U23163 (N_23163,N_20502,N_20929);
xnor U23164 (N_23164,N_20392,N_19258);
nand U23165 (N_23165,N_20239,N_20987);
xnor U23166 (N_23166,N_20693,N_21278);
xor U23167 (N_23167,N_21441,N_19154);
nor U23168 (N_23168,N_19158,N_18886);
nand U23169 (N_23169,N_21641,N_20916);
nand U23170 (N_23170,N_21230,N_19821);
or U23171 (N_23171,N_19452,N_19010);
or U23172 (N_23172,N_19510,N_18909);
or U23173 (N_23173,N_20023,N_20221);
nor U23174 (N_23174,N_19346,N_20529);
or U23175 (N_23175,N_19761,N_20583);
and U23176 (N_23176,N_21443,N_21149);
xor U23177 (N_23177,N_21042,N_19735);
or U23178 (N_23178,N_19635,N_19189);
xnor U23179 (N_23179,N_21583,N_21673);
or U23180 (N_23180,N_20364,N_21667);
and U23181 (N_23181,N_18882,N_20973);
and U23182 (N_23182,N_21635,N_21312);
nand U23183 (N_23183,N_19211,N_19861);
or U23184 (N_23184,N_19380,N_21289);
xor U23185 (N_23185,N_19040,N_20835);
nand U23186 (N_23186,N_19481,N_21684);
or U23187 (N_23187,N_20304,N_21724);
and U23188 (N_23188,N_19918,N_19144);
xnor U23189 (N_23189,N_20508,N_21775);
xnor U23190 (N_23190,N_21281,N_21064);
xor U23191 (N_23191,N_19533,N_19517);
nand U23192 (N_23192,N_20801,N_20497);
nand U23193 (N_23193,N_18935,N_21362);
nor U23194 (N_23194,N_20180,N_21017);
xnor U23195 (N_23195,N_20573,N_19002);
nor U23196 (N_23196,N_21073,N_21263);
xnor U23197 (N_23197,N_20490,N_21317);
or U23198 (N_23198,N_21303,N_19290);
or U23199 (N_23199,N_19122,N_20316);
nor U23200 (N_23200,N_21602,N_20062);
nor U23201 (N_23201,N_19554,N_20431);
nand U23202 (N_23202,N_20189,N_21294);
and U23203 (N_23203,N_20955,N_20390);
xnor U23204 (N_23204,N_21766,N_21014);
xor U23205 (N_23205,N_19224,N_19277);
nand U23206 (N_23206,N_19865,N_21729);
nor U23207 (N_23207,N_21810,N_21554);
nor U23208 (N_23208,N_20410,N_20881);
nor U23209 (N_23209,N_20799,N_19101);
and U23210 (N_23210,N_19470,N_19255);
xnor U23211 (N_23211,N_19541,N_20128);
and U23212 (N_23212,N_21066,N_20355);
nand U23213 (N_23213,N_19834,N_21543);
nor U23214 (N_23214,N_20172,N_18970);
or U23215 (N_23215,N_21080,N_20121);
and U23216 (N_23216,N_19931,N_20931);
nand U23217 (N_23217,N_18986,N_19849);
nand U23218 (N_23218,N_18870,N_19400);
and U23219 (N_23219,N_20986,N_21709);
or U23220 (N_23220,N_19487,N_21510);
nand U23221 (N_23221,N_21037,N_19460);
xor U23222 (N_23222,N_21705,N_20650);
or U23223 (N_23223,N_20864,N_21537);
and U23224 (N_23224,N_19658,N_20031);
nand U23225 (N_23225,N_20433,N_20888);
nor U23226 (N_23226,N_21496,N_19140);
xnor U23227 (N_23227,N_19856,N_20733);
and U23228 (N_23228,N_21221,N_19320);
nand U23229 (N_23229,N_21135,N_18987);
xor U23230 (N_23230,N_19081,N_21492);
and U23231 (N_23231,N_21354,N_19084);
xor U23232 (N_23232,N_21642,N_21604);
xnor U23233 (N_23233,N_18877,N_18997);
nand U23234 (N_23234,N_20461,N_21446);
or U23235 (N_23235,N_19442,N_20727);
nor U23236 (N_23236,N_19221,N_21077);
or U23237 (N_23237,N_21402,N_20695);
xnor U23238 (N_23238,N_19094,N_20409);
nor U23239 (N_23239,N_21491,N_20088);
or U23240 (N_23240,N_19210,N_21539);
or U23241 (N_23241,N_19961,N_21499);
nand U23242 (N_23242,N_20713,N_20066);
or U23243 (N_23243,N_19114,N_21872);
nand U23244 (N_23244,N_20301,N_19646);
nor U23245 (N_23245,N_20029,N_21660);
nor U23246 (N_23246,N_20077,N_18819);
nand U23247 (N_23247,N_21182,N_20667);
xor U23248 (N_23248,N_21616,N_20130);
nor U23249 (N_23249,N_19372,N_21428);
or U23250 (N_23250,N_19272,N_20145);
and U23251 (N_23251,N_20572,N_19753);
and U23252 (N_23252,N_18793,N_20742);
and U23253 (N_23253,N_21371,N_21674);
nor U23254 (N_23254,N_20758,N_20808);
and U23255 (N_23255,N_21012,N_21498);
and U23256 (N_23256,N_21819,N_19058);
nand U23257 (N_23257,N_19237,N_21433);
or U23258 (N_23258,N_20839,N_20703);
or U23259 (N_23259,N_19883,N_20036);
nand U23260 (N_23260,N_19242,N_19528);
or U23261 (N_23261,N_19061,N_20253);
xnor U23262 (N_23262,N_19466,N_19157);
and U23263 (N_23263,N_19959,N_20690);
nor U23264 (N_23264,N_19830,N_21549);
xnor U23265 (N_23265,N_21570,N_19143);
and U23266 (N_23266,N_21445,N_19110);
or U23267 (N_23267,N_21833,N_21577);
xnor U23268 (N_23268,N_20428,N_21416);
nor U23269 (N_23269,N_20157,N_21486);
and U23270 (N_23270,N_19607,N_20165);
and U23271 (N_23271,N_20144,N_20389);
and U23272 (N_23272,N_19204,N_20154);
or U23273 (N_23273,N_20134,N_20344);
and U23274 (N_23274,N_18784,N_20571);
or U23275 (N_23275,N_19066,N_19252);
and U23276 (N_23276,N_19128,N_19165);
nand U23277 (N_23277,N_21606,N_21200);
or U23278 (N_23278,N_21743,N_19925);
nand U23279 (N_23279,N_20674,N_20488);
or U23280 (N_23280,N_21173,N_20993);
xnor U23281 (N_23281,N_21124,N_19573);
or U23282 (N_23282,N_19929,N_21788);
xor U23283 (N_23283,N_19719,N_21346);
and U23284 (N_23284,N_20806,N_19922);
xnor U23285 (N_23285,N_19681,N_19271);
and U23286 (N_23286,N_20417,N_20943);
nor U23287 (N_23287,N_20483,N_21330);
nor U23288 (N_23288,N_19417,N_20011);
and U23289 (N_23289,N_21688,N_19488);
or U23290 (N_23290,N_21180,N_20763);
or U23291 (N_23291,N_20553,N_20617);
nand U23292 (N_23292,N_20089,N_21867);
xnor U23293 (N_23293,N_21115,N_19409);
xnor U23294 (N_23294,N_20689,N_20447);
nor U23295 (N_23295,N_19781,N_21316);
nor U23296 (N_23296,N_19284,N_21565);
xnor U23297 (N_23297,N_20774,N_21578);
or U23298 (N_23298,N_19524,N_21480);
and U23299 (N_23299,N_20629,N_20141);
nor U23300 (N_23300,N_18889,N_21216);
and U23301 (N_23301,N_21620,N_21476);
or U23302 (N_23302,N_18764,N_19809);
nand U23303 (N_23303,N_19772,N_21532);
or U23304 (N_23304,N_21104,N_20113);
or U23305 (N_23305,N_18921,N_19982);
and U23306 (N_23306,N_19353,N_20792);
nand U23307 (N_23307,N_19200,N_19758);
xnor U23308 (N_23308,N_20504,N_20985);
xor U23309 (N_23309,N_21007,N_19750);
and U23310 (N_23310,N_19051,N_21276);
xor U23311 (N_23311,N_20868,N_19115);
and U23312 (N_23312,N_21082,N_20959);
nand U23313 (N_23313,N_19828,N_19953);
nor U23314 (N_23314,N_21255,N_21426);
or U23315 (N_23315,N_20065,N_21351);
or U23316 (N_23316,N_21106,N_20046);
nor U23317 (N_23317,N_20735,N_19316);
nor U23318 (N_23318,N_21472,N_19513);
or U23319 (N_23319,N_21129,N_20726);
nand U23320 (N_23320,N_19103,N_21662);
or U23321 (N_23321,N_21450,N_21633);
and U23322 (N_23322,N_20757,N_19382);
or U23323 (N_23323,N_20394,N_19523);
nor U23324 (N_23324,N_19793,N_18904);
and U23325 (N_23325,N_21695,N_20599);
nand U23326 (N_23326,N_20858,N_21599);
xnor U23327 (N_23327,N_20420,N_18888);
or U23328 (N_23328,N_21184,N_20745);
nand U23329 (N_23329,N_21146,N_19124);
xnor U23330 (N_23330,N_19191,N_21421);
xor U23331 (N_23331,N_20279,N_20453);
xnor U23332 (N_23332,N_20559,N_20352);
xor U23333 (N_23333,N_19317,N_19399);
xnor U23334 (N_23334,N_21238,N_19304);
and U23335 (N_23335,N_19026,N_21291);
nand U23336 (N_23336,N_19873,N_18785);
nor U23337 (N_23337,N_19079,N_19483);
and U23338 (N_23338,N_19676,N_20913);
or U23339 (N_23339,N_20600,N_19710);
nor U23340 (N_23340,N_19744,N_21816);
or U23341 (N_23341,N_19226,N_20826);
xor U23342 (N_23342,N_20847,N_21183);
nor U23343 (N_23343,N_20201,N_21417);
or U23344 (N_23344,N_19478,N_20632);
and U23345 (N_23345,N_19765,N_21809);
or U23346 (N_23346,N_19815,N_20891);
nor U23347 (N_23347,N_19295,N_21301);
xor U23348 (N_23348,N_21236,N_19967);
nor U23349 (N_23349,N_21153,N_20770);
and U23350 (N_23350,N_20320,N_21348);
or U23351 (N_23351,N_20372,N_19556);
nor U23352 (N_23352,N_21260,N_21393);
and U23353 (N_23353,N_21045,N_20809);
nand U23354 (N_23354,N_18942,N_19313);
nor U23355 (N_23355,N_21415,N_19851);
nor U23356 (N_23356,N_19318,N_20524);
nor U23357 (N_23357,N_19129,N_20425);
xor U23358 (N_23358,N_20551,N_21690);
nand U23359 (N_23359,N_21630,N_19281);
xnor U23360 (N_23360,N_20116,N_21430);
or U23361 (N_23361,N_19866,N_19451);
nor U23362 (N_23362,N_20317,N_19276);
xor U23363 (N_23363,N_20308,N_21143);
or U23364 (N_23364,N_21678,N_20919);
and U23365 (N_23365,N_19414,N_19333);
nand U23366 (N_23366,N_19585,N_20196);
and U23367 (N_23367,N_18951,N_21637);
nor U23368 (N_23368,N_19438,N_18812);
xor U23369 (N_23369,N_21304,N_21521);
xnor U23370 (N_23370,N_21108,N_20615);
nor U23371 (N_23371,N_20569,N_20997);
and U23372 (N_23372,N_20578,N_19155);
xnor U23373 (N_23373,N_19104,N_19563);
nor U23374 (N_23374,N_21101,N_19286);
xor U23375 (N_23375,N_18883,N_20016);
nand U23376 (N_23376,N_21545,N_19491);
and U23377 (N_23377,N_20481,N_20220);
and U23378 (N_23378,N_19448,N_20591);
nor U23379 (N_23379,N_19769,N_19307);
and U23380 (N_23380,N_21841,N_20971);
or U23381 (N_23381,N_20823,N_21821);
and U23382 (N_23382,N_21832,N_21811);
xor U23383 (N_23383,N_21321,N_19450);
nor U23384 (N_23384,N_19369,N_18834);
nand U23385 (N_23385,N_18985,N_19596);
or U23386 (N_23386,N_21528,N_19751);
and U23387 (N_23387,N_20627,N_21639);
or U23388 (N_23388,N_20359,N_21136);
or U23389 (N_23389,N_21087,N_19615);
or U23390 (N_23390,N_21759,N_21477);
or U23391 (N_23391,N_18752,N_20580);
and U23392 (N_23392,N_20007,N_20645);
nor U23393 (N_23393,N_19334,N_20347);
nand U23394 (N_23394,N_19574,N_20748);
xor U23395 (N_23395,N_21300,N_20270);
or U23396 (N_23396,N_19963,N_20136);
nor U23397 (N_23397,N_21247,N_19678);
and U23398 (N_23398,N_19504,N_21170);
nor U23399 (N_23399,N_19263,N_19410);
and U23400 (N_23400,N_19936,N_19151);
nand U23401 (N_23401,N_20415,N_21585);
xor U23402 (N_23402,N_21535,N_19914);
nor U23403 (N_23403,N_21222,N_20885);
or U23404 (N_23404,N_19326,N_19309);
nor U23405 (N_23405,N_19300,N_19506);
nand U23406 (N_23406,N_20828,N_21127);
nor U23407 (N_23407,N_20791,N_21552);
nand U23408 (N_23408,N_19707,N_19132);
xnor U23409 (N_23409,N_19939,N_21600);
nor U23410 (N_23410,N_19391,N_19848);
nor U23411 (N_23411,N_21159,N_19505);
xnor U23412 (N_23412,N_20889,N_19053);
nor U23413 (N_23413,N_20900,N_20723);
or U23414 (N_23414,N_20053,N_20032);
xnor U23415 (N_23415,N_21784,N_21855);
xor U23416 (N_23416,N_21567,N_20259);
xnor U23417 (N_23417,N_19652,N_18916);
nand U23418 (N_23418,N_21659,N_20327);
and U23419 (N_23419,N_20638,N_20152);
or U23420 (N_23420,N_18867,N_18803);
or U23421 (N_23421,N_20222,N_21033);
nor U23422 (N_23422,N_20217,N_21791);
and U23423 (N_23423,N_21345,N_19198);
and U23424 (N_23424,N_19017,N_20471);
nand U23425 (N_23425,N_21691,N_21398);
or U23426 (N_23426,N_20000,N_20766);
xnor U23427 (N_23427,N_19653,N_19869);
nand U23428 (N_23428,N_20445,N_20277);
nor U23429 (N_23429,N_20854,N_18938);
nor U23430 (N_23430,N_20284,N_18897);
nor U23431 (N_23431,N_20915,N_21730);
xnor U23432 (N_23432,N_18963,N_20052);
nor U23433 (N_23433,N_20677,N_18810);
and U23434 (N_23434,N_19308,N_20250);
or U23435 (N_23435,N_20764,N_19282);
and U23436 (N_23436,N_20857,N_21288);
or U23437 (N_23437,N_19131,N_19587);
xnor U23438 (N_23438,N_19817,N_21781);
nand U23439 (N_23439,N_19386,N_21093);
nand U23440 (N_23440,N_19283,N_18867);
xor U23441 (N_23441,N_19094,N_20020);
and U23442 (N_23442,N_20466,N_19512);
nor U23443 (N_23443,N_21407,N_20956);
and U23444 (N_23444,N_19861,N_21311);
nor U23445 (N_23445,N_20612,N_21204);
xor U23446 (N_23446,N_19622,N_19331);
or U23447 (N_23447,N_21544,N_21537);
xnor U23448 (N_23448,N_19125,N_21560);
xor U23449 (N_23449,N_20804,N_18937);
and U23450 (N_23450,N_19213,N_18884);
or U23451 (N_23451,N_18935,N_19370);
nor U23452 (N_23452,N_21502,N_21396);
and U23453 (N_23453,N_20944,N_18856);
nor U23454 (N_23454,N_20656,N_21782);
nor U23455 (N_23455,N_18953,N_19478);
nor U23456 (N_23456,N_19768,N_19789);
xnor U23457 (N_23457,N_19523,N_21407);
and U23458 (N_23458,N_20756,N_19276);
and U23459 (N_23459,N_20236,N_19667);
and U23460 (N_23460,N_20105,N_18889);
nor U23461 (N_23461,N_18856,N_18958);
xnor U23462 (N_23462,N_20265,N_19251);
or U23463 (N_23463,N_19362,N_21316);
or U23464 (N_23464,N_19127,N_19200);
nand U23465 (N_23465,N_21600,N_20369);
xnor U23466 (N_23466,N_21860,N_19975);
nor U23467 (N_23467,N_21002,N_21235);
and U23468 (N_23468,N_19993,N_20911);
nand U23469 (N_23469,N_21377,N_20567);
nand U23470 (N_23470,N_21344,N_20157);
or U23471 (N_23471,N_20730,N_19399);
nand U23472 (N_23472,N_19031,N_20898);
and U23473 (N_23473,N_18890,N_19909);
or U23474 (N_23474,N_20710,N_18888);
and U23475 (N_23475,N_18814,N_19513);
or U23476 (N_23476,N_19860,N_20701);
xnor U23477 (N_23477,N_20028,N_19046);
and U23478 (N_23478,N_19933,N_20439);
or U23479 (N_23479,N_21491,N_18762);
or U23480 (N_23480,N_18946,N_20690);
nand U23481 (N_23481,N_21321,N_20828);
nand U23482 (N_23482,N_18831,N_20568);
and U23483 (N_23483,N_19171,N_19565);
xor U23484 (N_23484,N_19826,N_21519);
nand U23485 (N_23485,N_19096,N_20203);
nor U23486 (N_23486,N_20732,N_19097);
or U23487 (N_23487,N_20166,N_20928);
and U23488 (N_23488,N_20371,N_21489);
xnor U23489 (N_23489,N_21719,N_20353);
xnor U23490 (N_23490,N_21792,N_21611);
and U23491 (N_23491,N_20318,N_19084);
or U23492 (N_23492,N_19069,N_20023);
or U23493 (N_23493,N_21678,N_19576);
xor U23494 (N_23494,N_19359,N_19050);
xor U23495 (N_23495,N_21668,N_20146);
xor U23496 (N_23496,N_20791,N_21870);
or U23497 (N_23497,N_20923,N_20051);
nor U23498 (N_23498,N_21475,N_21423);
nor U23499 (N_23499,N_21383,N_21284);
nor U23500 (N_23500,N_20805,N_19324);
nor U23501 (N_23501,N_19982,N_21829);
and U23502 (N_23502,N_21642,N_20224);
nand U23503 (N_23503,N_19847,N_19000);
nor U23504 (N_23504,N_20915,N_19497);
nand U23505 (N_23505,N_20073,N_20194);
or U23506 (N_23506,N_21048,N_20657);
and U23507 (N_23507,N_20245,N_18953);
nor U23508 (N_23508,N_20878,N_20090);
xnor U23509 (N_23509,N_21785,N_20693);
nand U23510 (N_23510,N_20891,N_20310);
or U23511 (N_23511,N_19733,N_19630);
or U23512 (N_23512,N_20694,N_19350);
xor U23513 (N_23513,N_21118,N_21562);
nand U23514 (N_23514,N_19449,N_20761);
xnor U23515 (N_23515,N_19820,N_19918);
nor U23516 (N_23516,N_20711,N_21584);
nor U23517 (N_23517,N_21565,N_18878);
and U23518 (N_23518,N_21276,N_21787);
and U23519 (N_23519,N_21543,N_19959);
and U23520 (N_23520,N_21448,N_21455);
nand U23521 (N_23521,N_20935,N_20079);
and U23522 (N_23522,N_20839,N_21749);
or U23523 (N_23523,N_18812,N_19998);
nand U23524 (N_23524,N_20015,N_20229);
xnor U23525 (N_23525,N_21146,N_21866);
nand U23526 (N_23526,N_21005,N_21835);
and U23527 (N_23527,N_19348,N_21802);
and U23528 (N_23528,N_20103,N_20763);
nand U23529 (N_23529,N_20597,N_19507);
nor U23530 (N_23530,N_21220,N_20031);
nor U23531 (N_23531,N_21742,N_21490);
nand U23532 (N_23532,N_21864,N_20764);
nor U23533 (N_23533,N_21740,N_18844);
and U23534 (N_23534,N_21419,N_19424);
and U23535 (N_23535,N_21114,N_20039);
nor U23536 (N_23536,N_21498,N_19904);
or U23537 (N_23537,N_19547,N_20034);
nor U23538 (N_23538,N_19121,N_19003);
and U23539 (N_23539,N_21689,N_19388);
nand U23540 (N_23540,N_19318,N_19160);
nor U23541 (N_23541,N_19758,N_19359);
nor U23542 (N_23542,N_20734,N_21210);
and U23543 (N_23543,N_18764,N_19531);
nand U23544 (N_23544,N_19756,N_21394);
and U23545 (N_23545,N_21045,N_19010);
nand U23546 (N_23546,N_20034,N_20858);
xor U23547 (N_23547,N_19923,N_18826);
and U23548 (N_23548,N_19381,N_21326);
xor U23549 (N_23549,N_20403,N_21852);
or U23550 (N_23550,N_19339,N_20555);
nand U23551 (N_23551,N_19231,N_19397);
nor U23552 (N_23552,N_19399,N_21101);
xor U23553 (N_23553,N_19758,N_20088);
nand U23554 (N_23554,N_21258,N_18761);
nor U23555 (N_23555,N_19950,N_21189);
xor U23556 (N_23556,N_19213,N_20942);
xor U23557 (N_23557,N_20548,N_21562);
and U23558 (N_23558,N_18975,N_21644);
nor U23559 (N_23559,N_21515,N_20660);
xnor U23560 (N_23560,N_18762,N_19712);
nand U23561 (N_23561,N_19771,N_21227);
nor U23562 (N_23562,N_20576,N_20111);
nor U23563 (N_23563,N_21099,N_21592);
or U23564 (N_23564,N_19764,N_21299);
or U23565 (N_23565,N_19844,N_20705);
nor U23566 (N_23566,N_21005,N_19639);
or U23567 (N_23567,N_20985,N_21618);
nor U23568 (N_23568,N_19038,N_19196);
and U23569 (N_23569,N_18962,N_18928);
xnor U23570 (N_23570,N_21681,N_19463);
nand U23571 (N_23571,N_20688,N_18847);
nand U23572 (N_23572,N_20891,N_19203);
or U23573 (N_23573,N_20446,N_21126);
or U23574 (N_23574,N_18921,N_20962);
and U23575 (N_23575,N_19602,N_21553);
or U23576 (N_23576,N_21145,N_21198);
nor U23577 (N_23577,N_19651,N_21612);
and U23578 (N_23578,N_21114,N_21058);
nor U23579 (N_23579,N_20158,N_19443);
and U23580 (N_23580,N_21626,N_19773);
nor U23581 (N_23581,N_20719,N_20789);
xnor U23582 (N_23582,N_19448,N_21476);
nand U23583 (N_23583,N_21126,N_19397);
or U23584 (N_23584,N_21415,N_20189);
or U23585 (N_23585,N_21377,N_19403);
xor U23586 (N_23586,N_20909,N_18956);
and U23587 (N_23587,N_19435,N_20160);
xor U23588 (N_23588,N_20226,N_19486);
xnor U23589 (N_23589,N_20490,N_21656);
nor U23590 (N_23590,N_20968,N_19549);
or U23591 (N_23591,N_19515,N_20738);
nand U23592 (N_23592,N_19677,N_20277);
nand U23593 (N_23593,N_19918,N_20397);
or U23594 (N_23594,N_21629,N_19998);
nor U23595 (N_23595,N_19695,N_19136);
or U23596 (N_23596,N_20563,N_21054);
xnor U23597 (N_23597,N_21569,N_21465);
nor U23598 (N_23598,N_21389,N_19387);
nand U23599 (N_23599,N_20684,N_20692);
and U23600 (N_23600,N_19144,N_20843);
nor U23601 (N_23601,N_21608,N_21371);
nand U23602 (N_23602,N_19633,N_19387);
or U23603 (N_23603,N_20954,N_19250);
or U23604 (N_23604,N_20238,N_19686);
or U23605 (N_23605,N_20673,N_19081);
nand U23606 (N_23606,N_20131,N_20975);
nor U23607 (N_23607,N_19202,N_20785);
nand U23608 (N_23608,N_18847,N_20263);
and U23609 (N_23609,N_18887,N_18754);
and U23610 (N_23610,N_21698,N_21556);
or U23611 (N_23611,N_18768,N_21680);
nand U23612 (N_23612,N_20374,N_19095);
nor U23613 (N_23613,N_21549,N_21459);
nand U23614 (N_23614,N_19949,N_18999);
or U23615 (N_23615,N_20496,N_21627);
and U23616 (N_23616,N_20760,N_20821);
xnor U23617 (N_23617,N_19379,N_19042);
and U23618 (N_23618,N_18904,N_21841);
nand U23619 (N_23619,N_19141,N_19801);
and U23620 (N_23620,N_19322,N_20116);
or U23621 (N_23621,N_19065,N_20654);
or U23622 (N_23622,N_21743,N_20979);
nor U23623 (N_23623,N_18990,N_20142);
nand U23624 (N_23624,N_21388,N_19641);
and U23625 (N_23625,N_19882,N_20277);
nand U23626 (N_23626,N_19135,N_21261);
nor U23627 (N_23627,N_19359,N_19296);
or U23628 (N_23628,N_19378,N_21834);
nand U23629 (N_23629,N_21635,N_20100);
nand U23630 (N_23630,N_20462,N_21846);
xor U23631 (N_23631,N_19061,N_19474);
nand U23632 (N_23632,N_19804,N_18970);
or U23633 (N_23633,N_19005,N_18985);
xnor U23634 (N_23634,N_19329,N_20371);
xor U23635 (N_23635,N_19318,N_19215);
or U23636 (N_23636,N_18821,N_21327);
and U23637 (N_23637,N_19329,N_20617);
nand U23638 (N_23638,N_20415,N_21377);
nor U23639 (N_23639,N_20904,N_21601);
xnor U23640 (N_23640,N_21259,N_21720);
and U23641 (N_23641,N_19241,N_18807);
xnor U23642 (N_23642,N_21361,N_21532);
xnor U23643 (N_23643,N_19134,N_18954);
xor U23644 (N_23644,N_21729,N_21544);
or U23645 (N_23645,N_21106,N_19671);
nor U23646 (N_23646,N_21203,N_21473);
or U23647 (N_23647,N_20777,N_20623);
nand U23648 (N_23648,N_20971,N_18761);
xnor U23649 (N_23649,N_20527,N_21530);
or U23650 (N_23650,N_21341,N_19420);
xor U23651 (N_23651,N_20779,N_21612);
nand U23652 (N_23652,N_20625,N_21546);
and U23653 (N_23653,N_21532,N_20267);
or U23654 (N_23654,N_18941,N_21548);
and U23655 (N_23655,N_20375,N_19950);
nand U23656 (N_23656,N_21477,N_19731);
nor U23657 (N_23657,N_20145,N_19890);
and U23658 (N_23658,N_21686,N_20541);
nor U23659 (N_23659,N_21080,N_19258);
and U23660 (N_23660,N_20669,N_18843);
xor U23661 (N_23661,N_21495,N_21708);
or U23662 (N_23662,N_19467,N_21145);
nand U23663 (N_23663,N_19223,N_21268);
and U23664 (N_23664,N_21848,N_20535);
nor U23665 (N_23665,N_19546,N_20345);
or U23666 (N_23666,N_19433,N_21536);
and U23667 (N_23667,N_19652,N_19051);
or U23668 (N_23668,N_20573,N_19894);
nand U23669 (N_23669,N_20428,N_21643);
xor U23670 (N_23670,N_18853,N_19933);
xnor U23671 (N_23671,N_18924,N_21364);
nor U23672 (N_23672,N_20047,N_20264);
nor U23673 (N_23673,N_21450,N_21651);
nand U23674 (N_23674,N_21379,N_19438);
nand U23675 (N_23675,N_20858,N_19431);
xnor U23676 (N_23676,N_20396,N_20925);
xor U23677 (N_23677,N_21575,N_19472);
nor U23678 (N_23678,N_18793,N_18882);
or U23679 (N_23679,N_18769,N_21523);
nor U23680 (N_23680,N_21730,N_19844);
nor U23681 (N_23681,N_21048,N_21417);
or U23682 (N_23682,N_20127,N_20407);
or U23683 (N_23683,N_19403,N_19058);
nor U23684 (N_23684,N_20509,N_21198);
or U23685 (N_23685,N_19108,N_19336);
nand U23686 (N_23686,N_21026,N_21012);
or U23687 (N_23687,N_19470,N_21067);
or U23688 (N_23688,N_21058,N_19942);
xnor U23689 (N_23689,N_21144,N_19538);
nor U23690 (N_23690,N_21103,N_20308);
nand U23691 (N_23691,N_18781,N_21658);
xnor U23692 (N_23692,N_21445,N_21389);
or U23693 (N_23693,N_20801,N_21175);
nor U23694 (N_23694,N_19432,N_20843);
or U23695 (N_23695,N_20739,N_20570);
nor U23696 (N_23696,N_20874,N_21062);
nor U23697 (N_23697,N_21349,N_18936);
xnor U23698 (N_23698,N_21551,N_19188);
nor U23699 (N_23699,N_20680,N_20797);
xor U23700 (N_23700,N_21007,N_20665);
or U23701 (N_23701,N_21219,N_21283);
and U23702 (N_23702,N_19996,N_21691);
nor U23703 (N_23703,N_20151,N_20977);
or U23704 (N_23704,N_20239,N_20516);
nor U23705 (N_23705,N_21860,N_21133);
and U23706 (N_23706,N_19764,N_21223);
nor U23707 (N_23707,N_21712,N_19843);
xnor U23708 (N_23708,N_20846,N_20594);
and U23709 (N_23709,N_21599,N_19380);
nand U23710 (N_23710,N_20613,N_19174);
xor U23711 (N_23711,N_19646,N_20376);
and U23712 (N_23712,N_19864,N_20621);
nand U23713 (N_23713,N_20848,N_19249);
or U23714 (N_23714,N_20788,N_20695);
and U23715 (N_23715,N_20472,N_21321);
xor U23716 (N_23716,N_19484,N_20022);
or U23717 (N_23717,N_21052,N_20447);
nand U23718 (N_23718,N_20977,N_19754);
and U23719 (N_23719,N_20509,N_19429);
or U23720 (N_23720,N_21620,N_20665);
or U23721 (N_23721,N_21757,N_21065);
nand U23722 (N_23722,N_21715,N_20894);
xnor U23723 (N_23723,N_21350,N_19966);
nor U23724 (N_23724,N_20453,N_21760);
nand U23725 (N_23725,N_19905,N_18804);
xnor U23726 (N_23726,N_19832,N_19940);
nand U23727 (N_23727,N_21286,N_19861);
and U23728 (N_23728,N_21510,N_19409);
and U23729 (N_23729,N_20624,N_20979);
nand U23730 (N_23730,N_20535,N_21691);
and U23731 (N_23731,N_21398,N_21727);
xnor U23732 (N_23732,N_21227,N_19481);
or U23733 (N_23733,N_19392,N_18892);
and U23734 (N_23734,N_20360,N_19363);
or U23735 (N_23735,N_18889,N_19865);
and U23736 (N_23736,N_19818,N_20489);
or U23737 (N_23737,N_21082,N_21264);
xor U23738 (N_23738,N_19586,N_21526);
and U23739 (N_23739,N_18813,N_19534);
nand U23740 (N_23740,N_19046,N_20657);
xnor U23741 (N_23741,N_20958,N_19662);
xnor U23742 (N_23742,N_21260,N_19088);
or U23743 (N_23743,N_20093,N_20442);
nor U23744 (N_23744,N_20803,N_20778);
xnor U23745 (N_23745,N_21663,N_21395);
and U23746 (N_23746,N_21341,N_18833);
nor U23747 (N_23747,N_19906,N_19945);
nor U23748 (N_23748,N_19512,N_19820);
nand U23749 (N_23749,N_19227,N_21060);
nor U23750 (N_23750,N_21793,N_19006);
nand U23751 (N_23751,N_19410,N_20107);
or U23752 (N_23752,N_21178,N_20943);
nor U23753 (N_23753,N_20138,N_19201);
nand U23754 (N_23754,N_21135,N_19080);
and U23755 (N_23755,N_19551,N_19973);
and U23756 (N_23756,N_21378,N_18789);
or U23757 (N_23757,N_20101,N_19107);
nand U23758 (N_23758,N_21355,N_21295);
nor U23759 (N_23759,N_21629,N_19684);
nand U23760 (N_23760,N_19960,N_18765);
and U23761 (N_23761,N_20117,N_20034);
nor U23762 (N_23762,N_19181,N_21838);
or U23763 (N_23763,N_21362,N_18847);
nor U23764 (N_23764,N_19409,N_20966);
xor U23765 (N_23765,N_18771,N_20120);
xnor U23766 (N_23766,N_20970,N_20416);
and U23767 (N_23767,N_21495,N_21786);
nor U23768 (N_23768,N_19312,N_19419);
nor U23769 (N_23769,N_19167,N_20812);
and U23770 (N_23770,N_20829,N_19835);
nand U23771 (N_23771,N_19814,N_19025);
or U23772 (N_23772,N_19695,N_18795);
nand U23773 (N_23773,N_20169,N_19998);
and U23774 (N_23774,N_19422,N_20085);
nand U23775 (N_23775,N_20635,N_20259);
and U23776 (N_23776,N_20149,N_20868);
nand U23777 (N_23777,N_19112,N_20505);
nor U23778 (N_23778,N_21869,N_20015);
or U23779 (N_23779,N_19060,N_19822);
nand U23780 (N_23780,N_20812,N_21009);
xnor U23781 (N_23781,N_21154,N_21160);
and U23782 (N_23782,N_18845,N_21511);
nand U23783 (N_23783,N_20031,N_19287);
and U23784 (N_23784,N_20595,N_19427);
nor U23785 (N_23785,N_20497,N_19706);
nand U23786 (N_23786,N_19126,N_20082);
nand U23787 (N_23787,N_20094,N_21495);
nand U23788 (N_23788,N_19844,N_21178);
and U23789 (N_23789,N_19685,N_18832);
or U23790 (N_23790,N_18825,N_19779);
or U23791 (N_23791,N_18968,N_21166);
and U23792 (N_23792,N_19120,N_21638);
or U23793 (N_23793,N_19142,N_19956);
and U23794 (N_23794,N_19493,N_21232);
nand U23795 (N_23795,N_21227,N_19144);
xor U23796 (N_23796,N_21248,N_19418);
and U23797 (N_23797,N_20734,N_19772);
nor U23798 (N_23798,N_18864,N_20089);
or U23799 (N_23799,N_20320,N_21649);
nor U23800 (N_23800,N_21373,N_20684);
xnor U23801 (N_23801,N_21851,N_19250);
nand U23802 (N_23802,N_19988,N_19262);
and U23803 (N_23803,N_21517,N_20999);
or U23804 (N_23804,N_20310,N_19929);
nand U23805 (N_23805,N_21010,N_19263);
or U23806 (N_23806,N_20361,N_19489);
nor U23807 (N_23807,N_20560,N_21669);
xnor U23808 (N_23808,N_20749,N_20321);
nor U23809 (N_23809,N_20397,N_21788);
xnor U23810 (N_23810,N_19015,N_20899);
or U23811 (N_23811,N_21720,N_19519);
xnor U23812 (N_23812,N_20388,N_21532);
or U23813 (N_23813,N_19866,N_21229);
and U23814 (N_23814,N_21621,N_19729);
or U23815 (N_23815,N_20252,N_19000);
or U23816 (N_23816,N_20938,N_21476);
or U23817 (N_23817,N_19339,N_19475);
nand U23818 (N_23818,N_19890,N_19664);
xnor U23819 (N_23819,N_21743,N_21060);
and U23820 (N_23820,N_20996,N_20377);
and U23821 (N_23821,N_20641,N_21840);
or U23822 (N_23822,N_20554,N_19202);
nand U23823 (N_23823,N_21184,N_19820);
or U23824 (N_23824,N_21811,N_19394);
or U23825 (N_23825,N_20924,N_21309);
nand U23826 (N_23826,N_18805,N_19090);
nor U23827 (N_23827,N_19492,N_19644);
nor U23828 (N_23828,N_21041,N_21829);
or U23829 (N_23829,N_21812,N_19526);
and U23830 (N_23830,N_21305,N_21844);
nand U23831 (N_23831,N_19645,N_20054);
nor U23832 (N_23832,N_20061,N_21554);
nand U23833 (N_23833,N_19491,N_19936);
nand U23834 (N_23834,N_19420,N_21135);
or U23835 (N_23835,N_19996,N_19929);
xnor U23836 (N_23836,N_19876,N_20235);
xor U23837 (N_23837,N_21696,N_21207);
nand U23838 (N_23838,N_19710,N_21443);
nor U23839 (N_23839,N_20539,N_19332);
nand U23840 (N_23840,N_18877,N_18978);
or U23841 (N_23841,N_21088,N_18771);
or U23842 (N_23842,N_19538,N_20937);
xor U23843 (N_23843,N_19146,N_21256);
nand U23844 (N_23844,N_21046,N_19712);
or U23845 (N_23845,N_20885,N_19050);
xor U23846 (N_23846,N_18757,N_19407);
nor U23847 (N_23847,N_18977,N_19436);
nand U23848 (N_23848,N_20968,N_20479);
xnor U23849 (N_23849,N_20730,N_19197);
and U23850 (N_23850,N_21701,N_19232);
nor U23851 (N_23851,N_20703,N_20188);
and U23852 (N_23852,N_19288,N_19944);
or U23853 (N_23853,N_19209,N_19576);
nand U23854 (N_23854,N_20876,N_18817);
or U23855 (N_23855,N_20430,N_19718);
nand U23856 (N_23856,N_20488,N_18874);
or U23857 (N_23857,N_20996,N_20988);
and U23858 (N_23858,N_19676,N_19521);
nor U23859 (N_23859,N_19577,N_19958);
or U23860 (N_23860,N_20786,N_20483);
or U23861 (N_23861,N_20673,N_19283);
xnor U23862 (N_23862,N_20894,N_20727);
or U23863 (N_23863,N_21815,N_20126);
xor U23864 (N_23864,N_20467,N_20179);
or U23865 (N_23865,N_21492,N_19128);
nand U23866 (N_23866,N_19071,N_20200);
xnor U23867 (N_23867,N_18969,N_19289);
or U23868 (N_23868,N_19677,N_19243);
and U23869 (N_23869,N_21581,N_21739);
xnor U23870 (N_23870,N_21566,N_19177);
nand U23871 (N_23871,N_21135,N_21308);
or U23872 (N_23872,N_21569,N_20908);
or U23873 (N_23873,N_18990,N_19041);
or U23874 (N_23874,N_19538,N_20559);
xnor U23875 (N_23875,N_19467,N_21690);
and U23876 (N_23876,N_20182,N_21421);
nand U23877 (N_23877,N_20841,N_20942);
and U23878 (N_23878,N_19821,N_21083);
and U23879 (N_23879,N_19797,N_19851);
and U23880 (N_23880,N_19085,N_21674);
and U23881 (N_23881,N_21060,N_19942);
or U23882 (N_23882,N_21607,N_20082);
or U23883 (N_23883,N_18771,N_21294);
nand U23884 (N_23884,N_21150,N_21321);
or U23885 (N_23885,N_20344,N_20312);
xnor U23886 (N_23886,N_21418,N_20961);
xnor U23887 (N_23887,N_20525,N_19229);
or U23888 (N_23888,N_19971,N_20422);
nand U23889 (N_23889,N_21267,N_21207);
or U23890 (N_23890,N_21007,N_20925);
and U23891 (N_23891,N_21655,N_19236);
and U23892 (N_23892,N_19457,N_19458);
and U23893 (N_23893,N_18860,N_20725);
nand U23894 (N_23894,N_21400,N_21075);
and U23895 (N_23895,N_21169,N_19719);
or U23896 (N_23896,N_19403,N_19292);
and U23897 (N_23897,N_19164,N_18788);
nand U23898 (N_23898,N_18874,N_20219);
or U23899 (N_23899,N_20634,N_21287);
nand U23900 (N_23900,N_20613,N_20219);
xor U23901 (N_23901,N_18995,N_19574);
or U23902 (N_23902,N_20759,N_19414);
and U23903 (N_23903,N_19597,N_19875);
nand U23904 (N_23904,N_20064,N_19943);
nand U23905 (N_23905,N_19924,N_18939);
or U23906 (N_23906,N_21639,N_19831);
or U23907 (N_23907,N_21227,N_21001);
or U23908 (N_23908,N_18763,N_20074);
nand U23909 (N_23909,N_19649,N_19064);
nor U23910 (N_23910,N_20137,N_21195);
nor U23911 (N_23911,N_21838,N_19378);
and U23912 (N_23912,N_19077,N_19234);
nand U23913 (N_23913,N_19799,N_19490);
or U23914 (N_23914,N_19460,N_21544);
and U23915 (N_23915,N_20342,N_18871);
and U23916 (N_23916,N_20513,N_19327);
nor U23917 (N_23917,N_19075,N_20350);
and U23918 (N_23918,N_18826,N_20673);
nand U23919 (N_23919,N_20890,N_21115);
nand U23920 (N_23920,N_20918,N_18821);
or U23921 (N_23921,N_20673,N_19755);
and U23922 (N_23922,N_21089,N_21111);
nor U23923 (N_23923,N_21445,N_19858);
xnor U23924 (N_23924,N_18861,N_19543);
or U23925 (N_23925,N_19592,N_18960);
nand U23926 (N_23926,N_19592,N_19454);
xnor U23927 (N_23927,N_19368,N_18987);
nand U23928 (N_23928,N_20962,N_21004);
or U23929 (N_23929,N_18922,N_19332);
nor U23930 (N_23930,N_20943,N_21842);
xnor U23931 (N_23931,N_19377,N_21313);
and U23932 (N_23932,N_21556,N_19991);
and U23933 (N_23933,N_19986,N_18980);
and U23934 (N_23934,N_20446,N_20819);
nand U23935 (N_23935,N_19823,N_19004);
xor U23936 (N_23936,N_19919,N_20797);
nand U23937 (N_23937,N_20138,N_20624);
xnor U23938 (N_23938,N_18834,N_21222);
and U23939 (N_23939,N_21202,N_18806);
xor U23940 (N_23940,N_21305,N_19616);
or U23941 (N_23941,N_18834,N_20022);
nand U23942 (N_23942,N_19379,N_19631);
xor U23943 (N_23943,N_20080,N_21702);
nor U23944 (N_23944,N_20202,N_19337);
nor U23945 (N_23945,N_19764,N_21277);
nand U23946 (N_23946,N_19986,N_21535);
nand U23947 (N_23947,N_18990,N_19215);
and U23948 (N_23948,N_19591,N_21371);
nor U23949 (N_23949,N_19342,N_19561);
xor U23950 (N_23950,N_19094,N_21396);
or U23951 (N_23951,N_19052,N_21287);
nand U23952 (N_23952,N_21317,N_20472);
nor U23953 (N_23953,N_21088,N_20943);
and U23954 (N_23954,N_20711,N_21119);
or U23955 (N_23955,N_20349,N_21439);
nand U23956 (N_23956,N_21345,N_19532);
nor U23957 (N_23957,N_20774,N_20524);
and U23958 (N_23958,N_21140,N_19255);
xor U23959 (N_23959,N_20988,N_19179);
nor U23960 (N_23960,N_19233,N_20577);
nand U23961 (N_23961,N_21505,N_19878);
and U23962 (N_23962,N_21579,N_20241);
nand U23963 (N_23963,N_21448,N_21513);
or U23964 (N_23964,N_20382,N_20166);
nand U23965 (N_23965,N_19230,N_18771);
or U23966 (N_23966,N_18859,N_20540);
nand U23967 (N_23967,N_19364,N_19459);
or U23968 (N_23968,N_21448,N_19114);
and U23969 (N_23969,N_21369,N_19032);
and U23970 (N_23970,N_20178,N_21835);
nor U23971 (N_23971,N_19543,N_20030);
nor U23972 (N_23972,N_21816,N_21523);
or U23973 (N_23973,N_18878,N_19383);
or U23974 (N_23974,N_21481,N_18891);
and U23975 (N_23975,N_21095,N_19750);
and U23976 (N_23976,N_19837,N_20577);
nand U23977 (N_23977,N_20722,N_21566);
xnor U23978 (N_23978,N_19244,N_21227);
and U23979 (N_23979,N_20096,N_21265);
xnor U23980 (N_23980,N_20258,N_21504);
nor U23981 (N_23981,N_19928,N_19044);
xor U23982 (N_23982,N_20674,N_19493);
and U23983 (N_23983,N_20853,N_21292);
nand U23984 (N_23984,N_20341,N_20005);
xor U23985 (N_23985,N_21259,N_19668);
and U23986 (N_23986,N_20521,N_19991);
or U23987 (N_23987,N_18761,N_20580);
xor U23988 (N_23988,N_19143,N_19147);
and U23989 (N_23989,N_18752,N_19311);
nand U23990 (N_23990,N_19651,N_19545);
and U23991 (N_23991,N_21025,N_20147);
and U23992 (N_23992,N_20808,N_21442);
or U23993 (N_23993,N_20702,N_19513);
nor U23994 (N_23994,N_20890,N_21265);
nor U23995 (N_23995,N_20950,N_20617);
xor U23996 (N_23996,N_18959,N_18892);
or U23997 (N_23997,N_19013,N_21294);
xnor U23998 (N_23998,N_21774,N_21102);
and U23999 (N_23999,N_21837,N_20196);
xor U24000 (N_24000,N_19152,N_19765);
nand U24001 (N_24001,N_21017,N_19990);
nor U24002 (N_24002,N_20480,N_21550);
and U24003 (N_24003,N_18930,N_21510);
xor U24004 (N_24004,N_21734,N_18809);
or U24005 (N_24005,N_19916,N_20901);
and U24006 (N_24006,N_19132,N_20164);
xnor U24007 (N_24007,N_20991,N_18795);
and U24008 (N_24008,N_19560,N_21831);
nor U24009 (N_24009,N_18989,N_19171);
and U24010 (N_24010,N_19213,N_19824);
nand U24011 (N_24011,N_21537,N_21644);
nor U24012 (N_24012,N_19897,N_19456);
and U24013 (N_24013,N_19350,N_20190);
or U24014 (N_24014,N_20992,N_21573);
xnor U24015 (N_24015,N_19249,N_19799);
xor U24016 (N_24016,N_19522,N_21868);
nand U24017 (N_24017,N_19795,N_19047);
nand U24018 (N_24018,N_20694,N_19812);
nor U24019 (N_24019,N_21496,N_21811);
nor U24020 (N_24020,N_21409,N_19455);
xnor U24021 (N_24021,N_19763,N_19771);
and U24022 (N_24022,N_18963,N_20705);
xnor U24023 (N_24023,N_20388,N_20399);
nand U24024 (N_24024,N_18891,N_21117);
nand U24025 (N_24025,N_20556,N_20178);
nand U24026 (N_24026,N_19409,N_20287);
nand U24027 (N_24027,N_21660,N_19283);
nor U24028 (N_24028,N_21309,N_19489);
xnor U24029 (N_24029,N_19048,N_20015);
nor U24030 (N_24030,N_20085,N_19049);
and U24031 (N_24031,N_18768,N_20757);
or U24032 (N_24032,N_19589,N_21228);
and U24033 (N_24033,N_20380,N_20625);
nand U24034 (N_24034,N_20565,N_19211);
xor U24035 (N_24035,N_18934,N_19202);
nor U24036 (N_24036,N_21009,N_20598);
and U24037 (N_24037,N_20682,N_21034);
or U24038 (N_24038,N_18902,N_21332);
xor U24039 (N_24039,N_21087,N_20505);
nor U24040 (N_24040,N_20059,N_20756);
and U24041 (N_24041,N_18788,N_20858);
nand U24042 (N_24042,N_20009,N_21586);
xnor U24043 (N_24043,N_20971,N_21856);
nand U24044 (N_24044,N_21276,N_21601);
and U24045 (N_24045,N_20702,N_20088);
and U24046 (N_24046,N_20293,N_20114);
nand U24047 (N_24047,N_19674,N_18948);
xor U24048 (N_24048,N_21662,N_20334);
or U24049 (N_24049,N_18917,N_20550);
nor U24050 (N_24050,N_21164,N_20511);
or U24051 (N_24051,N_20611,N_19118);
and U24052 (N_24052,N_20406,N_19634);
nor U24053 (N_24053,N_19212,N_18894);
xnor U24054 (N_24054,N_21478,N_20346);
or U24055 (N_24055,N_20836,N_19781);
xnor U24056 (N_24056,N_19175,N_20895);
or U24057 (N_24057,N_21637,N_20948);
nor U24058 (N_24058,N_20543,N_19719);
xor U24059 (N_24059,N_20092,N_21301);
and U24060 (N_24060,N_21429,N_21009);
nor U24061 (N_24061,N_21393,N_20956);
and U24062 (N_24062,N_20121,N_19668);
and U24063 (N_24063,N_19988,N_20478);
nor U24064 (N_24064,N_19413,N_20509);
nand U24065 (N_24065,N_21088,N_18774);
nor U24066 (N_24066,N_20756,N_20057);
nand U24067 (N_24067,N_21506,N_21647);
xnor U24068 (N_24068,N_20992,N_19824);
nand U24069 (N_24069,N_20473,N_20729);
or U24070 (N_24070,N_20901,N_19096);
nor U24071 (N_24071,N_19805,N_21058);
nor U24072 (N_24072,N_19483,N_21758);
or U24073 (N_24073,N_20360,N_19778);
xor U24074 (N_24074,N_20567,N_21210);
nand U24075 (N_24075,N_20099,N_19684);
nor U24076 (N_24076,N_21539,N_20595);
nor U24077 (N_24077,N_19811,N_19983);
nor U24078 (N_24078,N_19853,N_18795);
and U24079 (N_24079,N_20436,N_21211);
nand U24080 (N_24080,N_20781,N_21359);
nor U24081 (N_24081,N_20633,N_20036);
nor U24082 (N_24082,N_20612,N_19592);
nand U24083 (N_24083,N_20640,N_19689);
nor U24084 (N_24084,N_18872,N_20390);
xnor U24085 (N_24085,N_19623,N_19027);
or U24086 (N_24086,N_20326,N_20984);
nand U24087 (N_24087,N_20837,N_21345);
or U24088 (N_24088,N_20400,N_20196);
or U24089 (N_24089,N_21231,N_19241);
nor U24090 (N_24090,N_20433,N_21393);
nor U24091 (N_24091,N_21529,N_19990);
xnor U24092 (N_24092,N_21053,N_20436);
nand U24093 (N_24093,N_20681,N_21759);
nor U24094 (N_24094,N_19474,N_18750);
nand U24095 (N_24095,N_20164,N_18978);
xnor U24096 (N_24096,N_19069,N_19512);
or U24097 (N_24097,N_20264,N_19933);
xor U24098 (N_24098,N_19589,N_18984);
or U24099 (N_24099,N_18873,N_20943);
xnor U24100 (N_24100,N_21414,N_19029);
nand U24101 (N_24101,N_20883,N_19233);
nor U24102 (N_24102,N_20570,N_20530);
nor U24103 (N_24103,N_20082,N_18993);
nor U24104 (N_24104,N_20400,N_19853);
or U24105 (N_24105,N_20353,N_21143);
nand U24106 (N_24106,N_21187,N_19646);
nand U24107 (N_24107,N_19743,N_19982);
nor U24108 (N_24108,N_21222,N_21192);
nand U24109 (N_24109,N_19461,N_19999);
nor U24110 (N_24110,N_19998,N_20758);
or U24111 (N_24111,N_20906,N_19083);
and U24112 (N_24112,N_21509,N_21445);
nor U24113 (N_24113,N_19994,N_21265);
nor U24114 (N_24114,N_21766,N_20809);
or U24115 (N_24115,N_21300,N_21592);
or U24116 (N_24116,N_21714,N_19498);
xor U24117 (N_24117,N_18901,N_20891);
xor U24118 (N_24118,N_20478,N_20918);
and U24119 (N_24119,N_21412,N_21511);
and U24120 (N_24120,N_21853,N_21712);
xor U24121 (N_24121,N_19969,N_21301);
or U24122 (N_24122,N_20278,N_19366);
nor U24123 (N_24123,N_19492,N_21250);
and U24124 (N_24124,N_20835,N_20142);
and U24125 (N_24125,N_21310,N_21644);
xor U24126 (N_24126,N_21277,N_21323);
xnor U24127 (N_24127,N_21790,N_18820);
xnor U24128 (N_24128,N_19941,N_21830);
or U24129 (N_24129,N_20777,N_18811);
nor U24130 (N_24130,N_21069,N_21558);
xor U24131 (N_24131,N_20323,N_20274);
nor U24132 (N_24132,N_19250,N_20025);
or U24133 (N_24133,N_20725,N_20653);
nand U24134 (N_24134,N_19294,N_18965);
nor U24135 (N_24135,N_19308,N_19560);
nor U24136 (N_24136,N_19619,N_19472);
nand U24137 (N_24137,N_20765,N_19024);
nor U24138 (N_24138,N_20782,N_18992);
xor U24139 (N_24139,N_19767,N_21090);
nand U24140 (N_24140,N_21705,N_20451);
nand U24141 (N_24141,N_21273,N_19490);
xnor U24142 (N_24142,N_19993,N_20323);
nand U24143 (N_24143,N_21378,N_18849);
and U24144 (N_24144,N_18848,N_20111);
or U24145 (N_24145,N_19190,N_21626);
nor U24146 (N_24146,N_19285,N_20120);
or U24147 (N_24147,N_20829,N_21471);
nor U24148 (N_24148,N_19654,N_21731);
nor U24149 (N_24149,N_19578,N_19929);
nand U24150 (N_24150,N_20623,N_18857);
nor U24151 (N_24151,N_19799,N_19977);
nor U24152 (N_24152,N_20275,N_20218);
nand U24153 (N_24153,N_21578,N_20671);
or U24154 (N_24154,N_21368,N_21502);
nand U24155 (N_24155,N_21281,N_19301);
and U24156 (N_24156,N_21055,N_19601);
or U24157 (N_24157,N_20259,N_21486);
nor U24158 (N_24158,N_21464,N_21746);
or U24159 (N_24159,N_19969,N_19175);
nand U24160 (N_24160,N_19849,N_20683);
xor U24161 (N_24161,N_20731,N_20774);
nor U24162 (N_24162,N_19242,N_20939);
nor U24163 (N_24163,N_20501,N_20977);
nand U24164 (N_24164,N_21817,N_21475);
nor U24165 (N_24165,N_20683,N_21516);
and U24166 (N_24166,N_19626,N_19396);
nor U24167 (N_24167,N_21250,N_20396);
xor U24168 (N_24168,N_21386,N_21644);
nand U24169 (N_24169,N_20581,N_20231);
and U24170 (N_24170,N_20056,N_21867);
and U24171 (N_24171,N_21282,N_21211);
or U24172 (N_24172,N_19311,N_20917);
xor U24173 (N_24173,N_21306,N_20102);
nor U24174 (N_24174,N_20402,N_19230);
or U24175 (N_24175,N_19881,N_20142);
xnor U24176 (N_24176,N_18892,N_21779);
and U24177 (N_24177,N_19093,N_21513);
and U24178 (N_24178,N_19755,N_21815);
nand U24179 (N_24179,N_19073,N_21038);
nor U24180 (N_24180,N_20102,N_19471);
xor U24181 (N_24181,N_20083,N_19630);
or U24182 (N_24182,N_21819,N_21780);
and U24183 (N_24183,N_19032,N_19994);
nand U24184 (N_24184,N_19007,N_19095);
and U24185 (N_24185,N_20173,N_21783);
nor U24186 (N_24186,N_21721,N_19012);
nand U24187 (N_24187,N_20620,N_19929);
and U24188 (N_24188,N_20909,N_20710);
xnor U24189 (N_24189,N_20051,N_21466);
or U24190 (N_24190,N_19415,N_19012);
nand U24191 (N_24191,N_20556,N_19821);
xor U24192 (N_24192,N_20912,N_21027);
and U24193 (N_24193,N_21570,N_20885);
nand U24194 (N_24194,N_20205,N_21306);
nor U24195 (N_24195,N_21680,N_20243);
nand U24196 (N_24196,N_21230,N_19524);
xnor U24197 (N_24197,N_19054,N_19515);
or U24198 (N_24198,N_20114,N_21810);
xnor U24199 (N_24199,N_19365,N_21794);
nand U24200 (N_24200,N_21298,N_21506);
nand U24201 (N_24201,N_19169,N_19223);
nor U24202 (N_24202,N_20037,N_19301);
nor U24203 (N_24203,N_19862,N_21009);
nor U24204 (N_24204,N_21469,N_20171);
xor U24205 (N_24205,N_19941,N_20094);
nor U24206 (N_24206,N_19922,N_21653);
nand U24207 (N_24207,N_19060,N_20883);
and U24208 (N_24208,N_21203,N_20090);
xor U24209 (N_24209,N_20436,N_21579);
xnor U24210 (N_24210,N_21242,N_20613);
and U24211 (N_24211,N_21446,N_19113);
or U24212 (N_24212,N_19758,N_19566);
xnor U24213 (N_24213,N_19403,N_19068);
nor U24214 (N_24214,N_18991,N_18960);
or U24215 (N_24215,N_21558,N_21447);
nor U24216 (N_24216,N_20860,N_20189);
nand U24217 (N_24217,N_19534,N_19148);
nor U24218 (N_24218,N_20035,N_19391);
xnor U24219 (N_24219,N_18832,N_19695);
and U24220 (N_24220,N_20540,N_19998);
xor U24221 (N_24221,N_20793,N_19100);
xor U24222 (N_24222,N_20528,N_20415);
and U24223 (N_24223,N_20874,N_19999);
xnor U24224 (N_24224,N_20539,N_18974);
and U24225 (N_24225,N_20836,N_19928);
nor U24226 (N_24226,N_20465,N_19745);
nor U24227 (N_24227,N_19186,N_21229);
nor U24228 (N_24228,N_20964,N_19702);
and U24229 (N_24229,N_20618,N_21660);
and U24230 (N_24230,N_21641,N_19913);
nor U24231 (N_24231,N_19103,N_19893);
or U24232 (N_24232,N_21104,N_21787);
and U24233 (N_24233,N_18934,N_20185);
xnor U24234 (N_24234,N_21316,N_21203);
nand U24235 (N_24235,N_21553,N_20286);
xor U24236 (N_24236,N_19247,N_20744);
and U24237 (N_24237,N_20591,N_19918);
nand U24238 (N_24238,N_21803,N_21367);
nand U24239 (N_24239,N_18796,N_20520);
nand U24240 (N_24240,N_20163,N_20991);
nand U24241 (N_24241,N_20894,N_20080);
and U24242 (N_24242,N_20495,N_21140);
xnor U24243 (N_24243,N_21597,N_19268);
xor U24244 (N_24244,N_19430,N_21736);
nor U24245 (N_24245,N_20116,N_18755);
nor U24246 (N_24246,N_19005,N_19998);
nand U24247 (N_24247,N_20042,N_19131);
nand U24248 (N_24248,N_20078,N_20029);
xnor U24249 (N_24249,N_20536,N_21670);
xnor U24250 (N_24250,N_19856,N_20291);
nor U24251 (N_24251,N_21779,N_21802);
nand U24252 (N_24252,N_19305,N_19207);
and U24253 (N_24253,N_21272,N_20334);
nor U24254 (N_24254,N_18833,N_21474);
and U24255 (N_24255,N_19365,N_19540);
xnor U24256 (N_24256,N_18826,N_19465);
nor U24257 (N_24257,N_19312,N_19662);
or U24258 (N_24258,N_19981,N_19214);
nor U24259 (N_24259,N_20046,N_21278);
nor U24260 (N_24260,N_19933,N_21533);
or U24261 (N_24261,N_19107,N_18831);
or U24262 (N_24262,N_19873,N_20771);
nand U24263 (N_24263,N_19085,N_20283);
xnor U24264 (N_24264,N_19437,N_19205);
nor U24265 (N_24265,N_21350,N_21221);
xnor U24266 (N_24266,N_20733,N_20832);
nand U24267 (N_24267,N_20282,N_18757);
and U24268 (N_24268,N_19953,N_19419);
xor U24269 (N_24269,N_20880,N_20574);
and U24270 (N_24270,N_19293,N_20217);
and U24271 (N_24271,N_19853,N_21226);
nor U24272 (N_24272,N_21528,N_21329);
xor U24273 (N_24273,N_20079,N_20568);
or U24274 (N_24274,N_21144,N_19764);
xor U24275 (N_24275,N_19821,N_19292);
nor U24276 (N_24276,N_21801,N_20405);
nand U24277 (N_24277,N_21234,N_19471);
and U24278 (N_24278,N_19102,N_19369);
and U24279 (N_24279,N_20636,N_20671);
and U24280 (N_24280,N_21740,N_19665);
nand U24281 (N_24281,N_18795,N_20113);
and U24282 (N_24282,N_19737,N_19271);
and U24283 (N_24283,N_21121,N_20118);
nand U24284 (N_24284,N_19303,N_20261);
nor U24285 (N_24285,N_20461,N_20983);
nand U24286 (N_24286,N_21863,N_21050);
or U24287 (N_24287,N_19057,N_19621);
nand U24288 (N_24288,N_19677,N_19064);
xnor U24289 (N_24289,N_21641,N_20735);
nor U24290 (N_24290,N_21561,N_21167);
xor U24291 (N_24291,N_20317,N_19395);
nand U24292 (N_24292,N_21618,N_19727);
nand U24293 (N_24293,N_19980,N_20967);
and U24294 (N_24294,N_20338,N_19505);
or U24295 (N_24295,N_21352,N_19303);
or U24296 (N_24296,N_19726,N_20270);
and U24297 (N_24297,N_21740,N_21632);
or U24298 (N_24298,N_19721,N_19348);
xnor U24299 (N_24299,N_21214,N_21053);
nor U24300 (N_24300,N_19456,N_21624);
or U24301 (N_24301,N_21033,N_21292);
nand U24302 (N_24302,N_20105,N_19882);
and U24303 (N_24303,N_21255,N_19950);
and U24304 (N_24304,N_21208,N_19252);
nand U24305 (N_24305,N_19653,N_21632);
and U24306 (N_24306,N_20967,N_21153);
or U24307 (N_24307,N_19337,N_19632);
nor U24308 (N_24308,N_20648,N_19282);
xor U24309 (N_24309,N_21524,N_20451);
xnor U24310 (N_24310,N_21649,N_21855);
nand U24311 (N_24311,N_20424,N_21575);
nand U24312 (N_24312,N_20118,N_19387);
xnor U24313 (N_24313,N_19920,N_19872);
nand U24314 (N_24314,N_21435,N_21307);
and U24315 (N_24315,N_20209,N_19195);
xnor U24316 (N_24316,N_21265,N_20512);
or U24317 (N_24317,N_20179,N_20585);
xor U24318 (N_24318,N_19220,N_19667);
or U24319 (N_24319,N_20406,N_20650);
xnor U24320 (N_24320,N_19390,N_20110);
nand U24321 (N_24321,N_19723,N_19545);
and U24322 (N_24322,N_19285,N_19609);
or U24323 (N_24323,N_21457,N_20048);
and U24324 (N_24324,N_21795,N_21333);
nand U24325 (N_24325,N_20325,N_20522);
nor U24326 (N_24326,N_21548,N_20570);
xor U24327 (N_24327,N_20973,N_20047);
or U24328 (N_24328,N_21635,N_20891);
nor U24329 (N_24329,N_18838,N_20317);
nand U24330 (N_24330,N_19503,N_21684);
nand U24331 (N_24331,N_19225,N_20502);
xor U24332 (N_24332,N_20597,N_20783);
nor U24333 (N_24333,N_21166,N_19151);
xor U24334 (N_24334,N_19084,N_19037);
and U24335 (N_24335,N_19533,N_20827);
and U24336 (N_24336,N_21219,N_19374);
or U24337 (N_24337,N_21744,N_21548);
xor U24338 (N_24338,N_19003,N_20617);
nand U24339 (N_24339,N_20872,N_20307);
xnor U24340 (N_24340,N_21468,N_21803);
nand U24341 (N_24341,N_19352,N_21162);
nand U24342 (N_24342,N_21621,N_18825);
nor U24343 (N_24343,N_19117,N_20128);
nand U24344 (N_24344,N_19582,N_20459);
xnor U24345 (N_24345,N_20939,N_19415);
nor U24346 (N_24346,N_21764,N_19769);
xor U24347 (N_24347,N_19175,N_20204);
xor U24348 (N_24348,N_18892,N_18899);
nor U24349 (N_24349,N_21307,N_21492);
nor U24350 (N_24350,N_19380,N_21624);
nor U24351 (N_24351,N_21522,N_19513);
and U24352 (N_24352,N_19769,N_20866);
and U24353 (N_24353,N_20862,N_18969);
or U24354 (N_24354,N_20969,N_21391);
xnor U24355 (N_24355,N_19577,N_19372);
and U24356 (N_24356,N_19755,N_21136);
and U24357 (N_24357,N_21503,N_19228);
nor U24358 (N_24358,N_21124,N_21145);
xor U24359 (N_24359,N_20312,N_20800);
nand U24360 (N_24360,N_18853,N_20160);
or U24361 (N_24361,N_20359,N_21088);
and U24362 (N_24362,N_19284,N_20576);
nand U24363 (N_24363,N_19180,N_21069);
or U24364 (N_24364,N_21029,N_21521);
xor U24365 (N_24365,N_20958,N_21051);
xnor U24366 (N_24366,N_19679,N_20855);
nand U24367 (N_24367,N_18781,N_19418);
nand U24368 (N_24368,N_21597,N_20713);
nor U24369 (N_24369,N_21464,N_19238);
nor U24370 (N_24370,N_19915,N_21232);
xnor U24371 (N_24371,N_19045,N_21638);
or U24372 (N_24372,N_20671,N_19240);
xnor U24373 (N_24373,N_19353,N_20393);
nand U24374 (N_24374,N_21447,N_20696);
or U24375 (N_24375,N_20281,N_19257);
nand U24376 (N_24376,N_20159,N_21757);
xor U24377 (N_24377,N_21619,N_20823);
or U24378 (N_24378,N_19321,N_19015);
xor U24379 (N_24379,N_19262,N_19783);
xor U24380 (N_24380,N_19748,N_19415);
or U24381 (N_24381,N_21608,N_20025);
and U24382 (N_24382,N_20968,N_18752);
or U24383 (N_24383,N_21628,N_21655);
xnor U24384 (N_24384,N_19151,N_20899);
nand U24385 (N_24385,N_20664,N_20558);
or U24386 (N_24386,N_21757,N_21284);
nor U24387 (N_24387,N_20167,N_20079);
xnor U24388 (N_24388,N_20392,N_20577);
xnor U24389 (N_24389,N_19118,N_21756);
nor U24390 (N_24390,N_19155,N_19254);
nand U24391 (N_24391,N_19245,N_19529);
xor U24392 (N_24392,N_21696,N_20710);
and U24393 (N_24393,N_19827,N_20839);
xor U24394 (N_24394,N_19498,N_18989);
nor U24395 (N_24395,N_21859,N_21025);
nor U24396 (N_24396,N_20154,N_21502);
or U24397 (N_24397,N_19039,N_19654);
nor U24398 (N_24398,N_21418,N_20022);
or U24399 (N_24399,N_21649,N_20665);
xor U24400 (N_24400,N_20935,N_19613);
or U24401 (N_24401,N_21483,N_19472);
nand U24402 (N_24402,N_20433,N_19737);
or U24403 (N_24403,N_20186,N_21836);
and U24404 (N_24404,N_18985,N_21636);
nand U24405 (N_24405,N_19047,N_20041);
nor U24406 (N_24406,N_20659,N_20611);
xor U24407 (N_24407,N_19305,N_20441);
nor U24408 (N_24408,N_20700,N_21238);
or U24409 (N_24409,N_20792,N_18886);
nor U24410 (N_24410,N_21665,N_19252);
xnor U24411 (N_24411,N_21041,N_21312);
nand U24412 (N_24412,N_21309,N_21662);
nor U24413 (N_24413,N_19052,N_21451);
nor U24414 (N_24414,N_19307,N_20743);
and U24415 (N_24415,N_19209,N_21736);
xnor U24416 (N_24416,N_21446,N_21661);
and U24417 (N_24417,N_21014,N_21499);
or U24418 (N_24418,N_20715,N_20420);
xor U24419 (N_24419,N_19150,N_21787);
or U24420 (N_24420,N_18910,N_21381);
and U24421 (N_24421,N_20829,N_20266);
xnor U24422 (N_24422,N_19720,N_18962);
nand U24423 (N_24423,N_21685,N_21415);
and U24424 (N_24424,N_19246,N_20206);
or U24425 (N_24425,N_19801,N_21296);
and U24426 (N_24426,N_19550,N_20204);
and U24427 (N_24427,N_20799,N_21002);
or U24428 (N_24428,N_21308,N_21795);
and U24429 (N_24429,N_20046,N_19240);
nand U24430 (N_24430,N_20516,N_21579);
nand U24431 (N_24431,N_21691,N_18849);
xnor U24432 (N_24432,N_19671,N_20869);
and U24433 (N_24433,N_20840,N_21636);
nor U24434 (N_24434,N_20088,N_20606);
xnor U24435 (N_24435,N_21266,N_19417);
and U24436 (N_24436,N_20992,N_21480);
xor U24437 (N_24437,N_19861,N_18885);
and U24438 (N_24438,N_19343,N_18785);
xor U24439 (N_24439,N_18841,N_19125);
nand U24440 (N_24440,N_18947,N_21410);
or U24441 (N_24441,N_21374,N_21157);
and U24442 (N_24442,N_18938,N_20145);
nand U24443 (N_24443,N_19709,N_20266);
nand U24444 (N_24444,N_21745,N_20260);
nor U24445 (N_24445,N_20686,N_19188);
or U24446 (N_24446,N_20850,N_21585);
nand U24447 (N_24447,N_19584,N_20631);
nand U24448 (N_24448,N_19561,N_21569);
xnor U24449 (N_24449,N_21862,N_19400);
xnor U24450 (N_24450,N_18865,N_21076);
nor U24451 (N_24451,N_20943,N_19390);
nand U24452 (N_24452,N_21655,N_21436);
and U24453 (N_24453,N_20499,N_21767);
or U24454 (N_24454,N_19286,N_20911);
and U24455 (N_24455,N_20742,N_20090);
nor U24456 (N_24456,N_19870,N_19942);
and U24457 (N_24457,N_20064,N_18984);
xor U24458 (N_24458,N_19374,N_20045);
and U24459 (N_24459,N_21220,N_20549);
nand U24460 (N_24460,N_19462,N_20432);
xnor U24461 (N_24461,N_19178,N_19609);
and U24462 (N_24462,N_20649,N_19287);
xor U24463 (N_24463,N_21132,N_21396);
xor U24464 (N_24464,N_19905,N_20302);
xor U24465 (N_24465,N_20704,N_20916);
nand U24466 (N_24466,N_19721,N_19603);
nand U24467 (N_24467,N_20346,N_18995);
or U24468 (N_24468,N_19775,N_18760);
xnor U24469 (N_24469,N_21841,N_19930);
xnor U24470 (N_24470,N_21653,N_20392);
and U24471 (N_24471,N_19891,N_21309);
nor U24472 (N_24472,N_18907,N_19413);
nor U24473 (N_24473,N_21318,N_21496);
or U24474 (N_24474,N_21400,N_21351);
and U24475 (N_24475,N_19365,N_19091);
nor U24476 (N_24476,N_20158,N_20501);
nor U24477 (N_24477,N_21729,N_21789);
nor U24478 (N_24478,N_20240,N_20552);
nand U24479 (N_24479,N_21004,N_19619);
xor U24480 (N_24480,N_21193,N_19946);
nand U24481 (N_24481,N_21213,N_20061);
nand U24482 (N_24482,N_20268,N_20113);
and U24483 (N_24483,N_20276,N_20245);
or U24484 (N_24484,N_19848,N_19450);
xnor U24485 (N_24485,N_19565,N_21726);
and U24486 (N_24486,N_19639,N_20666);
and U24487 (N_24487,N_21725,N_20120);
nor U24488 (N_24488,N_19181,N_21528);
nor U24489 (N_24489,N_18824,N_19447);
nor U24490 (N_24490,N_19253,N_19908);
xor U24491 (N_24491,N_21409,N_20290);
xnor U24492 (N_24492,N_19828,N_20742);
nand U24493 (N_24493,N_20725,N_19608);
or U24494 (N_24494,N_21292,N_19071);
nor U24495 (N_24495,N_20072,N_18939);
nor U24496 (N_24496,N_19937,N_18970);
nor U24497 (N_24497,N_19441,N_19638);
or U24498 (N_24498,N_18861,N_20569);
xor U24499 (N_24499,N_19529,N_20773);
or U24500 (N_24500,N_19944,N_21804);
and U24501 (N_24501,N_20045,N_19056);
nand U24502 (N_24502,N_20095,N_19408);
nand U24503 (N_24503,N_19291,N_19214);
or U24504 (N_24504,N_19608,N_20888);
xor U24505 (N_24505,N_21033,N_20643);
and U24506 (N_24506,N_20133,N_20393);
or U24507 (N_24507,N_20109,N_20229);
and U24508 (N_24508,N_19767,N_21687);
or U24509 (N_24509,N_21011,N_19627);
or U24510 (N_24510,N_18793,N_18937);
or U24511 (N_24511,N_21664,N_19633);
nor U24512 (N_24512,N_19840,N_19901);
nand U24513 (N_24513,N_20950,N_18948);
and U24514 (N_24514,N_19694,N_18829);
xor U24515 (N_24515,N_20630,N_21705);
nand U24516 (N_24516,N_18923,N_19504);
and U24517 (N_24517,N_21344,N_19255);
nand U24518 (N_24518,N_20225,N_19404);
nand U24519 (N_24519,N_19042,N_20209);
xnor U24520 (N_24520,N_19858,N_21094);
or U24521 (N_24521,N_19090,N_21313);
nand U24522 (N_24522,N_19926,N_19515);
nor U24523 (N_24523,N_21653,N_19212);
nand U24524 (N_24524,N_19487,N_18960);
nor U24525 (N_24525,N_20921,N_21250);
xor U24526 (N_24526,N_19901,N_19645);
or U24527 (N_24527,N_19971,N_20345);
or U24528 (N_24528,N_18802,N_21161);
xnor U24529 (N_24529,N_21716,N_19540);
nand U24530 (N_24530,N_21025,N_19254);
xor U24531 (N_24531,N_21753,N_19482);
and U24532 (N_24532,N_21127,N_20971);
or U24533 (N_24533,N_20824,N_21758);
xnor U24534 (N_24534,N_21331,N_19166);
and U24535 (N_24535,N_18929,N_20075);
and U24536 (N_24536,N_20444,N_19109);
or U24537 (N_24537,N_18825,N_19511);
or U24538 (N_24538,N_19305,N_20527);
and U24539 (N_24539,N_21401,N_19818);
xor U24540 (N_24540,N_21775,N_21302);
and U24541 (N_24541,N_21410,N_21484);
or U24542 (N_24542,N_19013,N_19283);
and U24543 (N_24543,N_21695,N_19167);
xnor U24544 (N_24544,N_19486,N_21608);
xnor U24545 (N_24545,N_21381,N_18911);
nand U24546 (N_24546,N_19812,N_20999);
or U24547 (N_24547,N_18818,N_19675);
or U24548 (N_24548,N_20464,N_19837);
xor U24549 (N_24549,N_20771,N_21426);
nor U24550 (N_24550,N_19787,N_20007);
or U24551 (N_24551,N_19712,N_18807);
and U24552 (N_24552,N_20230,N_19042);
or U24553 (N_24553,N_19853,N_20064);
nor U24554 (N_24554,N_20297,N_19044);
nor U24555 (N_24555,N_20693,N_19948);
nor U24556 (N_24556,N_18791,N_19606);
nor U24557 (N_24557,N_20135,N_21670);
nor U24558 (N_24558,N_21591,N_19735);
xor U24559 (N_24559,N_21209,N_20793);
xor U24560 (N_24560,N_21034,N_21437);
xor U24561 (N_24561,N_21624,N_19413);
or U24562 (N_24562,N_18824,N_20167);
or U24563 (N_24563,N_18815,N_21543);
or U24564 (N_24564,N_21162,N_20939);
nor U24565 (N_24565,N_19620,N_20133);
or U24566 (N_24566,N_19000,N_20800);
xor U24567 (N_24567,N_19441,N_19199);
nor U24568 (N_24568,N_19648,N_20585);
xnor U24569 (N_24569,N_19223,N_20476);
and U24570 (N_24570,N_20702,N_21160);
and U24571 (N_24571,N_21726,N_21760);
nand U24572 (N_24572,N_21358,N_18767);
and U24573 (N_24573,N_21555,N_19598);
nor U24574 (N_24574,N_19671,N_19081);
nor U24575 (N_24575,N_18777,N_19576);
and U24576 (N_24576,N_21587,N_19585);
xor U24577 (N_24577,N_20044,N_20684);
xor U24578 (N_24578,N_20581,N_20458);
nor U24579 (N_24579,N_19966,N_21058);
nand U24580 (N_24580,N_19895,N_21124);
and U24581 (N_24581,N_21041,N_19884);
xor U24582 (N_24582,N_19534,N_20596);
xnor U24583 (N_24583,N_20011,N_21166);
nand U24584 (N_24584,N_19138,N_21216);
or U24585 (N_24585,N_21827,N_21680);
nand U24586 (N_24586,N_20205,N_20833);
and U24587 (N_24587,N_20587,N_21210);
or U24588 (N_24588,N_20999,N_19041);
xor U24589 (N_24589,N_20585,N_21525);
xnor U24590 (N_24590,N_19484,N_19287);
nor U24591 (N_24591,N_21317,N_21318);
xnor U24592 (N_24592,N_19233,N_21753);
or U24593 (N_24593,N_21734,N_21653);
nand U24594 (N_24594,N_20293,N_21063);
or U24595 (N_24595,N_20009,N_21229);
xnor U24596 (N_24596,N_19798,N_19176);
xor U24597 (N_24597,N_21109,N_18812);
nor U24598 (N_24598,N_21747,N_20664);
nand U24599 (N_24599,N_19436,N_19744);
xor U24600 (N_24600,N_21048,N_18949);
nor U24601 (N_24601,N_21674,N_21660);
or U24602 (N_24602,N_20567,N_19137);
nand U24603 (N_24603,N_19414,N_20289);
and U24604 (N_24604,N_21553,N_20700);
nand U24605 (N_24605,N_19271,N_19633);
and U24606 (N_24606,N_21696,N_21586);
xnor U24607 (N_24607,N_19856,N_19973);
nand U24608 (N_24608,N_20789,N_20967);
and U24609 (N_24609,N_19884,N_21307);
nor U24610 (N_24610,N_20515,N_20182);
and U24611 (N_24611,N_21187,N_19533);
nand U24612 (N_24612,N_21023,N_20268);
nand U24613 (N_24613,N_20814,N_20031);
nor U24614 (N_24614,N_20106,N_21203);
nor U24615 (N_24615,N_19733,N_18911);
nand U24616 (N_24616,N_21313,N_18970);
nor U24617 (N_24617,N_20583,N_20308);
xnor U24618 (N_24618,N_21286,N_19038);
and U24619 (N_24619,N_20249,N_19593);
or U24620 (N_24620,N_19196,N_19238);
or U24621 (N_24621,N_19237,N_21333);
xnor U24622 (N_24622,N_20038,N_21391);
nor U24623 (N_24623,N_19626,N_21334);
xnor U24624 (N_24624,N_21211,N_19708);
and U24625 (N_24625,N_19740,N_20351);
nor U24626 (N_24626,N_19309,N_21739);
nand U24627 (N_24627,N_20566,N_20057);
nand U24628 (N_24628,N_20384,N_20130);
nor U24629 (N_24629,N_20770,N_21352);
and U24630 (N_24630,N_21505,N_19897);
nand U24631 (N_24631,N_18920,N_20109);
nor U24632 (N_24632,N_21649,N_18754);
and U24633 (N_24633,N_21393,N_20788);
nor U24634 (N_24634,N_18795,N_21212);
xnor U24635 (N_24635,N_21312,N_19779);
nand U24636 (N_24636,N_19431,N_20143);
and U24637 (N_24637,N_18867,N_18900);
xnor U24638 (N_24638,N_21475,N_19602);
xnor U24639 (N_24639,N_20585,N_19084);
or U24640 (N_24640,N_21416,N_19602);
nor U24641 (N_24641,N_19752,N_21388);
nand U24642 (N_24642,N_19354,N_19809);
nor U24643 (N_24643,N_21844,N_19131);
and U24644 (N_24644,N_19988,N_21214);
nor U24645 (N_24645,N_21146,N_19701);
nor U24646 (N_24646,N_20816,N_20108);
or U24647 (N_24647,N_19351,N_20567);
nand U24648 (N_24648,N_19326,N_20053);
or U24649 (N_24649,N_21638,N_21464);
xor U24650 (N_24650,N_20761,N_20030);
or U24651 (N_24651,N_19098,N_20446);
and U24652 (N_24652,N_18847,N_19222);
or U24653 (N_24653,N_21480,N_20591);
or U24654 (N_24654,N_20986,N_21264);
nand U24655 (N_24655,N_19101,N_20080);
xor U24656 (N_24656,N_19439,N_20597);
or U24657 (N_24657,N_19967,N_21163);
nor U24658 (N_24658,N_19703,N_21706);
nand U24659 (N_24659,N_19324,N_19224);
nand U24660 (N_24660,N_19289,N_20264);
xor U24661 (N_24661,N_21828,N_20494);
nor U24662 (N_24662,N_19253,N_19378);
nand U24663 (N_24663,N_21400,N_19046);
xnor U24664 (N_24664,N_20239,N_19433);
nor U24665 (N_24665,N_21068,N_18767);
and U24666 (N_24666,N_21019,N_21869);
nand U24667 (N_24667,N_19896,N_19425);
or U24668 (N_24668,N_20252,N_20086);
or U24669 (N_24669,N_21865,N_19351);
nor U24670 (N_24670,N_21111,N_20704);
nand U24671 (N_24671,N_18949,N_19193);
and U24672 (N_24672,N_20776,N_21690);
nand U24673 (N_24673,N_20500,N_19225);
and U24674 (N_24674,N_21133,N_20287);
xor U24675 (N_24675,N_21037,N_18798);
xnor U24676 (N_24676,N_20979,N_18905);
or U24677 (N_24677,N_18820,N_20105);
or U24678 (N_24678,N_18851,N_20451);
xnor U24679 (N_24679,N_20562,N_19737);
or U24680 (N_24680,N_19477,N_20943);
or U24681 (N_24681,N_20916,N_21493);
and U24682 (N_24682,N_18758,N_18940);
nand U24683 (N_24683,N_18892,N_20042);
or U24684 (N_24684,N_18818,N_20545);
and U24685 (N_24685,N_21273,N_21558);
xnor U24686 (N_24686,N_20513,N_20869);
and U24687 (N_24687,N_21842,N_21601);
xor U24688 (N_24688,N_18848,N_19695);
and U24689 (N_24689,N_21573,N_19485);
xor U24690 (N_24690,N_19139,N_19974);
and U24691 (N_24691,N_21488,N_20403);
and U24692 (N_24692,N_19754,N_19026);
and U24693 (N_24693,N_20963,N_21519);
and U24694 (N_24694,N_21302,N_20103);
and U24695 (N_24695,N_19016,N_20283);
nand U24696 (N_24696,N_21552,N_20370);
or U24697 (N_24697,N_21791,N_20821);
and U24698 (N_24698,N_20569,N_19420);
nor U24699 (N_24699,N_18980,N_20177);
and U24700 (N_24700,N_19274,N_21724);
xor U24701 (N_24701,N_19198,N_19728);
nor U24702 (N_24702,N_19313,N_20564);
or U24703 (N_24703,N_21004,N_20347);
nor U24704 (N_24704,N_21363,N_21242);
and U24705 (N_24705,N_18889,N_20707);
xnor U24706 (N_24706,N_19562,N_19499);
nand U24707 (N_24707,N_19082,N_20246);
and U24708 (N_24708,N_18886,N_20721);
nor U24709 (N_24709,N_21476,N_21386);
xor U24710 (N_24710,N_18840,N_20889);
xnor U24711 (N_24711,N_20376,N_20903);
and U24712 (N_24712,N_20646,N_19727);
xnor U24713 (N_24713,N_19622,N_19191);
nand U24714 (N_24714,N_21386,N_21706);
xnor U24715 (N_24715,N_20036,N_20229);
xor U24716 (N_24716,N_18829,N_20120);
nand U24717 (N_24717,N_20139,N_19968);
and U24718 (N_24718,N_20574,N_20206);
or U24719 (N_24719,N_20529,N_20160);
xnor U24720 (N_24720,N_20404,N_20145);
or U24721 (N_24721,N_19622,N_20695);
or U24722 (N_24722,N_20636,N_19887);
xnor U24723 (N_24723,N_19013,N_21132);
xor U24724 (N_24724,N_21784,N_18929);
or U24725 (N_24725,N_19087,N_20041);
and U24726 (N_24726,N_20818,N_20221);
nor U24727 (N_24727,N_21662,N_20226);
or U24728 (N_24728,N_18964,N_19939);
nand U24729 (N_24729,N_20001,N_20243);
nand U24730 (N_24730,N_20846,N_21205);
xor U24731 (N_24731,N_20009,N_21475);
xnor U24732 (N_24732,N_19766,N_20424);
xnor U24733 (N_24733,N_19863,N_18818);
or U24734 (N_24734,N_21083,N_19756);
or U24735 (N_24735,N_21135,N_18876);
nand U24736 (N_24736,N_21595,N_21146);
and U24737 (N_24737,N_19571,N_19271);
nor U24738 (N_24738,N_21048,N_20151);
xnor U24739 (N_24739,N_20396,N_19461);
nand U24740 (N_24740,N_21122,N_19015);
xor U24741 (N_24741,N_19920,N_19292);
nand U24742 (N_24742,N_19090,N_19577);
nor U24743 (N_24743,N_20030,N_21398);
nand U24744 (N_24744,N_20341,N_21125);
or U24745 (N_24745,N_20954,N_21523);
or U24746 (N_24746,N_20512,N_19713);
nand U24747 (N_24747,N_20237,N_20378);
or U24748 (N_24748,N_21213,N_21753);
nor U24749 (N_24749,N_19527,N_20904);
nor U24750 (N_24750,N_20497,N_20852);
nor U24751 (N_24751,N_18812,N_19418);
nor U24752 (N_24752,N_20913,N_19386);
nand U24753 (N_24753,N_20659,N_20756);
and U24754 (N_24754,N_20467,N_20523);
nand U24755 (N_24755,N_20217,N_19142);
and U24756 (N_24756,N_21459,N_21654);
and U24757 (N_24757,N_19893,N_19932);
nand U24758 (N_24758,N_20646,N_19198);
xnor U24759 (N_24759,N_19987,N_19793);
or U24760 (N_24760,N_20036,N_21705);
nand U24761 (N_24761,N_19634,N_21803);
nand U24762 (N_24762,N_21015,N_19830);
xnor U24763 (N_24763,N_19820,N_19344);
or U24764 (N_24764,N_21361,N_19106);
and U24765 (N_24765,N_18899,N_19646);
and U24766 (N_24766,N_19362,N_19034);
and U24767 (N_24767,N_19218,N_20236);
nand U24768 (N_24768,N_20812,N_19238);
or U24769 (N_24769,N_21616,N_19641);
nand U24770 (N_24770,N_19231,N_21582);
nand U24771 (N_24771,N_21835,N_20481);
or U24772 (N_24772,N_20798,N_20692);
xnor U24773 (N_24773,N_19136,N_21407);
or U24774 (N_24774,N_20170,N_18889);
and U24775 (N_24775,N_21264,N_19928);
xor U24776 (N_24776,N_20357,N_21402);
nor U24777 (N_24777,N_21099,N_20652);
nand U24778 (N_24778,N_19080,N_19149);
or U24779 (N_24779,N_19187,N_19025);
xor U24780 (N_24780,N_21162,N_21197);
nand U24781 (N_24781,N_20218,N_20923);
nand U24782 (N_24782,N_20520,N_20340);
nor U24783 (N_24783,N_21692,N_21529);
and U24784 (N_24784,N_19895,N_20247);
or U24785 (N_24785,N_20726,N_19449);
or U24786 (N_24786,N_19889,N_19863);
xor U24787 (N_24787,N_19025,N_19882);
or U24788 (N_24788,N_19153,N_21248);
nand U24789 (N_24789,N_21645,N_19582);
xnor U24790 (N_24790,N_20260,N_18829);
xor U24791 (N_24791,N_21825,N_21717);
nor U24792 (N_24792,N_19497,N_19805);
xnor U24793 (N_24793,N_21743,N_20849);
xor U24794 (N_24794,N_19787,N_20824);
nor U24795 (N_24795,N_18803,N_18892);
xor U24796 (N_24796,N_21500,N_19241);
or U24797 (N_24797,N_21613,N_21804);
nand U24798 (N_24798,N_20328,N_20419);
and U24799 (N_24799,N_20388,N_21148);
or U24800 (N_24800,N_20313,N_20098);
nand U24801 (N_24801,N_19183,N_20507);
nor U24802 (N_24802,N_20118,N_21690);
xnor U24803 (N_24803,N_19695,N_20899);
or U24804 (N_24804,N_20864,N_21378);
nand U24805 (N_24805,N_19742,N_18948);
and U24806 (N_24806,N_18752,N_19610);
xnor U24807 (N_24807,N_20610,N_19690);
nand U24808 (N_24808,N_19902,N_21091);
nand U24809 (N_24809,N_19661,N_20733);
or U24810 (N_24810,N_18902,N_18875);
nand U24811 (N_24811,N_20929,N_18844);
nor U24812 (N_24812,N_21351,N_18937);
nand U24813 (N_24813,N_19720,N_20808);
xnor U24814 (N_24814,N_21430,N_19287);
and U24815 (N_24815,N_21162,N_20631);
xor U24816 (N_24816,N_18877,N_21560);
xor U24817 (N_24817,N_18907,N_21251);
nand U24818 (N_24818,N_19326,N_20766);
xnor U24819 (N_24819,N_18954,N_19710);
nand U24820 (N_24820,N_19156,N_20250);
nand U24821 (N_24821,N_21815,N_20462);
xnor U24822 (N_24822,N_21465,N_21105);
nand U24823 (N_24823,N_21872,N_21768);
nor U24824 (N_24824,N_21019,N_20634);
nand U24825 (N_24825,N_19750,N_18853);
nand U24826 (N_24826,N_21240,N_20546);
nor U24827 (N_24827,N_21153,N_21370);
xor U24828 (N_24828,N_21528,N_20928);
nor U24829 (N_24829,N_18909,N_21247);
xnor U24830 (N_24830,N_19910,N_21040);
or U24831 (N_24831,N_21046,N_19286);
and U24832 (N_24832,N_20124,N_20291);
nor U24833 (N_24833,N_21105,N_20762);
xor U24834 (N_24834,N_20952,N_20498);
or U24835 (N_24835,N_21519,N_19637);
nor U24836 (N_24836,N_20511,N_21321);
and U24837 (N_24837,N_19403,N_20682);
nor U24838 (N_24838,N_20510,N_21588);
nor U24839 (N_24839,N_19490,N_19462);
and U24840 (N_24840,N_20593,N_20218);
and U24841 (N_24841,N_21623,N_19431);
nand U24842 (N_24842,N_19416,N_19078);
and U24843 (N_24843,N_20609,N_20251);
or U24844 (N_24844,N_20922,N_21860);
nand U24845 (N_24845,N_21427,N_18788);
nand U24846 (N_24846,N_21080,N_20777);
nor U24847 (N_24847,N_20406,N_19174);
nor U24848 (N_24848,N_20880,N_20577);
xnor U24849 (N_24849,N_20128,N_19427);
and U24850 (N_24850,N_20792,N_18984);
nor U24851 (N_24851,N_20494,N_21369);
nor U24852 (N_24852,N_21091,N_20130);
or U24853 (N_24853,N_19935,N_19641);
and U24854 (N_24854,N_20430,N_21619);
nand U24855 (N_24855,N_18842,N_19013);
or U24856 (N_24856,N_21602,N_20585);
or U24857 (N_24857,N_19611,N_21505);
or U24858 (N_24858,N_21658,N_20661);
nor U24859 (N_24859,N_20393,N_21210);
or U24860 (N_24860,N_19376,N_21638);
and U24861 (N_24861,N_21849,N_21503);
and U24862 (N_24862,N_19446,N_19568);
and U24863 (N_24863,N_19288,N_21330);
nor U24864 (N_24864,N_21040,N_19807);
and U24865 (N_24865,N_19061,N_19953);
xnor U24866 (N_24866,N_20634,N_20791);
nor U24867 (N_24867,N_18820,N_21591);
and U24868 (N_24868,N_21363,N_19867);
nand U24869 (N_24869,N_19082,N_21871);
nor U24870 (N_24870,N_19515,N_18821);
xor U24871 (N_24871,N_20246,N_21443);
or U24872 (N_24872,N_20637,N_19788);
nand U24873 (N_24873,N_18876,N_20729);
nor U24874 (N_24874,N_21509,N_18938);
nor U24875 (N_24875,N_19459,N_19520);
nand U24876 (N_24876,N_18999,N_21588);
xor U24877 (N_24877,N_19979,N_19503);
xnor U24878 (N_24878,N_19086,N_21649);
or U24879 (N_24879,N_20079,N_20413);
and U24880 (N_24880,N_21189,N_21183);
or U24881 (N_24881,N_20163,N_18831);
nor U24882 (N_24882,N_19476,N_20660);
nand U24883 (N_24883,N_20858,N_19993);
xnor U24884 (N_24884,N_20464,N_19231);
or U24885 (N_24885,N_20753,N_19998);
nand U24886 (N_24886,N_21343,N_20460);
nor U24887 (N_24887,N_19004,N_20909);
or U24888 (N_24888,N_20413,N_19933);
and U24889 (N_24889,N_19928,N_20259);
or U24890 (N_24890,N_19911,N_19587);
and U24891 (N_24891,N_21191,N_21059);
or U24892 (N_24892,N_20299,N_19332);
and U24893 (N_24893,N_19691,N_18980);
xnor U24894 (N_24894,N_21803,N_18786);
nand U24895 (N_24895,N_20460,N_19028);
xnor U24896 (N_24896,N_21209,N_20521);
or U24897 (N_24897,N_20192,N_21802);
nand U24898 (N_24898,N_20840,N_20148);
nand U24899 (N_24899,N_19597,N_21668);
nor U24900 (N_24900,N_20033,N_19772);
nand U24901 (N_24901,N_20826,N_20809);
or U24902 (N_24902,N_19872,N_21774);
xor U24903 (N_24903,N_21282,N_20569);
and U24904 (N_24904,N_21007,N_19204);
or U24905 (N_24905,N_20538,N_19198);
and U24906 (N_24906,N_21842,N_19229);
and U24907 (N_24907,N_21569,N_19572);
xor U24908 (N_24908,N_19174,N_21432);
and U24909 (N_24909,N_19448,N_19740);
nor U24910 (N_24910,N_21106,N_20533);
or U24911 (N_24911,N_21260,N_21341);
and U24912 (N_24912,N_20366,N_21108);
nand U24913 (N_24913,N_19055,N_21692);
nor U24914 (N_24914,N_19794,N_20963);
and U24915 (N_24915,N_19575,N_18828);
and U24916 (N_24916,N_20020,N_18845);
and U24917 (N_24917,N_18938,N_21730);
and U24918 (N_24918,N_21573,N_21657);
nand U24919 (N_24919,N_20640,N_20956);
nor U24920 (N_24920,N_18902,N_21532);
nor U24921 (N_24921,N_20839,N_21311);
nand U24922 (N_24922,N_18882,N_19531);
and U24923 (N_24923,N_19463,N_20913);
or U24924 (N_24924,N_21413,N_21313);
or U24925 (N_24925,N_21774,N_21555);
nand U24926 (N_24926,N_19141,N_20948);
nand U24927 (N_24927,N_20365,N_19440);
and U24928 (N_24928,N_21690,N_19608);
nand U24929 (N_24929,N_21867,N_19040);
xor U24930 (N_24930,N_18767,N_19292);
nand U24931 (N_24931,N_20674,N_20291);
nor U24932 (N_24932,N_19779,N_19873);
or U24933 (N_24933,N_21072,N_19845);
xor U24934 (N_24934,N_20341,N_19504);
and U24935 (N_24935,N_18795,N_21413);
or U24936 (N_24936,N_20438,N_19208);
nor U24937 (N_24937,N_21308,N_19001);
and U24938 (N_24938,N_21810,N_19985);
and U24939 (N_24939,N_20340,N_20539);
xor U24940 (N_24940,N_21701,N_21690);
and U24941 (N_24941,N_21422,N_21129);
nor U24942 (N_24942,N_19998,N_19900);
or U24943 (N_24943,N_19336,N_19275);
and U24944 (N_24944,N_19228,N_21816);
nand U24945 (N_24945,N_19308,N_20498);
xor U24946 (N_24946,N_21280,N_19448);
nor U24947 (N_24947,N_20126,N_19255);
xnor U24948 (N_24948,N_19168,N_21585);
nand U24949 (N_24949,N_21736,N_19690);
xnor U24950 (N_24950,N_20924,N_18822);
and U24951 (N_24951,N_21255,N_19860);
nand U24952 (N_24952,N_20390,N_21775);
xnor U24953 (N_24953,N_19921,N_20778);
nand U24954 (N_24954,N_20085,N_20806);
nand U24955 (N_24955,N_20236,N_21029);
xnor U24956 (N_24956,N_21044,N_21206);
and U24957 (N_24957,N_20148,N_20922);
nand U24958 (N_24958,N_20051,N_20694);
and U24959 (N_24959,N_19705,N_20424);
and U24960 (N_24960,N_20737,N_20998);
nor U24961 (N_24961,N_20435,N_21772);
and U24962 (N_24962,N_20430,N_19711);
or U24963 (N_24963,N_20975,N_21496);
nor U24964 (N_24964,N_20913,N_19240);
nand U24965 (N_24965,N_20016,N_20098);
and U24966 (N_24966,N_19637,N_20270);
xor U24967 (N_24967,N_21156,N_20972);
xnor U24968 (N_24968,N_19395,N_21806);
xor U24969 (N_24969,N_20341,N_19371);
nor U24970 (N_24970,N_19195,N_21153);
and U24971 (N_24971,N_21433,N_19210);
xor U24972 (N_24972,N_20808,N_19687);
nand U24973 (N_24973,N_21359,N_21719);
xor U24974 (N_24974,N_20171,N_19493);
xor U24975 (N_24975,N_19835,N_19747);
or U24976 (N_24976,N_20462,N_19421);
xnor U24977 (N_24977,N_21409,N_20635);
nor U24978 (N_24978,N_19254,N_20598);
and U24979 (N_24979,N_20476,N_20094);
xor U24980 (N_24980,N_21250,N_20492);
nand U24981 (N_24981,N_20632,N_20657);
nand U24982 (N_24982,N_20630,N_18983);
xor U24983 (N_24983,N_20165,N_21509);
or U24984 (N_24984,N_21487,N_21547);
and U24985 (N_24985,N_21793,N_20553);
or U24986 (N_24986,N_21713,N_20500);
or U24987 (N_24987,N_18967,N_20654);
nor U24988 (N_24988,N_20346,N_19187);
nand U24989 (N_24989,N_21758,N_19225);
or U24990 (N_24990,N_20513,N_18920);
or U24991 (N_24991,N_20303,N_21118);
xor U24992 (N_24992,N_18828,N_20526);
or U24993 (N_24993,N_20976,N_21695);
nand U24994 (N_24994,N_20770,N_20726);
and U24995 (N_24995,N_19657,N_21622);
or U24996 (N_24996,N_21411,N_20840);
nor U24997 (N_24997,N_19048,N_19544);
and U24998 (N_24998,N_21085,N_18857);
and U24999 (N_24999,N_19279,N_19959);
nor UO_0 (O_0,N_24491,N_23142);
nor UO_1 (O_1,N_24570,N_24766);
and UO_2 (O_2,N_23523,N_23086);
nor UO_3 (O_3,N_22762,N_23739);
nand UO_4 (O_4,N_24911,N_22459);
nand UO_5 (O_5,N_23177,N_24732);
or UO_6 (O_6,N_23561,N_24846);
nand UO_7 (O_7,N_23840,N_22768);
nand UO_8 (O_8,N_22991,N_22485);
nor UO_9 (O_9,N_22740,N_22515);
nand UO_10 (O_10,N_23853,N_23750);
and UO_11 (O_11,N_23205,N_24862);
nor UO_12 (O_12,N_24482,N_24559);
nor UO_13 (O_13,N_23902,N_24990);
nor UO_14 (O_14,N_24428,N_22390);
or UO_15 (O_15,N_24906,N_22670);
and UO_16 (O_16,N_24918,N_22508);
nand UO_17 (O_17,N_24313,N_23114);
nor UO_18 (O_18,N_22552,N_22081);
nor UO_19 (O_19,N_22152,N_24940);
or UO_20 (O_20,N_23039,N_24885);
nor UO_21 (O_21,N_24043,N_23600);
or UO_22 (O_22,N_22989,N_24873);
and UO_23 (O_23,N_23071,N_24996);
nand UO_24 (O_24,N_22141,N_22641);
nand UO_25 (O_25,N_23217,N_22329);
or UO_26 (O_26,N_22440,N_22422);
nor UO_27 (O_27,N_22662,N_24760);
nand UO_28 (O_28,N_23480,N_23216);
nand UO_29 (O_29,N_23966,N_22283);
xor UO_30 (O_30,N_24577,N_24196);
or UO_31 (O_31,N_23721,N_22623);
and UO_32 (O_32,N_22604,N_23028);
nor UO_33 (O_33,N_22476,N_22841);
xor UO_34 (O_34,N_22010,N_24876);
nand UO_35 (O_35,N_23378,N_24381);
xnor UO_36 (O_36,N_23295,N_24411);
nand UO_37 (O_37,N_22316,N_23711);
nor UO_38 (O_38,N_22062,N_23192);
and UO_39 (O_39,N_24441,N_24377);
or UO_40 (O_40,N_23947,N_23283);
and UO_41 (O_41,N_23377,N_23124);
nand UO_42 (O_42,N_23808,N_22253);
xnor UO_43 (O_43,N_24623,N_22842);
and UO_44 (O_44,N_23858,N_23695);
xnor UO_45 (O_45,N_24480,N_21888);
nor UO_46 (O_46,N_24517,N_24655);
and UO_47 (O_47,N_23030,N_21965);
and UO_48 (O_48,N_23131,N_23168);
and UO_49 (O_49,N_23343,N_22792);
and UO_50 (O_50,N_21886,N_22022);
nand UO_51 (O_51,N_24922,N_24342);
nor UO_52 (O_52,N_24265,N_22228);
xor UO_53 (O_53,N_22057,N_23149);
nor UO_54 (O_54,N_23341,N_23747);
xnor UO_55 (O_55,N_24405,N_22521);
nand UO_56 (O_56,N_24890,N_24057);
nor UO_57 (O_57,N_23171,N_24460);
nor UO_58 (O_58,N_24466,N_23802);
or UO_59 (O_59,N_24781,N_24206);
and UO_60 (O_60,N_22448,N_24029);
nor UO_61 (O_61,N_22318,N_22424);
and UO_62 (O_62,N_24030,N_23250);
nor UO_63 (O_63,N_21896,N_22950);
xor UO_64 (O_64,N_23745,N_24912);
or UO_65 (O_65,N_22649,N_24534);
nand UO_66 (O_66,N_23350,N_21955);
nand UO_67 (O_67,N_23683,N_22943);
or UO_68 (O_68,N_22277,N_23874);
and UO_69 (O_69,N_22583,N_24711);
or UO_70 (O_70,N_22666,N_23932);
nor UO_71 (O_71,N_24896,N_24737);
xor UO_72 (O_72,N_22749,N_22375);
or UO_73 (O_73,N_22890,N_24223);
and UO_74 (O_74,N_22857,N_24414);
xor UO_75 (O_75,N_24382,N_22076);
xor UO_76 (O_76,N_23896,N_24510);
nand UO_77 (O_77,N_24800,N_21884);
nand UO_78 (O_78,N_24602,N_22882);
and UO_79 (O_79,N_23676,N_22392);
nor UO_80 (O_80,N_24696,N_23460);
nor UO_81 (O_81,N_23094,N_22452);
nand UO_82 (O_82,N_22195,N_24391);
and UO_83 (O_83,N_23187,N_22952);
nor UO_84 (O_84,N_23167,N_24779);
nand UO_85 (O_85,N_24250,N_23338);
nor UO_86 (O_86,N_24692,N_23667);
nor UO_87 (O_87,N_23546,N_24677);
or UO_88 (O_88,N_23335,N_22914);
and UO_89 (O_89,N_22869,N_24437);
or UO_90 (O_90,N_22850,N_23985);
nor UO_91 (O_91,N_23627,N_22347);
nor UO_92 (O_92,N_22824,N_22093);
or UO_93 (O_93,N_23495,N_24881);
xnor UO_94 (O_94,N_22475,N_24593);
xnor UO_95 (O_95,N_21941,N_22874);
or UO_96 (O_96,N_24852,N_22721);
nand UO_97 (O_97,N_22285,N_23654);
nor UO_98 (O_98,N_22497,N_24281);
or UO_99 (O_99,N_22187,N_23520);
xnor UO_100 (O_100,N_24936,N_23307);
or UO_101 (O_101,N_23444,N_23281);
nor UO_102 (O_102,N_24955,N_24174);
or UO_103 (O_103,N_22578,N_22840);
or UO_104 (O_104,N_24739,N_21947);
or UO_105 (O_105,N_22105,N_24178);
xnor UO_106 (O_106,N_24993,N_22519);
or UO_107 (O_107,N_23605,N_22658);
or UO_108 (O_108,N_22673,N_24271);
nand UO_109 (O_109,N_22936,N_24248);
nor UO_110 (O_110,N_22160,N_24017);
and UO_111 (O_111,N_22432,N_22891);
or UO_112 (O_112,N_22610,N_23880);
or UO_113 (O_113,N_24130,N_24807);
nor UO_114 (O_114,N_21980,N_24447);
nor UO_115 (O_115,N_24679,N_24052);
and UO_116 (O_116,N_22083,N_22341);
and UO_117 (O_117,N_24791,N_24050);
and UO_118 (O_118,N_22225,N_24168);
nand UO_119 (O_119,N_24934,N_22844);
xor UO_120 (O_120,N_24670,N_24790);
and UO_121 (O_121,N_22102,N_21879);
or UO_122 (O_122,N_22117,N_22199);
nor UO_123 (O_123,N_23635,N_21966);
nand UO_124 (O_124,N_23119,N_24047);
nor UO_125 (O_125,N_24502,N_24855);
nor UO_126 (O_126,N_23972,N_23425);
and UO_127 (O_127,N_23263,N_24222);
and UO_128 (O_128,N_24835,N_22138);
and UO_129 (O_129,N_24180,N_23865);
xor UO_130 (O_130,N_23116,N_23956);
and UO_131 (O_131,N_22416,N_22617);
xor UO_132 (O_132,N_24601,N_24104);
nor UO_133 (O_133,N_24205,N_24118);
nor UO_134 (O_134,N_22180,N_23015);
or UO_135 (O_135,N_24945,N_23514);
nand UO_136 (O_136,N_22900,N_24953);
nand UO_137 (O_137,N_23780,N_24812);
and UO_138 (O_138,N_24660,N_23256);
xor UO_139 (O_139,N_24399,N_23121);
and UO_140 (O_140,N_23126,N_23506);
nor UO_141 (O_141,N_22602,N_22325);
and UO_142 (O_142,N_24340,N_24868);
nand UO_143 (O_143,N_22953,N_23696);
or UO_144 (O_144,N_23772,N_22363);
or UO_145 (O_145,N_22934,N_24645);
nor UO_146 (O_146,N_22132,N_22050);
and UO_147 (O_147,N_22637,N_21989);
nor UO_148 (O_148,N_22534,N_23306);
and UO_149 (O_149,N_24474,N_23839);
and UO_150 (O_150,N_22000,N_24471);
nor UO_151 (O_151,N_24236,N_24758);
xnor UO_152 (O_152,N_23395,N_22881);
nand UO_153 (O_153,N_22533,N_22429);
nand UO_154 (O_154,N_22974,N_24682);
or UO_155 (O_155,N_22605,N_22411);
xnor UO_156 (O_156,N_23007,N_24234);
or UO_157 (O_157,N_24803,N_22946);
xor UO_158 (O_158,N_23385,N_23313);
xor UO_159 (O_159,N_24432,N_23528);
nand UO_160 (O_160,N_23095,N_23438);
xor UO_161 (O_161,N_24869,N_22433);
xnor UO_162 (O_162,N_23861,N_22501);
nor UO_163 (O_163,N_21969,N_23678);
or UO_164 (O_164,N_22322,N_22524);
nand UO_165 (O_165,N_23541,N_22444);
or UO_166 (O_166,N_23580,N_24811);
nor UO_167 (O_167,N_22059,N_22486);
xnor UO_168 (O_168,N_24278,N_24794);
and UO_169 (O_169,N_23201,N_23038);
nor UO_170 (O_170,N_23628,N_24169);
xor UO_171 (O_171,N_24971,N_23286);
or UO_172 (O_172,N_24719,N_24767);
xnor UO_173 (O_173,N_22078,N_24170);
nor UO_174 (O_174,N_24082,N_23940);
and UO_175 (O_175,N_24435,N_23160);
nor UO_176 (O_176,N_23109,N_23558);
nand UO_177 (O_177,N_23310,N_23063);
nor UO_178 (O_178,N_22776,N_22818);
and UO_179 (O_179,N_23000,N_22743);
xor UO_180 (O_180,N_24998,N_24596);
or UO_181 (O_181,N_23420,N_24694);
nand UO_182 (O_182,N_23987,N_23782);
nor UO_183 (O_183,N_23887,N_22474);
or UO_184 (O_184,N_24200,N_24142);
and UO_185 (O_185,N_24233,N_23200);
and UO_186 (O_186,N_24663,N_23611);
xnor UO_187 (O_187,N_22420,N_24925);
nor UO_188 (O_188,N_22184,N_24628);
nor UO_189 (O_189,N_22833,N_24750);
or UO_190 (O_190,N_22150,N_21937);
or UO_191 (O_191,N_23097,N_22186);
and UO_192 (O_192,N_23686,N_24098);
nand UO_193 (O_193,N_22626,N_24635);
nand UO_194 (O_194,N_23869,N_23359);
nor UO_195 (O_195,N_22279,N_22599);
nand UO_196 (O_196,N_23001,N_23084);
and UO_197 (O_197,N_23741,N_24573);
nand UO_198 (O_198,N_23598,N_22977);
and UO_199 (O_199,N_22784,N_24806);
nor UO_200 (O_200,N_24454,N_24346);
nand UO_201 (O_201,N_23162,N_24423);
nor UO_202 (O_202,N_23464,N_21993);
and UO_203 (O_203,N_24121,N_23493);
nand UO_204 (O_204,N_22305,N_23459);
or UO_205 (O_205,N_24073,N_22729);
and UO_206 (O_206,N_24644,N_22115);
xor UO_207 (O_207,N_22876,N_24446);
nand UO_208 (O_208,N_23267,N_24989);
or UO_209 (O_209,N_24389,N_23065);
nor UO_210 (O_210,N_22082,N_22084);
or UO_211 (O_211,N_22229,N_23539);
xor UO_212 (O_212,N_23829,N_22509);
xnor UO_213 (O_213,N_23476,N_21913);
or UO_214 (O_214,N_23978,N_24282);
or UO_215 (O_215,N_24633,N_24796);
xor UO_216 (O_216,N_24544,N_23461);
nor UO_217 (O_217,N_21916,N_24283);
nor UO_218 (O_218,N_22568,N_22373);
and UO_219 (O_219,N_24436,N_24853);
nor UO_220 (O_220,N_22940,N_22997);
and UO_221 (O_221,N_23406,N_22383);
nand UO_222 (O_222,N_22308,N_22314);
xor UO_223 (O_223,N_21883,N_24563);
nor UO_224 (O_224,N_21983,N_24976);
and UO_225 (O_225,N_24429,N_23727);
or UO_226 (O_226,N_22087,N_23017);
nand UO_227 (O_227,N_23392,N_23178);
or UO_228 (O_228,N_23954,N_22008);
xnor UO_229 (O_229,N_24614,N_23404);
or UO_230 (O_230,N_24187,N_23156);
nand UO_231 (O_231,N_23994,N_24072);
or UO_232 (O_232,N_24484,N_23469);
nor UO_233 (O_233,N_22871,N_24009);
xor UO_234 (O_234,N_22919,N_22603);
nor UO_235 (O_235,N_24594,N_24287);
nor UO_236 (O_236,N_23342,N_23253);
and UO_237 (O_237,N_23401,N_23749);
xnor UO_238 (O_238,N_22713,N_22631);
and UO_239 (O_239,N_24603,N_24690);
nand UO_240 (O_240,N_23557,N_24861);
nor UO_241 (O_241,N_22031,N_22058);
nor UO_242 (O_242,N_22945,N_23908);
and UO_243 (O_243,N_24964,N_23308);
or UO_244 (O_244,N_22464,N_22636);
or UO_245 (O_245,N_24191,N_23516);
nor UO_246 (O_246,N_23836,N_24476);
and UO_247 (O_247,N_23530,N_21958);
and UO_248 (O_248,N_22757,N_22939);
nor UO_249 (O_249,N_23319,N_24152);
nand UO_250 (O_250,N_22100,N_23456);
and UO_251 (O_251,N_21986,N_23276);
xnor UO_252 (O_252,N_22302,N_22460);
or UO_253 (O_253,N_23744,N_22061);
or UO_254 (O_254,N_23878,N_24638);
or UO_255 (O_255,N_21882,N_22191);
and UO_256 (O_256,N_24725,N_23315);
nor UO_257 (O_257,N_23916,N_22335);
nor UO_258 (O_258,N_23883,N_24753);
nand UO_259 (O_259,N_22365,N_23662);
xnor UO_260 (O_260,N_24887,N_22517);
nand UO_261 (O_261,N_22979,N_23139);
nor UO_262 (O_262,N_21982,N_22136);
and UO_263 (O_263,N_23685,N_22600);
nand UO_264 (O_264,N_24744,N_22894);
or UO_265 (O_265,N_22790,N_22094);
and UO_266 (O_266,N_23052,N_22695);
nor UO_267 (O_267,N_24263,N_24515);
and UO_268 (O_268,N_24658,N_23413);
nor UO_269 (O_269,N_22553,N_21933);
nand UO_270 (O_270,N_24575,N_23230);
nor UO_271 (O_271,N_24108,N_23081);
xor UO_272 (O_272,N_22018,N_24727);
xnor UO_273 (O_273,N_23246,N_23176);
xor UO_274 (O_274,N_23435,N_23630);
nand UO_275 (O_275,N_22829,N_23353);
nand UO_276 (O_276,N_21875,N_24494);
nand UO_277 (O_277,N_23927,N_22613);
nor UO_278 (O_278,N_23213,N_22381);
nor UO_279 (O_279,N_24064,N_24465);
or UO_280 (O_280,N_24318,N_22851);
nor UO_281 (O_281,N_22520,N_24654);
nand UO_282 (O_282,N_24037,N_22689);
or UO_283 (O_283,N_24224,N_22069);
or UO_284 (O_284,N_22356,N_24189);
nor UO_285 (O_285,N_24897,N_24349);
nand UO_286 (O_286,N_22618,N_24330);
xnor UO_287 (O_287,N_24542,N_24828);
xnor UO_288 (O_288,N_22249,N_22633);
nor UO_289 (O_289,N_22539,N_22367);
nand UO_290 (O_290,N_22571,N_24505);
or UO_291 (O_291,N_23170,N_22708);
nor UO_292 (O_292,N_24207,N_22478);
or UO_293 (O_293,N_23781,N_23842);
xnor UO_294 (O_294,N_24260,N_23140);
nand UO_295 (O_295,N_23145,N_22343);
nand UO_296 (O_296,N_23963,N_23262);
nand UO_297 (O_297,N_22137,N_22358);
and UO_298 (O_298,N_23755,N_23365);
nand UO_299 (O_299,N_23374,N_24802);
or UO_300 (O_300,N_24583,N_23946);
nor UO_301 (O_301,N_24031,N_22039);
xnor UO_302 (O_302,N_24039,N_23542);
nand UO_303 (O_303,N_23285,N_23068);
xor UO_304 (O_304,N_24685,N_24345);
nor UO_305 (O_305,N_23364,N_21961);
nand UO_306 (O_306,N_24620,N_23926);
or UO_307 (O_307,N_22537,N_22742);
xor UO_308 (O_308,N_24228,N_22410);
xnor UO_309 (O_309,N_24536,N_22244);
nand UO_310 (O_310,N_24288,N_22906);
and UO_311 (O_311,N_23135,N_24089);
nor UO_312 (O_312,N_22024,N_23463);
nand UO_313 (O_313,N_22144,N_24388);
and UO_314 (O_314,N_24137,N_23606);
nand UO_315 (O_315,N_23161,N_22877);
and UO_316 (O_316,N_24571,N_24499);
xnor UO_317 (O_317,N_21954,N_22677);
nor UO_318 (O_318,N_23497,N_22070);
and UO_319 (O_319,N_22227,N_24456);
nand UO_320 (O_320,N_23673,N_22896);
or UO_321 (O_321,N_24924,N_22588);
nand UO_322 (O_322,N_24404,N_23958);
xnor UO_323 (O_323,N_22287,N_22415);
nand UO_324 (O_324,N_21971,N_21964);
and UO_325 (O_325,N_22660,N_23774);
xnor UO_326 (O_326,N_24935,N_23535);
or UO_327 (O_327,N_22458,N_24451);
xor UO_328 (O_328,N_21881,N_22006);
nand UO_329 (O_329,N_22053,N_24941);
xnor UO_330 (O_330,N_21877,N_24237);
nand UO_331 (O_331,N_23536,N_24400);
and UO_332 (O_332,N_23856,N_24386);
nor UO_333 (O_333,N_23921,N_22814);
or UO_334 (O_334,N_22854,N_22216);
and UO_335 (O_335,N_22931,N_23832);
nand UO_336 (O_336,N_22620,N_22699);
and UO_337 (O_337,N_22357,N_22988);
and UO_338 (O_338,N_22926,N_22212);
or UO_339 (O_339,N_23881,N_23659);
xnor UO_340 (O_340,N_24795,N_22525);
nand UO_341 (O_341,N_23043,N_23860);
and UO_342 (O_342,N_24858,N_23618);
and UO_343 (O_343,N_24167,N_22450);
nor UO_344 (O_344,N_24290,N_24680);
or UO_345 (O_345,N_23903,N_23826);
and UO_346 (O_346,N_22825,N_22858);
nand UO_347 (O_347,N_24041,N_22231);
nand UO_348 (O_348,N_23197,N_22513);
nand UO_349 (O_349,N_24119,N_22294);
and UO_350 (O_350,N_23701,N_22219);
xnor UO_351 (O_351,N_22860,N_24566);
xnor UO_352 (O_352,N_24392,N_22971);
nand UO_353 (O_353,N_24764,N_23393);
nand UO_354 (O_354,N_22108,N_24899);
xor UO_355 (O_355,N_24026,N_23675);
or UO_356 (O_356,N_23078,N_23723);
or UO_357 (O_357,N_23846,N_22387);
nor UO_358 (O_358,N_24341,N_23112);
and UO_359 (O_359,N_24155,N_22473);
and UO_360 (O_360,N_23834,N_22723);
nand UO_361 (O_361,N_23400,N_24621);
xnor UO_362 (O_362,N_24242,N_22516);
or UO_363 (O_363,N_24227,N_22601);
xnor UO_364 (O_364,N_24418,N_23157);
xor UO_365 (O_365,N_23762,N_23235);
and UO_366 (O_366,N_22169,N_23294);
nand UO_367 (O_367,N_22456,N_24141);
nand UO_368 (O_368,N_24561,N_22048);
nor UO_369 (O_369,N_24901,N_23754);
nand UO_370 (O_370,N_23025,N_21979);
nand UO_371 (O_371,N_23988,N_24303);
and UO_372 (O_372,N_24919,N_24259);
nand UO_373 (O_373,N_23202,N_23653);
nand UO_374 (O_374,N_22595,N_22077);
nor UO_375 (O_375,N_23348,N_22002);
and UO_376 (O_376,N_22795,N_23991);
xor UO_377 (O_377,N_22234,N_23284);
or UO_378 (O_378,N_22813,N_22849);
or UO_379 (O_379,N_24957,N_22344);
and UO_380 (O_380,N_24883,N_24933);
nand UO_381 (O_381,N_21960,N_24630);
and UO_382 (O_382,N_24019,N_22622);
or UO_383 (O_383,N_23641,N_24021);
xor UO_384 (O_384,N_24321,N_24642);
or UO_385 (O_385,N_24190,N_24493);
nor UO_386 (O_386,N_23417,N_22074);
or UO_387 (O_387,N_22379,N_22349);
nor UO_388 (O_388,N_24756,N_22674);
nand UO_389 (O_389,N_23871,N_23982);
nor UO_390 (O_390,N_22178,N_23505);
nor UO_391 (O_391,N_23472,N_24123);
nor UO_392 (O_392,N_24525,N_23233);
nand UO_393 (O_393,N_24643,N_23002);
or UO_394 (O_394,N_24212,N_22001);
nor UO_395 (O_395,N_24185,N_22457);
or UO_396 (O_396,N_22937,N_22042);
and UO_397 (O_397,N_23769,N_22856);
or UO_398 (O_398,N_23996,N_23527);
or UO_399 (O_399,N_24410,N_23031);
nand UO_400 (O_400,N_24361,N_22690);
nor UO_401 (O_401,N_23959,N_24095);
nor UO_402 (O_402,N_22238,N_23822);
xor UO_403 (O_403,N_23714,N_24421);
nor UO_404 (O_404,N_23713,N_23237);
xnor UO_405 (O_405,N_24289,N_23106);
xnor UO_406 (O_406,N_22013,N_23733);
and UO_407 (O_407,N_23525,N_23069);
and UO_408 (O_408,N_23273,N_23950);
nor UO_409 (O_409,N_22897,N_23941);
and UO_410 (O_410,N_23864,N_23984);
xnor UO_411 (O_411,N_24972,N_22959);
and UO_412 (O_412,N_24987,N_23934);
nor UO_413 (O_413,N_21957,N_23245);
nor UO_414 (O_414,N_23807,N_24668);
nand UO_415 (O_415,N_22331,N_24970);
nand UO_416 (O_416,N_24929,N_23003);
nor UO_417 (O_417,N_22598,N_24192);
nor UO_418 (O_418,N_23564,N_22656);
and UO_419 (O_419,N_23391,N_23613);
and UO_420 (O_420,N_23368,N_23324);
nor UO_421 (O_421,N_23886,N_24332);
nand UO_422 (O_422,N_23352,N_22451);
nand UO_423 (O_423,N_24818,N_22962);
xor UO_424 (O_424,N_24291,N_23055);
nand UO_425 (O_425,N_23997,N_23101);
or UO_426 (O_426,N_23153,N_24269);
nor UO_427 (O_427,N_23501,N_22301);
or UO_428 (O_428,N_23369,N_23214);
and UO_429 (O_429,N_23144,N_24409);
nand UO_430 (O_430,N_22399,N_22201);
nor UO_431 (O_431,N_22036,N_23023);
xnor UO_432 (O_432,N_22073,N_24698);
or UO_433 (O_433,N_24857,N_24847);
or UO_434 (O_434,N_24003,N_23843);
or UO_435 (O_435,N_24384,N_22175);
or UO_436 (O_436,N_24166,N_23234);
xor UO_437 (O_437,N_24979,N_23973);
or UO_438 (O_438,N_22886,N_24370);
nand UO_439 (O_439,N_22398,N_22046);
and UO_440 (O_440,N_23599,N_22867);
and UO_441 (O_441,N_24268,N_22586);
or UO_442 (O_442,N_24478,N_23643);
or UO_443 (O_443,N_23526,N_23266);
xor UO_444 (O_444,N_23346,N_22183);
xor UO_445 (O_445,N_22815,N_24626);
or UO_446 (O_446,N_23656,N_22007);
xor UO_447 (O_447,N_22467,N_24065);
nor UO_448 (O_448,N_21973,N_22430);
and UO_449 (O_449,N_24202,N_22819);
nor UO_450 (O_450,N_24986,N_22611);
nor UO_451 (O_451,N_24589,N_24210);
xor UO_452 (O_452,N_22655,N_22634);
and UO_453 (O_453,N_22382,N_22461);
and UO_454 (O_454,N_22413,N_23354);
xnor UO_455 (O_455,N_24353,N_22153);
and UO_456 (O_456,N_24742,N_24834);
nor UO_457 (O_457,N_22447,N_22134);
nor UO_458 (O_458,N_22135,N_24938);
nand UO_459 (O_459,N_22259,N_22208);
nand UO_460 (O_460,N_23876,N_23328);
or UO_461 (O_461,N_23298,N_23512);
or UO_462 (O_462,N_23898,N_22885);
nor UO_463 (O_463,N_23247,N_23154);
xor UO_464 (O_464,N_23625,N_24539);
or UO_465 (O_465,N_23798,N_24565);
and UO_466 (O_466,N_23809,N_22276);
or UO_467 (O_467,N_22254,N_21907);
nor UO_468 (O_468,N_23223,N_23243);
and UO_469 (O_469,N_22044,N_24535);
and UO_470 (O_470,N_22049,N_23793);
nor UO_471 (O_471,N_22507,N_24954);
xnor UO_472 (O_472,N_24298,N_22683);
nor UO_473 (O_473,N_21903,N_24163);
and UO_474 (O_474,N_24033,N_24787);
nand UO_475 (O_475,N_23566,N_24879);
and UO_476 (O_476,N_22916,N_24402);
xor UO_477 (O_477,N_22607,N_24352);
or UO_478 (O_478,N_23370,N_22330);
xor UO_479 (O_479,N_22481,N_23386);
nand UO_480 (O_480,N_22290,N_24366);
and UO_481 (O_481,N_23358,N_23347);
or UO_482 (O_482,N_22361,N_22288);
and UO_483 (O_483,N_23366,N_22127);
nand UO_484 (O_484,N_24090,N_24292);
or UO_485 (O_485,N_24467,N_23102);
xnor UO_486 (O_486,N_24075,N_22821);
nand UO_487 (O_487,N_21934,N_23492);
nand UO_488 (O_488,N_24443,N_22404);
or UO_489 (O_489,N_22263,N_22133);
or UO_490 (O_490,N_22720,N_24984);
xnor UO_491 (O_491,N_21949,N_24331);
nand UO_492 (O_492,N_23259,N_22651);
nand UO_493 (O_493,N_24982,N_24792);
and UO_494 (O_494,N_22555,N_24541);
or UO_495 (O_495,N_24173,N_24280);
xnor UO_496 (O_496,N_22671,N_24006);
nor UO_497 (O_497,N_23603,N_24301);
and UO_498 (O_498,N_23715,N_24556);
and UO_499 (O_499,N_24825,N_23848);
nand UO_500 (O_500,N_24179,N_23242);
xor UO_501 (O_501,N_24975,N_22947);
xor UO_502 (O_502,N_24849,N_24444);
xnor UO_503 (O_503,N_23041,N_23105);
nand UO_504 (O_504,N_24056,N_22233);
and UO_505 (O_505,N_23108,N_24475);
or UO_506 (O_506,N_23387,N_24761);
nor UO_507 (O_507,N_22865,N_24963);
nor UO_508 (O_508,N_23373,N_24365);
nor UO_509 (O_509,N_24182,N_22173);
xor UO_510 (O_510,N_23426,N_22676);
or UO_511 (O_511,N_22734,N_22368);
nor UO_512 (O_512,N_23033,N_23434);
nor UO_513 (O_513,N_22751,N_22146);
and UO_514 (O_514,N_22034,N_23917);
or UO_515 (O_515,N_22572,N_22808);
or UO_516 (O_516,N_24285,N_23212);
nand UO_517 (O_517,N_22038,N_24175);
and UO_518 (O_518,N_24531,N_22495);
nand UO_519 (O_519,N_23872,N_22992);
nand UO_520 (O_520,N_22561,N_22556);
xor UO_521 (O_521,N_23799,N_24208);
nor UO_522 (O_522,N_23302,N_23104);
and UO_523 (O_523,N_22128,N_22707);
nor UO_524 (O_524,N_23010,N_22903);
nor UO_525 (O_525,N_22893,N_22510);
nand UO_526 (O_526,N_23032,N_24789);
nor UO_527 (O_527,N_24904,N_24550);
or UO_528 (O_528,N_22804,N_22418);
xor UO_529 (O_529,N_22657,N_22987);
nand UO_530 (O_530,N_22640,N_23051);
nand UO_531 (O_531,N_21976,N_23968);
xor UO_532 (O_532,N_24077,N_21981);
or UO_533 (O_533,N_22438,N_24652);
xor UO_534 (O_534,N_23147,N_22140);
or UO_535 (O_535,N_23716,N_23445);
or UO_536 (O_536,N_23773,N_24942);
or UO_537 (O_537,N_24081,N_22691);
nor UO_538 (O_538,N_23827,N_21914);
or UO_539 (O_539,N_22733,N_23327);
nand UO_540 (O_540,N_23375,N_23828);
xor UO_541 (O_541,N_22627,N_22826);
or UO_542 (O_542,N_22628,N_24769);
nand UO_543 (O_543,N_21994,N_23638);
or UO_544 (O_544,N_22194,N_24691);
and UO_545 (O_545,N_22427,N_22221);
nand UO_546 (O_546,N_22193,N_22581);
nor UO_547 (O_547,N_24115,N_23614);
nand UO_548 (O_548,N_24558,N_23331);
or UO_549 (O_549,N_23951,N_22236);
and UO_550 (O_550,N_22748,N_22930);
nand UO_551 (O_551,N_24311,N_22158);
and UO_552 (O_552,N_24686,N_22727);
nand UO_553 (O_553,N_22593,N_23757);
nand UO_554 (O_554,N_24000,N_22615);
nand UO_555 (O_555,N_22585,N_24619);
and UO_556 (O_556,N_22261,N_24730);
or UO_557 (O_557,N_23819,N_24427);
and UO_558 (O_558,N_24279,N_23981);
xnor UO_559 (O_559,N_24249,N_23999);
xnor UO_560 (O_560,N_22468,N_24647);
and UO_561 (O_561,N_22224,N_21963);
nor UO_562 (O_562,N_22436,N_22337);
or UO_563 (O_563,N_21991,N_23082);
nand UO_564 (O_564,N_24143,N_22831);
nor UO_565 (O_565,N_22960,N_24841);
nand UO_566 (O_566,N_23920,N_24676);
xor UO_567 (O_567,N_24706,N_24914);
nand UO_568 (O_568,N_22296,N_23593);
nor UO_569 (O_569,N_22232,N_24864);
or UO_570 (O_570,N_22807,N_22827);
and UO_571 (O_571,N_22927,N_24569);
nor UO_572 (O_572,N_23491,N_22522);
xor UO_573 (O_573,N_23115,N_22345);
nor UO_574 (O_574,N_22580,N_24270);
xnor UO_575 (O_575,N_23009,N_23220);
xnor UO_576 (O_576,N_22340,N_22025);
nor UO_577 (O_577,N_22284,N_22995);
nor UO_578 (O_578,N_23892,N_23451);
and UO_579 (O_579,N_22498,N_22462);
nand UO_580 (O_580,N_23180,N_23026);
xor UO_581 (O_581,N_23050,N_22145);
nand UO_582 (O_582,N_23455,N_23150);
nand UO_583 (O_583,N_24665,N_23617);
or UO_584 (O_584,N_22577,N_22545);
nand UO_585 (O_585,N_23746,N_22397);
and UO_586 (O_586,N_24966,N_24132);
nor UO_587 (O_587,N_23024,N_23410);
nand UO_588 (O_588,N_23164,N_24995);
xnor UO_589 (O_589,N_24106,N_24748);
or UO_590 (O_590,N_24875,N_22801);
nand UO_591 (O_591,N_22116,N_24693);
nor UO_592 (O_592,N_24948,N_23190);
nor UO_593 (O_593,N_24829,N_24931);
xor UO_594 (O_594,N_22806,N_23899);
nand UO_595 (O_595,N_24856,N_22360);
or UO_596 (O_596,N_22864,N_22923);
xor UO_597 (O_597,N_24528,N_23691);
or UO_598 (O_598,N_24763,N_22226);
nand UO_599 (O_599,N_24592,N_24111);
or UO_600 (O_600,N_24859,N_24755);
and UO_601 (O_601,N_23468,N_22310);
nand UO_602 (O_602,N_24067,N_23334);
nor UO_603 (O_603,N_23014,N_24431);
or UO_604 (O_604,N_21906,N_24977);
or UO_605 (O_605,N_24889,N_23215);
nand UO_606 (O_606,N_24126,N_23742);
xor UO_607 (O_607,N_21876,N_22739);
nor UO_608 (O_608,N_23948,N_22624);
and UO_609 (O_609,N_23339,N_24576);
xnor UO_610 (O_610,N_22587,N_24662);
nand UO_611 (O_611,N_22338,N_23732);
nor UO_612 (O_612,N_23890,N_24253);
nand UO_613 (O_613,N_24203,N_23936);
xor UO_614 (O_614,N_22309,N_23579);
nor UO_615 (O_615,N_23875,N_24479);
nor UO_616 (O_616,N_22015,N_24054);
nand UO_617 (O_617,N_24369,N_22800);
nor UO_618 (O_618,N_24903,N_23107);
nor UO_619 (O_619,N_24981,N_24442);
or UO_620 (O_620,N_22080,N_22260);
nand UO_621 (O_621,N_22983,N_23575);
and UO_622 (O_622,N_23601,N_21927);
nand UO_623 (O_623,N_23665,N_22852);
nand UO_624 (O_624,N_23634,N_23553);
or UO_625 (O_625,N_23537,N_23743);
and UO_626 (O_626,N_22675,N_22455);
and UO_627 (O_627,N_24832,N_24092);
nand UO_628 (O_628,N_23394,N_23330);
nand UO_629 (O_629,N_24932,N_22986);
nand UO_630 (O_630,N_22780,N_24434);
and UO_631 (O_631,N_22514,N_23670);
nand UO_632 (O_632,N_23825,N_23844);
xor UO_633 (O_633,N_24994,N_23447);
xor UO_634 (O_634,N_24457,N_24125);
and UO_635 (O_635,N_23297,N_23709);
or UO_636 (O_636,N_24783,N_22911);
and UO_637 (O_637,N_22765,N_23710);
nand UO_638 (O_638,N_22570,N_24944);
xor UO_639 (O_639,N_22810,N_23693);
xnor UO_640 (O_640,N_24022,N_24681);
nor UO_641 (O_641,N_22889,N_24060);
and UO_642 (O_642,N_22981,N_22129);
nand UO_643 (O_643,N_22425,N_23609);
xor UO_644 (O_644,N_22705,N_23485);
or UO_645 (O_645,N_23228,N_22113);
xnor UO_646 (O_646,N_23123,N_24514);
nor UO_647 (O_647,N_24606,N_22567);
or UO_648 (O_648,N_23552,N_24518);
or UO_649 (O_649,N_23577,N_24516);
or UO_650 (O_650,N_24150,N_24424);
xnor UO_651 (O_651,N_24226,N_22407);
nand UO_652 (O_652,N_24751,N_22802);
xor UO_653 (O_653,N_22667,N_22718);
nor UO_654 (O_654,N_24776,N_22023);
xor UO_655 (O_655,N_24445,N_23067);
nor UO_656 (O_656,N_24615,N_23591);
or UO_657 (O_657,N_22596,N_23407);
nand UO_658 (O_658,N_22215,N_24997);
xor UO_659 (O_659,N_24080,N_23303);
and UO_660 (O_660,N_22921,N_22230);
nor UO_661 (O_661,N_22502,N_22465);
nor UO_662 (O_662,N_24158,N_24042);
nand UO_663 (O_663,N_23479,N_24209);
nor UO_664 (O_664,N_22421,N_23457);
nand UO_665 (O_665,N_24251,N_23964);
nor UO_666 (O_666,N_23048,N_21893);
nor UO_667 (O_667,N_23644,N_23428);
nand UO_668 (O_668,N_22817,N_23570);
nand UO_669 (O_669,N_22245,N_23314);
nand UO_670 (O_670,N_23879,N_22197);
and UO_671 (O_671,N_24070,N_23901);
nand UO_672 (O_672,N_22240,N_24634);
or UO_673 (O_673,N_23448,N_23186);
or UO_674 (O_674,N_22771,N_22439);
xnor UO_675 (O_675,N_22554,N_24325);
and UO_676 (O_676,N_22157,N_22530);
and UO_677 (O_677,N_23657,N_22925);
nand UO_678 (O_678,N_23900,N_23816);
nand UO_679 (O_679,N_24844,N_22887);
xor UO_680 (O_680,N_24612,N_22730);
or UO_681 (O_681,N_24329,N_22546);
or UO_682 (O_682,N_23198,N_23955);
and UO_683 (O_683,N_23127,N_22403);
nor UO_684 (O_684,N_22391,N_24091);
nor UO_685 (O_685,N_23588,N_23681);
nand UO_686 (O_686,N_23833,N_23111);
and UO_687 (O_687,N_23467,N_24165);
or UO_688 (O_688,N_24076,N_23045);
and UO_689 (O_689,N_22722,N_21924);
or UO_690 (O_690,N_24851,N_23529);
and UO_691 (O_691,N_23278,N_23759);
and UO_692 (O_692,N_23012,N_23592);
nor UO_693 (O_693,N_24220,N_24840);
or UO_694 (O_694,N_23735,N_23565);
or UO_695 (O_695,N_22542,N_23309);
nor UO_696 (O_696,N_23362,N_23640);
and UO_697 (O_697,N_24162,N_23522);
xor UO_698 (O_698,N_22118,N_21921);
or UO_699 (O_699,N_22020,N_24616);
xor UO_700 (O_700,N_22336,N_24378);
and UO_701 (O_701,N_22155,N_24112);
or UO_702 (O_702,N_24714,N_24598);
and UO_703 (O_703,N_24512,N_22861);
xnor UO_704 (O_704,N_22071,N_24845);
xnor UO_705 (O_705,N_22222,N_24653);
nand UO_706 (O_706,N_23726,N_22021);
nand UO_707 (O_707,N_23623,N_24962);
or UO_708 (O_708,N_24640,N_24215);
nand UO_709 (O_709,N_22999,N_23862);
nand UO_710 (O_710,N_23787,N_24472);
xnor UO_711 (O_711,N_24607,N_24532);
or UO_712 (O_712,N_22092,N_24562);
xor UO_713 (O_713,N_23034,N_23870);
and UO_714 (O_714,N_23943,N_24358);
and UO_715 (O_715,N_24231,N_24688);
and UO_716 (O_716,N_22270,N_23704);
nand UO_717 (O_717,N_24186,N_22863);
nand UO_718 (O_718,N_23036,N_22648);
nor UO_719 (O_719,N_22400,N_22879);
nor UO_720 (O_720,N_22033,N_22505);
nand UO_721 (O_721,N_24027,N_22003);
or UO_722 (O_722,N_23791,N_24498);
xor UO_723 (O_723,N_24646,N_23989);
xnor UO_724 (O_724,N_24005,N_22437);
xor UO_725 (O_725,N_24814,N_23022);
xnor UO_726 (O_726,N_24046,N_23572);
nor UO_727 (O_727,N_24778,N_21972);
nand UO_728 (O_728,N_24822,N_22179);
nor UO_729 (O_729,N_24567,N_22258);
and UO_730 (O_730,N_23454,N_22719);
xor UO_731 (O_731,N_24673,N_23970);
nor UO_732 (O_732,N_23470,N_24735);
and UO_733 (O_733,N_23312,N_22579);
xnor UO_734 (O_734,N_24772,N_24597);
or UO_735 (O_735,N_22778,N_24309);
nor UO_736 (O_736,N_22968,N_24622);
and UO_737 (O_737,N_24552,N_24557);
nand UO_738 (O_738,N_24310,N_23705);
and UO_739 (O_739,N_23680,N_22482);
nor UO_740 (O_740,N_24913,N_21968);
and UO_741 (O_741,N_23381,N_24413);
and UO_742 (O_742,N_24069,N_23274);
nand UO_743 (O_743,N_22731,N_24109);
xor UO_744 (O_744,N_24230,N_23057);
or UO_745 (O_745,N_21889,N_22299);
xor UO_746 (O_746,N_21992,N_22712);
xor UO_747 (O_747,N_23573,N_24216);
xnor UO_748 (O_748,N_22898,N_23408);
or UO_749 (O_749,N_22203,N_24943);
and UO_750 (O_750,N_23962,N_24871);
nand UO_751 (O_751,N_22786,N_21956);
xor UO_752 (O_752,N_22955,N_22441);
xor UO_753 (O_753,N_23877,N_23857);
nand UO_754 (O_754,N_24809,N_24759);
nand UO_755 (O_755,N_22273,N_22540);
nor UO_756 (O_756,N_23942,N_23806);
nand UO_757 (O_757,N_21977,N_23724);
and UO_758 (O_758,N_23134,N_21894);
and UO_759 (O_759,N_22646,N_22075);
or UO_760 (O_760,N_22239,N_23021);
and UO_761 (O_761,N_23288,N_24988);
or UO_762 (O_762,N_23053,N_23498);
nor UO_763 (O_763,N_23545,N_23775);
nor UO_764 (O_764,N_23770,N_24351);
nand UO_765 (O_765,N_22969,N_22111);
xnor UO_766 (O_766,N_24153,N_24385);
nand UO_767 (O_767,N_23938,N_22307);
nor UO_768 (O_768,N_24793,N_22011);
nand UO_769 (O_769,N_24743,N_24426);
xnor UO_770 (O_770,N_24015,N_22692);
nand UO_771 (O_771,N_23783,N_24160);
and UO_772 (O_772,N_23257,N_22716);
and UO_773 (O_773,N_24746,N_22774);
or UO_774 (O_774,N_22932,N_22592);
and UO_775 (O_775,N_24757,N_22782);
xnor UO_776 (O_776,N_24452,N_21922);
or UO_777 (O_777,N_24637,N_22242);
xnor UO_778 (O_778,N_24551,N_24316);
xnor UO_779 (O_779,N_24946,N_22315);
nand UO_780 (O_780,N_24580,N_22289);
xnor UO_781 (O_781,N_24302,N_23597);
nand UO_782 (O_782,N_23194,N_22174);
xor UO_783 (O_783,N_23906,N_22396);
nand UO_784 (O_784,N_24156,N_23199);
xor UO_785 (O_785,N_22875,N_24415);
and UO_786 (O_786,N_23289,N_24347);
or UO_787 (O_787,N_22332,N_24213);
nor UO_788 (O_788,N_23183,N_23211);
and UO_789 (O_789,N_23835,N_23549);
nand UO_790 (O_790,N_23687,N_23035);
and UO_791 (O_791,N_23703,N_24991);
nor UO_792 (O_792,N_24483,N_22326);
or UO_793 (O_793,N_24462,N_23543);
nor UO_794 (O_794,N_24266,N_24229);
xnor UO_795 (O_795,N_23576,N_22327);
and UO_796 (O_796,N_24320,N_24327);
or UO_797 (O_797,N_21943,N_22248);
or UO_798 (O_798,N_23889,N_22385);
nor UO_799 (O_799,N_24395,N_23503);
and UO_800 (O_800,N_22759,N_22684);
xor UO_801 (O_801,N_22766,N_21985);
and UO_802 (O_802,N_24117,N_22868);
nand UO_803 (O_803,N_23849,N_24773);
or UO_804 (O_804,N_23642,N_23188);
nand UO_805 (O_805,N_22256,N_22944);
or UO_806 (O_806,N_23452,N_23287);
xor UO_807 (O_807,N_24008,N_22755);
or UO_808 (O_808,N_22384,N_22538);
and UO_809 (O_809,N_24823,N_23712);
xnor UO_810 (O_810,N_22961,N_24350);
nand UO_811 (O_811,N_23818,N_23326);
nor UO_812 (O_812,N_22924,N_22255);
xnor UO_813 (O_813,N_22312,N_23953);
and UO_814 (O_814,N_23311,N_23939);
xnor UO_815 (O_815,N_22688,N_24749);
nand UO_816 (O_816,N_22453,N_22147);
nand UO_817 (O_817,N_22710,N_23152);
or UO_818 (O_818,N_24843,N_22463);
nor UO_819 (O_819,N_24171,N_23195);
or UO_820 (O_820,N_21890,N_24529);
and UO_821 (O_821,N_24338,N_23888);
xnor UO_822 (O_822,N_23396,N_23090);
and UO_823 (O_823,N_23986,N_23786);
nand UO_824 (O_824,N_23897,N_22619);
nand UO_825 (O_825,N_22687,N_23894);
and UO_826 (O_826,N_22032,N_22551);
and UO_827 (O_827,N_23684,N_24211);
nor UO_828 (O_828,N_24960,N_22725);
nand UO_829 (O_829,N_23992,N_23397);
or UO_830 (O_830,N_22697,N_22109);
and UO_831 (O_831,N_23087,N_22386);
nor UO_832 (O_832,N_23019,N_24584);
nor UO_833 (O_833,N_24605,N_23474);
and UO_834 (O_834,N_23648,N_22182);
and UO_835 (O_835,N_21978,N_23719);
or UO_836 (O_836,N_24838,N_24826);
nand UO_837 (O_837,N_22709,N_21959);
nand UO_838 (O_838,N_23254,N_23481);
and UO_839 (O_839,N_21929,N_21887);
xnor UO_840 (O_840,N_23133,N_22761);
and UO_841 (O_841,N_24579,N_24738);
xnor UO_842 (O_842,N_22012,N_22862);
nor UO_843 (O_843,N_22445,N_24380);
nor UO_844 (O_844,N_21945,N_24648);
or UO_845 (O_845,N_23502,N_21970);
xnor UO_846 (O_846,N_24771,N_24470);
nand UO_847 (O_847,N_23935,N_22642);
or UO_848 (O_848,N_22576,N_22122);
xor UO_849 (O_849,N_22805,N_24521);
and UO_850 (O_850,N_24372,N_23521);
or UO_851 (O_851,N_23388,N_24193);
xnor UO_852 (O_852,N_22756,N_24276);
and UO_853 (O_853,N_22223,N_24035);
nor UO_854 (O_854,N_24188,N_21900);
xor UO_855 (O_855,N_23221,N_22834);
xnor UO_856 (O_856,N_23753,N_24299);
and UO_857 (O_857,N_21951,N_24506);
and UO_858 (O_858,N_23416,N_23238);
xnor UO_859 (O_859,N_24002,N_24723);
xor UO_860 (O_860,N_23608,N_24905);
and UO_861 (O_861,N_24817,N_23868);
nand UO_862 (O_862,N_23866,N_24194);
nand UO_863 (O_863,N_22686,N_23018);
nor UO_864 (O_864,N_22489,N_22728);
nand UO_865 (O_865,N_21996,N_22635);
and UO_866 (O_866,N_22027,N_22777);
xor UO_867 (O_867,N_24705,N_23442);
nand UO_868 (O_868,N_24689,N_24958);
nand UO_869 (O_869,N_23582,N_22746);
nand UO_870 (O_870,N_22665,N_22275);
nand UO_871 (O_871,N_23767,N_24854);
nor UO_872 (O_872,N_22511,N_22292);
xor UO_873 (O_873,N_22353,N_24450);
nor UO_874 (O_874,N_22280,N_23688);
xnor UO_875 (O_875,N_24071,N_23867);
and UO_876 (O_876,N_22544,N_23619);
nand UO_877 (O_877,N_22750,N_24508);
and UO_878 (O_878,N_23692,N_24715);
xor UO_879 (O_879,N_22362,N_22394);
or UO_880 (O_880,N_24068,N_21899);
xnor UO_881 (O_881,N_23118,N_23029);
and UO_882 (O_882,N_23969,N_22099);
nand UO_883 (O_883,N_22004,N_23666);
nor UO_884 (O_884,N_24780,N_24201);
and UO_885 (O_885,N_22902,N_23091);
or UO_886 (O_886,N_24669,N_23453);
and UO_887 (O_887,N_23478,N_22142);
and UO_888 (O_888,N_21967,N_24649);
or UO_889 (O_889,N_24487,N_24140);
and UO_890 (O_890,N_24708,N_23587);
nor UO_891 (O_891,N_23507,N_23344);
and UO_892 (O_892,N_24217,N_21926);
and UO_893 (O_893,N_22218,N_22735);
nor UO_894 (O_894,N_23098,N_24886);
and UO_895 (O_895,N_22951,N_23363);
and UO_896 (O_896,N_24961,N_24798);
xor UO_897 (O_897,N_23569,N_22678);
or UO_898 (O_898,N_22278,N_24387);
nand UO_899 (O_899,N_24011,N_23544);
or UO_900 (O_900,N_23141,N_23891);
and UO_901 (O_901,N_22214,N_24600);
or UO_902 (O_902,N_24821,N_24218);
nor UO_903 (O_903,N_23292,N_24926);
and UO_904 (O_904,N_23423,N_23061);
nand UO_905 (O_905,N_24323,N_22878);
or UO_906 (O_906,N_21897,N_24980);
or UO_907 (O_907,N_24240,N_23046);
nor UO_908 (O_908,N_23624,N_24774);
nor UO_909 (O_909,N_21918,N_23255);
and UO_910 (O_910,N_24734,N_24636);
nor UO_911 (O_911,N_23821,N_22496);
or UO_912 (O_912,N_24074,N_24085);
nand UO_913 (O_913,N_24243,N_24564);
nor UO_914 (O_914,N_23929,N_22528);
or UO_915 (O_915,N_24860,N_23998);
xor UO_916 (O_916,N_23136,N_24745);
xor UO_917 (O_917,N_24937,N_23855);
nand UO_918 (O_918,N_22500,N_22741);
nand UO_919 (O_919,N_22908,N_24131);
nand UO_920 (O_920,N_24511,N_23854);
nand UO_921 (O_921,N_24430,N_22442);
xnor UO_922 (O_922,N_22492,N_24275);
nand UO_923 (O_923,N_24656,N_22682);
and UO_924 (O_924,N_22170,N_24221);
xor UO_925 (O_925,N_22414,N_22202);
nand UO_926 (O_926,N_24135,N_23040);
or UO_927 (O_927,N_24468,N_22063);
nor UO_928 (O_928,N_23961,N_23129);
nand UO_929 (O_929,N_21920,N_24928);
or UO_930 (O_930,N_22176,N_24401);
and UO_931 (O_931,N_22371,N_22479);
or UO_932 (O_932,N_23585,N_23475);
nand UO_933 (O_933,N_22164,N_22246);
nor UO_934 (O_934,N_22573,N_23291);
xnor UO_935 (O_935,N_22998,N_23430);
xnor UO_936 (O_936,N_24733,N_23013);
nand UO_937 (O_937,N_23458,N_21995);
nor UO_938 (O_938,N_21988,N_23884);
xor UO_939 (O_939,N_24819,N_22872);
nand UO_940 (O_940,N_24151,N_22333);
and UO_941 (O_941,N_24540,N_24425);
and UO_942 (O_942,N_22590,N_22910);
and UO_943 (O_943,N_22181,N_23380);
and UO_944 (O_944,N_24241,N_24895);
nand UO_945 (O_945,N_24144,N_23484);
nor UO_946 (O_946,N_24099,N_23429);
and UO_947 (O_947,N_22976,N_24393);
or UO_948 (O_948,N_21946,N_24902);
and UO_949 (O_949,N_22454,N_22306);
and UO_950 (O_950,N_23885,N_23594);
nand UO_951 (O_951,N_23914,N_22088);
or UO_952 (O_952,N_22098,N_22612);
nor UO_953 (O_953,N_23823,N_24560);
or UO_954 (O_954,N_23486,N_22839);
nand UO_955 (O_955,N_23179,N_22789);
xor UO_956 (O_956,N_22714,N_21895);
or UO_957 (O_957,N_24322,N_23477);
nor UO_958 (O_958,N_22188,N_22736);
nor UO_959 (O_959,N_22274,N_24088);
and UO_960 (O_960,N_22913,N_22772);
and UO_961 (O_961,N_22753,N_23928);
nor UO_962 (O_962,N_23158,N_23172);
nor UO_963 (O_963,N_23027,N_24831);
xor UO_964 (O_964,N_21952,N_24820);
nor UO_965 (O_965,N_22785,N_22529);
nand UO_966 (O_966,N_23236,N_24770);
nand UO_967 (O_967,N_24507,N_22388);
xor UO_968 (O_968,N_22095,N_22985);
and UO_969 (O_969,N_23677,N_23066);
nor UO_970 (O_970,N_22811,N_24877);
nor UO_971 (O_971,N_22217,N_22629);
and UO_972 (O_972,N_24496,N_23293);
nand UO_973 (O_973,N_23655,N_23316);
xnor UO_974 (O_974,N_22196,N_24463);
nand UO_975 (O_975,N_23383,N_23372);
nand UO_976 (O_976,N_24664,N_23551);
and UO_977 (O_977,N_24063,N_23805);
or UO_978 (O_978,N_24729,N_23804);
and UO_979 (O_979,N_23815,N_24214);
nor UO_980 (O_980,N_24124,N_22562);
nor UO_981 (O_981,N_23004,N_24286);
nand UO_982 (O_982,N_24827,N_22744);
or UO_983 (O_983,N_23208,N_23621);
nand UO_984 (O_984,N_22060,N_23103);
or UO_985 (O_985,N_22119,N_23225);
xnor UO_986 (O_986,N_23169,N_23515);
and UO_987 (O_987,N_22163,N_23616);
xor UO_988 (O_988,N_24138,N_24724);
or UO_989 (O_989,N_23099,N_23540);
or UO_990 (O_990,N_22148,N_24440);
nor UO_991 (O_991,N_23824,N_21930);
or UO_992 (O_992,N_22374,N_24956);
nand UO_993 (O_993,N_22342,N_22929);
or UO_994 (O_994,N_23707,N_24025);
nand UO_995 (O_995,N_24016,N_21987);
nand UO_996 (O_996,N_24830,N_23483);
and UO_997 (O_997,N_22773,N_23532);
nor UO_998 (O_998,N_24093,N_24524);
or UO_999 (O_999,N_22423,N_24582);
or UO_1000 (O_1000,N_23831,N_22663);
nand UO_1001 (O_1001,N_24718,N_23077);
or UO_1002 (O_1002,N_22653,N_24157);
nor UO_1003 (O_1003,N_22317,N_24034);
nor UO_1004 (O_1004,N_23037,N_23694);
and UO_1005 (O_1005,N_23604,N_22838);
nand UO_1006 (O_1006,N_24870,N_23062);
nor UO_1007 (O_1007,N_22028,N_23771);
nor UO_1008 (O_1008,N_23971,N_22506);
nand UO_1009 (O_1009,N_23513,N_22942);
or UO_1010 (O_1010,N_24284,N_24721);
xnor UO_1011 (O_1011,N_22724,N_23995);
xnor UO_1012 (O_1012,N_22487,N_22319);
xor UO_1013 (O_1013,N_23361,N_24252);
nor UO_1014 (O_1014,N_24639,N_23351);
or UO_1015 (O_1015,N_23509,N_23651);
and UO_1016 (O_1016,N_24459,N_22068);
nand UO_1017 (O_1017,N_23421,N_23290);
xnor UO_1018 (O_1018,N_22541,N_22401);
xor UO_1019 (O_1019,N_24900,N_22017);
or UO_1020 (O_1020,N_23706,N_24741);
or UO_1021 (O_1021,N_22668,N_24148);
or UO_1022 (O_1022,N_22738,N_23622);
xor UO_1023 (O_1023,N_24930,N_23499);
and UO_1024 (O_1024,N_22933,N_22958);
and UO_1025 (O_1025,N_23663,N_24526);
nor UO_1026 (O_1026,N_24406,N_24489);
or UO_1027 (O_1027,N_23143,N_23224);
and UO_1028 (O_1028,N_22171,N_24513);
and UO_1029 (O_1029,N_23252,N_24523);
nand UO_1030 (O_1030,N_24842,N_24461);
nor UO_1031 (O_1031,N_23059,N_24891);
nand UO_1032 (O_1032,N_21891,N_23130);
xnor UO_1033 (O_1033,N_24709,N_22304);
nor UO_1034 (O_1034,N_22406,N_24357);
nor UO_1035 (O_1035,N_24371,N_22469);
and UO_1036 (O_1036,N_24477,N_24147);
or UO_1037 (O_1037,N_23206,N_23776);
or UO_1038 (O_1038,N_23189,N_24547);
nor UO_1039 (O_1039,N_23909,N_23761);
nand UO_1040 (O_1040,N_24590,N_23433);
nand UO_1041 (O_1041,N_24509,N_23952);
or UO_1042 (O_1042,N_23207,N_21948);
nor UO_1043 (O_1043,N_23911,N_23251);
nand UO_1044 (O_1044,N_23664,N_24568);
nand UO_1045 (O_1045,N_24805,N_22645);
or UO_1046 (O_1046,N_22089,N_22466);
xor UO_1047 (O_1047,N_22957,N_24355);
nor UO_1048 (O_1048,N_23301,N_24604);
nor UO_1049 (O_1049,N_24973,N_24595);
and UO_1050 (O_1050,N_22085,N_24473);
nand UO_1051 (O_1051,N_22966,N_23439);
xor UO_1052 (O_1052,N_22954,N_24317);
and UO_1053 (O_1053,N_23738,N_22271);
xor UO_1054 (O_1054,N_22594,N_24740);
and UO_1055 (O_1055,N_22243,N_23519);
or UO_1056 (O_1056,N_24765,N_24172);
nand UO_1057 (O_1057,N_22575,N_24267);
and UO_1058 (O_1058,N_22518,N_23054);
and UO_1059 (O_1059,N_22779,N_22177);
and UO_1060 (O_1060,N_22694,N_24839);
and UO_1061 (O_1061,N_21925,N_22066);
xnor UO_1062 (O_1062,N_22832,N_23697);
or UO_1063 (O_1063,N_22472,N_24379);
and UO_1064 (O_1064,N_22200,N_24555);
or UO_1065 (O_1065,N_22715,N_22131);
or UO_1066 (O_1066,N_24128,N_22262);
or UO_1067 (O_1067,N_23931,N_22130);
nor UO_1068 (O_1068,N_23318,N_24333);
and UO_1069 (O_1069,N_24951,N_23649);
or UO_1070 (O_1070,N_22067,N_22419);
or UO_1071 (O_1071,N_23282,N_24334);
and UO_1072 (O_1072,N_22064,N_23011);
nand UO_1073 (O_1073,N_23837,N_22035);
xor UO_1074 (O_1074,N_24045,N_23717);
nand UO_1075 (O_1075,N_24578,N_22366);
and UO_1076 (O_1076,N_24195,N_22632);
nand UO_1077 (O_1077,N_24888,N_23271);
and UO_1078 (O_1078,N_22547,N_21962);
nor UO_1079 (O_1079,N_24713,N_21997);
nand UO_1080 (O_1080,N_24307,N_23431);
and UO_1081 (O_1081,N_23852,N_22282);
xnor UO_1082 (O_1082,N_24522,N_24650);
and UO_1083 (O_1083,N_22698,N_23933);
and UO_1084 (O_1084,N_23838,N_22747);
xor UO_1085 (O_1085,N_22884,N_22268);
or UO_1086 (O_1086,N_23589,N_23979);
nand UO_1087 (O_1087,N_22369,N_24374);
nor UO_1088 (O_1088,N_22405,N_23450);
nand UO_1089 (O_1089,N_22220,N_24920);
and UO_1090 (O_1090,N_22047,N_23645);
nand UO_1091 (O_1091,N_23722,N_23222);
nor UO_1092 (O_1092,N_23122,N_24294);
nor UO_1093 (O_1093,N_23056,N_21878);
xnor UO_1094 (O_1094,N_24417,N_23113);
xor UO_1095 (O_1095,N_24314,N_24611);
or UO_1096 (O_1096,N_23083,N_24985);
nand UO_1097 (O_1097,N_24262,N_22072);
xor UO_1098 (O_1098,N_22693,N_23260);
xor UO_1099 (O_1099,N_24554,N_22393);
and UO_1100 (O_1100,N_23006,N_24717);
or UO_1101 (O_1101,N_24588,N_23910);
nor UO_1102 (O_1102,N_22791,N_23414);
xnor UO_1103 (O_1103,N_21974,N_24519);
and UO_1104 (O_1104,N_22045,N_22948);
and UO_1105 (O_1105,N_24700,N_22198);
nand UO_1106 (O_1106,N_23560,N_24255);
xnor UO_1107 (O_1107,N_22717,N_24177);
nor UO_1108 (O_1108,N_24712,N_24572);
nand UO_1109 (O_1109,N_22650,N_23241);
nor UO_1110 (O_1110,N_24335,N_23080);
or UO_1111 (O_1111,N_22470,N_22471);
nor UO_1112 (O_1112,N_22297,N_24548);
and UO_1113 (O_1113,N_23626,N_23329);
and UO_1114 (O_1114,N_21912,N_23336);
and UO_1115 (O_1115,N_24863,N_22964);
xor UO_1116 (O_1116,N_24364,N_23249);
or UO_1117 (O_1117,N_24848,N_22029);
or UO_1118 (O_1118,N_22799,N_24362);
nor UO_1119 (O_1119,N_21898,N_24134);
or UO_1120 (O_1120,N_24254,N_22535);
nand UO_1121 (O_1121,N_23830,N_22125);
or UO_1122 (O_1122,N_21931,N_22836);
xnor UO_1123 (O_1123,N_24272,N_24710);
nor UO_1124 (O_1124,N_22809,N_22967);
or UO_1125 (O_1125,N_23734,N_23578);
nor UO_1126 (O_1126,N_24407,N_22395);
and UO_1127 (O_1127,N_23355,N_24884);
or UO_1128 (O_1128,N_22041,N_24136);
or UO_1129 (O_1129,N_23016,N_22126);
nor UO_1130 (O_1130,N_24609,N_23424);
or UO_1131 (O_1131,N_22643,N_24617);
nand UO_1132 (O_1132,N_23110,N_24087);
nor UO_1133 (O_1133,N_22159,N_22412);
nand UO_1134 (O_1134,N_24629,N_22770);
xor UO_1135 (O_1135,N_23277,N_23548);
nor UO_1136 (O_1136,N_24882,N_22354);
xnor UO_1137 (O_1137,N_22189,N_22798);
nand UO_1138 (O_1138,N_22167,N_22904);
xnor UO_1139 (O_1139,N_24359,N_24079);
xnor UO_1140 (O_1140,N_23138,N_23555);
nand UO_1141 (O_1141,N_24133,N_22848);
xor UO_1142 (O_1142,N_22970,N_22477);
xor UO_1143 (O_1143,N_24277,N_23072);
or UO_1144 (O_1144,N_23490,N_24799);
nand UO_1145 (O_1145,N_21939,N_24244);
or UO_1146 (O_1146,N_23765,N_23918);
and UO_1147 (O_1147,N_23731,N_21950);
or UO_1148 (O_1148,N_22935,N_24146);
nand UO_1149 (O_1149,N_22652,N_24326);
nand UO_1150 (O_1150,N_23210,N_24486);
and UO_1151 (O_1151,N_23554,N_24917);
nor UO_1152 (O_1152,N_24306,N_23064);
and UO_1153 (O_1153,N_22996,N_23768);
or UO_1154 (O_1154,N_23422,N_24293);
or UO_1155 (O_1155,N_23792,N_24788);
nand UO_1156 (O_1156,N_23174,N_23356);
nand UO_1157 (O_1157,N_24176,N_24149);
xnor UO_1158 (O_1158,N_24916,N_23231);
nor UO_1159 (O_1159,N_24246,N_22899);
or UO_1160 (O_1160,N_22843,N_24198);
xnor UO_1161 (O_1161,N_22172,N_22609);
or UO_1162 (O_1162,N_23304,N_23449);
nand UO_1163 (O_1163,N_23796,N_24574);
nand UO_1164 (O_1164,N_21932,N_22149);
xor UO_1165 (O_1165,N_24543,N_24659);
nor UO_1166 (O_1166,N_23487,N_22696);
or UO_1167 (O_1167,N_24094,N_22978);
xor UO_1168 (O_1168,N_22376,N_23132);
nor UO_1169 (O_1169,N_23272,N_22272);
and UO_1170 (O_1170,N_24546,N_23402);
xnor UO_1171 (O_1171,N_23155,N_24100);
and UO_1172 (O_1172,N_23305,N_24235);
nor UO_1173 (O_1173,N_22359,N_22162);
nor UO_1174 (O_1174,N_24018,N_23882);
xnor UO_1175 (O_1175,N_24549,N_22982);
or UO_1176 (O_1176,N_22775,N_24720);
nand UO_1177 (O_1177,N_23269,N_23584);
and UO_1178 (O_1178,N_24066,N_22014);
nand UO_1179 (O_1179,N_24497,N_24927);
or UO_1180 (O_1180,N_22569,N_22380);
nor UO_1181 (O_1181,N_22096,N_23367);
xor UO_1182 (O_1182,N_23740,N_24587);
and UO_1183 (O_1183,N_24501,N_24722);
nor UO_1184 (O_1184,N_24120,N_24768);
nor UO_1185 (O_1185,N_24258,N_21940);
nor UO_1186 (O_1186,N_23923,N_23473);
xor UO_1187 (O_1187,N_23049,N_22584);
or UO_1188 (O_1188,N_23567,N_24097);
nand UO_1189 (O_1189,N_22956,N_22892);
nand UO_1190 (O_1190,N_24398,N_24107);
nand UO_1191 (O_1191,N_24850,N_24319);
xnor UO_1192 (O_1192,N_22206,N_23088);
xor UO_1193 (O_1193,N_23814,N_24439);
xor UO_1194 (O_1194,N_23841,N_22606);
or UO_1195 (O_1195,N_24808,N_23586);
nor UO_1196 (O_1196,N_24801,N_23060);
and UO_1197 (O_1197,N_23020,N_22185);
nor UO_1198 (O_1198,N_23562,N_24538);
and UO_1199 (O_1199,N_22026,N_24867);
or UO_1200 (O_1200,N_22846,N_22672);
xor UO_1201 (O_1201,N_24495,N_22269);
or UO_1202 (O_1202,N_24585,N_24032);
or UO_1203 (O_1203,N_23800,N_22030);
or UO_1204 (O_1204,N_24704,N_23652);
xor UO_1205 (O_1205,N_24049,N_22975);
nand UO_1206 (O_1206,N_24784,N_22941);
or UO_1207 (O_1207,N_22993,N_22352);
xnor UO_1208 (O_1208,N_24731,N_23779);
nor UO_1209 (O_1209,N_22565,N_22503);
nand UO_1210 (O_1210,N_22334,N_23333);
xnor UO_1211 (O_1211,N_23390,N_22973);
nor UO_1212 (O_1212,N_22532,N_22112);
and UO_1213 (O_1213,N_23405,N_22855);
and UO_1214 (O_1214,N_24048,N_23096);
and UO_1215 (O_1215,N_21911,N_24959);
and UO_1216 (O_1216,N_22706,N_24974);
xnor UO_1217 (O_1217,N_23042,N_23398);
or UO_1218 (O_1218,N_24315,N_23137);
nand UO_1219 (O_1219,N_22293,N_23974);
xor UO_1220 (O_1220,N_24274,N_23270);
nand UO_1221 (O_1221,N_24304,N_23203);
nand UO_1222 (O_1222,N_23279,N_22123);
xor UO_1223 (O_1223,N_22760,N_23296);
or UO_1224 (O_1224,N_22531,N_24339);
xor UO_1225 (O_1225,N_24530,N_23845);
and UO_1226 (O_1226,N_22346,N_23280);
or UO_1227 (O_1227,N_22984,N_23322);
and UO_1228 (O_1228,N_23494,N_23788);
nand UO_1229 (O_1229,N_22654,N_23660);
nand UO_1230 (O_1230,N_22591,N_22557);
nand UO_1231 (O_1231,N_24952,N_24968);
xnor UO_1232 (O_1232,N_24898,N_24245);
xor UO_1233 (O_1233,N_22994,N_22266);
nand UO_1234 (O_1234,N_22560,N_23419);
nor UO_1235 (O_1235,N_24145,N_24683);
and UO_1236 (O_1236,N_23748,N_23668);
or UO_1237 (O_1237,N_23093,N_23547);
nor UO_1238 (O_1238,N_22484,N_23976);
xor UO_1239 (O_1239,N_22251,N_22311);
or UO_1240 (O_1240,N_23384,N_22250);
xor UO_1241 (O_1241,N_23092,N_24762);
or UO_1242 (O_1242,N_22549,N_22209);
xor UO_1243 (O_1243,N_24024,N_21975);
and UO_1244 (O_1244,N_23764,N_23275);
and UO_1245 (O_1245,N_21909,N_22252);
nor UO_1246 (O_1246,N_22847,N_23563);
or UO_1247 (O_1247,N_22625,N_23760);
nand UO_1248 (O_1248,N_23345,N_24004);
xnor UO_1249 (O_1249,N_24661,N_22139);
nand UO_1250 (O_1250,N_22491,N_24481);
nand UO_1251 (O_1251,N_23165,N_23008);
xor UO_1252 (O_1252,N_22377,N_23993);
or UO_1253 (O_1253,N_23508,N_24813);
xor UO_1254 (O_1254,N_24674,N_24373);
xnor UO_1255 (O_1255,N_23218,N_24247);
nor UO_1256 (O_1256,N_24308,N_23698);
and UO_1257 (O_1257,N_24702,N_22114);
and UO_1258 (O_1258,N_21910,N_23376);
and UO_1259 (O_1259,N_23184,N_22907);
nand UO_1260 (O_1260,N_24020,N_23432);
nor UO_1261 (O_1261,N_23639,N_22499);
xnor UO_1262 (O_1262,N_23674,N_21984);
xor UO_1263 (O_1263,N_22054,N_24999);
and UO_1264 (O_1264,N_24785,N_24113);
or UO_1265 (O_1265,N_24969,N_22661);
xor UO_1266 (O_1266,N_24375,N_23332);
or UO_1267 (O_1267,N_23794,N_23465);
nand UO_1268 (O_1268,N_24449,N_22638);
and UO_1269 (O_1269,N_24703,N_22630);
nor UO_1270 (O_1270,N_23446,N_23647);
and UO_1271 (O_1271,N_23682,N_22558);
or UO_1272 (O_1272,N_22097,N_23607);
nand UO_1273 (O_1273,N_24114,N_22845);
nand UO_1274 (O_1274,N_22681,N_24695);
xor UO_1275 (O_1275,N_24485,N_23248);
xnor UO_1276 (O_1276,N_23403,N_24553);
and UO_1277 (O_1277,N_23517,N_23851);
or UO_1278 (O_1278,N_23817,N_24599);
and UO_1279 (O_1279,N_24657,N_22052);
and UO_1280 (O_1280,N_23847,N_23227);
and UO_1281 (O_1281,N_23489,N_24950);
nand UO_1282 (O_1282,N_22965,N_23100);
or UO_1283 (O_1283,N_22812,N_23415);
nor UO_1284 (O_1284,N_24023,N_21901);
nand UO_1285 (O_1285,N_21905,N_23913);
nand UO_1286 (O_1286,N_22351,N_24701);
nor UO_1287 (O_1287,N_22597,N_24625);
nand UO_1288 (O_1288,N_22822,N_23785);
nand UO_1289 (O_1289,N_24343,N_23382);
and UO_1290 (O_1290,N_24038,N_24013);
nor UO_1291 (O_1291,N_22523,N_23912);
xnor UO_1292 (O_1292,N_22917,N_23340);
or UO_1293 (O_1293,N_22210,N_22483);
or UO_1294 (O_1294,N_22402,N_24420);
nand UO_1295 (O_1295,N_24014,N_24394);
nor UO_1296 (O_1296,N_22417,N_23229);
and UO_1297 (O_1297,N_22745,N_22370);
or UO_1298 (O_1298,N_21928,N_22372);
nand UO_1299 (O_1299,N_23895,N_23811);
nand UO_1300 (O_1300,N_24775,N_23763);
and UO_1301 (O_1301,N_22205,N_24300);
nand UO_1302 (O_1302,N_24527,N_22582);
xnor UO_1303 (O_1303,N_23196,N_22321);
xor UO_1304 (O_1304,N_23615,N_22211);
or UO_1305 (O_1305,N_23736,N_22859);
and UO_1306 (O_1306,N_23967,N_22866);
or UO_1307 (O_1307,N_22680,N_23323);
nand UO_1308 (O_1308,N_22664,N_23524);
nand UO_1309 (O_1309,N_23960,N_22355);
nand UO_1310 (O_1310,N_23128,N_22428);
xnor UO_1311 (O_1311,N_22107,N_24159);
xnor UO_1312 (O_1312,N_23325,N_24815);
nor UO_1313 (O_1313,N_21919,N_24403);
nand UO_1314 (O_1314,N_24012,N_23482);
and UO_1315 (O_1315,N_22527,N_22110);
nand UO_1316 (O_1316,N_22323,N_24360);
xor UO_1317 (O_1317,N_24295,N_23265);
nand UO_1318 (O_1318,N_24261,N_24396);
xnor UO_1319 (O_1319,N_23873,N_23471);
nor UO_1320 (O_1320,N_24992,N_23462);
or UO_1321 (O_1321,N_21917,N_24337);
xnor UO_1322 (O_1322,N_24608,N_23504);
nor UO_1323 (O_1323,N_24273,N_22151);
nand UO_1324 (O_1324,N_23360,N_23440);
and UO_1325 (O_1325,N_22350,N_22443);
xnor UO_1326 (O_1326,N_23650,N_23859);
xor UO_1327 (O_1327,N_23725,N_22548);
xnor UO_1328 (O_1328,N_23148,N_22787);
nand UO_1329 (O_1329,N_22679,N_22512);
and UO_1330 (O_1330,N_22915,N_24782);
xnor UO_1331 (O_1331,N_22895,N_24545);
nand UO_1332 (O_1332,N_24354,N_24312);
and UO_1333 (O_1333,N_24915,N_24040);
nor UO_1334 (O_1334,N_22435,N_24053);
and UO_1335 (O_1335,N_22574,N_24469);
and UO_1336 (O_1336,N_22621,N_22005);
or UO_1337 (O_1337,N_24624,N_23893);
or UO_1338 (O_1338,N_22190,N_23466);
xor UO_1339 (O_1339,N_22286,N_23983);
or UO_1340 (O_1340,N_23944,N_24641);
and UO_1341 (O_1341,N_23863,N_24161);
xnor UO_1342 (O_1342,N_24007,N_24257);
xor UO_1343 (O_1343,N_22659,N_22922);
nor UO_1344 (O_1344,N_23581,N_21923);
nor UO_1345 (O_1345,N_22168,N_24458);
or UO_1346 (O_1346,N_24010,N_23320);
nand UO_1347 (O_1347,N_24866,N_22504);
and UO_1348 (O_1348,N_22156,N_24865);
nor UO_1349 (O_1349,N_23488,N_23977);
xnor UO_1350 (O_1350,N_24225,N_23658);
or UO_1351 (O_1351,N_22769,N_23730);
xnor UO_1352 (O_1352,N_24618,N_23646);
and UO_1353 (O_1353,N_24296,N_23610);
nor UO_1354 (O_1354,N_22901,N_23568);
or UO_1355 (O_1355,N_23602,N_22409);
and UO_1356 (O_1356,N_22639,N_22348);
xor UO_1357 (O_1357,N_22928,N_22614);
xnor UO_1358 (O_1358,N_22647,N_22644);
nand UO_1359 (O_1359,N_22449,N_23766);
xnor UO_1360 (O_1360,N_22764,N_22237);
xnor UO_1361 (O_1361,N_22883,N_23590);
or UO_1362 (O_1362,N_24390,N_24103);
nor UO_1363 (O_1363,N_24059,N_24967);
or UO_1364 (O_1364,N_23166,N_23737);
or UO_1365 (O_1365,N_23636,N_22701);
or UO_1366 (O_1366,N_24631,N_23803);
nor UO_1367 (O_1367,N_22016,N_23631);
or UO_1368 (O_1368,N_24232,N_22550);
or UO_1369 (O_1369,N_22616,N_23412);
nand UO_1370 (O_1370,N_24736,N_24348);
xor UO_1371 (O_1371,N_24129,N_24893);
and UO_1372 (O_1372,N_22888,N_24520);
and UO_1373 (O_1373,N_22494,N_22566);
nor UO_1374 (O_1374,N_22589,N_24199);
xnor UO_1375 (O_1375,N_24036,N_23085);
and UO_1376 (O_1376,N_23399,N_24878);
nand UO_1377 (O_1377,N_23795,N_23812);
nor UO_1378 (O_1378,N_22161,N_24488);
or UO_1379 (O_1379,N_23191,N_23534);
and UO_1380 (O_1380,N_22265,N_23778);
xnor UO_1381 (O_1381,N_24455,N_22788);
or UO_1382 (O_1382,N_23690,N_22040);
and UO_1383 (O_1383,N_23975,N_24139);
and UO_1384 (O_1384,N_23163,N_22281);
and UO_1385 (O_1385,N_24051,N_22732);
xnor UO_1386 (O_1386,N_24102,N_24697);
and UO_1387 (O_1387,N_21885,N_23500);
nor UO_1388 (O_1388,N_24728,N_24978);
nand UO_1389 (O_1389,N_22702,N_24983);
nor UO_1390 (O_1390,N_24238,N_24305);
and UO_1391 (O_1391,N_22816,N_23583);
xor UO_1392 (O_1392,N_24383,N_24591);
or UO_1393 (O_1393,N_24632,N_22564);
nand UO_1394 (O_1394,N_24837,N_23729);
and UO_1395 (O_1395,N_24804,N_23371);
or UO_1396 (O_1396,N_23915,N_23120);
or UO_1397 (O_1397,N_23637,N_23193);
or UO_1398 (O_1398,N_23937,N_24101);
or UO_1399 (O_1399,N_21880,N_22295);
and UO_1400 (O_1400,N_23258,N_22963);
and UO_1401 (O_1401,N_22704,N_21953);
xor UO_1402 (O_1402,N_23268,N_22737);
xnor UO_1403 (O_1403,N_23850,N_24044);
nor UO_1404 (O_1404,N_23436,N_23699);
or UO_1405 (O_1405,N_21999,N_22711);
nor UO_1406 (O_1406,N_22431,N_23226);
xor UO_1407 (O_1407,N_23957,N_22767);
or UO_1408 (O_1408,N_22797,N_22493);
and UO_1409 (O_1409,N_22192,N_22378);
nand UO_1410 (O_1410,N_23990,N_21908);
and UO_1411 (O_1411,N_23784,N_24939);
nand UO_1412 (O_1412,N_23980,N_23574);
nor UO_1413 (O_1413,N_22536,N_23718);
and UO_1414 (O_1414,N_22121,N_22490);
or UO_1415 (O_1415,N_24716,N_23904);
and UO_1416 (O_1416,N_21892,N_24055);
xor UO_1417 (O_1417,N_22264,N_22051);
nand UO_1418 (O_1418,N_24367,N_24699);
xor UO_1419 (O_1419,N_22754,N_24613);
nor UO_1420 (O_1420,N_23550,N_24816);
and UO_1421 (O_1421,N_22783,N_24651);
nor UO_1422 (O_1422,N_23820,N_24907);
nand UO_1423 (O_1423,N_22920,N_23264);
nand UO_1424 (O_1424,N_23813,N_22938);
or UO_1425 (O_1425,N_22204,N_21942);
or UO_1426 (O_1426,N_23337,N_23146);
and UO_1427 (O_1427,N_21944,N_22241);
or UO_1428 (O_1428,N_24001,N_21990);
or UO_1429 (O_1429,N_24797,N_23185);
nand UO_1430 (O_1430,N_22758,N_23357);
xnor UO_1431 (O_1431,N_24586,N_22090);
nor UO_1432 (O_1432,N_23930,N_23073);
xor UO_1433 (O_1433,N_24880,N_21902);
nand UO_1434 (O_1434,N_23797,N_24627);
or UO_1435 (O_1435,N_24684,N_22166);
and UO_1436 (O_1436,N_24537,N_23595);
or UO_1437 (O_1437,N_23219,N_22320);
and UO_1438 (O_1438,N_23756,N_24836);
or UO_1439 (O_1439,N_24892,N_22752);
xor UO_1440 (O_1440,N_21938,N_22726);
nand UO_1441 (O_1441,N_23044,N_24181);
nand UO_1442 (O_1442,N_23728,N_23074);
or UO_1443 (O_1443,N_22873,N_22830);
nor UO_1444 (O_1444,N_22835,N_24453);
and UO_1445 (O_1445,N_21915,N_24154);
xnor UO_1446 (O_1446,N_22103,N_24297);
nor UO_1447 (O_1447,N_23379,N_22434);
nor UO_1448 (O_1448,N_24078,N_24061);
xor UO_1449 (O_1449,N_23047,N_23443);
nor UO_1450 (O_1450,N_24368,N_22880);
or UO_1451 (O_1451,N_23752,N_22143);
nand UO_1452 (O_1452,N_23175,N_24707);
or UO_1453 (O_1453,N_23801,N_24105);
xor UO_1454 (O_1454,N_22165,N_22905);
or UO_1455 (O_1455,N_24533,N_24581);
nand UO_1456 (O_1456,N_22870,N_23556);
xor UO_1457 (O_1457,N_24747,N_24336);
xnor UO_1458 (O_1458,N_24397,N_23299);
and UO_1459 (O_1459,N_23418,N_23633);
and UO_1460 (O_1460,N_23720,N_24096);
or UO_1461 (O_1461,N_22267,N_22364);
xnor UO_1462 (O_1462,N_24422,N_24910);
nor UO_1463 (O_1463,N_22608,N_23079);
nand UO_1464 (O_1464,N_24363,N_23538);
xor UO_1465 (O_1465,N_23777,N_22703);
or UO_1466 (O_1466,N_22324,N_22303);
xnor UO_1467 (O_1467,N_23700,N_23669);
and UO_1468 (O_1468,N_22339,N_23181);
xor UO_1469 (O_1469,N_22563,N_23629);
xor UO_1470 (O_1470,N_22781,N_23244);
and UO_1471 (O_1471,N_24824,N_23411);
and UO_1472 (O_1472,N_24110,N_24894);
nor UO_1473 (O_1473,N_24028,N_22803);
nor UO_1474 (O_1474,N_23702,N_22086);
nor UO_1475 (O_1475,N_22120,N_23511);
nor UO_1476 (O_1476,N_23240,N_23922);
nor UO_1477 (O_1477,N_24448,N_23151);
nor UO_1478 (O_1478,N_23571,N_22446);
nand UO_1479 (O_1479,N_24490,N_23533);
xor UO_1480 (O_1480,N_24752,N_24666);
and UO_1481 (O_1481,N_22912,N_23919);
xor UO_1482 (O_1482,N_24412,N_23209);
and UO_1483 (O_1483,N_24116,N_23117);
nor UO_1484 (O_1484,N_22793,N_24122);
or UO_1485 (O_1485,N_24949,N_24183);
nor UO_1486 (O_1486,N_22408,N_24833);
nand UO_1487 (O_1487,N_24324,N_22235);
nor UO_1488 (O_1488,N_23058,N_24874);
nor UO_1489 (O_1489,N_24675,N_23427);
nand UO_1490 (O_1490,N_23965,N_24671);
and UO_1491 (O_1491,N_22101,N_23204);
xor UO_1492 (O_1492,N_23751,N_22056);
and UO_1493 (O_1493,N_22065,N_23924);
and UO_1494 (O_1494,N_22526,N_22669);
or UO_1495 (O_1495,N_23173,N_22213);
or UO_1496 (O_1496,N_22091,N_22685);
or UO_1497 (O_1497,N_23182,N_23389);
xor UO_1498 (O_1498,N_23261,N_24184);
xnor UO_1499 (O_1499,N_23679,N_22559);
nand UO_1500 (O_1500,N_23089,N_22763);
or UO_1501 (O_1501,N_24197,N_22480);
or UO_1502 (O_1502,N_24610,N_24908);
or UO_1503 (O_1503,N_23409,N_24062);
xnor UO_1504 (O_1504,N_23441,N_22980);
nor UO_1505 (O_1505,N_22820,N_24419);
xnor UO_1506 (O_1506,N_21936,N_21904);
or UO_1507 (O_1507,N_23496,N_24328);
nand UO_1508 (O_1508,N_22918,N_23925);
nor UO_1509 (O_1509,N_22543,N_24127);
nor UO_1510 (O_1510,N_23005,N_22972);
and UO_1511 (O_1511,N_22019,N_21935);
nor UO_1512 (O_1512,N_23632,N_22300);
and UO_1513 (O_1513,N_23437,N_23789);
nand UO_1514 (O_1514,N_22389,N_24909);
nand UO_1515 (O_1515,N_22990,N_24777);
and UO_1516 (O_1516,N_24416,N_24084);
or UO_1517 (O_1517,N_22828,N_23531);
nand UO_1518 (O_1518,N_23689,N_24921);
nor UO_1519 (O_1519,N_24264,N_24726);
xnor UO_1520 (O_1520,N_23321,N_24083);
and UO_1521 (O_1521,N_24678,N_23612);
nand UO_1522 (O_1522,N_24500,N_23510);
and UO_1523 (O_1523,N_23790,N_24965);
and UO_1524 (O_1524,N_23239,N_22796);
xnor UO_1525 (O_1525,N_23317,N_22700);
xnor UO_1526 (O_1526,N_24058,N_22043);
and UO_1527 (O_1527,N_22313,N_24464);
or UO_1528 (O_1528,N_22257,N_23620);
xnor UO_1529 (O_1529,N_22837,N_24164);
and UO_1530 (O_1530,N_23672,N_22291);
nor UO_1531 (O_1531,N_24754,N_24438);
or UO_1532 (O_1532,N_23708,N_22009);
or UO_1533 (O_1533,N_24239,N_24256);
nor UO_1534 (O_1534,N_24872,N_22037);
and UO_1535 (O_1535,N_22247,N_22104);
nand UO_1536 (O_1536,N_24667,N_23075);
nand UO_1537 (O_1537,N_23070,N_23518);
nand UO_1538 (O_1538,N_23905,N_22823);
and UO_1539 (O_1539,N_24204,N_22909);
nand UO_1540 (O_1540,N_24923,N_23945);
and UO_1541 (O_1541,N_23159,N_24344);
or UO_1542 (O_1542,N_23949,N_22426);
and UO_1543 (O_1543,N_24672,N_24433);
or UO_1544 (O_1544,N_22124,N_23758);
xnor UO_1545 (O_1545,N_23300,N_24376);
xor UO_1546 (O_1546,N_22488,N_23349);
nand UO_1547 (O_1547,N_22794,N_23596);
or UO_1548 (O_1548,N_24786,N_23661);
nand UO_1549 (O_1549,N_24219,N_24492);
nor UO_1550 (O_1550,N_23125,N_22949);
and UO_1551 (O_1551,N_24408,N_24947);
or UO_1552 (O_1552,N_23232,N_21998);
or UO_1553 (O_1553,N_22055,N_22328);
and UO_1554 (O_1554,N_23559,N_23810);
nand UO_1555 (O_1555,N_24503,N_24810);
nor UO_1556 (O_1556,N_24086,N_22079);
or UO_1557 (O_1557,N_24687,N_23907);
nor UO_1558 (O_1558,N_23671,N_22106);
nand UO_1559 (O_1559,N_22853,N_22207);
xnor UO_1560 (O_1560,N_24504,N_22298);
or UO_1561 (O_1561,N_24356,N_22154);
nand UO_1562 (O_1562,N_23076,N_22068);
or UO_1563 (O_1563,N_23961,N_24320);
nand UO_1564 (O_1564,N_22745,N_23256);
nand UO_1565 (O_1565,N_23206,N_23224);
nand UO_1566 (O_1566,N_23861,N_22544);
nor UO_1567 (O_1567,N_22309,N_23337);
nand UO_1568 (O_1568,N_23011,N_23405);
or UO_1569 (O_1569,N_23430,N_22340);
xnor UO_1570 (O_1570,N_23549,N_23158);
nor UO_1571 (O_1571,N_21905,N_22971);
nor UO_1572 (O_1572,N_23031,N_22042);
and UO_1573 (O_1573,N_22408,N_24492);
nand UO_1574 (O_1574,N_23604,N_22100);
xor UO_1575 (O_1575,N_24376,N_22006);
or UO_1576 (O_1576,N_21914,N_22293);
or UO_1577 (O_1577,N_24479,N_22848);
xnor UO_1578 (O_1578,N_24989,N_22993);
or UO_1579 (O_1579,N_21909,N_22534);
nor UO_1580 (O_1580,N_23143,N_23715);
or UO_1581 (O_1581,N_24837,N_24060);
or UO_1582 (O_1582,N_22816,N_24111);
and UO_1583 (O_1583,N_24433,N_23554);
nand UO_1584 (O_1584,N_24359,N_23410);
nor UO_1585 (O_1585,N_22488,N_22877);
and UO_1586 (O_1586,N_23358,N_22627);
or UO_1587 (O_1587,N_23491,N_21998);
and UO_1588 (O_1588,N_22681,N_23301);
xor UO_1589 (O_1589,N_22699,N_23382);
nand UO_1590 (O_1590,N_22732,N_22018);
and UO_1591 (O_1591,N_22926,N_24460);
xor UO_1592 (O_1592,N_24419,N_23416);
nor UO_1593 (O_1593,N_22176,N_24260);
or UO_1594 (O_1594,N_21934,N_23002);
nand UO_1595 (O_1595,N_24779,N_24216);
nor UO_1596 (O_1596,N_23639,N_24936);
xnor UO_1597 (O_1597,N_23869,N_22107);
nor UO_1598 (O_1598,N_23469,N_24491);
xnor UO_1599 (O_1599,N_24557,N_24837);
or UO_1600 (O_1600,N_22422,N_22135);
nand UO_1601 (O_1601,N_22365,N_22166);
nand UO_1602 (O_1602,N_22159,N_24975);
nand UO_1603 (O_1603,N_22501,N_23717);
nor UO_1604 (O_1604,N_24044,N_22614);
and UO_1605 (O_1605,N_23597,N_23113);
xor UO_1606 (O_1606,N_22364,N_22583);
and UO_1607 (O_1607,N_22996,N_24111);
or UO_1608 (O_1608,N_23717,N_24144);
xnor UO_1609 (O_1609,N_23299,N_23558);
and UO_1610 (O_1610,N_22411,N_24451);
nand UO_1611 (O_1611,N_24675,N_24107);
xnor UO_1612 (O_1612,N_24433,N_24445);
or UO_1613 (O_1613,N_22626,N_22497);
nor UO_1614 (O_1614,N_22968,N_22917);
and UO_1615 (O_1615,N_23045,N_21956);
nor UO_1616 (O_1616,N_24404,N_24205);
nor UO_1617 (O_1617,N_24804,N_24329);
nor UO_1618 (O_1618,N_22524,N_22744);
and UO_1619 (O_1619,N_24126,N_22703);
nand UO_1620 (O_1620,N_22959,N_23226);
and UO_1621 (O_1621,N_23480,N_24748);
nand UO_1622 (O_1622,N_24265,N_24701);
nand UO_1623 (O_1623,N_24708,N_22103);
nand UO_1624 (O_1624,N_24683,N_22822);
xor UO_1625 (O_1625,N_24784,N_23591);
or UO_1626 (O_1626,N_24964,N_23857);
nand UO_1627 (O_1627,N_23020,N_24739);
xnor UO_1628 (O_1628,N_22537,N_21930);
or UO_1629 (O_1629,N_24307,N_22401);
nor UO_1630 (O_1630,N_22212,N_22726);
or UO_1631 (O_1631,N_23273,N_23393);
xor UO_1632 (O_1632,N_23908,N_22499);
xnor UO_1633 (O_1633,N_24022,N_23185);
xor UO_1634 (O_1634,N_23985,N_23549);
or UO_1635 (O_1635,N_23502,N_22844);
nand UO_1636 (O_1636,N_23633,N_23087);
nand UO_1637 (O_1637,N_24721,N_22094);
and UO_1638 (O_1638,N_24151,N_23596);
or UO_1639 (O_1639,N_23578,N_22776);
nor UO_1640 (O_1640,N_22980,N_24529);
nand UO_1641 (O_1641,N_24332,N_24471);
nor UO_1642 (O_1642,N_23695,N_23370);
xnor UO_1643 (O_1643,N_24673,N_23945);
xor UO_1644 (O_1644,N_23678,N_22351);
or UO_1645 (O_1645,N_24137,N_23406);
nor UO_1646 (O_1646,N_22567,N_24200);
nor UO_1647 (O_1647,N_24464,N_22868);
nor UO_1648 (O_1648,N_22465,N_23878);
or UO_1649 (O_1649,N_23035,N_24349);
and UO_1650 (O_1650,N_23650,N_23218);
and UO_1651 (O_1651,N_24379,N_24505);
or UO_1652 (O_1652,N_22445,N_23024);
nand UO_1653 (O_1653,N_22949,N_24226);
or UO_1654 (O_1654,N_24640,N_24538);
nand UO_1655 (O_1655,N_24975,N_22264);
nor UO_1656 (O_1656,N_23272,N_24315);
and UO_1657 (O_1657,N_23666,N_23770);
nor UO_1658 (O_1658,N_23660,N_24881);
and UO_1659 (O_1659,N_22790,N_22018);
or UO_1660 (O_1660,N_24701,N_23101);
xor UO_1661 (O_1661,N_23455,N_22920);
xor UO_1662 (O_1662,N_24192,N_23942);
xor UO_1663 (O_1663,N_22096,N_24142);
and UO_1664 (O_1664,N_22289,N_23737);
nand UO_1665 (O_1665,N_24919,N_23228);
or UO_1666 (O_1666,N_22864,N_23832);
nor UO_1667 (O_1667,N_24191,N_22030);
or UO_1668 (O_1668,N_24666,N_23166);
nor UO_1669 (O_1669,N_22208,N_24183);
and UO_1670 (O_1670,N_22909,N_22652);
xnor UO_1671 (O_1671,N_24232,N_22176);
nor UO_1672 (O_1672,N_22866,N_22420);
and UO_1673 (O_1673,N_22873,N_23027);
nor UO_1674 (O_1674,N_24490,N_23661);
nand UO_1675 (O_1675,N_22752,N_23911);
xor UO_1676 (O_1676,N_24781,N_23735);
and UO_1677 (O_1677,N_22953,N_23749);
xnor UO_1678 (O_1678,N_23909,N_23269);
xor UO_1679 (O_1679,N_23645,N_22648);
nand UO_1680 (O_1680,N_24148,N_23208);
or UO_1681 (O_1681,N_22781,N_23965);
or UO_1682 (O_1682,N_23283,N_22990);
or UO_1683 (O_1683,N_22665,N_23740);
nor UO_1684 (O_1684,N_21971,N_23543);
nand UO_1685 (O_1685,N_23829,N_23975);
xor UO_1686 (O_1686,N_21982,N_23768);
xnor UO_1687 (O_1687,N_24797,N_22687);
xor UO_1688 (O_1688,N_22497,N_23633);
xnor UO_1689 (O_1689,N_23022,N_24080);
or UO_1690 (O_1690,N_24995,N_21911);
xor UO_1691 (O_1691,N_24732,N_23435);
nor UO_1692 (O_1692,N_24120,N_21887);
xor UO_1693 (O_1693,N_22520,N_24417);
and UO_1694 (O_1694,N_23054,N_24940);
nand UO_1695 (O_1695,N_23954,N_23609);
nor UO_1696 (O_1696,N_24950,N_23057);
or UO_1697 (O_1697,N_23959,N_22232);
xnor UO_1698 (O_1698,N_22159,N_23689);
nand UO_1699 (O_1699,N_22029,N_22410);
and UO_1700 (O_1700,N_22578,N_22036);
or UO_1701 (O_1701,N_24550,N_23237);
or UO_1702 (O_1702,N_24767,N_24738);
or UO_1703 (O_1703,N_22797,N_21953);
and UO_1704 (O_1704,N_23990,N_23188);
nor UO_1705 (O_1705,N_22527,N_24664);
and UO_1706 (O_1706,N_23277,N_22233);
xor UO_1707 (O_1707,N_24988,N_24646);
xnor UO_1708 (O_1708,N_23352,N_24907);
nand UO_1709 (O_1709,N_22874,N_23895);
nand UO_1710 (O_1710,N_22142,N_22893);
nor UO_1711 (O_1711,N_24290,N_23451);
and UO_1712 (O_1712,N_23004,N_24974);
and UO_1713 (O_1713,N_24523,N_22730);
xor UO_1714 (O_1714,N_23994,N_23682);
nor UO_1715 (O_1715,N_22830,N_22931);
nand UO_1716 (O_1716,N_22284,N_24096);
nand UO_1717 (O_1717,N_24405,N_22932);
nand UO_1718 (O_1718,N_22103,N_22671);
or UO_1719 (O_1719,N_23903,N_22054);
and UO_1720 (O_1720,N_23723,N_22518);
xor UO_1721 (O_1721,N_23756,N_24423);
nand UO_1722 (O_1722,N_22912,N_23370);
nor UO_1723 (O_1723,N_23882,N_23649);
nor UO_1724 (O_1724,N_22069,N_24036);
nor UO_1725 (O_1725,N_23917,N_24477);
or UO_1726 (O_1726,N_21923,N_24527);
nor UO_1727 (O_1727,N_22606,N_22260);
or UO_1728 (O_1728,N_23695,N_23067);
nand UO_1729 (O_1729,N_23822,N_24613);
xor UO_1730 (O_1730,N_23984,N_24146);
or UO_1731 (O_1731,N_22705,N_23030);
or UO_1732 (O_1732,N_24076,N_24859);
or UO_1733 (O_1733,N_23007,N_22108);
nand UO_1734 (O_1734,N_23980,N_22684);
xor UO_1735 (O_1735,N_23693,N_22379);
xor UO_1736 (O_1736,N_24896,N_22433);
or UO_1737 (O_1737,N_22842,N_24052);
and UO_1738 (O_1738,N_23187,N_24246);
xor UO_1739 (O_1739,N_23851,N_23270);
xnor UO_1740 (O_1740,N_23759,N_22169);
and UO_1741 (O_1741,N_24359,N_22616);
and UO_1742 (O_1742,N_22175,N_23786);
nor UO_1743 (O_1743,N_22694,N_22963);
or UO_1744 (O_1744,N_22862,N_24061);
nand UO_1745 (O_1745,N_22056,N_22813);
or UO_1746 (O_1746,N_23179,N_23195);
xnor UO_1747 (O_1747,N_22003,N_22027);
and UO_1748 (O_1748,N_24601,N_23963);
or UO_1749 (O_1749,N_24988,N_24311);
or UO_1750 (O_1750,N_23967,N_22722);
nand UO_1751 (O_1751,N_23421,N_22225);
nand UO_1752 (O_1752,N_23516,N_22190);
nand UO_1753 (O_1753,N_24199,N_22890);
and UO_1754 (O_1754,N_22534,N_22322);
nor UO_1755 (O_1755,N_23750,N_22594);
and UO_1756 (O_1756,N_22700,N_22832);
nand UO_1757 (O_1757,N_23085,N_23255);
nand UO_1758 (O_1758,N_23930,N_22512);
nor UO_1759 (O_1759,N_24212,N_22403);
nand UO_1760 (O_1760,N_23649,N_23062);
and UO_1761 (O_1761,N_23114,N_23842);
xor UO_1762 (O_1762,N_23113,N_23245);
nor UO_1763 (O_1763,N_21961,N_23058);
and UO_1764 (O_1764,N_24195,N_23702);
or UO_1765 (O_1765,N_22337,N_23529);
and UO_1766 (O_1766,N_24653,N_22905);
xor UO_1767 (O_1767,N_23605,N_23946);
or UO_1768 (O_1768,N_24751,N_23693);
and UO_1769 (O_1769,N_23186,N_23090);
nand UO_1770 (O_1770,N_22840,N_22488);
or UO_1771 (O_1771,N_23504,N_24655);
xor UO_1772 (O_1772,N_23067,N_24118);
xnor UO_1773 (O_1773,N_22525,N_24881);
and UO_1774 (O_1774,N_22861,N_24357);
nor UO_1775 (O_1775,N_24509,N_24482);
nand UO_1776 (O_1776,N_22261,N_22725);
nor UO_1777 (O_1777,N_22870,N_24068);
or UO_1778 (O_1778,N_24607,N_23797);
nor UO_1779 (O_1779,N_24339,N_24950);
nor UO_1780 (O_1780,N_22901,N_23649);
nor UO_1781 (O_1781,N_23589,N_22041);
or UO_1782 (O_1782,N_22288,N_21964);
and UO_1783 (O_1783,N_22024,N_24283);
and UO_1784 (O_1784,N_22580,N_22513);
xnor UO_1785 (O_1785,N_24455,N_23834);
xor UO_1786 (O_1786,N_24454,N_22783);
nand UO_1787 (O_1787,N_23859,N_22968);
nand UO_1788 (O_1788,N_22727,N_23585);
xor UO_1789 (O_1789,N_23829,N_22851);
nand UO_1790 (O_1790,N_23426,N_23751);
and UO_1791 (O_1791,N_24249,N_24756);
nor UO_1792 (O_1792,N_23333,N_23730);
or UO_1793 (O_1793,N_24993,N_22460);
nor UO_1794 (O_1794,N_22758,N_21909);
nor UO_1795 (O_1795,N_23481,N_23868);
nand UO_1796 (O_1796,N_23860,N_23596);
nand UO_1797 (O_1797,N_22840,N_22406);
nand UO_1798 (O_1798,N_21909,N_22918);
xor UO_1799 (O_1799,N_24260,N_23563);
xor UO_1800 (O_1800,N_22090,N_23124);
and UO_1801 (O_1801,N_22627,N_23514);
xor UO_1802 (O_1802,N_24228,N_22267);
xor UO_1803 (O_1803,N_22207,N_22197);
nor UO_1804 (O_1804,N_22743,N_22304);
or UO_1805 (O_1805,N_23974,N_23115);
nand UO_1806 (O_1806,N_23751,N_22978);
and UO_1807 (O_1807,N_24286,N_23312);
xor UO_1808 (O_1808,N_23936,N_24680);
xnor UO_1809 (O_1809,N_22459,N_23292);
nor UO_1810 (O_1810,N_23766,N_24029);
nand UO_1811 (O_1811,N_22021,N_24189);
or UO_1812 (O_1812,N_21979,N_22806);
nand UO_1813 (O_1813,N_23067,N_22562);
and UO_1814 (O_1814,N_22642,N_22514);
and UO_1815 (O_1815,N_23946,N_23375);
nor UO_1816 (O_1816,N_22238,N_24595);
and UO_1817 (O_1817,N_24789,N_23868);
and UO_1818 (O_1818,N_23474,N_22278);
and UO_1819 (O_1819,N_22902,N_23057);
or UO_1820 (O_1820,N_22707,N_22891);
nand UO_1821 (O_1821,N_24754,N_22471);
or UO_1822 (O_1822,N_22936,N_22526);
or UO_1823 (O_1823,N_23143,N_24223);
and UO_1824 (O_1824,N_24098,N_23621);
and UO_1825 (O_1825,N_24721,N_22748);
xor UO_1826 (O_1826,N_24012,N_23222);
and UO_1827 (O_1827,N_22406,N_23646);
or UO_1828 (O_1828,N_23788,N_24765);
nand UO_1829 (O_1829,N_23805,N_24691);
or UO_1830 (O_1830,N_23823,N_24747);
and UO_1831 (O_1831,N_23512,N_23218);
xor UO_1832 (O_1832,N_23851,N_23940);
and UO_1833 (O_1833,N_23046,N_23349);
or UO_1834 (O_1834,N_24164,N_23734);
or UO_1835 (O_1835,N_23414,N_23943);
nand UO_1836 (O_1836,N_22727,N_23856);
xnor UO_1837 (O_1837,N_24571,N_24187);
xnor UO_1838 (O_1838,N_22172,N_22269);
and UO_1839 (O_1839,N_23119,N_22122);
or UO_1840 (O_1840,N_24303,N_23419);
nor UO_1841 (O_1841,N_24510,N_22475);
xor UO_1842 (O_1842,N_22685,N_22154);
nand UO_1843 (O_1843,N_22870,N_22358);
xor UO_1844 (O_1844,N_22800,N_22937);
and UO_1845 (O_1845,N_22007,N_23366);
or UO_1846 (O_1846,N_24162,N_22766);
or UO_1847 (O_1847,N_22974,N_24592);
nand UO_1848 (O_1848,N_23681,N_23337);
nand UO_1849 (O_1849,N_23000,N_24132);
or UO_1850 (O_1850,N_23917,N_24377);
nor UO_1851 (O_1851,N_24729,N_22214);
and UO_1852 (O_1852,N_22339,N_24911);
nand UO_1853 (O_1853,N_22231,N_23246);
xor UO_1854 (O_1854,N_24009,N_24649);
and UO_1855 (O_1855,N_22801,N_23740);
nor UO_1856 (O_1856,N_24648,N_22978);
nor UO_1857 (O_1857,N_23167,N_23246);
xnor UO_1858 (O_1858,N_23541,N_23315);
nor UO_1859 (O_1859,N_24627,N_23121);
nand UO_1860 (O_1860,N_23149,N_23453);
nor UO_1861 (O_1861,N_22303,N_23567);
nand UO_1862 (O_1862,N_22163,N_23388);
xor UO_1863 (O_1863,N_22666,N_24443);
nand UO_1864 (O_1864,N_24894,N_24225);
nand UO_1865 (O_1865,N_24940,N_23373);
and UO_1866 (O_1866,N_22723,N_23146);
or UO_1867 (O_1867,N_22390,N_22140);
nand UO_1868 (O_1868,N_24744,N_24691);
nor UO_1869 (O_1869,N_24627,N_22696);
nand UO_1870 (O_1870,N_24367,N_24916);
nand UO_1871 (O_1871,N_24839,N_22726);
and UO_1872 (O_1872,N_23842,N_22518);
nor UO_1873 (O_1873,N_23355,N_22933);
nor UO_1874 (O_1874,N_22084,N_21999);
nand UO_1875 (O_1875,N_21961,N_24913);
nor UO_1876 (O_1876,N_22128,N_21928);
nor UO_1877 (O_1877,N_23648,N_22619);
or UO_1878 (O_1878,N_23717,N_24476);
or UO_1879 (O_1879,N_22728,N_22898);
nor UO_1880 (O_1880,N_23626,N_24571);
nor UO_1881 (O_1881,N_24579,N_24103);
xor UO_1882 (O_1882,N_23176,N_24637);
or UO_1883 (O_1883,N_24912,N_23768);
xnor UO_1884 (O_1884,N_23282,N_22242);
or UO_1885 (O_1885,N_22907,N_22844);
xnor UO_1886 (O_1886,N_23023,N_22264);
nand UO_1887 (O_1887,N_24610,N_24557);
xnor UO_1888 (O_1888,N_24066,N_22839);
and UO_1889 (O_1889,N_24773,N_22665);
xnor UO_1890 (O_1890,N_22486,N_22871);
and UO_1891 (O_1891,N_22672,N_24111);
nand UO_1892 (O_1892,N_23439,N_23558);
nand UO_1893 (O_1893,N_23185,N_22235);
nor UO_1894 (O_1894,N_22107,N_22034);
xor UO_1895 (O_1895,N_24994,N_23781);
and UO_1896 (O_1896,N_23050,N_23150);
nor UO_1897 (O_1897,N_24039,N_23935);
and UO_1898 (O_1898,N_22068,N_22655);
nor UO_1899 (O_1899,N_24288,N_22514);
xnor UO_1900 (O_1900,N_24794,N_22271);
and UO_1901 (O_1901,N_22918,N_23038);
and UO_1902 (O_1902,N_22465,N_23430);
xnor UO_1903 (O_1903,N_22656,N_23762);
nor UO_1904 (O_1904,N_22903,N_22568);
or UO_1905 (O_1905,N_24789,N_22313);
xor UO_1906 (O_1906,N_22858,N_24061);
nor UO_1907 (O_1907,N_23002,N_22308);
and UO_1908 (O_1908,N_23575,N_22041);
nand UO_1909 (O_1909,N_23154,N_21875);
and UO_1910 (O_1910,N_23241,N_24956);
and UO_1911 (O_1911,N_23860,N_23743);
or UO_1912 (O_1912,N_24868,N_23313);
nor UO_1913 (O_1913,N_22418,N_23448);
nor UO_1914 (O_1914,N_23918,N_22656);
nor UO_1915 (O_1915,N_23503,N_23980);
and UO_1916 (O_1916,N_22255,N_23319);
nor UO_1917 (O_1917,N_23699,N_23833);
xnor UO_1918 (O_1918,N_23827,N_23159);
nor UO_1919 (O_1919,N_22533,N_24405);
nor UO_1920 (O_1920,N_24447,N_22287);
xor UO_1921 (O_1921,N_23040,N_24771);
xnor UO_1922 (O_1922,N_23930,N_23533);
nand UO_1923 (O_1923,N_21976,N_24670);
nor UO_1924 (O_1924,N_22795,N_23129);
or UO_1925 (O_1925,N_23455,N_24594);
nand UO_1926 (O_1926,N_23160,N_23288);
nor UO_1927 (O_1927,N_22681,N_22010);
nor UO_1928 (O_1928,N_23803,N_24024);
or UO_1929 (O_1929,N_24280,N_22128);
xnor UO_1930 (O_1930,N_22135,N_22753);
and UO_1931 (O_1931,N_22748,N_23957);
or UO_1932 (O_1932,N_24311,N_24173);
nand UO_1933 (O_1933,N_23924,N_23329);
nor UO_1934 (O_1934,N_22059,N_22964);
and UO_1935 (O_1935,N_22712,N_22322);
and UO_1936 (O_1936,N_23666,N_23415);
and UO_1937 (O_1937,N_24603,N_23890);
xor UO_1938 (O_1938,N_23190,N_23331);
or UO_1939 (O_1939,N_22454,N_22861);
xor UO_1940 (O_1940,N_23333,N_23146);
nor UO_1941 (O_1941,N_24017,N_22535);
xnor UO_1942 (O_1942,N_22412,N_21905);
and UO_1943 (O_1943,N_23462,N_22242);
and UO_1944 (O_1944,N_23206,N_24135);
or UO_1945 (O_1945,N_22553,N_22376);
nand UO_1946 (O_1946,N_23186,N_23612);
xor UO_1947 (O_1947,N_22089,N_23148);
and UO_1948 (O_1948,N_21919,N_23832);
and UO_1949 (O_1949,N_23070,N_22013);
and UO_1950 (O_1950,N_24585,N_23838);
or UO_1951 (O_1951,N_22822,N_24570);
or UO_1952 (O_1952,N_22696,N_24018);
nor UO_1953 (O_1953,N_22610,N_22377);
or UO_1954 (O_1954,N_23219,N_22200);
xor UO_1955 (O_1955,N_24251,N_22099);
nor UO_1956 (O_1956,N_22822,N_24949);
and UO_1957 (O_1957,N_22326,N_24318);
nand UO_1958 (O_1958,N_22990,N_22826);
or UO_1959 (O_1959,N_24677,N_24313);
and UO_1960 (O_1960,N_24269,N_23591);
xor UO_1961 (O_1961,N_23382,N_22898);
nor UO_1962 (O_1962,N_21888,N_24743);
xnor UO_1963 (O_1963,N_22649,N_24741);
or UO_1964 (O_1964,N_22325,N_24684);
xor UO_1965 (O_1965,N_22094,N_22256);
nor UO_1966 (O_1966,N_23091,N_22945);
xor UO_1967 (O_1967,N_23807,N_24616);
xor UO_1968 (O_1968,N_22102,N_24945);
nand UO_1969 (O_1969,N_23088,N_21918);
nor UO_1970 (O_1970,N_24487,N_24505);
nor UO_1971 (O_1971,N_22134,N_24726);
nand UO_1972 (O_1972,N_23387,N_23571);
and UO_1973 (O_1973,N_22263,N_24439);
nor UO_1974 (O_1974,N_22679,N_23425);
nor UO_1975 (O_1975,N_22925,N_22334);
or UO_1976 (O_1976,N_22831,N_23105);
nand UO_1977 (O_1977,N_24029,N_24756);
nand UO_1978 (O_1978,N_24032,N_23686);
nand UO_1979 (O_1979,N_21901,N_22604);
xnor UO_1980 (O_1980,N_23556,N_23703);
and UO_1981 (O_1981,N_22272,N_24079);
and UO_1982 (O_1982,N_22336,N_23869);
nor UO_1983 (O_1983,N_22767,N_22686);
or UO_1984 (O_1984,N_23664,N_24481);
nor UO_1985 (O_1985,N_23859,N_24716);
nor UO_1986 (O_1986,N_23218,N_22659);
xnor UO_1987 (O_1987,N_24531,N_24353);
xnor UO_1988 (O_1988,N_24930,N_24369);
nand UO_1989 (O_1989,N_22188,N_22002);
and UO_1990 (O_1990,N_22334,N_23026);
xor UO_1991 (O_1991,N_24660,N_24366);
xnor UO_1992 (O_1992,N_24981,N_23018);
nand UO_1993 (O_1993,N_24416,N_22292);
nor UO_1994 (O_1994,N_24256,N_24627);
or UO_1995 (O_1995,N_22259,N_22019);
nor UO_1996 (O_1996,N_24701,N_24256);
xnor UO_1997 (O_1997,N_22071,N_22463);
nor UO_1998 (O_1998,N_24357,N_24051);
nor UO_1999 (O_1999,N_22152,N_22555);
and UO_2000 (O_2000,N_24887,N_22673);
nand UO_2001 (O_2001,N_24364,N_23187);
nor UO_2002 (O_2002,N_24556,N_23070);
nand UO_2003 (O_2003,N_22879,N_23350);
xnor UO_2004 (O_2004,N_22687,N_24093);
nand UO_2005 (O_2005,N_24424,N_22243);
nand UO_2006 (O_2006,N_24416,N_23390);
nor UO_2007 (O_2007,N_22988,N_23366);
and UO_2008 (O_2008,N_24943,N_23522);
or UO_2009 (O_2009,N_23728,N_22302);
nor UO_2010 (O_2010,N_22607,N_24876);
xor UO_2011 (O_2011,N_24022,N_24850);
or UO_2012 (O_2012,N_22198,N_24902);
xnor UO_2013 (O_2013,N_23324,N_24116);
xnor UO_2014 (O_2014,N_24651,N_21912);
nor UO_2015 (O_2015,N_22474,N_24571);
nand UO_2016 (O_2016,N_24160,N_23267);
or UO_2017 (O_2017,N_23165,N_24721);
and UO_2018 (O_2018,N_24987,N_23918);
nand UO_2019 (O_2019,N_23957,N_23563);
xor UO_2020 (O_2020,N_24490,N_24626);
or UO_2021 (O_2021,N_23889,N_23896);
or UO_2022 (O_2022,N_23896,N_22488);
and UO_2023 (O_2023,N_23618,N_23435);
nor UO_2024 (O_2024,N_23493,N_23421);
nand UO_2025 (O_2025,N_22356,N_23081);
or UO_2026 (O_2026,N_22356,N_24044);
nand UO_2027 (O_2027,N_24484,N_23824);
nor UO_2028 (O_2028,N_22193,N_24198);
and UO_2029 (O_2029,N_24804,N_23210);
xor UO_2030 (O_2030,N_23660,N_24356);
or UO_2031 (O_2031,N_24365,N_24391);
nand UO_2032 (O_2032,N_23846,N_23071);
and UO_2033 (O_2033,N_24810,N_21972);
xnor UO_2034 (O_2034,N_24158,N_22370);
or UO_2035 (O_2035,N_23728,N_21924);
nand UO_2036 (O_2036,N_22374,N_24328);
nand UO_2037 (O_2037,N_21917,N_22149);
nand UO_2038 (O_2038,N_24416,N_22548);
nand UO_2039 (O_2039,N_24040,N_22766);
nand UO_2040 (O_2040,N_22440,N_22514);
or UO_2041 (O_2041,N_22440,N_22300);
nand UO_2042 (O_2042,N_24800,N_22570);
nor UO_2043 (O_2043,N_21960,N_23642);
xnor UO_2044 (O_2044,N_24981,N_24712);
and UO_2045 (O_2045,N_24441,N_23875);
nand UO_2046 (O_2046,N_24137,N_22988);
nand UO_2047 (O_2047,N_24557,N_22596);
nand UO_2048 (O_2048,N_24542,N_24105);
or UO_2049 (O_2049,N_21977,N_23939);
and UO_2050 (O_2050,N_24910,N_23239);
and UO_2051 (O_2051,N_24917,N_23406);
nand UO_2052 (O_2052,N_21935,N_23446);
and UO_2053 (O_2053,N_24132,N_23133);
nor UO_2054 (O_2054,N_23077,N_24056);
xnor UO_2055 (O_2055,N_23773,N_22990);
nand UO_2056 (O_2056,N_24677,N_24033);
xor UO_2057 (O_2057,N_23065,N_22492);
or UO_2058 (O_2058,N_24709,N_22720);
and UO_2059 (O_2059,N_23973,N_22247);
xor UO_2060 (O_2060,N_23612,N_24679);
and UO_2061 (O_2061,N_23576,N_24642);
xnor UO_2062 (O_2062,N_24884,N_24389);
and UO_2063 (O_2063,N_22283,N_22657);
xor UO_2064 (O_2064,N_22357,N_24845);
and UO_2065 (O_2065,N_24597,N_24855);
nor UO_2066 (O_2066,N_24028,N_24705);
nor UO_2067 (O_2067,N_23102,N_24394);
xnor UO_2068 (O_2068,N_23231,N_24414);
nand UO_2069 (O_2069,N_23665,N_23516);
and UO_2070 (O_2070,N_22790,N_23315);
xor UO_2071 (O_2071,N_23395,N_23012);
nor UO_2072 (O_2072,N_23815,N_22798);
nand UO_2073 (O_2073,N_23627,N_24119);
or UO_2074 (O_2074,N_24300,N_24390);
nor UO_2075 (O_2075,N_24380,N_23653);
xor UO_2076 (O_2076,N_23443,N_21970);
nor UO_2077 (O_2077,N_22310,N_22659);
xnor UO_2078 (O_2078,N_22873,N_24191);
nor UO_2079 (O_2079,N_23975,N_22251);
nand UO_2080 (O_2080,N_24220,N_22206);
or UO_2081 (O_2081,N_22705,N_22012);
nand UO_2082 (O_2082,N_23126,N_24591);
nand UO_2083 (O_2083,N_22566,N_22304);
xor UO_2084 (O_2084,N_24483,N_24591);
nor UO_2085 (O_2085,N_22700,N_24469);
xnor UO_2086 (O_2086,N_23722,N_24190);
xor UO_2087 (O_2087,N_22107,N_22644);
nor UO_2088 (O_2088,N_22180,N_22709);
or UO_2089 (O_2089,N_22413,N_23892);
nand UO_2090 (O_2090,N_23465,N_24565);
and UO_2091 (O_2091,N_22458,N_23759);
xor UO_2092 (O_2092,N_24958,N_21933);
nand UO_2093 (O_2093,N_24076,N_22107);
and UO_2094 (O_2094,N_24052,N_24719);
nor UO_2095 (O_2095,N_23200,N_24787);
or UO_2096 (O_2096,N_23675,N_23203);
or UO_2097 (O_2097,N_24234,N_23962);
and UO_2098 (O_2098,N_22305,N_23591);
or UO_2099 (O_2099,N_22537,N_23034);
xor UO_2100 (O_2100,N_22608,N_22132);
and UO_2101 (O_2101,N_23258,N_24070);
or UO_2102 (O_2102,N_24105,N_22380);
nand UO_2103 (O_2103,N_23029,N_23843);
and UO_2104 (O_2104,N_23075,N_22897);
nand UO_2105 (O_2105,N_22282,N_24142);
and UO_2106 (O_2106,N_24726,N_23183);
xnor UO_2107 (O_2107,N_24244,N_23320);
nor UO_2108 (O_2108,N_22398,N_24901);
or UO_2109 (O_2109,N_23708,N_24358);
or UO_2110 (O_2110,N_22108,N_24600);
nor UO_2111 (O_2111,N_24013,N_22387);
xnor UO_2112 (O_2112,N_23391,N_22816);
nor UO_2113 (O_2113,N_24942,N_22481);
nor UO_2114 (O_2114,N_24442,N_23257);
or UO_2115 (O_2115,N_22657,N_24108);
nand UO_2116 (O_2116,N_24746,N_23633);
or UO_2117 (O_2117,N_24894,N_23296);
xor UO_2118 (O_2118,N_23616,N_24137);
or UO_2119 (O_2119,N_23176,N_24054);
nand UO_2120 (O_2120,N_23863,N_24545);
xnor UO_2121 (O_2121,N_23220,N_23283);
nand UO_2122 (O_2122,N_22956,N_24011);
nor UO_2123 (O_2123,N_23396,N_23072);
nand UO_2124 (O_2124,N_24641,N_22619);
and UO_2125 (O_2125,N_22976,N_24761);
or UO_2126 (O_2126,N_22899,N_22084);
or UO_2127 (O_2127,N_21938,N_22990);
or UO_2128 (O_2128,N_24213,N_24542);
and UO_2129 (O_2129,N_23204,N_23171);
nand UO_2130 (O_2130,N_22085,N_23360);
nand UO_2131 (O_2131,N_22271,N_22728);
nor UO_2132 (O_2132,N_23977,N_23426);
nand UO_2133 (O_2133,N_23480,N_23705);
nand UO_2134 (O_2134,N_22981,N_24143);
nor UO_2135 (O_2135,N_23377,N_22601);
nor UO_2136 (O_2136,N_22290,N_24365);
and UO_2137 (O_2137,N_23884,N_22966);
nand UO_2138 (O_2138,N_22731,N_22713);
xor UO_2139 (O_2139,N_23333,N_23064);
nand UO_2140 (O_2140,N_24265,N_23564);
nor UO_2141 (O_2141,N_23409,N_24026);
or UO_2142 (O_2142,N_22601,N_23976);
xnor UO_2143 (O_2143,N_23551,N_24188);
or UO_2144 (O_2144,N_24002,N_21953);
nand UO_2145 (O_2145,N_24103,N_24491);
xor UO_2146 (O_2146,N_24346,N_24785);
nor UO_2147 (O_2147,N_22483,N_23083);
xor UO_2148 (O_2148,N_23213,N_22789);
xor UO_2149 (O_2149,N_23770,N_22126);
nand UO_2150 (O_2150,N_22437,N_24277);
and UO_2151 (O_2151,N_22018,N_24854);
or UO_2152 (O_2152,N_23558,N_24927);
or UO_2153 (O_2153,N_24501,N_21910);
xnor UO_2154 (O_2154,N_22548,N_23898);
and UO_2155 (O_2155,N_22748,N_23448);
nor UO_2156 (O_2156,N_22781,N_24040);
nand UO_2157 (O_2157,N_24560,N_24884);
nand UO_2158 (O_2158,N_22685,N_23425);
nor UO_2159 (O_2159,N_23592,N_24308);
and UO_2160 (O_2160,N_22454,N_22593);
or UO_2161 (O_2161,N_22592,N_23348);
or UO_2162 (O_2162,N_22981,N_22408);
xnor UO_2163 (O_2163,N_22956,N_24704);
and UO_2164 (O_2164,N_24594,N_22492);
nand UO_2165 (O_2165,N_24590,N_23813);
xor UO_2166 (O_2166,N_24019,N_24167);
and UO_2167 (O_2167,N_24099,N_23672);
nand UO_2168 (O_2168,N_24239,N_22730);
nor UO_2169 (O_2169,N_22026,N_24278);
nor UO_2170 (O_2170,N_23085,N_24538);
xor UO_2171 (O_2171,N_24126,N_22847);
xor UO_2172 (O_2172,N_22404,N_23483);
xnor UO_2173 (O_2173,N_23406,N_22096);
xnor UO_2174 (O_2174,N_24475,N_23337);
xor UO_2175 (O_2175,N_23978,N_22807);
nand UO_2176 (O_2176,N_22646,N_24262);
xor UO_2177 (O_2177,N_23774,N_22892);
and UO_2178 (O_2178,N_23033,N_23302);
nor UO_2179 (O_2179,N_22584,N_23024);
or UO_2180 (O_2180,N_22381,N_22309);
or UO_2181 (O_2181,N_24973,N_24335);
xor UO_2182 (O_2182,N_23925,N_24259);
nand UO_2183 (O_2183,N_24719,N_22094);
or UO_2184 (O_2184,N_22431,N_23770);
xor UO_2185 (O_2185,N_24374,N_23541);
and UO_2186 (O_2186,N_22552,N_24333);
xor UO_2187 (O_2187,N_22223,N_24717);
xor UO_2188 (O_2188,N_22613,N_24523);
and UO_2189 (O_2189,N_23925,N_22682);
nor UO_2190 (O_2190,N_22171,N_22991);
and UO_2191 (O_2191,N_24940,N_23736);
nor UO_2192 (O_2192,N_24553,N_21934);
nand UO_2193 (O_2193,N_23675,N_23578);
xor UO_2194 (O_2194,N_24812,N_22772);
nor UO_2195 (O_2195,N_22242,N_22493);
nand UO_2196 (O_2196,N_24748,N_24730);
nor UO_2197 (O_2197,N_21892,N_22629);
nor UO_2198 (O_2198,N_23308,N_24768);
xnor UO_2199 (O_2199,N_22437,N_24758);
or UO_2200 (O_2200,N_24900,N_22990);
nor UO_2201 (O_2201,N_22207,N_24436);
nand UO_2202 (O_2202,N_22654,N_23657);
xnor UO_2203 (O_2203,N_24340,N_22741);
nand UO_2204 (O_2204,N_24124,N_23014);
and UO_2205 (O_2205,N_22457,N_24720);
nand UO_2206 (O_2206,N_24020,N_22884);
or UO_2207 (O_2207,N_22390,N_24371);
xor UO_2208 (O_2208,N_23975,N_24191);
nor UO_2209 (O_2209,N_24898,N_23213);
nor UO_2210 (O_2210,N_24039,N_22706);
or UO_2211 (O_2211,N_22867,N_23378);
nor UO_2212 (O_2212,N_23805,N_22667);
and UO_2213 (O_2213,N_22967,N_24853);
nor UO_2214 (O_2214,N_22989,N_24907);
and UO_2215 (O_2215,N_23820,N_24113);
and UO_2216 (O_2216,N_23206,N_22723);
nand UO_2217 (O_2217,N_23600,N_22411);
or UO_2218 (O_2218,N_23576,N_24735);
xor UO_2219 (O_2219,N_23020,N_23952);
or UO_2220 (O_2220,N_22628,N_24604);
nor UO_2221 (O_2221,N_22624,N_23191);
nand UO_2222 (O_2222,N_24143,N_23880);
xnor UO_2223 (O_2223,N_23772,N_23387);
nor UO_2224 (O_2224,N_24234,N_24215);
xnor UO_2225 (O_2225,N_24370,N_23099);
or UO_2226 (O_2226,N_24424,N_23949);
nor UO_2227 (O_2227,N_24876,N_23257);
or UO_2228 (O_2228,N_22302,N_22199);
and UO_2229 (O_2229,N_22188,N_22303);
or UO_2230 (O_2230,N_21955,N_22894);
nor UO_2231 (O_2231,N_23334,N_24756);
xnor UO_2232 (O_2232,N_24065,N_24003);
or UO_2233 (O_2233,N_23810,N_23824);
nor UO_2234 (O_2234,N_24171,N_23877);
nor UO_2235 (O_2235,N_24886,N_24020);
nand UO_2236 (O_2236,N_24189,N_22753);
and UO_2237 (O_2237,N_24898,N_23474);
nor UO_2238 (O_2238,N_22191,N_22991);
nor UO_2239 (O_2239,N_22972,N_22391);
nand UO_2240 (O_2240,N_23846,N_22409);
nand UO_2241 (O_2241,N_24028,N_22249);
and UO_2242 (O_2242,N_23484,N_23961);
or UO_2243 (O_2243,N_23755,N_23610);
xor UO_2244 (O_2244,N_23370,N_23292);
xnor UO_2245 (O_2245,N_24353,N_22148);
nand UO_2246 (O_2246,N_23186,N_23413);
xnor UO_2247 (O_2247,N_23586,N_23374);
nor UO_2248 (O_2248,N_21901,N_22978);
nand UO_2249 (O_2249,N_23921,N_23844);
and UO_2250 (O_2250,N_22970,N_22860);
xor UO_2251 (O_2251,N_24854,N_24219);
xor UO_2252 (O_2252,N_22913,N_23345);
xor UO_2253 (O_2253,N_23463,N_23709);
nor UO_2254 (O_2254,N_23150,N_24342);
nor UO_2255 (O_2255,N_23965,N_24294);
xor UO_2256 (O_2256,N_24162,N_23200);
nand UO_2257 (O_2257,N_23484,N_23653);
nand UO_2258 (O_2258,N_24892,N_22026);
nand UO_2259 (O_2259,N_24835,N_22769);
xor UO_2260 (O_2260,N_24505,N_24423);
or UO_2261 (O_2261,N_24767,N_24451);
xor UO_2262 (O_2262,N_22153,N_22832);
and UO_2263 (O_2263,N_24809,N_22135);
nand UO_2264 (O_2264,N_24689,N_24864);
and UO_2265 (O_2265,N_24374,N_24165);
nand UO_2266 (O_2266,N_23933,N_22712);
nor UO_2267 (O_2267,N_22426,N_23229);
and UO_2268 (O_2268,N_22321,N_24145);
nor UO_2269 (O_2269,N_24014,N_23217);
nor UO_2270 (O_2270,N_22933,N_22908);
nand UO_2271 (O_2271,N_22942,N_22882);
nand UO_2272 (O_2272,N_23001,N_23613);
nor UO_2273 (O_2273,N_22050,N_23233);
nand UO_2274 (O_2274,N_24951,N_23503);
xor UO_2275 (O_2275,N_23761,N_24180);
nand UO_2276 (O_2276,N_21953,N_24500);
or UO_2277 (O_2277,N_22751,N_24215);
xnor UO_2278 (O_2278,N_23340,N_22893);
xnor UO_2279 (O_2279,N_22443,N_21916);
nand UO_2280 (O_2280,N_24255,N_22231);
and UO_2281 (O_2281,N_24244,N_22287);
nand UO_2282 (O_2282,N_24066,N_24177);
nand UO_2283 (O_2283,N_22038,N_21978);
xnor UO_2284 (O_2284,N_24203,N_23913);
xnor UO_2285 (O_2285,N_24549,N_24249);
xnor UO_2286 (O_2286,N_22246,N_22181);
or UO_2287 (O_2287,N_22636,N_23811);
nand UO_2288 (O_2288,N_22347,N_24949);
xor UO_2289 (O_2289,N_23793,N_23821);
nor UO_2290 (O_2290,N_22781,N_24266);
and UO_2291 (O_2291,N_24275,N_21989);
xnor UO_2292 (O_2292,N_22483,N_23442);
nor UO_2293 (O_2293,N_22448,N_24637);
nor UO_2294 (O_2294,N_24527,N_24594);
or UO_2295 (O_2295,N_24426,N_24893);
or UO_2296 (O_2296,N_22383,N_22157);
or UO_2297 (O_2297,N_24387,N_24565);
nor UO_2298 (O_2298,N_23714,N_23511);
and UO_2299 (O_2299,N_22854,N_22004);
xor UO_2300 (O_2300,N_23647,N_22102);
and UO_2301 (O_2301,N_24702,N_22634);
or UO_2302 (O_2302,N_24654,N_23600);
xor UO_2303 (O_2303,N_23203,N_23796);
or UO_2304 (O_2304,N_24757,N_22523);
and UO_2305 (O_2305,N_24927,N_24594);
xor UO_2306 (O_2306,N_23668,N_23156);
and UO_2307 (O_2307,N_24675,N_23884);
or UO_2308 (O_2308,N_23888,N_24074);
or UO_2309 (O_2309,N_24182,N_24803);
or UO_2310 (O_2310,N_24022,N_24991);
nand UO_2311 (O_2311,N_24208,N_23302);
and UO_2312 (O_2312,N_23470,N_22829);
nor UO_2313 (O_2313,N_22374,N_23125);
xnor UO_2314 (O_2314,N_24938,N_24523);
nor UO_2315 (O_2315,N_24417,N_24178);
xor UO_2316 (O_2316,N_23291,N_23601);
and UO_2317 (O_2317,N_22393,N_24865);
nand UO_2318 (O_2318,N_23171,N_24879);
nor UO_2319 (O_2319,N_21904,N_24369);
and UO_2320 (O_2320,N_24708,N_23257);
and UO_2321 (O_2321,N_23295,N_23539);
or UO_2322 (O_2322,N_24733,N_24473);
or UO_2323 (O_2323,N_23256,N_24809);
nor UO_2324 (O_2324,N_23606,N_23613);
nor UO_2325 (O_2325,N_24501,N_22917);
nand UO_2326 (O_2326,N_23707,N_24034);
xor UO_2327 (O_2327,N_23825,N_23584);
or UO_2328 (O_2328,N_22689,N_23657);
nor UO_2329 (O_2329,N_24132,N_24750);
nand UO_2330 (O_2330,N_24061,N_23165);
nand UO_2331 (O_2331,N_24832,N_23026);
and UO_2332 (O_2332,N_22633,N_23965);
nand UO_2333 (O_2333,N_22432,N_22654);
nor UO_2334 (O_2334,N_24986,N_24662);
and UO_2335 (O_2335,N_24658,N_24151);
nand UO_2336 (O_2336,N_22648,N_23423);
nor UO_2337 (O_2337,N_22248,N_23354);
xnor UO_2338 (O_2338,N_23174,N_22698);
nor UO_2339 (O_2339,N_23818,N_24284);
nand UO_2340 (O_2340,N_24095,N_23217);
xor UO_2341 (O_2341,N_23973,N_24254);
and UO_2342 (O_2342,N_24516,N_22335);
nor UO_2343 (O_2343,N_24390,N_24514);
nand UO_2344 (O_2344,N_23876,N_22203);
nor UO_2345 (O_2345,N_24102,N_23497);
and UO_2346 (O_2346,N_22135,N_22768);
and UO_2347 (O_2347,N_22725,N_24436);
nand UO_2348 (O_2348,N_22107,N_22193);
nand UO_2349 (O_2349,N_24758,N_21999);
xor UO_2350 (O_2350,N_23166,N_23720);
nand UO_2351 (O_2351,N_24876,N_23663);
xor UO_2352 (O_2352,N_24415,N_22004);
nand UO_2353 (O_2353,N_22425,N_22175);
nor UO_2354 (O_2354,N_24626,N_23268);
or UO_2355 (O_2355,N_22554,N_21965);
nand UO_2356 (O_2356,N_23793,N_24586);
xor UO_2357 (O_2357,N_24083,N_24074);
or UO_2358 (O_2358,N_24481,N_24242);
nand UO_2359 (O_2359,N_24455,N_24442);
nor UO_2360 (O_2360,N_23741,N_24315);
nor UO_2361 (O_2361,N_24961,N_23251);
xor UO_2362 (O_2362,N_22648,N_24380);
or UO_2363 (O_2363,N_24181,N_23067);
nor UO_2364 (O_2364,N_24793,N_22866);
nor UO_2365 (O_2365,N_22801,N_23499);
or UO_2366 (O_2366,N_22566,N_24155);
nor UO_2367 (O_2367,N_23293,N_23173);
xor UO_2368 (O_2368,N_22021,N_22518);
and UO_2369 (O_2369,N_24160,N_24940);
or UO_2370 (O_2370,N_22102,N_21963);
or UO_2371 (O_2371,N_24468,N_23622);
xnor UO_2372 (O_2372,N_23347,N_22262);
nor UO_2373 (O_2373,N_23225,N_22482);
or UO_2374 (O_2374,N_22623,N_23410);
or UO_2375 (O_2375,N_21993,N_23870);
and UO_2376 (O_2376,N_21989,N_22332);
and UO_2377 (O_2377,N_23741,N_22508);
or UO_2378 (O_2378,N_22480,N_22548);
xor UO_2379 (O_2379,N_24824,N_23864);
nand UO_2380 (O_2380,N_22663,N_22097);
nor UO_2381 (O_2381,N_24734,N_24598);
nor UO_2382 (O_2382,N_24754,N_21946);
or UO_2383 (O_2383,N_22610,N_23751);
and UO_2384 (O_2384,N_23745,N_22576);
nand UO_2385 (O_2385,N_22298,N_22152);
and UO_2386 (O_2386,N_23266,N_23577);
nand UO_2387 (O_2387,N_23321,N_21968);
and UO_2388 (O_2388,N_23238,N_24327);
xnor UO_2389 (O_2389,N_23973,N_22811);
and UO_2390 (O_2390,N_24032,N_22162);
xor UO_2391 (O_2391,N_23596,N_22773);
or UO_2392 (O_2392,N_23697,N_22175);
nand UO_2393 (O_2393,N_24289,N_24217);
or UO_2394 (O_2394,N_24707,N_24133);
xor UO_2395 (O_2395,N_23991,N_24103);
or UO_2396 (O_2396,N_22298,N_22710);
and UO_2397 (O_2397,N_23162,N_23998);
xnor UO_2398 (O_2398,N_22668,N_23241);
or UO_2399 (O_2399,N_22268,N_22416);
and UO_2400 (O_2400,N_22136,N_22367);
and UO_2401 (O_2401,N_22820,N_22381);
nand UO_2402 (O_2402,N_24106,N_24720);
or UO_2403 (O_2403,N_24655,N_23438);
nor UO_2404 (O_2404,N_24354,N_23986);
and UO_2405 (O_2405,N_24228,N_23891);
or UO_2406 (O_2406,N_23434,N_22678);
nor UO_2407 (O_2407,N_24153,N_22795);
nand UO_2408 (O_2408,N_22344,N_24659);
and UO_2409 (O_2409,N_21927,N_23827);
nand UO_2410 (O_2410,N_22219,N_22676);
nor UO_2411 (O_2411,N_24496,N_23547);
and UO_2412 (O_2412,N_22639,N_23366);
xor UO_2413 (O_2413,N_24480,N_24758);
or UO_2414 (O_2414,N_24133,N_22718);
or UO_2415 (O_2415,N_22247,N_22800);
or UO_2416 (O_2416,N_24365,N_22058);
xor UO_2417 (O_2417,N_23065,N_22082);
or UO_2418 (O_2418,N_23900,N_23699);
or UO_2419 (O_2419,N_21928,N_24816);
nand UO_2420 (O_2420,N_22693,N_23079);
xnor UO_2421 (O_2421,N_22803,N_23132);
xnor UO_2422 (O_2422,N_23303,N_23012);
xor UO_2423 (O_2423,N_23684,N_23218);
nor UO_2424 (O_2424,N_23419,N_23272);
nor UO_2425 (O_2425,N_23194,N_23647);
nor UO_2426 (O_2426,N_24625,N_22757);
nor UO_2427 (O_2427,N_23846,N_23763);
and UO_2428 (O_2428,N_24906,N_24176);
xor UO_2429 (O_2429,N_24582,N_24254);
or UO_2430 (O_2430,N_23116,N_23735);
and UO_2431 (O_2431,N_21935,N_24798);
nand UO_2432 (O_2432,N_23573,N_22509);
or UO_2433 (O_2433,N_22291,N_24449);
or UO_2434 (O_2434,N_22976,N_22154);
xor UO_2435 (O_2435,N_24301,N_22856);
nor UO_2436 (O_2436,N_24258,N_23664);
and UO_2437 (O_2437,N_22978,N_22748);
nand UO_2438 (O_2438,N_24066,N_23135);
nand UO_2439 (O_2439,N_23339,N_24974);
xnor UO_2440 (O_2440,N_24133,N_24055);
nor UO_2441 (O_2441,N_22859,N_24834);
nor UO_2442 (O_2442,N_24927,N_22060);
nand UO_2443 (O_2443,N_23015,N_24856);
and UO_2444 (O_2444,N_23058,N_22561);
xor UO_2445 (O_2445,N_22130,N_24779);
nand UO_2446 (O_2446,N_22419,N_22344);
or UO_2447 (O_2447,N_23470,N_22203);
nor UO_2448 (O_2448,N_24689,N_23721);
xnor UO_2449 (O_2449,N_22499,N_22836);
and UO_2450 (O_2450,N_23469,N_24992);
nand UO_2451 (O_2451,N_24801,N_24939);
nor UO_2452 (O_2452,N_23966,N_24799);
or UO_2453 (O_2453,N_22191,N_22201);
and UO_2454 (O_2454,N_24442,N_24632);
nor UO_2455 (O_2455,N_22329,N_21988);
nand UO_2456 (O_2456,N_23740,N_23743);
and UO_2457 (O_2457,N_22190,N_24792);
nand UO_2458 (O_2458,N_22324,N_24802);
xnor UO_2459 (O_2459,N_21906,N_23441);
xnor UO_2460 (O_2460,N_24407,N_24666);
xnor UO_2461 (O_2461,N_24945,N_23420);
nor UO_2462 (O_2462,N_22939,N_24468);
nor UO_2463 (O_2463,N_22447,N_23272);
nand UO_2464 (O_2464,N_23440,N_24576);
nand UO_2465 (O_2465,N_22508,N_23078);
xor UO_2466 (O_2466,N_23283,N_22125);
and UO_2467 (O_2467,N_22972,N_24009);
nand UO_2468 (O_2468,N_24238,N_23084);
xnor UO_2469 (O_2469,N_23707,N_23265);
xnor UO_2470 (O_2470,N_22225,N_23501);
nor UO_2471 (O_2471,N_23087,N_22952);
xnor UO_2472 (O_2472,N_23015,N_24485);
nor UO_2473 (O_2473,N_24352,N_22271);
nor UO_2474 (O_2474,N_24768,N_24933);
and UO_2475 (O_2475,N_22137,N_23650);
or UO_2476 (O_2476,N_23176,N_23571);
and UO_2477 (O_2477,N_23439,N_23389);
and UO_2478 (O_2478,N_24842,N_24737);
nand UO_2479 (O_2479,N_21918,N_23086);
and UO_2480 (O_2480,N_23245,N_22273);
or UO_2481 (O_2481,N_23437,N_24457);
nand UO_2482 (O_2482,N_22473,N_21976);
or UO_2483 (O_2483,N_24227,N_23271);
or UO_2484 (O_2484,N_23737,N_23271);
nor UO_2485 (O_2485,N_24785,N_24266);
and UO_2486 (O_2486,N_22571,N_24600);
xnor UO_2487 (O_2487,N_21936,N_23179);
nor UO_2488 (O_2488,N_23751,N_23445);
xnor UO_2489 (O_2489,N_23883,N_22607);
xnor UO_2490 (O_2490,N_23640,N_21880);
nor UO_2491 (O_2491,N_24664,N_22856);
nor UO_2492 (O_2492,N_22075,N_24720);
or UO_2493 (O_2493,N_23605,N_24592);
nor UO_2494 (O_2494,N_22855,N_22647);
and UO_2495 (O_2495,N_22976,N_22813);
nand UO_2496 (O_2496,N_24379,N_24143);
or UO_2497 (O_2497,N_23775,N_21970);
nand UO_2498 (O_2498,N_24496,N_22603);
and UO_2499 (O_2499,N_22821,N_22339);
nor UO_2500 (O_2500,N_22999,N_23966);
nor UO_2501 (O_2501,N_22732,N_23266);
nor UO_2502 (O_2502,N_22426,N_23907);
nor UO_2503 (O_2503,N_23843,N_23621);
or UO_2504 (O_2504,N_23132,N_23046);
nand UO_2505 (O_2505,N_22008,N_23164);
nor UO_2506 (O_2506,N_23603,N_22279);
or UO_2507 (O_2507,N_21960,N_21930);
and UO_2508 (O_2508,N_24196,N_22809);
or UO_2509 (O_2509,N_24668,N_24851);
and UO_2510 (O_2510,N_22565,N_22743);
or UO_2511 (O_2511,N_22867,N_23580);
nor UO_2512 (O_2512,N_22840,N_24809);
or UO_2513 (O_2513,N_24290,N_24453);
xnor UO_2514 (O_2514,N_22736,N_23563);
nand UO_2515 (O_2515,N_24154,N_22535);
or UO_2516 (O_2516,N_22822,N_23535);
and UO_2517 (O_2517,N_24762,N_22504);
and UO_2518 (O_2518,N_24988,N_22235);
nor UO_2519 (O_2519,N_24684,N_23593);
xor UO_2520 (O_2520,N_22596,N_24326);
or UO_2521 (O_2521,N_24860,N_23905);
nand UO_2522 (O_2522,N_22306,N_23085);
or UO_2523 (O_2523,N_22746,N_24137);
nand UO_2524 (O_2524,N_24811,N_22469);
nor UO_2525 (O_2525,N_23364,N_22881);
xnor UO_2526 (O_2526,N_24059,N_22737);
or UO_2527 (O_2527,N_23618,N_22849);
and UO_2528 (O_2528,N_22883,N_22906);
and UO_2529 (O_2529,N_24168,N_23197);
nand UO_2530 (O_2530,N_22862,N_23966);
or UO_2531 (O_2531,N_23773,N_24854);
and UO_2532 (O_2532,N_23550,N_23688);
or UO_2533 (O_2533,N_22016,N_24894);
nand UO_2534 (O_2534,N_24598,N_23804);
or UO_2535 (O_2535,N_24880,N_21993);
or UO_2536 (O_2536,N_22644,N_23983);
and UO_2537 (O_2537,N_22513,N_23334);
nand UO_2538 (O_2538,N_22741,N_24049);
nand UO_2539 (O_2539,N_23553,N_24092);
nand UO_2540 (O_2540,N_23203,N_24268);
nor UO_2541 (O_2541,N_23187,N_22515);
nand UO_2542 (O_2542,N_23031,N_23219);
nor UO_2543 (O_2543,N_23427,N_21958);
nand UO_2544 (O_2544,N_22458,N_24321);
and UO_2545 (O_2545,N_23798,N_22142);
xor UO_2546 (O_2546,N_22013,N_24729);
nand UO_2547 (O_2547,N_24747,N_23621);
nor UO_2548 (O_2548,N_24999,N_24454);
and UO_2549 (O_2549,N_22389,N_24366);
xor UO_2550 (O_2550,N_21892,N_24415);
or UO_2551 (O_2551,N_22968,N_22391);
nor UO_2552 (O_2552,N_24935,N_23549);
nor UO_2553 (O_2553,N_23027,N_23823);
or UO_2554 (O_2554,N_24119,N_22064);
or UO_2555 (O_2555,N_21939,N_22786);
xor UO_2556 (O_2556,N_23326,N_23592);
nor UO_2557 (O_2557,N_23298,N_23836);
or UO_2558 (O_2558,N_22109,N_22260);
nand UO_2559 (O_2559,N_24514,N_22434);
or UO_2560 (O_2560,N_24430,N_22940);
or UO_2561 (O_2561,N_24851,N_22305);
or UO_2562 (O_2562,N_23114,N_23176);
or UO_2563 (O_2563,N_22280,N_23844);
nor UO_2564 (O_2564,N_23937,N_23180);
and UO_2565 (O_2565,N_22084,N_24618);
or UO_2566 (O_2566,N_23676,N_23941);
and UO_2567 (O_2567,N_22278,N_24315);
xor UO_2568 (O_2568,N_23021,N_23287);
nand UO_2569 (O_2569,N_23839,N_24377);
nand UO_2570 (O_2570,N_22784,N_22261);
nor UO_2571 (O_2571,N_24071,N_23629);
nor UO_2572 (O_2572,N_24413,N_23346);
xor UO_2573 (O_2573,N_22463,N_23918);
and UO_2574 (O_2574,N_24993,N_23709);
nand UO_2575 (O_2575,N_23891,N_23338);
or UO_2576 (O_2576,N_22437,N_24229);
nor UO_2577 (O_2577,N_21908,N_23994);
nand UO_2578 (O_2578,N_24134,N_22429);
nor UO_2579 (O_2579,N_23155,N_24154);
xnor UO_2580 (O_2580,N_23896,N_23510);
and UO_2581 (O_2581,N_23967,N_22589);
nand UO_2582 (O_2582,N_22527,N_22967);
or UO_2583 (O_2583,N_23824,N_23367);
xor UO_2584 (O_2584,N_22147,N_23998);
or UO_2585 (O_2585,N_24657,N_23926);
nor UO_2586 (O_2586,N_22424,N_22104);
xor UO_2587 (O_2587,N_22780,N_24795);
or UO_2588 (O_2588,N_22073,N_21979);
nor UO_2589 (O_2589,N_24042,N_24618);
or UO_2590 (O_2590,N_22295,N_22010);
or UO_2591 (O_2591,N_24151,N_23119);
or UO_2592 (O_2592,N_23087,N_24194);
and UO_2593 (O_2593,N_22070,N_22289);
xnor UO_2594 (O_2594,N_23390,N_23699);
and UO_2595 (O_2595,N_24136,N_21942);
or UO_2596 (O_2596,N_23140,N_23965);
and UO_2597 (O_2597,N_24803,N_22101);
xor UO_2598 (O_2598,N_23000,N_24911);
xor UO_2599 (O_2599,N_24762,N_22840);
and UO_2600 (O_2600,N_21973,N_22648);
and UO_2601 (O_2601,N_24375,N_22292);
nor UO_2602 (O_2602,N_22307,N_24317);
xor UO_2603 (O_2603,N_23110,N_23192);
and UO_2604 (O_2604,N_24653,N_23700);
or UO_2605 (O_2605,N_23660,N_24402);
and UO_2606 (O_2606,N_24274,N_22091);
xnor UO_2607 (O_2607,N_23621,N_24028);
and UO_2608 (O_2608,N_22200,N_23056);
nand UO_2609 (O_2609,N_24507,N_24353);
nand UO_2610 (O_2610,N_22289,N_24430);
and UO_2611 (O_2611,N_22398,N_23160);
xnor UO_2612 (O_2612,N_22142,N_22951);
nor UO_2613 (O_2613,N_24391,N_23507);
nand UO_2614 (O_2614,N_22777,N_24355);
nor UO_2615 (O_2615,N_23412,N_23281);
nand UO_2616 (O_2616,N_22377,N_22097);
nor UO_2617 (O_2617,N_22510,N_23281);
xnor UO_2618 (O_2618,N_23199,N_21945);
xor UO_2619 (O_2619,N_24988,N_24033);
xnor UO_2620 (O_2620,N_23258,N_22085);
nand UO_2621 (O_2621,N_22390,N_22465);
nand UO_2622 (O_2622,N_22737,N_23769);
and UO_2623 (O_2623,N_22969,N_22011);
nand UO_2624 (O_2624,N_23851,N_23282);
nand UO_2625 (O_2625,N_24708,N_23304);
nor UO_2626 (O_2626,N_24898,N_22902);
and UO_2627 (O_2627,N_22010,N_24290);
xor UO_2628 (O_2628,N_22782,N_23184);
and UO_2629 (O_2629,N_23267,N_24659);
or UO_2630 (O_2630,N_22994,N_22518);
or UO_2631 (O_2631,N_24318,N_22665);
xor UO_2632 (O_2632,N_23853,N_22241);
nand UO_2633 (O_2633,N_22005,N_23534);
or UO_2634 (O_2634,N_22089,N_23944);
and UO_2635 (O_2635,N_24035,N_22368);
nand UO_2636 (O_2636,N_22316,N_23657);
or UO_2637 (O_2637,N_24886,N_24667);
and UO_2638 (O_2638,N_23047,N_22193);
or UO_2639 (O_2639,N_23563,N_22133);
and UO_2640 (O_2640,N_24156,N_23934);
nor UO_2641 (O_2641,N_23250,N_24753);
xor UO_2642 (O_2642,N_23184,N_24578);
nand UO_2643 (O_2643,N_23715,N_24033);
nand UO_2644 (O_2644,N_22189,N_24430);
nor UO_2645 (O_2645,N_23350,N_24731);
or UO_2646 (O_2646,N_24279,N_23970);
or UO_2647 (O_2647,N_23623,N_24531);
nand UO_2648 (O_2648,N_24350,N_22444);
nand UO_2649 (O_2649,N_23223,N_23151);
nand UO_2650 (O_2650,N_22379,N_22077);
xor UO_2651 (O_2651,N_23347,N_24169);
and UO_2652 (O_2652,N_22396,N_24417);
or UO_2653 (O_2653,N_24297,N_24347);
or UO_2654 (O_2654,N_22640,N_22238);
and UO_2655 (O_2655,N_24234,N_23319);
and UO_2656 (O_2656,N_24869,N_24742);
or UO_2657 (O_2657,N_24175,N_24729);
nor UO_2658 (O_2658,N_24052,N_21984);
xnor UO_2659 (O_2659,N_23406,N_23437);
nand UO_2660 (O_2660,N_23473,N_23946);
nand UO_2661 (O_2661,N_22419,N_23813);
xnor UO_2662 (O_2662,N_24736,N_23249);
and UO_2663 (O_2663,N_24911,N_22827);
and UO_2664 (O_2664,N_22890,N_22205);
xor UO_2665 (O_2665,N_23047,N_23614);
and UO_2666 (O_2666,N_22792,N_24984);
nand UO_2667 (O_2667,N_22974,N_23416);
nor UO_2668 (O_2668,N_22436,N_23825);
and UO_2669 (O_2669,N_23065,N_23458);
nand UO_2670 (O_2670,N_24770,N_23375);
xnor UO_2671 (O_2671,N_22685,N_22061);
nand UO_2672 (O_2672,N_22732,N_22713);
or UO_2673 (O_2673,N_23182,N_22419);
xor UO_2674 (O_2674,N_23878,N_22890);
xnor UO_2675 (O_2675,N_22848,N_24538);
nand UO_2676 (O_2676,N_23291,N_24347);
or UO_2677 (O_2677,N_23452,N_23137);
or UO_2678 (O_2678,N_22659,N_22420);
xnor UO_2679 (O_2679,N_21937,N_22578);
xor UO_2680 (O_2680,N_23953,N_23883);
nand UO_2681 (O_2681,N_23404,N_22160);
nor UO_2682 (O_2682,N_22228,N_22852);
or UO_2683 (O_2683,N_22190,N_24962);
nand UO_2684 (O_2684,N_24345,N_24078);
and UO_2685 (O_2685,N_24111,N_24347);
or UO_2686 (O_2686,N_23977,N_21929);
and UO_2687 (O_2687,N_24315,N_23991);
and UO_2688 (O_2688,N_22117,N_23945);
nand UO_2689 (O_2689,N_23864,N_23204);
and UO_2690 (O_2690,N_24959,N_22695);
nand UO_2691 (O_2691,N_23499,N_22214);
xnor UO_2692 (O_2692,N_22944,N_22373);
and UO_2693 (O_2693,N_24701,N_24140);
xnor UO_2694 (O_2694,N_23634,N_22540);
or UO_2695 (O_2695,N_24950,N_23494);
or UO_2696 (O_2696,N_23775,N_23422);
nor UO_2697 (O_2697,N_24572,N_23035);
and UO_2698 (O_2698,N_24135,N_24479);
and UO_2699 (O_2699,N_23628,N_22882);
or UO_2700 (O_2700,N_22599,N_22295);
xnor UO_2701 (O_2701,N_24182,N_23750);
nor UO_2702 (O_2702,N_23604,N_22223);
nor UO_2703 (O_2703,N_24787,N_23088);
xnor UO_2704 (O_2704,N_24038,N_24206);
or UO_2705 (O_2705,N_23102,N_22057);
nand UO_2706 (O_2706,N_22290,N_21916);
and UO_2707 (O_2707,N_23221,N_24625);
and UO_2708 (O_2708,N_23168,N_22684);
and UO_2709 (O_2709,N_23156,N_23646);
and UO_2710 (O_2710,N_23580,N_24122);
or UO_2711 (O_2711,N_24656,N_23506);
nand UO_2712 (O_2712,N_23487,N_22449);
nor UO_2713 (O_2713,N_24364,N_24874);
nor UO_2714 (O_2714,N_24389,N_22814);
and UO_2715 (O_2715,N_22316,N_23831);
and UO_2716 (O_2716,N_24850,N_23456);
or UO_2717 (O_2717,N_22088,N_22965);
xor UO_2718 (O_2718,N_22701,N_22006);
nor UO_2719 (O_2719,N_22165,N_22922);
nor UO_2720 (O_2720,N_24323,N_22787);
and UO_2721 (O_2721,N_23452,N_23732);
and UO_2722 (O_2722,N_24818,N_24951);
nand UO_2723 (O_2723,N_24808,N_22135);
nand UO_2724 (O_2724,N_23633,N_22942);
or UO_2725 (O_2725,N_23505,N_24112);
xor UO_2726 (O_2726,N_22486,N_22348);
xnor UO_2727 (O_2727,N_23279,N_23530);
or UO_2728 (O_2728,N_24294,N_22306);
and UO_2729 (O_2729,N_23081,N_22121);
or UO_2730 (O_2730,N_22789,N_24453);
xnor UO_2731 (O_2731,N_23700,N_22418);
nor UO_2732 (O_2732,N_22945,N_22494);
nor UO_2733 (O_2733,N_23385,N_24643);
nor UO_2734 (O_2734,N_24540,N_23435);
or UO_2735 (O_2735,N_24617,N_22203);
nor UO_2736 (O_2736,N_22712,N_23801);
xor UO_2737 (O_2737,N_24244,N_22751);
nor UO_2738 (O_2738,N_24313,N_23028);
xor UO_2739 (O_2739,N_24952,N_22779);
or UO_2740 (O_2740,N_22898,N_22605);
nor UO_2741 (O_2741,N_22741,N_24809);
or UO_2742 (O_2742,N_22823,N_23663);
nand UO_2743 (O_2743,N_22245,N_24198);
xor UO_2744 (O_2744,N_23822,N_24334);
or UO_2745 (O_2745,N_22299,N_23540);
xnor UO_2746 (O_2746,N_22186,N_22944);
nor UO_2747 (O_2747,N_23422,N_23113);
or UO_2748 (O_2748,N_22152,N_24026);
xor UO_2749 (O_2749,N_22815,N_23927);
xnor UO_2750 (O_2750,N_23736,N_23938);
or UO_2751 (O_2751,N_23205,N_24498);
and UO_2752 (O_2752,N_24489,N_24052);
nand UO_2753 (O_2753,N_22819,N_22132);
nor UO_2754 (O_2754,N_22217,N_23127);
or UO_2755 (O_2755,N_24796,N_23759);
nor UO_2756 (O_2756,N_22532,N_23996);
and UO_2757 (O_2757,N_24024,N_24200);
xor UO_2758 (O_2758,N_24781,N_24306);
and UO_2759 (O_2759,N_22727,N_22896);
or UO_2760 (O_2760,N_23089,N_24205);
or UO_2761 (O_2761,N_22443,N_22360);
nand UO_2762 (O_2762,N_24400,N_24350);
xor UO_2763 (O_2763,N_24989,N_24892);
nand UO_2764 (O_2764,N_23926,N_24436);
xnor UO_2765 (O_2765,N_23147,N_22161);
xor UO_2766 (O_2766,N_24813,N_23258);
nor UO_2767 (O_2767,N_23516,N_23818);
or UO_2768 (O_2768,N_22288,N_24428);
nand UO_2769 (O_2769,N_21892,N_24565);
nand UO_2770 (O_2770,N_23115,N_22720);
nand UO_2771 (O_2771,N_24254,N_22135);
and UO_2772 (O_2772,N_22295,N_23486);
nor UO_2773 (O_2773,N_23402,N_22298);
or UO_2774 (O_2774,N_23901,N_24062);
xor UO_2775 (O_2775,N_23857,N_22447);
nor UO_2776 (O_2776,N_23504,N_23253);
or UO_2777 (O_2777,N_23277,N_24614);
or UO_2778 (O_2778,N_22616,N_23886);
and UO_2779 (O_2779,N_24451,N_23115);
and UO_2780 (O_2780,N_23100,N_22534);
or UO_2781 (O_2781,N_22175,N_23503);
nand UO_2782 (O_2782,N_22497,N_22949);
or UO_2783 (O_2783,N_23509,N_22582);
nor UO_2784 (O_2784,N_23267,N_24688);
or UO_2785 (O_2785,N_23103,N_22930);
and UO_2786 (O_2786,N_23815,N_22338);
nand UO_2787 (O_2787,N_22515,N_24848);
nand UO_2788 (O_2788,N_23709,N_22172);
or UO_2789 (O_2789,N_24917,N_22483);
and UO_2790 (O_2790,N_24623,N_22639);
xnor UO_2791 (O_2791,N_24808,N_22124);
xor UO_2792 (O_2792,N_22480,N_22238);
nand UO_2793 (O_2793,N_22567,N_22081);
and UO_2794 (O_2794,N_24364,N_24784);
nor UO_2795 (O_2795,N_22431,N_22267);
and UO_2796 (O_2796,N_24461,N_24831);
nor UO_2797 (O_2797,N_22425,N_23080);
and UO_2798 (O_2798,N_24463,N_24708);
xnor UO_2799 (O_2799,N_24591,N_22712);
or UO_2800 (O_2800,N_23106,N_22527);
or UO_2801 (O_2801,N_24155,N_22004);
or UO_2802 (O_2802,N_22021,N_23270);
or UO_2803 (O_2803,N_23133,N_24085);
xnor UO_2804 (O_2804,N_22617,N_22796);
nand UO_2805 (O_2805,N_24636,N_21945);
or UO_2806 (O_2806,N_22900,N_24655);
and UO_2807 (O_2807,N_23106,N_22869);
nand UO_2808 (O_2808,N_24929,N_23815);
xor UO_2809 (O_2809,N_22536,N_24618);
xor UO_2810 (O_2810,N_22026,N_24151);
or UO_2811 (O_2811,N_24526,N_22689);
nor UO_2812 (O_2812,N_22960,N_22898);
or UO_2813 (O_2813,N_24815,N_23746);
and UO_2814 (O_2814,N_23624,N_22419);
xor UO_2815 (O_2815,N_22303,N_23900);
or UO_2816 (O_2816,N_23805,N_22475);
nand UO_2817 (O_2817,N_22866,N_24899);
nand UO_2818 (O_2818,N_23657,N_22119);
xor UO_2819 (O_2819,N_22900,N_22949);
xnor UO_2820 (O_2820,N_23965,N_24961);
and UO_2821 (O_2821,N_24070,N_22132);
or UO_2822 (O_2822,N_22274,N_23186);
and UO_2823 (O_2823,N_24861,N_23472);
nor UO_2824 (O_2824,N_24731,N_22861);
nand UO_2825 (O_2825,N_22143,N_22442);
and UO_2826 (O_2826,N_24179,N_23311);
nand UO_2827 (O_2827,N_22873,N_22703);
and UO_2828 (O_2828,N_22922,N_24347);
or UO_2829 (O_2829,N_23416,N_24807);
nand UO_2830 (O_2830,N_23022,N_22087);
and UO_2831 (O_2831,N_24922,N_22298);
and UO_2832 (O_2832,N_23342,N_23093);
and UO_2833 (O_2833,N_22276,N_23557);
nor UO_2834 (O_2834,N_22156,N_22845);
nand UO_2835 (O_2835,N_22775,N_23733);
and UO_2836 (O_2836,N_22718,N_24244);
nor UO_2837 (O_2837,N_22978,N_24502);
nand UO_2838 (O_2838,N_24238,N_22681);
nor UO_2839 (O_2839,N_22724,N_24534);
and UO_2840 (O_2840,N_22308,N_23681);
and UO_2841 (O_2841,N_24069,N_22511);
or UO_2842 (O_2842,N_23873,N_23796);
nand UO_2843 (O_2843,N_22798,N_23263);
and UO_2844 (O_2844,N_22709,N_24006);
xor UO_2845 (O_2845,N_22728,N_22184);
or UO_2846 (O_2846,N_24285,N_23640);
xnor UO_2847 (O_2847,N_22027,N_24931);
nand UO_2848 (O_2848,N_22856,N_24423);
nor UO_2849 (O_2849,N_24174,N_23663);
or UO_2850 (O_2850,N_24622,N_24704);
xnor UO_2851 (O_2851,N_22156,N_23289);
or UO_2852 (O_2852,N_24571,N_23641);
nand UO_2853 (O_2853,N_22433,N_23206);
nand UO_2854 (O_2854,N_23224,N_24775);
or UO_2855 (O_2855,N_23309,N_22339);
and UO_2856 (O_2856,N_24104,N_22799);
or UO_2857 (O_2857,N_22837,N_23818);
nand UO_2858 (O_2858,N_23918,N_22484);
or UO_2859 (O_2859,N_24089,N_23379);
and UO_2860 (O_2860,N_24990,N_23957);
nor UO_2861 (O_2861,N_23759,N_23179);
xor UO_2862 (O_2862,N_22303,N_24062);
nand UO_2863 (O_2863,N_22046,N_22259);
nor UO_2864 (O_2864,N_22238,N_23479);
or UO_2865 (O_2865,N_22573,N_22872);
nand UO_2866 (O_2866,N_24037,N_23899);
nor UO_2867 (O_2867,N_23487,N_23332);
nand UO_2868 (O_2868,N_22337,N_23356);
xor UO_2869 (O_2869,N_23034,N_22496);
xnor UO_2870 (O_2870,N_24320,N_22291);
and UO_2871 (O_2871,N_23071,N_24133);
and UO_2872 (O_2872,N_24612,N_22162);
and UO_2873 (O_2873,N_24713,N_22791);
xnor UO_2874 (O_2874,N_24561,N_22711);
nor UO_2875 (O_2875,N_22431,N_24153);
or UO_2876 (O_2876,N_22646,N_24950);
nand UO_2877 (O_2877,N_24753,N_21911);
or UO_2878 (O_2878,N_24373,N_24698);
and UO_2879 (O_2879,N_24075,N_24790);
or UO_2880 (O_2880,N_24989,N_23067);
nand UO_2881 (O_2881,N_24543,N_22253);
nand UO_2882 (O_2882,N_23209,N_23762);
xnor UO_2883 (O_2883,N_24842,N_23936);
xnor UO_2884 (O_2884,N_23276,N_24640);
xnor UO_2885 (O_2885,N_22775,N_24862);
nand UO_2886 (O_2886,N_24737,N_23182);
xnor UO_2887 (O_2887,N_23744,N_23360);
and UO_2888 (O_2888,N_23286,N_22970);
or UO_2889 (O_2889,N_23046,N_24788);
or UO_2890 (O_2890,N_22681,N_22669);
or UO_2891 (O_2891,N_24267,N_24020);
nor UO_2892 (O_2892,N_24477,N_23717);
xor UO_2893 (O_2893,N_22782,N_24826);
or UO_2894 (O_2894,N_22148,N_23502);
xor UO_2895 (O_2895,N_23865,N_22836);
nand UO_2896 (O_2896,N_23949,N_24827);
nand UO_2897 (O_2897,N_23606,N_22258);
or UO_2898 (O_2898,N_24912,N_22781);
nand UO_2899 (O_2899,N_24177,N_22505);
nor UO_2900 (O_2900,N_22197,N_24842);
and UO_2901 (O_2901,N_23573,N_23759);
or UO_2902 (O_2902,N_22497,N_22360);
nand UO_2903 (O_2903,N_22460,N_23496);
xor UO_2904 (O_2904,N_24067,N_24995);
nand UO_2905 (O_2905,N_22231,N_22104);
or UO_2906 (O_2906,N_22728,N_22631);
nand UO_2907 (O_2907,N_24100,N_22458);
xnor UO_2908 (O_2908,N_23218,N_24902);
nor UO_2909 (O_2909,N_23082,N_23423);
and UO_2910 (O_2910,N_22405,N_23296);
and UO_2911 (O_2911,N_22719,N_23810);
nand UO_2912 (O_2912,N_23792,N_22237);
and UO_2913 (O_2913,N_23689,N_23971);
xnor UO_2914 (O_2914,N_24240,N_23337);
and UO_2915 (O_2915,N_22832,N_22611);
or UO_2916 (O_2916,N_23159,N_24441);
or UO_2917 (O_2917,N_22172,N_24829);
or UO_2918 (O_2918,N_23570,N_24994);
nand UO_2919 (O_2919,N_21910,N_24445);
nand UO_2920 (O_2920,N_24682,N_24561);
and UO_2921 (O_2921,N_21903,N_22661);
nor UO_2922 (O_2922,N_23973,N_23722);
or UO_2923 (O_2923,N_24460,N_23793);
nor UO_2924 (O_2924,N_22548,N_24401);
xnor UO_2925 (O_2925,N_23412,N_22570);
or UO_2926 (O_2926,N_22859,N_24156);
or UO_2927 (O_2927,N_22503,N_23010);
xor UO_2928 (O_2928,N_23299,N_24375);
nor UO_2929 (O_2929,N_23072,N_23286);
nor UO_2930 (O_2930,N_22940,N_22494);
nand UO_2931 (O_2931,N_24955,N_22918);
nand UO_2932 (O_2932,N_22854,N_23766);
nor UO_2933 (O_2933,N_24802,N_22597);
xor UO_2934 (O_2934,N_24796,N_22588);
and UO_2935 (O_2935,N_24762,N_24752);
xnor UO_2936 (O_2936,N_24988,N_24483);
or UO_2937 (O_2937,N_24797,N_24414);
and UO_2938 (O_2938,N_24112,N_23025);
and UO_2939 (O_2939,N_23313,N_23956);
and UO_2940 (O_2940,N_23380,N_22036);
or UO_2941 (O_2941,N_23168,N_22121);
nor UO_2942 (O_2942,N_21908,N_22621);
xor UO_2943 (O_2943,N_24257,N_22370);
and UO_2944 (O_2944,N_22039,N_21987);
xnor UO_2945 (O_2945,N_22784,N_22062);
or UO_2946 (O_2946,N_24395,N_24639);
nor UO_2947 (O_2947,N_24390,N_23112);
xnor UO_2948 (O_2948,N_24654,N_23918);
nand UO_2949 (O_2949,N_22173,N_23003);
or UO_2950 (O_2950,N_24166,N_24320);
nand UO_2951 (O_2951,N_23782,N_24263);
xor UO_2952 (O_2952,N_24389,N_22494);
or UO_2953 (O_2953,N_21921,N_24556);
nand UO_2954 (O_2954,N_22340,N_23494);
and UO_2955 (O_2955,N_22895,N_22614);
nor UO_2956 (O_2956,N_24262,N_22652);
and UO_2957 (O_2957,N_23720,N_24575);
nor UO_2958 (O_2958,N_24829,N_24192);
and UO_2959 (O_2959,N_22678,N_21947);
and UO_2960 (O_2960,N_22225,N_22175);
xnor UO_2961 (O_2961,N_24902,N_23340);
or UO_2962 (O_2962,N_23469,N_24846);
xor UO_2963 (O_2963,N_22133,N_23644);
xor UO_2964 (O_2964,N_23621,N_22321);
nand UO_2965 (O_2965,N_24998,N_22925);
nand UO_2966 (O_2966,N_24034,N_23471);
nor UO_2967 (O_2967,N_22210,N_23916);
xor UO_2968 (O_2968,N_23571,N_22715);
and UO_2969 (O_2969,N_22505,N_24499);
and UO_2970 (O_2970,N_23066,N_23142);
or UO_2971 (O_2971,N_22713,N_23747);
or UO_2972 (O_2972,N_22284,N_24082);
xnor UO_2973 (O_2973,N_24271,N_23036);
or UO_2974 (O_2974,N_24274,N_24735);
nor UO_2975 (O_2975,N_24461,N_22749);
and UO_2976 (O_2976,N_22056,N_21908);
nand UO_2977 (O_2977,N_24371,N_24849);
nand UO_2978 (O_2978,N_22776,N_24226);
nor UO_2979 (O_2979,N_24338,N_22374);
or UO_2980 (O_2980,N_22992,N_23991);
xor UO_2981 (O_2981,N_24465,N_22954);
nor UO_2982 (O_2982,N_24915,N_23462);
and UO_2983 (O_2983,N_24408,N_24926);
nor UO_2984 (O_2984,N_21895,N_22428);
or UO_2985 (O_2985,N_22249,N_23018);
xnor UO_2986 (O_2986,N_24231,N_23499);
or UO_2987 (O_2987,N_21952,N_24372);
xnor UO_2988 (O_2988,N_24378,N_23109);
xnor UO_2989 (O_2989,N_24459,N_22940);
xor UO_2990 (O_2990,N_24999,N_24356);
nor UO_2991 (O_2991,N_23830,N_23001);
nand UO_2992 (O_2992,N_22468,N_24341);
xnor UO_2993 (O_2993,N_24472,N_24953);
nor UO_2994 (O_2994,N_23438,N_22849);
and UO_2995 (O_2995,N_23012,N_21906);
nor UO_2996 (O_2996,N_22039,N_23547);
nor UO_2997 (O_2997,N_22581,N_24427);
and UO_2998 (O_2998,N_24905,N_24737);
xnor UO_2999 (O_2999,N_23631,N_24815);
endmodule