module basic_500_3000_500_15_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_236,In_180);
or U1 (N_1,In_448,In_199);
nand U2 (N_2,In_261,In_463);
nand U3 (N_3,In_240,In_206);
nand U4 (N_4,In_499,In_410);
and U5 (N_5,In_406,In_347);
nand U6 (N_6,In_132,In_229);
and U7 (N_7,In_461,In_320);
nand U8 (N_8,In_210,In_85);
nand U9 (N_9,In_83,In_327);
nand U10 (N_10,In_198,In_262);
nor U11 (N_11,In_148,In_248);
nor U12 (N_12,In_219,In_93);
nand U13 (N_13,In_189,In_196);
nor U14 (N_14,In_481,In_170);
xor U15 (N_15,In_111,In_444);
and U16 (N_16,In_187,In_139);
nand U17 (N_17,In_264,In_204);
nand U18 (N_18,In_119,In_355);
nor U19 (N_19,In_422,In_354);
nand U20 (N_20,In_97,In_98);
nor U21 (N_21,In_321,In_177);
nor U22 (N_22,In_122,In_82);
nor U23 (N_23,In_245,In_62);
and U24 (N_24,In_446,In_226);
nand U25 (N_25,In_358,In_183);
or U26 (N_26,In_175,In_53);
or U27 (N_27,In_151,In_263);
nand U28 (N_28,In_441,In_471);
or U29 (N_29,In_389,In_84);
nand U30 (N_30,In_49,In_468);
nand U31 (N_31,In_457,In_173);
nor U32 (N_32,In_246,In_150);
and U33 (N_33,In_96,In_87);
xor U34 (N_34,In_144,In_393);
nand U35 (N_35,In_5,In_75);
nand U36 (N_36,In_54,In_202);
or U37 (N_37,In_162,In_216);
or U38 (N_38,In_88,In_214);
nand U39 (N_39,In_312,In_67);
nor U40 (N_40,In_369,In_290);
and U41 (N_41,In_419,In_424);
and U42 (N_42,In_326,In_439);
xnor U43 (N_43,In_351,In_251);
and U44 (N_44,In_69,In_318);
or U45 (N_45,In_239,In_495);
nand U46 (N_46,In_357,In_185);
or U47 (N_47,In_108,In_466);
nand U48 (N_48,In_449,In_141);
and U49 (N_49,In_287,In_137);
and U50 (N_50,In_138,In_257);
and U51 (N_51,In_1,In_289);
nand U52 (N_52,In_277,In_160);
or U53 (N_53,In_403,In_135);
and U54 (N_54,In_109,In_184);
or U55 (N_55,In_303,In_456);
and U56 (N_56,In_314,In_21);
nand U57 (N_57,In_417,In_102);
nor U58 (N_58,In_193,In_55);
nor U59 (N_59,In_285,In_411);
and U60 (N_60,In_498,In_294);
nor U61 (N_61,In_359,In_352);
and U62 (N_62,In_408,In_415);
nand U63 (N_63,In_483,In_68);
nand U64 (N_64,In_100,In_3);
and U65 (N_65,In_366,In_43);
nand U66 (N_66,In_372,In_26);
and U67 (N_67,In_61,In_433);
and U68 (N_68,In_258,In_301);
or U69 (N_69,In_434,In_377);
or U70 (N_70,In_237,In_106);
and U71 (N_71,In_371,In_390);
or U72 (N_72,In_348,In_392);
or U73 (N_73,In_267,In_440);
and U74 (N_74,In_38,In_281);
and U75 (N_75,In_121,In_306);
nor U76 (N_76,In_126,In_117);
xor U77 (N_77,In_33,In_191);
nand U78 (N_78,In_201,In_208);
nand U79 (N_79,In_315,In_101);
and U80 (N_80,In_10,In_431);
nand U81 (N_81,In_114,In_316);
nand U82 (N_82,In_309,In_167);
and U83 (N_83,In_0,In_15);
nor U84 (N_84,In_59,In_271);
and U85 (N_85,In_266,In_493);
nor U86 (N_86,In_460,In_274);
nor U87 (N_87,In_455,In_194);
and U88 (N_88,In_472,In_243);
nor U89 (N_89,In_291,In_491);
nand U90 (N_90,In_116,In_35);
nand U91 (N_91,In_496,In_399);
nand U92 (N_92,In_418,In_242);
nor U93 (N_93,In_211,In_79);
nand U94 (N_94,In_334,In_70);
and U95 (N_95,In_335,In_22);
nor U96 (N_96,In_401,In_385);
nand U97 (N_97,In_473,In_400);
nand U98 (N_98,In_368,In_325);
nor U99 (N_99,In_273,In_272);
and U100 (N_100,In_293,In_310);
xnor U101 (N_101,In_171,In_421);
nor U102 (N_102,In_60,In_428);
nand U103 (N_103,In_124,In_45);
or U104 (N_104,In_343,In_395);
and U105 (N_105,In_91,In_65);
nand U106 (N_106,In_423,In_174);
nand U107 (N_107,In_345,In_292);
nor U108 (N_108,In_182,In_129);
nor U109 (N_109,In_131,In_249);
xnor U110 (N_110,In_11,In_76);
or U111 (N_111,In_299,In_169);
and U112 (N_112,In_391,In_346);
nand U113 (N_113,In_228,In_95);
and U114 (N_114,In_213,In_497);
nor U115 (N_115,In_488,In_103);
nand U116 (N_116,In_373,In_450);
xnor U117 (N_117,In_381,In_247);
and U118 (N_118,In_244,In_110);
nand U119 (N_119,In_363,In_32);
nand U120 (N_120,In_64,In_149);
and U121 (N_121,In_23,In_307);
and U122 (N_122,In_74,In_313);
nand U123 (N_123,In_476,In_232);
xnor U124 (N_124,In_238,In_487);
nand U125 (N_125,In_250,In_28);
nor U126 (N_126,In_337,In_426);
and U127 (N_127,In_482,In_462);
and U128 (N_128,In_402,In_298);
or U129 (N_129,In_397,In_259);
nand U130 (N_130,In_13,In_143);
and U131 (N_131,In_374,In_179);
or U132 (N_132,In_470,In_25);
or U133 (N_133,In_12,In_178);
or U134 (N_134,In_147,In_380);
or U135 (N_135,In_81,In_447);
nor U136 (N_136,In_370,In_207);
xnor U137 (N_137,In_252,In_467);
nor U138 (N_138,In_458,In_378);
nor U139 (N_139,In_4,In_112);
nand U140 (N_140,In_104,In_99);
nor U141 (N_141,In_331,In_490);
nor U142 (N_142,In_24,In_157);
and U143 (N_143,In_19,In_477);
nand U144 (N_144,In_276,In_145);
xnor U145 (N_145,In_73,In_71);
nand U146 (N_146,In_63,In_494);
nand U147 (N_147,In_161,In_376);
or U148 (N_148,In_156,In_452);
or U149 (N_149,In_155,In_361);
nor U150 (N_150,In_14,In_115);
and U151 (N_151,In_260,In_414);
and U152 (N_152,In_459,In_474);
and U153 (N_153,In_52,In_47);
or U154 (N_154,In_77,In_158);
nor U155 (N_155,In_396,In_296);
xor U156 (N_156,In_383,In_323);
and U157 (N_157,In_308,In_31);
nand U158 (N_158,In_479,In_443);
or U159 (N_159,In_270,In_492);
or U160 (N_160,In_225,In_136);
and U161 (N_161,In_478,In_432);
and U162 (N_162,In_279,In_218);
or U163 (N_163,In_409,In_486);
nand U164 (N_164,In_379,In_34);
and U165 (N_165,In_300,In_280);
nor U166 (N_166,In_329,In_107);
or U167 (N_167,In_58,In_420);
and U168 (N_168,In_436,In_367);
and U169 (N_169,In_319,In_235);
or U170 (N_170,In_89,In_181);
or U171 (N_171,In_269,In_453);
nand U172 (N_172,In_27,In_451);
nor U173 (N_173,In_134,In_195);
or U174 (N_174,In_154,In_118);
nand U175 (N_175,In_176,In_283);
nor U176 (N_176,In_407,In_288);
or U177 (N_177,In_317,In_18);
xnor U178 (N_178,In_234,In_442);
nand U179 (N_179,In_253,In_128);
or U180 (N_180,In_212,In_469);
nor U181 (N_181,In_153,In_360);
or U182 (N_182,In_333,In_209);
and U183 (N_183,In_80,In_413);
and U184 (N_184,In_140,In_105);
nor U185 (N_185,In_429,In_278);
and U186 (N_186,In_416,In_336);
or U187 (N_187,In_412,In_480);
nor U188 (N_188,In_230,In_454);
or U189 (N_189,In_36,In_2);
nor U190 (N_190,In_51,In_465);
and U191 (N_191,In_123,In_39);
and U192 (N_192,In_255,In_311);
and U193 (N_193,In_425,In_305);
nor U194 (N_194,In_203,In_215);
nand U195 (N_195,In_254,In_241);
and U196 (N_196,In_6,In_324);
xnor U197 (N_197,In_332,In_437);
nand U198 (N_198,In_7,In_438);
and U199 (N_199,In_17,In_304);
xnor U200 (N_200,N_61,N_32);
and U201 (N_201,N_188,N_97);
or U202 (N_202,In_130,N_74);
or U203 (N_203,N_19,N_11);
and U204 (N_204,In_268,In_286);
xnor U205 (N_205,N_182,N_168);
nor U206 (N_206,N_69,N_174);
or U207 (N_207,N_141,In_265);
nor U208 (N_208,N_180,N_41);
nor U209 (N_209,N_190,In_133);
or U210 (N_210,In_223,In_217);
nand U211 (N_211,In_20,In_398);
nor U212 (N_212,N_30,In_192);
or U213 (N_213,N_139,N_118);
or U214 (N_214,In_42,In_344);
nor U215 (N_215,N_136,N_179);
nor U216 (N_216,In_165,In_220);
and U217 (N_217,N_143,In_375);
and U218 (N_218,N_149,In_29);
or U219 (N_219,N_103,N_7);
nand U220 (N_220,N_132,In_275);
nor U221 (N_221,N_157,In_57);
and U222 (N_222,N_28,N_116);
and U223 (N_223,In_127,N_85);
or U224 (N_224,In_435,N_155);
and U225 (N_225,N_16,N_195);
and U226 (N_226,N_17,In_302);
or U227 (N_227,N_77,In_349);
and U228 (N_228,N_126,N_31);
nor U229 (N_229,In_94,In_342);
nor U230 (N_230,In_164,N_183);
and U231 (N_231,N_8,In_364);
and U232 (N_232,In_384,In_394);
and U233 (N_233,N_1,N_163);
nand U234 (N_234,In_224,N_192);
or U235 (N_235,In_464,In_489);
xnor U236 (N_236,In_9,In_341);
nor U237 (N_237,N_67,N_14);
and U238 (N_238,In_205,N_145);
nand U239 (N_239,N_64,In_475);
or U240 (N_240,N_146,N_47);
nand U241 (N_241,N_18,N_176);
nor U242 (N_242,N_60,N_33);
or U243 (N_243,In_90,N_43);
nand U244 (N_244,In_44,N_73);
or U245 (N_245,N_95,N_184);
xor U246 (N_246,N_127,N_71);
and U247 (N_247,N_86,N_181);
or U248 (N_248,N_37,N_81);
and U249 (N_249,N_102,N_99);
nor U250 (N_250,N_65,N_117);
and U251 (N_251,N_36,N_87);
xor U252 (N_252,In_163,In_233);
nand U253 (N_253,In_484,N_52);
nor U254 (N_254,In_72,N_76);
and U255 (N_255,N_137,N_129);
nor U256 (N_256,N_135,N_185);
or U257 (N_257,N_94,N_113);
nor U258 (N_258,N_6,N_170);
nand U259 (N_259,In_295,N_111);
and U260 (N_260,In_405,N_125);
nor U261 (N_261,N_165,N_120);
or U262 (N_262,In_113,N_130);
nor U263 (N_263,In_297,In_221);
nor U264 (N_264,N_152,In_125);
xor U265 (N_265,In_365,N_148);
nand U266 (N_266,N_29,In_445);
and U267 (N_267,N_24,In_40);
or U268 (N_268,N_175,N_101);
nand U269 (N_269,N_100,N_107);
xor U270 (N_270,N_80,In_37);
nor U271 (N_271,N_9,N_172);
and U272 (N_272,N_196,N_25);
nor U273 (N_273,In_92,In_120);
nor U274 (N_274,N_128,In_338);
and U275 (N_275,In_387,N_75);
or U276 (N_276,In_56,In_172);
xnor U277 (N_277,N_22,In_227);
and U278 (N_278,In_86,N_48);
xor U279 (N_279,N_199,N_173);
and U280 (N_280,In_222,N_54);
or U281 (N_281,N_142,N_171);
and U282 (N_282,N_10,In_142);
or U283 (N_283,N_53,In_382);
or U284 (N_284,N_159,N_122);
nand U285 (N_285,N_197,N_84);
nor U286 (N_286,N_13,N_46);
and U287 (N_287,In_256,In_30);
or U288 (N_288,N_23,In_339);
xor U289 (N_289,N_56,N_138);
nand U290 (N_290,N_144,In_146);
or U291 (N_291,In_159,N_40);
or U292 (N_292,N_49,In_200);
or U293 (N_293,N_198,N_164);
nor U294 (N_294,N_108,N_191);
and U295 (N_295,N_154,N_45);
or U296 (N_296,N_15,N_134);
or U297 (N_297,In_41,N_194);
and U298 (N_298,N_177,N_106);
and U299 (N_299,In_186,N_82);
and U300 (N_300,N_2,In_16);
nor U301 (N_301,In_353,In_190);
or U302 (N_302,N_131,N_78);
xor U303 (N_303,N_167,N_34);
xor U304 (N_304,N_189,N_66);
nor U305 (N_305,N_90,In_485);
nand U306 (N_306,In_350,N_68);
nor U307 (N_307,N_193,N_140);
nand U308 (N_308,In_50,In_356);
nand U309 (N_309,N_58,In_340);
nand U310 (N_310,In_168,In_66);
nor U311 (N_311,N_105,In_404);
nand U312 (N_312,N_72,N_35);
nand U313 (N_313,N_124,N_27);
nor U314 (N_314,In_386,N_123);
xor U315 (N_315,N_20,N_50);
nand U316 (N_316,N_156,N_59);
nor U317 (N_317,In_231,N_166);
xnor U318 (N_318,N_96,In_282);
or U319 (N_319,In_48,N_21);
nand U320 (N_320,N_51,N_161);
and U321 (N_321,N_79,In_78);
nor U322 (N_322,N_112,N_186);
and U323 (N_323,N_169,N_119);
and U324 (N_324,N_158,N_5);
xor U325 (N_325,N_44,N_38);
and U326 (N_326,N_57,N_147);
nor U327 (N_327,N_93,In_427);
nand U328 (N_328,In_152,N_133);
and U329 (N_329,N_83,In_328);
nor U330 (N_330,N_12,N_42);
nand U331 (N_331,N_92,N_160);
nand U332 (N_332,N_109,In_197);
or U333 (N_333,In_330,N_151);
nand U334 (N_334,N_3,N_150);
nand U335 (N_335,In_188,N_98);
or U336 (N_336,N_63,N_55);
nand U337 (N_337,N_178,N_39);
nor U338 (N_338,In_362,In_430);
nor U339 (N_339,N_89,In_46);
and U340 (N_340,N_4,In_166);
or U341 (N_341,In_8,N_121);
and U342 (N_342,N_26,In_322);
and U343 (N_343,N_70,N_187);
nor U344 (N_344,N_88,N_110);
and U345 (N_345,N_104,In_388);
nor U346 (N_346,N_162,In_284);
nand U347 (N_347,N_0,N_91);
or U348 (N_348,N_114,N_153);
xnor U349 (N_349,N_62,N_115);
and U350 (N_350,In_56,N_104);
or U351 (N_351,In_163,N_34);
and U352 (N_352,In_127,N_135);
nor U353 (N_353,N_82,In_330);
nor U354 (N_354,N_12,In_384);
or U355 (N_355,N_113,In_66);
xnor U356 (N_356,N_179,N_123);
nand U357 (N_357,N_7,N_162);
or U358 (N_358,N_5,In_78);
or U359 (N_359,In_445,N_99);
nand U360 (N_360,N_93,N_146);
nor U361 (N_361,N_41,N_119);
nor U362 (N_362,N_56,In_142);
or U363 (N_363,N_52,N_181);
nand U364 (N_364,N_64,N_84);
and U365 (N_365,N_164,N_147);
nand U366 (N_366,N_113,N_126);
nand U367 (N_367,N_76,N_105);
xor U368 (N_368,N_68,N_28);
or U369 (N_369,N_74,In_485);
xor U370 (N_370,In_302,In_146);
xor U371 (N_371,In_282,In_328);
nor U372 (N_372,N_98,In_386);
nor U373 (N_373,N_131,N_138);
or U374 (N_374,N_175,N_182);
nand U375 (N_375,In_364,N_93);
and U376 (N_376,In_382,In_188);
nand U377 (N_377,N_0,N_74);
and U378 (N_378,N_10,In_20);
or U379 (N_379,N_83,In_168);
or U380 (N_380,N_168,N_97);
nor U381 (N_381,N_176,N_2);
nand U382 (N_382,N_85,N_39);
nand U383 (N_383,N_182,In_9);
xor U384 (N_384,N_140,In_190);
nand U385 (N_385,N_77,N_131);
and U386 (N_386,N_169,N_52);
nor U387 (N_387,N_30,N_46);
or U388 (N_388,N_32,N_43);
and U389 (N_389,N_98,N_161);
xor U390 (N_390,N_4,N_146);
nand U391 (N_391,N_149,N_125);
nand U392 (N_392,In_227,In_41);
nor U393 (N_393,N_124,N_153);
xor U394 (N_394,In_330,N_146);
nand U395 (N_395,N_117,N_134);
xnor U396 (N_396,In_221,In_125);
xor U397 (N_397,N_1,In_382);
and U398 (N_398,In_46,N_167);
and U399 (N_399,N_52,In_20);
or U400 (N_400,N_240,N_205);
or U401 (N_401,N_376,N_301);
and U402 (N_402,N_233,N_356);
or U403 (N_403,N_277,N_334);
nor U404 (N_404,N_299,N_394);
xnor U405 (N_405,N_249,N_278);
or U406 (N_406,N_265,N_257);
nor U407 (N_407,N_369,N_202);
xnor U408 (N_408,N_255,N_262);
and U409 (N_409,N_387,N_384);
and U410 (N_410,N_217,N_361);
nor U411 (N_411,N_309,N_377);
nor U412 (N_412,N_296,N_386);
or U413 (N_413,N_341,N_381);
nand U414 (N_414,N_370,N_312);
nand U415 (N_415,N_360,N_207);
xnor U416 (N_416,N_298,N_342);
nand U417 (N_417,N_297,N_289);
or U418 (N_418,N_317,N_378);
nor U419 (N_419,N_391,N_306);
nand U420 (N_420,N_211,N_285);
nor U421 (N_421,N_243,N_343);
or U422 (N_422,N_208,N_282);
nor U423 (N_423,N_252,N_286);
and U424 (N_424,N_284,N_399);
nor U425 (N_425,N_398,N_396);
xnor U426 (N_426,N_373,N_337);
or U427 (N_427,N_264,N_272);
nor U428 (N_428,N_310,N_215);
or U429 (N_429,N_332,N_273);
or U430 (N_430,N_222,N_328);
nand U431 (N_431,N_220,N_279);
nand U432 (N_432,N_358,N_280);
nand U433 (N_433,N_375,N_340);
nand U434 (N_434,N_379,N_363);
nand U435 (N_435,N_253,N_256);
and U436 (N_436,N_216,N_366);
and U437 (N_437,N_234,N_389);
or U438 (N_438,N_287,N_260);
xnor U439 (N_439,N_364,N_347);
or U440 (N_440,N_271,N_241);
nor U441 (N_441,N_350,N_321);
nand U442 (N_442,N_263,N_380);
nor U443 (N_443,N_248,N_201);
or U444 (N_444,N_314,N_318);
nand U445 (N_445,N_345,N_325);
xnor U446 (N_446,N_275,N_228);
or U447 (N_447,N_242,N_392);
nor U448 (N_448,N_368,N_230);
and U449 (N_449,N_294,N_258);
and U450 (N_450,N_352,N_372);
nor U451 (N_451,N_339,N_238);
and U452 (N_452,N_388,N_266);
and U453 (N_453,N_232,N_357);
and U454 (N_454,N_291,N_393);
nor U455 (N_455,N_212,N_374);
xor U456 (N_456,N_367,N_331);
nor U457 (N_457,N_200,N_307);
xnor U458 (N_458,N_313,N_270);
nand U459 (N_459,N_259,N_290);
or U460 (N_460,N_210,N_204);
nor U461 (N_461,N_371,N_338);
or U462 (N_462,N_326,N_288);
nand U463 (N_463,N_327,N_221);
or U464 (N_464,N_353,N_308);
nor U465 (N_465,N_382,N_333);
and U466 (N_466,N_303,N_349);
xnor U467 (N_467,N_362,N_267);
nor U468 (N_468,N_219,N_274);
or U469 (N_469,N_320,N_229);
nand U470 (N_470,N_223,N_344);
and U471 (N_471,N_330,N_359);
nor U472 (N_472,N_336,N_283);
and U473 (N_473,N_244,N_329);
or U474 (N_474,N_348,N_383);
nor U475 (N_475,N_227,N_335);
nor U476 (N_476,N_246,N_237);
and U477 (N_477,N_292,N_236);
nor U478 (N_478,N_224,N_323);
and U479 (N_479,N_235,N_295);
and U480 (N_480,N_276,N_311);
nand U481 (N_481,N_351,N_316);
and U482 (N_482,N_305,N_322);
nand U483 (N_483,N_213,N_251);
nand U484 (N_484,N_395,N_269);
xnor U485 (N_485,N_300,N_390);
or U486 (N_486,N_304,N_203);
nand U487 (N_487,N_261,N_293);
xnor U488 (N_488,N_254,N_245);
nor U489 (N_489,N_250,N_397);
or U490 (N_490,N_206,N_209);
nand U491 (N_491,N_281,N_355);
xor U492 (N_492,N_231,N_302);
or U493 (N_493,N_218,N_239);
nor U494 (N_494,N_225,N_365);
and U495 (N_495,N_214,N_346);
or U496 (N_496,N_324,N_315);
nor U497 (N_497,N_247,N_268);
nor U498 (N_498,N_226,N_319);
nor U499 (N_499,N_354,N_385);
and U500 (N_500,N_355,N_363);
nor U501 (N_501,N_239,N_203);
nor U502 (N_502,N_203,N_330);
or U503 (N_503,N_279,N_293);
and U504 (N_504,N_375,N_304);
nand U505 (N_505,N_264,N_337);
nand U506 (N_506,N_330,N_293);
nand U507 (N_507,N_233,N_299);
nand U508 (N_508,N_296,N_250);
or U509 (N_509,N_259,N_303);
or U510 (N_510,N_388,N_281);
nand U511 (N_511,N_329,N_350);
nand U512 (N_512,N_307,N_242);
or U513 (N_513,N_371,N_386);
xnor U514 (N_514,N_275,N_391);
and U515 (N_515,N_325,N_239);
nand U516 (N_516,N_264,N_202);
and U517 (N_517,N_228,N_330);
nor U518 (N_518,N_378,N_303);
and U519 (N_519,N_243,N_396);
and U520 (N_520,N_264,N_200);
or U521 (N_521,N_251,N_212);
and U522 (N_522,N_299,N_334);
nand U523 (N_523,N_284,N_369);
nor U524 (N_524,N_240,N_329);
or U525 (N_525,N_298,N_236);
or U526 (N_526,N_321,N_339);
nand U527 (N_527,N_254,N_375);
nand U528 (N_528,N_293,N_324);
or U529 (N_529,N_220,N_367);
xor U530 (N_530,N_246,N_397);
nor U531 (N_531,N_345,N_269);
nand U532 (N_532,N_218,N_263);
nand U533 (N_533,N_335,N_360);
and U534 (N_534,N_267,N_374);
xnor U535 (N_535,N_354,N_275);
xor U536 (N_536,N_219,N_367);
nor U537 (N_537,N_276,N_388);
nand U538 (N_538,N_286,N_292);
xor U539 (N_539,N_263,N_307);
nor U540 (N_540,N_328,N_228);
or U541 (N_541,N_336,N_252);
nand U542 (N_542,N_337,N_303);
and U543 (N_543,N_214,N_261);
nand U544 (N_544,N_338,N_226);
nand U545 (N_545,N_218,N_209);
nor U546 (N_546,N_321,N_271);
nand U547 (N_547,N_249,N_216);
or U548 (N_548,N_287,N_353);
nor U549 (N_549,N_282,N_362);
xor U550 (N_550,N_222,N_209);
and U551 (N_551,N_295,N_330);
nor U552 (N_552,N_324,N_306);
nor U553 (N_553,N_368,N_276);
or U554 (N_554,N_342,N_223);
and U555 (N_555,N_231,N_362);
and U556 (N_556,N_205,N_226);
and U557 (N_557,N_269,N_285);
and U558 (N_558,N_312,N_384);
or U559 (N_559,N_219,N_361);
or U560 (N_560,N_295,N_335);
or U561 (N_561,N_212,N_245);
or U562 (N_562,N_233,N_385);
nand U563 (N_563,N_274,N_276);
or U564 (N_564,N_205,N_333);
xor U565 (N_565,N_259,N_279);
xnor U566 (N_566,N_384,N_221);
nor U567 (N_567,N_309,N_342);
and U568 (N_568,N_248,N_353);
nand U569 (N_569,N_292,N_361);
nor U570 (N_570,N_301,N_362);
nand U571 (N_571,N_384,N_263);
and U572 (N_572,N_345,N_389);
nor U573 (N_573,N_356,N_247);
or U574 (N_574,N_383,N_322);
nand U575 (N_575,N_250,N_272);
and U576 (N_576,N_210,N_339);
nand U577 (N_577,N_324,N_390);
nand U578 (N_578,N_330,N_223);
and U579 (N_579,N_354,N_327);
or U580 (N_580,N_207,N_316);
and U581 (N_581,N_387,N_335);
nand U582 (N_582,N_292,N_297);
nand U583 (N_583,N_249,N_275);
xor U584 (N_584,N_386,N_331);
xor U585 (N_585,N_256,N_383);
nand U586 (N_586,N_245,N_210);
and U587 (N_587,N_370,N_358);
or U588 (N_588,N_221,N_289);
nor U589 (N_589,N_267,N_298);
nand U590 (N_590,N_218,N_203);
or U591 (N_591,N_262,N_395);
and U592 (N_592,N_221,N_391);
xor U593 (N_593,N_247,N_362);
or U594 (N_594,N_300,N_307);
xor U595 (N_595,N_267,N_256);
and U596 (N_596,N_268,N_261);
or U597 (N_597,N_384,N_326);
and U598 (N_598,N_218,N_368);
nand U599 (N_599,N_240,N_272);
or U600 (N_600,N_539,N_471);
or U601 (N_601,N_401,N_508);
nor U602 (N_602,N_467,N_547);
or U603 (N_603,N_543,N_469);
and U604 (N_604,N_589,N_512);
nand U605 (N_605,N_492,N_534);
and U606 (N_606,N_504,N_519);
and U607 (N_607,N_556,N_437);
nor U608 (N_608,N_483,N_551);
or U609 (N_609,N_456,N_497);
nand U610 (N_610,N_453,N_515);
and U611 (N_611,N_489,N_536);
nand U612 (N_612,N_465,N_540);
or U613 (N_613,N_413,N_448);
nand U614 (N_614,N_546,N_440);
and U615 (N_615,N_498,N_501);
or U616 (N_616,N_499,N_578);
nand U617 (N_617,N_463,N_407);
or U618 (N_618,N_435,N_550);
nand U619 (N_619,N_445,N_466);
and U620 (N_620,N_464,N_450);
or U621 (N_621,N_532,N_549);
nor U622 (N_622,N_455,N_449);
and U623 (N_623,N_416,N_461);
and U624 (N_624,N_487,N_502);
or U625 (N_625,N_484,N_475);
and U626 (N_626,N_506,N_432);
and U627 (N_627,N_422,N_439);
xnor U628 (N_628,N_429,N_485);
nand U629 (N_629,N_554,N_414);
nor U630 (N_630,N_548,N_518);
xnor U631 (N_631,N_470,N_477);
nand U632 (N_632,N_482,N_562);
nand U633 (N_633,N_565,N_421);
nand U634 (N_634,N_509,N_412);
nor U635 (N_635,N_577,N_468);
nor U636 (N_636,N_527,N_496);
or U637 (N_637,N_472,N_520);
or U638 (N_638,N_410,N_528);
xor U639 (N_639,N_579,N_598);
nor U640 (N_640,N_402,N_553);
or U641 (N_641,N_571,N_516);
and U642 (N_642,N_529,N_507);
nand U643 (N_643,N_561,N_573);
or U644 (N_644,N_576,N_428);
or U645 (N_645,N_533,N_493);
or U646 (N_646,N_503,N_490);
and U647 (N_647,N_521,N_405);
and U648 (N_648,N_486,N_426);
nand U649 (N_649,N_481,N_434);
and U650 (N_650,N_542,N_593);
xnor U651 (N_651,N_411,N_535);
or U652 (N_652,N_591,N_569);
and U653 (N_653,N_478,N_587);
nand U654 (N_654,N_473,N_403);
nor U655 (N_655,N_572,N_599);
nand U656 (N_656,N_566,N_457);
xor U657 (N_657,N_526,N_552);
and U658 (N_658,N_530,N_415);
and U659 (N_659,N_418,N_537);
nand U660 (N_660,N_424,N_558);
nor U661 (N_661,N_568,N_594);
nand U662 (N_662,N_458,N_560);
nor U663 (N_663,N_523,N_581);
xnor U664 (N_664,N_557,N_592);
nand U665 (N_665,N_479,N_408);
or U666 (N_666,N_524,N_531);
nor U667 (N_667,N_417,N_505);
nand U668 (N_668,N_442,N_425);
xor U669 (N_669,N_511,N_513);
or U670 (N_670,N_419,N_420);
and U671 (N_671,N_588,N_559);
nand U672 (N_672,N_541,N_454);
and U673 (N_673,N_596,N_446);
nand U674 (N_674,N_474,N_480);
nand U675 (N_675,N_491,N_514);
nand U676 (N_676,N_582,N_404);
or U677 (N_677,N_430,N_431);
or U678 (N_678,N_563,N_476);
nor U679 (N_679,N_575,N_436);
nor U680 (N_680,N_400,N_522);
or U681 (N_681,N_545,N_488);
and U682 (N_682,N_495,N_441);
and U683 (N_683,N_459,N_586);
nor U684 (N_684,N_590,N_409);
nor U685 (N_685,N_517,N_597);
or U686 (N_686,N_447,N_544);
nand U687 (N_687,N_570,N_406);
or U688 (N_688,N_574,N_462);
and U689 (N_689,N_443,N_580);
or U690 (N_690,N_510,N_423);
nand U691 (N_691,N_494,N_585);
and U692 (N_692,N_583,N_595);
xor U693 (N_693,N_451,N_564);
nand U694 (N_694,N_538,N_500);
nand U695 (N_695,N_555,N_584);
nor U696 (N_696,N_433,N_427);
or U697 (N_697,N_452,N_438);
nor U698 (N_698,N_460,N_444);
xor U699 (N_699,N_525,N_567);
nand U700 (N_700,N_585,N_481);
xor U701 (N_701,N_473,N_496);
and U702 (N_702,N_574,N_552);
or U703 (N_703,N_408,N_464);
xor U704 (N_704,N_411,N_564);
and U705 (N_705,N_511,N_516);
nor U706 (N_706,N_463,N_532);
nand U707 (N_707,N_456,N_401);
and U708 (N_708,N_540,N_406);
nor U709 (N_709,N_450,N_497);
nand U710 (N_710,N_458,N_585);
and U711 (N_711,N_534,N_432);
nor U712 (N_712,N_513,N_571);
or U713 (N_713,N_492,N_589);
or U714 (N_714,N_559,N_465);
or U715 (N_715,N_419,N_516);
xnor U716 (N_716,N_508,N_587);
nor U717 (N_717,N_442,N_423);
nand U718 (N_718,N_449,N_448);
xor U719 (N_719,N_467,N_457);
nor U720 (N_720,N_443,N_560);
or U721 (N_721,N_411,N_581);
nor U722 (N_722,N_480,N_549);
and U723 (N_723,N_516,N_505);
and U724 (N_724,N_475,N_494);
and U725 (N_725,N_566,N_406);
and U726 (N_726,N_588,N_498);
nand U727 (N_727,N_587,N_586);
or U728 (N_728,N_537,N_405);
or U729 (N_729,N_488,N_406);
nor U730 (N_730,N_478,N_549);
nand U731 (N_731,N_567,N_452);
or U732 (N_732,N_446,N_512);
xor U733 (N_733,N_408,N_543);
or U734 (N_734,N_534,N_444);
nor U735 (N_735,N_480,N_496);
or U736 (N_736,N_569,N_433);
nand U737 (N_737,N_408,N_534);
nand U738 (N_738,N_446,N_563);
and U739 (N_739,N_532,N_455);
or U740 (N_740,N_582,N_405);
and U741 (N_741,N_415,N_571);
or U742 (N_742,N_565,N_510);
nor U743 (N_743,N_458,N_545);
or U744 (N_744,N_477,N_570);
xnor U745 (N_745,N_431,N_536);
nand U746 (N_746,N_425,N_542);
or U747 (N_747,N_403,N_423);
or U748 (N_748,N_475,N_456);
xnor U749 (N_749,N_505,N_584);
nand U750 (N_750,N_504,N_455);
nor U751 (N_751,N_406,N_413);
nand U752 (N_752,N_429,N_563);
nand U753 (N_753,N_466,N_412);
nor U754 (N_754,N_408,N_519);
nand U755 (N_755,N_569,N_595);
nor U756 (N_756,N_458,N_450);
nor U757 (N_757,N_422,N_507);
nor U758 (N_758,N_576,N_591);
nand U759 (N_759,N_593,N_504);
nor U760 (N_760,N_422,N_425);
nand U761 (N_761,N_541,N_570);
xor U762 (N_762,N_530,N_596);
or U763 (N_763,N_481,N_510);
or U764 (N_764,N_502,N_419);
nor U765 (N_765,N_577,N_594);
or U766 (N_766,N_492,N_592);
and U767 (N_767,N_566,N_471);
nand U768 (N_768,N_445,N_590);
xor U769 (N_769,N_504,N_569);
or U770 (N_770,N_502,N_441);
and U771 (N_771,N_445,N_430);
nor U772 (N_772,N_447,N_445);
and U773 (N_773,N_435,N_499);
nand U774 (N_774,N_555,N_540);
and U775 (N_775,N_528,N_513);
nor U776 (N_776,N_586,N_548);
nor U777 (N_777,N_500,N_598);
and U778 (N_778,N_503,N_564);
and U779 (N_779,N_437,N_515);
xor U780 (N_780,N_541,N_400);
or U781 (N_781,N_552,N_461);
or U782 (N_782,N_412,N_536);
and U783 (N_783,N_571,N_494);
and U784 (N_784,N_549,N_533);
nor U785 (N_785,N_472,N_538);
nand U786 (N_786,N_535,N_445);
xor U787 (N_787,N_439,N_521);
and U788 (N_788,N_594,N_449);
or U789 (N_789,N_504,N_475);
nor U790 (N_790,N_528,N_555);
nand U791 (N_791,N_474,N_484);
nand U792 (N_792,N_421,N_456);
nor U793 (N_793,N_401,N_448);
and U794 (N_794,N_554,N_574);
nand U795 (N_795,N_521,N_484);
nor U796 (N_796,N_544,N_415);
xnor U797 (N_797,N_444,N_425);
xor U798 (N_798,N_589,N_480);
and U799 (N_799,N_523,N_585);
or U800 (N_800,N_790,N_651);
nand U801 (N_801,N_799,N_603);
nand U802 (N_802,N_668,N_662);
nand U803 (N_803,N_696,N_664);
or U804 (N_804,N_766,N_618);
nor U805 (N_805,N_638,N_627);
xor U806 (N_806,N_713,N_666);
or U807 (N_807,N_770,N_785);
nand U808 (N_808,N_721,N_763);
xor U809 (N_809,N_743,N_680);
nor U810 (N_810,N_748,N_720);
nor U811 (N_811,N_742,N_728);
nand U812 (N_812,N_787,N_739);
xnor U813 (N_813,N_635,N_736);
nor U814 (N_814,N_794,N_671);
nor U815 (N_815,N_726,N_754);
nor U816 (N_816,N_774,N_789);
nand U817 (N_817,N_791,N_777);
nor U818 (N_818,N_675,N_780);
nand U819 (N_819,N_692,N_691);
and U820 (N_820,N_768,N_765);
nand U821 (N_821,N_631,N_628);
xnor U822 (N_822,N_712,N_673);
or U823 (N_823,N_606,N_633);
and U824 (N_824,N_601,N_613);
or U825 (N_825,N_687,N_672);
nor U826 (N_826,N_661,N_655);
nor U827 (N_827,N_650,N_667);
nand U828 (N_828,N_756,N_632);
and U829 (N_829,N_641,N_795);
and U830 (N_830,N_622,N_630);
and U831 (N_831,N_783,N_644);
nand U832 (N_832,N_750,N_683);
and U833 (N_833,N_718,N_733);
and U834 (N_834,N_698,N_634);
xor U835 (N_835,N_620,N_693);
xor U836 (N_836,N_663,N_652);
xnor U837 (N_837,N_615,N_719);
nand U838 (N_838,N_647,N_772);
and U839 (N_839,N_679,N_788);
and U840 (N_840,N_600,N_643);
xor U841 (N_841,N_755,N_796);
nand U842 (N_842,N_769,N_752);
xnor U843 (N_843,N_625,N_745);
or U844 (N_844,N_757,N_705);
and U845 (N_845,N_686,N_674);
and U846 (N_846,N_729,N_751);
nor U847 (N_847,N_759,N_708);
nor U848 (N_848,N_732,N_731);
nand U849 (N_849,N_709,N_704);
or U850 (N_850,N_798,N_792);
and U851 (N_851,N_747,N_706);
nand U852 (N_852,N_699,N_670);
and U853 (N_853,N_734,N_658);
xnor U854 (N_854,N_730,N_694);
nand U855 (N_855,N_681,N_677);
or U856 (N_856,N_727,N_659);
xnor U857 (N_857,N_758,N_778);
or U858 (N_858,N_797,N_689);
or U859 (N_859,N_612,N_723);
nand U860 (N_860,N_646,N_660);
xnor U861 (N_861,N_724,N_609);
nand U862 (N_862,N_657,N_623);
xnor U863 (N_863,N_654,N_746);
nand U864 (N_864,N_775,N_707);
nand U865 (N_865,N_669,N_678);
or U866 (N_866,N_716,N_614);
nor U867 (N_867,N_610,N_793);
and U868 (N_868,N_741,N_722);
and U869 (N_869,N_702,N_771);
nor U870 (N_870,N_784,N_607);
nor U871 (N_871,N_640,N_715);
or U872 (N_872,N_636,N_786);
nand U873 (N_873,N_779,N_695);
and U874 (N_874,N_717,N_605);
and U875 (N_875,N_737,N_645);
or U876 (N_876,N_602,N_611);
nor U877 (N_877,N_649,N_749);
nand U878 (N_878,N_776,N_629);
or U879 (N_879,N_781,N_700);
nor U880 (N_880,N_656,N_714);
nand U881 (N_881,N_710,N_608);
nand U882 (N_882,N_617,N_685);
nor U883 (N_883,N_616,N_653);
or U884 (N_884,N_684,N_725);
nor U885 (N_885,N_697,N_624);
nand U886 (N_886,N_703,N_738);
or U887 (N_887,N_676,N_711);
and U888 (N_888,N_740,N_642);
nor U889 (N_889,N_637,N_762);
or U890 (N_890,N_690,N_621);
and U891 (N_891,N_760,N_639);
or U892 (N_892,N_665,N_701);
or U893 (N_893,N_604,N_626);
nand U894 (N_894,N_764,N_782);
nand U895 (N_895,N_753,N_688);
and U896 (N_896,N_761,N_648);
and U897 (N_897,N_682,N_767);
or U898 (N_898,N_744,N_619);
or U899 (N_899,N_773,N_735);
or U900 (N_900,N_783,N_726);
nand U901 (N_901,N_697,N_737);
and U902 (N_902,N_628,N_733);
xor U903 (N_903,N_724,N_628);
nand U904 (N_904,N_613,N_699);
or U905 (N_905,N_653,N_677);
nor U906 (N_906,N_647,N_732);
nand U907 (N_907,N_624,N_635);
or U908 (N_908,N_638,N_745);
or U909 (N_909,N_744,N_607);
and U910 (N_910,N_623,N_704);
nor U911 (N_911,N_729,N_610);
or U912 (N_912,N_779,N_618);
xor U913 (N_913,N_737,N_634);
and U914 (N_914,N_730,N_680);
or U915 (N_915,N_779,N_691);
and U916 (N_916,N_764,N_615);
nand U917 (N_917,N_626,N_671);
or U918 (N_918,N_621,N_622);
and U919 (N_919,N_700,N_756);
nor U920 (N_920,N_613,N_628);
and U921 (N_921,N_672,N_683);
nor U922 (N_922,N_676,N_672);
or U923 (N_923,N_767,N_688);
xnor U924 (N_924,N_721,N_640);
xnor U925 (N_925,N_781,N_612);
nor U926 (N_926,N_748,N_689);
and U927 (N_927,N_656,N_688);
or U928 (N_928,N_737,N_672);
nand U929 (N_929,N_676,N_630);
and U930 (N_930,N_646,N_630);
and U931 (N_931,N_777,N_618);
and U932 (N_932,N_600,N_710);
nor U933 (N_933,N_726,N_684);
nand U934 (N_934,N_765,N_791);
xnor U935 (N_935,N_758,N_652);
or U936 (N_936,N_741,N_651);
nor U937 (N_937,N_673,N_669);
nand U938 (N_938,N_678,N_760);
nor U939 (N_939,N_654,N_763);
nor U940 (N_940,N_733,N_662);
and U941 (N_941,N_799,N_652);
nand U942 (N_942,N_614,N_620);
or U943 (N_943,N_781,N_754);
nor U944 (N_944,N_776,N_703);
nor U945 (N_945,N_662,N_763);
or U946 (N_946,N_646,N_704);
or U947 (N_947,N_793,N_688);
nor U948 (N_948,N_619,N_710);
or U949 (N_949,N_711,N_607);
and U950 (N_950,N_662,N_618);
nand U951 (N_951,N_726,N_748);
or U952 (N_952,N_792,N_769);
xor U953 (N_953,N_775,N_752);
and U954 (N_954,N_627,N_759);
nand U955 (N_955,N_730,N_615);
and U956 (N_956,N_747,N_653);
and U957 (N_957,N_702,N_670);
or U958 (N_958,N_690,N_695);
nand U959 (N_959,N_622,N_624);
or U960 (N_960,N_768,N_785);
xnor U961 (N_961,N_717,N_785);
or U962 (N_962,N_673,N_798);
xor U963 (N_963,N_706,N_746);
and U964 (N_964,N_675,N_688);
xnor U965 (N_965,N_608,N_782);
nand U966 (N_966,N_703,N_672);
nor U967 (N_967,N_724,N_684);
nand U968 (N_968,N_708,N_711);
nor U969 (N_969,N_773,N_636);
xnor U970 (N_970,N_601,N_649);
and U971 (N_971,N_675,N_659);
nor U972 (N_972,N_708,N_600);
nor U973 (N_973,N_785,N_608);
nand U974 (N_974,N_778,N_613);
and U975 (N_975,N_610,N_648);
nor U976 (N_976,N_622,N_626);
nand U977 (N_977,N_754,N_646);
and U978 (N_978,N_730,N_653);
xor U979 (N_979,N_628,N_727);
nor U980 (N_980,N_631,N_646);
nand U981 (N_981,N_657,N_685);
or U982 (N_982,N_707,N_730);
nand U983 (N_983,N_665,N_711);
nor U984 (N_984,N_646,N_612);
nand U985 (N_985,N_675,N_603);
or U986 (N_986,N_671,N_743);
and U987 (N_987,N_605,N_612);
and U988 (N_988,N_724,N_799);
or U989 (N_989,N_706,N_648);
or U990 (N_990,N_719,N_705);
or U991 (N_991,N_689,N_716);
and U992 (N_992,N_710,N_606);
nor U993 (N_993,N_602,N_722);
nand U994 (N_994,N_762,N_732);
nand U995 (N_995,N_719,N_632);
nand U996 (N_996,N_629,N_664);
nor U997 (N_997,N_711,N_613);
xor U998 (N_998,N_609,N_616);
or U999 (N_999,N_656,N_604);
nand U1000 (N_1000,N_979,N_917);
and U1001 (N_1001,N_859,N_897);
or U1002 (N_1002,N_883,N_861);
or U1003 (N_1003,N_830,N_870);
nand U1004 (N_1004,N_912,N_804);
nand U1005 (N_1005,N_879,N_933);
xor U1006 (N_1006,N_927,N_822);
nand U1007 (N_1007,N_821,N_990);
nor U1008 (N_1008,N_940,N_946);
xnor U1009 (N_1009,N_969,N_975);
and U1010 (N_1010,N_824,N_941);
nand U1011 (N_1011,N_867,N_913);
nand U1012 (N_1012,N_828,N_907);
and U1013 (N_1013,N_998,N_832);
and U1014 (N_1014,N_973,N_872);
and U1015 (N_1015,N_928,N_855);
nor U1016 (N_1016,N_947,N_831);
xor U1017 (N_1017,N_955,N_978);
nand U1018 (N_1018,N_962,N_869);
and U1019 (N_1019,N_930,N_838);
nor U1020 (N_1020,N_991,N_891);
or U1021 (N_1021,N_906,N_850);
nor U1022 (N_1022,N_968,N_819);
or U1023 (N_1023,N_890,N_818);
nand U1024 (N_1024,N_915,N_853);
or U1025 (N_1025,N_977,N_842);
or U1026 (N_1026,N_800,N_892);
and U1027 (N_1027,N_984,N_936);
and U1028 (N_1028,N_837,N_888);
nand U1029 (N_1029,N_865,N_988);
and U1030 (N_1030,N_843,N_908);
or U1031 (N_1031,N_812,N_981);
and U1032 (N_1032,N_961,N_847);
xor U1033 (N_1033,N_854,N_881);
and U1034 (N_1034,N_987,N_976);
xor U1035 (N_1035,N_806,N_801);
xor U1036 (N_1036,N_989,N_956);
nor U1037 (N_1037,N_816,N_918);
and U1038 (N_1038,N_809,N_845);
xor U1039 (N_1039,N_937,N_840);
and U1040 (N_1040,N_957,N_885);
and U1041 (N_1041,N_935,N_919);
nor U1042 (N_1042,N_871,N_954);
or U1043 (N_1043,N_810,N_911);
and U1044 (N_1044,N_958,N_894);
nand U1045 (N_1045,N_826,N_993);
nor U1046 (N_1046,N_982,N_959);
or U1047 (N_1047,N_898,N_924);
nand U1048 (N_1048,N_948,N_803);
and U1049 (N_1049,N_802,N_805);
nand U1050 (N_1050,N_916,N_886);
nor U1051 (N_1051,N_932,N_900);
nor U1052 (N_1052,N_972,N_808);
nand U1053 (N_1053,N_903,N_995);
nor U1054 (N_1054,N_971,N_942);
and U1055 (N_1055,N_874,N_905);
nand U1056 (N_1056,N_851,N_852);
and U1057 (N_1057,N_846,N_827);
nand U1058 (N_1058,N_920,N_902);
or U1059 (N_1059,N_960,N_914);
or U1060 (N_1060,N_833,N_943);
and U1061 (N_1061,N_866,N_893);
and U1062 (N_1062,N_967,N_910);
and U1063 (N_1063,N_929,N_844);
nand U1064 (N_1064,N_901,N_952);
or U1065 (N_1065,N_863,N_980);
and U1066 (N_1066,N_899,N_896);
and U1067 (N_1067,N_875,N_953);
and U1068 (N_1068,N_820,N_965);
nand U1069 (N_1069,N_887,N_839);
nand U1070 (N_1070,N_814,N_925);
and U1071 (N_1071,N_882,N_815);
nor U1072 (N_1072,N_868,N_922);
nor U1073 (N_1073,N_841,N_877);
nor U1074 (N_1074,N_873,N_983);
nand U1075 (N_1075,N_966,N_921);
and U1076 (N_1076,N_849,N_950);
and U1077 (N_1077,N_834,N_964);
xnor U1078 (N_1078,N_926,N_974);
and U1079 (N_1079,N_945,N_817);
nor U1080 (N_1080,N_923,N_856);
or U1081 (N_1081,N_857,N_938);
nor U1082 (N_1082,N_876,N_811);
and U1083 (N_1083,N_996,N_986);
nor U1084 (N_1084,N_949,N_939);
or U1085 (N_1085,N_999,N_860);
xnor U1086 (N_1086,N_931,N_835);
nand U1087 (N_1087,N_825,N_934);
nand U1088 (N_1088,N_997,N_992);
and U1089 (N_1089,N_889,N_823);
and U1090 (N_1090,N_904,N_994);
nand U1091 (N_1091,N_985,N_858);
or U1092 (N_1092,N_963,N_944);
and U1093 (N_1093,N_829,N_884);
and U1094 (N_1094,N_951,N_848);
nand U1095 (N_1095,N_895,N_807);
and U1096 (N_1096,N_878,N_864);
nor U1097 (N_1097,N_970,N_909);
or U1098 (N_1098,N_880,N_813);
and U1099 (N_1099,N_862,N_836);
or U1100 (N_1100,N_828,N_929);
xor U1101 (N_1101,N_936,N_883);
or U1102 (N_1102,N_891,N_854);
nor U1103 (N_1103,N_977,N_984);
nor U1104 (N_1104,N_913,N_969);
and U1105 (N_1105,N_910,N_958);
or U1106 (N_1106,N_803,N_931);
and U1107 (N_1107,N_898,N_936);
nor U1108 (N_1108,N_895,N_935);
nand U1109 (N_1109,N_833,N_905);
or U1110 (N_1110,N_878,N_801);
and U1111 (N_1111,N_943,N_968);
and U1112 (N_1112,N_959,N_885);
nand U1113 (N_1113,N_915,N_913);
nand U1114 (N_1114,N_901,N_981);
nor U1115 (N_1115,N_987,N_834);
nand U1116 (N_1116,N_959,N_877);
nand U1117 (N_1117,N_820,N_817);
and U1118 (N_1118,N_920,N_809);
nand U1119 (N_1119,N_911,N_855);
xnor U1120 (N_1120,N_895,N_846);
or U1121 (N_1121,N_996,N_826);
or U1122 (N_1122,N_828,N_843);
nand U1123 (N_1123,N_825,N_891);
xnor U1124 (N_1124,N_808,N_864);
and U1125 (N_1125,N_913,N_827);
and U1126 (N_1126,N_845,N_964);
or U1127 (N_1127,N_818,N_834);
xnor U1128 (N_1128,N_803,N_801);
nor U1129 (N_1129,N_918,N_956);
or U1130 (N_1130,N_886,N_932);
or U1131 (N_1131,N_972,N_897);
xnor U1132 (N_1132,N_821,N_930);
xor U1133 (N_1133,N_852,N_991);
and U1134 (N_1134,N_977,N_970);
or U1135 (N_1135,N_961,N_842);
nand U1136 (N_1136,N_835,N_950);
or U1137 (N_1137,N_853,N_883);
nor U1138 (N_1138,N_864,N_813);
or U1139 (N_1139,N_838,N_867);
nor U1140 (N_1140,N_829,N_927);
or U1141 (N_1141,N_899,N_822);
xnor U1142 (N_1142,N_831,N_997);
or U1143 (N_1143,N_931,N_859);
nand U1144 (N_1144,N_950,N_807);
and U1145 (N_1145,N_943,N_902);
nand U1146 (N_1146,N_818,N_968);
nor U1147 (N_1147,N_806,N_841);
or U1148 (N_1148,N_823,N_902);
nor U1149 (N_1149,N_896,N_861);
nor U1150 (N_1150,N_940,N_971);
xnor U1151 (N_1151,N_883,N_866);
nor U1152 (N_1152,N_961,N_996);
xnor U1153 (N_1153,N_876,N_817);
or U1154 (N_1154,N_974,N_909);
nand U1155 (N_1155,N_854,N_928);
nand U1156 (N_1156,N_807,N_808);
nand U1157 (N_1157,N_911,N_979);
and U1158 (N_1158,N_941,N_958);
and U1159 (N_1159,N_927,N_994);
nand U1160 (N_1160,N_804,N_849);
nand U1161 (N_1161,N_828,N_995);
nor U1162 (N_1162,N_857,N_858);
and U1163 (N_1163,N_951,N_990);
or U1164 (N_1164,N_822,N_829);
or U1165 (N_1165,N_884,N_984);
nand U1166 (N_1166,N_912,N_899);
xor U1167 (N_1167,N_942,N_941);
xnor U1168 (N_1168,N_870,N_833);
or U1169 (N_1169,N_946,N_843);
and U1170 (N_1170,N_809,N_951);
or U1171 (N_1171,N_893,N_945);
or U1172 (N_1172,N_875,N_945);
and U1173 (N_1173,N_846,N_829);
or U1174 (N_1174,N_939,N_892);
nor U1175 (N_1175,N_879,N_961);
nor U1176 (N_1176,N_882,N_957);
nor U1177 (N_1177,N_832,N_887);
or U1178 (N_1178,N_934,N_957);
or U1179 (N_1179,N_978,N_800);
nand U1180 (N_1180,N_970,N_923);
and U1181 (N_1181,N_985,N_855);
or U1182 (N_1182,N_964,N_901);
or U1183 (N_1183,N_939,N_873);
or U1184 (N_1184,N_819,N_994);
or U1185 (N_1185,N_847,N_980);
and U1186 (N_1186,N_857,N_972);
nor U1187 (N_1187,N_983,N_840);
nand U1188 (N_1188,N_912,N_921);
and U1189 (N_1189,N_879,N_963);
and U1190 (N_1190,N_800,N_986);
xor U1191 (N_1191,N_942,N_983);
and U1192 (N_1192,N_805,N_935);
and U1193 (N_1193,N_861,N_928);
nor U1194 (N_1194,N_995,N_818);
or U1195 (N_1195,N_927,N_859);
and U1196 (N_1196,N_915,N_989);
nand U1197 (N_1197,N_982,N_920);
or U1198 (N_1198,N_990,N_887);
or U1199 (N_1199,N_891,N_867);
or U1200 (N_1200,N_1162,N_1049);
and U1201 (N_1201,N_1156,N_1048);
nor U1202 (N_1202,N_1061,N_1131);
nand U1203 (N_1203,N_1003,N_1173);
nand U1204 (N_1204,N_1110,N_1054);
nand U1205 (N_1205,N_1152,N_1118);
nor U1206 (N_1206,N_1033,N_1084);
nor U1207 (N_1207,N_1085,N_1028);
nor U1208 (N_1208,N_1042,N_1143);
nand U1209 (N_1209,N_1171,N_1081);
or U1210 (N_1210,N_1062,N_1023);
and U1211 (N_1211,N_1117,N_1004);
and U1212 (N_1212,N_1080,N_1009);
or U1213 (N_1213,N_1195,N_1198);
or U1214 (N_1214,N_1140,N_1076);
nor U1215 (N_1215,N_1178,N_1130);
nor U1216 (N_1216,N_1000,N_1026);
nand U1217 (N_1217,N_1119,N_1055);
nor U1218 (N_1218,N_1043,N_1176);
nand U1219 (N_1219,N_1116,N_1190);
or U1220 (N_1220,N_1147,N_1005);
or U1221 (N_1221,N_1101,N_1007);
nor U1222 (N_1222,N_1024,N_1107);
nor U1223 (N_1223,N_1070,N_1059);
nor U1224 (N_1224,N_1160,N_1180);
nand U1225 (N_1225,N_1072,N_1077);
or U1226 (N_1226,N_1108,N_1175);
and U1227 (N_1227,N_1006,N_1010);
or U1228 (N_1228,N_1193,N_1057);
xor U1229 (N_1229,N_1058,N_1002);
xnor U1230 (N_1230,N_1078,N_1083);
and U1231 (N_1231,N_1136,N_1090);
or U1232 (N_1232,N_1185,N_1089);
nor U1233 (N_1233,N_1105,N_1188);
and U1234 (N_1234,N_1041,N_1184);
nor U1235 (N_1235,N_1016,N_1050);
nor U1236 (N_1236,N_1031,N_1148);
nand U1237 (N_1237,N_1191,N_1124);
and U1238 (N_1238,N_1121,N_1038);
and U1239 (N_1239,N_1123,N_1027);
or U1240 (N_1240,N_1093,N_1075);
nand U1241 (N_1241,N_1199,N_1164);
nor U1242 (N_1242,N_1096,N_1167);
nand U1243 (N_1243,N_1032,N_1091);
nand U1244 (N_1244,N_1127,N_1145);
nand U1245 (N_1245,N_1040,N_1088);
nor U1246 (N_1246,N_1120,N_1079);
and U1247 (N_1247,N_1071,N_1183);
or U1248 (N_1248,N_1144,N_1019);
xnor U1249 (N_1249,N_1182,N_1053);
and U1250 (N_1250,N_1129,N_1022);
or U1251 (N_1251,N_1068,N_1044);
nand U1252 (N_1252,N_1161,N_1065);
and U1253 (N_1253,N_1150,N_1014);
xnor U1254 (N_1254,N_1039,N_1064);
or U1255 (N_1255,N_1106,N_1138);
nand U1256 (N_1256,N_1149,N_1056);
nand U1257 (N_1257,N_1139,N_1189);
xor U1258 (N_1258,N_1047,N_1034);
xor U1259 (N_1259,N_1151,N_1035);
nand U1260 (N_1260,N_1155,N_1086);
nand U1261 (N_1261,N_1045,N_1114);
and U1262 (N_1262,N_1008,N_1133);
and U1263 (N_1263,N_1017,N_1001);
nor U1264 (N_1264,N_1099,N_1113);
xnor U1265 (N_1265,N_1122,N_1146);
nor U1266 (N_1266,N_1046,N_1128);
and U1267 (N_1267,N_1087,N_1196);
nand U1268 (N_1268,N_1125,N_1170);
xor U1269 (N_1269,N_1095,N_1063);
nor U1270 (N_1270,N_1094,N_1069);
nand U1271 (N_1271,N_1115,N_1154);
and U1272 (N_1272,N_1181,N_1111);
or U1273 (N_1273,N_1174,N_1067);
or U1274 (N_1274,N_1082,N_1011);
or U1275 (N_1275,N_1194,N_1060);
xnor U1276 (N_1276,N_1172,N_1051);
and U1277 (N_1277,N_1073,N_1166);
nand U1278 (N_1278,N_1112,N_1098);
or U1279 (N_1279,N_1126,N_1030);
nand U1280 (N_1280,N_1179,N_1163);
nand U1281 (N_1281,N_1092,N_1192);
nand U1282 (N_1282,N_1100,N_1186);
nor U1283 (N_1283,N_1187,N_1137);
or U1284 (N_1284,N_1157,N_1021);
or U1285 (N_1285,N_1141,N_1102);
nor U1286 (N_1286,N_1012,N_1153);
nand U1287 (N_1287,N_1109,N_1135);
or U1288 (N_1288,N_1074,N_1037);
and U1289 (N_1289,N_1158,N_1134);
and U1290 (N_1290,N_1025,N_1142);
nand U1291 (N_1291,N_1169,N_1029);
or U1292 (N_1292,N_1018,N_1104);
nand U1293 (N_1293,N_1015,N_1197);
nand U1294 (N_1294,N_1036,N_1020);
xor U1295 (N_1295,N_1103,N_1168);
and U1296 (N_1296,N_1177,N_1132);
and U1297 (N_1297,N_1159,N_1097);
or U1298 (N_1298,N_1013,N_1066);
nor U1299 (N_1299,N_1165,N_1052);
nor U1300 (N_1300,N_1131,N_1016);
and U1301 (N_1301,N_1135,N_1075);
or U1302 (N_1302,N_1133,N_1011);
nor U1303 (N_1303,N_1149,N_1041);
or U1304 (N_1304,N_1194,N_1093);
nor U1305 (N_1305,N_1182,N_1181);
nor U1306 (N_1306,N_1032,N_1072);
or U1307 (N_1307,N_1091,N_1059);
or U1308 (N_1308,N_1167,N_1051);
and U1309 (N_1309,N_1000,N_1103);
or U1310 (N_1310,N_1043,N_1077);
nand U1311 (N_1311,N_1020,N_1074);
nand U1312 (N_1312,N_1089,N_1193);
and U1313 (N_1313,N_1094,N_1045);
or U1314 (N_1314,N_1035,N_1056);
nand U1315 (N_1315,N_1171,N_1134);
and U1316 (N_1316,N_1028,N_1037);
or U1317 (N_1317,N_1172,N_1156);
and U1318 (N_1318,N_1172,N_1035);
nor U1319 (N_1319,N_1058,N_1158);
or U1320 (N_1320,N_1172,N_1065);
nand U1321 (N_1321,N_1071,N_1152);
and U1322 (N_1322,N_1060,N_1168);
nor U1323 (N_1323,N_1142,N_1169);
and U1324 (N_1324,N_1096,N_1179);
or U1325 (N_1325,N_1165,N_1070);
nand U1326 (N_1326,N_1121,N_1157);
nand U1327 (N_1327,N_1152,N_1105);
or U1328 (N_1328,N_1114,N_1062);
and U1329 (N_1329,N_1163,N_1196);
nor U1330 (N_1330,N_1022,N_1061);
and U1331 (N_1331,N_1002,N_1174);
nand U1332 (N_1332,N_1125,N_1153);
and U1333 (N_1333,N_1004,N_1059);
nand U1334 (N_1334,N_1124,N_1166);
nor U1335 (N_1335,N_1184,N_1150);
nand U1336 (N_1336,N_1012,N_1174);
nor U1337 (N_1337,N_1139,N_1193);
or U1338 (N_1338,N_1177,N_1040);
or U1339 (N_1339,N_1146,N_1154);
and U1340 (N_1340,N_1040,N_1120);
and U1341 (N_1341,N_1100,N_1079);
or U1342 (N_1342,N_1194,N_1135);
or U1343 (N_1343,N_1019,N_1193);
or U1344 (N_1344,N_1090,N_1005);
nand U1345 (N_1345,N_1052,N_1120);
nand U1346 (N_1346,N_1185,N_1167);
nand U1347 (N_1347,N_1047,N_1118);
or U1348 (N_1348,N_1172,N_1103);
or U1349 (N_1349,N_1156,N_1072);
nor U1350 (N_1350,N_1154,N_1064);
nand U1351 (N_1351,N_1096,N_1070);
nand U1352 (N_1352,N_1053,N_1172);
nor U1353 (N_1353,N_1123,N_1162);
nor U1354 (N_1354,N_1101,N_1159);
nand U1355 (N_1355,N_1074,N_1080);
and U1356 (N_1356,N_1014,N_1072);
nor U1357 (N_1357,N_1043,N_1102);
and U1358 (N_1358,N_1070,N_1119);
nand U1359 (N_1359,N_1101,N_1036);
and U1360 (N_1360,N_1046,N_1066);
or U1361 (N_1361,N_1015,N_1014);
nand U1362 (N_1362,N_1078,N_1075);
and U1363 (N_1363,N_1184,N_1106);
nor U1364 (N_1364,N_1030,N_1040);
xor U1365 (N_1365,N_1063,N_1070);
nor U1366 (N_1366,N_1003,N_1021);
nand U1367 (N_1367,N_1129,N_1161);
nor U1368 (N_1368,N_1119,N_1080);
and U1369 (N_1369,N_1161,N_1017);
nor U1370 (N_1370,N_1147,N_1132);
or U1371 (N_1371,N_1140,N_1025);
nand U1372 (N_1372,N_1193,N_1072);
xnor U1373 (N_1373,N_1181,N_1133);
nand U1374 (N_1374,N_1194,N_1045);
nand U1375 (N_1375,N_1085,N_1001);
and U1376 (N_1376,N_1150,N_1149);
nor U1377 (N_1377,N_1070,N_1102);
nand U1378 (N_1378,N_1106,N_1149);
and U1379 (N_1379,N_1026,N_1118);
or U1380 (N_1380,N_1100,N_1151);
nor U1381 (N_1381,N_1182,N_1054);
nor U1382 (N_1382,N_1046,N_1149);
nand U1383 (N_1383,N_1042,N_1167);
and U1384 (N_1384,N_1152,N_1022);
nand U1385 (N_1385,N_1159,N_1046);
and U1386 (N_1386,N_1095,N_1013);
nand U1387 (N_1387,N_1109,N_1057);
nor U1388 (N_1388,N_1139,N_1081);
nand U1389 (N_1389,N_1120,N_1148);
nand U1390 (N_1390,N_1135,N_1111);
or U1391 (N_1391,N_1182,N_1026);
xnor U1392 (N_1392,N_1142,N_1008);
nand U1393 (N_1393,N_1003,N_1160);
nand U1394 (N_1394,N_1027,N_1164);
nor U1395 (N_1395,N_1114,N_1127);
nand U1396 (N_1396,N_1156,N_1195);
and U1397 (N_1397,N_1051,N_1058);
nor U1398 (N_1398,N_1044,N_1059);
xnor U1399 (N_1399,N_1072,N_1008);
nand U1400 (N_1400,N_1368,N_1397);
nand U1401 (N_1401,N_1239,N_1284);
or U1402 (N_1402,N_1281,N_1370);
nand U1403 (N_1403,N_1264,N_1265);
xnor U1404 (N_1404,N_1396,N_1294);
nor U1405 (N_1405,N_1325,N_1361);
nor U1406 (N_1406,N_1387,N_1324);
nand U1407 (N_1407,N_1214,N_1238);
and U1408 (N_1408,N_1381,N_1274);
nor U1409 (N_1409,N_1316,N_1250);
xor U1410 (N_1410,N_1348,N_1386);
nor U1411 (N_1411,N_1272,N_1300);
nor U1412 (N_1412,N_1280,N_1201);
or U1413 (N_1413,N_1277,N_1352);
nand U1414 (N_1414,N_1353,N_1333);
nand U1415 (N_1415,N_1232,N_1362);
nor U1416 (N_1416,N_1251,N_1234);
nor U1417 (N_1417,N_1295,N_1240);
xnor U1418 (N_1418,N_1221,N_1313);
or U1419 (N_1419,N_1327,N_1303);
nor U1420 (N_1420,N_1395,N_1304);
or U1421 (N_1421,N_1331,N_1377);
or U1422 (N_1422,N_1227,N_1389);
or U1423 (N_1423,N_1311,N_1245);
and U1424 (N_1424,N_1371,N_1243);
nor U1425 (N_1425,N_1342,N_1210);
or U1426 (N_1426,N_1350,N_1322);
and U1427 (N_1427,N_1317,N_1246);
nand U1428 (N_1428,N_1207,N_1205);
and U1429 (N_1429,N_1283,N_1335);
or U1430 (N_1430,N_1261,N_1372);
nor U1431 (N_1431,N_1336,N_1388);
and U1432 (N_1432,N_1218,N_1332);
and U1433 (N_1433,N_1393,N_1259);
or U1434 (N_1434,N_1288,N_1291);
or U1435 (N_1435,N_1321,N_1363);
nor U1436 (N_1436,N_1229,N_1206);
nand U1437 (N_1437,N_1334,N_1209);
nand U1438 (N_1438,N_1219,N_1337);
and U1439 (N_1439,N_1282,N_1262);
nand U1440 (N_1440,N_1223,N_1319);
nor U1441 (N_1441,N_1399,N_1338);
and U1442 (N_1442,N_1326,N_1286);
or U1443 (N_1443,N_1241,N_1297);
and U1444 (N_1444,N_1275,N_1320);
nand U1445 (N_1445,N_1383,N_1345);
and U1446 (N_1446,N_1255,N_1374);
nand U1447 (N_1447,N_1301,N_1365);
nor U1448 (N_1448,N_1236,N_1271);
nand U1449 (N_1449,N_1364,N_1216);
and U1450 (N_1450,N_1252,N_1351);
nand U1451 (N_1451,N_1384,N_1305);
xor U1452 (N_1452,N_1289,N_1314);
nor U1453 (N_1453,N_1228,N_1330);
xor U1454 (N_1454,N_1254,N_1308);
nor U1455 (N_1455,N_1266,N_1248);
or U1456 (N_1456,N_1315,N_1309);
xnor U1457 (N_1457,N_1356,N_1204);
nand U1458 (N_1458,N_1298,N_1285);
and U1459 (N_1459,N_1260,N_1273);
and U1460 (N_1460,N_1390,N_1378);
or U1461 (N_1461,N_1247,N_1222);
nand U1462 (N_1462,N_1341,N_1346);
and U1463 (N_1463,N_1367,N_1257);
nor U1464 (N_1464,N_1318,N_1203);
or U1465 (N_1465,N_1376,N_1385);
and U1466 (N_1466,N_1296,N_1217);
and U1467 (N_1467,N_1230,N_1237);
nor U1468 (N_1468,N_1213,N_1263);
xnor U1469 (N_1469,N_1306,N_1231);
or U1470 (N_1470,N_1310,N_1258);
or U1471 (N_1471,N_1375,N_1242);
nor U1472 (N_1472,N_1358,N_1279);
nor U1473 (N_1473,N_1392,N_1249);
xor U1474 (N_1474,N_1224,N_1200);
xnor U1475 (N_1475,N_1256,N_1349);
xor U1476 (N_1476,N_1270,N_1347);
nor U1477 (N_1477,N_1340,N_1215);
xor U1478 (N_1478,N_1312,N_1369);
nand U1479 (N_1479,N_1226,N_1357);
nor U1480 (N_1480,N_1359,N_1307);
or U1481 (N_1481,N_1344,N_1328);
nor U1482 (N_1482,N_1398,N_1380);
xor U1483 (N_1483,N_1394,N_1366);
nand U1484 (N_1484,N_1323,N_1211);
or U1485 (N_1485,N_1202,N_1379);
xnor U1486 (N_1486,N_1299,N_1278);
nor U1487 (N_1487,N_1220,N_1292);
or U1488 (N_1488,N_1287,N_1212);
and U1489 (N_1489,N_1290,N_1373);
xor U1490 (N_1490,N_1225,N_1276);
or U1491 (N_1491,N_1235,N_1253);
nor U1492 (N_1492,N_1208,N_1329);
or U1493 (N_1493,N_1293,N_1343);
and U1494 (N_1494,N_1268,N_1302);
or U1495 (N_1495,N_1244,N_1269);
or U1496 (N_1496,N_1354,N_1360);
nor U1497 (N_1497,N_1382,N_1391);
xnor U1498 (N_1498,N_1355,N_1339);
or U1499 (N_1499,N_1267,N_1233);
nor U1500 (N_1500,N_1376,N_1336);
and U1501 (N_1501,N_1380,N_1327);
xnor U1502 (N_1502,N_1273,N_1206);
nand U1503 (N_1503,N_1359,N_1333);
nor U1504 (N_1504,N_1233,N_1351);
and U1505 (N_1505,N_1201,N_1396);
and U1506 (N_1506,N_1380,N_1304);
nor U1507 (N_1507,N_1316,N_1334);
nor U1508 (N_1508,N_1286,N_1371);
or U1509 (N_1509,N_1215,N_1394);
nand U1510 (N_1510,N_1243,N_1299);
nor U1511 (N_1511,N_1291,N_1326);
nand U1512 (N_1512,N_1208,N_1217);
nor U1513 (N_1513,N_1283,N_1292);
xnor U1514 (N_1514,N_1302,N_1294);
xor U1515 (N_1515,N_1309,N_1313);
or U1516 (N_1516,N_1275,N_1204);
nand U1517 (N_1517,N_1380,N_1391);
and U1518 (N_1518,N_1316,N_1217);
or U1519 (N_1519,N_1311,N_1231);
xor U1520 (N_1520,N_1327,N_1268);
xor U1521 (N_1521,N_1279,N_1383);
or U1522 (N_1522,N_1390,N_1350);
nor U1523 (N_1523,N_1233,N_1219);
and U1524 (N_1524,N_1252,N_1372);
or U1525 (N_1525,N_1274,N_1340);
or U1526 (N_1526,N_1395,N_1232);
nor U1527 (N_1527,N_1321,N_1385);
or U1528 (N_1528,N_1345,N_1235);
nand U1529 (N_1529,N_1228,N_1332);
xnor U1530 (N_1530,N_1232,N_1294);
or U1531 (N_1531,N_1240,N_1227);
nor U1532 (N_1532,N_1274,N_1339);
or U1533 (N_1533,N_1227,N_1371);
or U1534 (N_1534,N_1321,N_1311);
xor U1535 (N_1535,N_1205,N_1277);
and U1536 (N_1536,N_1341,N_1280);
nor U1537 (N_1537,N_1304,N_1316);
nand U1538 (N_1538,N_1201,N_1298);
xnor U1539 (N_1539,N_1249,N_1345);
xnor U1540 (N_1540,N_1396,N_1229);
nand U1541 (N_1541,N_1260,N_1223);
xor U1542 (N_1542,N_1257,N_1237);
nor U1543 (N_1543,N_1305,N_1234);
nand U1544 (N_1544,N_1326,N_1357);
nor U1545 (N_1545,N_1329,N_1205);
or U1546 (N_1546,N_1304,N_1344);
or U1547 (N_1547,N_1326,N_1265);
and U1548 (N_1548,N_1336,N_1325);
nand U1549 (N_1549,N_1252,N_1277);
or U1550 (N_1550,N_1345,N_1323);
or U1551 (N_1551,N_1205,N_1311);
or U1552 (N_1552,N_1303,N_1215);
and U1553 (N_1553,N_1349,N_1368);
or U1554 (N_1554,N_1367,N_1275);
or U1555 (N_1555,N_1370,N_1378);
nand U1556 (N_1556,N_1226,N_1279);
xnor U1557 (N_1557,N_1233,N_1245);
and U1558 (N_1558,N_1294,N_1309);
xor U1559 (N_1559,N_1233,N_1363);
or U1560 (N_1560,N_1304,N_1274);
nand U1561 (N_1561,N_1390,N_1208);
nand U1562 (N_1562,N_1391,N_1231);
nand U1563 (N_1563,N_1239,N_1365);
nand U1564 (N_1564,N_1317,N_1234);
nand U1565 (N_1565,N_1296,N_1215);
and U1566 (N_1566,N_1341,N_1217);
nor U1567 (N_1567,N_1234,N_1278);
nand U1568 (N_1568,N_1350,N_1394);
nand U1569 (N_1569,N_1396,N_1210);
or U1570 (N_1570,N_1317,N_1239);
nand U1571 (N_1571,N_1349,N_1378);
or U1572 (N_1572,N_1320,N_1353);
and U1573 (N_1573,N_1220,N_1268);
and U1574 (N_1574,N_1369,N_1366);
and U1575 (N_1575,N_1337,N_1205);
nor U1576 (N_1576,N_1328,N_1228);
nor U1577 (N_1577,N_1242,N_1234);
nor U1578 (N_1578,N_1214,N_1280);
or U1579 (N_1579,N_1395,N_1255);
xor U1580 (N_1580,N_1331,N_1226);
xnor U1581 (N_1581,N_1331,N_1370);
or U1582 (N_1582,N_1217,N_1344);
or U1583 (N_1583,N_1314,N_1269);
nand U1584 (N_1584,N_1251,N_1279);
nor U1585 (N_1585,N_1376,N_1333);
nor U1586 (N_1586,N_1231,N_1329);
nand U1587 (N_1587,N_1284,N_1207);
and U1588 (N_1588,N_1240,N_1228);
nor U1589 (N_1589,N_1391,N_1311);
or U1590 (N_1590,N_1209,N_1242);
or U1591 (N_1591,N_1246,N_1337);
or U1592 (N_1592,N_1263,N_1238);
nand U1593 (N_1593,N_1236,N_1295);
xnor U1594 (N_1594,N_1239,N_1381);
nand U1595 (N_1595,N_1283,N_1353);
and U1596 (N_1596,N_1367,N_1201);
xnor U1597 (N_1597,N_1366,N_1370);
nor U1598 (N_1598,N_1323,N_1367);
nand U1599 (N_1599,N_1389,N_1295);
nor U1600 (N_1600,N_1489,N_1581);
xnor U1601 (N_1601,N_1437,N_1404);
or U1602 (N_1602,N_1469,N_1414);
nor U1603 (N_1603,N_1523,N_1506);
and U1604 (N_1604,N_1569,N_1532);
and U1605 (N_1605,N_1521,N_1421);
nand U1606 (N_1606,N_1564,N_1560);
nand U1607 (N_1607,N_1443,N_1471);
xor U1608 (N_1608,N_1552,N_1522);
or U1609 (N_1609,N_1446,N_1490);
nand U1610 (N_1610,N_1500,N_1566);
or U1611 (N_1611,N_1432,N_1586);
or U1612 (N_1612,N_1553,N_1587);
nor U1613 (N_1613,N_1557,N_1418);
nand U1614 (N_1614,N_1538,N_1431);
or U1615 (N_1615,N_1461,N_1579);
or U1616 (N_1616,N_1515,N_1485);
or U1617 (N_1617,N_1424,N_1573);
and U1618 (N_1618,N_1466,N_1595);
and U1619 (N_1619,N_1492,N_1533);
nand U1620 (N_1620,N_1453,N_1462);
and U1621 (N_1621,N_1435,N_1496);
nor U1622 (N_1622,N_1572,N_1436);
nor U1623 (N_1623,N_1537,N_1577);
nand U1624 (N_1624,N_1576,N_1501);
and U1625 (N_1625,N_1513,N_1434);
nand U1626 (N_1626,N_1519,N_1464);
or U1627 (N_1627,N_1530,N_1463);
or U1628 (N_1628,N_1447,N_1561);
and U1629 (N_1629,N_1548,N_1465);
or U1630 (N_1630,N_1508,N_1428);
nor U1631 (N_1631,N_1440,N_1419);
and U1632 (N_1632,N_1547,N_1574);
or U1633 (N_1633,N_1427,N_1535);
nand U1634 (N_1634,N_1512,N_1417);
nor U1635 (N_1635,N_1413,N_1441);
nor U1636 (N_1636,N_1596,N_1438);
nor U1637 (N_1637,N_1531,N_1423);
and U1638 (N_1638,N_1592,N_1481);
nand U1639 (N_1639,N_1470,N_1559);
nor U1640 (N_1640,N_1520,N_1475);
xnor U1641 (N_1641,N_1497,N_1562);
or U1642 (N_1642,N_1402,N_1509);
and U1643 (N_1643,N_1468,N_1477);
or U1644 (N_1644,N_1456,N_1498);
and U1645 (N_1645,N_1433,N_1526);
nand U1646 (N_1646,N_1594,N_1504);
nand U1647 (N_1647,N_1510,N_1426);
xor U1648 (N_1648,N_1529,N_1458);
xnor U1649 (N_1649,N_1478,N_1451);
or U1650 (N_1650,N_1582,N_1439);
and U1651 (N_1651,N_1429,N_1568);
nand U1652 (N_1652,N_1480,N_1400);
xor U1653 (N_1653,N_1597,N_1422);
nand U1654 (N_1654,N_1503,N_1476);
or U1655 (N_1655,N_1405,N_1450);
nand U1656 (N_1656,N_1445,N_1525);
nand U1657 (N_1657,N_1411,N_1407);
nand U1658 (N_1658,N_1543,N_1412);
nand U1659 (N_1659,N_1457,N_1516);
or U1660 (N_1660,N_1449,N_1459);
or U1661 (N_1661,N_1554,N_1416);
nand U1662 (N_1662,N_1565,N_1563);
and U1663 (N_1663,N_1483,N_1408);
nor U1664 (N_1664,N_1585,N_1507);
or U1665 (N_1665,N_1544,N_1495);
nand U1666 (N_1666,N_1420,N_1491);
and U1667 (N_1667,N_1578,N_1590);
nor U1668 (N_1668,N_1486,N_1534);
or U1669 (N_1669,N_1406,N_1545);
and U1670 (N_1670,N_1472,N_1455);
or U1671 (N_1671,N_1502,N_1514);
or U1672 (N_1672,N_1528,N_1415);
and U1673 (N_1673,N_1558,N_1473);
nand U1674 (N_1674,N_1403,N_1484);
nor U1675 (N_1675,N_1588,N_1567);
or U1676 (N_1676,N_1599,N_1401);
nor U1677 (N_1677,N_1410,N_1448);
xnor U1678 (N_1678,N_1430,N_1555);
and U1679 (N_1679,N_1524,N_1546);
nor U1680 (N_1680,N_1580,N_1584);
and U1681 (N_1681,N_1540,N_1539);
and U1682 (N_1682,N_1493,N_1570);
or U1683 (N_1683,N_1593,N_1425);
and U1684 (N_1684,N_1551,N_1549);
and U1685 (N_1685,N_1511,N_1591);
nand U1686 (N_1686,N_1583,N_1474);
or U1687 (N_1687,N_1482,N_1589);
xor U1688 (N_1688,N_1467,N_1494);
or U1689 (N_1689,N_1454,N_1598);
nand U1690 (N_1690,N_1499,N_1517);
and U1691 (N_1691,N_1518,N_1541);
nand U1692 (N_1692,N_1550,N_1527);
and U1693 (N_1693,N_1505,N_1575);
nor U1694 (N_1694,N_1460,N_1452);
nor U1695 (N_1695,N_1409,N_1479);
nor U1696 (N_1696,N_1556,N_1442);
nor U1697 (N_1697,N_1487,N_1488);
nand U1698 (N_1698,N_1542,N_1444);
or U1699 (N_1699,N_1536,N_1571);
nor U1700 (N_1700,N_1537,N_1415);
nor U1701 (N_1701,N_1501,N_1533);
xor U1702 (N_1702,N_1567,N_1461);
nand U1703 (N_1703,N_1468,N_1508);
xor U1704 (N_1704,N_1510,N_1532);
nand U1705 (N_1705,N_1432,N_1434);
nand U1706 (N_1706,N_1450,N_1567);
nor U1707 (N_1707,N_1411,N_1466);
xor U1708 (N_1708,N_1576,N_1423);
and U1709 (N_1709,N_1465,N_1409);
or U1710 (N_1710,N_1485,N_1431);
and U1711 (N_1711,N_1484,N_1450);
nand U1712 (N_1712,N_1566,N_1470);
nand U1713 (N_1713,N_1547,N_1517);
or U1714 (N_1714,N_1586,N_1460);
nand U1715 (N_1715,N_1511,N_1488);
nand U1716 (N_1716,N_1584,N_1461);
xor U1717 (N_1717,N_1483,N_1592);
or U1718 (N_1718,N_1476,N_1498);
and U1719 (N_1719,N_1453,N_1476);
and U1720 (N_1720,N_1535,N_1475);
xor U1721 (N_1721,N_1572,N_1434);
or U1722 (N_1722,N_1497,N_1597);
and U1723 (N_1723,N_1425,N_1439);
or U1724 (N_1724,N_1456,N_1566);
and U1725 (N_1725,N_1407,N_1431);
or U1726 (N_1726,N_1542,N_1501);
nor U1727 (N_1727,N_1496,N_1540);
nand U1728 (N_1728,N_1560,N_1430);
nor U1729 (N_1729,N_1503,N_1487);
or U1730 (N_1730,N_1490,N_1406);
or U1731 (N_1731,N_1506,N_1539);
and U1732 (N_1732,N_1517,N_1455);
or U1733 (N_1733,N_1594,N_1456);
and U1734 (N_1734,N_1430,N_1540);
or U1735 (N_1735,N_1410,N_1561);
or U1736 (N_1736,N_1492,N_1567);
nor U1737 (N_1737,N_1448,N_1492);
nor U1738 (N_1738,N_1525,N_1581);
nand U1739 (N_1739,N_1550,N_1448);
and U1740 (N_1740,N_1567,N_1423);
and U1741 (N_1741,N_1514,N_1582);
nor U1742 (N_1742,N_1407,N_1474);
xnor U1743 (N_1743,N_1405,N_1505);
or U1744 (N_1744,N_1490,N_1456);
nand U1745 (N_1745,N_1570,N_1590);
xor U1746 (N_1746,N_1483,N_1597);
xnor U1747 (N_1747,N_1594,N_1488);
xnor U1748 (N_1748,N_1434,N_1510);
nor U1749 (N_1749,N_1592,N_1412);
nand U1750 (N_1750,N_1565,N_1548);
and U1751 (N_1751,N_1562,N_1511);
xnor U1752 (N_1752,N_1427,N_1542);
and U1753 (N_1753,N_1486,N_1580);
xnor U1754 (N_1754,N_1490,N_1553);
and U1755 (N_1755,N_1571,N_1561);
xnor U1756 (N_1756,N_1592,N_1519);
xor U1757 (N_1757,N_1444,N_1426);
nand U1758 (N_1758,N_1527,N_1580);
nor U1759 (N_1759,N_1440,N_1581);
nand U1760 (N_1760,N_1499,N_1407);
or U1761 (N_1761,N_1416,N_1580);
xor U1762 (N_1762,N_1472,N_1489);
xnor U1763 (N_1763,N_1488,N_1430);
and U1764 (N_1764,N_1422,N_1488);
xor U1765 (N_1765,N_1546,N_1498);
nand U1766 (N_1766,N_1416,N_1500);
xor U1767 (N_1767,N_1518,N_1468);
nand U1768 (N_1768,N_1431,N_1522);
nor U1769 (N_1769,N_1496,N_1596);
nand U1770 (N_1770,N_1454,N_1453);
or U1771 (N_1771,N_1467,N_1408);
or U1772 (N_1772,N_1477,N_1483);
nand U1773 (N_1773,N_1535,N_1500);
xor U1774 (N_1774,N_1458,N_1419);
nand U1775 (N_1775,N_1578,N_1585);
xnor U1776 (N_1776,N_1446,N_1599);
and U1777 (N_1777,N_1507,N_1454);
nand U1778 (N_1778,N_1413,N_1581);
or U1779 (N_1779,N_1543,N_1496);
nor U1780 (N_1780,N_1454,N_1488);
xor U1781 (N_1781,N_1488,N_1514);
or U1782 (N_1782,N_1566,N_1520);
nor U1783 (N_1783,N_1423,N_1503);
nor U1784 (N_1784,N_1583,N_1526);
nand U1785 (N_1785,N_1570,N_1475);
or U1786 (N_1786,N_1484,N_1591);
xor U1787 (N_1787,N_1537,N_1592);
nand U1788 (N_1788,N_1412,N_1485);
nor U1789 (N_1789,N_1506,N_1422);
nand U1790 (N_1790,N_1516,N_1445);
and U1791 (N_1791,N_1565,N_1569);
and U1792 (N_1792,N_1431,N_1457);
nand U1793 (N_1793,N_1502,N_1471);
and U1794 (N_1794,N_1527,N_1493);
nor U1795 (N_1795,N_1416,N_1465);
or U1796 (N_1796,N_1584,N_1426);
or U1797 (N_1797,N_1591,N_1482);
nor U1798 (N_1798,N_1417,N_1502);
or U1799 (N_1799,N_1568,N_1575);
or U1800 (N_1800,N_1797,N_1677);
or U1801 (N_1801,N_1627,N_1744);
nor U1802 (N_1802,N_1661,N_1723);
or U1803 (N_1803,N_1764,N_1650);
or U1804 (N_1804,N_1630,N_1607);
and U1805 (N_1805,N_1737,N_1732);
nand U1806 (N_1806,N_1686,N_1740);
nand U1807 (N_1807,N_1705,N_1711);
nand U1808 (N_1808,N_1758,N_1713);
or U1809 (N_1809,N_1783,N_1657);
or U1810 (N_1810,N_1785,N_1731);
and U1811 (N_1811,N_1793,N_1761);
nor U1812 (N_1812,N_1605,N_1707);
or U1813 (N_1813,N_1695,N_1739);
xor U1814 (N_1814,N_1609,N_1610);
nand U1815 (N_1815,N_1690,N_1637);
or U1816 (N_1816,N_1670,N_1694);
nand U1817 (N_1817,N_1666,N_1780);
and U1818 (N_1818,N_1614,N_1619);
nand U1819 (N_1819,N_1623,N_1682);
nor U1820 (N_1820,N_1645,N_1617);
xnor U1821 (N_1821,N_1728,N_1791);
nand U1822 (N_1822,N_1691,N_1699);
and U1823 (N_1823,N_1628,N_1649);
xnor U1824 (N_1824,N_1778,N_1646);
or U1825 (N_1825,N_1712,N_1678);
or U1826 (N_1826,N_1684,N_1603);
or U1827 (N_1827,N_1715,N_1643);
or U1828 (N_1828,N_1710,N_1719);
nand U1829 (N_1829,N_1716,N_1629);
nor U1830 (N_1830,N_1671,N_1679);
and U1831 (N_1831,N_1773,N_1796);
and U1832 (N_1832,N_1634,N_1620);
or U1833 (N_1833,N_1784,N_1703);
nor U1834 (N_1834,N_1604,N_1786);
and U1835 (N_1835,N_1751,N_1743);
nor U1836 (N_1836,N_1663,N_1633);
nor U1837 (N_1837,N_1790,N_1748);
nand U1838 (N_1838,N_1681,N_1789);
xnor U1839 (N_1839,N_1706,N_1641);
or U1840 (N_1840,N_1722,N_1729);
nand U1841 (N_1841,N_1704,N_1765);
nand U1842 (N_1842,N_1733,N_1745);
nor U1843 (N_1843,N_1755,N_1769);
and U1844 (N_1844,N_1798,N_1753);
nand U1845 (N_1845,N_1611,N_1680);
and U1846 (N_1846,N_1652,N_1763);
and U1847 (N_1847,N_1792,N_1606);
nand U1848 (N_1848,N_1735,N_1782);
and U1849 (N_1849,N_1726,N_1701);
nand U1850 (N_1850,N_1613,N_1777);
nor U1851 (N_1851,N_1766,N_1647);
and U1852 (N_1852,N_1635,N_1659);
and U1853 (N_1853,N_1781,N_1741);
nor U1854 (N_1854,N_1724,N_1721);
nor U1855 (N_1855,N_1602,N_1616);
or U1856 (N_1856,N_1717,N_1709);
and U1857 (N_1857,N_1655,N_1720);
nor U1858 (N_1858,N_1654,N_1693);
xnor U1859 (N_1859,N_1636,N_1752);
nor U1860 (N_1860,N_1759,N_1618);
and U1861 (N_1861,N_1658,N_1794);
nor U1862 (N_1862,N_1668,N_1696);
nor U1863 (N_1863,N_1676,N_1688);
or U1864 (N_1864,N_1644,N_1767);
nor U1865 (N_1865,N_1600,N_1775);
nor U1866 (N_1866,N_1714,N_1612);
nor U1867 (N_1867,N_1648,N_1700);
nand U1868 (N_1868,N_1626,N_1673);
nor U1869 (N_1869,N_1795,N_1738);
and U1870 (N_1870,N_1687,N_1674);
nor U1871 (N_1871,N_1669,N_1656);
nor U1872 (N_1872,N_1750,N_1698);
nor U1873 (N_1873,N_1651,N_1702);
and U1874 (N_1874,N_1725,N_1754);
and U1875 (N_1875,N_1760,N_1697);
and U1876 (N_1876,N_1771,N_1736);
nor U1877 (N_1877,N_1727,N_1757);
or U1878 (N_1878,N_1640,N_1770);
and U1879 (N_1879,N_1692,N_1718);
and U1880 (N_1880,N_1787,N_1730);
or U1881 (N_1881,N_1624,N_1746);
nor U1882 (N_1882,N_1660,N_1734);
nand U1883 (N_1883,N_1756,N_1776);
and U1884 (N_1884,N_1642,N_1762);
or U1885 (N_1885,N_1742,N_1708);
or U1886 (N_1886,N_1689,N_1638);
nand U1887 (N_1887,N_1747,N_1685);
nor U1888 (N_1888,N_1625,N_1774);
xor U1889 (N_1889,N_1675,N_1639);
and U1890 (N_1890,N_1662,N_1665);
xor U1891 (N_1891,N_1608,N_1768);
and U1892 (N_1892,N_1601,N_1621);
nand U1893 (N_1893,N_1632,N_1672);
or U1894 (N_1894,N_1615,N_1622);
nor U1895 (N_1895,N_1779,N_1799);
nand U1896 (N_1896,N_1653,N_1683);
and U1897 (N_1897,N_1788,N_1667);
and U1898 (N_1898,N_1664,N_1772);
and U1899 (N_1899,N_1631,N_1749);
nor U1900 (N_1900,N_1661,N_1645);
or U1901 (N_1901,N_1788,N_1763);
nor U1902 (N_1902,N_1620,N_1703);
and U1903 (N_1903,N_1777,N_1647);
nand U1904 (N_1904,N_1769,N_1643);
nand U1905 (N_1905,N_1626,N_1757);
nand U1906 (N_1906,N_1630,N_1709);
nor U1907 (N_1907,N_1698,N_1733);
or U1908 (N_1908,N_1784,N_1735);
nor U1909 (N_1909,N_1730,N_1799);
nand U1910 (N_1910,N_1623,N_1725);
nor U1911 (N_1911,N_1663,N_1740);
nor U1912 (N_1912,N_1678,N_1650);
and U1913 (N_1913,N_1619,N_1759);
xor U1914 (N_1914,N_1721,N_1774);
or U1915 (N_1915,N_1756,N_1615);
nor U1916 (N_1916,N_1755,N_1635);
nand U1917 (N_1917,N_1759,N_1641);
or U1918 (N_1918,N_1726,N_1747);
nand U1919 (N_1919,N_1622,N_1695);
and U1920 (N_1920,N_1613,N_1728);
and U1921 (N_1921,N_1704,N_1605);
nor U1922 (N_1922,N_1701,N_1720);
and U1923 (N_1923,N_1726,N_1684);
xnor U1924 (N_1924,N_1611,N_1796);
nor U1925 (N_1925,N_1664,N_1661);
nor U1926 (N_1926,N_1706,N_1788);
or U1927 (N_1927,N_1704,N_1600);
or U1928 (N_1928,N_1606,N_1719);
and U1929 (N_1929,N_1723,N_1604);
nor U1930 (N_1930,N_1772,N_1649);
nor U1931 (N_1931,N_1772,N_1728);
nand U1932 (N_1932,N_1718,N_1634);
nand U1933 (N_1933,N_1797,N_1622);
or U1934 (N_1934,N_1630,N_1664);
nand U1935 (N_1935,N_1789,N_1799);
or U1936 (N_1936,N_1731,N_1740);
or U1937 (N_1937,N_1639,N_1646);
or U1938 (N_1938,N_1794,N_1714);
or U1939 (N_1939,N_1662,N_1681);
xnor U1940 (N_1940,N_1780,N_1728);
and U1941 (N_1941,N_1776,N_1740);
nor U1942 (N_1942,N_1731,N_1631);
nor U1943 (N_1943,N_1640,N_1719);
xor U1944 (N_1944,N_1629,N_1686);
nor U1945 (N_1945,N_1745,N_1688);
and U1946 (N_1946,N_1736,N_1606);
and U1947 (N_1947,N_1786,N_1764);
xnor U1948 (N_1948,N_1790,N_1727);
xnor U1949 (N_1949,N_1630,N_1632);
nand U1950 (N_1950,N_1678,N_1626);
nand U1951 (N_1951,N_1711,N_1776);
nor U1952 (N_1952,N_1612,N_1776);
and U1953 (N_1953,N_1658,N_1753);
nor U1954 (N_1954,N_1606,N_1709);
and U1955 (N_1955,N_1772,N_1773);
nand U1956 (N_1956,N_1704,N_1777);
and U1957 (N_1957,N_1725,N_1689);
nand U1958 (N_1958,N_1736,N_1615);
nand U1959 (N_1959,N_1646,N_1669);
nor U1960 (N_1960,N_1798,N_1623);
nor U1961 (N_1961,N_1638,N_1649);
and U1962 (N_1962,N_1707,N_1776);
or U1963 (N_1963,N_1622,N_1788);
nand U1964 (N_1964,N_1705,N_1723);
and U1965 (N_1965,N_1606,N_1652);
nor U1966 (N_1966,N_1624,N_1698);
nand U1967 (N_1967,N_1770,N_1637);
and U1968 (N_1968,N_1761,N_1629);
nor U1969 (N_1969,N_1770,N_1610);
nor U1970 (N_1970,N_1741,N_1676);
nor U1971 (N_1971,N_1710,N_1751);
nand U1972 (N_1972,N_1725,N_1608);
and U1973 (N_1973,N_1657,N_1627);
nor U1974 (N_1974,N_1614,N_1618);
or U1975 (N_1975,N_1666,N_1697);
or U1976 (N_1976,N_1764,N_1694);
or U1977 (N_1977,N_1760,N_1751);
and U1978 (N_1978,N_1797,N_1639);
or U1979 (N_1979,N_1708,N_1660);
nor U1980 (N_1980,N_1608,N_1758);
xor U1981 (N_1981,N_1711,N_1655);
nor U1982 (N_1982,N_1757,N_1610);
nor U1983 (N_1983,N_1793,N_1752);
and U1984 (N_1984,N_1607,N_1755);
nor U1985 (N_1985,N_1792,N_1679);
xnor U1986 (N_1986,N_1715,N_1671);
nor U1987 (N_1987,N_1786,N_1732);
nor U1988 (N_1988,N_1796,N_1640);
and U1989 (N_1989,N_1606,N_1799);
nand U1990 (N_1990,N_1736,N_1655);
or U1991 (N_1991,N_1761,N_1680);
and U1992 (N_1992,N_1726,N_1717);
and U1993 (N_1993,N_1721,N_1647);
and U1994 (N_1994,N_1650,N_1770);
nor U1995 (N_1995,N_1724,N_1739);
xor U1996 (N_1996,N_1720,N_1654);
and U1997 (N_1997,N_1739,N_1735);
and U1998 (N_1998,N_1740,N_1789);
nand U1999 (N_1999,N_1683,N_1650);
nor U2000 (N_2000,N_1900,N_1820);
and U2001 (N_2001,N_1842,N_1831);
and U2002 (N_2002,N_1975,N_1817);
or U2003 (N_2003,N_1938,N_1993);
xor U2004 (N_2004,N_1876,N_1874);
nand U2005 (N_2005,N_1880,N_1833);
nand U2006 (N_2006,N_1855,N_1877);
nand U2007 (N_2007,N_1854,N_1872);
nand U2008 (N_2008,N_1819,N_1963);
and U2009 (N_2009,N_1934,N_1861);
or U2010 (N_2010,N_1837,N_1944);
or U2011 (N_2011,N_1950,N_1864);
or U2012 (N_2012,N_1912,N_1826);
nand U2013 (N_2013,N_1888,N_1964);
xnor U2014 (N_2014,N_1839,N_1850);
nand U2015 (N_2015,N_1980,N_1935);
or U2016 (N_2016,N_1985,N_1942);
nor U2017 (N_2017,N_1945,N_1914);
and U2018 (N_2018,N_1885,N_1869);
nand U2019 (N_2019,N_1960,N_1970);
or U2020 (N_2020,N_1919,N_1859);
nand U2021 (N_2021,N_1862,N_1917);
and U2022 (N_2022,N_1816,N_1903);
nor U2023 (N_2023,N_1966,N_1858);
nor U2024 (N_2024,N_1807,N_1961);
nor U2025 (N_2025,N_1882,N_1927);
nand U2026 (N_2026,N_1863,N_1846);
or U2027 (N_2027,N_1968,N_1986);
nand U2028 (N_2028,N_1867,N_1892);
nand U2029 (N_2029,N_1937,N_1998);
or U2030 (N_2030,N_1875,N_1948);
and U2031 (N_2031,N_1881,N_1959);
or U2032 (N_2032,N_1838,N_1922);
nor U2033 (N_2033,N_1982,N_1893);
or U2034 (N_2034,N_1990,N_1887);
and U2035 (N_2035,N_1891,N_1840);
nor U2036 (N_2036,N_1916,N_1984);
xnor U2037 (N_2037,N_1886,N_1977);
and U2038 (N_2038,N_1847,N_1987);
or U2039 (N_2039,N_1971,N_1871);
nor U2040 (N_2040,N_1953,N_1878);
nand U2041 (N_2041,N_1805,N_1992);
nand U2042 (N_2042,N_1815,N_1883);
xor U2043 (N_2043,N_1907,N_1997);
and U2044 (N_2044,N_1921,N_1910);
nand U2045 (N_2045,N_1849,N_1909);
nor U2046 (N_2046,N_1821,N_1940);
nand U2047 (N_2047,N_1889,N_1979);
or U2048 (N_2048,N_1829,N_1870);
or U2049 (N_2049,N_1943,N_1905);
or U2050 (N_2050,N_1834,N_1879);
xnor U2051 (N_2051,N_1845,N_1811);
or U2052 (N_2052,N_1824,N_1902);
xor U2053 (N_2053,N_1852,N_1976);
nand U2054 (N_2054,N_1808,N_1956);
nand U2055 (N_2055,N_1936,N_1955);
nor U2056 (N_2056,N_1822,N_1809);
nor U2057 (N_2057,N_1929,N_1920);
nor U2058 (N_2058,N_1894,N_1967);
and U2059 (N_2059,N_1974,N_1931);
nor U2060 (N_2060,N_1973,N_1813);
nand U2061 (N_2061,N_1926,N_1962);
nor U2062 (N_2062,N_1951,N_1918);
nor U2063 (N_2063,N_1853,N_1895);
xnor U2064 (N_2064,N_1983,N_1954);
and U2065 (N_2065,N_1806,N_1901);
nand U2066 (N_2066,N_1965,N_1949);
or U2067 (N_2067,N_1915,N_1856);
nand U2068 (N_2068,N_1841,N_1930);
and U2069 (N_2069,N_1988,N_1827);
or U2070 (N_2070,N_1939,N_1941);
nor U2071 (N_2071,N_1828,N_1851);
nor U2072 (N_2072,N_1947,N_1946);
nand U2073 (N_2073,N_1814,N_1957);
nand U2074 (N_2074,N_1981,N_1835);
nor U2075 (N_2075,N_1924,N_1801);
xnor U2076 (N_2076,N_1890,N_1810);
and U2077 (N_2077,N_1844,N_1995);
nand U2078 (N_2078,N_1836,N_1843);
or U2079 (N_2079,N_1991,N_1978);
nor U2080 (N_2080,N_1899,N_1818);
nor U2081 (N_2081,N_1932,N_1952);
or U2082 (N_2082,N_1804,N_1911);
nand U2083 (N_2083,N_1823,N_1933);
nand U2084 (N_2084,N_1898,N_1868);
nand U2085 (N_2085,N_1896,N_1857);
and U2086 (N_2086,N_1803,N_1928);
nand U2087 (N_2087,N_1866,N_1908);
nand U2088 (N_2088,N_1906,N_1860);
and U2089 (N_2089,N_1865,N_1830);
nand U2090 (N_2090,N_1800,N_1848);
xor U2091 (N_2091,N_1897,N_1873);
nor U2092 (N_2092,N_1972,N_1802);
and U2093 (N_2093,N_1994,N_1996);
xnor U2094 (N_2094,N_1904,N_1989);
nor U2095 (N_2095,N_1832,N_1925);
or U2096 (N_2096,N_1958,N_1969);
nand U2097 (N_2097,N_1913,N_1884);
nand U2098 (N_2098,N_1812,N_1923);
nand U2099 (N_2099,N_1999,N_1825);
nand U2100 (N_2100,N_1851,N_1928);
nand U2101 (N_2101,N_1897,N_1885);
or U2102 (N_2102,N_1842,N_1998);
xor U2103 (N_2103,N_1857,N_1908);
or U2104 (N_2104,N_1941,N_1884);
nand U2105 (N_2105,N_1992,N_1810);
xnor U2106 (N_2106,N_1891,N_1928);
or U2107 (N_2107,N_1838,N_1987);
and U2108 (N_2108,N_1897,N_1868);
and U2109 (N_2109,N_1860,N_1876);
and U2110 (N_2110,N_1963,N_1840);
nor U2111 (N_2111,N_1947,N_1883);
nor U2112 (N_2112,N_1950,N_1973);
nand U2113 (N_2113,N_1960,N_1952);
nand U2114 (N_2114,N_1914,N_1919);
nand U2115 (N_2115,N_1984,N_1989);
and U2116 (N_2116,N_1882,N_1876);
nor U2117 (N_2117,N_1822,N_1980);
nor U2118 (N_2118,N_1931,N_1932);
or U2119 (N_2119,N_1995,N_1885);
and U2120 (N_2120,N_1975,N_1873);
or U2121 (N_2121,N_1863,N_1941);
or U2122 (N_2122,N_1801,N_1961);
and U2123 (N_2123,N_1983,N_1980);
xnor U2124 (N_2124,N_1917,N_1888);
nor U2125 (N_2125,N_1857,N_1997);
or U2126 (N_2126,N_1841,N_1880);
and U2127 (N_2127,N_1962,N_1945);
or U2128 (N_2128,N_1917,N_1949);
nand U2129 (N_2129,N_1957,N_1825);
xnor U2130 (N_2130,N_1980,N_1859);
nor U2131 (N_2131,N_1955,N_1875);
xor U2132 (N_2132,N_1981,N_1846);
nand U2133 (N_2133,N_1855,N_1833);
xor U2134 (N_2134,N_1901,N_1908);
nor U2135 (N_2135,N_1990,N_1803);
xor U2136 (N_2136,N_1965,N_1924);
nor U2137 (N_2137,N_1880,N_1849);
or U2138 (N_2138,N_1819,N_1990);
xnor U2139 (N_2139,N_1852,N_1828);
and U2140 (N_2140,N_1864,N_1922);
nand U2141 (N_2141,N_1856,N_1805);
nand U2142 (N_2142,N_1816,N_1827);
nor U2143 (N_2143,N_1858,N_1992);
and U2144 (N_2144,N_1840,N_1863);
nor U2145 (N_2145,N_1972,N_1803);
nand U2146 (N_2146,N_1891,N_1956);
nand U2147 (N_2147,N_1800,N_1963);
nor U2148 (N_2148,N_1951,N_1892);
and U2149 (N_2149,N_1989,N_1933);
xnor U2150 (N_2150,N_1958,N_1999);
nor U2151 (N_2151,N_1933,N_1843);
nor U2152 (N_2152,N_1813,N_1979);
and U2153 (N_2153,N_1855,N_1812);
nor U2154 (N_2154,N_1869,N_1983);
or U2155 (N_2155,N_1916,N_1966);
xnor U2156 (N_2156,N_1967,N_1908);
nor U2157 (N_2157,N_1916,N_1862);
nor U2158 (N_2158,N_1842,N_1887);
xor U2159 (N_2159,N_1840,N_1882);
or U2160 (N_2160,N_1821,N_1878);
or U2161 (N_2161,N_1870,N_1951);
nand U2162 (N_2162,N_1970,N_1974);
or U2163 (N_2163,N_1914,N_1880);
xnor U2164 (N_2164,N_1960,N_1879);
nor U2165 (N_2165,N_1983,N_1998);
and U2166 (N_2166,N_1968,N_1829);
nor U2167 (N_2167,N_1896,N_1956);
or U2168 (N_2168,N_1901,N_1894);
xnor U2169 (N_2169,N_1816,N_1818);
nand U2170 (N_2170,N_1926,N_1953);
nand U2171 (N_2171,N_1947,N_1842);
nand U2172 (N_2172,N_1825,N_1800);
and U2173 (N_2173,N_1866,N_1841);
or U2174 (N_2174,N_1870,N_1938);
or U2175 (N_2175,N_1897,N_1838);
or U2176 (N_2176,N_1909,N_1862);
and U2177 (N_2177,N_1898,N_1924);
or U2178 (N_2178,N_1999,N_1997);
and U2179 (N_2179,N_1905,N_1907);
and U2180 (N_2180,N_1950,N_1974);
or U2181 (N_2181,N_1980,N_1805);
or U2182 (N_2182,N_1863,N_1877);
nand U2183 (N_2183,N_1855,N_1982);
or U2184 (N_2184,N_1866,N_1845);
or U2185 (N_2185,N_1869,N_1947);
and U2186 (N_2186,N_1886,N_1857);
xor U2187 (N_2187,N_1862,N_1827);
nor U2188 (N_2188,N_1957,N_1980);
xnor U2189 (N_2189,N_1802,N_1821);
nor U2190 (N_2190,N_1985,N_1851);
or U2191 (N_2191,N_1876,N_1814);
nand U2192 (N_2192,N_1818,N_1823);
and U2193 (N_2193,N_1859,N_1884);
nor U2194 (N_2194,N_1937,N_1956);
and U2195 (N_2195,N_1980,N_1873);
nand U2196 (N_2196,N_1895,N_1970);
and U2197 (N_2197,N_1808,N_1827);
and U2198 (N_2198,N_1875,N_1978);
nand U2199 (N_2199,N_1810,N_1959);
nor U2200 (N_2200,N_2107,N_2067);
nand U2201 (N_2201,N_2196,N_2122);
nor U2202 (N_2202,N_2194,N_2025);
and U2203 (N_2203,N_2034,N_2002);
and U2204 (N_2204,N_2033,N_2080);
or U2205 (N_2205,N_2073,N_2129);
or U2206 (N_2206,N_2123,N_2050);
nor U2207 (N_2207,N_2181,N_2051);
nand U2208 (N_2208,N_2147,N_2057);
nor U2209 (N_2209,N_2044,N_2005);
nand U2210 (N_2210,N_2108,N_2008);
nor U2211 (N_2211,N_2141,N_2156);
xnor U2212 (N_2212,N_2182,N_2151);
and U2213 (N_2213,N_2039,N_2017);
or U2214 (N_2214,N_2176,N_2171);
nand U2215 (N_2215,N_2105,N_2028);
nor U2216 (N_2216,N_2072,N_2082);
and U2217 (N_2217,N_2098,N_2099);
and U2218 (N_2218,N_2116,N_2012);
nand U2219 (N_2219,N_2081,N_2078);
nand U2220 (N_2220,N_2024,N_2112);
nand U2221 (N_2221,N_2053,N_2007);
nor U2222 (N_2222,N_2027,N_2134);
nor U2223 (N_2223,N_2075,N_2135);
nor U2224 (N_2224,N_2140,N_2093);
nand U2225 (N_2225,N_2056,N_2113);
or U2226 (N_2226,N_2037,N_2029);
or U2227 (N_2227,N_2136,N_2199);
or U2228 (N_2228,N_2168,N_2074);
and U2229 (N_2229,N_2069,N_2126);
and U2230 (N_2230,N_2010,N_2085);
or U2231 (N_2231,N_2009,N_2094);
or U2232 (N_2232,N_2106,N_2132);
xnor U2233 (N_2233,N_2054,N_2131);
or U2234 (N_2234,N_2114,N_2117);
or U2235 (N_2235,N_2128,N_2097);
nor U2236 (N_2236,N_2011,N_2162);
or U2237 (N_2237,N_2018,N_2020);
and U2238 (N_2238,N_2137,N_2143);
and U2239 (N_2239,N_2150,N_2148);
nor U2240 (N_2240,N_2120,N_2102);
nor U2241 (N_2241,N_2086,N_2042);
and U2242 (N_2242,N_2088,N_2071);
nand U2243 (N_2243,N_2124,N_2026);
nand U2244 (N_2244,N_2019,N_2160);
and U2245 (N_2245,N_2153,N_2161);
or U2246 (N_2246,N_2096,N_2188);
and U2247 (N_2247,N_2164,N_2154);
or U2248 (N_2248,N_2159,N_2142);
xor U2249 (N_2249,N_2041,N_2193);
nand U2250 (N_2250,N_2004,N_2197);
or U2251 (N_2251,N_2163,N_2121);
or U2252 (N_2252,N_2092,N_2187);
nor U2253 (N_2253,N_2145,N_2065);
or U2254 (N_2254,N_2152,N_2127);
nand U2255 (N_2255,N_2047,N_2158);
nand U2256 (N_2256,N_2003,N_2023);
nor U2257 (N_2257,N_2125,N_2046);
nand U2258 (N_2258,N_2119,N_2035);
nor U2259 (N_2259,N_2058,N_2090);
or U2260 (N_2260,N_2149,N_2070);
nor U2261 (N_2261,N_2104,N_2014);
or U2262 (N_2262,N_2083,N_2022);
and U2263 (N_2263,N_2180,N_2006);
and U2264 (N_2264,N_2174,N_2061);
nor U2265 (N_2265,N_2016,N_2190);
nor U2266 (N_2266,N_2048,N_2144);
nor U2267 (N_2267,N_2178,N_2084);
nand U2268 (N_2268,N_2043,N_2169);
and U2269 (N_2269,N_2064,N_2192);
nand U2270 (N_2270,N_2191,N_2103);
nor U2271 (N_2271,N_2179,N_2100);
xnor U2272 (N_2272,N_2189,N_2165);
or U2273 (N_2273,N_2167,N_2089);
nor U2274 (N_2274,N_2166,N_2038);
and U2275 (N_2275,N_2045,N_2077);
and U2276 (N_2276,N_2172,N_2052);
or U2277 (N_2277,N_2138,N_2000);
nand U2278 (N_2278,N_2021,N_2133);
nor U2279 (N_2279,N_2109,N_2184);
and U2280 (N_2280,N_2040,N_2087);
nor U2281 (N_2281,N_2155,N_2062);
nor U2282 (N_2282,N_2115,N_2091);
or U2283 (N_2283,N_2063,N_2055);
xnor U2284 (N_2284,N_2195,N_2013);
and U2285 (N_2285,N_2076,N_2031);
nor U2286 (N_2286,N_2095,N_2139);
and U2287 (N_2287,N_2049,N_2157);
and U2288 (N_2288,N_2177,N_2066);
xnor U2289 (N_2289,N_2079,N_2059);
nor U2290 (N_2290,N_2068,N_2111);
nand U2291 (N_2291,N_2030,N_2198);
or U2292 (N_2292,N_2185,N_2175);
and U2293 (N_2293,N_2015,N_2001);
xnor U2294 (N_2294,N_2130,N_2173);
and U2295 (N_2295,N_2101,N_2060);
and U2296 (N_2296,N_2186,N_2118);
and U2297 (N_2297,N_2110,N_2036);
nor U2298 (N_2298,N_2170,N_2183);
and U2299 (N_2299,N_2032,N_2146);
nor U2300 (N_2300,N_2018,N_2179);
or U2301 (N_2301,N_2110,N_2007);
and U2302 (N_2302,N_2184,N_2003);
nor U2303 (N_2303,N_2128,N_2162);
nand U2304 (N_2304,N_2088,N_2110);
and U2305 (N_2305,N_2039,N_2031);
or U2306 (N_2306,N_2060,N_2108);
or U2307 (N_2307,N_2081,N_2047);
xnor U2308 (N_2308,N_2037,N_2134);
nor U2309 (N_2309,N_2178,N_2102);
nor U2310 (N_2310,N_2152,N_2095);
nand U2311 (N_2311,N_2001,N_2153);
or U2312 (N_2312,N_2191,N_2119);
or U2313 (N_2313,N_2080,N_2057);
nor U2314 (N_2314,N_2083,N_2045);
nor U2315 (N_2315,N_2149,N_2044);
nor U2316 (N_2316,N_2117,N_2196);
nor U2317 (N_2317,N_2119,N_2196);
nor U2318 (N_2318,N_2006,N_2164);
and U2319 (N_2319,N_2097,N_2174);
nand U2320 (N_2320,N_2155,N_2017);
xor U2321 (N_2321,N_2041,N_2126);
and U2322 (N_2322,N_2172,N_2089);
and U2323 (N_2323,N_2191,N_2027);
xnor U2324 (N_2324,N_2182,N_2143);
or U2325 (N_2325,N_2020,N_2015);
nand U2326 (N_2326,N_2122,N_2098);
xnor U2327 (N_2327,N_2055,N_2053);
nor U2328 (N_2328,N_2009,N_2190);
nor U2329 (N_2329,N_2184,N_2122);
and U2330 (N_2330,N_2078,N_2013);
and U2331 (N_2331,N_2128,N_2192);
nor U2332 (N_2332,N_2150,N_2196);
nor U2333 (N_2333,N_2187,N_2120);
nor U2334 (N_2334,N_2112,N_2185);
nand U2335 (N_2335,N_2063,N_2141);
or U2336 (N_2336,N_2044,N_2113);
nand U2337 (N_2337,N_2065,N_2029);
or U2338 (N_2338,N_2172,N_2141);
and U2339 (N_2339,N_2020,N_2014);
nor U2340 (N_2340,N_2093,N_2159);
or U2341 (N_2341,N_2108,N_2119);
and U2342 (N_2342,N_2149,N_2045);
and U2343 (N_2343,N_2160,N_2193);
and U2344 (N_2344,N_2095,N_2049);
xor U2345 (N_2345,N_2148,N_2087);
nand U2346 (N_2346,N_2181,N_2072);
or U2347 (N_2347,N_2171,N_2101);
nand U2348 (N_2348,N_2109,N_2163);
or U2349 (N_2349,N_2145,N_2059);
nor U2350 (N_2350,N_2000,N_2011);
nor U2351 (N_2351,N_2052,N_2027);
and U2352 (N_2352,N_2107,N_2019);
nor U2353 (N_2353,N_2121,N_2172);
or U2354 (N_2354,N_2178,N_2165);
and U2355 (N_2355,N_2150,N_2018);
nand U2356 (N_2356,N_2150,N_2068);
nand U2357 (N_2357,N_2053,N_2012);
nor U2358 (N_2358,N_2123,N_2098);
nand U2359 (N_2359,N_2114,N_2144);
and U2360 (N_2360,N_2138,N_2159);
or U2361 (N_2361,N_2166,N_2013);
nand U2362 (N_2362,N_2094,N_2128);
or U2363 (N_2363,N_2008,N_2117);
nand U2364 (N_2364,N_2075,N_2148);
nor U2365 (N_2365,N_2087,N_2083);
or U2366 (N_2366,N_2184,N_2031);
nand U2367 (N_2367,N_2110,N_2144);
nand U2368 (N_2368,N_2149,N_2141);
or U2369 (N_2369,N_2093,N_2158);
nor U2370 (N_2370,N_2198,N_2142);
and U2371 (N_2371,N_2020,N_2101);
nor U2372 (N_2372,N_2044,N_2110);
or U2373 (N_2373,N_2126,N_2110);
and U2374 (N_2374,N_2176,N_2004);
nor U2375 (N_2375,N_2179,N_2050);
nand U2376 (N_2376,N_2133,N_2192);
and U2377 (N_2377,N_2001,N_2119);
xnor U2378 (N_2378,N_2110,N_2104);
nand U2379 (N_2379,N_2131,N_2010);
or U2380 (N_2380,N_2017,N_2173);
or U2381 (N_2381,N_2180,N_2173);
nor U2382 (N_2382,N_2085,N_2178);
nor U2383 (N_2383,N_2133,N_2061);
nand U2384 (N_2384,N_2055,N_2015);
nand U2385 (N_2385,N_2062,N_2125);
nor U2386 (N_2386,N_2032,N_2013);
nand U2387 (N_2387,N_2130,N_2127);
and U2388 (N_2388,N_2107,N_2086);
and U2389 (N_2389,N_2169,N_2180);
and U2390 (N_2390,N_2108,N_2031);
nor U2391 (N_2391,N_2134,N_2091);
nor U2392 (N_2392,N_2162,N_2120);
or U2393 (N_2393,N_2077,N_2140);
or U2394 (N_2394,N_2159,N_2104);
or U2395 (N_2395,N_2089,N_2028);
nand U2396 (N_2396,N_2162,N_2199);
nor U2397 (N_2397,N_2112,N_2039);
nor U2398 (N_2398,N_2010,N_2195);
and U2399 (N_2399,N_2025,N_2126);
or U2400 (N_2400,N_2287,N_2309);
or U2401 (N_2401,N_2235,N_2241);
nand U2402 (N_2402,N_2387,N_2252);
xnor U2403 (N_2403,N_2391,N_2229);
nand U2404 (N_2404,N_2389,N_2340);
or U2405 (N_2405,N_2376,N_2293);
and U2406 (N_2406,N_2201,N_2210);
nor U2407 (N_2407,N_2351,N_2356);
nor U2408 (N_2408,N_2276,N_2240);
nor U2409 (N_2409,N_2226,N_2335);
nand U2410 (N_2410,N_2336,N_2251);
and U2411 (N_2411,N_2237,N_2326);
and U2412 (N_2412,N_2219,N_2374);
and U2413 (N_2413,N_2362,N_2332);
nor U2414 (N_2414,N_2382,N_2386);
and U2415 (N_2415,N_2259,N_2242);
nand U2416 (N_2416,N_2277,N_2288);
and U2417 (N_2417,N_2290,N_2263);
nor U2418 (N_2418,N_2346,N_2325);
and U2419 (N_2419,N_2261,N_2212);
and U2420 (N_2420,N_2239,N_2268);
nand U2421 (N_2421,N_2398,N_2305);
or U2422 (N_2422,N_2352,N_2255);
nor U2423 (N_2423,N_2397,N_2365);
xor U2424 (N_2424,N_2223,N_2321);
nor U2425 (N_2425,N_2303,N_2214);
xor U2426 (N_2426,N_2316,N_2218);
xor U2427 (N_2427,N_2289,N_2300);
and U2428 (N_2428,N_2361,N_2301);
nor U2429 (N_2429,N_2298,N_2227);
nor U2430 (N_2430,N_2260,N_2215);
and U2431 (N_2431,N_2370,N_2209);
nor U2432 (N_2432,N_2393,N_2249);
and U2433 (N_2433,N_2334,N_2314);
and U2434 (N_2434,N_2394,N_2299);
nor U2435 (N_2435,N_2354,N_2367);
nand U2436 (N_2436,N_2312,N_2269);
xor U2437 (N_2437,N_2317,N_2294);
nand U2438 (N_2438,N_2205,N_2375);
nand U2439 (N_2439,N_2328,N_2228);
or U2440 (N_2440,N_2270,N_2272);
and U2441 (N_2441,N_2213,N_2322);
and U2442 (N_2442,N_2379,N_2265);
or U2443 (N_2443,N_2246,N_2230);
and U2444 (N_2444,N_2368,N_2324);
nor U2445 (N_2445,N_2355,N_2337);
nand U2446 (N_2446,N_2345,N_2318);
nand U2447 (N_2447,N_2378,N_2264);
and U2448 (N_2448,N_2392,N_2281);
and U2449 (N_2449,N_2286,N_2206);
nor U2450 (N_2450,N_2248,N_2307);
and U2451 (N_2451,N_2285,N_2359);
or U2452 (N_2452,N_2258,N_2310);
or U2453 (N_2453,N_2384,N_2211);
or U2454 (N_2454,N_2304,N_2256);
and U2455 (N_2455,N_2247,N_2347);
nand U2456 (N_2456,N_2262,N_2279);
or U2457 (N_2457,N_2253,N_2331);
or U2458 (N_2458,N_2296,N_2373);
or U2459 (N_2459,N_2369,N_2364);
or U2460 (N_2460,N_2372,N_2250);
or U2461 (N_2461,N_2280,N_2327);
nand U2462 (N_2462,N_2366,N_2399);
or U2463 (N_2463,N_2202,N_2254);
and U2464 (N_2464,N_2319,N_2315);
or U2465 (N_2465,N_2274,N_2353);
xnor U2466 (N_2466,N_2360,N_2395);
and U2467 (N_2467,N_2313,N_2232);
and U2468 (N_2468,N_2377,N_2349);
nor U2469 (N_2469,N_2200,N_2302);
or U2470 (N_2470,N_2284,N_2390);
and U2471 (N_2471,N_2363,N_2297);
nor U2472 (N_2472,N_2341,N_2231);
nor U2473 (N_2473,N_2343,N_2245);
or U2474 (N_2474,N_2308,N_2385);
nor U2475 (N_2475,N_2339,N_2207);
nand U2476 (N_2476,N_2233,N_2323);
xor U2477 (N_2477,N_2380,N_2338);
nand U2478 (N_2478,N_2273,N_2311);
nand U2479 (N_2479,N_2381,N_2291);
and U2480 (N_2480,N_2266,N_2220);
or U2481 (N_2481,N_2221,N_2383);
nor U2482 (N_2482,N_2282,N_2204);
or U2483 (N_2483,N_2234,N_2224);
or U2484 (N_2484,N_2243,N_2357);
nor U2485 (N_2485,N_2271,N_2217);
nand U2486 (N_2486,N_2342,N_2216);
and U2487 (N_2487,N_2236,N_2358);
nand U2488 (N_2488,N_2267,N_2329);
or U2489 (N_2489,N_2275,N_2344);
and U2490 (N_2490,N_2306,N_2208);
or U2491 (N_2491,N_2350,N_2283);
xor U2492 (N_2492,N_2244,N_2225);
nor U2493 (N_2493,N_2371,N_2348);
or U2494 (N_2494,N_2257,N_2333);
and U2495 (N_2495,N_2320,N_2396);
or U2496 (N_2496,N_2203,N_2388);
and U2497 (N_2497,N_2278,N_2222);
and U2498 (N_2498,N_2292,N_2330);
or U2499 (N_2499,N_2238,N_2295);
or U2500 (N_2500,N_2201,N_2313);
and U2501 (N_2501,N_2258,N_2349);
nand U2502 (N_2502,N_2251,N_2280);
nand U2503 (N_2503,N_2377,N_2212);
xor U2504 (N_2504,N_2231,N_2272);
nor U2505 (N_2505,N_2219,N_2247);
nor U2506 (N_2506,N_2320,N_2253);
nand U2507 (N_2507,N_2252,N_2263);
or U2508 (N_2508,N_2328,N_2311);
xnor U2509 (N_2509,N_2335,N_2310);
and U2510 (N_2510,N_2302,N_2369);
nand U2511 (N_2511,N_2280,N_2390);
nand U2512 (N_2512,N_2248,N_2296);
or U2513 (N_2513,N_2212,N_2336);
nand U2514 (N_2514,N_2219,N_2390);
xor U2515 (N_2515,N_2238,N_2203);
or U2516 (N_2516,N_2231,N_2375);
and U2517 (N_2517,N_2327,N_2210);
and U2518 (N_2518,N_2351,N_2313);
and U2519 (N_2519,N_2287,N_2370);
xnor U2520 (N_2520,N_2398,N_2306);
nor U2521 (N_2521,N_2229,N_2209);
and U2522 (N_2522,N_2333,N_2378);
nor U2523 (N_2523,N_2347,N_2216);
or U2524 (N_2524,N_2374,N_2276);
nor U2525 (N_2525,N_2215,N_2267);
nand U2526 (N_2526,N_2358,N_2204);
and U2527 (N_2527,N_2306,N_2299);
xnor U2528 (N_2528,N_2239,N_2392);
nor U2529 (N_2529,N_2346,N_2315);
or U2530 (N_2530,N_2389,N_2314);
and U2531 (N_2531,N_2340,N_2361);
and U2532 (N_2532,N_2382,N_2388);
xor U2533 (N_2533,N_2277,N_2389);
nand U2534 (N_2534,N_2310,N_2288);
or U2535 (N_2535,N_2389,N_2310);
or U2536 (N_2536,N_2312,N_2277);
and U2537 (N_2537,N_2397,N_2233);
or U2538 (N_2538,N_2202,N_2207);
nor U2539 (N_2539,N_2300,N_2332);
or U2540 (N_2540,N_2287,N_2304);
or U2541 (N_2541,N_2281,N_2322);
and U2542 (N_2542,N_2246,N_2336);
nand U2543 (N_2543,N_2265,N_2250);
or U2544 (N_2544,N_2296,N_2317);
or U2545 (N_2545,N_2217,N_2314);
xor U2546 (N_2546,N_2334,N_2218);
xnor U2547 (N_2547,N_2248,N_2316);
nand U2548 (N_2548,N_2242,N_2212);
nand U2549 (N_2549,N_2273,N_2262);
or U2550 (N_2550,N_2347,N_2329);
nor U2551 (N_2551,N_2308,N_2357);
nor U2552 (N_2552,N_2323,N_2204);
nor U2553 (N_2553,N_2220,N_2201);
and U2554 (N_2554,N_2316,N_2241);
nand U2555 (N_2555,N_2329,N_2354);
nor U2556 (N_2556,N_2310,N_2350);
nand U2557 (N_2557,N_2315,N_2366);
nor U2558 (N_2558,N_2330,N_2376);
xor U2559 (N_2559,N_2369,N_2360);
xor U2560 (N_2560,N_2210,N_2288);
nand U2561 (N_2561,N_2223,N_2366);
nor U2562 (N_2562,N_2305,N_2245);
nor U2563 (N_2563,N_2348,N_2293);
and U2564 (N_2564,N_2375,N_2303);
nor U2565 (N_2565,N_2291,N_2326);
and U2566 (N_2566,N_2221,N_2253);
or U2567 (N_2567,N_2219,N_2379);
nor U2568 (N_2568,N_2210,N_2357);
xnor U2569 (N_2569,N_2226,N_2263);
xor U2570 (N_2570,N_2397,N_2232);
xnor U2571 (N_2571,N_2275,N_2221);
or U2572 (N_2572,N_2286,N_2264);
and U2573 (N_2573,N_2231,N_2216);
or U2574 (N_2574,N_2291,N_2270);
xor U2575 (N_2575,N_2272,N_2313);
nor U2576 (N_2576,N_2298,N_2343);
or U2577 (N_2577,N_2239,N_2312);
or U2578 (N_2578,N_2229,N_2363);
nor U2579 (N_2579,N_2389,N_2239);
nand U2580 (N_2580,N_2303,N_2344);
and U2581 (N_2581,N_2368,N_2349);
nand U2582 (N_2582,N_2278,N_2302);
nor U2583 (N_2583,N_2388,N_2266);
nand U2584 (N_2584,N_2272,N_2200);
or U2585 (N_2585,N_2218,N_2203);
nor U2586 (N_2586,N_2231,N_2327);
nor U2587 (N_2587,N_2202,N_2201);
or U2588 (N_2588,N_2278,N_2290);
nand U2589 (N_2589,N_2222,N_2370);
nand U2590 (N_2590,N_2370,N_2203);
nor U2591 (N_2591,N_2248,N_2253);
or U2592 (N_2592,N_2355,N_2331);
and U2593 (N_2593,N_2339,N_2204);
and U2594 (N_2594,N_2335,N_2265);
xor U2595 (N_2595,N_2237,N_2270);
and U2596 (N_2596,N_2362,N_2231);
and U2597 (N_2597,N_2269,N_2366);
nor U2598 (N_2598,N_2288,N_2256);
and U2599 (N_2599,N_2396,N_2292);
nor U2600 (N_2600,N_2518,N_2581);
nand U2601 (N_2601,N_2499,N_2587);
and U2602 (N_2602,N_2456,N_2495);
or U2603 (N_2603,N_2452,N_2457);
nor U2604 (N_2604,N_2554,N_2486);
xnor U2605 (N_2605,N_2543,N_2591);
xor U2606 (N_2606,N_2563,N_2586);
or U2607 (N_2607,N_2509,N_2411);
nand U2608 (N_2608,N_2467,N_2445);
nor U2609 (N_2609,N_2590,N_2559);
and U2610 (N_2610,N_2402,N_2502);
nor U2611 (N_2611,N_2498,N_2464);
xor U2612 (N_2612,N_2484,N_2419);
nor U2613 (N_2613,N_2597,N_2531);
nor U2614 (N_2614,N_2507,N_2596);
or U2615 (N_2615,N_2482,N_2497);
nor U2616 (N_2616,N_2517,N_2583);
nand U2617 (N_2617,N_2501,N_2442);
and U2618 (N_2618,N_2567,N_2435);
nand U2619 (N_2619,N_2440,N_2454);
or U2620 (N_2620,N_2471,N_2431);
nand U2621 (N_2621,N_2585,N_2429);
or U2622 (N_2622,N_2468,N_2438);
or U2623 (N_2623,N_2463,N_2422);
nor U2624 (N_2624,N_2552,N_2423);
xor U2625 (N_2625,N_2539,N_2489);
or U2626 (N_2626,N_2416,N_2459);
or U2627 (N_2627,N_2520,N_2549);
or U2628 (N_2628,N_2446,N_2528);
xor U2629 (N_2629,N_2481,N_2546);
nor U2630 (N_2630,N_2493,N_2455);
nand U2631 (N_2631,N_2475,N_2580);
and U2632 (N_2632,N_2503,N_2526);
and U2633 (N_2633,N_2473,N_2415);
nor U2634 (N_2634,N_2511,N_2557);
nor U2635 (N_2635,N_2523,N_2485);
and U2636 (N_2636,N_2564,N_2448);
or U2637 (N_2637,N_2444,N_2451);
or U2638 (N_2638,N_2414,N_2521);
or U2639 (N_2639,N_2584,N_2479);
and U2640 (N_2640,N_2558,N_2515);
nor U2641 (N_2641,N_2408,N_2418);
nor U2642 (N_2642,N_2568,N_2400);
or U2643 (N_2643,N_2469,N_2465);
nor U2644 (N_2644,N_2578,N_2529);
and U2645 (N_2645,N_2466,N_2548);
xor U2646 (N_2646,N_2434,N_2426);
nand U2647 (N_2647,N_2439,N_2404);
nor U2648 (N_2648,N_2537,N_2405);
or U2649 (N_2649,N_2565,N_2472);
and U2650 (N_2650,N_2538,N_2589);
nor U2651 (N_2651,N_2576,N_2532);
and U2652 (N_2652,N_2421,N_2535);
nand U2653 (N_2653,N_2478,N_2570);
nand U2654 (N_2654,N_2410,N_2460);
xnor U2655 (N_2655,N_2401,N_2477);
and U2656 (N_2656,N_2447,N_2595);
nor U2657 (N_2657,N_2417,N_2571);
nor U2658 (N_2658,N_2533,N_2593);
nand U2659 (N_2659,N_2491,N_2594);
nand U2660 (N_2660,N_2504,N_2437);
and U2661 (N_2661,N_2407,N_2492);
or U2662 (N_2662,N_2449,N_2433);
nand U2663 (N_2663,N_2427,N_2406);
nand U2664 (N_2664,N_2579,N_2506);
nand U2665 (N_2665,N_2510,N_2540);
and U2666 (N_2666,N_2514,N_2458);
and U2667 (N_2667,N_2409,N_2547);
nor U2668 (N_2668,N_2566,N_2490);
or U2669 (N_2669,N_2474,N_2575);
nand U2670 (N_2670,N_2572,N_2592);
nor U2671 (N_2671,N_2441,N_2462);
and U2672 (N_2672,N_2476,N_2577);
nand U2673 (N_2673,N_2544,N_2500);
nor U2674 (N_2674,N_2403,N_2519);
nor U2675 (N_2675,N_2599,N_2480);
and U2676 (N_2676,N_2420,N_2527);
nand U2677 (N_2677,N_2551,N_2534);
nor U2678 (N_2678,N_2582,N_2562);
or U2679 (N_2679,N_2508,N_2496);
and U2680 (N_2680,N_2487,N_2424);
nor U2681 (N_2681,N_2494,N_2453);
nor U2682 (N_2682,N_2425,N_2461);
or U2683 (N_2683,N_2412,N_2450);
nand U2684 (N_2684,N_2560,N_2574);
or U2685 (N_2685,N_2536,N_2569);
or U2686 (N_2686,N_2555,N_2522);
nand U2687 (N_2687,N_2436,N_2443);
or U2688 (N_2688,N_2470,N_2525);
nand U2689 (N_2689,N_2430,N_2573);
nand U2690 (N_2690,N_2413,N_2432);
or U2691 (N_2691,N_2561,N_2516);
or U2692 (N_2692,N_2598,N_2530);
and U2693 (N_2693,N_2556,N_2483);
and U2694 (N_2694,N_2550,N_2553);
nand U2695 (N_2695,N_2488,N_2505);
or U2696 (N_2696,N_2545,N_2542);
and U2697 (N_2697,N_2512,N_2541);
and U2698 (N_2698,N_2513,N_2588);
or U2699 (N_2699,N_2524,N_2428);
and U2700 (N_2700,N_2426,N_2524);
or U2701 (N_2701,N_2475,N_2504);
or U2702 (N_2702,N_2579,N_2499);
and U2703 (N_2703,N_2567,N_2533);
xor U2704 (N_2704,N_2578,N_2542);
nor U2705 (N_2705,N_2489,N_2508);
and U2706 (N_2706,N_2413,N_2497);
or U2707 (N_2707,N_2592,N_2576);
or U2708 (N_2708,N_2552,N_2527);
nand U2709 (N_2709,N_2520,N_2472);
or U2710 (N_2710,N_2434,N_2520);
or U2711 (N_2711,N_2564,N_2538);
or U2712 (N_2712,N_2528,N_2439);
nor U2713 (N_2713,N_2561,N_2409);
nor U2714 (N_2714,N_2575,N_2426);
and U2715 (N_2715,N_2568,N_2540);
xor U2716 (N_2716,N_2453,N_2571);
nand U2717 (N_2717,N_2565,N_2499);
and U2718 (N_2718,N_2471,N_2588);
and U2719 (N_2719,N_2557,N_2419);
nand U2720 (N_2720,N_2474,N_2444);
nor U2721 (N_2721,N_2564,N_2455);
and U2722 (N_2722,N_2561,N_2477);
and U2723 (N_2723,N_2568,N_2589);
nor U2724 (N_2724,N_2502,N_2407);
nor U2725 (N_2725,N_2413,N_2534);
or U2726 (N_2726,N_2539,N_2460);
nand U2727 (N_2727,N_2431,N_2451);
xnor U2728 (N_2728,N_2479,N_2432);
nand U2729 (N_2729,N_2483,N_2487);
nand U2730 (N_2730,N_2551,N_2547);
and U2731 (N_2731,N_2482,N_2529);
nand U2732 (N_2732,N_2475,N_2450);
nor U2733 (N_2733,N_2412,N_2587);
nor U2734 (N_2734,N_2502,N_2463);
nand U2735 (N_2735,N_2553,N_2531);
nor U2736 (N_2736,N_2485,N_2513);
nand U2737 (N_2737,N_2576,N_2521);
or U2738 (N_2738,N_2540,N_2532);
nand U2739 (N_2739,N_2488,N_2551);
and U2740 (N_2740,N_2451,N_2588);
or U2741 (N_2741,N_2507,N_2524);
and U2742 (N_2742,N_2456,N_2422);
nor U2743 (N_2743,N_2424,N_2557);
xnor U2744 (N_2744,N_2487,N_2566);
nor U2745 (N_2745,N_2541,N_2438);
and U2746 (N_2746,N_2435,N_2463);
nand U2747 (N_2747,N_2548,N_2585);
and U2748 (N_2748,N_2547,N_2425);
and U2749 (N_2749,N_2455,N_2574);
or U2750 (N_2750,N_2579,N_2420);
xor U2751 (N_2751,N_2448,N_2435);
xor U2752 (N_2752,N_2439,N_2498);
nor U2753 (N_2753,N_2406,N_2589);
nor U2754 (N_2754,N_2435,N_2562);
nand U2755 (N_2755,N_2598,N_2403);
or U2756 (N_2756,N_2486,N_2480);
nand U2757 (N_2757,N_2430,N_2563);
nand U2758 (N_2758,N_2512,N_2582);
nor U2759 (N_2759,N_2438,N_2551);
xnor U2760 (N_2760,N_2590,N_2546);
or U2761 (N_2761,N_2576,N_2445);
nand U2762 (N_2762,N_2526,N_2551);
and U2763 (N_2763,N_2461,N_2530);
nor U2764 (N_2764,N_2538,N_2497);
xnor U2765 (N_2765,N_2482,N_2455);
or U2766 (N_2766,N_2547,N_2579);
and U2767 (N_2767,N_2409,N_2420);
or U2768 (N_2768,N_2480,N_2526);
or U2769 (N_2769,N_2572,N_2549);
nor U2770 (N_2770,N_2536,N_2551);
xor U2771 (N_2771,N_2466,N_2583);
or U2772 (N_2772,N_2423,N_2474);
or U2773 (N_2773,N_2479,N_2448);
and U2774 (N_2774,N_2473,N_2421);
nor U2775 (N_2775,N_2515,N_2539);
nand U2776 (N_2776,N_2452,N_2513);
and U2777 (N_2777,N_2590,N_2501);
xor U2778 (N_2778,N_2521,N_2439);
or U2779 (N_2779,N_2474,N_2449);
and U2780 (N_2780,N_2414,N_2427);
and U2781 (N_2781,N_2531,N_2451);
nand U2782 (N_2782,N_2574,N_2457);
nand U2783 (N_2783,N_2538,N_2587);
xor U2784 (N_2784,N_2430,N_2488);
nor U2785 (N_2785,N_2459,N_2478);
nand U2786 (N_2786,N_2428,N_2528);
nor U2787 (N_2787,N_2456,N_2563);
and U2788 (N_2788,N_2598,N_2441);
nand U2789 (N_2789,N_2570,N_2400);
nor U2790 (N_2790,N_2431,N_2403);
or U2791 (N_2791,N_2520,N_2552);
nand U2792 (N_2792,N_2488,N_2447);
nor U2793 (N_2793,N_2426,N_2560);
nor U2794 (N_2794,N_2577,N_2508);
and U2795 (N_2795,N_2478,N_2522);
nand U2796 (N_2796,N_2538,N_2487);
or U2797 (N_2797,N_2424,N_2515);
nor U2798 (N_2798,N_2469,N_2530);
and U2799 (N_2799,N_2443,N_2476);
or U2800 (N_2800,N_2741,N_2646);
xnor U2801 (N_2801,N_2652,N_2727);
or U2802 (N_2802,N_2726,N_2684);
nor U2803 (N_2803,N_2740,N_2743);
nand U2804 (N_2804,N_2709,N_2619);
xor U2805 (N_2805,N_2655,N_2681);
nand U2806 (N_2806,N_2617,N_2706);
and U2807 (N_2807,N_2779,N_2679);
nor U2808 (N_2808,N_2725,N_2644);
and U2809 (N_2809,N_2624,N_2680);
nor U2810 (N_2810,N_2641,N_2775);
and U2811 (N_2811,N_2688,N_2798);
or U2812 (N_2812,N_2794,N_2653);
nor U2813 (N_2813,N_2772,N_2643);
nand U2814 (N_2814,N_2745,N_2777);
and U2815 (N_2815,N_2654,N_2728);
and U2816 (N_2816,N_2712,N_2778);
and U2817 (N_2817,N_2666,N_2734);
and U2818 (N_2818,N_2671,N_2698);
nand U2819 (N_2819,N_2786,N_2760);
or U2820 (N_2820,N_2754,N_2766);
and U2821 (N_2821,N_2708,N_2776);
nor U2822 (N_2822,N_2642,N_2763);
and U2823 (N_2823,N_2699,N_2748);
nand U2824 (N_2824,N_2773,N_2636);
or U2825 (N_2825,N_2761,N_2612);
nand U2826 (N_2826,N_2675,N_2720);
nor U2827 (N_2827,N_2735,N_2659);
nor U2828 (N_2828,N_2780,N_2660);
xnor U2829 (N_2829,N_2759,N_2625);
nand U2830 (N_2830,N_2755,N_2685);
nand U2831 (N_2831,N_2647,N_2781);
nor U2832 (N_2832,N_2724,N_2694);
nor U2833 (N_2833,N_2610,N_2715);
or U2834 (N_2834,N_2795,N_2791);
or U2835 (N_2835,N_2613,N_2656);
or U2836 (N_2836,N_2606,N_2731);
nand U2837 (N_2837,N_2645,N_2723);
or U2838 (N_2838,N_2651,N_2722);
and U2839 (N_2839,N_2672,N_2600);
nor U2840 (N_2840,N_2609,N_2769);
nor U2841 (N_2841,N_2792,N_2718);
nand U2842 (N_2842,N_2733,N_2785);
and U2843 (N_2843,N_2782,N_2607);
nand U2844 (N_2844,N_2605,N_2742);
and U2845 (N_2845,N_2788,N_2611);
nand U2846 (N_2846,N_2604,N_2602);
nand U2847 (N_2847,N_2623,N_2616);
nand U2848 (N_2848,N_2774,N_2627);
and U2849 (N_2849,N_2736,N_2753);
and U2850 (N_2850,N_2670,N_2686);
or U2851 (N_2851,N_2667,N_2690);
xnor U2852 (N_2852,N_2710,N_2658);
nor U2853 (N_2853,N_2799,N_2716);
nor U2854 (N_2854,N_2637,N_2783);
xnor U2855 (N_2855,N_2707,N_2657);
xnor U2856 (N_2856,N_2676,N_2770);
nor U2857 (N_2857,N_2749,N_2750);
or U2858 (N_2858,N_2633,N_2704);
nor U2859 (N_2859,N_2664,N_2649);
or U2860 (N_2860,N_2677,N_2752);
xnor U2861 (N_2861,N_2638,N_2608);
nand U2862 (N_2862,N_2719,N_2758);
or U2863 (N_2863,N_2635,N_2618);
or U2864 (N_2864,N_2762,N_2797);
or U2865 (N_2865,N_2738,N_2687);
nor U2866 (N_2866,N_2757,N_2692);
or U2867 (N_2867,N_2665,N_2668);
nor U2868 (N_2868,N_2737,N_2730);
nor U2869 (N_2869,N_2793,N_2683);
and U2870 (N_2870,N_2601,N_2650);
or U2871 (N_2871,N_2703,N_2639);
and U2872 (N_2872,N_2771,N_2603);
or U2873 (N_2873,N_2717,N_2767);
or U2874 (N_2874,N_2705,N_2663);
nor U2875 (N_2875,N_2622,N_2751);
nand U2876 (N_2876,N_2695,N_2693);
or U2877 (N_2877,N_2732,N_2701);
or U2878 (N_2878,N_2661,N_2739);
xnor U2879 (N_2879,N_2669,N_2630);
or U2880 (N_2880,N_2765,N_2689);
and U2881 (N_2881,N_2634,N_2629);
and U2882 (N_2882,N_2784,N_2620);
nand U2883 (N_2883,N_2768,N_2747);
xnor U2884 (N_2884,N_2632,N_2721);
nor U2885 (N_2885,N_2682,N_2764);
nor U2886 (N_2886,N_2614,N_2696);
or U2887 (N_2887,N_2640,N_2648);
or U2888 (N_2888,N_2787,N_2673);
and U2889 (N_2889,N_2744,N_2621);
nand U2890 (N_2890,N_2628,N_2702);
and U2891 (N_2891,N_2729,N_2631);
nand U2892 (N_2892,N_2711,N_2756);
nor U2893 (N_2893,N_2789,N_2678);
xor U2894 (N_2894,N_2662,N_2697);
nand U2895 (N_2895,N_2790,N_2796);
nand U2896 (N_2896,N_2700,N_2615);
nor U2897 (N_2897,N_2626,N_2746);
and U2898 (N_2898,N_2713,N_2691);
nor U2899 (N_2899,N_2674,N_2714);
and U2900 (N_2900,N_2771,N_2722);
and U2901 (N_2901,N_2779,N_2796);
nand U2902 (N_2902,N_2741,N_2715);
or U2903 (N_2903,N_2651,N_2780);
xor U2904 (N_2904,N_2710,N_2669);
and U2905 (N_2905,N_2609,N_2755);
nor U2906 (N_2906,N_2757,N_2683);
and U2907 (N_2907,N_2737,N_2673);
and U2908 (N_2908,N_2732,N_2707);
nand U2909 (N_2909,N_2797,N_2728);
nor U2910 (N_2910,N_2739,N_2740);
nand U2911 (N_2911,N_2760,N_2660);
nor U2912 (N_2912,N_2665,N_2736);
nand U2913 (N_2913,N_2724,N_2772);
and U2914 (N_2914,N_2662,N_2652);
or U2915 (N_2915,N_2777,N_2740);
or U2916 (N_2916,N_2631,N_2669);
or U2917 (N_2917,N_2657,N_2608);
nand U2918 (N_2918,N_2670,N_2629);
or U2919 (N_2919,N_2759,N_2630);
and U2920 (N_2920,N_2616,N_2645);
nand U2921 (N_2921,N_2755,N_2670);
or U2922 (N_2922,N_2634,N_2690);
nor U2923 (N_2923,N_2771,N_2745);
nand U2924 (N_2924,N_2655,N_2708);
nor U2925 (N_2925,N_2760,N_2763);
nand U2926 (N_2926,N_2796,N_2653);
and U2927 (N_2927,N_2724,N_2726);
nor U2928 (N_2928,N_2782,N_2792);
and U2929 (N_2929,N_2605,N_2645);
xor U2930 (N_2930,N_2734,N_2764);
nand U2931 (N_2931,N_2669,N_2723);
or U2932 (N_2932,N_2677,N_2762);
and U2933 (N_2933,N_2600,N_2616);
nor U2934 (N_2934,N_2709,N_2681);
or U2935 (N_2935,N_2704,N_2611);
nor U2936 (N_2936,N_2781,N_2635);
nand U2937 (N_2937,N_2682,N_2734);
or U2938 (N_2938,N_2658,N_2620);
nor U2939 (N_2939,N_2658,N_2605);
and U2940 (N_2940,N_2730,N_2755);
or U2941 (N_2941,N_2694,N_2604);
nor U2942 (N_2942,N_2772,N_2653);
and U2943 (N_2943,N_2736,N_2752);
and U2944 (N_2944,N_2727,N_2747);
and U2945 (N_2945,N_2674,N_2768);
and U2946 (N_2946,N_2600,N_2787);
or U2947 (N_2947,N_2777,N_2700);
or U2948 (N_2948,N_2748,N_2636);
nand U2949 (N_2949,N_2744,N_2606);
nand U2950 (N_2950,N_2678,N_2703);
and U2951 (N_2951,N_2796,N_2655);
or U2952 (N_2952,N_2798,N_2732);
nor U2953 (N_2953,N_2600,N_2757);
nor U2954 (N_2954,N_2765,N_2711);
or U2955 (N_2955,N_2627,N_2660);
nor U2956 (N_2956,N_2700,N_2799);
and U2957 (N_2957,N_2774,N_2680);
xor U2958 (N_2958,N_2796,N_2798);
nor U2959 (N_2959,N_2734,N_2642);
nand U2960 (N_2960,N_2602,N_2784);
nand U2961 (N_2961,N_2779,N_2675);
nand U2962 (N_2962,N_2609,N_2640);
and U2963 (N_2963,N_2618,N_2749);
xor U2964 (N_2964,N_2778,N_2629);
nor U2965 (N_2965,N_2654,N_2681);
nand U2966 (N_2966,N_2657,N_2746);
nor U2967 (N_2967,N_2609,N_2797);
nand U2968 (N_2968,N_2610,N_2612);
nor U2969 (N_2969,N_2649,N_2785);
nand U2970 (N_2970,N_2771,N_2608);
or U2971 (N_2971,N_2768,N_2664);
nand U2972 (N_2972,N_2793,N_2752);
or U2973 (N_2973,N_2610,N_2777);
nor U2974 (N_2974,N_2776,N_2715);
nor U2975 (N_2975,N_2663,N_2617);
and U2976 (N_2976,N_2730,N_2622);
or U2977 (N_2977,N_2704,N_2602);
nand U2978 (N_2978,N_2777,N_2637);
nor U2979 (N_2979,N_2621,N_2797);
nand U2980 (N_2980,N_2675,N_2701);
nand U2981 (N_2981,N_2783,N_2748);
nor U2982 (N_2982,N_2717,N_2718);
nand U2983 (N_2983,N_2670,N_2688);
nor U2984 (N_2984,N_2603,N_2757);
nor U2985 (N_2985,N_2701,N_2609);
and U2986 (N_2986,N_2744,N_2694);
and U2987 (N_2987,N_2667,N_2605);
nor U2988 (N_2988,N_2759,N_2627);
nor U2989 (N_2989,N_2672,N_2625);
xor U2990 (N_2990,N_2704,N_2673);
or U2991 (N_2991,N_2784,N_2741);
and U2992 (N_2992,N_2798,N_2675);
and U2993 (N_2993,N_2791,N_2623);
or U2994 (N_2994,N_2734,N_2614);
nor U2995 (N_2995,N_2612,N_2626);
or U2996 (N_2996,N_2734,N_2718);
nor U2997 (N_2997,N_2733,N_2631);
or U2998 (N_2998,N_2632,N_2708);
nor U2999 (N_2999,N_2701,N_2688);
and UO_0 (O_0,N_2908,N_2807);
or UO_1 (O_1,N_2985,N_2830);
and UO_2 (O_2,N_2942,N_2883);
nand UO_3 (O_3,N_2916,N_2845);
or UO_4 (O_4,N_2804,N_2971);
nor UO_5 (O_5,N_2816,N_2988);
or UO_6 (O_6,N_2854,N_2912);
or UO_7 (O_7,N_2968,N_2800);
or UO_8 (O_8,N_2866,N_2842);
nand UO_9 (O_9,N_2928,N_2899);
or UO_10 (O_10,N_2833,N_2978);
nor UO_11 (O_11,N_2900,N_2917);
nor UO_12 (O_12,N_2951,N_2814);
nor UO_13 (O_13,N_2825,N_2998);
or UO_14 (O_14,N_2945,N_2984);
nand UO_15 (O_15,N_2808,N_2818);
or UO_16 (O_16,N_2875,N_2817);
xnor UO_17 (O_17,N_2958,N_2884);
or UO_18 (O_18,N_2893,N_2805);
or UO_19 (O_19,N_2931,N_2994);
xor UO_20 (O_20,N_2809,N_2961);
and UO_21 (O_21,N_2801,N_2839);
or UO_22 (O_22,N_2891,N_2925);
or UO_23 (O_23,N_2837,N_2901);
nand UO_24 (O_24,N_2956,N_2803);
or UO_25 (O_25,N_2834,N_2911);
and UO_26 (O_26,N_2841,N_2836);
nand UO_27 (O_27,N_2895,N_2936);
and UO_28 (O_28,N_2829,N_2976);
or UO_29 (O_29,N_2959,N_2941);
and UO_30 (O_30,N_2947,N_2950);
or UO_31 (O_31,N_2880,N_2877);
or UO_32 (O_32,N_2930,N_2828);
nor UO_33 (O_33,N_2843,N_2944);
nor UO_34 (O_34,N_2937,N_2896);
nor UO_35 (O_35,N_2894,N_2914);
nand UO_36 (O_36,N_2915,N_2962);
or UO_37 (O_37,N_2887,N_2977);
nor UO_38 (O_38,N_2850,N_2851);
nand UO_39 (O_39,N_2993,N_2873);
or UO_40 (O_40,N_2860,N_2870);
nor UO_41 (O_41,N_2822,N_2989);
nand UO_42 (O_42,N_2960,N_2810);
or UO_43 (O_43,N_2935,N_2859);
nand UO_44 (O_44,N_2926,N_2840);
or UO_45 (O_45,N_2923,N_2835);
xor UO_46 (O_46,N_2946,N_2980);
and UO_47 (O_47,N_2847,N_2878);
or UO_48 (O_48,N_2943,N_2806);
nand UO_49 (O_49,N_2927,N_2987);
nand UO_50 (O_50,N_2913,N_2813);
xnor UO_51 (O_51,N_2922,N_2802);
xnor UO_52 (O_52,N_2991,N_2972);
and UO_53 (O_53,N_2827,N_2905);
nand UO_54 (O_54,N_2932,N_2955);
and UO_55 (O_55,N_2846,N_2819);
and UO_56 (O_56,N_2876,N_2995);
and UO_57 (O_57,N_2957,N_2852);
nand UO_58 (O_58,N_2907,N_2832);
or UO_59 (O_59,N_2939,N_2865);
and UO_60 (O_60,N_2969,N_2924);
xnor UO_61 (O_61,N_2903,N_2869);
xnor UO_62 (O_62,N_2862,N_2996);
and UO_63 (O_63,N_2910,N_2871);
xor UO_64 (O_64,N_2898,N_2967);
and UO_65 (O_65,N_2983,N_2858);
or UO_66 (O_66,N_2921,N_2933);
or UO_67 (O_67,N_2815,N_2975);
xor UO_68 (O_68,N_2823,N_2929);
nor UO_69 (O_69,N_2879,N_2868);
nand UO_70 (O_70,N_2963,N_2909);
xor UO_71 (O_71,N_2953,N_2864);
or UO_72 (O_72,N_2890,N_2979);
and UO_73 (O_73,N_2853,N_2952);
xor UO_74 (O_74,N_2826,N_2999);
xor UO_75 (O_75,N_2821,N_2966);
and UO_76 (O_76,N_2918,N_2970);
and UO_77 (O_77,N_2888,N_2986);
and UO_78 (O_78,N_2934,N_2982);
nor UO_79 (O_79,N_2973,N_2990);
or UO_80 (O_80,N_2811,N_2863);
xnor UO_81 (O_81,N_2949,N_2881);
nand UO_82 (O_82,N_2992,N_2856);
nand UO_83 (O_83,N_2974,N_2954);
nand UO_84 (O_84,N_2981,N_2861);
and UO_85 (O_85,N_2964,N_2857);
or UO_86 (O_86,N_2897,N_2997);
nor UO_87 (O_87,N_2855,N_2920);
nor UO_88 (O_88,N_2867,N_2906);
and UO_89 (O_89,N_2882,N_2948);
nor UO_90 (O_90,N_2874,N_2820);
and UO_91 (O_91,N_2848,N_2824);
and UO_92 (O_92,N_2938,N_2904);
nor UO_93 (O_93,N_2831,N_2940);
nor UO_94 (O_94,N_2838,N_2885);
nand UO_95 (O_95,N_2889,N_2965);
nand UO_96 (O_96,N_2892,N_2919);
and UO_97 (O_97,N_2844,N_2812);
and UO_98 (O_98,N_2872,N_2886);
nor UO_99 (O_99,N_2902,N_2849);
nor UO_100 (O_100,N_2955,N_2864);
and UO_101 (O_101,N_2860,N_2851);
nand UO_102 (O_102,N_2938,N_2843);
and UO_103 (O_103,N_2957,N_2941);
xnor UO_104 (O_104,N_2806,N_2843);
nand UO_105 (O_105,N_2861,N_2979);
nand UO_106 (O_106,N_2927,N_2848);
nand UO_107 (O_107,N_2967,N_2956);
or UO_108 (O_108,N_2835,N_2819);
or UO_109 (O_109,N_2970,N_2982);
nand UO_110 (O_110,N_2961,N_2814);
or UO_111 (O_111,N_2979,N_2973);
nand UO_112 (O_112,N_2979,N_2995);
xor UO_113 (O_113,N_2932,N_2806);
nor UO_114 (O_114,N_2870,N_2813);
or UO_115 (O_115,N_2917,N_2808);
nand UO_116 (O_116,N_2851,N_2810);
nor UO_117 (O_117,N_2885,N_2990);
and UO_118 (O_118,N_2859,N_2974);
and UO_119 (O_119,N_2801,N_2822);
xnor UO_120 (O_120,N_2950,N_2920);
nand UO_121 (O_121,N_2893,N_2831);
nand UO_122 (O_122,N_2968,N_2964);
or UO_123 (O_123,N_2896,N_2863);
nor UO_124 (O_124,N_2903,N_2823);
and UO_125 (O_125,N_2825,N_2864);
or UO_126 (O_126,N_2970,N_2934);
and UO_127 (O_127,N_2888,N_2833);
and UO_128 (O_128,N_2819,N_2820);
and UO_129 (O_129,N_2932,N_2946);
nor UO_130 (O_130,N_2897,N_2965);
and UO_131 (O_131,N_2835,N_2824);
and UO_132 (O_132,N_2969,N_2816);
or UO_133 (O_133,N_2868,N_2890);
and UO_134 (O_134,N_2984,N_2850);
and UO_135 (O_135,N_2895,N_2839);
and UO_136 (O_136,N_2942,N_2980);
nand UO_137 (O_137,N_2932,N_2833);
nor UO_138 (O_138,N_2946,N_2931);
nor UO_139 (O_139,N_2872,N_2891);
nor UO_140 (O_140,N_2901,N_2904);
and UO_141 (O_141,N_2829,N_2943);
or UO_142 (O_142,N_2971,N_2938);
or UO_143 (O_143,N_2940,N_2932);
and UO_144 (O_144,N_2972,N_2820);
and UO_145 (O_145,N_2983,N_2958);
nand UO_146 (O_146,N_2973,N_2820);
nand UO_147 (O_147,N_2804,N_2976);
and UO_148 (O_148,N_2977,N_2922);
or UO_149 (O_149,N_2826,N_2970);
nand UO_150 (O_150,N_2920,N_2929);
nor UO_151 (O_151,N_2950,N_2808);
or UO_152 (O_152,N_2859,N_2889);
or UO_153 (O_153,N_2945,N_2888);
nor UO_154 (O_154,N_2835,N_2955);
nor UO_155 (O_155,N_2849,N_2847);
or UO_156 (O_156,N_2906,N_2942);
or UO_157 (O_157,N_2896,N_2956);
nand UO_158 (O_158,N_2804,N_2849);
and UO_159 (O_159,N_2890,N_2804);
and UO_160 (O_160,N_2944,N_2831);
xor UO_161 (O_161,N_2808,N_2988);
xnor UO_162 (O_162,N_2986,N_2863);
nor UO_163 (O_163,N_2883,N_2908);
or UO_164 (O_164,N_2929,N_2890);
nand UO_165 (O_165,N_2909,N_2823);
nor UO_166 (O_166,N_2873,N_2824);
or UO_167 (O_167,N_2969,N_2865);
nand UO_168 (O_168,N_2918,N_2996);
nor UO_169 (O_169,N_2939,N_2996);
nand UO_170 (O_170,N_2896,N_2932);
nor UO_171 (O_171,N_2886,N_2900);
nand UO_172 (O_172,N_2810,N_2811);
nand UO_173 (O_173,N_2989,N_2994);
or UO_174 (O_174,N_2802,N_2946);
nor UO_175 (O_175,N_2924,N_2963);
and UO_176 (O_176,N_2930,N_2877);
and UO_177 (O_177,N_2916,N_2810);
and UO_178 (O_178,N_2992,N_2820);
nand UO_179 (O_179,N_2931,N_2975);
nand UO_180 (O_180,N_2870,N_2920);
xnor UO_181 (O_181,N_2922,N_2856);
xor UO_182 (O_182,N_2988,N_2845);
nor UO_183 (O_183,N_2958,N_2878);
nand UO_184 (O_184,N_2979,N_2809);
and UO_185 (O_185,N_2884,N_2909);
or UO_186 (O_186,N_2871,N_2819);
or UO_187 (O_187,N_2829,N_2962);
and UO_188 (O_188,N_2829,N_2919);
or UO_189 (O_189,N_2989,N_2882);
and UO_190 (O_190,N_2843,N_2955);
nand UO_191 (O_191,N_2998,N_2919);
or UO_192 (O_192,N_2863,N_2912);
nor UO_193 (O_193,N_2986,N_2814);
nor UO_194 (O_194,N_2822,N_2889);
and UO_195 (O_195,N_2905,N_2970);
or UO_196 (O_196,N_2953,N_2888);
or UO_197 (O_197,N_2830,N_2844);
nor UO_198 (O_198,N_2947,N_2899);
and UO_199 (O_199,N_2856,N_2919);
xor UO_200 (O_200,N_2865,N_2909);
or UO_201 (O_201,N_2974,N_2819);
nor UO_202 (O_202,N_2830,N_2939);
or UO_203 (O_203,N_2808,N_2837);
or UO_204 (O_204,N_2845,N_2919);
and UO_205 (O_205,N_2917,N_2871);
nor UO_206 (O_206,N_2846,N_2830);
xnor UO_207 (O_207,N_2985,N_2860);
and UO_208 (O_208,N_2930,N_2842);
nor UO_209 (O_209,N_2804,N_2973);
or UO_210 (O_210,N_2826,N_2902);
or UO_211 (O_211,N_2959,N_2803);
and UO_212 (O_212,N_2947,N_2845);
nand UO_213 (O_213,N_2978,N_2923);
nor UO_214 (O_214,N_2911,N_2838);
nand UO_215 (O_215,N_2928,N_2842);
and UO_216 (O_216,N_2969,N_2809);
nor UO_217 (O_217,N_2908,N_2835);
xor UO_218 (O_218,N_2873,N_2901);
nand UO_219 (O_219,N_2968,N_2892);
and UO_220 (O_220,N_2859,N_2980);
or UO_221 (O_221,N_2897,N_2910);
or UO_222 (O_222,N_2841,N_2882);
xor UO_223 (O_223,N_2859,N_2951);
or UO_224 (O_224,N_2977,N_2907);
or UO_225 (O_225,N_2847,N_2988);
nand UO_226 (O_226,N_2976,N_2907);
nand UO_227 (O_227,N_2830,N_2973);
and UO_228 (O_228,N_2870,N_2940);
and UO_229 (O_229,N_2922,N_2861);
or UO_230 (O_230,N_2807,N_2909);
or UO_231 (O_231,N_2944,N_2812);
nor UO_232 (O_232,N_2949,N_2888);
or UO_233 (O_233,N_2883,N_2944);
nor UO_234 (O_234,N_2865,N_2908);
nor UO_235 (O_235,N_2978,N_2928);
nor UO_236 (O_236,N_2981,N_2870);
nor UO_237 (O_237,N_2991,N_2936);
nand UO_238 (O_238,N_2967,N_2935);
nand UO_239 (O_239,N_2876,N_2831);
and UO_240 (O_240,N_2868,N_2986);
nor UO_241 (O_241,N_2954,N_2955);
and UO_242 (O_242,N_2931,N_2932);
nand UO_243 (O_243,N_2992,N_2998);
and UO_244 (O_244,N_2921,N_2811);
or UO_245 (O_245,N_2981,N_2966);
nor UO_246 (O_246,N_2852,N_2813);
nor UO_247 (O_247,N_2882,N_2902);
and UO_248 (O_248,N_2847,N_2992);
and UO_249 (O_249,N_2810,N_2920);
nand UO_250 (O_250,N_2808,N_2921);
xnor UO_251 (O_251,N_2842,N_2867);
and UO_252 (O_252,N_2899,N_2875);
nand UO_253 (O_253,N_2980,N_2987);
or UO_254 (O_254,N_2971,N_2984);
or UO_255 (O_255,N_2802,N_2888);
nand UO_256 (O_256,N_2805,N_2862);
or UO_257 (O_257,N_2801,N_2813);
and UO_258 (O_258,N_2991,N_2995);
nor UO_259 (O_259,N_2992,N_2994);
nor UO_260 (O_260,N_2814,N_2909);
nand UO_261 (O_261,N_2858,N_2862);
nor UO_262 (O_262,N_2861,N_2966);
or UO_263 (O_263,N_2923,N_2872);
and UO_264 (O_264,N_2986,N_2939);
nor UO_265 (O_265,N_2811,N_2964);
nor UO_266 (O_266,N_2836,N_2933);
nand UO_267 (O_267,N_2988,N_2825);
nor UO_268 (O_268,N_2941,N_2810);
nand UO_269 (O_269,N_2862,N_2875);
xnor UO_270 (O_270,N_2810,N_2872);
nand UO_271 (O_271,N_2924,N_2911);
nand UO_272 (O_272,N_2800,N_2839);
and UO_273 (O_273,N_2861,N_2996);
and UO_274 (O_274,N_2997,N_2950);
nor UO_275 (O_275,N_2982,N_2879);
and UO_276 (O_276,N_2905,N_2985);
or UO_277 (O_277,N_2836,N_2839);
or UO_278 (O_278,N_2822,N_2955);
and UO_279 (O_279,N_2865,N_2837);
nor UO_280 (O_280,N_2922,N_2882);
xor UO_281 (O_281,N_2811,N_2878);
nand UO_282 (O_282,N_2844,N_2864);
or UO_283 (O_283,N_2817,N_2933);
and UO_284 (O_284,N_2993,N_2816);
nor UO_285 (O_285,N_2901,N_2866);
or UO_286 (O_286,N_2931,N_2809);
and UO_287 (O_287,N_2990,N_2850);
and UO_288 (O_288,N_2932,N_2924);
nand UO_289 (O_289,N_2932,N_2911);
and UO_290 (O_290,N_2963,N_2815);
nor UO_291 (O_291,N_2888,N_2910);
or UO_292 (O_292,N_2959,N_2835);
or UO_293 (O_293,N_2830,N_2891);
nand UO_294 (O_294,N_2981,N_2964);
nor UO_295 (O_295,N_2930,N_2889);
nand UO_296 (O_296,N_2890,N_2881);
or UO_297 (O_297,N_2998,N_2803);
nor UO_298 (O_298,N_2804,N_2826);
nor UO_299 (O_299,N_2811,N_2975);
nor UO_300 (O_300,N_2958,N_2907);
or UO_301 (O_301,N_2907,N_2975);
nand UO_302 (O_302,N_2970,N_2981);
or UO_303 (O_303,N_2951,N_2812);
and UO_304 (O_304,N_2879,N_2887);
or UO_305 (O_305,N_2899,N_2948);
and UO_306 (O_306,N_2981,N_2868);
or UO_307 (O_307,N_2993,N_2951);
or UO_308 (O_308,N_2861,N_2925);
xnor UO_309 (O_309,N_2816,N_2837);
nand UO_310 (O_310,N_2983,N_2874);
and UO_311 (O_311,N_2875,N_2888);
or UO_312 (O_312,N_2891,N_2847);
or UO_313 (O_313,N_2825,N_2960);
or UO_314 (O_314,N_2900,N_2983);
nor UO_315 (O_315,N_2834,N_2813);
nor UO_316 (O_316,N_2830,N_2822);
nand UO_317 (O_317,N_2879,N_2998);
xor UO_318 (O_318,N_2972,N_2982);
nand UO_319 (O_319,N_2959,N_2851);
nor UO_320 (O_320,N_2860,N_2801);
nor UO_321 (O_321,N_2994,N_2976);
and UO_322 (O_322,N_2800,N_2814);
and UO_323 (O_323,N_2932,N_2943);
nor UO_324 (O_324,N_2980,N_2808);
or UO_325 (O_325,N_2916,N_2901);
nor UO_326 (O_326,N_2986,N_2877);
or UO_327 (O_327,N_2838,N_2859);
or UO_328 (O_328,N_2992,N_2911);
or UO_329 (O_329,N_2861,N_2982);
nor UO_330 (O_330,N_2928,N_2871);
or UO_331 (O_331,N_2869,N_2945);
nand UO_332 (O_332,N_2841,N_2812);
or UO_333 (O_333,N_2996,N_2988);
xor UO_334 (O_334,N_2924,N_2915);
and UO_335 (O_335,N_2870,N_2895);
or UO_336 (O_336,N_2825,N_2994);
nor UO_337 (O_337,N_2850,N_2865);
xnor UO_338 (O_338,N_2987,N_2813);
nor UO_339 (O_339,N_2902,N_2993);
or UO_340 (O_340,N_2802,N_2996);
and UO_341 (O_341,N_2824,N_2938);
and UO_342 (O_342,N_2939,N_2814);
nor UO_343 (O_343,N_2950,N_2956);
and UO_344 (O_344,N_2858,N_2977);
or UO_345 (O_345,N_2869,N_2806);
nor UO_346 (O_346,N_2827,N_2860);
nor UO_347 (O_347,N_2985,N_2886);
nand UO_348 (O_348,N_2979,N_2899);
and UO_349 (O_349,N_2896,N_2856);
nand UO_350 (O_350,N_2953,N_2840);
and UO_351 (O_351,N_2800,N_2977);
nand UO_352 (O_352,N_2806,N_2968);
xor UO_353 (O_353,N_2918,N_2840);
or UO_354 (O_354,N_2852,N_2935);
nand UO_355 (O_355,N_2895,N_2808);
or UO_356 (O_356,N_2925,N_2818);
or UO_357 (O_357,N_2868,N_2958);
and UO_358 (O_358,N_2906,N_2802);
nor UO_359 (O_359,N_2833,N_2859);
and UO_360 (O_360,N_2801,N_2994);
and UO_361 (O_361,N_2824,N_2909);
or UO_362 (O_362,N_2903,N_2849);
or UO_363 (O_363,N_2913,N_2900);
or UO_364 (O_364,N_2834,N_2935);
nor UO_365 (O_365,N_2958,N_2912);
and UO_366 (O_366,N_2891,N_2908);
nand UO_367 (O_367,N_2880,N_2902);
or UO_368 (O_368,N_2866,N_2896);
nor UO_369 (O_369,N_2828,N_2971);
and UO_370 (O_370,N_2875,N_2969);
xor UO_371 (O_371,N_2885,N_2820);
nand UO_372 (O_372,N_2910,N_2885);
nor UO_373 (O_373,N_2980,N_2809);
nand UO_374 (O_374,N_2962,N_2891);
nor UO_375 (O_375,N_2980,N_2884);
or UO_376 (O_376,N_2879,N_2977);
xnor UO_377 (O_377,N_2913,N_2853);
and UO_378 (O_378,N_2963,N_2978);
and UO_379 (O_379,N_2896,N_2987);
and UO_380 (O_380,N_2977,N_2903);
nor UO_381 (O_381,N_2938,N_2841);
nand UO_382 (O_382,N_2904,N_2828);
nor UO_383 (O_383,N_2875,N_2962);
nor UO_384 (O_384,N_2911,N_2940);
or UO_385 (O_385,N_2984,N_2882);
nor UO_386 (O_386,N_2966,N_2877);
xor UO_387 (O_387,N_2928,N_2800);
nor UO_388 (O_388,N_2872,N_2867);
nand UO_389 (O_389,N_2967,N_2970);
and UO_390 (O_390,N_2964,N_2893);
and UO_391 (O_391,N_2822,N_2995);
and UO_392 (O_392,N_2854,N_2839);
xor UO_393 (O_393,N_2995,N_2923);
or UO_394 (O_394,N_2953,N_2962);
nor UO_395 (O_395,N_2966,N_2897);
nand UO_396 (O_396,N_2964,N_2835);
and UO_397 (O_397,N_2840,N_2819);
or UO_398 (O_398,N_2806,N_2865);
or UO_399 (O_399,N_2808,N_2884);
and UO_400 (O_400,N_2997,N_2866);
or UO_401 (O_401,N_2990,N_2883);
xor UO_402 (O_402,N_2840,N_2830);
and UO_403 (O_403,N_2854,N_2978);
nand UO_404 (O_404,N_2947,N_2978);
or UO_405 (O_405,N_2863,N_2989);
nor UO_406 (O_406,N_2968,N_2979);
nand UO_407 (O_407,N_2810,N_2959);
and UO_408 (O_408,N_2812,N_2930);
nand UO_409 (O_409,N_2984,N_2905);
nor UO_410 (O_410,N_2875,N_2820);
or UO_411 (O_411,N_2865,N_2925);
or UO_412 (O_412,N_2896,N_2963);
and UO_413 (O_413,N_2900,N_2999);
nand UO_414 (O_414,N_2982,N_2974);
nand UO_415 (O_415,N_2899,N_2931);
nor UO_416 (O_416,N_2920,N_2911);
xor UO_417 (O_417,N_2823,N_2819);
and UO_418 (O_418,N_2944,N_2963);
or UO_419 (O_419,N_2946,N_2825);
nor UO_420 (O_420,N_2970,N_2957);
and UO_421 (O_421,N_2911,N_2927);
nor UO_422 (O_422,N_2987,N_2810);
and UO_423 (O_423,N_2980,N_2913);
nor UO_424 (O_424,N_2859,N_2943);
or UO_425 (O_425,N_2941,N_2943);
nor UO_426 (O_426,N_2836,N_2885);
nor UO_427 (O_427,N_2972,N_2981);
xor UO_428 (O_428,N_2885,N_2991);
and UO_429 (O_429,N_2972,N_2994);
or UO_430 (O_430,N_2873,N_2883);
or UO_431 (O_431,N_2811,N_2950);
or UO_432 (O_432,N_2907,N_2843);
nand UO_433 (O_433,N_2863,N_2868);
and UO_434 (O_434,N_2889,N_2951);
nand UO_435 (O_435,N_2864,N_2920);
nor UO_436 (O_436,N_2932,N_2820);
xor UO_437 (O_437,N_2932,N_2814);
or UO_438 (O_438,N_2884,N_2801);
and UO_439 (O_439,N_2862,N_2933);
nor UO_440 (O_440,N_2999,N_2830);
xor UO_441 (O_441,N_2845,N_2888);
or UO_442 (O_442,N_2987,N_2831);
nand UO_443 (O_443,N_2915,N_2828);
nor UO_444 (O_444,N_2870,N_2823);
or UO_445 (O_445,N_2822,N_2846);
nor UO_446 (O_446,N_2933,N_2945);
or UO_447 (O_447,N_2991,N_2887);
or UO_448 (O_448,N_2810,N_2977);
or UO_449 (O_449,N_2818,N_2989);
nor UO_450 (O_450,N_2913,N_2862);
nor UO_451 (O_451,N_2907,N_2867);
and UO_452 (O_452,N_2853,N_2944);
and UO_453 (O_453,N_2841,N_2969);
or UO_454 (O_454,N_2864,N_2872);
xnor UO_455 (O_455,N_2916,N_2831);
or UO_456 (O_456,N_2883,N_2938);
and UO_457 (O_457,N_2885,N_2933);
nand UO_458 (O_458,N_2843,N_2845);
and UO_459 (O_459,N_2937,N_2906);
nor UO_460 (O_460,N_2843,N_2887);
nand UO_461 (O_461,N_2837,N_2929);
or UO_462 (O_462,N_2803,N_2975);
or UO_463 (O_463,N_2825,N_2891);
nor UO_464 (O_464,N_2953,N_2964);
nor UO_465 (O_465,N_2898,N_2938);
nor UO_466 (O_466,N_2887,N_2964);
and UO_467 (O_467,N_2955,N_2974);
nand UO_468 (O_468,N_2867,N_2891);
nor UO_469 (O_469,N_2906,N_2966);
xnor UO_470 (O_470,N_2869,N_2970);
nand UO_471 (O_471,N_2988,N_2906);
or UO_472 (O_472,N_2951,N_2978);
or UO_473 (O_473,N_2860,N_2874);
and UO_474 (O_474,N_2870,N_2807);
nor UO_475 (O_475,N_2949,N_2928);
nand UO_476 (O_476,N_2923,N_2819);
nand UO_477 (O_477,N_2924,N_2998);
and UO_478 (O_478,N_2908,N_2884);
nor UO_479 (O_479,N_2860,N_2850);
and UO_480 (O_480,N_2853,N_2937);
or UO_481 (O_481,N_2847,N_2932);
nor UO_482 (O_482,N_2938,N_2818);
and UO_483 (O_483,N_2904,N_2979);
nand UO_484 (O_484,N_2827,N_2954);
and UO_485 (O_485,N_2897,N_2826);
or UO_486 (O_486,N_2974,N_2948);
nand UO_487 (O_487,N_2926,N_2864);
or UO_488 (O_488,N_2859,N_2805);
or UO_489 (O_489,N_2878,N_2955);
and UO_490 (O_490,N_2904,N_2881);
nor UO_491 (O_491,N_2928,N_2922);
and UO_492 (O_492,N_2867,N_2965);
xnor UO_493 (O_493,N_2942,N_2981);
nand UO_494 (O_494,N_2893,N_2941);
xnor UO_495 (O_495,N_2989,N_2936);
nor UO_496 (O_496,N_2886,N_2881);
nor UO_497 (O_497,N_2864,N_2886);
nor UO_498 (O_498,N_2880,N_2961);
and UO_499 (O_499,N_2886,N_2997);
endmodule